
module auction_BMR_N7_W32 ( p_input, o );
  input [4095:0] p_input;
  output [38:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408;

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(o[6]), .B(n3), .Z(n1) );
  XOR U3 ( .A(n2), .B(n4), .Z(n3) );
  XOR U4 ( .A(n5), .B(n6), .Z(o[8]) );
  AND U5 ( .A(o[6]), .B(n7), .Z(n5) );
  XOR U6 ( .A(n8), .B(n9), .Z(n7) );
  XNOR U7 ( .A(n10), .B(n11), .Z(o[7]) );
  AND U8 ( .A(o[6]), .B(n12), .Z(n10) );
  XNOR U9 ( .A(n13), .B(n11), .Z(n12) );
  XOR U10 ( .A(n14), .B(n15), .Z(o[38]) );
  AND U11 ( .A(o[6]), .B(n16), .Z(n14) );
  XOR U12 ( .A(n17), .B(n18), .Z(n16) );
  XOR U13 ( .A(n19), .B(n20), .Z(o[37]) );
  AND U14 ( .A(o[6]), .B(n21), .Z(n19) );
  XOR U15 ( .A(n22), .B(n23), .Z(n21) );
  XOR U16 ( .A(n24), .B(n25), .Z(o[36]) );
  AND U17 ( .A(o[6]), .B(n26), .Z(n24) );
  XOR U18 ( .A(n27), .B(n28), .Z(n26) );
  XOR U19 ( .A(n29), .B(n30), .Z(o[35]) );
  AND U20 ( .A(o[6]), .B(n31), .Z(n29) );
  XOR U21 ( .A(n32), .B(n33), .Z(n31) );
  XOR U22 ( .A(n34), .B(n35), .Z(o[34]) );
  AND U23 ( .A(o[6]), .B(n36), .Z(n34) );
  XOR U24 ( .A(n37), .B(n38), .Z(n36) );
  XOR U25 ( .A(n39), .B(n40), .Z(o[33]) );
  AND U26 ( .A(o[6]), .B(n41), .Z(n39) );
  XOR U27 ( .A(n42), .B(n43), .Z(n41) );
  XOR U28 ( .A(n44), .B(n45), .Z(o[32]) );
  AND U29 ( .A(o[6]), .B(n46), .Z(n44) );
  XOR U30 ( .A(n47), .B(n48), .Z(n46) );
  XOR U31 ( .A(n49), .B(n50), .Z(o[31]) );
  AND U32 ( .A(o[6]), .B(n51), .Z(n49) );
  XOR U33 ( .A(n52), .B(n53), .Z(n51) );
  XOR U34 ( .A(n54), .B(n55), .Z(o[30]) );
  AND U35 ( .A(o[6]), .B(n56), .Z(n54) );
  XOR U36 ( .A(n57), .B(n58), .Z(n56) );
  XOR U37 ( .A(n59), .B(n60), .Z(o[29]) );
  AND U38 ( .A(o[6]), .B(n61), .Z(n59) );
  XOR U39 ( .A(n62), .B(n63), .Z(n61) );
  XOR U40 ( .A(n64), .B(n65), .Z(o[28]) );
  AND U41 ( .A(o[6]), .B(n66), .Z(n64) );
  XOR U42 ( .A(n67), .B(n68), .Z(n66) );
  XOR U43 ( .A(n69), .B(n70), .Z(o[27]) );
  AND U44 ( .A(o[6]), .B(n71), .Z(n69) );
  XOR U45 ( .A(n72), .B(n73), .Z(n71) );
  XOR U46 ( .A(n74), .B(n75), .Z(o[26]) );
  AND U47 ( .A(o[6]), .B(n76), .Z(n74) );
  XOR U48 ( .A(n77), .B(n78), .Z(n76) );
  XOR U49 ( .A(n79), .B(n80), .Z(o[25]) );
  AND U50 ( .A(o[6]), .B(n81), .Z(n79) );
  XOR U51 ( .A(n82), .B(n83), .Z(n81) );
  XOR U52 ( .A(n84), .B(n85), .Z(o[24]) );
  AND U53 ( .A(o[6]), .B(n86), .Z(n84) );
  XOR U54 ( .A(n87), .B(n88), .Z(n86) );
  XOR U55 ( .A(n89), .B(n90), .Z(o[23]) );
  AND U56 ( .A(o[6]), .B(n91), .Z(n89) );
  XOR U57 ( .A(n92), .B(n93), .Z(n91) );
  XOR U58 ( .A(n94), .B(n95), .Z(o[22]) );
  AND U59 ( .A(o[6]), .B(n96), .Z(n94) );
  XOR U60 ( .A(n97), .B(n98), .Z(n96) );
  XOR U61 ( .A(n99), .B(n100), .Z(o[21]) );
  AND U62 ( .A(o[6]), .B(n101), .Z(n99) );
  XOR U63 ( .A(n102), .B(n103), .Z(n101) );
  XOR U64 ( .A(n104), .B(n105), .Z(o[20]) );
  AND U65 ( .A(o[6]), .B(n106), .Z(n104) );
  XOR U66 ( .A(n107), .B(n108), .Z(n106) );
  XOR U67 ( .A(n109), .B(n110), .Z(o[19]) );
  AND U68 ( .A(o[6]), .B(n111), .Z(n109) );
  XOR U69 ( .A(n112), .B(n113), .Z(n111) );
  XOR U70 ( .A(n114), .B(n115), .Z(o[18]) );
  AND U71 ( .A(o[6]), .B(n116), .Z(n114) );
  XOR U72 ( .A(n117), .B(n118), .Z(n116) );
  XOR U73 ( .A(n119), .B(n120), .Z(o[17]) );
  AND U74 ( .A(o[6]), .B(n121), .Z(n119) );
  XOR U75 ( .A(n122), .B(n123), .Z(n121) );
  XOR U76 ( .A(n124), .B(n125), .Z(o[16]) );
  AND U77 ( .A(o[6]), .B(n126), .Z(n124) );
  XOR U78 ( .A(n127), .B(n128), .Z(n126) );
  XOR U79 ( .A(n129), .B(n130), .Z(o[15]) );
  AND U80 ( .A(o[6]), .B(n131), .Z(n129) );
  XOR U81 ( .A(n132), .B(n133), .Z(n131) );
  XOR U82 ( .A(n134), .B(n135), .Z(o[14]) );
  AND U83 ( .A(o[6]), .B(n136), .Z(n134) );
  XOR U84 ( .A(n137), .B(n138), .Z(n136) );
  XOR U85 ( .A(n139), .B(n140), .Z(o[13]) );
  AND U86 ( .A(o[6]), .B(n141), .Z(n139) );
  XOR U87 ( .A(n142), .B(n143), .Z(n141) );
  XOR U88 ( .A(n144), .B(n145), .Z(o[12]) );
  AND U89 ( .A(o[6]), .B(n146), .Z(n144) );
  XOR U90 ( .A(n147), .B(n148), .Z(n146) );
  XOR U91 ( .A(n149), .B(n150), .Z(o[11]) );
  AND U92 ( .A(o[6]), .B(n151), .Z(n149) );
  XOR U93 ( .A(n152), .B(n153), .Z(n151) );
  XOR U94 ( .A(n154), .B(n155), .Z(o[10]) );
  AND U95 ( .A(o[6]), .B(n156), .Z(n154) );
  XOR U96 ( .A(n157), .B(n158), .Z(n156) );
  XOR U97 ( .A(n159), .B(n160), .Z(o[0]) );
  AND U98 ( .A(o[1]), .B(n161), .Z(n160) );
  XNOR U99 ( .A(n162), .B(n163), .Z(n161) );
  XNOR U100 ( .A(n164), .B(n159), .Z(n163) );
  AND U101 ( .A(o[2]), .B(n165), .Z(n164) );
  XNOR U102 ( .A(n166), .B(n167), .Z(n165) );
  XNOR U103 ( .A(n168), .B(n162), .Z(n167) );
  AND U104 ( .A(o[3]), .B(n169), .Z(n168) );
  XNOR U105 ( .A(n170), .B(n171), .Z(n169) );
  XNOR U106 ( .A(n172), .B(n166), .Z(n171) );
  AND U107 ( .A(o[4]), .B(n173), .Z(n172) );
  XNOR U108 ( .A(n174), .B(n175), .Z(n173) );
  XNOR U109 ( .A(n176), .B(n170), .Z(n175) );
  AND U110 ( .A(o[5]), .B(n177), .Z(n176) );
  XNOR U111 ( .A(n174), .B(n178), .Z(n177) );
  XNOR U112 ( .A(n179), .B(n180), .Z(n178) );
  AND U113 ( .A(o[6]), .B(n181), .Z(n179) );
  XOR U114 ( .A(n180), .B(n182), .Z(n181) );
  XOR U115 ( .A(n183), .B(n184), .Z(n174) );
  AND U116 ( .A(o[6]), .B(n185), .Z(n184) );
  XOR U117 ( .A(n183), .B(n186), .Z(n185) );
  XOR U118 ( .A(n187), .B(n188), .Z(n170) );
  AND U119 ( .A(o[5]), .B(n189), .Z(n188) );
  XNOR U120 ( .A(n187), .B(n190), .Z(n189) );
  XNOR U121 ( .A(n191), .B(n192), .Z(n190) );
  AND U122 ( .A(o[6]), .B(n193), .Z(n191) );
  XOR U123 ( .A(n192), .B(n194), .Z(n193) );
  XOR U124 ( .A(n195), .B(n196), .Z(n187) );
  AND U125 ( .A(o[6]), .B(n197), .Z(n196) );
  XOR U126 ( .A(n195), .B(n198), .Z(n197) );
  XOR U127 ( .A(n199), .B(n200), .Z(n166) );
  AND U128 ( .A(o[4]), .B(n201), .Z(n200) );
  XNOR U129 ( .A(n202), .B(n203), .Z(n201) );
  XNOR U130 ( .A(n204), .B(n199), .Z(n203) );
  AND U131 ( .A(o[5]), .B(n205), .Z(n204) );
  XNOR U132 ( .A(n202), .B(n206), .Z(n205) );
  XNOR U133 ( .A(n207), .B(n208), .Z(n206) );
  AND U134 ( .A(o[6]), .B(n209), .Z(n207) );
  XOR U135 ( .A(n208), .B(n210), .Z(n209) );
  XOR U136 ( .A(n211), .B(n212), .Z(n202) );
  AND U137 ( .A(o[6]), .B(n213), .Z(n212) );
  XOR U138 ( .A(n211), .B(n214), .Z(n213) );
  XOR U139 ( .A(n215), .B(n216), .Z(n199) );
  AND U140 ( .A(o[5]), .B(n217), .Z(n216) );
  XNOR U141 ( .A(n215), .B(n218), .Z(n217) );
  XNOR U142 ( .A(n219), .B(n220), .Z(n218) );
  AND U143 ( .A(o[6]), .B(n221), .Z(n219) );
  XOR U144 ( .A(n220), .B(n222), .Z(n221) );
  XOR U145 ( .A(n223), .B(n224), .Z(n215) );
  AND U146 ( .A(o[6]), .B(n225), .Z(n224) );
  XOR U147 ( .A(n223), .B(n226), .Z(n225) );
  XOR U148 ( .A(n227), .B(n228), .Z(n162) );
  AND U149 ( .A(o[3]), .B(n229), .Z(n228) );
  XNOR U150 ( .A(n230), .B(n231), .Z(n229) );
  XNOR U151 ( .A(n232), .B(n227), .Z(n231) );
  AND U152 ( .A(o[4]), .B(n233), .Z(n232) );
  XNOR U153 ( .A(n234), .B(n235), .Z(n233) );
  XNOR U154 ( .A(n236), .B(n230), .Z(n235) );
  AND U155 ( .A(o[5]), .B(n237), .Z(n236) );
  XNOR U156 ( .A(n234), .B(n238), .Z(n237) );
  XNOR U157 ( .A(n239), .B(n240), .Z(n238) );
  AND U158 ( .A(o[6]), .B(n241), .Z(n239) );
  XOR U159 ( .A(n240), .B(n242), .Z(n241) );
  XOR U160 ( .A(n243), .B(n244), .Z(n234) );
  AND U161 ( .A(o[6]), .B(n245), .Z(n244) );
  XOR U162 ( .A(n243), .B(n246), .Z(n245) );
  XOR U163 ( .A(n247), .B(n248), .Z(n230) );
  AND U164 ( .A(o[5]), .B(n249), .Z(n248) );
  XNOR U165 ( .A(n247), .B(n250), .Z(n249) );
  XNOR U166 ( .A(n251), .B(n252), .Z(n250) );
  AND U167 ( .A(o[6]), .B(n253), .Z(n251) );
  XOR U168 ( .A(n252), .B(n254), .Z(n253) );
  XOR U169 ( .A(n255), .B(n256), .Z(n247) );
  AND U170 ( .A(o[6]), .B(n257), .Z(n256) );
  XOR U171 ( .A(n255), .B(n258), .Z(n257) );
  XOR U172 ( .A(n259), .B(n260), .Z(n227) );
  AND U173 ( .A(o[4]), .B(n261), .Z(n260) );
  XNOR U174 ( .A(n262), .B(n263), .Z(n261) );
  XNOR U175 ( .A(n264), .B(n259), .Z(n263) );
  AND U176 ( .A(o[5]), .B(n265), .Z(n264) );
  XNOR U177 ( .A(n262), .B(n266), .Z(n265) );
  XNOR U178 ( .A(n267), .B(n268), .Z(n266) );
  AND U179 ( .A(o[6]), .B(n269), .Z(n267) );
  XOR U180 ( .A(n268), .B(n270), .Z(n269) );
  XOR U181 ( .A(n271), .B(n272), .Z(n262) );
  AND U182 ( .A(o[6]), .B(n273), .Z(n272) );
  XOR U183 ( .A(n271), .B(n274), .Z(n273) );
  XOR U184 ( .A(n275), .B(n276), .Z(n259) );
  AND U185 ( .A(o[5]), .B(n277), .Z(n276) );
  XNOR U186 ( .A(n275), .B(n278), .Z(n277) );
  XNOR U187 ( .A(n279), .B(n280), .Z(n278) );
  AND U188 ( .A(o[6]), .B(n281), .Z(n279) );
  XOR U189 ( .A(n280), .B(n282), .Z(n281) );
  XOR U190 ( .A(n283), .B(n284), .Z(n275) );
  AND U191 ( .A(o[6]), .B(n285), .Z(n284) );
  XOR U192 ( .A(n283), .B(n286), .Z(n285) );
  XOR U193 ( .A(n287), .B(n288), .Z(o[1]) );
  AND U194 ( .A(o[2]), .B(n289), .Z(n288) );
  XNOR U195 ( .A(n290), .B(n291), .Z(n289) );
  XNOR U196 ( .A(n292), .B(n287), .Z(n291) );
  AND U197 ( .A(o[3]), .B(n293), .Z(n292) );
  XNOR U198 ( .A(n294), .B(n295), .Z(n293) );
  XNOR U199 ( .A(n296), .B(n290), .Z(n295) );
  AND U200 ( .A(o[4]), .B(n297), .Z(n296) );
  XNOR U201 ( .A(n298), .B(n299), .Z(n297) );
  XNOR U202 ( .A(n300), .B(n294), .Z(n299) );
  AND U203 ( .A(o[5]), .B(n301), .Z(n300) );
  XNOR U204 ( .A(n298), .B(n302), .Z(n301) );
  XNOR U205 ( .A(n303), .B(n304), .Z(n302) );
  AND U206 ( .A(o[6]), .B(n305), .Z(n303) );
  XOR U207 ( .A(n304), .B(n306), .Z(n305) );
  XOR U208 ( .A(n307), .B(n308), .Z(n298) );
  AND U209 ( .A(o[6]), .B(n309), .Z(n308) );
  XOR U210 ( .A(n307), .B(n310), .Z(n309) );
  XOR U211 ( .A(n311), .B(n312), .Z(n294) );
  AND U212 ( .A(o[5]), .B(n313), .Z(n312) );
  XNOR U213 ( .A(n311), .B(n314), .Z(n313) );
  XNOR U214 ( .A(n315), .B(n316), .Z(n314) );
  AND U215 ( .A(o[6]), .B(n317), .Z(n315) );
  XOR U216 ( .A(n316), .B(n318), .Z(n317) );
  XOR U217 ( .A(n319), .B(n320), .Z(n311) );
  AND U218 ( .A(o[6]), .B(n321), .Z(n320) );
  XOR U219 ( .A(n319), .B(n322), .Z(n321) );
  XOR U220 ( .A(n323), .B(n324), .Z(n290) );
  AND U221 ( .A(o[4]), .B(n325), .Z(n324) );
  XNOR U222 ( .A(n326), .B(n327), .Z(n325) );
  XNOR U223 ( .A(n328), .B(n323), .Z(n327) );
  AND U224 ( .A(o[5]), .B(n329), .Z(n328) );
  XNOR U225 ( .A(n326), .B(n330), .Z(n329) );
  XNOR U226 ( .A(n331), .B(n332), .Z(n330) );
  AND U227 ( .A(o[6]), .B(n333), .Z(n331) );
  XOR U228 ( .A(n332), .B(n334), .Z(n333) );
  XOR U229 ( .A(n335), .B(n336), .Z(n326) );
  AND U230 ( .A(o[6]), .B(n337), .Z(n336) );
  XOR U231 ( .A(n335), .B(n338), .Z(n337) );
  XOR U232 ( .A(n339), .B(n340), .Z(n323) );
  AND U233 ( .A(o[5]), .B(n341), .Z(n340) );
  XNOR U234 ( .A(n339), .B(n342), .Z(n341) );
  XNOR U235 ( .A(n343), .B(n344), .Z(n342) );
  AND U236 ( .A(o[6]), .B(n345), .Z(n343) );
  XOR U237 ( .A(n344), .B(n346), .Z(n345) );
  XOR U238 ( .A(n347), .B(n348), .Z(n339) );
  AND U239 ( .A(o[6]), .B(n349), .Z(n348) );
  XOR U240 ( .A(n347), .B(n350), .Z(n349) );
  XOR U241 ( .A(n351), .B(n352), .Z(n287) );
  AND U242 ( .A(o[3]), .B(n353), .Z(n352) );
  XNOR U243 ( .A(n354), .B(n355), .Z(n353) );
  XNOR U244 ( .A(n356), .B(n351), .Z(n355) );
  AND U245 ( .A(o[4]), .B(n357), .Z(n356) );
  XNOR U246 ( .A(n358), .B(n359), .Z(n357) );
  XNOR U247 ( .A(n360), .B(n354), .Z(n359) );
  AND U248 ( .A(o[5]), .B(n361), .Z(n360) );
  XNOR U249 ( .A(n358), .B(n362), .Z(n361) );
  XNOR U250 ( .A(n363), .B(n364), .Z(n362) );
  AND U251 ( .A(o[6]), .B(n365), .Z(n363) );
  XOR U252 ( .A(n364), .B(n366), .Z(n365) );
  XOR U253 ( .A(n367), .B(n368), .Z(n358) );
  AND U254 ( .A(o[6]), .B(n369), .Z(n368) );
  XOR U255 ( .A(n367), .B(n370), .Z(n369) );
  XOR U256 ( .A(n371), .B(n372), .Z(n354) );
  AND U257 ( .A(o[5]), .B(n373), .Z(n372) );
  XNOR U258 ( .A(n371), .B(n374), .Z(n373) );
  XNOR U259 ( .A(n375), .B(n376), .Z(n374) );
  AND U260 ( .A(o[6]), .B(n377), .Z(n375) );
  XOR U261 ( .A(n376), .B(n378), .Z(n377) );
  XOR U262 ( .A(n379), .B(n380), .Z(n371) );
  AND U263 ( .A(o[6]), .B(n381), .Z(n380) );
  XOR U264 ( .A(n379), .B(n382), .Z(n381) );
  XOR U265 ( .A(n383), .B(n384), .Z(n351) );
  AND U266 ( .A(o[4]), .B(n385), .Z(n384) );
  XNOR U267 ( .A(n386), .B(n387), .Z(n385) );
  XNOR U268 ( .A(n388), .B(n383), .Z(n387) );
  AND U269 ( .A(o[5]), .B(n389), .Z(n388) );
  XNOR U270 ( .A(n386), .B(n390), .Z(n389) );
  XNOR U271 ( .A(n391), .B(n392), .Z(n390) );
  AND U272 ( .A(o[6]), .B(n393), .Z(n391) );
  XOR U273 ( .A(n392), .B(n394), .Z(n393) );
  XOR U274 ( .A(n395), .B(n396), .Z(n386) );
  AND U275 ( .A(o[6]), .B(n397), .Z(n396) );
  XOR U276 ( .A(n395), .B(n398), .Z(n397) );
  XOR U277 ( .A(n399), .B(n400), .Z(n383) );
  AND U278 ( .A(o[5]), .B(n401), .Z(n400) );
  XNOR U279 ( .A(n399), .B(n402), .Z(n401) );
  XNOR U280 ( .A(n403), .B(n404), .Z(n402) );
  AND U281 ( .A(o[6]), .B(n405), .Z(n403) );
  XOR U282 ( .A(n404), .B(n406), .Z(n405) );
  XOR U283 ( .A(n407), .B(n408), .Z(n399) );
  AND U284 ( .A(o[6]), .B(n409), .Z(n408) );
  XOR U285 ( .A(n407), .B(n410), .Z(n409) );
  XOR U286 ( .A(n411), .B(n412), .Z(n159) );
  AND U287 ( .A(o[2]), .B(n413), .Z(n412) );
  XNOR U288 ( .A(n414), .B(n415), .Z(n413) );
  XNOR U289 ( .A(n416), .B(n411), .Z(n415) );
  AND U290 ( .A(o[3]), .B(n417), .Z(n416) );
  XNOR U291 ( .A(n418), .B(n419), .Z(n417) );
  XNOR U292 ( .A(n420), .B(n414), .Z(n419) );
  AND U293 ( .A(o[4]), .B(n421), .Z(n420) );
  XNOR U294 ( .A(n422), .B(n423), .Z(n421) );
  XNOR U295 ( .A(n424), .B(n418), .Z(n423) );
  AND U296 ( .A(o[5]), .B(n425), .Z(n424) );
  XNOR U297 ( .A(n422), .B(n426), .Z(n425) );
  XNOR U298 ( .A(n427), .B(n428), .Z(n426) );
  AND U299 ( .A(o[6]), .B(n429), .Z(n427) );
  XOR U300 ( .A(n428), .B(n430), .Z(n429) );
  XOR U301 ( .A(n431), .B(n432), .Z(n422) );
  AND U302 ( .A(o[6]), .B(n433), .Z(n432) );
  XOR U303 ( .A(n431), .B(n434), .Z(n433) );
  XOR U304 ( .A(n435), .B(n436), .Z(n418) );
  AND U305 ( .A(o[5]), .B(n437), .Z(n436) );
  XNOR U306 ( .A(n435), .B(n438), .Z(n437) );
  XNOR U307 ( .A(n439), .B(n440), .Z(n438) );
  AND U308 ( .A(o[6]), .B(n441), .Z(n439) );
  XOR U309 ( .A(n440), .B(n442), .Z(n441) );
  XOR U310 ( .A(n443), .B(n444), .Z(n435) );
  AND U311 ( .A(o[6]), .B(n445), .Z(n444) );
  XOR U312 ( .A(n443), .B(n446), .Z(n445) );
  XOR U313 ( .A(n447), .B(n448), .Z(n414) );
  AND U314 ( .A(o[4]), .B(n449), .Z(n448) );
  XNOR U315 ( .A(n450), .B(n451), .Z(n449) );
  XNOR U316 ( .A(n452), .B(n447), .Z(n451) );
  AND U317 ( .A(o[5]), .B(n453), .Z(n452) );
  XNOR U318 ( .A(n450), .B(n454), .Z(n453) );
  XNOR U319 ( .A(n455), .B(n456), .Z(n454) );
  AND U320 ( .A(o[6]), .B(n457), .Z(n455) );
  XOR U321 ( .A(n456), .B(n458), .Z(n457) );
  XOR U322 ( .A(n459), .B(n460), .Z(n450) );
  AND U323 ( .A(o[6]), .B(n461), .Z(n460) );
  XOR U324 ( .A(n459), .B(n462), .Z(n461) );
  XOR U325 ( .A(n463), .B(n464), .Z(n447) );
  AND U326 ( .A(o[5]), .B(n465), .Z(n464) );
  XNOR U327 ( .A(n463), .B(n466), .Z(n465) );
  XNOR U328 ( .A(n467), .B(n468), .Z(n466) );
  AND U329 ( .A(o[6]), .B(n469), .Z(n467) );
  XOR U330 ( .A(n468), .B(n470), .Z(n469) );
  XOR U331 ( .A(n471), .B(n472), .Z(n463) );
  AND U332 ( .A(o[6]), .B(n473), .Z(n472) );
  XOR U333 ( .A(n471), .B(n474), .Z(n473) );
  XOR U334 ( .A(n475), .B(n476), .Z(o[2]) );
  AND U335 ( .A(o[3]), .B(n477), .Z(n476) );
  XNOR U336 ( .A(n478), .B(n479), .Z(n477) );
  XNOR U337 ( .A(n480), .B(n475), .Z(n479) );
  AND U338 ( .A(o[4]), .B(n481), .Z(n480) );
  XNOR U339 ( .A(n482), .B(n483), .Z(n481) );
  XNOR U340 ( .A(n484), .B(n478), .Z(n483) );
  AND U341 ( .A(o[5]), .B(n485), .Z(n484) );
  XNOR U342 ( .A(n482), .B(n486), .Z(n485) );
  XNOR U343 ( .A(n487), .B(n488), .Z(n486) );
  AND U344 ( .A(o[6]), .B(n489), .Z(n487) );
  XOR U345 ( .A(n488), .B(n490), .Z(n489) );
  XOR U346 ( .A(n491), .B(n492), .Z(n482) );
  AND U347 ( .A(o[6]), .B(n493), .Z(n492) );
  XOR U348 ( .A(n491), .B(n494), .Z(n493) );
  XOR U349 ( .A(n495), .B(n496), .Z(n478) );
  AND U350 ( .A(o[5]), .B(n497), .Z(n496) );
  XNOR U351 ( .A(n495), .B(n498), .Z(n497) );
  XNOR U352 ( .A(n499), .B(n500), .Z(n498) );
  AND U353 ( .A(o[6]), .B(n501), .Z(n499) );
  XOR U354 ( .A(n500), .B(n502), .Z(n501) );
  XOR U355 ( .A(n503), .B(n504), .Z(n495) );
  AND U356 ( .A(o[6]), .B(n505), .Z(n504) );
  XOR U357 ( .A(n503), .B(n506), .Z(n505) );
  XOR U358 ( .A(n507), .B(n508), .Z(n475) );
  AND U359 ( .A(o[4]), .B(n509), .Z(n508) );
  XNOR U360 ( .A(n510), .B(n511), .Z(n509) );
  XNOR U361 ( .A(n512), .B(n507), .Z(n511) );
  AND U362 ( .A(o[5]), .B(n513), .Z(n512) );
  XNOR U363 ( .A(n510), .B(n514), .Z(n513) );
  XNOR U364 ( .A(n515), .B(n516), .Z(n514) );
  AND U365 ( .A(o[6]), .B(n517), .Z(n515) );
  XOR U366 ( .A(n516), .B(n518), .Z(n517) );
  XOR U367 ( .A(n519), .B(n520), .Z(n510) );
  AND U368 ( .A(o[6]), .B(n521), .Z(n520) );
  XOR U369 ( .A(n519), .B(n522), .Z(n521) );
  XOR U370 ( .A(n523), .B(n524), .Z(n507) );
  AND U371 ( .A(o[5]), .B(n525), .Z(n524) );
  XNOR U372 ( .A(n523), .B(n526), .Z(n525) );
  XNOR U373 ( .A(n527), .B(n528), .Z(n526) );
  AND U374 ( .A(o[6]), .B(n529), .Z(n527) );
  XOR U375 ( .A(n528), .B(n530), .Z(n529) );
  XOR U376 ( .A(n531), .B(n532), .Z(n523) );
  AND U377 ( .A(o[6]), .B(n533), .Z(n532) );
  XOR U378 ( .A(n531), .B(n534), .Z(n533) );
  XOR U379 ( .A(n535), .B(n536), .Z(n411) );
  AND U380 ( .A(o[3]), .B(n537), .Z(n536) );
  XNOR U381 ( .A(n538), .B(n539), .Z(n537) );
  XNOR U382 ( .A(n540), .B(n535), .Z(n539) );
  AND U383 ( .A(o[4]), .B(n541), .Z(n540) );
  XNOR U384 ( .A(n542), .B(n543), .Z(n541) );
  XNOR U385 ( .A(n544), .B(n538), .Z(n543) );
  AND U386 ( .A(o[5]), .B(n545), .Z(n544) );
  XNOR U387 ( .A(n542), .B(n546), .Z(n545) );
  XNOR U388 ( .A(n547), .B(n548), .Z(n546) );
  AND U389 ( .A(o[6]), .B(n549), .Z(n547) );
  XOR U390 ( .A(n548), .B(n550), .Z(n549) );
  XOR U391 ( .A(n551), .B(n552), .Z(n542) );
  AND U392 ( .A(o[6]), .B(n553), .Z(n552) );
  XOR U393 ( .A(n551), .B(n554), .Z(n553) );
  XOR U394 ( .A(n555), .B(n556), .Z(n538) );
  AND U395 ( .A(o[5]), .B(n557), .Z(n556) );
  XNOR U396 ( .A(n555), .B(n558), .Z(n557) );
  XNOR U397 ( .A(n559), .B(n560), .Z(n558) );
  AND U398 ( .A(o[6]), .B(n561), .Z(n559) );
  XOR U399 ( .A(n560), .B(n562), .Z(n561) );
  XOR U400 ( .A(n563), .B(n564), .Z(n555) );
  AND U401 ( .A(o[6]), .B(n565), .Z(n564) );
  XOR U402 ( .A(n563), .B(n566), .Z(n565) );
  XOR U403 ( .A(n567), .B(n568), .Z(o[3]) );
  AND U404 ( .A(o[4]), .B(n569), .Z(n568) );
  XNOR U405 ( .A(n570), .B(n571), .Z(n569) );
  XNOR U406 ( .A(n572), .B(n567), .Z(n571) );
  AND U407 ( .A(o[5]), .B(n573), .Z(n572) );
  XNOR U408 ( .A(n570), .B(n574), .Z(n573) );
  XNOR U409 ( .A(n575), .B(n576), .Z(n574) );
  AND U410 ( .A(o[6]), .B(n577), .Z(n575) );
  XOR U411 ( .A(n576), .B(n578), .Z(n577) );
  XOR U412 ( .A(n579), .B(n580), .Z(n570) );
  AND U413 ( .A(o[6]), .B(n581), .Z(n580) );
  XOR U414 ( .A(n579), .B(n582), .Z(n581) );
  XOR U415 ( .A(n583), .B(n584), .Z(n567) );
  AND U416 ( .A(o[5]), .B(n585), .Z(n584) );
  XNOR U417 ( .A(n583), .B(n586), .Z(n585) );
  XNOR U418 ( .A(n587), .B(n588), .Z(n586) );
  AND U419 ( .A(o[6]), .B(n589), .Z(n587) );
  XOR U420 ( .A(n588), .B(n590), .Z(n589) );
  XOR U421 ( .A(n591), .B(n592), .Z(n583) );
  AND U422 ( .A(o[6]), .B(n593), .Z(n592) );
  XOR U423 ( .A(n591), .B(n594), .Z(n593) );
  XOR U424 ( .A(n595), .B(n596), .Z(n535) );
  AND U425 ( .A(o[4]), .B(n597), .Z(n596) );
  XNOR U426 ( .A(n598), .B(n599), .Z(n597) );
  XNOR U427 ( .A(n600), .B(n595), .Z(n599) );
  AND U428 ( .A(o[5]), .B(n601), .Z(n600) );
  XNOR U429 ( .A(n598), .B(n602), .Z(n601) );
  XNOR U430 ( .A(n603), .B(n604), .Z(n602) );
  AND U431 ( .A(o[6]), .B(n605), .Z(n603) );
  XOR U432 ( .A(n604), .B(n606), .Z(n605) );
  XOR U433 ( .A(n607), .B(n608), .Z(n598) );
  AND U434 ( .A(o[6]), .B(n609), .Z(n608) );
  XOR U435 ( .A(n607), .B(n610), .Z(n609) );
  XOR U436 ( .A(n611), .B(n612), .Z(o[4]) );
  AND U437 ( .A(o[5]), .B(n613), .Z(n612) );
  XNOR U438 ( .A(n611), .B(n614), .Z(n613) );
  XNOR U439 ( .A(n615), .B(n616), .Z(n614) );
  AND U440 ( .A(o[6]), .B(n617), .Z(n615) );
  XOR U441 ( .A(n616), .B(n618), .Z(n617) );
  XOR U442 ( .A(n619), .B(n620), .Z(n611) );
  AND U443 ( .A(o[6]), .B(n621), .Z(n620) );
  XOR U444 ( .A(n619), .B(n622), .Z(n621) );
  XOR U445 ( .A(n623), .B(n624), .Z(n595) );
  AND U446 ( .A(o[5]), .B(n625), .Z(n624) );
  XNOR U447 ( .A(n623), .B(n626), .Z(n625) );
  XNOR U448 ( .A(n627), .B(n628), .Z(n626) );
  AND U449 ( .A(o[6]), .B(n629), .Z(n627) );
  XOR U450 ( .A(n628), .B(n630), .Z(n629) );
  XOR U451 ( .A(n631), .B(n632), .Z(o[5]) );
  AND U452 ( .A(o[6]), .B(n633), .Z(n632) );
  XOR U453 ( .A(n631), .B(n634), .Z(n633) );
  XOR U454 ( .A(n635), .B(n636), .Z(n623) );
  AND U455 ( .A(o[6]), .B(n637), .Z(n636) );
  XOR U456 ( .A(n635), .B(n638), .Z(n637) );
  XOR U457 ( .A(n639), .B(n640), .Z(o[6]) );
  AND U458 ( .A(n641), .B(n642), .Z(n640) );
  XOR U459 ( .A(n639), .B(n17), .Z(n642) );
  XOR U460 ( .A(n643), .B(n644), .Z(n17) );
  AND U461 ( .A(n634), .B(n645), .Z(n644) );
  XOR U462 ( .A(n646), .B(n643), .Z(n645) );
  XNOR U463 ( .A(n18), .B(n639), .Z(n641) );
  IV U464 ( .A(n15), .Z(n18) );
  XNOR U465 ( .A(n647), .B(n648), .Z(n15) );
  AND U466 ( .A(n631), .B(n649), .Z(n648) );
  XOR U467 ( .A(n650), .B(n647), .Z(n649) );
  XOR U468 ( .A(n651), .B(n652), .Z(n639) );
  AND U469 ( .A(n653), .B(n654), .Z(n652) );
  XOR U470 ( .A(n651), .B(n22), .Z(n654) );
  XOR U471 ( .A(n655), .B(n656), .Z(n22) );
  AND U472 ( .A(n634), .B(n657), .Z(n656) );
  XOR U473 ( .A(n658), .B(n655), .Z(n657) );
  XNOR U474 ( .A(n23), .B(n651), .Z(n653) );
  IV U475 ( .A(n20), .Z(n23) );
  XNOR U476 ( .A(n659), .B(n660), .Z(n20) );
  AND U477 ( .A(n631), .B(n661), .Z(n660) );
  XOR U478 ( .A(n662), .B(n659), .Z(n661) );
  XOR U479 ( .A(n663), .B(n664), .Z(n651) );
  AND U480 ( .A(n665), .B(n666), .Z(n664) );
  XOR U481 ( .A(n663), .B(n27), .Z(n666) );
  XOR U482 ( .A(n667), .B(n668), .Z(n27) );
  AND U483 ( .A(n634), .B(n669), .Z(n668) );
  XOR U484 ( .A(n670), .B(n667), .Z(n669) );
  XNOR U485 ( .A(n28), .B(n663), .Z(n665) );
  IV U486 ( .A(n25), .Z(n28) );
  XNOR U487 ( .A(n671), .B(n672), .Z(n25) );
  AND U488 ( .A(n631), .B(n673), .Z(n672) );
  XOR U489 ( .A(n674), .B(n671), .Z(n673) );
  XOR U490 ( .A(n675), .B(n676), .Z(n663) );
  AND U491 ( .A(n677), .B(n678), .Z(n676) );
  XOR U492 ( .A(n675), .B(n32), .Z(n678) );
  XOR U493 ( .A(n679), .B(n680), .Z(n32) );
  AND U494 ( .A(n634), .B(n681), .Z(n680) );
  XOR U495 ( .A(n682), .B(n679), .Z(n681) );
  XNOR U496 ( .A(n33), .B(n675), .Z(n677) );
  IV U497 ( .A(n30), .Z(n33) );
  XNOR U498 ( .A(n683), .B(n684), .Z(n30) );
  AND U499 ( .A(n631), .B(n685), .Z(n684) );
  XOR U500 ( .A(n686), .B(n683), .Z(n685) );
  XOR U501 ( .A(n687), .B(n688), .Z(n675) );
  AND U502 ( .A(n689), .B(n690), .Z(n688) );
  XOR U503 ( .A(n687), .B(n37), .Z(n690) );
  XOR U504 ( .A(n691), .B(n692), .Z(n37) );
  AND U505 ( .A(n634), .B(n693), .Z(n692) );
  XOR U506 ( .A(n694), .B(n691), .Z(n693) );
  XNOR U507 ( .A(n38), .B(n687), .Z(n689) );
  IV U508 ( .A(n35), .Z(n38) );
  XNOR U509 ( .A(n695), .B(n696), .Z(n35) );
  AND U510 ( .A(n631), .B(n697), .Z(n696) );
  XOR U511 ( .A(n698), .B(n695), .Z(n697) );
  XOR U512 ( .A(n699), .B(n700), .Z(n687) );
  AND U513 ( .A(n701), .B(n702), .Z(n700) );
  XOR U514 ( .A(n699), .B(n42), .Z(n702) );
  XOR U515 ( .A(n703), .B(n704), .Z(n42) );
  AND U516 ( .A(n634), .B(n705), .Z(n704) );
  XOR U517 ( .A(n706), .B(n703), .Z(n705) );
  XNOR U518 ( .A(n43), .B(n699), .Z(n701) );
  IV U519 ( .A(n40), .Z(n43) );
  XNOR U520 ( .A(n707), .B(n708), .Z(n40) );
  AND U521 ( .A(n631), .B(n709), .Z(n708) );
  XOR U522 ( .A(n710), .B(n707), .Z(n709) );
  XOR U523 ( .A(n711), .B(n712), .Z(n699) );
  AND U524 ( .A(n713), .B(n714), .Z(n712) );
  XOR U525 ( .A(n711), .B(n47), .Z(n714) );
  XOR U526 ( .A(n715), .B(n716), .Z(n47) );
  AND U527 ( .A(n634), .B(n717), .Z(n716) );
  XOR U528 ( .A(n718), .B(n715), .Z(n717) );
  XNOR U529 ( .A(n48), .B(n711), .Z(n713) );
  IV U530 ( .A(n45), .Z(n48) );
  XNOR U531 ( .A(n719), .B(n720), .Z(n45) );
  AND U532 ( .A(n631), .B(n721), .Z(n720) );
  XOR U533 ( .A(n722), .B(n719), .Z(n721) );
  XOR U534 ( .A(n723), .B(n724), .Z(n711) );
  AND U535 ( .A(n725), .B(n726), .Z(n724) );
  XOR U536 ( .A(n723), .B(n52), .Z(n726) );
  XOR U537 ( .A(n727), .B(n728), .Z(n52) );
  AND U538 ( .A(n634), .B(n729), .Z(n728) );
  XOR U539 ( .A(n730), .B(n727), .Z(n729) );
  XNOR U540 ( .A(n53), .B(n723), .Z(n725) );
  IV U541 ( .A(n50), .Z(n53) );
  XNOR U542 ( .A(n731), .B(n732), .Z(n50) );
  AND U543 ( .A(n631), .B(n733), .Z(n732) );
  XOR U544 ( .A(n734), .B(n731), .Z(n733) );
  XOR U545 ( .A(n735), .B(n736), .Z(n723) );
  AND U546 ( .A(n737), .B(n738), .Z(n736) );
  XOR U547 ( .A(n735), .B(n57), .Z(n738) );
  XOR U548 ( .A(n739), .B(n740), .Z(n57) );
  AND U549 ( .A(n634), .B(n741), .Z(n740) );
  XOR U550 ( .A(n742), .B(n739), .Z(n741) );
  XNOR U551 ( .A(n58), .B(n735), .Z(n737) );
  IV U552 ( .A(n55), .Z(n58) );
  XNOR U553 ( .A(n743), .B(n744), .Z(n55) );
  AND U554 ( .A(n631), .B(n745), .Z(n744) );
  XOR U555 ( .A(n746), .B(n743), .Z(n745) );
  XOR U556 ( .A(n747), .B(n748), .Z(n735) );
  AND U557 ( .A(n749), .B(n750), .Z(n748) );
  XOR U558 ( .A(n747), .B(n62), .Z(n750) );
  XOR U559 ( .A(n751), .B(n752), .Z(n62) );
  AND U560 ( .A(n634), .B(n753), .Z(n752) );
  XOR U561 ( .A(n754), .B(n751), .Z(n753) );
  XNOR U562 ( .A(n63), .B(n747), .Z(n749) );
  IV U563 ( .A(n60), .Z(n63) );
  XNOR U564 ( .A(n755), .B(n756), .Z(n60) );
  AND U565 ( .A(n631), .B(n757), .Z(n756) );
  XOR U566 ( .A(n758), .B(n755), .Z(n757) );
  XOR U567 ( .A(n759), .B(n760), .Z(n747) );
  AND U568 ( .A(n761), .B(n762), .Z(n760) );
  XOR U569 ( .A(n759), .B(n67), .Z(n762) );
  XOR U570 ( .A(n763), .B(n764), .Z(n67) );
  AND U571 ( .A(n634), .B(n765), .Z(n764) );
  XOR U572 ( .A(n766), .B(n763), .Z(n765) );
  XNOR U573 ( .A(n68), .B(n759), .Z(n761) );
  IV U574 ( .A(n65), .Z(n68) );
  XNOR U575 ( .A(n767), .B(n768), .Z(n65) );
  AND U576 ( .A(n631), .B(n769), .Z(n768) );
  XOR U577 ( .A(n770), .B(n767), .Z(n769) );
  XOR U578 ( .A(n771), .B(n772), .Z(n759) );
  AND U579 ( .A(n773), .B(n774), .Z(n772) );
  XOR U580 ( .A(n771), .B(n72), .Z(n774) );
  XOR U581 ( .A(n775), .B(n776), .Z(n72) );
  AND U582 ( .A(n634), .B(n777), .Z(n776) );
  XOR U583 ( .A(n778), .B(n775), .Z(n777) );
  XNOR U584 ( .A(n73), .B(n771), .Z(n773) );
  IV U585 ( .A(n70), .Z(n73) );
  XNOR U586 ( .A(n779), .B(n780), .Z(n70) );
  AND U587 ( .A(n631), .B(n781), .Z(n780) );
  XOR U588 ( .A(n782), .B(n779), .Z(n781) );
  XOR U589 ( .A(n783), .B(n784), .Z(n771) );
  AND U590 ( .A(n785), .B(n786), .Z(n784) );
  XOR U591 ( .A(n783), .B(n77), .Z(n786) );
  XOR U592 ( .A(n787), .B(n788), .Z(n77) );
  AND U593 ( .A(n634), .B(n789), .Z(n788) );
  XOR U594 ( .A(n790), .B(n787), .Z(n789) );
  XNOR U595 ( .A(n78), .B(n783), .Z(n785) );
  IV U596 ( .A(n75), .Z(n78) );
  XNOR U597 ( .A(n791), .B(n792), .Z(n75) );
  AND U598 ( .A(n631), .B(n793), .Z(n792) );
  XOR U599 ( .A(n794), .B(n791), .Z(n793) );
  XOR U600 ( .A(n795), .B(n796), .Z(n783) );
  AND U601 ( .A(n797), .B(n798), .Z(n796) );
  XOR U602 ( .A(n795), .B(n82), .Z(n798) );
  XOR U603 ( .A(n799), .B(n800), .Z(n82) );
  AND U604 ( .A(n634), .B(n801), .Z(n800) );
  XOR U605 ( .A(n802), .B(n799), .Z(n801) );
  XNOR U606 ( .A(n83), .B(n795), .Z(n797) );
  IV U607 ( .A(n80), .Z(n83) );
  XNOR U608 ( .A(n803), .B(n804), .Z(n80) );
  AND U609 ( .A(n631), .B(n805), .Z(n804) );
  XOR U610 ( .A(n806), .B(n803), .Z(n805) );
  XOR U611 ( .A(n807), .B(n808), .Z(n795) );
  AND U612 ( .A(n809), .B(n810), .Z(n808) );
  XOR U613 ( .A(n807), .B(n87), .Z(n810) );
  XOR U614 ( .A(n811), .B(n812), .Z(n87) );
  AND U615 ( .A(n634), .B(n813), .Z(n812) );
  XOR U616 ( .A(n814), .B(n811), .Z(n813) );
  XNOR U617 ( .A(n88), .B(n807), .Z(n809) );
  IV U618 ( .A(n85), .Z(n88) );
  XNOR U619 ( .A(n815), .B(n816), .Z(n85) );
  AND U620 ( .A(n631), .B(n817), .Z(n816) );
  XOR U621 ( .A(n818), .B(n815), .Z(n817) );
  XOR U622 ( .A(n819), .B(n820), .Z(n807) );
  AND U623 ( .A(n821), .B(n822), .Z(n820) );
  XOR U624 ( .A(n819), .B(n92), .Z(n822) );
  XOR U625 ( .A(n823), .B(n824), .Z(n92) );
  AND U626 ( .A(n634), .B(n825), .Z(n824) );
  XOR U627 ( .A(n826), .B(n823), .Z(n825) );
  XNOR U628 ( .A(n93), .B(n819), .Z(n821) );
  IV U629 ( .A(n90), .Z(n93) );
  XNOR U630 ( .A(n827), .B(n828), .Z(n90) );
  AND U631 ( .A(n631), .B(n829), .Z(n828) );
  XOR U632 ( .A(n830), .B(n827), .Z(n829) );
  XOR U633 ( .A(n831), .B(n832), .Z(n819) );
  AND U634 ( .A(n833), .B(n834), .Z(n832) );
  XOR U635 ( .A(n831), .B(n97), .Z(n834) );
  XOR U636 ( .A(n835), .B(n836), .Z(n97) );
  AND U637 ( .A(n634), .B(n837), .Z(n836) );
  XOR U638 ( .A(n838), .B(n835), .Z(n837) );
  XNOR U639 ( .A(n98), .B(n831), .Z(n833) );
  IV U640 ( .A(n95), .Z(n98) );
  XNOR U641 ( .A(n839), .B(n840), .Z(n95) );
  AND U642 ( .A(n631), .B(n841), .Z(n840) );
  XOR U643 ( .A(n842), .B(n839), .Z(n841) );
  XOR U644 ( .A(n843), .B(n844), .Z(n831) );
  AND U645 ( .A(n845), .B(n846), .Z(n844) );
  XOR U646 ( .A(n843), .B(n102), .Z(n846) );
  XOR U647 ( .A(n847), .B(n848), .Z(n102) );
  AND U648 ( .A(n634), .B(n849), .Z(n848) );
  XOR U649 ( .A(n850), .B(n847), .Z(n849) );
  XNOR U650 ( .A(n103), .B(n843), .Z(n845) );
  IV U651 ( .A(n100), .Z(n103) );
  XNOR U652 ( .A(n851), .B(n852), .Z(n100) );
  AND U653 ( .A(n631), .B(n853), .Z(n852) );
  XOR U654 ( .A(n854), .B(n851), .Z(n853) );
  XOR U655 ( .A(n855), .B(n856), .Z(n843) );
  AND U656 ( .A(n857), .B(n858), .Z(n856) );
  XOR U657 ( .A(n855), .B(n107), .Z(n858) );
  XOR U658 ( .A(n859), .B(n860), .Z(n107) );
  AND U659 ( .A(n634), .B(n861), .Z(n860) );
  XOR U660 ( .A(n862), .B(n859), .Z(n861) );
  XNOR U661 ( .A(n108), .B(n855), .Z(n857) );
  IV U662 ( .A(n105), .Z(n108) );
  XNOR U663 ( .A(n863), .B(n864), .Z(n105) );
  AND U664 ( .A(n631), .B(n865), .Z(n864) );
  XOR U665 ( .A(n866), .B(n863), .Z(n865) );
  XOR U666 ( .A(n867), .B(n868), .Z(n855) );
  AND U667 ( .A(n869), .B(n870), .Z(n868) );
  XOR U668 ( .A(n867), .B(n112), .Z(n870) );
  XOR U669 ( .A(n871), .B(n872), .Z(n112) );
  AND U670 ( .A(n634), .B(n873), .Z(n872) );
  XOR U671 ( .A(n874), .B(n871), .Z(n873) );
  XNOR U672 ( .A(n113), .B(n867), .Z(n869) );
  IV U673 ( .A(n110), .Z(n113) );
  XNOR U674 ( .A(n875), .B(n876), .Z(n110) );
  AND U675 ( .A(n631), .B(n877), .Z(n876) );
  XOR U676 ( .A(n878), .B(n875), .Z(n877) );
  XOR U677 ( .A(n879), .B(n880), .Z(n867) );
  AND U678 ( .A(n881), .B(n882), .Z(n880) );
  XOR U679 ( .A(n879), .B(n117), .Z(n882) );
  XOR U680 ( .A(n883), .B(n884), .Z(n117) );
  AND U681 ( .A(n634), .B(n885), .Z(n884) );
  XOR U682 ( .A(n886), .B(n883), .Z(n885) );
  XNOR U683 ( .A(n118), .B(n879), .Z(n881) );
  IV U684 ( .A(n115), .Z(n118) );
  XNOR U685 ( .A(n887), .B(n888), .Z(n115) );
  AND U686 ( .A(n631), .B(n889), .Z(n888) );
  XOR U687 ( .A(n890), .B(n887), .Z(n889) );
  XOR U688 ( .A(n891), .B(n892), .Z(n879) );
  AND U689 ( .A(n893), .B(n894), .Z(n892) );
  XOR U690 ( .A(n891), .B(n122), .Z(n894) );
  XOR U691 ( .A(n895), .B(n896), .Z(n122) );
  AND U692 ( .A(n634), .B(n897), .Z(n896) );
  XOR U693 ( .A(n898), .B(n895), .Z(n897) );
  XNOR U694 ( .A(n123), .B(n891), .Z(n893) );
  IV U695 ( .A(n120), .Z(n123) );
  XNOR U696 ( .A(n899), .B(n900), .Z(n120) );
  AND U697 ( .A(n631), .B(n901), .Z(n900) );
  XOR U698 ( .A(n902), .B(n899), .Z(n901) );
  XOR U699 ( .A(n903), .B(n904), .Z(n891) );
  AND U700 ( .A(n905), .B(n906), .Z(n904) );
  XOR U701 ( .A(n903), .B(n127), .Z(n906) );
  XOR U702 ( .A(n907), .B(n908), .Z(n127) );
  AND U703 ( .A(n634), .B(n909), .Z(n908) );
  XOR U704 ( .A(n910), .B(n907), .Z(n909) );
  XNOR U705 ( .A(n128), .B(n903), .Z(n905) );
  IV U706 ( .A(n125), .Z(n128) );
  XNOR U707 ( .A(n911), .B(n912), .Z(n125) );
  AND U708 ( .A(n631), .B(n913), .Z(n912) );
  XOR U709 ( .A(n914), .B(n911), .Z(n913) );
  XOR U710 ( .A(n915), .B(n916), .Z(n903) );
  AND U711 ( .A(n917), .B(n918), .Z(n916) );
  XOR U712 ( .A(n915), .B(n132), .Z(n918) );
  XOR U713 ( .A(n919), .B(n920), .Z(n132) );
  AND U714 ( .A(n634), .B(n921), .Z(n920) );
  XOR U715 ( .A(n922), .B(n919), .Z(n921) );
  XNOR U716 ( .A(n133), .B(n915), .Z(n917) );
  IV U717 ( .A(n130), .Z(n133) );
  XNOR U718 ( .A(n923), .B(n924), .Z(n130) );
  AND U719 ( .A(n631), .B(n925), .Z(n924) );
  XOR U720 ( .A(n926), .B(n923), .Z(n925) );
  XOR U721 ( .A(n927), .B(n928), .Z(n915) );
  AND U722 ( .A(n929), .B(n930), .Z(n928) );
  XOR U723 ( .A(n927), .B(n137), .Z(n930) );
  XOR U724 ( .A(n931), .B(n932), .Z(n137) );
  AND U725 ( .A(n634), .B(n933), .Z(n932) );
  XOR U726 ( .A(n934), .B(n931), .Z(n933) );
  XNOR U727 ( .A(n138), .B(n927), .Z(n929) );
  IV U728 ( .A(n135), .Z(n138) );
  XNOR U729 ( .A(n935), .B(n936), .Z(n135) );
  AND U730 ( .A(n631), .B(n937), .Z(n936) );
  XOR U731 ( .A(n938), .B(n935), .Z(n937) );
  XOR U732 ( .A(n939), .B(n940), .Z(n927) );
  AND U733 ( .A(n941), .B(n942), .Z(n940) );
  XOR U734 ( .A(n939), .B(n142), .Z(n942) );
  XOR U735 ( .A(n943), .B(n944), .Z(n142) );
  AND U736 ( .A(n634), .B(n945), .Z(n944) );
  XOR U737 ( .A(n946), .B(n943), .Z(n945) );
  XNOR U738 ( .A(n143), .B(n939), .Z(n941) );
  IV U739 ( .A(n140), .Z(n143) );
  XNOR U740 ( .A(n947), .B(n948), .Z(n140) );
  AND U741 ( .A(n631), .B(n949), .Z(n948) );
  XOR U742 ( .A(n950), .B(n947), .Z(n949) );
  XOR U743 ( .A(n951), .B(n952), .Z(n939) );
  AND U744 ( .A(n953), .B(n954), .Z(n952) );
  XOR U745 ( .A(n951), .B(n147), .Z(n954) );
  XOR U746 ( .A(n955), .B(n956), .Z(n147) );
  AND U747 ( .A(n634), .B(n957), .Z(n956) );
  XOR U748 ( .A(n958), .B(n955), .Z(n957) );
  XNOR U749 ( .A(n148), .B(n951), .Z(n953) );
  IV U750 ( .A(n145), .Z(n148) );
  XNOR U751 ( .A(n959), .B(n960), .Z(n145) );
  AND U752 ( .A(n631), .B(n961), .Z(n960) );
  XOR U753 ( .A(n962), .B(n959), .Z(n961) );
  XOR U754 ( .A(n963), .B(n964), .Z(n951) );
  AND U755 ( .A(n965), .B(n966), .Z(n964) );
  XOR U756 ( .A(n963), .B(n152), .Z(n966) );
  XOR U757 ( .A(n967), .B(n968), .Z(n152) );
  AND U758 ( .A(n634), .B(n969), .Z(n968) );
  XOR U759 ( .A(n970), .B(n967), .Z(n969) );
  XNOR U760 ( .A(n153), .B(n963), .Z(n965) );
  IV U761 ( .A(n150), .Z(n153) );
  XNOR U762 ( .A(n971), .B(n972), .Z(n150) );
  AND U763 ( .A(n631), .B(n973), .Z(n972) );
  XOR U764 ( .A(n974), .B(n971), .Z(n973) );
  XOR U765 ( .A(n975), .B(n976), .Z(n963) );
  AND U766 ( .A(n977), .B(n978), .Z(n976) );
  XOR U767 ( .A(n975), .B(n157), .Z(n978) );
  XOR U768 ( .A(n979), .B(n980), .Z(n157) );
  AND U769 ( .A(n634), .B(n981), .Z(n980) );
  XOR U770 ( .A(n982), .B(n979), .Z(n981) );
  XNOR U771 ( .A(n158), .B(n975), .Z(n977) );
  IV U772 ( .A(n155), .Z(n158) );
  XNOR U773 ( .A(n983), .B(n984), .Z(n155) );
  AND U774 ( .A(n631), .B(n985), .Z(n984) );
  XOR U775 ( .A(n986), .B(n983), .Z(n985) );
  XOR U776 ( .A(n987), .B(n988), .Z(n975) );
  AND U777 ( .A(n989), .B(n990), .Z(n988) );
  XOR U778 ( .A(n4), .B(n987), .Z(n990) );
  XOR U779 ( .A(n991), .B(n992), .Z(n4) );
  AND U780 ( .A(n634), .B(n993), .Z(n992) );
  XOR U781 ( .A(n991), .B(n994), .Z(n993) );
  XNOR U782 ( .A(n987), .B(n2), .Z(n989) );
  XOR U783 ( .A(n995), .B(n996), .Z(n2) );
  AND U784 ( .A(n631), .B(n997), .Z(n996) );
  XOR U785 ( .A(n995), .B(n998), .Z(n997) );
  XNOR U786 ( .A(n999), .B(n1000), .Z(n987) );
  AND U787 ( .A(n1001), .B(n1002), .Z(n1000) );
  XNOR U788 ( .A(n999), .B(n8), .Z(n1002) );
  XOR U789 ( .A(n1003), .B(n1004), .Z(n8) );
  AND U790 ( .A(n634), .B(n1005), .Z(n1004) );
  XOR U791 ( .A(n1006), .B(n1003), .Z(n1005) );
  XOR U792 ( .A(n9), .B(n999), .Z(n1001) );
  IV U793 ( .A(n6), .Z(n9) );
  XNOR U794 ( .A(n1007), .B(n1008), .Z(n6) );
  AND U795 ( .A(n631), .B(n1009), .Z(n1008) );
  XOR U796 ( .A(n1010), .B(n1007), .Z(n1009) );
  AND U797 ( .A(n11), .B(n13), .Z(n999) );
  XNOR U798 ( .A(n1011), .B(n1012), .Z(n13) );
  AND U799 ( .A(n634), .B(n1013), .Z(n1012) );
  XNOR U800 ( .A(n1014), .B(n1011), .Z(n1013) );
  XOR U801 ( .A(n1015), .B(n1016), .Z(n634) );
  AND U802 ( .A(n1017), .B(n1018), .Z(n1016) );
  XOR U803 ( .A(n1015), .B(n646), .Z(n1018) );
  XOR U804 ( .A(n1019), .B(n1020), .Z(n646) );
  AND U805 ( .A(n618), .B(n1021), .Z(n1020) );
  XOR U806 ( .A(n1022), .B(n1019), .Z(n1021) );
  XNOR U807 ( .A(n643), .B(n1015), .Z(n1017) );
  XOR U808 ( .A(n1023), .B(n1024), .Z(n643) );
  AND U809 ( .A(n616), .B(n1025), .Z(n1024) );
  XOR U810 ( .A(n1026), .B(n1023), .Z(n1025) );
  XOR U811 ( .A(n1027), .B(n1028), .Z(n1015) );
  AND U812 ( .A(n1029), .B(n1030), .Z(n1028) );
  XOR U813 ( .A(n1027), .B(n658), .Z(n1030) );
  XOR U814 ( .A(n1031), .B(n1032), .Z(n658) );
  AND U815 ( .A(n618), .B(n1033), .Z(n1032) );
  XOR U816 ( .A(n1034), .B(n1031), .Z(n1033) );
  XNOR U817 ( .A(n655), .B(n1027), .Z(n1029) );
  XOR U818 ( .A(n1035), .B(n1036), .Z(n655) );
  AND U819 ( .A(n616), .B(n1037), .Z(n1036) );
  XOR U820 ( .A(n1038), .B(n1035), .Z(n1037) );
  XOR U821 ( .A(n1039), .B(n1040), .Z(n1027) );
  AND U822 ( .A(n1041), .B(n1042), .Z(n1040) );
  XOR U823 ( .A(n1039), .B(n670), .Z(n1042) );
  XOR U824 ( .A(n1043), .B(n1044), .Z(n670) );
  AND U825 ( .A(n618), .B(n1045), .Z(n1044) );
  XOR U826 ( .A(n1046), .B(n1043), .Z(n1045) );
  XNOR U827 ( .A(n667), .B(n1039), .Z(n1041) );
  XOR U828 ( .A(n1047), .B(n1048), .Z(n667) );
  AND U829 ( .A(n616), .B(n1049), .Z(n1048) );
  XOR U830 ( .A(n1050), .B(n1047), .Z(n1049) );
  XOR U831 ( .A(n1051), .B(n1052), .Z(n1039) );
  AND U832 ( .A(n1053), .B(n1054), .Z(n1052) );
  XOR U833 ( .A(n1051), .B(n682), .Z(n1054) );
  XOR U834 ( .A(n1055), .B(n1056), .Z(n682) );
  AND U835 ( .A(n618), .B(n1057), .Z(n1056) );
  XOR U836 ( .A(n1058), .B(n1055), .Z(n1057) );
  XNOR U837 ( .A(n679), .B(n1051), .Z(n1053) );
  XOR U838 ( .A(n1059), .B(n1060), .Z(n679) );
  AND U839 ( .A(n616), .B(n1061), .Z(n1060) );
  XOR U840 ( .A(n1062), .B(n1059), .Z(n1061) );
  XOR U841 ( .A(n1063), .B(n1064), .Z(n1051) );
  AND U842 ( .A(n1065), .B(n1066), .Z(n1064) );
  XOR U843 ( .A(n1063), .B(n694), .Z(n1066) );
  XOR U844 ( .A(n1067), .B(n1068), .Z(n694) );
  AND U845 ( .A(n618), .B(n1069), .Z(n1068) );
  XOR U846 ( .A(n1070), .B(n1067), .Z(n1069) );
  XNOR U847 ( .A(n691), .B(n1063), .Z(n1065) );
  XOR U848 ( .A(n1071), .B(n1072), .Z(n691) );
  AND U849 ( .A(n616), .B(n1073), .Z(n1072) );
  XOR U850 ( .A(n1074), .B(n1071), .Z(n1073) );
  XOR U851 ( .A(n1075), .B(n1076), .Z(n1063) );
  AND U852 ( .A(n1077), .B(n1078), .Z(n1076) );
  XOR U853 ( .A(n1075), .B(n706), .Z(n1078) );
  XOR U854 ( .A(n1079), .B(n1080), .Z(n706) );
  AND U855 ( .A(n618), .B(n1081), .Z(n1080) );
  XOR U856 ( .A(n1082), .B(n1079), .Z(n1081) );
  XNOR U857 ( .A(n703), .B(n1075), .Z(n1077) );
  XOR U858 ( .A(n1083), .B(n1084), .Z(n703) );
  AND U859 ( .A(n616), .B(n1085), .Z(n1084) );
  XOR U860 ( .A(n1086), .B(n1083), .Z(n1085) );
  XOR U861 ( .A(n1087), .B(n1088), .Z(n1075) );
  AND U862 ( .A(n1089), .B(n1090), .Z(n1088) );
  XOR U863 ( .A(n1087), .B(n718), .Z(n1090) );
  XOR U864 ( .A(n1091), .B(n1092), .Z(n718) );
  AND U865 ( .A(n618), .B(n1093), .Z(n1092) );
  XOR U866 ( .A(n1094), .B(n1091), .Z(n1093) );
  XNOR U867 ( .A(n715), .B(n1087), .Z(n1089) );
  XOR U868 ( .A(n1095), .B(n1096), .Z(n715) );
  AND U869 ( .A(n616), .B(n1097), .Z(n1096) );
  XOR U870 ( .A(n1098), .B(n1095), .Z(n1097) );
  XOR U871 ( .A(n1099), .B(n1100), .Z(n1087) );
  AND U872 ( .A(n1101), .B(n1102), .Z(n1100) );
  XOR U873 ( .A(n1099), .B(n730), .Z(n1102) );
  XOR U874 ( .A(n1103), .B(n1104), .Z(n730) );
  AND U875 ( .A(n618), .B(n1105), .Z(n1104) );
  XOR U876 ( .A(n1106), .B(n1103), .Z(n1105) );
  XNOR U877 ( .A(n727), .B(n1099), .Z(n1101) );
  XOR U878 ( .A(n1107), .B(n1108), .Z(n727) );
  AND U879 ( .A(n616), .B(n1109), .Z(n1108) );
  XOR U880 ( .A(n1110), .B(n1107), .Z(n1109) );
  XOR U881 ( .A(n1111), .B(n1112), .Z(n1099) );
  AND U882 ( .A(n1113), .B(n1114), .Z(n1112) );
  XOR U883 ( .A(n1111), .B(n742), .Z(n1114) );
  XOR U884 ( .A(n1115), .B(n1116), .Z(n742) );
  AND U885 ( .A(n618), .B(n1117), .Z(n1116) );
  XOR U886 ( .A(n1118), .B(n1115), .Z(n1117) );
  XNOR U887 ( .A(n739), .B(n1111), .Z(n1113) );
  XOR U888 ( .A(n1119), .B(n1120), .Z(n739) );
  AND U889 ( .A(n616), .B(n1121), .Z(n1120) );
  XOR U890 ( .A(n1122), .B(n1119), .Z(n1121) );
  XOR U891 ( .A(n1123), .B(n1124), .Z(n1111) );
  AND U892 ( .A(n1125), .B(n1126), .Z(n1124) );
  XOR U893 ( .A(n1123), .B(n754), .Z(n1126) );
  XOR U894 ( .A(n1127), .B(n1128), .Z(n754) );
  AND U895 ( .A(n618), .B(n1129), .Z(n1128) );
  XOR U896 ( .A(n1130), .B(n1127), .Z(n1129) );
  XNOR U897 ( .A(n751), .B(n1123), .Z(n1125) );
  XOR U898 ( .A(n1131), .B(n1132), .Z(n751) );
  AND U899 ( .A(n616), .B(n1133), .Z(n1132) );
  XOR U900 ( .A(n1134), .B(n1131), .Z(n1133) );
  XOR U901 ( .A(n1135), .B(n1136), .Z(n1123) );
  AND U902 ( .A(n1137), .B(n1138), .Z(n1136) );
  XOR U903 ( .A(n1135), .B(n766), .Z(n1138) );
  XOR U904 ( .A(n1139), .B(n1140), .Z(n766) );
  AND U905 ( .A(n618), .B(n1141), .Z(n1140) );
  XOR U906 ( .A(n1142), .B(n1139), .Z(n1141) );
  XNOR U907 ( .A(n763), .B(n1135), .Z(n1137) );
  XOR U908 ( .A(n1143), .B(n1144), .Z(n763) );
  AND U909 ( .A(n616), .B(n1145), .Z(n1144) );
  XOR U910 ( .A(n1146), .B(n1143), .Z(n1145) );
  XOR U911 ( .A(n1147), .B(n1148), .Z(n1135) );
  AND U912 ( .A(n1149), .B(n1150), .Z(n1148) );
  XOR U913 ( .A(n1147), .B(n778), .Z(n1150) );
  XOR U914 ( .A(n1151), .B(n1152), .Z(n778) );
  AND U915 ( .A(n618), .B(n1153), .Z(n1152) );
  XOR U916 ( .A(n1154), .B(n1151), .Z(n1153) );
  XNOR U917 ( .A(n775), .B(n1147), .Z(n1149) );
  XOR U918 ( .A(n1155), .B(n1156), .Z(n775) );
  AND U919 ( .A(n616), .B(n1157), .Z(n1156) );
  XOR U920 ( .A(n1158), .B(n1155), .Z(n1157) );
  XOR U921 ( .A(n1159), .B(n1160), .Z(n1147) );
  AND U922 ( .A(n1161), .B(n1162), .Z(n1160) );
  XOR U923 ( .A(n1159), .B(n790), .Z(n1162) );
  XOR U924 ( .A(n1163), .B(n1164), .Z(n790) );
  AND U925 ( .A(n618), .B(n1165), .Z(n1164) );
  XOR U926 ( .A(n1166), .B(n1163), .Z(n1165) );
  XNOR U927 ( .A(n787), .B(n1159), .Z(n1161) );
  XOR U928 ( .A(n1167), .B(n1168), .Z(n787) );
  AND U929 ( .A(n616), .B(n1169), .Z(n1168) );
  XOR U930 ( .A(n1170), .B(n1167), .Z(n1169) );
  XOR U931 ( .A(n1171), .B(n1172), .Z(n1159) );
  AND U932 ( .A(n1173), .B(n1174), .Z(n1172) );
  XOR U933 ( .A(n1171), .B(n802), .Z(n1174) );
  XOR U934 ( .A(n1175), .B(n1176), .Z(n802) );
  AND U935 ( .A(n618), .B(n1177), .Z(n1176) );
  XOR U936 ( .A(n1178), .B(n1175), .Z(n1177) );
  XNOR U937 ( .A(n799), .B(n1171), .Z(n1173) );
  XOR U938 ( .A(n1179), .B(n1180), .Z(n799) );
  AND U939 ( .A(n616), .B(n1181), .Z(n1180) );
  XOR U940 ( .A(n1182), .B(n1179), .Z(n1181) );
  XOR U941 ( .A(n1183), .B(n1184), .Z(n1171) );
  AND U942 ( .A(n1185), .B(n1186), .Z(n1184) );
  XOR U943 ( .A(n1183), .B(n814), .Z(n1186) );
  XOR U944 ( .A(n1187), .B(n1188), .Z(n814) );
  AND U945 ( .A(n618), .B(n1189), .Z(n1188) );
  XOR U946 ( .A(n1190), .B(n1187), .Z(n1189) );
  XNOR U947 ( .A(n811), .B(n1183), .Z(n1185) );
  XOR U948 ( .A(n1191), .B(n1192), .Z(n811) );
  AND U949 ( .A(n616), .B(n1193), .Z(n1192) );
  XOR U950 ( .A(n1194), .B(n1191), .Z(n1193) );
  XOR U951 ( .A(n1195), .B(n1196), .Z(n1183) );
  AND U952 ( .A(n1197), .B(n1198), .Z(n1196) );
  XOR U953 ( .A(n1195), .B(n826), .Z(n1198) );
  XOR U954 ( .A(n1199), .B(n1200), .Z(n826) );
  AND U955 ( .A(n618), .B(n1201), .Z(n1200) );
  XOR U956 ( .A(n1202), .B(n1199), .Z(n1201) );
  XNOR U957 ( .A(n823), .B(n1195), .Z(n1197) );
  XOR U958 ( .A(n1203), .B(n1204), .Z(n823) );
  AND U959 ( .A(n616), .B(n1205), .Z(n1204) );
  XOR U960 ( .A(n1206), .B(n1203), .Z(n1205) );
  XOR U961 ( .A(n1207), .B(n1208), .Z(n1195) );
  AND U962 ( .A(n1209), .B(n1210), .Z(n1208) );
  XOR U963 ( .A(n1207), .B(n838), .Z(n1210) );
  XOR U964 ( .A(n1211), .B(n1212), .Z(n838) );
  AND U965 ( .A(n618), .B(n1213), .Z(n1212) );
  XOR U966 ( .A(n1214), .B(n1211), .Z(n1213) );
  XNOR U967 ( .A(n835), .B(n1207), .Z(n1209) );
  XOR U968 ( .A(n1215), .B(n1216), .Z(n835) );
  AND U969 ( .A(n616), .B(n1217), .Z(n1216) );
  XOR U970 ( .A(n1218), .B(n1215), .Z(n1217) );
  XOR U971 ( .A(n1219), .B(n1220), .Z(n1207) );
  AND U972 ( .A(n1221), .B(n1222), .Z(n1220) );
  XOR U973 ( .A(n1219), .B(n850), .Z(n1222) );
  XOR U974 ( .A(n1223), .B(n1224), .Z(n850) );
  AND U975 ( .A(n618), .B(n1225), .Z(n1224) );
  XOR U976 ( .A(n1226), .B(n1223), .Z(n1225) );
  XNOR U977 ( .A(n847), .B(n1219), .Z(n1221) );
  XOR U978 ( .A(n1227), .B(n1228), .Z(n847) );
  AND U979 ( .A(n616), .B(n1229), .Z(n1228) );
  XOR U980 ( .A(n1230), .B(n1227), .Z(n1229) );
  XOR U981 ( .A(n1231), .B(n1232), .Z(n1219) );
  AND U982 ( .A(n1233), .B(n1234), .Z(n1232) );
  XOR U983 ( .A(n1231), .B(n862), .Z(n1234) );
  XOR U984 ( .A(n1235), .B(n1236), .Z(n862) );
  AND U985 ( .A(n618), .B(n1237), .Z(n1236) );
  XOR U986 ( .A(n1238), .B(n1235), .Z(n1237) );
  XNOR U987 ( .A(n859), .B(n1231), .Z(n1233) );
  XOR U988 ( .A(n1239), .B(n1240), .Z(n859) );
  AND U989 ( .A(n616), .B(n1241), .Z(n1240) );
  XOR U990 ( .A(n1242), .B(n1239), .Z(n1241) );
  XOR U991 ( .A(n1243), .B(n1244), .Z(n1231) );
  AND U992 ( .A(n1245), .B(n1246), .Z(n1244) );
  XOR U993 ( .A(n1243), .B(n874), .Z(n1246) );
  XOR U994 ( .A(n1247), .B(n1248), .Z(n874) );
  AND U995 ( .A(n618), .B(n1249), .Z(n1248) );
  XOR U996 ( .A(n1250), .B(n1247), .Z(n1249) );
  XNOR U997 ( .A(n871), .B(n1243), .Z(n1245) );
  XOR U998 ( .A(n1251), .B(n1252), .Z(n871) );
  AND U999 ( .A(n616), .B(n1253), .Z(n1252) );
  XOR U1000 ( .A(n1254), .B(n1251), .Z(n1253) );
  XOR U1001 ( .A(n1255), .B(n1256), .Z(n1243) );
  AND U1002 ( .A(n1257), .B(n1258), .Z(n1256) );
  XOR U1003 ( .A(n1255), .B(n886), .Z(n1258) );
  XOR U1004 ( .A(n1259), .B(n1260), .Z(n886) );
  AND U1005 ( .A(n618), .B(n1261), .Z(n1260) );
  XOR U1006 ( .A(n1262), .B(n1259), .Z(n1261) );
  XNOR U1007 ( .A(n883), .B(n1255), .Z(n1257) );
  XOR U1008 ( .A(n1263), .B(n1264), .Z(n883) );
  AND U1009 ( .A(n616), .B(n1265), .Z(n1264) );
  XOR U1010 ( .A(n1266), .B(n1263), .Z(n1265) );
  XOR U1011 ( .A(n1267), .B(n1268), .Z(n1255) );
  AND U1012 ( .A(n1269), .B(n1270), .Z(n1268) );
  XOR U1013 ( .A(n1267), .B(n898), .Z(n1270) );
  XOR U1014 ( .A(n1271), .B(n1272), .Z(n898) );
  AND U1015 ( .A(n618), .B(n1273), .Z(n1272) );
  XOR U1016 ( .A(n1274), .B(n1271), .Z(n1273) );
  XNOR U1017 ( .A(n895), .B(n1267), .Z(n1269) );
  XOR U1018 ( .A(n1275), .B(n1276), .Z(n895) );
  AND U1019 ( .A(n616), .B(n1277), .Z(n1276) );
  XOR U1020 ( .A(n1278), .B(n1275), .Z(n1277) );
  XOR U1021 ( .A(n1279), .B(n1280), .Z(n1267) );
  AND U1022 ( .A(n1281), .B(n1282), .Z(n1280) );
  XOR U1023 ( .A(n1279), .B(n910), .Z(n1282) );
  XOR U1024 ( .A(n1283), .B(n1284), .Z(n910) );
  AND U1025 ( .A(n618), .B(n1285), .Z(n1284) );
  XOR U1026 ( .A(n1286), .B(n1283), .Z(n1285) );
  XNOR U1027 ( .A(n907), .B(n1279), .Z(n1281) );
  XOR U1028 ( .A(n1287), .B(n1288), .Z(n907) );
  AND U1029 ( .A(n616), .B(n1289), .Z(n1288) );
  XOR U1030 ( .A(n1290), .B(n1287), .Z(n1289) );
  XOR U1031 ( .A(n1291), .B(n1292), .Z(n1279) );
  AND U1032 ( .A(n1293), .B(n1294), .Z(n1292) );
  XOR U1033 ( .A(n1291), .B(n922), .Z(n1294) );
  XOR U1034 ( .A(n1295), .B(n1296), .Z(n922) );
  AND U1035 ( .A(n618), .B(n1297), .Z(n1296) );
  XOR U1036 ( .A(n1298), .B(n1295), .Z(n1297) );
  XNOR U1037 ( .A(n919), .B(n1291), .Z(n1293) );
  XOR U1038 ( .A(n1299), .B(n1300), .Z(n919) );
  AND U1039 ( .A(n616), .B(n1301), .Z(n1300) );
  XOR U1040 ( .A(n1302), .B(n1299), .Z(n1301) );
  XOR U1041 ( .A(n1303), .B(n1304), .Z(n1291) );
  AND U1042 ( .A(n1305), .B(n1306), .Z(n1304) );
  XOR U1043 ( .A(n1303), .B(n934), .Z(n1306) );
  XOR U1044 ( .A(n1307), .B(n1308), .Z(n934) );
  AND U1045 ( .A(n618), .B(n1309), .Z(n1308) );
  XOR U1046 ( .A(n1310), .B(n1307), .Z(n1309) );
  XNOR U1047 ( .A(n931), .B(n1303), .Z(n1305) );
  XOR U1048 ( .A(n1311), .B(n1312), .Z(n931) );
  AND U1049 ( .A(n616), .B(n1313), .Z(n1312) );
  XOR U1050 ( .A(n1314), .B(n1311), .Z(n1313) );
  XOR U1051 ( .A(n1315), .B(n1316), .Z(n1303) );
  AND U1052 ( .A(n1317), .B(n1318), .Z(n1316) );
  XOR U1053 ( .A(n1315), .B(n946), .Z(n1318) );
  XOR U1054 ( .A(n1319), .B(n1320), .Z(n946) );
  AND U1055 ( .A(n618), .B(n1321), .Z(n1320) );
  XOR U1056 ( .A(n1322), .B(n1319), .Z(n1321) );
  XNOR U1057 ( .A(n943), .B(n1315), .Z(n1317) );
  XOR U1058 ( .A(n1323), .B(n1324), .Z(n943) );
  AND U1059 ( .A(n616), .B(n1325), .Z(n1324) );
  XOR U1060 ( .A(n1326), .B(n1323), .Z(n1325) );
  XOR U1061 ( .A(n1327), .B(n1328), .Z(n1315) );
  AND U1062 ( .A(n1329), .B(n1330), .Z(n1328) );
  XOR U1063 ( .A(n1327), .B(n958), .Z(n1330) );
  XOR U1064 ( .A(n1331), .B(n1332), .Z(n958) );
  AND U1065 ( .A(n618), .B(n1333), .Z(n1332) );
  XOR U1066 ( .A(n1334), .B(n1331), .Z(n1333) );
  XNOR U1067 ( .A(n955), .B(n1327), .Z(n1329) );
  XOR U1068 ( .A(n1335), .B(n1336), .Z(n955) );
  AND U1069 ( .A(n616), .B(n1337), .Z(n1336) );
  XOR U1070 ( .A(n1338), .B(n1335), .Z(n1337) );
  XOR U1071 ( .A(n1339), .B(n1340), .Z(n1327) );
  AND U1072 ( .A(n1341), .B(n1342), .Z(n1340) );
  XOR U1073 ( .A(n1339), .B(n970), .Z(n1342) );
  XOR U1074 ( .A(n1343), .B(n1344), .Z(n970) );
  AND U1075 ( .A(n618), .B(n1345), .Z(n1344) );
  XOR U1076 ( .A(n1346), .B(n1343), .Z(n1345) );
  XNOR U1077 ( .A(n967), .B(n1339), .Z(n1341) );
  XOR U1078 ( .A(n1347), .B(n1348), .Z(n967) );
  AND U1079 ( .A(n616), .B(n1349), .Z(n1348) );
  XOR U1080 ( .A(n1350), .B(n1347), .Z(n1349) );
  XOR U1081 ( .A(n1351), .B(n1352), .Z(n1339) );
  AND U1082 ( .A(n1353), .B(n1354), .Z(n1352) );
  XOR U1083 ( .A(n1351), .B(n982), .Z(n1354) );
  XOR U1084 ( .A(n1355), .B(n1356), .Z(n982) );
  AND U1085 ( .A(n618), .B(n1357), .Z(n1356) );
  XOR U1086 ( .A(n1358), .B(n1355), .Z(n1357) );
  XNOR U1087 ( .A(n979), .B(n1351), .Z(n1353) );
  XOR U1088 ( .A(n1359), .B(n1360), .Z(n979) );
  AND U1089 ( .A(n616), .B(n1361), .Z(n1360) );
  XOR U1090 ( .A(n1362), .B(n1359), .Z(n1361) );
  XOR U1091 ( .A(n1363), .B(n1364), .Z(n1351) );
  AND U1092 ( .A(n1365), .B(n1366), .Z(n1364) );
  XOR U1093 ( .A(n994), .B(n1363), .Z(n1366) );
  XOR U1094 ( .A(n1367), .B(n1368), .Z(n994) );
  AND U1095 ( .A(n618), .B(n1369), .Z(n1368) );
  XOR U1096 ( .A(n1367), .B(n1370), .Z(n1369) );
  XNOR U1097 ( .A(n1363), .B(n991), .Z(n1365) );
  XOR U1098 ( .A(n1371), .B(n1372), .Z(n991) );
  AND U1099 ( .A(n616), .B(n1373), .Z(n1372) );
  XOR U1100 ( .A(n1371), .B(n1374), .Z(n1373) );
  XOR U1101 ( .A(n1375), .B(n1376), .Z(n1363) );
  AND U1102 ( .A(n1377), .B(n1378), .Z(n1376) );
  XNOR U1103 ( .A(n1379), .B(n1006), .Z(n1378) );
  XOR U1104 ( .A(n1380), .B(n1381), .Z(n1006) );
  AND U1105 ( .A(n618), .B(n1382), .Z(n1381) );
  XOR U1106 ( .A(n1383), .B(n1380), .Z(n1382) );
  XNOR U1107 ( .A(n1003), .B(n1375), .Z(n1377) );
  XOR U1108 ( .A(n1384), .B(n1385), .Z(n1003) );
  AND U1109 ( .A(n616), .B(n1386), .Z(n1385) );
  XOR U1110 ( .A(n1387), .B(n1384), .Z(n1386) );
  IV U1111 ( .A(n1379), .Z(n1375) );
  AND U1112 ( .A(n1011), .B(n1014), .Z(n1379) );
  XNOR U1113 ( .A(n1388), .B(n1389), .Z(n1014) );
  AND U1114 ( .A(n618), .B(n1390), .Z(n1389) );
  XNOR U1115 ( .A(n1391), .B(n1388), .Z(n1390) );
  XOR U1116 ( .A(n1392), .B(n1393), .Z(n618) );
  AND U1117 ( .A(n1394), .B(n1395), .Z(n1393) );
  XOR U1118 ( .A(n1392), .B(n1022), .Z(n1395) );
  XOR U1119 ( .A(n1396), .B(n1397), .Z(n1022) );
  AND U1120 ( .A(n578), .B(n1398), .Z(n1397) );
  XOR U1121 ( .A(n1399), .B(n1396), .Z(n1398) );
  XNOR U1122 ( .A(n1019), .B(n1392), .Z(n1394) );
  XOR U1123 ( .A(n1400), .B(n1401), .Z(n1019) );
  AND U1124 ( .A(n576), .B(n1402), .Z(n1401) );
  XOR U1125 ( .A(n1403), .B(n1400), .Z(n1402) );
  XOR U1126 ( .A(n1404), .B(n1405), .Z(n1392) );
  AND U1127 ( .A(n1406), .B(n1407), .Z(n1405) );
  XOR U1128 ( .A(n1404), .B(n1034), .Z(n1407) );
  XOR U1129 ( .A(n1408), .B(n1409), .Z(n1034) );
  AND U1130 ( .A(n578), .B(n1410), .Z(n1409) );
  XOR U1131 ( .A(n1411), .B(n1408), .Z(n1410) );
  XNOR U1132 ( .A(n1031), .B(n1404), .Z(n1406) );
  XOR U1133 ( .A(n1412), .B(n1413), .Z(n1031) );
  AND U1134 ( .A(n576), .B(n1414), .Z(n1413) );
  XOR U1135 ( .A(n1415), .B(n1412), .Z(n1414) );
  XOR U1136 ( .A(n1416), .B(n1417), .Z(n1404) );
  AND U1137 ( .A(n1418), .B(n1419), .Z(n1417) );
  XOR U1138 ( .A(n1416), .B(n1046), .Z(n1419) );
  XOR U1139 ( .A(n1420), .B(n1421), .Z(n1046) );
  AND U1140 ( .A(n578), .B(n1422), .Z(n1421) );
  XOR U1141 ( .A(n1423), .B(n1420), .Z(n1422) );
  XNOR U1142 ( .A(n1043), .B(n1416), .Z(n1418) );
  XOR U1143 ( .A(n1424), .B(n1425), .Z(n1043) );
  AND U1144 ( .A(n576), .B(n1426), .Z(n1425) );
  XOR U1145 ( .A(n1427), .B(n1424), .Z(n1426) );
  XOR U1146 ( .A(n1428), .B(n1429), .Z(n1416) );
  AND U1147 ( .A(n1430), .B(n1431), .Z(n1429) );
  XOR U1148 ( .A(n1428), .B(n1058), .Z(n1431) );
  XOR U1149 ( .A(n1432), .B(n1433), .Z(n1058) );
  AND U1150 ( .A(n578), .B(n1434), .Z(n1433) );
  XOR U1151 ( .A(n1435), .B(n1432), .Z(n1434) );
  XNOR U1152 ( .A(n1055), .B(n1428), .Z(n1430) );
  XOR U1153 ( .A(n1436), .B(n1437), .Z(n1055) );
  AND U1154 ( .A(n576), .B(n1438), .Z(n1437) );
  XOR U1155 ( .A(n1439), .B(n1436), .Z(n1438) );
  XOR U1156 ( .A(n1440), .B(n1441), .Z(n1428) );
  AND U1157 ( .A(n1442), .B(n1443), .Z(n1441) );
  XOR U1158 ( .A(n1440), .B(n1070), .Z(n1443) );
  XOR U1159 ( .A(n1444), .B(n1445), .Z(n1070) );
  AND U1160 ( .A(n578), .B(n1446), .Z(n1445) );
  XOR U1161 ( .A(n1447), .B(n1444), .Z(n1446) );
  XNOR U1162 ( .A(n1067), .B(n1440), .Z(n1442) );
  XOR U1163 ( .A(n1448), .B(n1449), .Z(n1067) );
  AND U1164 ( .A(n576), .B(n1450), .Z(n1449) );
  XOR U1165 ( .A(n1451), .B(n1448), .Z(n1450) );
  XOR U1166 ( .A(n1452), .B(n1453), .Z(n1440) );
  AND U1167 ( .A(n1454), .B(n1455), .Z(n1453) );
  XOR U1168 ( .A(n1452), .B(n1082), .Z(n1455) );
  XOR U1169 ( .A(n1456), .B(n1457), .Z(n1082) );
  AND U1170 ( .A(n578), .B(n1458), .Z(n1457) );
  XOR U1171 ( .A(n1459), .B(n1456), .Z(n1458) );
  XNOR U1172 ( .A(n1079), .B(n1452), .Z(n1454) );
  XOR U1173 ( .A(n1460), .B(n1461), .Z(n1079) );
  AND U1174 ( .A(n576), .B(n1462), .Z(n1461) );
  XOR U1175 ( .A(n1463), .B(n1460), .Z(n1462) );
  XOR U1176 ( .A(n1464), .B(n1465), .Z(n1452) );
  AND U1177 ( .A(n1466), .B(n1467), .Z(n1465) );
  XOR U1178 ( .A(n1464), .B(n1094), .Z(n1467) );
  XOR U1179 ( .A(n1468), .B(n1469), .Z(n1094) );
  AND U1180 ( .A(n578), .B(n1470), .Z(n1469) );
  XOR U1181 ( .A(n1471), .B(n1468), .Z(n1470) );
  XNOR U1182 ( .A(n1091), .B(n1464), .Z(n1466) );
  XOR U1183 ( .A(n1472), .B(n1473), .Z(n1091) );
  AND U1184 ( .A(n576), .B(n1474), .Z(n1473) );
  XOR U1185 ( .A(n1475), .B(n1472), .Z(n1474) );
  XOR U1186 ( .A(n1476), .B(n1477), .Z(n1464) );
  AND U1187 ( .A(n1478), .B(n1479), .Z(n1477) );
  XOR U1188 ( .A(n1476), .B(n1106), .Z(n1479) );
  XOR U1189 ( .A(n1480), .B(n1481), .Z(n1106) );
  AND U1190 ( .A(n578), .B(n1482), .Z(n1481) );
  XOR U1191 ( .A(n1483), .B(n1480), .Z(n1482) );
  XNOR U1192 ( .A(n1103), .B(n1476), .Z(n1478) );
  XOR U1193 ( .A(n1484), .B(n1485), .Z(n1103) );
  AND U1194 ( .A(n576), .B(n1486), .Z(n1485) );
  XOR U1195 ( .A(n1487), .B(n1484), .Z(n1486) );
  XOR U1196 ( .A(n1488), .B(n1489), .Z(n1476) );
  AND U1197 ( .A(n1490), .B(n1491), .Z(n1489) );
  XOR U1198 ( .A(n1488), .B(n1118), .Z(n1491) );
  XOR U1199 ( .A(n1492), .B(n1493), .Z(n1118) );
  AND U1200 ( .A(n578), .B(n1494), .Z(n1493) );
  XOR U1201 ( .A(n1495), .B(n1492), .Z(n1494) );
  XNOR U1202 ( .A(n1115), .B(n1488), .Z(n1490) );
  XOR U1203 ( .A(n1496), .B(n1497), .Z(n1115) );
  AND U1204 ( .A(n576), .B(n1498), .Z(n1497) );
  XOR U1205 ( .A(n1499), .B(n1496), .Z(n1498) );
  XOR U1206 ( .A(n1500), .B(n1501), .Z(n1488) );
  AND U1207 ( .A(n1502), .B(n1503), .Z(n1501) );
  XOR U1208 ( .A(n1500), .B(n1130), .Z(n1503) );
  XOR U1209 ( .A(n1504), .B(n1505), .Z(n1130) );
  AND U1210 ( .A(n578), .B(n1506), .Z(n1505) );
  XOR U1211 ( .A(n1507), .B(n1504), .Z(n1506) );
  XNOR U1212 ( .A(n1127), .B(n1500), .Z(n1502) );
  XOR U1213 ( .A(n1508), .B(n1509), .Z(n1127) );
  AND U1214 ( .A(n576), .B(n1510), .Z(n1509) );
  XOR U1215 ( .A(n1511), .B(n1508), .Z(n1510) );
  XOR U1216 ( .A(n1512), .B(n1513), .Z(n1500) );
  AND U1217 ( .A(n1514), .B(n1515), .Z(n1513) );
  XOR U1218 ( .A(n1512), .B(n1142), .Z(n1515) );
  XOR U1219 ( .A(n1516), .B(n1517), .Z(n1142) );
  AND U1220 ( .A(n578), .B(n1518), .Z(n1517) );
  XOR U1221 ( .A(n1519), .B(n1516), .Z(n1518) );
  XNOR U1222 ( .A(n1139), .B(n1512), .Z(n1514) );
  XOR U1223 ( .A(n1520), .B(n1521), .Z(n1139) );
  AND U1224 ( .A(n576), .B(n1522), .Z(n1521) );
  XOR U1225 ( .A(n1523), .B(n1520), .Z(n1522) );
  XOR U1226 ( .A(n1524), .B(n1525), .Z(n1512) );
  AND U1227 ( .A(n1526), .B(n1527), .Z(n1525) );
  XOR U1228 ( .A(n1524), .B(n1154), .Z(n1527) );
  XOR U1229 ( .A(n1528), .B(n1529), .Z(n1154) );
  AND U1230 ( .A(n578), .B(n1530), .Z(n1529) );
  XOR U1231 ( .A(n1531), .B(n1528), .Z(n1530) );
  XNOR U1232 ( .A(n1151), .B(n1524), .Z(n1526) );
  XOR U1233 ( .A(n1532), .B(n1533), .Z(n1151) );
  AND U1234 ( .A(n576), .B(n1534), .Z(n1533) );
  XOR U1235 ( .A(n1535), .B(n1532), .Z(n1534) );
  XOR U1236 ( .A(n1536), .B(n1537), .Z(n1524) );
  AND U1237 ( .A(n1538), .B(n1539), .Z(n1537) );
  XOR U1238 ( .A(n1536), .B(n1166), .Z(n1539) );
  XOR U1239 ( .A(n1540), .B(n1541), .Z(n1166) );
  AND U1240 ( .A(n578), .B(n1542), .Z(n1541) );
  XOR U1241 ( .A(n1543), .B(n1540), .Z(n1542) );
  XNOR U1242 ( .A(n1163), .B(n1536), .Z(n1538) );
  XOR U1243 ( .A(n1544), .B(n1545), .Z(n1163) );
  AND U1244 ( .A(n576), .B(n1546), .Z(n1545) );
  XOR U1245 ( .A(n1547), .B(n1544), .Z(n1546) );
  XOR U1246 ( .A(n1548), .B(n1549), .Z(n1536) );
  AND U1247 ( .A(n1550), .B(n1551), .Z(n1549) );
  XOR U1248 ( .A(n1548), .B(n1178), .Z(n1551) );
  XOR U1249 ( .A(n1552), .B(n1553), .Z(n1178) );
  AND U1250 ( .A(n578), .B(n1554), .Z(n1553) );
  XOR U1251 ( .A(n1555), .B(n1552), .Z(n1554) );
  XNOR U1252 ( .A(n1175), .B(n1548), .Z(n1550) );
  XOR U1253 ( .A(n1556), .B(n1557), .Z(n1175) );
  AND U1254 ( .A(n576), .B(n1558), .Z(n1557) );
  XOR U1255 ( .A(n1559), .B(n1556), .Z(n1558) );
  XOR U1256 ( .A(n1560), .B(n1561), .Z(n1548) );
  AND U1257 ( .A(n1562), .B(n1563), .Z(n1561) );
  XOR U1258 ( .A(n1560), .B(n1190), .Z(n1563) );
  XOR U1259 ( .A(n1564), .B(n1565), .Z(n1190) );
  AND U1260 ( .A(n578), .B(n1566), .Z(n1565) );
  XOR U1261 ( .A(n1567), .B(n1564), .Z(n1566) );
  XNOR U1262 ( .A(n1187), .B(n1560), .Z(n1562) );
  XOR U1263 ( .A(n1568), .B(n1569), .Z(n1187) );
  AND U1264 ( .A(n576), .B(n1570), .Z(n1569) );
  XOR U1265 ( .A(n1571), .B(n1568), .Z(n1570) );
  XOR U1266 ( .A(n1572), .B(n1573), .Z(n1560) );
  AND U1267 ( .A(n1574), .B(n1575), .Z(n1573) );
  XOR U1268 ( .A(n1572), .B(n1202), .Z(n1575) );
  XOR U1269 ( .A(n1576), .B(n1577), .Z(n1202) );
  AND U1270 ( .A(n578), .B(n1578), .Z(n1577) );
  XOR U1271 ( .A(n1579), .B(n1576), .Z(n1578) );
  XNOR U1272 ( .A(n1199), .B(n1572), .Z(n1574) );
  XOR U1273 ( .A(n1580), .B(n1581), .Z(n1199) );
  AND U1274 ( .A(n576), .B(n1582), .Z(n1581) );
  XOR U1275 ( .A(n1583), .B(n1580), .Z(n1582) );
  XOR U1276 ( .A(n1584), .B(n1585), .Z(n1572) );
  AND U1277 ( .A(n1586), .B(n1587), .Z(n1585) );
  XOR U1278 ( .A(n1584), .B(n1214), .Z(n1587) );
  XOR U1279 ( .A(n1588), .B(n1589), .Z(n1214) );
  AND U1280 ( .A(n578), .B(n1590), .Z(n1589) );
  XOR U1281 ( .A(n1591), .B(n1588), .Z(n1590) );
  XNOR U1282 ( .A(n1211), .B(n1584), .Z(n1586) );
  XOR U1283 ( .A(n1592), .B(n1593), .Z(n1211) );
  AND U1284 ( .A(n576), .B(n1594), .Z(n1593) );
  XOR U1285 ( .A(n1595), .B(n1592), .Z(n1594) );
  XOR U1286 ( .A(n1596), .B(n1597), .Z(n1584) );
  AND U1287 ( .A(n1598), .B(n1599), .Z(n1597) );
  XOR U1288 ( .A(n1596), .B(n1226), .Z(n1599) );
  XOR U1289 ( .A(n1600), .B(n1601), .Z(n1226) );
  AND U1290 ( .A(n578), .B(n1602), .Z(n1601) );
  XOR U1291 ( .A(n1603), .B(n1600), .Z(n1602) );
  XNOR U1292 ( .A(n1223), .B(n1596), .Z(n1598) );
  XOR U1293 ( .A(n1604), .B(n1605), .Z(n1223) );
  AND U1294 ( .A(n576), .B(n1606), .Z(n1605) );
  XOR U1295 ( .A(n1607), .B(n1604), .Z(n1606) );
  XOR U1296 ( .A(n1608), .B(n1609), .Z(n1596) );
  AND U1297 ( .A(n1610), .B(n1611), .Z(n1609) );
  XOR U1298 ( .A(n1608), .B(n1238), .Z(n1611) );
  XOR U1299 ( .A(n1612), .B(n1613), .Z(n1238) );
  AND U1300 ( .A(n578), .B(n1614), .Z(n1613) );
  XOR U1301 ( .A(n1615), .B(n1612), .Z(n1614) );
  XNOR U1302 ( .A(n1235), .B(n1608), .Z(n1610) );
  XOR U1303 ( .A(n1616), .B(n1617), .Z(n1235) );
  AND U1304 ( .A(n576), .B(n1618), .Z(n1617) );
  XOR U1305 ( .A(n1619), .B(n1616), .Z(n1618) );
  XOR U1306 ( .A(n1620), .B(n1621), .Z(n1608) );
  AND U1307 ( .A(n1622), .B(n1623), .Z(n1621) );
  XOR U1308 ( .A(n1620), .B(n1250), .Z(n1623) );
  XOR U1309 ( .A(n1624), .B(n1625), .Z(n1250) );
  AND U1310 ( .A(n578), .B(n1626), .Z(n1625) );
  XOR U1311 ( .A(n1627), .B(n1624), .Z(n1626) );
  XNOR U1312 ( .A(n1247), .B(n1620), .Z(n1622) );
  XOR U1313 ( .A(n1628), .B(n1629), .Z(n1247) );
  AND U1314 ( .A(n576), .B(n1630), .Z(n1629) );
  XOR U1315 ( .A(n1631), .B(n1628), .Z(n1630) );
  XOR U1316 ( .A(n1632), .B(n1633), .Z(n1620) );
  AND U1317 ( .A(n1634), .B(n1635), .Z(n1633) );
  XOR U1318 ( .A(n1632), .B(n1262), .Z(n1635) );
  XOR U1319 ( .A(n1636), .B(n1637), .Z(n1262) );
  AND U1320 ( .A(n578), .B(n1638), .Z(n1637) );
  XOR U1321 ( .A(n1639), .B(n1636), .Z(n1638) );
  XNOR U1322 ( .A(n1259), .B(n1632), .Z(n1634) );
  XOR U1323 ( .A(n1640), .B(n1641), .Z(n1259) );
  AND U1324 ( .A(n576), .B(n1642), .Z(n1641) );
  XOR U1325 ( .A(n1643), .B(n1640), .Z(n1642) );
  XOR U1326 ( .A(n1644), .B(n1645), .Z(n1632) );
  AND U1327 ( .A(n1646), .B(n1647), .Z(n1645) );
  XOR U1328 ( .A(n1644), .B(n1274), .Z(n1647) );
  XOR U1329 ( .A(n1648), .B(n1649), .Z(n1274) );
  AND U1330 ( .A(n578), .B(n1650), .Z(n1649) );
  XOR U1331 ( .A(n1651), .B(n1648), .Z(n1650) );
  XNOR U1332 ( .A(n1271), .B(n1644), .Z(n1646) );
  XOR U1333 ( .A(n1652), .B(n1653), .Z(n1271) );
  AND U1334 ( .A(n576), .B(n1654), .Z(n1653) );
  XOR U1335 ( .A(n1655), .B(n1652), .Z(n1654) );
  XOR U1336 ( .A(n1656), .B(n1657), .Z(n1644) );
  AND U1337 ( .A(n1658), .B(n1659), .Z(n1657) );
  XOR U1338 ( .A(n1656), .B(n1286), .Z(n1659) );
  XOR U1339 ( .A(n1660), .B(n1661), .Z(n1286) );
  AND U1340 ( .A(n578), .B(n1662), .Z(n1661) );
  XOR U1341 ( .A(n1663), .B(n1660), .Z(n1662) );
  XNOR U1342 ( .A(n1283), .B(n1656), .Z(n1658) );
  XOR U1343 ( .A(n1664), .B(n1665), .Z(n1283) );
  AND U1344 ( .A(n576), .B(n1666), .Z(n1665) );
  XOR U1345 ( .A(n1667), .B(n1664), .Z(n1666) );
  XOR U1346 ( .A(n1668), .B(n1669), .Z(n1656) );
  AND U1347 ( .A(n1670), .B(n1671), .Z(n1669) );
  XOR U1348 ( .A(n1668), .B(n1298), .Z(n1671) );
  XOR U1349 ( .A(n1672), .B(n1673), .Z(n1298) );
  AND U1350 ( .A(n578), .B(n1674), .Z(n1673) );
  XOR U1351 ( .A(n1675), .B(n1672), .Z(n1674) );
  XNOR U1352 ( .A(n1295), .B(n1668), .Z(n1670) );
  XOR U1353 ( .A(n1676), .B(n1677), .Z(n1295) );
  AND U1354 ( .A(n576), .B(n1678), .Z(n1677) );
  XOR U1355 ( .A(n1679), .B(n1676), .Z(n1678) );
  XOR U1356 ( .A(n1680), .B(n1681), .Z(n1668) );
  AND U1357 ( .A(n1682), .B(n1683), .Z(n1681) );
  XOR U1358 ( .A(n1680), .B(n1310), .Z(n1683) );
  XOR U1359 ( .A(n1684), .B(n1685), .Z(n1310) );
  AND U1360 ( .A(n578), .B(n1686), .Z(n1685) );
  XOR U1361 ( .A(n1687), .B(n1684), .Z(n1686) );
  XNOR U1362 ( .A(n1307), .B(n1680), .Z(n1682) );
  XOR U1363 ( .A(n1688), .B(n1689), .Z(n1307) );
  AND U1364 ( .A(n576), .B(n1690), .Z(n1689) );
  XOR U1365 ( .A(n1691), .B(n1688), .Z(n1690) );
  XOR U1366 ( .A(n1692), .B(n1693), .Z(n1680) );
  AND U1367 ( .A(n1694), .B(n1695), .Z(n1693) );
  XOR U1368 ( .A(n1692), .B(n1322), .Z(n1695) );
  XOR U1369 ( .A(n1696), .B(n1697), .Z(n1322) );
  AND U1370 ( .A(n578), .B(n1698), .Z(n1697) );
  XOR U1371 ( .A(n1699), .B(n1696), .Z(n1698) );
  XNOR U1372 ( .A(n1319), .B(n1692), .Z(n1694) );
  XOR U1373 ( .A(n1700), .B(n1701), .Z(n1319) );
  AND U1374 ( .A(n576), .B(n1702), .Z(n1701) );
  XOR U1375 ( .A(n1703), .B(n1700), .Z(n1702) );
  XOR U1376 ( .A(n1704), .B(n1705), .Z(n1692) );
  AND U1377 ( .A(n1706), .B(n1707), .Z(n1705) );
  XOR U1378 ( .A(n1704), .B(n1334), .Z(n1707) );
  XOR U1379 ( .A(n1708), .B(n1709), .Z(n1334) );
  AND U1380 ( .A(n578), .B(n1710), .Z(n1709) );
  XOR U1381 ( .A(n1711), .B(n1708), .Z(n1710) );
  XNOR U1382 ( .A(n1331), .B(n1704), .Z(n1706) );
  XOR U1383 ( .A(n1712), .B(n1713), .Z(n1331) );
  AND U1384 ( .A(n576), .B(n1714), .Z(n1713) );
  XOR U1385 ( .A(n1715), .B(n1712), .Z(n1714) );
  XOR U1386 ( .A(n1716), .B(n1717), .Z(n1704) );
  AND U1387 ( .A(n1718), .B(n1719), .Z(n1717) );
  XOR U1388 ( .A(n1716), .B(n1346), .Z(n1719) );
  XOR U1389 ( .A(n1720), .B(n1721), .Z(n1346) );
  AND U1390 ( .A(n578), .B(n1722), .Z(n1721) );
  XOR U1391 ( .A(n1723), .B(n1720), .Z(n1722) );
  XNOR U1392 ( .A(n1343), .B(n1716), .Z(n1718) );
  XOR U1393 ( .A(n1724), .B(n1725), .Z(n1343) );
  AND U1394 ( .A(n576), .B(n1726), .Z(n1725) );
  XOR U1395 ( .A(n1727), .B(n1724), .Z(n1726) );
  XOR U1396 ( .A(n1728), .B(n1729), .Z(n1716) );
  AND U1397 ( .A(n1730), .B(n1731), .Z(n1729) );
  XOR U1398 ( .A(n1728), .B(n1358), .Z(n1731) );
  XOR U1399 ( .A(n1732), .B(n1733), .Z(n1358) );
  AND U1400 ( .A(n578), .B(n1734), .Z(n1733) );
  XOR U1401 ( .A(n1735), .B(n1732), .Z(n1734) );
  XNOR U1402 ( .A(n1355), .B(n1728), .Z(n1730) );
  XOR U1403 ( .A(n1736), .B(n1737), .Z(n1355) );
  AND U1404 ( .A(n576), .B(n1738), .Z(n1737) );
  XOR U1405 ( .A(n1739), .B(n1736), .Z(n1738) );
  XOR U1406 ( .A(n1740), .B(n1741), .Z(n1728) );
  AND U1407 ( .A(n1742), .B(n1743), .Z(n1741) );
  XOR U1408 ( .A(n1370), .B(n1740), .Z(n1743) );
  XOR U1409 ( .A(n1744), .B(n1745), .Z(n1370) );
  AND U1410 ( .A(n578), .B(n1746), .Z(n1745) );
  XOR U1411 ( .A(n1744), .B(n1747), .Z(n1746) );
  XNOR U1412 ( .A(n1740), .B(n1367), .Z(n1742) );
  XOR U1413 ( .A(n1748), .B(n1749), .Z(n1367) );
  AND U1414 ( .A(n576), .B(n1750), .Z(n1749) );
  XOR U1415 ( .A(n1748), .B(n1751), .Z(n1750) );
  XOR U1416 ( .A(n1752), .B(n1753), .Z(n1740) );
  AND U1417 ( .A(n1754), .B(n1755), .Z(n1753) );
  XNOR U1418 ( .A(n1756), .B(n1383), .Z(n1755) );
  XOR U1419 ( .A(n1757), .B(n1758), .Z(n1383) );
  AND U1420 ( .A(n578), .B(n1759), .Z(n1758) );
  XOR U1421 ( .A(n1760), .B(n1757), .Z(n1759) );
  XNOR U1422 ( .A(n1380), .B(n1752), .Z(n1754) );
  XOR U1423 ( .A(n1761), .B(n1762), .Z(n1380) );
  AND U1424 ( .A(n576), .B(n1763), .Z(n1762) );
  XOR U1425 ( .A(n1764), .B(n1761), .Z(n1763) );
  IV U1426 ( .A(n1756), .Z(n1752) );
  AND U1427 ( .A(n1388), .B(n1391), .Z(n1756) );
  XNOR U1428 ( .A(n1765), .B(n1766), .Z(n1391) );
  AND U1429 ( .A(n578), .B(n1767), .Z(n1766) );
  XNOR U1430 ( .A(n1768), .B(n1765), .Z(n1767) );
  XOR U1431 ( .A(n1769), .B(n1770), .Z(n578) );
  AND U1432 ( .A(n1771), .B(n1772), .Z(n1770) );
  XOR U1433 ( .A(n1769), .B(n1399), .Z(n1772) );
  XOR U1434 ( .A(n1773), .B(n1774), .Z(n1399) );
  AND U1435 ( .A(n490), .B(n1775), .Z(n1774) );
  XOR U1436 ( .A(n1776), .B(n1773), .Z(n1775) );
  XNOR U1437 ( .A(n1396), .B(n1769), .Z(n1771) );
  XOR U1438 ( .A(n1777), .B(n1778), .Z(n1396) );
  AND U1439 ( .A(n488), .B(n1779), .Z(n1778) );
  XOR U1440 ( .A(n1780), .B(n1777), .Z(n1779) );
  XOR U1441 ( .A(n1781), .B(n1782), .Z(n1769) );
  AND U1442 ( .A(n1783), .B(n1784), .Z(n1782) );
  XOR U1443 ( .A(n1781), .B(n1411), .Z(n1784) );
  XOR U1444 ( .A(n1785), .B(n1786), .Z(n1411) );
  AND U1445 ( .A(n490), .B(n1787), .Z(n1786) );
  XOR U1446 ( .A(n1788), .B(n1785), .Z(n1787) );
  XNOR U1447 ( .A(n1408), .B(n1781), .Z(n1783) );
  XOR U1448 ( .A(n1789), .B(n1790), .Z(n1408) );
  AND U1449 ( .A(n488), .B(n1791), .Z(n1790) );
  XOR U1450 ( .A(n1792), .B(n1789), .Z(n1791) );
  XOR U1451 ( .A(n1793), .B(n1794), .Z(n1781) );
  AND U1452 ( .A(n1795), .B(n1796), .Z(n1794) );
  XOR U1453 ( .A(n1793), .B(n1423), .Z(n1796) );
  XOR U1454 ( .A(n1797), .B(n1798), .Z(n1423) );
  AND U1455 ( .A(n490), .B(n1799), .Z(n1798) );
  XOR U1456 ( .A(n1800), .B(n1797), .Z(n1799) );
  XNOR U1457 ( .A(n1420), .B(n1793), .Z(n1795) );
  XOR U1458 ( .A(n1801), .B(n1802), .Z(n1420) );
  AND U1459 ( .A(n488), .B(n1803), .Z(n1802) );
  XOR U1460 ( .A(n1804), .B(n1801), .Z(n1803) );
  XOR U1461 ( .A(n1805), .B(n1806), .Z(n1793) );
  AND U1462 ( .A(n1807), .B(n1808), .Z(n1806) );
  XOR U1463 ( .A(n1805), .B(n1435), .Z(n1808) );
  XOR U1464 ( .A(n1809), .B(n1810), .Z(n1435) );
  AND U1465 ( .A(n490), .B(n1811), .Z(n1810) );
  XOR U1466 ( .A(n1812), .B(n1809), .Z(n1811) );
  XNOR U1467 ( .A(n1432), .B(n1805), .Z(n1807) );
  XOR U1468 ( .A(n1813), .B(n1814), .Z(n1432) );
  AND U1469 ( .A(n488), .B(n1815), .Z(n1814) );
  XOR U1470 ( .A(n1816), .B(n1813), .Z(n1815) );
  XOR U1471 ( .A(n1817), .B(n1818), .Z(n1805) );
  AND U1472 ( .A(n1819), .B(n1820), .Z(n1818) );
  XOR U1473 ( .A(n1817), .B(n1447), .Z(n1820) );
  XOR U1474 ( .A(n1821), .B(n1822), .Z(n1447) );
  AND U1475 ( .A(n490), .B(n1823), .Z(n1822) );
  XOR U1476 ( .A(n1824), .B(n1821), .Z(n1823) );
  XNOR U1477 ( .A(n1444), .B(n1817), .Z(n1819) );
  XOR U1478 ( .A(n1825), .B(n1826), .Z(n1444) );
  AND U1479 ( .A(n488), .B(n1827), .Z(n1826) );
  XOR U1480 ( .A(n1828), .B(n1825), .Z(n1827) );
  XOR U1481 ( .A(n1829), .B(n1830), .Z(n1817) );
  AND U1482 ( .A(n1831), .B(n1832), .Z(n1830) );
  XOR U1483 ( .A(n1829), .B(n1459), .Z(n1832) );
  XOR U1484 ( .A(n1833), .B(n1834), .Z(n1459) );
  AND U1485 ( .A(n490), .B(n1835), .Z(n1834) );
  XOR U1486 ( .A(n1836), .B(n1833), .Z(n1835) );
  XNOR U1487 ( .A(n1456), .B(n1829), .Z(n1831) );
  XOR U1488 ( .A(n1837), .B(n1838), .Z(n1456) );
  AND U1489 ( .A(n488), .B(n1839), .Z(n1838) );
  XOR U1490 ( .A(n1840), .B(n1837), .Z(n1839) );
  XOR U1491 ( .A(n1841), .B(n1842), .Z(n1829) );
  AND U1492 ( .A(n1843), .B(n1844), .Z(n1842) );
  XOR U1493 ( .A(n1841), .B(n1471), .Z(n1844) );
  XOR U1494 ( .A(n1845), .B(n1846), .Z(n1471) );
  AND U1495 ( .A(n490), .B(n1847), .Z(n1846) );
  XOR U1496 ( .A(n1848), .B(n1845), .Z(n1847) );
  XNOR U1497 ( .A(n1468), .B(n1841), .Z(n1843) );
  XOR U1498 ( .A(n1849), .B(n1850), .Z(n1468) );
  AND U1499 ( .A(n488), .B(n1851), .Z(n1850) );
  XOR U1500 ( .A(n1852), .B(n1849), .Z(n1851) );
  XOR U1501 ( .A(n1853), .B(n1854), .Z(n1841) );
  AND U1502 ( .A(n1855), .B(n1856), .Z(n1854) );
  XOR U1503 ( .A(n1853), .B(n1483), .Z(n1856) );
  XOR U1504 ( .A(n1857), .B(n1858), .Z(n1483) );
  AND U1505 ( .A(n490), .B(n1859), .Z(n1858) );
  XOR U1506 ( .A(n1860), .B(n1857), .Z(n1859) );
  XNOR U1507 ( .A(n1480), .B(n1853), .Z(n1855) );
  XOR U1508 ( .A(n1861), .B(n1862), .Z(n1480) );
  AND U1509 ( .A(n488), .B(n1863), .Z(n1862) );
  XOR U1510 ( .A(n1864), .B(n1861), .Z(n1863) );
  XOR U1511 ( .A(n1865), .B(n1866), .Z(n1853) );
  AND U1512 ( .A(n1867), .B(n1868), .Z(n1866) );
  XOR U1513 ( .A(n1865), .B(n1495), .Z(n1868) );
  XOR U1514 ( .A(n1869), .B(n1870), .Z(n1495) );
  AND U1515 ( .A(n490), .B(n1871), .Z(n1870) );
  XOR U1516 ( .A(n1872), .B(n1869), .Z(n1871) );
  XNOR U1517 ( .A(n1492), .B(n1865), .Z(n1867) );
  XOR U1518 ( .A(n1873), .B(n1874), .Z(n1492) );
  AND U1519 ( .A(n488), .B(n1875), .Z(n1874) );
  XOR U1520 ( .A(n1876), .B(n1873), .Z(n1875) );
  XOR U1521 ( .A(n1877), .B(n1878), .Z(n1865) );
  AND U1522 ( .A(n1879), .B(n1880), .Z(n1878) );
  XOR U1523 ( .A(n1877), .B(n1507), .Z(n1880) );
  XOR U1524 ( .A(n1881), .B(n1882), .Z(n1507) );
  AND U1525 ( .A(n490), .B(n1883), .Z(n1882) );
  XOR U1526 ( .A(n1884), .B(n1881), .Z(n1883) );
  XNOR U1527 ( .A(n1504), .B(n1877), .Z(n1879) );
  XOR U1528 ( .A(n1885), .B(n1886), .Z(n1504) );
  AND U1529 ( .A(n488), .B(n1887), .Z(n1886) );
  XOR U1530 ( .A(n1888), .B(n1885), .Z(n1887) );
  XOR U1531 ( .A(n1889), .B(n1890), .Z(n1877) );
  AND U1532 ( .A(n1891), .B(n1892), .Z(n1890) );
  XOR U1533 ( .A(n1889), .B(n1519), .Z(n1892) );
  XOR U1534 ( .A(n1893), .B(n1894), .Z(n1519) );
  AND U1535 ( .A(n490), .B(n1895), .Z(n1894) );
  XOR U1536 ( .A(n1896), .B(n1893), .Z(n1895) );
  XNOR U1537 ( .A(n1516), .B(n1889), .Z(n1891) );
  XOR U1538 ( .A(n1897), .B(n1898), .Z(n1516) );
  AND U1539 ( .A(n488), .B(n1899), .Z(n1898) );
  XOR U1540 ( .A(n1900), .B(n1897), .Z(n1899) );
  XOR U1541 ( .A(n1901), .B(n1902), .Z(n1889) );
  AND U1542 ( .A(n1903), .B(n1904), .Z(n1902) );
  XOR U1543 ( .A(n1901), .B(n1531), .Z(n1904) );
  XOR U1544 ( .A(n1905), .B(n1906), .Z(n1531) );
  AND U1545 ( .A(n490), .B(n1907), .Z(n1906) );
  XOR U1546 ( .A(n1908), .B(n1905), .Z(n1907) );
  XNOR U1547 ( .A(n1528), .B(n1901), .Z(n1903) );
  XOR U1548 ( .A(n1909), .B(n1910), .Z(n1528) );
  AND U1549 ( .A(n488), .B(n1911), .Z(n1910) );
  XOR U1550 ( .A(n1912), .B(n1909), .Z(n1911) );
  XOR U1551 ( .A(n1913), .B(n1914), .Z(n1901) );
  AND U1552 ( .A(n1915), .B(n1916), .Z(n1914) );
  XOR U1553 ( .A(n1913), .B(n1543), .Z(n1916) );
  XOR U1554 ( .A(n1917), .B(n1918), .Z(n1543) );
  AND U1555 ( .A(n490), .B(n1919), .Z(n1918) );
  XOR U1556 ( .A(n1920), .B(n1917), .Z(n1919) );
  XNOR U1557 ( .A(n1540), .B(n1913), .Z(n1915) );
  XOR U1558 ( .A(n1921), .B(n1922), .Z(n1540) );
  AND U1559 ( .A(n488), .B(n1923), .Z(n1922) );
  XOR U1560 ( .A(n1924), .B(n1921), .Z(n1923) );
  XOR U1561 ( .A(n1925), .B(n1926), .Z(n1913) );
  AND U1562 ( .A(n1927), .B(n1928), .Z(n1926) );
  XOR U1563 ( .A(n1925), .B(n1555), .Z(n1928) );
  XOR U1564 ( .A(n1929), .B(n1930), .Z(n1555) );
  AND U1565 ( .A(n490), .B(n1931), .Z(n1930) );
  XOR U1566 ( .A(n1932), .B(n1929), .Z(n1931) );
  XNOR U1567 ( .A(n1552), .B(n1925), .Z(n1927) );
  XOR U1568 ( .A(n1933), .B(n1934), .Z(n1552) );
  AND U1569 ( .A(n488), .B(n1935), .Z(n1934) );
  XOR U1570 ( .A(n1936), .B(n1933), .Z(n1935) );
  XOR U1571 ( .A(n1937), .B(n1938), .Z(n1925) );
  AND U1572 ( .A(n1939), .B(n1940), .Z(n1938) );
  XOR U1573 ( .A(n1937), .B(n1567), .Z(n1940) );
  XOR U1574 ( .A(n1941), .B(n1942), .Z(n1567) );
  AND U1575 ( .A(n490), .B(n1943), .Z(n1942) );
  XOR U1576 ( .A(n1944), .B(n1941), .Z(n1943) );
  XNOR U1577 ( .A(n1564), .B(n1937), .Z(n1939) );
  XOR U1578 ( .A(n1945), .B(n1946), .Z(n1564) );
  AND U1579 ( .A(n488), .B(n1947), .Z(n1946) );
  XOR U1580 ( .A(n1948), .B(n1945), .Z(n1947) );
  XOR U1581 ( .A(n1949), .B(n1950), .Z(n1937) );
  AND U1582 ( .A(n1951), .B(n1952), .Z(n1950) );
  XOR U1583 ( .A(n1949), .B(n1579), .Z(n1952) );
  XOR U1584 ( .A(n1953), .B(n1954), .Z(n1579) );
  AND U1585 ( .A(n490), .B(n1955), .Z(n1954) );
  XOR U1586 ( .A(n1956), .B(n1953), .Z(n1955) );
  XNOR U1587 ( .A(n1576), .B(n1949), .Z(n1951) );
  XOR U1588 ( .A(n1957), .B(n1958), .Z(n1576) );
  AND U1589 ( .A(n488), .B(n1959), .Z(n1958) );
  XOR U1590 ( .A(n1960), .B(n1957), .Z(n1959) );
  XOR U1591 ( .A(n1961), .B(n1962), .Z(n1949) );
  AND U1592 ( .A(n1963), .B(n1964), .Z(n1962) );
  XOR U1593 ( .A(n1961), .B(n1591), .Z(n1964) );
  XOR U1594 ( .A(n1965), .B(n1966), .Z(n1591) );
  AND U1595 ( .A(n490), .B(n1967), .Z(n1966) );
  XOR U1596 ( .A(n1968), .B(n1965), .Z(n1967) );
  XNOR U1597 ( .A(n1588), .B(n1961), .Z(n1963) );
  XOR U1598 ( .A(n1969), .B(n1970), .Z(n1588) );
  AND U1599 ( .A(n488), .B(n1971), .Z(n1970) );
  XOR U1600 ( .A(n1972), .B(n1969), .Z(n1971) );
  XOR U1601 ( .A(n1973), .B(n1974), .Z(n1961) );
  AND U1602 ( .A(n1975), .B(n1976), .Z(n1974) );
  XOR U1603 ( .A(n1973), .B(n1603), .Z(n1976) );
  XOR U1604 ( .A(n1977), .B(n1978), .Z(n1603) );
  AND U1605 ( .A(n490), .B(n1979), .Z(n1978) );
  XOR U1606 ( .A(n1980), .B(n1977), .Z(n1979) );
  XNOR U1607 ( .A(n1600), .B(n1973), .Z(n1975) );
  XOR U1608 ( .A(n1981), .B(n1982), .Z(n1600) );
  AND U1609 ( .A(n488), .B(n1983), .Z(n1982) );
  XOR U1610 ( .A(n1984), .B(n1981), .Z(n1983) );
  XOR U1611 ( .A(n1985), .B(n1986), .Z(n1973) );
  AND U1612 ( .A(n1987), .B(n1988), .Z(n1986) );
  XOR U1613 ( .A(n1985), .B(n1615), .Z(n1988) );
  XOR U1614 ( .A(n1989), .B(n1990), .Z(n1615) );
  AND U1615 ( .A(n490), .B(n1991), .Z(n1990) );
  XOR U1616 ( .A(n1992), .B(n1989), .Z(n1991) );
  XNOR U1617 ( .A(n1612), .B(n1985), .Z(n1987) );
  XOR U1618 ( .A(n1993), .B(n1994), .Z(n1612) );
  AND U1619 ( .A(n488), .B(n1995), .Z(n1994) );
  XOR U1620 ( .A(n1996), .B(n1993), .Z(n1995) );
  XOR U1621 ( .A(n1997), .B(n1998), .Z(n1985) );
  AND U1622 ( .A(n1999), .B(n2000), .Z(n1998) );
  XOR U1623 ( .A(n1997), .B(n1627), .Z(n2000) );
  XOR U1624 ( .A(n2001), .B(n2002), .Z(n1627) );
  AND U1625 ( .A(n490), .B(n2003), .Z(n2002) );
  XOR U1626 ( .A(n2004), .B(n2001), .Z(n2003) );
  XNOR U1627 ( .A(n1624), .B(n1997), .Z(n1999) );
  XOR U1628 ( .A(n2005), .B(n2006), .Z(n1624) );
  AND U1629 ( .A(n488), .B(n2007), .Z(n2006) );
  XOR U1630 ( .A(n2008), .B(n2005), .Z(n2007) );
  XOR U1631 ( .A(n2009), .B(n2010), .Z(n1997) );
  AND U1632 ( .A(n2011), .B(n2012), .Z(n2010) );
  XOR U1633 ( .A(n2009), .B(n1639), .Z(n2012) );
  XOR U1634 ( .A(n2013), .B(n2014), .Z(n1639) );
  AND U1635 ( .A(n490), .B(n2015), .Z(n2014) );
  XOR U1636 ( .A(n2016), .B(n2013), .Z(n2015) );
  XNOR U1637 ( .A(n1636), .B(n2009), .Z(n2011) );
  XOR U1638 ( .A(n2017), .B(n2018), .Z(n1636) );
  AND U1639 ( .A(n488), .B(n2019), .Z(n2018) );
  XOR U1640 ( .A(n2020), .B(n2017), .Z(n2019) );
  XOR U1641 ( .A(n2021), .B(n2022), .Z(n2009) );
  AND U1642 ( .A(n2023), .B(n2024), .Z(n2022) );
  XOR U1643 ( .A(n2021), .B(n1651), .Z(n2024) );
  XOR U1644 ( .A(n2025), .B(n2026), .Z(n1651) );
  AND U1645 ( .A(n490), .B(n2027), .Z(n2026) );
  XOR U1646 ( .A(n2028), .B(n2025), .Z(n2027) );
  XNOR U1647 ( .A(n1648), .B(n2021), .Z(n2023) );
  XOR U1648 ( .A(n2029), .B(n2030), .Z(n1648) );
  AND U1649 ( .A(n488), .B(n2031), .Z(n2030) );
  XOR U1650 ( .A(n2032), .B(n2029), .Z(n2031) );
  XOR U1651 ( .A(n2033), .B(n2034), .Z(n2021) );
  AND U1652 ( .A(n2035), .B(n2036), .Z(n2034) );
  XOR U1653 ( .A(n2033), .B(n1663), .Z(n2036) );
  XOR U1654 ( .A(n2037), .B(n2038), .Z(n1663) );
  AND U1655 ( .A(n490), .B(n2039), .Z(n2038) );
  XOR U1656 ( .A(n2040), .B(n2037), .Z(n2039) );
  XNOR U1657 ( .A(n1660), .B(n2033), .Z(n2035) );
  XOR U1658 ( .A(n2041), .B(n2042), .Z(n1660) );
  AND U1659 ( .A(n488), .B(n2043), .Z(n2042) );
  XOR U1660 ( .A(n2044), .B(n2041), .Z(n2043) );
  XOR U1661 ( .A(n2045), .B(n2046), .Z(n2033) );
  AND U1662 ( .A(n2047), .B(n2048), .Z(n2046) );
  XOR U1663 ( .A(n2045), .B(n1675), .Z(n2048) );
  XOR U1664 ( .A(n2049), .B(n2050), .Z(n1675) );
  AND U1665 ( .A(n490), .B(n2051), .Z(n2050) );
  XOR U1666 ( .A(n2052), .B(n2049), .Z(n2051) );
  XNOR U1667 ( .A(n1672), .B(n2045), .Z(n2047) );
  XOR U1668 ( .A(n2053), .B(n2054), .Z(n1672) );
  AND U1669 ( .A(n488), .B(n2055), .Z(n2054) );
  XOR U1670 ( .A(n2056), .B(n2053), .Z(n2055) );
  XOR U1671 ( .A(n2057), .B(n2058), .Z(n2045) );
  AND U1672 ( .A(n2059), .B(n2060), .Z(n2058) );
  XOR U1673 ( .A(n2057), .B(n1687), .Z(n2060) );
  XOR U1674 ( .A(n2061), .B(n2062), .Z(n1687) );
  AND U1675 ( .A(n490), .B(n2063), .Z(n2062) );
  XOR U1676 ( .A(n2064), .B(n2061), .Z(n2063) );
  XNOR U1677 ( .A(n1684), .B(n2057), .Z(n2059) );
  XOR U1678 ( .A(n2065), .B(n2066), .Z(n1684) );
  AND U1679 ( .A(n488), .B(n2067), .Z(n2066) );
  XOR U1680 ( .A(n2068), .B(n2065), .Z(n2067) );
  XOR U1681 ( .A(n2069), .B(n2070), .Z(n2057) );
  AND U1682 ( .A(n2071), .B(n2072), .Z(n2070) );
  XOR U1683 ( .A(n2069), .B(n1699), .Z(n2072) );
  XOR U1684 ( .A(n2073), .B(n2074), .Z(n1699) );
  AND U1685 ( .A(n490), .B(n2075), .Z(n2074) );
  XOR U1686 ( .A(n2076), .B(n2073), .Z(n2075) );
  XNOR U1687 ( .A(n1696), .B(n2069), .Z(n2071) );
  XOR U1688 ( .A(n2077), .B(n2078), .Z(n1696) );
  AND U1689 ( .A(n488), .B(n2079), .Z(n2078) );
  XOR U1690 ( .A(n2080), .B(n2077), .Z(n2079) );
  XOR U1691 ( .A(n2081), .B(n2082), .Z(n2069) );
  AND U1692 ( .A(n2083), .B(n2084), .Z(n2082) );
  XOR U1693 ( .A(n2081), .B(n1711), .Z(n2084) );
  XOR U1694 ( .A(n2085), .B(n2086), .Z(n1711) );
  AND U1695 ( .A(n490), .B(n2087), .Z(n2086) );
  XOR U1696 ( .A(n2088), .B(n2085), .Z(n2087) );
  XNOR U1697 ( .A(n1708), .B(n2081), .Z(n2083) );
  XOR U1698 ( .A(n2089), .B(n2090), .Z(n1708) );
  AND U1699 ( .A(n488), .B(n2091), .Z(n2090) );
  XOR U1700 ( .A(n2092), .B(n2089), .Z(n2091) );
  XOR U1701 ( .A(n2093), .B(n2094), .Z(n2081) );
  AND U1702 ( .A(n2095), .B(n2096), .Z(n2094) );
  XOR U1703 ( .A(n2093), .B(n1723), .Z(n2096) );
  XOR U1704 ( .A(n2097), .B(n2098), .Z(n1723) );
  AND U1705 ( .A(n490), .B(n2099), .Z(n2098) );
  XOR U1706 ( .A(n2100), .B(n2097), .Z(n2099) );
  XNOR U1707 ( .A(n1720), .B(n2093), .Z(n2095) );
  XOR U1708 ( .A(n2101), .B(n2102), .Z(n1720) );
  AND U1709 ( .A(n488), .B(n2103), .Z(n2102) );
  XOR U1710 ( .A(n2104), .B(n2101), .Z(n2103) );
  XOR U1711 ( .A(n2105), .B(n2106), .Z(n2093) );
  AND U1712 ( .A(n2107), .B(n2108), .Z(n2106) );
  XOR U1713 ( .A(n2105), .B(n1735), .Z(n2108) );
  XOR U1714 ( .A(n2109), .B(n2110), .Z(n1735) );
  AND U1715 ( .A(n490), .B(n2111), .Z(n2110) );
  XOR U1716 ( .A(n2112), .B(n2109), .Z(n2111) );
  XNOR U1717 ( .A(n1732), .B(n2105), .Z(n2107) );
  XOR U1718 ( .A(n2113), .B(n2114), .Z(n1732) );
  AND U1719 ( .A(n488), .B(n2115), .Z(n2114) );
  XOR U1720 ( .A(n2116), .B(n2113), .Z(n2115) );
  XOR U1721 ( .A(n2117), .B(n2118), .Z(n2105) );
  AND U1722 ( .A(n2119), .B(n2120), .Z(n2118) );
  XOR U1723 ( .A(n1747), .B(n2117), .Z(n2120) );
  XOR U1724 ( .A(n2121), .B(n2122), .Z(n1747) );
  AND U1725 ( .A(n490), .B(n2123), .Z(n2122) );
  XOR U1726 ( .A(n2121), .B(n2124), .Z(n2123) );
  XNOR U1727 ( .A(n2117), .B(n1744), .Z(n2119) );
  XOR U1728 ( .A(n2125), .B(n2126), .Z(n1744) );
  AND U1729 ( .A(n488), .B(n2127), .Z(n2126) );
  XOR U1730 ( .A(n2125), .B(n2128), .Z(n2127) );
  XOR U1731 ( .A(n2129), .B(n2130), .Z(n2117) );
  AND U1732 ( .A(n2131), .B(n2132), .Z(n2130) );
  XNOR U1733 ( .A(n2133), .B(n1760), .Z(n2132) );
  XOR U1734 ( .A(n2134), .B(n2135), .Z(n1760) );
  AND U1735 ( .A(n490), .B(n2136), .Z(n2135) );
  XOR U1736 ( .A(n2137), .B(n2134), .Z(n2136) );
  XNOR U1737 ( .A(n1757), .B(n2129), .Z(n2131) );
  XOR U1738 ( .A(n2138), .B(n2139), .Z(n1757) );
  AND U1739 ( .A(n488), .B(n2140), .Z(n2139) );
  XOR U1740 ( .A(n2141), .B(n2138), .Z(n2140) );
  IV U1741 ( .A(n2133), .Z(n2129) );
  AND U1742 ( .A(n1765), .B(n1768), .Z(n2133) );
  XNOR U1743 ( .A(n2142), .B(n2143), .Z(n1768) );
  AND U1744 ( .A(n490), .B(n2144), .Z(n2143) );
  XNOR U1745 ( .A(n2145), .B(n2142), .Z(n2144) );
  XOR U1746 ( .A(n2146), .B(n2147), .Z(n490) );
  AND U1747 ( .A(n2148), .B(n2149), .Z(n2147) );
  XOR U1748 ( .A(n2146), .B(n1776), .Z(n2149) );
  XNOR U1749 ( .A(n2150), .B(n2151), .Z(n1776) );
  AND U1750 ( .A(n2152), .B(n306), .Z(n2151) );
  AND U1751 ( .A(n2150), .B(n2153), .Z(n2152) );
  XNOR U1752 ( .A(n1773), .B(n2146), .Z(n2148) );
  XOR U1753 ( .A(n2154), .B(n2155), .Z(n1773) );
  AND U1754 ( .A(n2156), .B(n304), .Z(n2155) );
  NOR U1755 ( .A(n2154), .B(n2157), .Z(n2156) );
  XOR U1756 ( .A(n2158), .B(n2159), .Z(n2146) );
  AND U1757 ( .A(n2160), .B(n2161), .Z(n2159) );
  XOR U1758 ( .A(n2158), .B(n1788), .Z(n2161) );
  XOR U1759 ( .A(n2162), .B(n2163), .Z(n1788) );
  AND U1760 ( .A(n306), .B(n2164), .Z(n2163) );
  XOR U1761 ( .A(n2165), .B(n2162), .Z(n2164) );
  XNOR U1762 ( .A(n1785), .B(n2158), .Z(n2160) );
  XOR U1763 ( .A(n2166), .B(n2167), .Z(n1785) );
  AND U1764 ( .A(n304), .B(n2168), .Z(n2167) );
  XOR U1765 ( .A(n2169), .B(n2166), .Z(n2168) );
  XOR U1766 ( .A(n2170), .B(n2171), .Z(n2158) );
  AND U1767 ( .A(n2172), .B(n2173), .Z(n2171) );
  XOR U1768 ( .A(n2170), .B(n1800), .Z(n2173) );
  XOR U1769 ( .A(n2174), .B(n2175), .Z(n1800) );
  AND U1770 ( .A(n306), .B(n2176), .Z(n2175) );
  XOR U1771 ( .A(n2177), .B(n2174), .Z(n2176) );
  XNOR U1772 ( .A(n1797), .B(n2170), .Z(n2172) );
  XOR U1773 ( .A(n2178), .B(n2179), .Z(n1797) );
  AND U1774 ( .A(n304), .B(n2180), .Z(n2179) );
  XOR U1775 ( .A(n2181), .B(n2178), .Z(n2180) );
  XOR U1776 ( .A(n2182), .B(n2183), .Z(n2170) );
  AND U1777 ( .A(n2184), .B(n2185), .Z(n2183) );
  XOR U1778 ( .A(n2182), .B(n1812), .Z(n2185) );
  XOR U1779 ( .A(n2186), .B(n2187), .Z(n1812) );
  AND U1780 ( .A(n306), .B(n2188), .Z(n2187) );
  XOR U1781 ( .A(n2189), .B(n2186), .Z(n2188) );
  XNOR U1782 ( .A(n1809), .B(n2182), .Z(n2184) );
  XOR U1783 ( .A(n2190), .B(n2191), .Z(n1809) );
  AND U1784 ( .A(n304), .B(n2192), .Z(n2191) );
  XOR U1785 ( .A(n2193), .B(n2190), .Z(n2192) );
  XOR U1786 ( .A(n2194), .B(n2195), .Z(n2182) );
  AND U1787 ( .A(n2196), .B(n2197), .Z(n2195) );
  XOR U1788 ( .A(n2194), .B(n1824), .Z(n2197) );
  XOR U1789 ( .A(n2198), .B(n2199), .Z(n1824) );
  AND U1790 ( .A(n306), .B(n2200), .Z(n2199) );
  XOR U1791 ( .A(n2201), .B(n2198), .Z(n2200) );
  XNOR U1792 ( .A(n1821), .B(n2194), .Z(n2196) );
  XOR U1793 ( .A(n2202), .B(n2203), .Z(n1821) );
  AND U1794 ( .A(n304), .B(n2204), .Z(n2203) );
  XOR U1795 ( .A(n2205), .B(n2202), .Z(n2204) );
  XOR U1796 ( .A(n2206), .B(n2207), .Z(n2194) );
  AND U1797 ( .A(n2208), .B(n2209), .Z(n2207) );
  XOR U1798 ( .A(n2206), .B(n1836), .Z(n2209) );
  XOR U1799 ( .A(n2210), .B(n2211), .Z(n1836) );
  AND U1800 ( .A(n306), .B(n2212), .Z(n2211) );
  XOR U1801 ( .A(n2213), .B(n2210), .Z(n2212) );
  XNOR U1802 ( .A(n1833), .B(n2206), .Z(n2208) );
  XOR U1803 ( .A(n2214), .B(n2215), .Z(n1833) );
  AND U1804 ( .A(n304), .B(n2216), .Z(n2215) );
  XOR U1805 ( .A(n2217), .B(n2214), .Z(n2216) );
  XOR U1806 ( .A(n2218), .B(n2219), .Z(n2206) );
  AND U1807 ( .A(n2220), .B(n2221), .Z(n2219) );
  XOR U1808 ( .A(n2218), .B(n1848), .Z(n2221) );
  XOR U1809 ( .A(n2222), .B(n2223), .Z(n1848) );
  AND U1810 ( .A(n306), .B(n2224), .Z(n2223) );
  XOR U1811 ( .A(n2225), .B(n2222), .Z(n2224) );
  XNOR U1812 ( .A(n1845), .B(n2218), .Z(n2220) );
  XOR U1813 ( .A(n2226), .B(n2227), .Z(n1845) );
  AND U1814 ( .A(n304), .B(n2228), .Z(n2227) );
  XOR U1815 ( .A(n2229), .B(n2226), .Z(n2228) );
  XOR U1816 ( .A(n2230), .B(n2231), .Z(n2218) );
  AND U1817 ( .A(n2232), .B(n2233), .Z(n2231) );
  XOR U1818 ( .A(n2230), .B(n1860), .Z(n2233) );
  XOR U1819 ( .A(n2234), .B(n2235), .Z(n1860) );
  AND U1820 ( .A(n306), .B(n2236), .Z(n2235) );
  XOR U1821 ( .A(n2237), .B(n2234), .Z(n2236) );
  XNOR U1822 ( .A(n1857), .B(n2230), .Z(n2232) );
  XOR U1823 ( .A(n2238), .B(n2239), .Z(n1857) );
  AND U1824 ( .A(n304), .B(n2240), .Z(n2239) );
  XOR U1825 ( .A(n2241), .B(n2238), .Z(n2240) );
  XOR U1826 ( .A(n2242), .B(n2243), .Z(n2230) );
  AND U1827 ( .A(n2244), .B(n2245), .Z(n2243) );
  XOR U1828 ( .A(n2242), .B(n1872), .Z(n2245) );
  XOR U1829 ( .A(n2246), .B(n2247), .Z(n1872) );
  AND U1830 ( .A(n306), .B(n2248), .Z(n2247) );
  XOR U1831 ( .A(n2249), .B(n2246), .Z(n2248) );
  XNOR U1832 ( .A(n1869), .B(n2242), .Z(n2244) );
  XOR U1833 ( .A(n2250), .B(n2251), .Z(n1869) );
  AND U1834 ( .A(n304), .B(n2252), .Z(n2251) );
  XOR U1835 ( .A(n2253), .B(n2250), .Z(n2252) );
  XOR U1836 ( .A(n2254), .B(n2255), .Z(n2242) );
  AND U1837 ( .A(n2256), .B(n2257), .Z(n2255) );
  XOR U1838 ( .A(n2254), .B(n1884), .Z(n2257) );
  XOR U1839 ( .A(n2258), .B(n2259), .Z(n1884) );
  AND U1840 ( .A(n306), .B(n2260), .Z(n2259) );
  XOR U1841 ( .A(n2261), .B(n2258), .Z(n2260) );
  XNOR U1842 ( .A(n1881), .B(n2254), .Z(n2256) );
  XOR U1843 ( .A(n2262), .B(n2263), .Z(n1881) );
  AND U1844 ( .A(n304), .B(n2264), .Z(n2263) );
  XOR U1845 ( .A(n2265), .B(n2262), .Z(n2264) );
  XOR U1846 ( .A(n2266), .B(n2267), .Z(n2254) );
  AND U1847 ( .A(n2268), .B(n2269), .Z(n2267) );
  XOR U1848 ( .A(n2266), .B(n1896), .Z(n2269) );
  XOR U1849 ( .A(n2270), .B(n2271), .Z(n1896) );
  AND U1850 ( .A(n306), .B(n2272), .Z(n2271) );
  XOR U1851 ( .A(n2273), .B(n2270), .Z(n2272) );
  XNOR U1852 ( .A(n1893), .B(n2266), .Z(n2268) );
  XOR U1853 ( .A(n2274), .B(n2275), .Z(n1893) );
  AND U1854 ( .A(n304), .B(n2276), .Z(n2275) );
  XOR U1855 ( .A(n2277), .B(n2274), .Z(n2276) );
  XOR U1856 ( .A(n2278), .B(n2279), .Z(n2266) );
  AND U1857 ( .A(n2280), .B(n2281), .Z(n2279) );
  XOR U1858 ( .A(n2278), .B(n1908), .Z(n2281) );
  XOR U1859 ( .A(n2282), .B(n2283), .Z(n1908) );
  AND U1860 ( .A(n306), .B(n2284), .Z(n2283) );
  XOR U1861 ( .A(n2285), .B(n2282), .Z(n2284) );
  XNOR U1862 ( .A(n1905), .B(n2278), .Z(n2280) );
  XOR U1863 ( .A(n2286), .B(n2287), .Z(n1905) );
  AND U1864 ( .A(n304), .B(n2288), .Z(n2287) );
  XOR U1865 ( .A(n2289), .B(n2286), .Z(n2288) );
  XOR U1866 ( .A(n2290), .B(n2291), .Z(n2278) );
  AND U1867 ( .A(n2292), .B(n2293), .Z(n2291) );
  XOR U1868 ( .A(n2290), .B(n1920), .Z(n2293) );
  XOR U1869 ( .A(n2294), .B(n2295), .Z(n1920) );
  AND U1870 ( .A(n306), .B(n2296), .Z(n2295) );
  XOR U1871 ( .A(n2297), .B(n2294), .Z(n2296) );
  XNOR U1872 ( .A(n1917), .B(n2290), .Z(n2292) );
  XOR U1873 ( .A(n2298), .B(n2299), .Z(n1917) );
  AND U1874 ( .A(n304), .B(n2300), .Z(n2299) );
  XOR U1875 ( .A(n2301), .B(n2298), .Z(n2300) );
  XOR U1876 ( .A(n2302), .B(n2303), .Z(n2290) );
  AND U1877 ( .A(n2304), .B(n2305), .Z(n2303) );
  XOR U1878 ( .A(n2302), .B(n1932), .Z(n2305) );
  XOR U1879 ( .A(n2306), .B(n2307), .Z(n1932) );
  AND U1880 ( .A(n306), .B(n2308), .Z(n2307) );
  XOR U1881 ( .A(n2309), .B(n2306), .Z(n2308) );
  XNOR U1882 ( .A(n1929), .B(n2302), .Z(n2304) );
  XOR U1883 ( .A(n2310), .B(n2311), .Z(n1929) );
  AND U1884 ( .A(n304), .B(n2312), .Z(n2311) );
  XOR U1885 ( .A(n2313), .B(n2310), .Z(n2312) );
  XOR U1886 ( .A(n2314), .B(n2315), .Z(n2302) );
  AND U1887 ( .A(n2316), .B(n2317), .Z(n2315) );
  XOR U1888 ( .A(n2314), .B(n1944), .Z(n2317) );
  XOR U1889 ( .A(n2318), .B(n2319), .Z(n1944) );
  AND U1890 ( .A(n306), .B(n2320), .Z(n2319) );
  XOR U1891 ( .A(n2321), .B(n2318), .Z(n2320) );
  XNOR U1892 ( .A(n1941), .B(n2314), .Z(n2316) );
  XOR U1893 ( .A(n2322), .B(n2323), .Z(n1941) );
  AND U1894 ( .A(n304), .B(n2324), .Z(n2323) );
  XOR U1895 ( .A(n2325), .B(n2322), .Z(n2324) );
  XOR U1896 ( .A(n2326), .B(n2327), .Z(n2314) );
  AND U1897 ( .A(n2328), .B(n2329), .Z(n2327) );
  XOR U1898 ( .A(n2326), .B(n1956), .Z(n2329) );
  XOR U1899 ( .A(n2330), .B(n2331), .Z(n1956) );
  AND U1900 ( .A(n306), .B(n2332), .Z(n2331) );
  XOR U1901 ( .A(n2333), .B(n2330), .Z(n2332) );
  XNOR U1902 ( .A(n1953), .B(n2326), .Z(n2328) );
  XOR U1903 ( .A(n2334), .B(n2335), .Z(n1953) );
  AND U1904 ( .A(n304), .B(n2336), .Z(n2335) );
  XOR U1905 ( .A(n2337), .B(n2334), .Z(n2336) );
  XOR U1906 ( .A(n2338), .B(n2339), .Z(n2326) );
  AND U1907 ( .A(n2340), .B(n2341), .Z(n2339) );
  XOR U1908 ( .A(n2338), .B(n1968), .Z(n2341) );
  XOR U1909 ( .A(n2342), .B(n2343), .Z(n1968) );
  AND U1910 ( .A(n306), .B(n2344), .Z(n2343) );
  XOR U1911 ( .A(n2345), .B(n2342), .Z(n2344) );
  XNOR U1912 ( .A(n1965), .B(n2338), .Z(n2340) );
  XOR U1913 ( .A(n2346), .B(n2347), .Z(n1965) );
  AND U1914 ( .A(n304), .B(n2348), .Z(n2347) );
  XOR U1915 ( .A(n2349), .B(n2346), .Z(n2348) );
  XOR U1916 ( .A(n2350), .B(n2351), .Z(n2338) );
  AND U1917 ( .A(n2352), .B(n2353), .Z(n2351) );
  XOR U1918 ( .A(n2350), .B(n1980), .Z(n2353) );
  XOR U1919 ( .A(n2354), .B(n2355), .Z(n1980) );
  AND U1920 ( .A(n306), .B(n2356), .Z(n2355) );
  XOR U1921 ( .A(n2357), .B(n2354), .Z(n2356) );
  XNOR U1922 ( .A(n1977), .B(n2350), .Z(n2352) );
  XOR U1923 ( .A(n2358), .B(n2359), .Z(n1977) );
  AND U1924 ( .A(n304), .B(n2360), .Z(n2359) );
  XOR U1925 ( .A(n2361), .B(n2358), .Z(n2360) );
  XOR U1926 ( .A(n2362), .B(n2363), .Z(n2350) );
  AND U1927 ( .A(n2364), .B(n2365), .Z(n2363) );
  XOR U1928 ( .A(n2362), .B(n1992), .Z(n2365) );
  XOR U1929 ( .A(n2366), .B(n2367), .Z(n1992) );
  AND U1930 ( .A(n306), .B(n2368), .Z(n2367) );
  XOR U1931 ( .A(n2369), .B(n2366), .Z(n2368) );
  XNOR U1932 ( .A(n1989), .B(n2362), .Z(n2364) );
  XOR U1933 ( .A(n2370), .B(n2371), .Z(n1989) );
  AND U1934 ( .A(n304), .B(n2372), .Z(n2371) );
  XOR U1935 ( .A(n2373), .B(n2370), .Z(n2372) );
  XOR U1936 ( .A(n2374), .B(n2375), .Z(n2362) );
  AND U1937 ( .A(n2376), .B(n2377), .Z(n2375) );
  XOR U1938 ( .A(n2374), .B(n2004), .Z(n2377) );
  XOR U1939 ( .A(n2378), .B(n2379), .Z(n2004) );
  AND U1940 ( .A(n306), .B(n2380), .Z(n2379) );
  XOR U1941 ( .A(n2381), .B(n2378), .Z(n2380) );
  XNOR U1942 ( .A(n2001), .B(n2374), .Z(n2376) );
  XOR U1943 ( .A(n2382), .B(n2383), .Z(n2001) );
  AND U1944 ( .A(n304), .B(n2384), .Z(n2383) );
  XOR U1945 ( .A(n2385), .B(n2382), .Z(n2384) );
  XOR U1946 ( .A(n2386), .B(n2387), .Z(n2374) );
  AND U1947 ( .A(n2388), .B(n2389), .Z(n2387) );
  XOR U1948 ( .A(n2386), .B(n2016), .Z(n2389) );
  XOR U1949 ( .A(n2390), .B(n2391), .Z(n2016) );
  AND U1950 ( .A(n306), .B(n2392), .Z(n2391) );
  XOR U1951 ( .A(n2393), .B(n2390), .Z(n2392) );
  XNOR U1952 ( .A(n2013), .B(n2386), .Z(n2388) );
  XOR U1953 ( .A(n2394), .B(n2395), .Z(n2013) );
  AND U1954 ( .A(n304), .B(n2396), .Z(n2395) );
  XOR U1955 ( .A(n2397), .B(n2394), .Z(n2396) );
  XOR U1956 ( .A(n2398), .B(n2399), .Z(n2386) );
  AND U1957 ( .A(n2400), .B(n2401), .Z(n2399) );
  XOR U1958 ( .A(n2398), .B(n2028), .Z(n2401) );
  XOR U1959 ( .A(n2402), .B(n2403), .Z(n2028) );
  AND U1960 ( .A(n306), .B(n2404), .Z(n2403) );
  XOR U1961 ( .A(n2405), .B(n2402), .Z(n2404) );
  XNOR U1962 ( .A(n2025), .B(n2398), .Z(n2400) );
  XOR U1963 ( .A(n2406), .B(n2407), .Z(n2025) );
  AND U1964 ( .A(n304), .B(n2408), .Z(n2407) );
  XOR U1965 ( .A(n2409), .B(n2406), .Z(n2408) );
  XOR U1966 ( .A(n2410), .B(n2411), .Z(n2398) );
  AND U1967 ( .A(n2412), .B(n2413), .Z(n2411) );
  XOR U1968 ( .A(n2410), .B(n2040), .Z(n2413) );
  XOR U1969 ( .A(n2414), .B(n2415), .Z(n2040) );
  AND U1970 ( .A(n306), .B(n2416), .Z(n2415) );
  XOR U1971 ( .A(n2417), .B(n2414), .Z(n2416) );
  XNOR U1972 ( .A(n2037), .B(n2410), .Z(n2412) );
  XOR U1973 ( .A(n2418), .B(n2419), .Z(n2037) );
  AND U1974 ( .A(n304), .B(n2420), .Z(n2419) );
  XOR U1975 ( .A(n2421), .B(n2418), .Z(n2420) );
  XOR U1976 ( .A(n2422), .B(n2423), .Z(n2410) );
  AND U1977 ( .A(n2424), .B(n2425), .Z(n2423) );
  XOR U1978 ( .A(n2422), .B(n2052), .Z(n2425) );
  XOR U1979 ( .A(n2426), .B(n2427), .Z(n2052) );
  AND U1980 ( .A(n306), .B(n2428), .Z(n2427) );
  XOR U1981 ( .A(n2429), .B(n2426), .Z(n2428) );
  XNOR U1982 ( .A(n2049), .B(n2422), .Z(n2424) );
  XOR U1983 ( .A(n2430), .B(n2431), .Z(n2049) );
  AND U1984 ( .A(n304), .B(n2432), .Z(n2431) );
  XOR U1985 ( .A(n2433), .B(n2430), .Z(n2432) );
  XOR U1986 ( .A(n2434), .B(n2435), .Z(n2422) );
  AND U1987 ( .A(n2436), .B(n2437), .Z(n2435) );
  XOR U1988 ( .A(n2434), .B(n2064), .Z(n2437) );
  XOR U1989 ( .A(n2438), .B(n2439), .Z(n2064) );
  AND U1990 ( .A(n306), .B(n2440), .Z(n2439) );
  XOR U1991 ( .A(n2441), .B(n2438), .Z(n2440) );
  XNOR U1992 ( .A(n2061), .B(n2434), .Z(n2436) );
  XOR U1993 ( .A(n2442), .B(n2443), .Z(n2061) );
  AND U1994 ( .A(n304), .B(n2444), .Z(n2443) );
  XOR U1995 ( .A(n2445), .B(n2442), .Z(n2444) );
  XOR U1996 ( .A(n2446), .B(n2447), .Z(n2434) );
  AND U1997 ( .A(n2448), .B(n2449), .Z(n2447) );
  XOR U1998 ( .A(n2446), .B(n2076), .Z(n2449) );
  XOR U1999 ( .A(n2450), .B(n2451), .Z(n2076) );
  AND U2000 ( .A(n306), .B(n2452), .Z(n2451) );
  XOR U2001 ( .A(n2453), .B(n2450), .Z(n2452) );
  XNOR U2002 ( .A(n2073), .B(n2446), .Z(n2448) );
  XOR U2003 ( .A(n2454), .B(n2455), .Z(n2073) );
  AND U2004 ( .A(n304), .B(n2456), .Z(n2455) );
  XOR U2005 ( .A(n2457), .B(n2454), .Z(n2456) );
  XOR U2006 ( .A(n2458), .B(n2459), .Z(n2446) );
  AND U2007 ( .A(n2460), .B(n2461), .Z(n2459) );
  XOR U2008 ( .A(n2458), .B(n2088), .Z(n2461) );
  XOR U2009 ( .A(n2462), .B(n2463), .Z(n2088) );
  AND U2010 ( .A(n306), .B(n2464), .Z(n2463) );
  XOR U2011 ( .A(n2465), .B(n2462), .Z(n2464) );
  XNOR U2012 ( .A(n2085), .B(n2458), .Z(n2460) );
  XOR U2013 ( .A(n2466), .B(n2467), .Z(n2085) );
  AND U2014 ( .A(n304), .B(n2468), .Z(n2467) );
  XOR U2015 ( .A(n2469), .B(n2466), .Z(n2468) );
  XOR U2016 ( .A(n2470), .B(n2471), .Z(n2458) );
  AND U2017 ( .A(n2472), .B(n2473), .Z(n2471) );
  XOR U2018 ( .A(n2470), .B(n2100), .Z(n2473) );
  XOR U2019 ( .A(n2474), .B(n2475), .Z(n2100) );
  AND U2020 ( .A(n306), .B(n2476), .Z(n2475) );
  XOR U2021 ( .A(n2477), .B(n2474), .Z(n2476) );
  XNOR U2022 ( .A(n2097), .B(n2470), .Z(n2472) );
  XOR U2023 ( .A(n2478), .B(n2479), .Z(n2097) );
  AND U2024 ( .A(n304), .B(n2480), .Z(n2479) );
  XOR U2025 ( .A(n2481), .B(n2478), .Z(n2480) );
  XOR U2026 ( .A(n2482), .B(n2483), .Z(n2470) );
  AND U2027 ( .A(n2484), .B(n2485), .Z(n2483) );
  XOR U2028 ( .A(n2482), .B(n2112), .Z(n2485) );
  XOR U2029 ( .A(n2486), .B(n2487), .Z(n2112) );
  AND U2030 ( .A(n306), .B(n2488), .Z(n2487) );
  XOR U2031 ( .A(n2489), .B(n2486), .Z(n2488) );
  XNOR U2032 ( .A(n2109), .B(n2482), .Z(n2484) );
  XOR U2033 ( .A(n2490), .B(n2491), .Z(n2109) );
  AND U2034 ( .A(n304), .B(n2492), .Z(n2491) );
  XOR U2035 ( .A(n2493), .B(n2490), .Z(n2492) );
  XOR U2036 ( .A(n2494), .B(n2495), .Z(n2482) );
  AND U2037 ( .A(n2496), .B(n2497), .Z(n2495) );
  XOR U2038 ( .A(n2124), .B(n2494), .Z(n2497) );
  XOR U2039 ( .A(n2498), .B(n2499), .Z(n2124) );
  AND U2040 ( .A(n306), .B(n2500), .Z(n2499) );
  XOR U2041 ( .A(n2498), .B(n2501), .Z(n2500) );
  XNOR U2042 ( .A(n2494), .B(n2121), .Z(n2496) );
  XOR U2043 ( .A(n2502), .B(n2503), .Z(n2121) );
  AND U2044 ( .A(n304), .B(n2504), .Z(n2503) );
  XOR U2045 ( .A(n2502), .B(n2505), .Z(n2504) );
  XOR U2046 ( .A(n2506), .B(n2507), .Z(n2494) );
  AND U2047 ( .A(n2508), .B(n2509), .Z(n2507) );
  XNOR U2048 ( .A(n2510), .B(n2137), .Z(n2509) );
  XOR U2049 ( .A(n2511), .B(n2512), .Z(n2137) );
  AND U2050 ( .A(n306), .B(n2513), .Z(n2512) );
  XOR U2051 ( .A(n2514), .B(n2511), .Z(n2513) );
  XNOR U2052 ( .A(n2134), .B(n2506), .Z(n2508) );
  XOR U2053 ( .A(n2515), .B(n2516), .Z(n2134) );
  AND U2054 ( .A(n304), .B(n2517), .Z(n2516) );
  XOR U2055 ( .A(n2518), .B(n2515), .Z(n2517) );
  IV U2056 ( .A(n2510), .Z(n2506) );
  AND U2057 ( .A(n2142), .B(n2145), .Z(n2510) );
  XNOR U2058 ( .A(n2519), .B(n2520), .Z(n2145) );
  AND U2059 ( .A(n306), .B(n2521), .Z(n2520) );
  XNOR U2060 ( .A(n2522), .B(n2519), .Z(n2521) );
  XOR U2061 ( .A(n2523), .B(n2524), .Z(n306) );
  AND U2062 ( .A(n2525), .B(n2526), .Z(n2524) );
  XOR U2063 ( .A(n2153), .B(n2523), .Z(n2526) );
  IV U2064 ( .A(n2527), .Z(n2153) );
  AND U2065 ( .A(p_input[4095]), .B(p_input[4063]), .Z(n2527) );
  XOR U2066 ( .A(n2523), .B(n2150), .Z(n2525) );
  AND U2067 ( .A(p_input[3999]), .B(p_input[4031]), .Z(n2150) );
  XOR U2068 ( .A(n2528), .B(n2529), .Z(n2523) );
  AND U2069 ( .A(n2530), .B(n2531), .Z(n2529) );
  XOR U2070 ( .A(n2528), .B(n2165), .Z(n2531) );
  XNOR U2071 ( .A(p_input[4062]), .B(n2532), .Z(n2165) );
  AND U2072 ( .A(n182), .B(n2533), .Z(n2532) );
  XOR U2073 ( .A(p_input[4094]), .B(p_input[4062]), .Z(n2533) );
  XNOR U2074 ( .A(n2162), .B(n2528), .Z(n2530) );
  XOR U2075 ( .A(n2534), .B(n2535), .Z(n2162) );
  AND U2076 ( .A(n180), .B(n2536), .Z(n2535) );
  XOR U2077 ( .A(p_input[4030]), .B(p_input[3998]), .Z(n2536) );
  XOR U2078 ( .A(n2537), .B(n2538), .Z(n2528) );
  AND U2079 ( .A(n2539), .B(n2540), .Z(n2538) );
  XOR U2080 ( .A(n2537), .B(n2177), .Z(n2540) );
  XNOR U2081 ( .A(p_input[4061]), .B(n2541), .Z(n2177) );
  AND U2082 ( .A(n182), .B(n2542), .Z(n2541) );
  XOR U2083 ( .A(p_input[4093]), .B(p_input[4061]), .Z(n2542) );
  XNOR U2084 ( .A(n2174), .B(n2537), .Z(n2539) );
  XOR U2085 ( .A(n2543), .B(n2544), .Z(n2174) );
  AND U2086 ( .A(n180), .B(n2545), .Z(n2544) );
  XOR U2087 ( .A(p_input[4029]), .B(p_input[3997]), .Z(n2545) );
  XOR U2088 ( .A(n2546), .B(n2547), .Z(n2537) );
  AND U2089 ( .A(n2548), .B(n2549), .Z(n2547) );
  XOR U2090 ( .A(n2546), .B(n2189), .Z(n2549) );
  XNOR U2091 ( .A(p_input[4060]), .B(n2550), .Z(n2189) );
  AND U2092 ( .A(n182), .B(n2551), .Z(n2550) );
  XOR U2093 ( .A(p_input[4092]), .B(p_input[4060]), .Z(n2551) );
  XNOR U2094 ( .A(n2186), .B(n2546), .Z(n2548) );
  XOR U2095 ( .A(n2552), .B(n2553), .Z(n2186) );
  AND U2096 ( .A(n180), .B(n2554), .Z(n2553) );
  XOR U2097 ( .A(p_input[4028]), .B(p_input[3996]), .Z(n2554) );
  XOR U2098 ( .A(n2555), .B(n2556), .Z(n2546) );
  AND U2099 ( .A(n2557), .B(n2558), .Z(n2556) );
  XOR U2100 ( .A(n2555), .B(n2201), .Z(n2558) );
  XNOR U2101 ( .A(p_input[4059]), .B(n2559), .Z(n2201) );
  AND U2102 ( .A(n182), .B(n2560), .Z(n2559) );
  XOR U2103 ( .A(p_input[4091]), .B(p_input[4059]), .Z(n2560) );
  XNOR U2104 ( .A(n2198), .B(n2555), .Z(n2557) );
  XOR U2105 ( .A(n2561), .B(n2562), .Z(n2198) );
  AND U2106 ( .A(n180), .B(n2563), .Z(n2562) );
  XOR U2107 ( .A(p_input[4027]), .B(p_input[3995]), .Z(n2563) );
  XOR U2108 ( .A(n2564), .B(n2565), .Z(n2555) );
  AND U2109 ( .A(n2566), .B(n2567), .Z(n2565) );
  XOR U2110 ( .A(n2564), .B(n2213), .Z(n2567) );
  XNOR U2111 ( .A(p_input[4058]), .B(n2568), .Z(n2213) );
  AND U2112 ( .A(n182), .B(n2569), .Z(n2568) );
  XOR U2113 ( .A(p_input[4090]), .B(p_input[4058]), .Z(n2569) );
  XNOR U2114 ( .A(n2210), .B(n2564), .Z(n2566) );
  XOR U2115 ( .A(n2570), .B(n2571), .Z(n2210) );
  AND U2116 ( .A(n180), .B(n2572), .Z(n2571) );
  XOR U2117 ( .A(p_input[4026]), .B(p_input[3994]), .Z(n2572) );
  XOR U2118 ( .A(n2573), .B(n2574), .Z(n2564) );
  AND U2119 ( .A(n2575), .B(n2576), .Z(n2574) );
  XOR U2120 ( .A(n2573), .B(n2225), .Z(n2576) );
  XNOR U2121 ( .A(p_input[4057]), .B(n2577), .Z(n2225) );
  AND U2122 ( .A(n182), .B(n2578), .Z(n2577) );
  XOR U2123 ( .A(p_input[4089]), .B(p_input[4057]), .Z(n2578) );
  XNOR U2124 ( .A(n2222), .B(n2573), .Z(n2575) );
  XOR U2125 ( .A(n2579), .B(n2580), .Z(n2222) );
  AND U2126 ( .A(n180), .B(n2581), .Z(n2580) );
  XOR U2127 ( .A(p_input[4025]), .B(p_input[3993]), .Z(n2581) );
  XOR U2128 ( .A(n2582), .B(n2583), .Z(n2573) );
  AND U2129 ( .A(n2584), .B(n2585), .Z(n2583) );
  XOR U2130 ( .A(n2582), .B(n2237), .Z(n2585) );
  XNOR U2131 ( .A(p_input[4056]), .B(n2586), .Z(n2237) );
  AND U2132 ( .A(n182), .B(n2587), .Z(n2586) );
  XOR U2133 ( .A(p_input[4088]), .B(p_input[4056]), .Z(n2587) );
  XNOR U2134 ( .A(n2234), .B(n2582), .Z(n2584) );
  XOR U2135 ( .A(n2588), .B(n2589), .Z(n2234) );
  AND U2136 ( .A(n180), .B(n2590), .Z(n2589) );
  XOR U2137 ( .A(p_input[4024]), .B(p_input[3992]), .Z(n2590) );
  XOR U2138 ( .A(n2591), .B(n2592), .Z(n2582) );
  AND U2139 ( .A(n2593), .B(n2594), .Z(n2592) );
  XOR U2140 ( .A(n2591), .B(n2249), .Z(n2594) );
  XNOR U2141 ( .A(p_input[4055]), .B(n2595), .Z(n2249) );
  AND U2142 ( .A(n182), .B(n2596), .Z(n2595) );
  XOR U2143 ( .A(p_input[4087]), .B(p_input[4055]), .Z(n2596) );
  XNOR U2144 ( .A(n2246), .B(n2591), .Z(n2593) );
  XOR U2145 ( .A(n2597), .B(n2598), .Z(n2246) );
  AND U2146 ( .A(n180), .B(n2599), .Z(n2598) );
  XOR U2147 ( .A(p_input[4023]), .B(p_input[3991]), .Z(n2599) );
  XOR U2148 ( .A(n2600), .B(n2601), .Z(n2591) );
  AND U2149 ( .A(n2602), .B(n2603), .Z(n2601) );
  XOR U2150 ( .A(n2600), .B(n2261), .Z(n2603) );
  XNOR U2151 ( .A(p_input[4054]), .B(n2604), .Z(n2261) );
  AND U2152 ( .A(n182), .B(n2605), .Z(n2604) );
  XOR U2153 ( .A(p_input[4086]), .B(p_input[4054]), .Z(n2605) );
  XNOR U2154 ( .A(n2258), .B(n2600), .Z(n2602) );
  XOR U2155 ( .A(n2606), .B(n2607), .Z(n2258) );
  AND U2156 ( .A(n180), .B(n2608), .Z(n2607) );
  XOR U2157 ( .A(p_input[4022]), .B(p_input[3990]), .Z(n2608) );
  XOR U2158 ( .A(n2609), .B(n2610), .Z(n2600) );
  AND U2159 ( .A(n2611), .B(n2612), .Z(n2610) );
  XOR U2160 ( .A(n2609), .B(n2273), .Z(n2612) );
  XNOR U2161 ( .A(p_input[4053]), .B(n2613), .Z(n2273) );
  AND U2162 ( .A(n182), .B(n2614), .Z(n2613) );
  XOR U2163 ( .A(p_input[4085]), .B(p_input[4053]), .Z(n2614) );
  XNOR U2164 ( .A(n2270), .B(n2609), .Z(n2611) );
  XOR U2165 ( .A(n2615), .B(n2616), .Z(n2270) );
  AND U2166 ( .A(n180), .B(n2617), .Z(n2616) );
  XOR U2167 ( .A(p_input[4021]), .B(p_input[3989]), .Z(n2617) );
  XOR U2168 ( .A(n2618), .B(n2619), .Z(n2609) );
  AND U2169 ( .A(n2620), .B(n2621), .Z(n2619) );
  XOR U2170 ( .A(n2618), .B(n2285), .Z(n2621) );
  XNOR U2171 ( .A(p_input[4052]), .B(n2622), .Z(n2285) );
  AND U2172 ( .A(n182), .B(n2623), .Z(n2622) );
  XOR U2173 ( .A(p_input[4084]), .B(p_input[4052]), .Z(n2623) );
  XNOR U2174 ( .A(n2282), .B(n2618), .Z(n2620) );
  XOR U2175 ( .A(n2624), .B(n2625), .Z(n2282) );
  AND U2176 ( .A(n180), .B(n2626), .Z(n2625) );
  XOR U2177 ( .A(p_input[4020]), .B(p_input[3988]), .Z(n2626) );
  XOR U2178 ( .A(n2627), .B(n2628), .Z(n2618) );
  AND U2179 ( .A(n2629), .B(n2630), .Z(n2628) );
  XOR U2180 ( .A(n2627), .B(n2297), .Z(n2630) );
  XNOR U2181 ( .A(p_input[4051]), .B(n2631), .Z(n2297) );
  AND U2182 ( .A(n182), .B(n2632), .Z(n2631) );
  XOR U2183 ( .A(p_input[4083]), .B(p_input[4051]), .Z(n2632) );
  XNOR U2184 ( .A(n2294), .B(n2627), .Z(n2629) );
  XOR U2185 ( .A(n2633), .B(n2634), .Z(n2294) );
  AND U2186 ( .A(n180), .B(n2635), .Z(n2634) );
  XOR U2187 ( .A(p_input[4019]), .B(p_input[3987]), .Z(n2635) );
  XOR U2188 ( .A(n2636), .B(n2637), .Z(n2627) );
  AND U2189 ( .A(n2638), .B(n2639), .Z(n2637) );
  XOR U2190 ( .A(n2636), .B(n2309), .Z(n2639) );
  XNOR U2191 ( .A(p_input[4050]), .B(n2640), .Z(n2309) );
  AND U2192 ( .A(n182), .B(n2641), .Z(n2640) );
  XOR U2193 ( .A(p_input[4082]), .B(p_input[4050]), .Z(n2641) );
  XNOR U2194 ( .A(n2306), .B(n2636), .Z(n2638) );
  XOR U2195 ( .A(n2642), .B(n2643), .Z(n2306) );
  AND U2196 ( .A(n180), .B(n2644), .Z(n2643) );
  XOR U2197 ( .A(p_input[4018]), .B(p_input[3986]), .Z(n2644) );
  XOR U2198 ( .A(n2645), .B(n2646), .Z(n2636) );
  AND U2199 ( .A(n2647), .B(n2648), .Z(n2646) );
  XOR U2200 ( .A(n2645), .B(n2321), .Z(n2648) );
  XNOR U2201 ( .A(p_input[4049]), .B(n2649), .Z(n2321) );
  AND U2202 ( .A(n182), .B(n2650), .Z(n2649) );
  XOR U2203 ( .A(p_input[4081]), .B(p_input[4049]), .Z(n2650) );
  XNOR U2204 ( .A(n2318), .B(n2645), .Z(n2647) );
  XOR U2205 ( .A(n2651), .B(n2652), .Z(n2318) );
  AND U2206 ( .A(n180), .B(n2653), .Z(n2652) );
  XOR U2207 ( .A(p_input[4017]), .B(p_input[3985]), .Z(n2653) );
  XOR U2208 ( .A(n2654), .B(n2655), .Z(n2645) );
  AND U2209 ( .A(n2656), .B(n2657), .Z(n2655) );
  XOR U2210 ( .A(n2654), .B(n2333), .Z(n2657) );
  XNOR U2211 ( .A(p_input[4048]), .B(n2658), .Z(n2333) );
  AND U2212 ( .A(n182), .B(n2659), .Z(n2658) );
  XOR U2213 ( .A(p_input[4080]), .B(p_input[4048]), .Z(n2659) );
  XNOR U2214 ( .A(n2330), .B(n2654), .Z(n2656) );
  XOR U2215 ( .A(n2660), .B(n2661), .Z(n2330) );
  AND U2216 ( .A(n180), .B(n2662), .Z(n2661) );
  XOR U2217 ( .A(p_input[4016]), .B(p_input[3984]), .Z(n2662) );
  XOR U2218 ( .A(n2663), .B(n2664), .Z(n2654) );
  AND U2219 ( .A(n2665), .B(n2666), .Z(n2664) );
  XOR U2220 ( .A(n2663), .B(n2345), .Z(n2666) );
  XNOR U2221 ( .A(p_input[4047]), .B(n2667), .Z(n2345) );
  AND U2222 ( .A(n182), .B(n2668), .Z(n2667) );
  XOR U2223 ( .A(p_input[4079]), .B(p_input[4047]), .Z(n2668) );
  XNOR U2224 ( .A(n2342), .B(n2663), .Z(n2665) );
  XOR U2225 ( .A(n2669), .B(n2670), .Z(n2342) );
  AND U2226 ( .A(n180), .B(n2671), .Z(n2670) );
  XOR U2227 ( .A(p_input[4015]), .B(p_input[3983]), .Z(n2671) );
  XOR U2228 ( .A(n2672), .B(n2673), .Z(n2663) );
  AND U2229 ( .A(n2674), .B(n2675), .Z(n2673) );
  XOR U2230 ( .A(n2672), .B(n2357), .Z(n2675) );
  XNOR U2231 ( .A(p_input[4046]), .B(n2676), .Z(n2357) );
  AND U2232 ( .A(n182), .B(n2677), .Z(n2676) );
  XOR U2233 ( .A(p_input[4078]), .B(p_input[4046]), .Z(n2677) );
  XNOR U2234 ( .A(n2354), .B(n2672), .Z(n2674) );
  XOR U2235 ( .A(n2678), .B(n2679), .Z(n2354) );
  AND U2236 ( .A(n180), .B(n2680), .Z(n2679) );
  XOR U2237 ( .A(p_input[4014]), .B(p_input[3982]), .Z(n2680) );
  XOR U2238 ( .A(n2681), .B(n2682), .Z(n2672) );
  AND U2239 ( .A(n2683), .B(n2684), .Z(n2682) );
  XOR U2240 ( .A(n2681), .B(n2369), .Z(n2684) );
  XNOR U2241 ( .A(p_input[4045]), .B(n2685), .Z(n2369) );
  AND U2242 ( .A(n182), .B(n2686), .Z(n2685) );
  XOR U2243 ( .A(p_input[4077]), .B(p_input[4045]), .Z(n2686) );
  XNOR U2244 ( .A(n2366), .B(n2681), .Z(n2683) );
  XOR U2245 ( .A(n2687), .B(n2688), .Z(n2366) );
  AND U2246 ( .A(n180), .B(n2689), .Z(n2688) );
  XOR U2247 ( .A(p_input[4013]), .B(p_input[3981]), .Z(n2689) );
  XOR U2248 ( .A(n2690), .B(n2691), .Z(n2681) );
  AND U2249 ( .A(n2692), .B(n2693), .Z(n2691) );
  XOR U2250 ( .A(n2690), .B(n2381), .Z(n2693) );
  XNOR U2251 ( .A(p_input[4044]), .B(n2694), .Z(n2381) );
  AND U2252 ( .A(n182), .B(n2695), .Z(n2694) );
  XOR U2253 ( .A(p_input[4076]), .B(p_input[4044]), .Z(n2695) );
  XNOR U2254 ( .A(n2378), .B(n2690), .Z(n2692) );
  XOR U2255 ( .A(n2696), .B(n2697), .Z(n2378) );
  AND U2256 ( .A(n180), .B(n2698), .Z(n2697) );
  XOR U2257 ( .A(p_input[4012]), .B(p_input[3980]), .Z(n2698) );
  XOR U2258 ( .A(n2699), .B(n2700), .Z(n2690) );
  AND U2259 ( .A(n2701), .B(n2702), .Z(n2700) );
  XOR U2260 ( .A(n2699), .B(n2393), .Z(n2702) );
  XNOR U2261 ( .A(p_input[4043]), .B(n2703), .Z(n2393) );
  AND U2262 ( .A(n182), .B(n2704), .Z(n2703) );
  XOR U2263 ( .A(p_input[4075]), .B(p_input[4043]), .Z(n2704) );
  XNOR U2264 ( .A(n2390), .B(n2699), .Z(n2701) );
  XOR U2265 ( .A(n2705), .B(n2706), .Z(n2390) );
  AND U2266 ( .A(n180), .B(n2707), .Z(n2706) );
  XOR U2267 ( .A(p_input[4011]), .B(p_input[3979]), .Z(n2707) );
  XOR U2268 ( .A(n2708), .B(n2709), .Z(n2699) );
  AND U2269 ( .A(n2710), .B(n2711), .Z(n2709) );
  XOR U2270 ( .A(n2708), .B(n2405), .Z(n2711) );
  XNOR U2271 ( .A(p_input[4042]), .B(n2712), .Z(n2405) );
  AND U2272 ( .A(n182), .B(n2713), .Z(n2712) );
  XOR U2273 ( .A(p_input[4074]), .B(p_input[4042]), .Z(n2713) );
  XNOR U2274 ( .A(n2402), .B(n2708), .Z(n2710) );
  XOR U2275 ( .A(n2714), .B(n2715), .Z(n2402) );
  AND U2276 ( .A(n180), .B(n2716), .Z(n2715) );
  XOR U2277 ( .A(p_input[4010]), .B(p_input[3978]), .Z(n2716) );
  XOR U2278 ( .A(n2717), .B(n2718), .Z(n2708) );
  AND U2279 ( .A(n2719), .B(n2720), .Z(n2718) );
  XOR U2280 ( .A(n2717), .B(n2417), .Z(n2720) );
  XNOR U2281 ( .A(p_input[4041]), .B(n2721), .Z(n2417) );
  AND U2282 ( .A(n182), .B(n2722), .Z(n2721) );
  XOR U2283 ( .A(p_input[4073]), .B(p_input[4041]), .Z(n2722) );
  XNOR U2284 ( .A(n2414), .B(n2717), .Z(n2719) );
  XOR U2285 ( .A(n2723), .B(n2724), .Z(n2414) );
  AND U2286 ( .A(n180), .B(n2725), .Z(n2724) );
  XOR U2287 ( .A(p_input[4009]), .B(p_input[3977]), .Z(n2725) );
  XOR U2288 ( .A(n2726), .B(n2727), .Z(n2717) );
  AND U2289 ( .A(n2728), .B(n2729), .Z(n2727) );
  XOR U2290 ( .A(n2726), .B(n2429), .Z(n2729) );
  XNOR U2291 ( .A(p_input[4040]), .B(n2730), .Z(n2429) );
  AND U2292 ( .A(n182), .B(n2731), .Z(n2730) );
  XOR U2293 ( .A(p_input[4072]), .B(p_input[4040]), .Z(n2731) );
  XNOR U2294 ( .A(n2426), .B(n2726), .Z(n2728) );
  XOR U2295 ( .A(n2732), .B(n2733), .Z(n2426) );
  AND U2296 ( .A(n180), .B(n2734), .Z(n2733) );
  XOR U2297 ( .A(p_input[4008]), .B(p_input[3976]), .Z(n2734) );
  XOR U2298 ( .A(n2735), .B(n2736), .Z(n2726) );
  AND U2299 ( .A(n2737), .B(n2738), .Z(n2736) );
  XOR U2300 ( .A(n2735), .B(n2441), .Z(n2738) );
  XNOR U2301 ( .A(p_input[4039]), .B(n2739), .Z(n2441) );
  AND U2302 ( .A(n182), .B(n2740), .Z(n2739) );
  XOR U2303 ( .A(p_input[4071]), .B(p_input[4039]), .Z(n2740) );
  XNOR U2304 ( .A(n2438), .B(n2735), .Z(n2737) );
  XOR U2305 ( .A(n2741), .B(n2742), .Z(n2438) );
  AND U2306 ( .A(n180), .B(n2743), .Z(n2742) );
  XOR U2307 ( .A(p_input[4007]), .B(p_input[3975]), .Z(n2743) );
  XOR U2308 ( .A(n2744), .B(n2745), .Z(n2735) );
  AND U2309 ( .A(n2746), .B(n2747), .Z(n2745) );
  XOR U2310 ( .A(n2744), .B(n2453), .Z(n2747) );
  XNOR U2311 ( .A(p_input[4038]), .B(n2748), .Z(n2453) );
  AND U2312 ( .A(n182), .B(n2749), .Z(n2748) );
  XOR U2313 ( .A(p_input[4070]), .B(p_input[4038]), .Z(n2749) );
  XNOR U2314 ( .A(n2450), .B(n2744), .Z(n2746) );
  XOR U2315 ( .A(n2750), .B(n2751), .Z(n2450) );
  AND U2316 ( .A(n180), .B(n2752), .Z(n2751) );
  XOR U2317 ( .A(p_input[4006]), .B(p_input[3974]), .Z(n2752) );
  XOR U2318 ( .A(n2753), .B(n2754), .Z(n2744) );
  AND U2319 ( .A(n2755), .B(n2756), .Z(n2754) );
  XOR U2320 ( .A(n2753), .B(n2465), .Z(n2756) );
  XNOR U2321 ( .A(p_input[4037]), .B(n2757), .Z(n2465) );
  AND U2322 ( .A(n182), .B(n2758), .Z(n2757) );
  XOR U2323 ( .A(p_input[4069]), .B(p_input[4037]), .Z(n2758) );
  XNOR U2324 ( .A(n2462), .B(n2753), .Z(n2755) );
  XOR U2325 ( .A(n2759), .B(n2760), .Z(n2462) );
  AND U2326 ( .A(n180), .B(n2761), .Z(n2760) );
  XOR U2327 ( .A(p_input[4005]), .B(p_input[3973]), .Z(n2761) );
  XOR U2328 ( .A(n2762), .B(n2763), .Z(n2753) );
  AND U2329 ( .A(n2764), .B(n2765), .Z(n2763) );
  XOR U2330 ( .A(n2762), .B(n2477), .Z(n2765) );
  XNOR U2331 ( .A(p_input[4036]), .B(n2766), .Z(n2477) );
  AND U2332 ( .A(n182), .B(n2767), .Z(n2766) );
  XOR U2333 ( .A(p_input[4068]), .B(p_input[4036]), .Z(n2767) );
  XNOR U2334 ( .A(n2474), .B(n2762), .Z(n2764) );
  XOR U2335 ( .A(n2768), .B(n2769), .Z(n2474) );
  AND U2336 ( .A(n180), .B(n2770), .Z(n2769) );
  XOR U2337 ( .A(p_input[4004]), .B(p_input[3972]), .Z(n2770) );
  XOR U2338 ( .A(n2771), .B(n2772), .Z(n2762) );
  AND U2339 ( .A(n2773), .B(n2774), .Z(n2772) );
  XOR U2340 ( .A(n2771), .B(n2489), .Z(n2774) );
  XNOR U2341 ( .A(p_input[4035]), .B(n2775), .Z(n2489) );
  AND U2342 ( .A(n182), .B(n2776), .Z(n2775) );
  XOR U2343 ( .A(p_input[4067]), .B(p_input[4035]), .Z(n2776) );
  XNOR U2344 ( .A(n2486), .B(n2771), .Z(n2773) );
  XOR U2345 ( .A(n2777), .B(n2778), .Z(n2486) );
  AND U2346 ( .A(n180), .B(n2779), .Z(n2778) );
  XOR U2347 ( .A(p_input[4003]), .B(p_input[3971]), .Z(n2779) );
  XOR U2348 ( .A(n2780), .B(n2781), .Z(n2771) );
  AND U2349 ( .A(n2782), .B(n2783), .Z(n2781) );
  XOR U2350 ( .A(n2501), .B(n2780), .Z(n2783) );
  XNOR U2351 ( .A(p_input[4034]), .B(n2784), .Z(n2501) );
  AND U2352 ( .A(n182), .B(n2785), .Z(n2784) );
  XOR U2353 ( .A(p_input[4066]), .B(p_input[4034]), .Z(n2785) );
  XNOR U2354 ( .A(n2780), .B(n2498), .Z(n2782) );
  XOR U2355 ( .A(n2786), .B(n2787), .Z(n2498) );
  AND U2356 ( .A(n180), .B(n2788), .Z(n2787) );
  XOR U2357 ( .A(p_input[4002]), .B(p_input[3970]), .Z(n2788) );
  XOR U2358 ( .A(n2789), .B(n2790), .Z(n2780) );
  AND U2359 ( .A(n2791), .B(n2792), .Z(n2790) );
  XNOR U2360 ( .A(n2793), .B(n2514), .Z(n2792) );
  XNOR U2361 ( .A(p_input[4033]), .B(n2794), .Z(n2514) );
  AND U2362 ( .A(n182), .B(n2795), .Z(n2794) );
  XNOR U2363 ( .A(p_input[4065]), .B(n2796), .Z(n2795) );
  IV U2364 ( .A(p_input[4033]), .Z(n2796) );
  XNOR U2365 ( .A(n2511), .B(n2789), .Z(n2791) );
  XNOR U2366 ( .A(p_input[3969]), .B(n2797), .Z(n2511) );
  AND U2367 ( .A(n180), .B(n2798), .Z(n2797) );
  XOR U2368 ( .A(p_input[4001]), .B(p_input[3969]), .Z(n2798) );
  IV U2369 ( .A(n2793), .Z(n2789) );
  AND U2370 ( .A(n2519), .B(n2522), .Z(n2793) );
  XOR U2371 ( .A(p_input[4032]), .B(n2799), .Z(n2522) );
  AND U2372 ( .A(n182), .B(n2800), .Z(n2799) );
  XOR U2373 ( .A(p_input[4064]), .B(p_input[4032]), .Z(n2800) );
  XOR U2374 ( .A(n2801), .B(n2802), .Z(n182) );
  AND U2375 ( .A(n2803), .B(n2804), .Z(n2802) );
  XNOR U2376 ( .A(p_input[4095]), .B(n2801), .Z(n2804) );
  XOR U2377 ( .A(n2801), .B(p_input[4063]), .Z(n2803) );
  XOR U2378 ( .A(n2805), .B(n2806), .Z(n2801) );
  AND U2379 ( .A(n2807), .B(n2808), .Z(n2806) );
  XNOR U2380 ( .A(p_input[4094]), .B(n2805), .Z(n2808) );
  XOR U2381 ( .A(n2805), .B(p_input[4062]), .Z(n2807) );
  XOR U2382 ( .A(n2809), .B(n2810), .Z(n2805) );
  AND U2383 ( .A(n2811), .B(n2812), .Z(n2810) );
  XNOR U2384 ( .A(p_input[4093]), .B(n2809), .Z(n2812) );
  XOR U2385 ( .A(n2809), .B(p_input[4061]), .Z(n2811) );
  XOR U2386 ( .A(n2813), .B(n2814), .Z(n2809) );
  AND U2387 ( .A(n2815), .B(n2816), .Z(n2814) );
  XNOR U2388 ( .A(p_input[4092]), .B(n2813), .Z(n2816) );
  XOR U2389 ( .A(n2813), .B(p_input[4060]), .Z(n2815) );
  XOR U2390 ( .A(n2817), .B(n2818), .Z(n2813) );
  AND U2391 ( .A(n2819), .B(n2820), .Z(n2818) );
  XNOR U2392 ( .A(p_input[4091]), .B(n2817), .Z(n2820) );
  XOR U2393 ( .A(n2817), .B(p_input[4059]), .Z(n2819) );
  XOR U2394 ( .A(n2821), .B(n2822), .Z(n2817) );
  AND U2395 ( .A(n2823), .B(n2824), .Z(n2822) );
  XNOR U2396 ( .A(p_input[4090]), .B(n2821), .Z(n2824) );
  XOR U2397 ( .A(n2821), .B(p_input[4058]), .Z(n2823) );
  XOR U2398 ( .A(n2825), .B(n2826), .Z(n2821) );
  AND U2399 ( .A(n2827), .B(n2828), .Z(n2826) );
  XNOR U2400 ( .A(p_input[4089]), .B(n2825), .Z(n2828) );
  XOR U2401 ( .A(n2825), .B(p_input[4057]), .Z(n2827) );
  XOR U2402 ( .A(n2829), .B(n2830), .Z(n2825) );
  AND U2403 ( .A(n2831), .B(n2832), .Z(n2830) );
  XNOR U2404 ( .A(p_input[4088]), .B(n2829), .Z(n2832) );
  XOR U2405 ( .A(n2829), .B(p_input[4056]), .Z(n2831) );
  XOR U2406 ( .A(n2833), .B(n2834), .Z(n2829) );
  AND U2407 ( .A(n2835), .B(n2836), .Z(n2834) );
  XNOR U2408 ( .A(p_input[4087]), .B(n2833), .Z(n2836) );
  XOR U2409 ( .A(n2833), .B(p_input[4055]), .Z(n2835) );
  XOR U2410 ( .A(n2837), .B(n2838), .Z(n2833) );
  AND U2411 ( .A(n2839), .B(n2840), .Z(n2838) );
  XNOR U2412 ( .A(p_input[4086]), .B(n2837), .Z(n2840) );
  XOR U2413 ( .A(n2837), .B(p_input[4054]), .Z(n2839) );
  XOR U2414 ( .A(n2841), .B(n2842), .Z(n2837) );
  AND U2415 ( .A(n2843), .B(n2844), .Z(n2842) );
  XNOR U2416 ( .A(p_input[4085]), .B(n2841), .Z(n2844) );
  XOR U2417 ( .A(n2841), .B(p_input[4053]), .Z(n2843) );
  XOR U2418 ( .A(n2845), .B(n2846), .Z(n2841) );
  AND U2419 ( .A(n2847), .B(n2848), .Z(n2846) );
  XNOR U2420 ( .A(p_input[4084]), .B(n2845), .Z(n2848) );
  XOR U2421 ( .A(n2845), .B(p_input[4052]), .Z(n2847) );
  XOR U2422 ( .A(n2849), .B(n2850), .Z(n2845) );
  AND U2423 ( .A(n2851), .B(n2852), .Z(n2850) );
  XNOR U2424 ( .A(p_input[4083]), .B(n2849), .Z(n2852) );
  XOR U2425 ( .A(n2849), .B(p_input[4051]), .Z(n2851) );
  XOR U2426 ( .A(n2853), .B(n2854), .Z(n2849) );
  AND U2427 ( .A(n2855), .B(n2856), .Z(n2854) );
  XNOR U2428 ( .A(p_input[4082]), .B(n2853), .Z(n2856) );
  XOR U2429 ( .A(n2853), .B(p_input[4050]), .Z(n2855) );
  XOR U2430 ( .A(n2857), .B(n2858), .Z(n2853) );
  AND U2431 ( .A(n2859), .B(n2860), .Z(n2858) );
  XNOR U2432 ( .A(p_input[4081]), .B(n2857), .Z(n2860) );
  XOR U2433 ( .A(n2857), .B(p_input[4049]), .Z(n2859) );
  XOR U2434 ( .A(n2861), .B(n2862), .Z(n2857) );
  AND U2435 ( .A(n2863), .B(n2864), .Z(n2862) );
  XNOR U2436 ( .A(p_input[4080]), .B(n2861), .Z(n2864) );
  XOR U2437 ( .A(n2861), .B(p_input[4048]), .Z(n2863) );
  XOR U2438 ( .A(n2865), .B(n2866), .Z(n2861) );
  AND U2439 ( .A(n2867), .B(n2868), .Z(n2866) );
  XNOR U2440 ( .A(p_input[4079]), .B(n2865), .Z(n2868) );
  XOR U2441 ( .A(n2865), .B(p_input[4047]), .Z(n2867) );
  XOR U2442 ( .A(n2869), .B(n2870), .Z(n2865) );
  AND U2443 ( .A(n2871), .B(n2872), .Z(n2870) );
  XNOR U2444 ( .A(p_input[4078]), .B(n2869), .Z(n2872) );
  XOR U2445 ( .A(n2869), .B(p_input[4046]), .Z(n2871) );
  XOR U2446 ( .A(n2873), .B(n2874), .Z(n2869) );
  AND U2447 ( .A(n2875), .B(n2876), .Z(n2874) );
  XNOR U2448 ( .A(p_input[4077]), .B(n2873), .Z(n2876) );
  XOR U2449 ( .A(n2873), .B(p_input[4045]), .Z(n2875) );
  XOR U2450 ( .A(n2877), .B(n2878), .Z(n2873) );
  AND U2451 ( .A(n2879), .B(n2880), .Z(n2878) );
  XNOR U2452 ( .A(p_input[4076]), .B(n2877), .Z(n2880) );
  XOR U2453 ( .A(n2877), .B(p_input[4044]), .Z(n2879) );
  XOR U2454 ( .A(n2881), .B(n2882), .Z(n2877) );
  AND U2455 ( .A(n2883), .B(n2884), .Z(n2882) );
  XNOR U2456 ( .A(p_input[4075]), .B(n2881), .Z(n2884) );
  XOR U2457 ( .A(n2881), .B(p_input[4043]), .Z(n2883) );
  XOR U2458 ( .A(n2885), .B(n2886), .Z(n2881) );
  AND U2459 ( .A(n2887), .B(n2888), .Z(n2886) );
  XNOR U2460 ( .A(p_input[4074]), .B(n2885), .Z(n2888) );
  XOR U2461 ( .A(n2885), .B(p_input[4042]), .Z(n2887) );
  XOR U2462 ( .A(n2889), .B(n2890), .Z(n2885) );
  AND U2463 ( .A(n2891), .B(n2892), .Z(n2890) );
  XNOR U2464 ( .A(p_input[4073]), .B(n2889), .Z(n2892) );
  XOR U2465 ( .A(n2889), .B(p_input[4041]), .Z(n2891) );
  XOR U2466 ( .A(n2893), .B(n2894), .Z(n2889) );
  AND U2467 ( .A(n2895), .B(n2896), .Z(n2894) );
  XNOR U2468 ( .A(p_input[4072]), .B(n2893), .Z(n2896) );
  XOR U2469 ( .A(n2893), .B(p_input[4040]), .Z(n2895) );
  XOR U2470 ( .A(n2897), .B(n2898), .Z(n2893) );
  AND U2471 ( .A(n2899), .B(n2900), .Z(n2898) );
  XNOR U2472 ( .A(p_input[4071]), .B(n2897), .Z(n2900) );
  XOR U2473 ( .A(n2897), .B(p_input[4039]), .Z(n2899) );
  XOR U2474 ( .A(n2901), .B(n2902), .Z(n2897) );
  AND U2475 ( .A(n2903), .B(n2904), .Z(n2902) );
  XNOR U2476 ( .A(p_input[4070]), .B(n2901), .Z(n2904) );
  XOR U2477 ( .A(n2901), .B(p_input[4038]), .Z(n2903) );
  XOR U2478 ( .A(n2905), .B(n2906), .Z(n2901) );
  AND U2479 ( .A(n2907), .B(n2908), .Z(n2906) );
  XNOR U2480 ( .A(p_input[4069]), .B(n2905), .Z(n2908) );
  XOR U2481 ( .A(n2905), .B(p_input[4037]), .Z(n2907) );
  XOR U2482 ( .A(n2909), .B(n2910), .Z(n2905) );
  AND U2483 ( .A(n2911), .B(n2912), .Z(n2910) );
  XNOR U2484 ( .A(p_input[4068]), .B(n2909), .Z(n2912) );
  XOR U2485 ( .A(n2909), .B(p_input[4036]), .Z(n2911) );
  XOR U2486 ( .A(n2913), .B(n2914), .Z(n2909) );
  AND U2487 ( .A(n2915), .B(n2916), .Z(n2914) );
  XNOR U2488 ( .A(p_input[4067]), .B(n2913), .Z(n2916) );
  XOR U2489 ( .A(n2913), .B(p_input[4035]), .Z(n2915) );
  XOR U2490 ( .A(n2917), .B(n2918), .Z(n2913) );
  AND U2491 ( .A(n2919), .B(n2920), .Z(n2918) );
  XNOR U2492 ( .A(p_input[4066]), .B(n2917), .Z(n2920) );
  XOR U2493 ( .A(n2917), .B(p_input[4034]), .Z(n2919) );
  XNOR U2494 ( .A(n2921), .B(n2922), .Z(n2917) );
  AND U2495 ( .A(n2923), .B(n2924), .Z(n2922) );
  XOR U2496 ( .A(p_input[4065]), .B(n2921), .Z(n2924) );
  XNOR U2497 ( .A(p_input[4033]), .B(n2921), .Z(n2923) );
  AND U2498 ( .A(p_input[4064]), .B(n2925), .Z(n2921) );
  IV U2499 ( .A(p_input[4032]), .Z(n2925) );
  XNOR U2500 ( .A(p_input[3968]), .B(n2926), .Z(n2519) );
  AND U2501 ( .A(n180), .B(n2927), .Z(n2926) );
  XOR U2502 ( .A(p_input[4000]), .B(p_input[3968]), .Z(n2927) );
  XOR U2503 ( .A(n2928), .B(n2929), .Z(n180) );
  AND U2504 ( .A(n2930), .B(n2931), .Z(n2929) );
  XNOR U2505 ( .A(p_input[4031]), .B(n2928), .Z(n2931) );
  XOR U2506 ( .A(n2928), .B(p_input[3999]), .Z(n2930) );
  XOR U2507 ( .A(n2932), .B(n2933), .Z(n2928) );
  AND U2508 ( .A(n2934), .B(n2935), .Z(n2933) );
  XNOR U2509 ( .A(p_input[4030]), .B(n2932), .Z(n2935) );
  XNOR U2510 ( .A(n2932), .B(n2534), .Z(n2934) );
  IV U2511 ( .A(p_input[3998]), .Z(n2534) );
  XOR U2512 ( .A(n2936), .B(n2937), .Z(n2932) );
  AND U2513 ( .A(n2938), .B(n2939), .Z(n2937) );
  XNOR U2514 ( .A(p_input[4029]), .B(n2936), .Z(n2939) );
  XNOR U2515 ( .A(n2936), .B(n2543), .Z(n2938) );
  IV U2516 ( .A(p_input[3997]), .Z(n2543) );
  XOR U2517 ( .A(n2940), .B(n2941), .Z(n2936) );
  AND U2518 ( .A(n2942), .B(n2943), .Z(n2941) );
  XNOR U2519 ( .A(p_input[4028]), .B(n2940), .Z(n2943) );
  XNOR U2520 ( .A(n2940), .B(n2552), .Z(n2942) );
  IV U2521 ( .A(p_input[3996]), .Z(n2552) );
  XOR U2522 ( .A(n2944), .B(n2945), .Z(n2940) );
  AND U2523 ( .A(n2946), .B(n2947), .Z(n2945) );
  XNOR U2524 ( .A(p_input[4027]), .B(n2944), .Z(n2947) );
  XNOR U2525 ( .A(n2944), .B(n2561), .Z(n2946) );
  IV U2526 ( .A(p_input[3995]), .Z(n2561) );
  XOR U2527 ( .A(n2948), .B(n2949), .Z(n2944) );
  AND U2528 ( .A(n2950), .B(n2951), .Z(n2949) );
  XNOR U2529 ( .A(p_input[4026]), .B(n2948), .Z(n2951) );
  XNOR U2530 ( .A(n2948), .B(n2570), .Z(n2950) );
  IV U2531 ( .A(p_input[3994]), .Z(n2570) );
  XOR U2532 ( .A(n2952), .B(n2953), .Z(n2948) );
  AND U2533 ( .A(n2954), .B(n2955), .Z(n2953) );
  XNOR U2534 ( .A(p_input[4025]), .B(n2952), .Z(n2955) );
  XNOR U2535 ( .A(n2952), .B(n2579), .Z(n2954) );
  IV U2536 ( .A(p_input[3993]), .Z(n2579) );
  XOR U2537 ( .A(n2956), .B(n2957), .Z(n2952) );
  AND U2538 ( .A(n2958), .B(n2959), .Z(n2957) );
  XNOR U2539 ( .A(p_input[4024]), .B(n2956), .Z(n2959) );
  XNOR U2540 ( .A(n2956), .B(n2588), .Z(n2958) );
  IV U2541 ( .A(p_input[3992]), .Z(n2588) );
  XOR U2542 ( .A(n2960), .B(n2961), .Z(n2956) );
  AND U2543 ( .A(n2962), .B(n2963), .Z(n2961) );
  XNOR U2544 ( .A(p_input[4023]), .B(n2960), .Z(n2963) );
  XNOR U2545 ( .A(n2960), .B(n2597), .Z(n2962) );
  IV U2546 ( .A(p_input[3991]), .Z(n2597) );
  XOR U2547 ( .A(n2964), .B(n2965), .Z(n2960) );
  AND U2548 ( .A(n2966), .B(n2967), .Z(n2965) );
  XNOR U2549 ( .A(p_input[4022]), .B(n2964), .Z(n2967) );
  XNOR U2550 ( .A(n2964), .B(n2606), .Z(n2966) );
  IV U2551 ( .A(p_input[3990]), .Z(n2606) );
  XOR U2552 ( .A(n2968), .B(n2969), .Z(n2964) );
  AND U2553 ( .A(n2970), .B(n2971), .Z(n2969) );
  XNOR U2554 ( .A(p_input[4021]), .B(n2968), .Z(n2971) );
  XNOR U2555 ( .A(n2968), .B(n2615), .Z(n2970) );
  IV U2556 ( .A(p_input[3989]), .Z(n2615) );
  XOR U2557 ( .A(n2972), .B(n2973), .Z(n2968) );
  AND U2558 ( .A(n2974), .B(n2975), .Z(n2973) );
  XNOR U2559 ( .A(p_input[4020]), .B(n2972), .Z(n2975) );
  XNOR U2560 ( .A(n2972), .B(n2624), .Z(n2974) );
  IV U2561 ( .A(p_input[3988]), .Z(n2624) );
  XOR U2562 ( .A(n2976), .B(n2977), .Z(n2972) );
  AND U2563 ( .A(n2978), .B(n2979), .Z(n2977) );
  XNOR U2564 ( .A(p_input[4019]), .B(n2976), .Z(n2979) );
  XNOR U2565 ( .A(n2976), .B(n2633), .Z(n2978) );
  IV U2566 ( .A(p_input[3987]), .Z(n2633) );
  XOR U2567 ( .A(n2980), .B(n2981), .Z(n2976) );
  AND U2568 ( .A(n2982), .B(n2983), .Z(n2981) );
  XNOR U2569 ( .A(p_input[4018]), .B(n2980), .Z(n2983) );
  XNOR U2570 ( .A(n2980), .B(n2642), .Z(n2982) );
  IV U2571 ( .A(p_input[3986]), .Z(n2642) );
  XOR U2572 ( .A(n2984), .B(n2985), .Z(n2980) );
  AND U2573 ( .A(n2986), .B(n2987), .Z(n2985) );
  XNOR U2574 ( .A(p_input[4017]), .B(n2984), .Z(n2987) );
  XNOR U2575 ( .A(n2984), .B(n2651), .Z(n2986) );
  IV U2576 ( .A(p_input[3985]), .Z(n2651) );
  XOR U2577 ( .A(n2988), .B(n2989), .Z(n2984) );
  AND U2578 ( .A(n2990), .B(n2991), .Z(n2989) );
  XNOR U2579 ( .A(p_input[4016]), .B(n2988), .Z(n2991) );
  XNOR U2580 ( .A(n2988), .B(n2660), .Z(n2990) );
  IV U2581 ( .A(p_input[3984]), .Z(n2660) );
  XOR U2582 ( .A(n2992), .B(n2993), .Z(n2988) );
  AND U2583 ( .A(n2994), .B(n2995), .Z(n2993) );
  XNOR U2584 ( .A(p_input[4015]), .B(n2992), .Z(n2995) );
  XNOR U2585 ( .A(n2992), .B(n2669), .Z(n2994) );
  IV U2586 ( .A(p_input[3983]), .Z(n2669) );
  XOR U2587 ( .A(n2996), .B(n2997), .Z(n2992) );
  AND U2588 ( .A(n2998), .B(n2999), .Z(n2997) );
  XNOR U2589 ( .A(p_input[4014]), .B(n2996), .Z(n2999) );
  XNOR U2590 ( .A(n2996), .B(n2678), .Z(n2998) );
  IV U2591 ( .A(p_input[3982]), .Z(n2678) );
  XOR U2592 ( .A(n3000), .B(n3001), .Z(n2996) );
  AND U2593 ( .A(n3002), .B(n3003), .Z(n3001) );
  XNOR U2594 ( .A(p_input[4013]), .B(n3000), .Z(n3003) );
  XNOR U2595 ( .A(n3000), .B(n2687), .Z(n3002) );
  IV U2596 ( .A(p_input[3981]), .Z(n2687) );
  XOR U2597 ( .A(n3004), .B(n3005), .Z(n3000) );
  AND U2598 ( .A(n3006), .B(n3007), .Z(n3005) );
  XNOR U2599 ( .A(p_input[4012]), .B(n3004), .Z(n3007) );
  XNOR U2600 ( .A(n3004), .B(n2696), .Z(n3006) );
  IV U2601 ( .A(p_input[3980]), .Z(n2696) );
  XOR U2602 ( .A(n3008), .B(n3009), .Z(n3004) );
  AND U2603 ( .A(n3010), .B(n3011), .Z(n3009) );
  XNOR U2604 ( .A(p_input[4011]), .B(n3008), .Z(n3011) );
  XNOR U2605 ( .A(n3008), .B(n2705), .Z(n3010) );
  IV U2606 ( .A(p_input[3979]), .Z(n2705) );
  XOR U2607 ( .A(n3012), .B(n3013), .Z(n3008) );
  AND U2608 ( .A(n3014), .B(n3015), .Z(n3013) );
  XNOR U2609 ( .A(p_input[4010]), .B(n3012), .Z(n3015) );
  XNOR U2610 ( .A(n3012), .B(n2714), .Z(n3014) );
  IV U2611 ( .A(p_input[3978]), .Z(n2714) );
  XOR U2612 ( .A(n3016), .B(n3017), .Z(n3012) );
  AND U2613 ( .A(n3018), .B(n3019), .Z(n3017) );
  XNOR U2614 ( .A(p_input[4009]), .B(n3016), .Z(n3019) );
  XNOR U2615 ( .A(n3016), .B(n2723), .Z(n3018) );
  IV U2616 ( .A(p_input[3977]), .Z(n2723) );
  XOR U2617 ( .A(n3020), .B(n3021), .Z(n3016) );
  AND U2618 ( .A(n3022), .B(n3023), .Z(n3021) );
  XNOR U2619 ( .A(p_input[4008]), .B(n3020), .Z(n3023) );
  XNOR U2620 ( .A(n3020), .B(n2732), .Z(n3022) );
  IV U2621 ( .A(p_input[3976]), .Z(n2732) );
  XOR U2622 ( .A(n3024), .B(n3025), .Z(n3020) );
  AND U2623 ( .A(n3026), .B(n3027), .Z(n3025) );
  XNOR U2624 ( .A(p_input[4007]), .B(n3024), .Z(n3027) );
  XNOR U2625 ( .A(n3024), .B(n2741), .Z(n3026) );
  IV U2626 ( .A(p_input[3975]), .Z(n2741) );
  XOR U2627 ( .A(n3028), .B(n3029), .Z(n3024) );
  AND U2628 ( .A(n3030), .B(n3031), .Z(n3029) );
  XNOR U2629 ( .A(p_input[4006]), .B(n3028), .Z(n3031) );
  XNOR U2630 ( .A(n3028), .B(n2750), .Z(n3030) );
  IV U2631 ( .A(p_input[3974]), .Z(n2750) );
  XOR U2632 ( .A(n3032), .B(n3033), .Z(n3028) );
  AND U2633 ( .A(n3034), .B(n3035), .Z(n3033) );
  XNOR U2634 ( .A(p_input[4005]), .B(n3032), .Z(n3035) );
  XNOR U2635 ( .A(n3032), .B(n2759), .Z(n3034) );
  IV U2636 ( .A(p_input[3973]), .Z(n2759) );
  XOR U2637 ( .A(n3036), .B(n3037), .Z(n3032) );
  AND U2638 ( .A(n3038), .B(n3039), .Z(n3037) );
  XNOR U2639 ( .A(p_input[4004]), .B(n3036), .Z(n3039) );
  XNOR U2640 ( .A(n3036), .B(n2768), .Z(n3038) );
  IV U2641 ( .A(p_input[3972]), .Z(n2768) );
  XOR U2642 ( .A(n3040), .B(n3041), .Z(n3036) );
  AND U2643 ( .A(n3042), .B(n3043), .Z(n3041) );
  XNOR U2644 ( .A(p_input[4003]), .B(n3040), .Z(n3043) );
  XNOR U2645 ( .A(n3040), .B(n2777), .Z(n3042) );
  IV U2646 ( .A(p_input[3971]), .Z(n2777) );
  XOR U2647 ( .A(n3044), .B(n3045), .Z(n3040) );
  AND U2648 ( .A(n3046), .B(n3047), .Z(n3045) );
  XNOR U2649 ( .A(p_input[4002]), .B(n3044), .Z(n3047) );
  XNOR U2650 ( .A(n3044), .B(n2786), .Z(n3046) );
  IV U2651 ( .A(p_input[3970]), .Z(n2786) );
  XNOR U2652 ( .A(n3048), .B(n3049), .Z(n3044) );
  AND U2653 ( .A(n3050), .B(n3051), .Z(n3049) );
  XOR U2654 ( .A(p_input[4001]), .B(n3048), .Z(n3051) );
  XNOR U2655 ( .A(p_input[3969]), .B(n3048), .Z(n3050) );
  AND U2656 ( .A(p_input[4000]), .B(n3052), .Z(n3048) );
  IV U2657 ( .A(p_input[3968]), .Z(n3052) );
  XOR U2658 ( .A(n3053), .B(n3054), .Z(n2142) );
  AND U2659 ( .A(n304), .B(n3055), .Z(n3054) );
  XNOR U2660 ( .A(n3056), .B(n3053), .Z(n3055) );
  XOR U2661 ( .A(n3057), .B(n3058), .Z(n304) );
  AND U2662 ( .A(n3059), .B(n3060), .Z(n3058) );
  XNOR U2663 ( .A(n2157), .B(n3057), .Z(n3060) );
  AND U2664 ( .A(p_input[3967]), .B(p_input[3935]), .Z(n2157) );
  XNOR U2665 ( .A(n3057), .B(n2154), .Z(n3059) );
  IV U2666 ( .A(n3061), .Z(n2154) );
  AND U2667 ( .A(p_input[3871]), .B(p_input[3903]), .Z(n3061) );
  XOR U2668 ( .A(n3062), .B(n3063), .Z(n3057) );
  AND U2669 ( .A(n3064), .B(n3065), .Z(n3063) );
  XOR U2670 ( .A(n3062), .B(n2169), .Z(n3065) );
  XNOR U2671 ( .A(p_input[3934]), .B(n3066), .Z(n2169) );
  AND U2672 ( .A(n186), .B(n3067), .Z(n3066) );
  XOR U2673 ( .A(p_input[3966]), .B(p_input[3934]), .Z(n3067) );
  XNOR U2674 ( .A(n2166), .B(n3062), .Z(n3064) );
  XOR U2675 ( .A(n3068), .B(n3069), .Z(n2166) );
  AND U2676 ( .A(n183), .B(n3070), .Z(n3069) );
  XOR U2677 ( .A(p_input[3902]), .B(p_input[3870]), .Z(n3070) );
  XOR U2678 ( .A(n3071), .B(n3072), .Z(n3062) );
  AND U2679 ( .A(n3073), .B(n3074), .Z(n3072) );
  XOR U2680 ( .A(n3071), .B(n2181), .Z(n3074) );
  XNOR U2681 ( .A(p_input[3933]), .B(n3075), .Z(n2181) );
  AND U2682 ( .A(n186), .B(n3076), .Z(n3075) );
  XOR U2683 ( .A(p_input[3965]), .B(p_input[3933]), .Z(n3076) );
  XNOR U2684 ( .A(n2178), .B(n3071), .Z(n3073) );
  XOR U2685 ( .A(n3077), .B(n3078), .Z(n2178) );
  AND U2686 ( .A(n183), .B(n3079), .Z(n3078) );
  XOR U2687 ( .A(p_input[3901]), .B(p_input[3869]), .Z(n3079) );
  XOR U2688 ( .A(n3080), .B(n3081), .Z(n3071) );
  AND U2689 ( .A(n3082), .B(n3083), .Z(n3081) );
  XOR U2690 ( .A(n3080), .B(n2193), .Z(n3083) );
  XNOR U2691 ( .A(p_input[3932]), .B(n3084), .Z(n2193) );
  AND U2692 ( .A(n186), .B(n3085), .Z(n3084) );
  XOR U2693 ( .A(p_input[3964]), .B(p_input[3932]), .Z(n3085) );
  XNOR U2694 ( .A(n2190), .B(n3080), .Z(n3082) );
  XOR U2695 ( .A(n3086), .B(n3087), .Z(n2190) );
  AND U2696 ( .A(n183), .B(n3088), .Z(n3087) );
  XOR U2697 ( .A(p_input[3900]), .B(p_input[3868]), .Z(n3088) );
  XOR U2698 ( .A(n3089), .B(n3090), .Z(n3080) );
  AND U2699 ( .A(n3091), .B(n3092), .Z(n3090) );
  XOR U2700 ( .A(n3089), .B(n2205), .Z(n3092) );
  XNOR U2701 ( .A(p_input[3931]), .B(n3093), .Z(n2205) );
  AND U2702 ( .A(n186), .B(n3094), .Z(n3093) );
  XOR U2703 ( .A(p_input[3963]), .B(p_input[3931]), .Z(n3094) );
  XNOR U2704 ( .A(n2202), .B(n3089), .Z(n3091) );
  XOR U2705 ( .A(n3095), .B(n3096), .Z(n2202) );
  AND U2706 ( .A(n183), .B(n3097), .Z(n3096) );
  XOR U2707 ( .A(p_input[3899]), .B(p_input[3867]), .Z(n3097) );
  XOR U2708 ( .A(n3098), .B(n3099), .Z(n3089) );
  AND U2709 ( .A(n3100), .B(n3101), .Z(n3099) );
  XOR U2710 ( .A(n3098), .B(n2217), .Z(n3101) );
  XNOR U2711 ( .A(p_input[3930]), .B(n3102), .Z(n2217) );
  AND U2712 ( .A(n186), .B(n3103), .Z(n3102) );
  XOR U2713 ( .A(p_input[3962]), .B(p_input[3930]), .Z(n3103) );
  XNOR U2714 ( .A(n2214), .B(n3098), .Z(n3100) );
  XOR U2715 ( .A(n3104), .B(n3105), .Z(n2214) );
  AND U2716 ( .A(n183), .B(n3106), .Z(n3105) );
  XOR U2717 ( .A(p_input[3898]), .B(p_input[3866]), .Z(n3106) );
  XOR U2718 ( .A(n3107), .B(n3108), .Z(n3098) );
  AND U2719 ( .A(n3109), .B(n3110), .Z(n3108) );
  XOR U2720 ( .A(n3107), .B(n2229), .Z(n3110) );
  XNOR U2721 ( .A(p_input[3929]), .B(n3111), .Z(n2229) );
  AND U2722 ( .A(n186), .B(n3112), .Z(n3111) );
  XOR U2723 ( .A(p_input[3961]), .B(p_input[3929]), .Z(n3112) );
  XNOR U2724 ( .A(n2226), .B(n3107), .Z(n3109) );
  XOR U2725 ( .A(n3113), .B(n3114), .Z(n2226) );
  AND U2726 ( .A(n183), .B(n3115), .Z(n3114) );
  XOR U2727 ( .A(p_input[3897]), .B(p_input[3865]), .Z(n3115) );
  XOR U2728 ( .A(n3116), .B(n3117), .Z(n3107) );
  AND U2729 ( .A(n3118), .B(n3119), .Z(n3117) );
  XOR U2730 ( .A(n3116), .B(n2241), .Z(n3119) );
  XNOR U2731 ( .A(p_input[3928]), .B(n3120), .Z(n2241) );
  AND U2732 ( .A(n186), .B(n3121), .Z(n3120) );
  XOR U2733 ( .A(p_input[3960]), .B(p_input[3928]), .Z(n3121) );
  XNOR U2734 ( .A(n2238), .B(n3116), .Z(n3118) );
  XOR U2735 ( .A(n3122), .B(n3123), .Z(n2238) );
  AND U2736 ( .A(n183), .B(n3124), .Z(n3123) );
  XOR U2737 ( .A(p_input[3896]), .B(p_input[3864]), .Z(n3124) );
  XOR U2738 ( .A(n3125), .B(n3126), .Z(n3116) );
  AND U2739 ( .A(n3127), .B(n3128), .Z(n3126) );
  XOR U2740 ( .A(n3125), .B(n2253), .Z(n3128) );
  XNOR U2741 ( .A(p_input[3927]), .B(n3129), .Z(n2253) );
  AND U2742 ( .A(n186), .B(n3130), .Z(n3129) );
  XOR U2743 ( .A(p_input[3959]), .B(p_input[3927]), .Z(n3130) );
  XNOR U2744 ( .A(n2250), .B(n3125), .Z(n3127) );
  XOR U2745 ( .A(n3131), .B(n3132), .Z(n2250) );
  AND U2746 ( .A(n183), .B(n3133), .Z(n3132) );
  XOR U2747 ( .A(p_input[3895]), .B(p_input[3863]), .Z(n3133) );
  XOR U2748 ( .A(n3134), .B(n3135), .Z(n3125) );
  AND U2749 ( .A(n3136), .B(n3137), .Z(n3135) );
  XOR U2750 ( .A(n3134), .B(n2265), .Z(n3137) );
  XNOR U2751 ( .A(p_input[3926]), .B(n3138), .Z(n2265) );
  AND U2752 ( .A(n186), .B(n3139), .Z(n3138) );
  XOR U2753 ( .A(p_input[3958]), .B(p_input[3926]), .Z(n3139) );
  XNOR U2754 ( .A(n2262), .B(n3134), .Z(n3136) );
  XOR U2755 ( .A(n3140), .B(n3141), .Z(n2262) );
  AND U2756 ( .A(n183), .B(n3142), .Z(n3141) );
  XOR U2757 ( .A(p_input[3894]), .B(p_input[3862]), .Z(n3142) );
  XOR U2758 ( .A(n3143), .B(n3144), .Z(n3134) );
  AND U2759 ( .A(n3145), .B(n3146), .Z(n3144) );
  XOR U2760 ( .A(n3143), .B(n2277), .Z(n3146) );
  XNOR U2761 ( .A(p_input[3925]), .B(n3147), .Z(n2277) );
  AND U2762 ( .A(n186), .B(n3148), .Z(n3147) );
  XOR U2763 ( .A(p_input[3957]), .B(p_input[3925]), .Z(n3148) );
  XNOR U2764 ( .A(n2274), .B(n3143), .Z(n3145) );
  XOR U2765 ( .A(n3149), .B(n3150), .Z(n2274) );
  AND U2766 ( .A(n183), .B(n3151), .Z(n3150) );
  XOR U2767 ( .A(p_input[3893]), .B(p_input[3861]), .Z(n3151) );
  XOR U2768 ( .A(n3152), .B(n3153), .Z(n3143) );
  AND U2769 ( .A(n3154), .B(n3155), .Z(n3153) );
  XOR U2770 ( .A(n3152), .B(n2289), .Z(n3155) );
  XNOR U2771 ( .A(p_input[3924]), .B(n3156), .Z(n2289) );
  AND U2772 ( .A(n186), .B(n3157), .Z(n3156) );
  XOR U2773 ( .A(p_input[3956]), .B(p_input[3924]), .Z(n3157) );
  XNOR U2774 ( .A(n2286), .B(n3152), .Z(n3154) );
  XOR U2775 ( .A(n3158), .B(n3159), .Z(n2286) );
  AND U2776 ( .A(n183), .B(n3160), .Z(n3159) );
  XOR U2777 ( .A(p_input[3892]), .B(p_input[3860]), .Z(n3160) );
  XOR U2778 ( .A(n3161), .B(n3162), .Z(n3152) );
  AND U2779 ( .A(n3163), .B(n3164), .Z(n3162) );
  XOR U2780 ( .A(n3161), .B(n2301), .Z(n3164) );
  XNOR U2781 ( .A(p_input[3923]), .B(n3165), .Z(n2301) );
  AND U2782 ( .A(n186), .B(n3166), .Z(n3165) );
  XOR U2783 ( .A(p_input[3955]), .B(p_input[3923]), .Z(n3166) );
  XNOR U2784 ( .A(n2298), .B(n3161), .Z(n3163) );
  XOR U2785 ( .A(n3167), .B(n3168), .Z(n2298) );
  AND U2786 ( .A(n183), .B(n3169), .Z(n3168) );
  XOR U2787 ( .A(p_input[3891]), .B(p_input[3859]), .Z(n3169) );
  XOR U2788 ( .A(n3170), .B(n3171), .Z(n3161) );
  AND U2789 ( .A(n3172), .B(n3173), .Z(n3171) );
  XOR U2790 ( .A(n3170), .B(n2313), .Z(n3173) );
  XNOR U2791 ( .A(p_input[3922]), .B(n3174), .Z(n2313) );
  AND U2792 ( .A(n186), .B(n3175), .Z(n3174) );
  XOR U2793 ( .A(p_input[3954]), .B(p_input[3922]), .Z(n3175) );
  XNOR U2794 ( .A(n2310), .B(n3170), .Z(n3172) );
  XOR U2795 ( .A(n3176), .B(n3177), .Z(n2310) );
  AND U2796 ( .A(n183), .B(n3178), .Z(n3177) );
  XOR U2797 ( .A(p_input[3890]), .B(p_input[3858]), .Z(n3178) );
  XOR U2798 ( .A(n3179), .B(n3180), .Z(n3170) );
  AND U2799 ( .A(n3181), .B(n3182), .Z(n3180) );
  XOR U2800 ( .A(n3179), .B(n2325), .Z(n3182) );
  XNOR U2801 ( .A(p_input[3921]), .B(n3183), .Z(n2325) );
  AND U2802 ( .A(n186), .B(n3184), .Z(n3183) );
  XOR U2803 ( .A(p_input[3953]), .B(p_input[3921]), .Z(n3184) );
  XNOR U2804 ( .A(n2322), .B(n3179), .Z(n3181) );
  XOR U2805 ( .A(n3185), .B(n3186), .Z(n2322) );
  AND U2806 ( .A(n183), .B(n3187), .Z(n3186) );
  XOR U2807 ( .A(p_input[3889]), .B(p_input[3857]), .Z(n3187) );
  XOR U2808 ( .A(n3188), .B(n3189), .Z(n3179) );
  AND U2809 ( .A(n3190), .B(n3191), .Z(n3189) );
  XOR U2810 ( .A(n3188), .B(n2337), .Z(n3191) );
  XNOR U2811 ( .A(p_input[3920]), .B(n3192), .Z(n2337) );
  AND U2812 ( .A(n186), .B(n3193), .Z(n3192) );
  XOR U2813 ( .A(p_input[3952]), .B(p_input[3920]), .Z(n3193) );
  XNOR U2814 ( .A(n2334), .B(n3188), .Z(n3190) );
  XOR U2815 ( .A(n3194), .B(n3195), .Z(n2334) );
  AND U2816 ( .A(n183), .B(n3196), .Z(n3195) );
  XOR U2817 ( .A(p_input[3888]), .B(p_input[3856]), .Z(n3196) );
  XOR U2818 ( .A(n3197), .B(n3198), .Z(n3188) );
  AND U2819 ( .A(n3199), .B(n3200), .Z(n3198) );
  XOR U2820 ( .A(n3197), .B(n2349), .Z(n3200) );
  XNOR U2821 ( .A(p_input[3919]), .B(n3201), .Z(n2349) );
  AND U2822 ( .A(n186), .B(n3202), .Z(n3201) );
  XOR U2823 ( .A(p_input[3951]), .B(p_input[3919]), .Z(n3202) );
  XNOR U2824 ( .A(n2346), .B(n3197), .Z(n3199) );
  XOR U2825 ( .A(n3203), .B(n3204), .Z(n2346) );
  AND U2826 ( .A(n183), .B(n3205), .Z(n3204) );
  XOR U2827 ( .A(p_input[3887]), .B(p_input[3855]), .Z(n3205) );
  XOR U2828 ( .A(n3206), .B(n3207), .Z(n3197) );
  AND U2829 ( .A(n3208), .B(n3209), .Z(n3207) );
  XOR U2830 ( .A(n3206), .B(n2361), .Z(n3209) );
  XNOR U2831 ( .A(p_input[3918]), .B(n3210), .Z(n2361) );
  AND U2832 ( .A(n186), .B(n3211), .Z(n3210) );
  XOR U2833 ( .A(p_input[3950]), .B(p_input[3918]), .Z(n3211) );
  XNOR U2834 ( .A(n2358), .B(n3206), .Z(n3208) );
  XOR U2835 ( .A(n3212), .B(n3213), .Z(n2358) );
  AND U2836 ( .A(n183), .B(n3214), .Z(n3213) );
  XOR U2837 ( .A(p_input[3886]), .B(p_input[3854]), .Z(n3214) );
  XOR U2838 ( .A(n3215), .B(n3216), .Z(n3206) );
  AND U2839 ( .A(n3217), .B(n3218), .Z(n3216) );
  XOR U2840 ( .A(n3215), .B(n2373), .Z(n3218) );
  XNOR U2841 ( .A(p_input[3917]), .B(n3219), .Z(n2373) );
  AND U2842 ( .A(n186), .B(n3220), .Z(n3219) );
  XOR U2843 ( .A(p_input[3949]), .B(p_input[3917]), .Z(n3220) );
  XNOR U2844 ( .A(n2370), .B(n3215), .Z(n3217) );
  XOR U2845 ( .A(n3221), .B(n3222), .Z(n2370) );
  AND U2846 ( .A(n183), .B(n3223), .Z(n3222) );
  XOR U2847 ( .A(p_input[3885]), .B(p_input[3853]), .Z(n3223) );
  XOR U2848 ( .A(n3224), .B(n3225), .Z(n3215) );
  AND U2849 ( .A(n3226), .B(n3227), .Z(n3225) );
  XOR U2850 ( .A(n3224), .B(n2385), .Z(n3227) );
  XNOR U2851 ( .A(p_input[3916]), .B(n3228), .Z(n2385) );
  AND U2852 ( .A(n186), .B(n3229), .Z(n3228) );
  XOR U2853 ( .A(p_input[3948]), .B(p_input[3916]), .Z(n3229) );
  XNOR U2854 ( .A(n2382), .B(n3224), .Z(n3226) );
  XOR U2855 ( .A(n3230), .B(n3231), .Z(n2382) );
  AND U2856 ( .A(n183), .B(n3232), .Z(n3231) );
  XOR U2857 ( .A(p_input[3884]), .B(p_input[3852]), .Z(n3232) );
  XOR U2858 ( .A(n3233), .B(n3234), .Z(n3224) );
  AND U2859 ( .A(n3235), .B(n3236), .Z(n3234) );
  XOR U2860 ( .A(n3233), .B(n2397), .Z(n3236) );
  XNOR U2861 ( .A(p_input[3915]), .B(n3237), .Z(n2397) );
  AND U2862 ( .A(n186), .B(n3238), .Z(n3237) );
  XOR U2863 ( .A(p_input[3947]), .B(p_input[3915]), .Z(n3238) );
  XNOR U2864 ( .A(n2394), .B(n3233), .Z(n3235) );
  XOR U2865 ( .A(n3239), .B(n3240), .Z(n2394) );
  AND U2866 ( .A(n183), .B(n3241), .Z(n3240) );
  XOR U2867 ( .A(p_input[3883]), .B(p_input[3851]), .Z(n3241) );
  XOR U2868 ( .A(n3242), .B(n3243), .Z(n3233) );
  AND U2869 ( .A(n3244), .B(n3245), .Z(n3243) );
  XOR U2870 ( .A(n3242), .B(n2409), .Z(n3245) );
  XNOR U2871 ( .A(p_input[3914]), .B(n3246), .Z(n2409) );
  AND U2872 ( .A(n186), .B(n3247), .Z(n3246) );
  XOR U2873 ( .A(p_input[3946]), .B(p_input[3914]), .Z(n3247) );
  XNOR U2874 ( .A(n2406), .B(n3242), .Z(n3244) );
  XOR U2875 ( .A(n3248), .B(n3249), .Z(n2406) );
  AND U2876 ( .A(n183), .B(n3250), .Z(n3249) );
  XOR U2877 ( .A(p_input[3882]), .B(p_input[3850]), .Z(n3250) );
  XOR U2878 ( .A(n3251), .B(n3252), .Z(n3242) );
  AND U2879 ( .A(n3253), .B(n3254), .Z(n3252) );
  XOR U2880 ( .A(n3251), .B(n2421), .Z(n3254) );
  XNOR U2881 ( .A(p_input[3913]), .B(n3255), .Z(n2421) );
  AND U2882 ( .A(n186), .B(n3256), .Z(n3255) );
  XOR U2883 ( .A(p_input[3945]), .B(p_input[3913]), .Z(n3256) );
  XNOR U2884 ( .A(n2418), .B(n3251), .Z(n3253) );
  XOR U2885 ( .A(n3257), .B(n3258), .Z(n2418) );
  AND U2886 ( .A(n183), .B(n3259), .Z(n3258) );
  XOR U2887 ( .A(p_input[3881]), .B(p_input[3849]), .Z(n3259) );
  XOR U2888 ( .A(n3260), .B(n3261), .Z(n3251) );
  AND U2889 ( .A(n3262), .B(n3263), .Z(n3261) );
  XOR U2890 ( .A(n3260), .B(n2433), .Z(n3263) );
  XNOR U2891 ( .A(p_input[3912]), .B(n3264), .Z(n2433) );
  AND U2892 ( .A(n186), .B(n3265), .Z(n3264) );
  XOR U2893 ( .A(p_input[3944]), .B(p_input[3912]), .Z(n3265) );
  XNOR U2894 ( .A(n2430), .B(n3260), .Z(n3262) );
  XOR U2895 ( .A(n3266), .B(n3267), .Z(n2430) );
  AND U2896 ( .A(n183), .B(n3268), .Z(n3267) );
  XOR U2897 ( .A(p_input[3880]), .B(p_input[3848]), .Z(n3268) );
  XOR U2898 ( .A(n3269), .B(n3270), .Z(n3260) );
  AND U2899 ( .A(n3271), .B(n3272), .Z(n3270) );
  XOR U2900 ( .A(n3269), .B(n2445), .Z(n3272) );
  XNOR U2901 ( .A(p_input[3911]), .B(n3273), .Z(n2445) );
  AND U2902 ( .A(n186), .B(n3274), .Z(n3273) );
  XOR U2903 ( .A(p_input[3943]), .B(p_input[3911]), .Z(n3274) );
  XNOR U2904 ( .A(n2442), .B(n3269), .Z(n3271) );
  XOR U2905 ( .A(n3275), .B(n3276), .Z(n2442) );
  AND U2906 ( .A(n183), .B(n3277), .Z(n3276) );
  XOR U2907 ( .A(p_input[3879]), .B(p_input[3847]), .Z(n3277) );
  XOR U2908 ( .A(n3278), .B(n3279), .Z(n3269) );
  AND U2909 ( .A(n3280), .B(n3281), .Z(n3279) );
  XOR U2910 ( .A(n3278), .B(n2457), .Z(n3281) );
  XNOR U2911 ( .A(p_input[3910]), .B(n3282), .Z(n2457) );
  AND U2912 ( .A(n186), .B(n3283), .Z(n3282) );
  XOR U2913 ( .A(p_input[3942]), .B(p_input[3910]), .Z(n3283) );
  XNOR U2914 ( .A(n2454), .B(n3278), .Z(n3280) );
  XOR U2915 ( .A(n3284), .B(n3285), .Z(n2454) );
  AND U2916 ( .A(n183), .B(n3286), .Z(n3285) );
  XOR U2917 ( .A(p_input[3878]), .B(p_input[3846]), .Z(n3286) );
  XOR U2918 ( .A(n3287), .B(n3288), .Z(n3278) );
  AND U2919 ( .A(n3289), .B(n3290), .Z(n3288) );
  XOR U2920 ( .A(n3287), .B(n2469), .Z(n3290) );
  XNOR U2921 ( .A(p_input[3909]), .B(n3291), .Z(n2469) );
  AND U2922 ( .A(n186), .B(n3292), .Z(n3291) );
  XOR U2923 ( .A(p_input[3941]), .B(p_input[3909]), .Z(n3292) );
  XNOR U2924 ( .A(n2466), .B(n3287), .Z(n3289) );
  XOR U2925 ( .A(n3293), .B(n3294), .Z(n2466) );
  AND U2926 ( .A(n183), .B(n3295), .Z(n3294) );
  XOR U2927 ( .A(p_input[3877]), .B(p_input[3845]), .Z(n3295) );
  XOR U2928 ( .A(n3296), .B(n3297), .Z(n3287) );
  AND U2929 ( .A(n3298), .B(n3299), .Z(n3297) );
  XOR U2930 ( .A(n3296), .B(n2481), .Z(n3299) );
  XNOR U2931 ( .A(p_input[3908]), .B(n3300), .Z(n2481) );
  AND U2932 ( .A(n186), .B(n3301), .Z(n3300) );
  XOR U2933 ( .A(p_input[3940]), .B(p_input[3908]), .Z(n3301) );
  XNOR U2934 ( .A(n2478), .B(n3296), .Z(n3298) );
  XOR U2935 ( .A(n3302), .B(n3303), .Z(n2478) );
  AND U2936 ( .A(n183), .B(n3304), .Z(n3303) );
  XOR U2937 ( .A(p_input[3876]), .B(p_input[3844]), .Z(n3304) );
  XOR U2938 ( .A(n3305), .B(n3306), .Z(n3296) );
  AND U2939 ( .A(n3307), .B(n3308), .Z(n3306) );
  XOR U2940 ( .A(n3305), .B(n2493), .Z(n3308) );
  XNOR U2941 ( .A(p_input[3907]), .B(n3309), .Z(n2493) );
  AND U2942 ( .A(n186), .B(n3310), .Z(n3309) );
  XOR U2943 ( .A(p_input[3939]), .B(p_input[3907]), .Z(n3310) );
  XNOR U2944 ( .A(n2490), .B(n3305), .Z(n3307) );
  XOR U2945 ( .A(n3311), .B(n3312), .Z(n2490) );
  AND U2946 ( .A(n183), .B(n3313), .Z(n3312) );
  XOR U2947 ( .A(p_input[3875]), .B(p_input[3843]), .Z(n3313) );
  XOR U2948 ( .A(n3314), .B(n3315), .Z(n3305) );
  AND U2949 ( .A(n3316), .B(n3317), .Z(n3315) );
  XOR U2950 ( .A(n2505), .B(n3314), .Z(n3317) );
  XNOR U2951 ( .A(p_input[3906]), .B(n3318), .Z(n2505) );
  AND U2952 ( .A(n186), .B(n3319), .Z(n3318) );
  XOR U2953 ( .A(p_input[3938]), .B(p_input[3906]), .Z(n3319) );
  XNOR U2954 ( .A(n3314), .B(n2502), .Z(n3316) );
  XOR U2955 ( .A(n3320), .B(n3321), .Z(n2502) );
  AND U2956 ( .A(n183), .B(n3322), .Z(n3321) );
  XOR U2957 ( .A(p_input[3874]), .B(p_input[3842]), .Z(n3322) );
  XOR U2958 ( .A(n3323), .B(n3324), .Z(n3314) );
  AND U2959 ( .A(n3325), .B(n3326), .Z(n3324) );
  XNOR U2960 ( .A(n3327), .B(n2518), .Z(n3326) );
  XNOR U2961 ( .A(p_input[3905]), .B(n3328), .Z(n2518) );
  AND U2962 ( .A(n186), .B(n3329), .Z(n3328) );
  XNOR U2963 ( .A(p_input[3937]), .B(n3330), .Z(n3329) );
  IV U2964 ( .A(p_input[3905]), .Z(n3330) );
  XNOR U2965 ( .A(n2515), .B(n3323), .Z(n3325) );
  XNOR U2966 ( .A(p_input[3841]), .B(n3331), .Z(n2515) );
  AND U2967 ( .A(n183), .B(n3332), .Z(n3331) );
  XOR U2968 ( .A(p_input[3873]), .B(p_input[3841]), .Z(n3332) );
  IV U2969 ( .A(n3327), .Z(n3323) );
  AND U2970 ( .A(n3053), .B(n3056), .Z(n3327) );
  XOR U2971 ( .A(p_input[3904]), .B(n3333), .Z(n3056) );
  AND U2972 ( .A(n186), .B(n3334), .Z(n3333) );
  XOR U2973 ( .A(p_input[3936]), .B(p_input[3904]), .Z(n3334) );
  XOR U2974 ( .A(n3335), .B(n3336), .Z(n186) );
  AND U2975 ( .A(n3337), .B(n3338), .Z(n3336) );
  XNOR U2976 ( .A(p_input[3967]), .B(n3335), .Z(n3338) );
  XOR U2977 ( .A(n3335), .B(p_input[3935]), .Z(n3337) );
  XOR U2978 ( .A(n3339), .B(n3340), .Z(n3335) );
  AND U2979 ( .A(n3341), .B(n3342), .Z(n3340) );
  XNOR U2980 ( .A(p_input[3966]), .B(n3339), .Z(n3342) );
  XOR U2981 ( .A(n3339), .B(p_input[3934]), .Z(n3341) );
  XOR U2982 ( .A(n3343), .B(n3344), .Z(n3339) );
  AND U2983 ( .A(n3345), .B(n3346), .Z(n3344) );
  XNOR U2984 ( .A(p_input[3965]), .B(n3343), .Z(n3346) );
  XOR U2985 ( .A(n3343), .B(p_input[3933]), .Z(n3345) );
  XOR U2986 ( .A(n3347), .B(n3348), .Z(n3343) );
  AND U2987 ( .A(n3349), .B(n3350), .Z(n3348) );
  XNOR U2988 ( .A(p_input[3964]), .B(n3347), .Z(n3350) );
  XOR U2989 ( .A(n3347), .B(p_input[3932]), .Z(n3349) );
  XOR U2990 ( .A(n3351), .B(n3352), .Z(n3347) );
  AND U2991 ( .A(n3353), .B(n3354), .Z(n3352) );
  XNOR U2992 ( .A(p_input[3963]), .B(n3351), .Z(n3354) );
  XOR U2993 ( .A(n3351), .B(p_input[3931]), .Z(n3353) );
  XOR U2994 ( .A(n3355), .B(n3356), .Z(n3351) );
  AND U2995 ( .A(n3357), .B(n3358), .Z(n3356) );
  XNOR U2996 ( .A(p_input[3962]), .B(n3355), .Z(n3358) );
  XOR U2997 ( .A(n3355), .B(p_input[3930]), .Z(n3357) );
  XOR U2998 ( .A(n3359), .B(n3360), .Z(n3355) );
  AND U2999 ( .A(n3361), .B(n3362), .Z(n3360) );
  XNOR U3000 ( .A(p_input[3961]), .B(n3359), .Z(n3362) );
  XOR U3001 ( .A(n3359), .B(p_input[3929]), .Z(n3361) );
  XOR U3002 ( .A(n3363), .B(n3364), .Z(n3359) );
  AND U3003 ( .A(n3365), .B(n3366), .Z(n3364) );
  XNOR U3004 ( .A(p_input[3960]), .B(n3363), .Z(n3366) );
  XOR U3005 ( .A(n3363), .B(p_input[3928]), .Z(n3365) );
  XOR U3006 ( .A(n3367), .B(n3368), .Z(n3363) );
  AND U3007 ( .A(n3369), .B(n3370), .Z(n3368) );
  XNOR U3008 ( .A(p_input[3959]), .B(n3367), .Z(n3370) );
  XOR U3009 ( .A(n3367), .B(p_input[3927]), .Z(n3369) );
  XOR U3010 ( .A(n3371), .B(n3372), .Z(n3367) );
  AND U3011 ( .A(n3373), .B(n3374), .Z(n3372) );
  XNOR U3012 ( .A(p_input[3958]), .B(n3371), .Z(n3374) );
  XOR U3013 ( .A(n3371), .B(p_input[3926]), .Z(n3373) );
  XOR U3014 ( .A(n3375), .B(n3376), .Z(n3371) );
  AND U3015 ( .A(n3377), .B(n3378), .Z(n3376) );
  XNOR U3016 ( .A(p_input[3957]), .B(n3375), .Z(n3378) );
  XOR U3017 ( .A(n3375), .B(p_input[3925]), .Z(n3377) );
  XOR U3018 ( .A(n3379), .B(n3380), .Z(n3375) );
  AND U3019 ( .A(n3381), .B(n3382), .Z(n3380) );
  XNOR U3020 ( .A(p_input[3956]), .B(n3379), .Z(n3382) );
  XOR U3021 ( .A(n3379), .B(p_input[3924]), .Z(n3381) );
  XOR U3022 ( .A(n3383), .B(n3384), .Z(n3379) );
  AND U3023 ( .A(n3385), .B(n3386), .Z(n3384) );
  XNOR U3024 ( .A(p_input[3955]), .B(n3383), .Z(n3386) );
  XOR U3025 ( .A(n3383), .B(p_input[3923]), .Z(n3385) );
  XOR U3026 ( .A(n3387), .B(n3388), .Z(n3383) );
  AND U3027 ( .A(n3389), .B(n3390), .Z(n3388) );
  XNOR U3028 ( .A(p_input[3954]), .B(n3387), .Z(n3390) );
  XOR U3029 ( .A(n3387), .B(p_input[3922]), .Z(n3389) );
  XOR U3030 ( .A(n3391), .B(n3392), .Z(n3387) );
  AND U3031 ( .A(n3393), .B(n3394), .Z(n3392) );
  XNOR U3032 ( .A(p_input[3953]), .B(n3391), .Z(n3394) );
  XOR U3033 ( .A(n3391), .B(p_input[3921]), .Z(n3393) );
  XOR U3034 ( .A(n3395), .B(n3396), .Z(n3391) );
  AND U3035 ( .A(n3397), .B(n3398), .Z(n3396) );
  XNOR U3036 ( .A(p_input[3952]), .B(n3395), .Z(n3398) );
  XOR U3037 ( .A(n3395), .B(p_input[3920]), .Z(n3397) );
  XOR U3038 ( .A(n3399), .B(n3400), .Z(n3395) );
  AND U3039 ( .A(n3401), .B(n3402), .Z(n3400) );
  XNOR U3040 ( .A(p_input[3951]), .B(n3399), .Z(n3402) );
  XOR U3041 ( .A(n3399), .B(p_input[3919]), .Z(n3401) );
  XOR U3042 ( .A(n3403), .B(n3404), .Z(n3399) );
  AND U3043 ( .A(n3405), .B(n3406), .Z(n3404) );
  XNOR U3044 ( .A(p_input[3950]), .B(n3403), .Z(n3406) );
  XOR U3045 ( .A(n3403), .B(p_input[3918]), .Z(n3405) );
  XOR U3046 ( .A(n3407), .B(n3408), .Z(n3403) );
  AND U3047 ( .A(n3409), .B(n3410), .Z(n3408) );
  XNOR U3048 ( .A(p_input[3949]), .B(n3407), .Z(n3410) );
  XOR U3049 ( .A(n3407), .B(p_input[3917]), .Z(n3409) );
  XOR U3050 ( .A(n3411), .B(n3412), .Z(n3407) );
  AND U3051 ( .A(n3413), .B(n3414), .Z(n3412) );
  XNOR U3052 ( .A(p_input[3948]), .B(n3411), .Z(n3414) );
  XOR U3053 ( .A(n3411), .B(p_input[3916]), .Z(n3413) );
  XOR U3054 ( .A(n3415), .B(n3416), .Z(n3411) );
  AND U3055 ( .A(n3417), .B(n3418), .Z(n3416) );
  XNOR U3056 ( .A(p_input[3947]), .B(n3415), .Z(n3418) );
  XOR U3057 ( .A(n3415), .B(p_input[3915]), .Z(n3417) );
  XOR U3058 ( .A(n3419), .B(n3420), .Z(n3415) );
  AND U3059 ( .A(n3421), .B(n3422), .Z(n3420) );
  XNOR U3060 ( .A(p_input[3946]), .B(n3419), .Z(n3422) );
  XOR U3061 ( .A(n3419), .B(p_input[3914]), .Z(n3421) );
  XOR U3062 ( .A(n3423), .B(n3424), .Z(n3419) );
  AND U3063 ( .A(n3425), .B(n3426), .Z(n3424) );
  XNOR U3064 ( .A(p_input[3945]), .B(n3423), .Z(n3426) );
  XOR U3065 ( .A(n3423), .B(p_input[3913]), .Z(n3425) );
  XOR U3066 ( .A(n3427), .B(n3428), .Z(n3423) );
  AND U3067 ( .A(n3429), .B(n3430), .Z(n3428) );
  XNOR U3068 ( .A(p_input[3944]), .B(n3427), .Z(n3430) );
  XOR U3069 ( .A(n3427), .B(p_input[3912]), .Z(n3429) );
  XOR U3070 ( .A(n3431), .B(n3432), .Z(n3427) );
  AND U3071 ( .A(n3433), .B(n3434), .Z(n3432) );
  XNOR U3072 ( .A(p_input[3943]), .B(n3431), .Z(n3434) );
  XOR U3073 ( .A(n3431), .B(p_input[3911]), .Z(n3433) );
  XOR U3074 ( .A(n3435), .B(n3436), .Z(n3431) );
  AND U3075 ( .A(n3437), .B(n3438), .Z(n3436) );
  XNOR U3076 ( .A(p_input[3942]), .B(n3435), .Z(n3438) );
  XOR U3077 ( .A(n3435), .B(p_input[3910]), .Z(n3437) );
  XOR U3078 ( .A(n3439), .B(n3440), .Z(n3435) );
  AND U3079 ( .A(n3441), .B(n3442), .Z(n3440) );
  XNOR U3080 ( .A(p_input[3941]), .B(n3439), .Z(n3442) );
  XOR U3081 ( .A(n3439), .B(p_input[3909]), .Z(n3441) );
  XOR U3082 ( .A(n3443), .B(n3444), .Z(n3439) );
  AND U3083 ( .A(n3445), .B(n3446), .Z(n3444) );
  XNOR U3084 ( .A(p_input[3940]), .B(n3443), .Z(n3446) );
  XOR U3085 ( .A(n3443), .B(p_input[3908]), .Z(n3445) );
  XOR U3086 ( .A(n3447), .B(n3448), .Z(n3443) );
  AND U3087 ( .A(n3449), .B(n3450), .Z(n3448) );
  XNOR U3088 ( .A(p_input[3939]), .B(n3447), .Z(n3450) );
  XOR U3089 ( .A(n3447), .B(p_input[3907]), .Z(n3449) );
  XOR U3090 ( .A(n3451), .B(n3452), .Z(n3447) );
  AND U3091 ( .A(n3453), .B(n3454), .Z(n3452) );
  XNOR U3092 ( .A(p_input[3938]), .B(n3451), .Z(n3454) );
  XOR U3093 ( .A(n3451), .B(p_input[3906]), .Z(n3453) );
  XNOR U3094 ( .A(n3455), .B(n3456), .Z(n3451) );
  AND U3095 ( .A(n3457), .B(n3458), .Z(n3456) );
  XOR U3096 ( .A(p_input[3937]), .B(n3455), .Z(n3458) );
  XNOR U3097 ( .A(p_input[3905]), .B(n3455), .Z(n3457) );
  AND U3098 ( .A(p_input[3936]), .B(n3459), .Z(n3455) );
  IV U3099 ( .A(p_input[3904]), .Z(n3459) );
  XNOR U3100 ( .A(p_input[3840]), .B(n3460), .Z(n3053) );
  AND U3101 ( .A(n183), .B(n3461), .Z(n3460) );
  XOR U3102 ( .A(p_input[3872]), .B(p_input[3840]), .Z(n3461) );
  XOR U3103 ( .A(n3462), .B(n3463), .Z(n183) );
  AND U3104 ( .A(n3464), .B(n3465), .Z(n3463) );
  XNOR U3105 ( .A(p_input[3903]), .B(n3462), .Z(n3465) );
  XOR U3106 ( .A(n3462), .B(p_input[3871]), .Z(n3464) );
  XOR U3107 ( .A(n3466), .B(n3467), .Z(n3462) );
  AND U3108 ( .A(n3468), .B(n3469), .Z(n3467) );
  XNOR U3109 ( .A(p_input[3902]), .B(n3466), .Z(n3469) );
  XNOR U3110 ( .A(n3466), .B(n3068), .Z(n3468) );
  IV U3111 ( .A(p_input[3870]), .Z(n3068) );
  XOR U3112 ( .A(n3470), .B(n3471), .Z(n3466) );
  AND U3113 ( .A(n3472), .B(n3473), .Z(n3471) );
  XNOR U3114 ( .A(p_input[3901]), .B(n3470), .Z(n3473) );
  XNOR U3115 ( .A(n3470), .B(n3077), .Z(n3472) );
  IV U3116 ( .A(p_input[3869]), .Z(n3077) );
  XOR U3117 ( .A(n3474), .B(n3475), .Z(n3470) );
  AND U3118 ( .A(n3476), .B(n3477), .Z(n3475) );
  XNOR U3119 ( .A(p_input[3900]), .B(n3474), .Z(n3477) );
  XNOR U3120 ( .A(n3474), .B(n3086), .Z(n3476) );
  IV U3121 ( .A(p_input[3868]), .Z(n3086) );
  XOR U3122 ( .A(n3478), .B(n3479), .Z(n3474) );
  AND U3123 ( .A(n3480), .B(n3481), .Z(n3479) );
  XNOR U3124 ( .A(p_input[3899]), .B(n3478), .Z(n3481) );
  XNOR U3125 ( .A(n3478), .B(n3095), .Z(n3480) );
  IV U3126 ( .A(p_input[3867]), .Z(n3095) );
  XOR U3127 ( .A(n3482), .B(n3483), .Z(n3478) );
  AND U3128 ( .A(n3484), .B(n3485), .Z(n3483) );
  XNOR U3129 ( .A(p_input[3898]), .B(n3482), .Z(n3485) );
  XNOR U3130 ( .A(n3482), .B(n3104), .Z(n3484) );
  IV U3131 ( .A(p_input[3866]), .Z(n3104) );
  XOR U3132 ( .A(n3486), .B(n3487), .Z(n3482) );
  AND U3133 ( .A(n3488), .B(n3489), .Z(n3487) );
  XNOR U3134 ( .A(p_input[3897]), .B(n3486), .Z(n3489) );
  XNOR U3135 ( .A(n3486), .B(n3113), .Z(n3488) );
  IV U3136 ( .A(p_input[3865]), .Z(n3113) );
  XOR U3137 ( .A(n3490), .B(n3491), .Z(n3486) );
  AND U3138 ( .A(n3492), .B(n3493), .Z(n3491) );
  XNOR U3139 ( .A(p_input[3896]), .B(n3490), .Z(n3493) );
  XNOR U3140 ( .A(n3490), .B(n3122), .Z(n3492) );
  IV U3141 ( .A(p_input[3864]), .Z(n3122) );
  XOR U3142 ( .A(n3494), .B(n3495), .Z(n3490) );
  AND U3143 ( .A(n3496), .B(n3497), .Z(n3495) );
  XNOR U3144 ( .A(p_input[3895]), .B(n3494), .Z(n3497) );
  XNOR U3145 ( .A(n3494), .B(n3131), .Z(n3496) );
  IV U3146 ( .A(p_input[3863]), .Z(n3131) );
  XOR U3147 ( .A(n3498), .B(n3499), .Z(n3494) );
  AND U3148 ( .A(n3500), .B(n3501), .Z(n3499) );
  XNOR U3149 ( .A(p_input[3894]), .B(n3498), .Z(n3501) );
  XNOR U3150 ( .A(n3498), .B(n3140), .Z(n3500) );
  IV U3151 ( .A(p_input[3862]), .Z(n3140) );
  XOR U3152 ( .A(n3502), .B(n3503), .Z(n3498) );
  AND U3153 ( .A(n3504), .B(n3505), .Z(n3503) );
  XNOR U3154 ( .A(p_input[3893]), .B(n3502), .Z(n3505) );
  XNOR U3155 ( .A(n3502), .B(n3149), .Z(n3504) );
  IV U3156 ( .A(p_input[3861]), .Z(n3149) );
  XOR U3157 ( .A(n3506), .B(n3507), .Z(n3502) );
  AND U3158 ( .A(n3508), .B(n3509), .Z(n3507) );
  XNOR U3159 ( .A(p_input[3892]), .B(n3506), .Z(n3509) );
  XNOR U3160 ( .A(n3506), .B(n3158), .Z(n3508) );
  IV U3161 ( .A(p_input[3860]), .Z(n3158) );
  XOR U3162 ( .A(n3510), .B(n3511), .Z(n3506) );
  AND U3163 ( .A(n3512), .B(n3513), .Z(n3511) );
  XNOR U3164 ( .A(p_input[3891]), .B(n3510), .Z(n3513) );
  XNOR U3165 ( .A(n3510), .B(n3167), .Z(n3512) );
  IV U3166 ( .A(p_input[3859]), .Z(n3167) );
  XOR U3167 ( .A(n3514), .B(n3515), .Z(n3510) );
  AND U3168 ( .A(n3516), .B(n3517), .Z(n3515) );
  XNOR U3169 ( .A(p_input[3890]), .B(n3514), .Z(n3517) );
  XNOR U3170 ( .A(n3514), .B(n3176), .Z(n3516) );
  IV U3171 ( .A(p_input[3858]), .Z(n3176) );
  XOR U3172 ( .A(n3518), .B(n3519), .Z(n3514) );
  AND U3173 ( .A(n3520), .B(n3521), .Z(n3519) );
  XNOR U3174 ( .A(p_input[3889]), .B(n3518), .Z(n3521) );
  XNOR U3175 ( .A(n3518), .B(n3185), .Z(n3520) );
  IV U3176 ( .A(p_input[3857]), .Z(n3185) );
  XOR U3177 ( .A(n3522), .B(n3523), .Z(n3518) );
  AND U3178 ( .A(n3524), .B(n3525), .Z(n3523) );
  XNOR U3179 ( .A(p_input[3888]), .B(n3522), .Z(n3525) );
  XNOR U3180 ( .A(n3522), .B(n3194), .Z(n3524) );
  IV U3181 ( .A(p_input[3856]), .Z(n3194) );
  XOR U3182 ( .A(n3526), .B(n3527), .Z(n3522) );
  AND U3183 ( .A(n3528), .B(n3529), .Z(n3527) );
  XNOR U3184 ( .A(p_input[3887]), .B(n3526), .Z(n3529) );
  XNOR U3185 ( .A(n3526), .B(n3203), .Z(n3528) );
  IV U3186 ( .A(p_input[3855]), .Z(n3203) );
  XOR U3187 ( .A(n3530), .B(n3531), .Z(n3526) );
  AND U3188 ( .A(n3532), .B(n3533), .Z(n3531) );
  XNOR U3189 ( .A(p_input[3886]), .B(n3530), .Z(n3533) );
  XNOR U3190 ( .A(n3530), .B(n3212), .Z(n3532) );
  IV U3191 ( .A(p_input[3854]), .Z(n3212) );
  XOR U3192 ( .A(n3534), .B(n3535), .Z(n3530) );
  AND U3193 ( .A(n3536), .B(n3537), .Z(n3535) );
  XNOR U3194 ( .A(p_input[3885]), .B(n3534), .Z(n3537) );
  XNOR U3195 ( .A(n3534), .B(n3221), .Z(n3536) );
  IV U3196 ( .A(p_input[3853]), .Z(n3221) );
  XOR U3197 ( .A(n3538), .B(n3539), .Z(n3534) );
  AND U3198 ( .A(n3540), .B(n3541), .Z(n3539) );
  XNOR U3199 ( .A(p_input[3884]), .B(n3538), .Z(n3541) );
  XNOR U3200 ( .A(n3538), .B(n3230), .Z(n3540) );
  IV U3201 ( .A(p_input[3852]), .Z(n3230) );
  XOR U3202 ( .A(n3542), .B(n3543), .Z(n3538) );
  AND U3203 ( .A(n3544), .B(n3545), .Z(n3543) );
  XNOR U3204 ( .A(p_input[3883]), .B(n3542), .Z(n3545) );
  XNOR U3205 ( .A(n3542), .B(n3239), .Z(n3544) );
  IV U3206 ( .A(p_input[3851]), .Z(n3239) );
  XOR U3207 ( .A(n3546), .B(n3547), .Z(n3542) );
  AND U3208 ( .A(n3548), .B(n3549), .Z(n3547) );
  XNOR U3209 ( .A(p_input[3882]), .B(n3546), .Z(n3549) );
  XNOR U3210 ( .A(n3546), .B(n3248), .Z(n3548) );
  IV U3211 ( .A(p_input[3850]), .Z(n3248) );
  XOR U3212 ( .A(n3550), .B(n3551), .Z(n3546) );
  AND U3213 ( .A(n3552), .B(n3553), .Z(n3551) );
  XNOR U3214 ( .A(p_input[3881]), .B(n3550), .Z(n3553) );
  XNOR U3215 ( .A(n3550), .B(n3257), .Z(n3552) );
  IV U3216 ( .A(p_input[3849]), .Z(n3257) );
  XOR U3217 ( .A(n3554), .B(n3555), .Z(n3550) );
  AND U3218 ( .A(n3556), .B(n3557), .Z(n3555) );
  XNOR U3219 ( .A(p_input[3880]), .B(n3554), .Z(n3557) );
  XNOR U3220 ( .A(n3554), .B(n3266), .Z(n3556) );
  IV U3221 ( .A(p_input[3848]), .Z(n3266) );
  XOR U3222 ( .A(n3558), .B(n3559), .Z(n3554) );
  AND U3223 ( .A(n3560), .B(n3561), .Z(n3559) );
  XNOR U3224 ( .A(p_input[3879]), .B(n3558), .Z(n3561) );
  XNOR U3225 ( .A(n3558), .B(n3275), .Z(n3560) );
  IV U3226 ( .A(p_input[3847]), .Z(n3275) );
  XOR U3227 ( .A(n3562), .B(n3563), .Z(n3558) );
  AND U3228 ( .A(n3564), .B(n3565), .Z(n3563) );
  XNOR U3229 ( .A(p_input[3878]), .B(n3562), .Z(n3565) );
  XNOR U3230 ( .A(n3562), .B(n3284), .Z(n3564) );
  IV U3231 ( .A(p_input[3846]), .Z(n3284) );
  XOR U3232 ( .A(n3566), .B(n3567), .Z(n3562) );
  AND U3233 ( .A(n3568), .B(n3569), .Z(n3567) );
  XNOR U3234 ( .A(p_input[3877]), .B(n3566), .Z(n3569) );
  XNOR U3235 ( .A(n3566), .B(n3293), .Z(n3568) );
  IV U3236 ( .A(p_input[3845]), .Z(n3293) );
  XOR U3237 ( .A(n3570), .B(n3571), .Z(n3566) );
  AND U3238 ( .A(n3572), .B(n3573), .Z(n3571) );
  XNOR U3239 ( .A(p_input[3876]), .B(n3570), .Z(n3573) );
  XNOR U3240 ( .A(n3570), .B(n3302), .Z(n3572) );
  IV U3241 ( .A(p_input[3844]), .Z(n3302) );
  XOR U3242 ( .A(n3574), .B(n3575), .Z(n3570) );
  AND U3243 ( .A(n3576), .B(n3577), .Z(n3575) );
  XNOR U3244 ( .A(p_input[3875]), .B(n3574), .Z(n3577) );
  XNOR U3245 ( .A(n3574), .B(n3311), .Z(n3576) );
  IV U3246 ( .A(p_input[3843]), .Z(n3311) );
  XOR U3247 ( .A(n3578), .B(n3579), .Z(n3574) );
  AND U3248 ( .A(n3580), .B(n3581), .Z(n3579) );
  XNOR U3249 ( .A(p_input[3874]), .B(n3578), .Z(n3581) );
  XNOR U3250 ( .A(n3578), .B(n3320), .Z(n3580) );
  IV U3251 ( .A(p_input[3842]), .Z(n3320) );
  XNOR U3252 ( .A(n3582), .B(n3583), .Z(n3578) );
  AND U3253 ( .A(n3584), .B(n3585), .Z(n3583) );
  XOR U3254 ( .A(p_input[3873]), .B(n3582), .Z(n3585) );
  XNOR U3255 ( .A(p_input[3841]), .B(n3582), .Z(n3584) );
  AND U3256 ( .A(p_input[3872]), .B(n3586), .Z(n3582) );
  IV U3257 ( .A(p_input[3840]), .Z(n3586) );
  XOR U3258 ( .A(n3587), .B(n3588), .Z(n1765) );
  AND U3259 ( .A(n488), .B(n3589), .Z(n3588) );
  XNOR U3260 ( .A(n3590), .B(n3587), .Z(n3589) );
  XOR U3261 ( .A(n3591), .B(n3592), .Z(n488) );
  AND U3262 ( .A(n3593), .B(n3594), .Z(n3592) );
  XOR U3263 ( .A(n3591), .B(n1780), .Z(n3594) );
  XNOR U3264 ( .A(n3595), .B(n3596), .Z(n1780) );
  AND U3265 ( .A(n3597), .B(n310), .Z(n3596) );
  AND U3266 ( .A(n3595), .B(n3598), .Z(n3597) );
  XNOR U3267 ( .A(n1777), .B(n3591), .Z(n3593) );
  XOR U3268 ( .A(n3599), .B(n3600), .Z(n1777) );
  AND U3269 ( .A(n3601), .B(n307), .Z(n3600) );
  NOR U3270 ( .A(n3599), .B(n3602), .Z(n3601) );
  XOR U3271 ( .A(n3603), .B(n3604), .Z(n3591) );
  AND U3272 ( .A(n3605), .B(n3606), .Z(n3604) );
  XOR U3273 ( .A(n3603), .B(n1792), .Z(n3606) );
  XOR U3274 ( .A(n3607), .B(n3608), .Z(n1792) );
  AND U3275 ( .A(n310), .B(n3609), .Z(n3608) );
  XOR U3276 ( .A(n3610), .B(n3607), .Z(n3609) );
  XNOR U3277 ( .A(n1789), .B(n3603), .Z(n3605) );
  XOR U3278 ( .A(n3611), .B(n3612), .Z(n1789) );
  AND U3279 ( .A(n307), .B(n3613), .Z(n3612) );
  XOR U3280 ( .A(n3614), .B(n3611), .Z(n3613) );
  XOR U3281 ( .A(n3615), .B(n3616), .Z(n3603) );
  AND U3282 ( .A(n3617), .B(n3618), .Z(n3616) );
  XOR U3283 ( .A(n3615), .B(n1804), .Z(n3618) );
  XOR U3284 ( .A(n3619), .B(n3620), .Z(n1804) );
  AND U3285 ( .A(n310), .B(n3621), .Z(n3620) );
  XOR U3286 ( .A(n3622), .B(n3619), .Z(n3621) );
  XNOR U3287 ( .A(n1801), .B(n3615), .Z(n3617) );
  XOR U3288 ( .A(n3623), .B(n3624), .Z(n1801) );
  AND U3289 ( .A(n307), .B(n3625), .Z(n3624) );
  XOR U3290 ( .A(n3626), .B(n3623), .Z(n3625) );
  XOR U3291 ( .A(n3627), .B(n3628), .Z(n3615) );
  AND U3292 ( .A(n3629), .B(n3630), .Z(n3628) );
  XOR U3293 ( .A(n3627), .B(n1816), .Z(n3630) );
  XOR U3294 ( .A(n3631), .B(n3632), .Z(n1816) );
  AND U3295 ( .A(n310), .B(n3633), .Z(n3632) );
  XOR U3296 ( .A(n3634), .B(n3631), .Z(n3633) );
  XNOR U3297 ( .A(n1813), .B(n3627), .Z(n3629) );
  XOR U3298 ( .A(n3635), .B(n3636), .Z(n1813) );
  AND U3299 ( .A(n307), .B(n3637), .Z(n3636) );
  XOR U3300 ( .A(n3638), .B(n3635), .Z(n3637) );
  XOR U3301 ( .A(n3639), .B(n3640), .Z(n3627) );
  AND U3302 ( .A(n3641), .B(n3642), .Z(n3640) );
  XOR U3303 ( .A(n3639), .B(n1828), .Z(n3642) );
  XOR U3304 ( .A(n3643), .B(n3644), .Z(n1828) );
  AND U3305 ( .A(n310), .B(n3645), .Z(n3644) );
  XOR U3306 ( .A(n3646), .B(n3643), .Z(n3645) );
  XNOR U3307 ( .A(n1825), .B(n3639), .Z(n3641) );
  XOR U3308 ( .A(n3647), .B(n3648), .Z(n1825) );
  AND U3309 ( .A(n307), .B(n3649), .Z(n3648) );
  XOR U3310 ( .A(n3650), .B(n3647), .Z(n3649) );
  XOR U3311 ( .A(n3651), .B(n3652), .Z(n3639) );
  AND U3312 ( .A(n3653), .B(n3654), .Z(n3652) );
  XOR U3313 ( .A(n3651), .B(n1840), .Z(n3654) );
  XOR U3314 ( .A(n3655), .B(n3656), .Z(n1840) );
  AND U3315 ( .A(n310), .B(n3657), .Z(n3656) );
  XOR U3316 ( .A(n3658), .B(n3655), .Z(n3657) );
  XNOR U3317 ( .A(n1837), .B(n3651), .Z(n3653) );
  XOR U3318 ( .A(n3659), .B(n3660), .Z(n1837) );
  AND U3319 ( .A(n307), .B(n3661), .Z(n3660) );
  XOR U3320 ( .A(n3662), .B(n3659), .Z(n3661) );
  XOR U3321 ( .A(n3663), .B(n3664), .Z(n3651) );
  AND U3322 ( .A(n3665), .B(n3666), .Z(n3664) );
  XOR U3323 ( .A(n3663), .B(n1852), .Z(n3666) );
  XOR U3324 ( .A(n3667), .B(n3668), .Z(n1852) );
  AND U3325 ( .A(n310), .B(n3669), .Z(n3668) );
  XOR U3326 ( .A(n3670), .B(n3667), .Z(n3669) );
  XNOR U3327 ( .A(n1849), .B(n3663), .Z(n3665) );
  XOR U3328 ( .A(n3671), .B(n3672), .Z(n1849) );
  AND U3329 ( .A(n307), .B(n3673), .Z(n3672) );
  XOR U3330 ( .A(n3674), .B(n3671), .Z(n3673) );
  XOR U3331 ( .A(n3675), .B(n3676), .Z(n3663) );
  AND U3332 ( .A(n3677), .B(n3678), .Z(n3676) );
  XOR U3333 ( .A(n3675), .B(n1864), .Z(n3678) );
  XOR U3334 ( .A(n3679), .B(n3680), .Z(n1864) );
  AND U3335 ( .A(n310), .B(n3681), .Z(n3680) );
  XOR U3336 ( .A(n3682), .B(n3679), .Z(n3681) );
  XNOR U3337 ( .A(n1861), .B(n3675), .Z(n3677) );
  XOR U3338 ( .A(n3683), .B(n3684), .Z(n1861) );
  AND U3339 ( .A(n307), .B(n3685), .Z(n3684) );
  XOR U3340 ( .A(n3686), .B(n3683), .Z(n3685) );
  XOR U3341 ( .A(n3687), .B(n3688), .Z(n3675) );
  AND U3342 ( .A(n3689), .B(n3690), .Z(n3688) );
  XOR U3343 ( .A(n3687), .B(n1876), .Z(n3690) );
  XOR U3344 ( .A(n3691), .B(n3692), .Z(n1876) );
  AND U3345 ( .A(n310), .B(n3693), .Z(n3692) );
  XOR U3346 ( .A(n3694), .B(n3691), .Z(n3693) );
  XNOR U3347 ( .A(n1873), .B(n3687), .Z(n3689) );
  XOR U3348 ( .A(n3695), .B(n3696), .Z(n1873) );
  AND U3349 ( .A(n307), .B(n3697), .Z(n3696) );
  XOR U3350 ( .A(n3698), .B(n3695), .Z(n3697) );
  XOR U3351 ( .A(n3699), .B(n3700), .Z(n3687) );
  AND U3352 ( .A(n3701), .B(n3702), .Z(n3700) );
  XOR U3353 ( .A(n3699), .B(n1888), .Z(n3702) );
  XOR U3354 ( .A(n3703), .B(n3704), .Z(n1888) );
  AND U3355 ( .A(n310), .B(n3705), .Z(n3704) );
  XOR U3356 ( .A(n3706), .B(n3703), .Z(n3705) );
  XNOR U3357 ( .A(n1885), .B(n3699), .Z(n3701) );
  XOR U3358 ( .A(n3707), .B(n3708), .Z(n1885) );
  AND U3359 ( .A(n307), .B(n3709), .Z(n3708) );
  XOR U3360 ( .A(n3710), .B(n3707), .Z(n3709) );
  XOR U3361 ( .A(n3711), .B(n3712), .Z(n3699) );
  AND U3362 ( .A(n3713), .B(n3714), .Z(n3712) );
  XOR U3363 ( .A(n3711), .B(n1900), .Z(n3714) );
  XOR U3364 ( .A(n3715), .B(n3716), .Z(n1900) );
  AND U3365 ( .A(n310), .B(n3717), .Z(n3716) );
  XOR U3366 ( .A(n3718), .B(n3715), .Z(n3717) );
  XNOR U3367 ( .A(n1897), .B(n3711), .Z(n3713) );
  XOR U3368 ( .A(n3719), .B(n3720), .Z(n1897) );
  AND U3369 ( .A(n307), .B(n3721), .Z(n3720) );
  XOR U3370 ( .A(n3722), .B(n3719), .Z(n3721) );
  XOR U3371 ( .A(n3723), .B(n3724), .Z(n3711) );
  AND U3372 ( .A(n3725), .B(n3726), .Z(n3724) );
  XOR U3373 ( .A(n3723), .B(n1912), .Z(n3726) );
  XOR U3374 ( .A(n3727), .B(n3728), .Z(n1912) );
  AND U3375 ( .A(n310), .B(n3729), .Z(n3728) );
  XOR U3376 ( .A(n3730), .B(n3727), .Z(n3729) );
  XNOR U3377 ( .A(n1909), .B(n3723), .Z(n3725) );
  XOR U3378 ( .A(n3731), .B(n3732), .Z(n1909) );
  AND U3379 ( .A(n307), .B(n3733), .Z(n3732) );
  XOR U3380 ( .A(n3734), .B(n3731), .Z(n3733) );
  XOR U3381 ( .A(n3735), .B(n3736), .Z(n3723) );
  AND U3382 ( .A(n3737), .B(n3738), .Z(n3736) );
  XOR U3383 ( .A(n3735), .B(n1924), .Z(n3738) );
  XOR U3384 ( .A(n3739), .B(n3740), .Z(n1924) );
  AND U3385 ( .A(n310), .B(n3741), .Z(n3740) );
  XOR U3386 ( .A(n3742), .B(n3739), .Z(n3741) );
  XNOR U3387 ( .A(n1921), .B(n3735), .Z(n3737) );
  XOR U3388 ( .A(n3743), .B(n3744), .Z(n1921) );
  AND U3389 ( .A(n307), .B(n3745), .Z(n3744) );
  XOR U3390 ( .A(n3746), .B(n3743), .Z(n3745) );
  XOR U3391 ( .A(n3747), .B(n3748), .Z(n3735) );
  AND U3392 ( .A(n3749), .B(n3750), .Z(n3748) );
  XOR U3393 ( .A(n3747), .B(n1936), .Z(n3750) );
  XOR U3394 ( .A(n3751), .B(n3752), .Z(n1936) );
  AND U3395 ( .A(n310), .B(n3753), .Z(n3752) );
  XOR U3396 ( .A(n3754), .B(n3751), .Z(n3753) );
  XNOR U3397 ( .A(n1933), .B(n3747), .Z(n3749) );
  XOR U3398 ( .A(n3755), .B(n3756), .Z(n1933) );
  AND U3399 ( .A(n307), .B(n3757), .Z(n3756) );
  XOR U3400 ( .A(n3758), .B(n3755), .Z(n3757) );
  XOR U3401 ( .A(n3759), .B(n3760), .Z(n3747) );
  AND U3402 ( .A(n3761), .B(n3762), .Z(n3760) );
  XOR U3403 ( .A(n3759), .B(n1948), .Z(n3762) );
  XOR U3404 ( .A(n3763), .B(n3764), .Z(n1948) );
  AND U3405 ( .A(n310), .B(n3765), .Z(n3764) );
  XOR U3406 ( .A(n3766), .B(n3763), .Z(n3765) );
  XNOR U3407 ( .A(n1945), .B(n3759), .Z(n3761) );
  XOR U3408 ( .A(n3767), .B(n3768), .Z(n1945) );
  AND U3409 ( .A(n307), .B(n3769), .Z(n3768) );
  XOR U3410 ( .A(n3770), .B(n3767), .Z(n3769) );
  XOR U3411 ( .A(n3771), .B(n3772), .Z(n3759) );
  AND U3412 ( .A(n3773), .B(n3774), .Z(n3772) );
  XOR U3413 ( .A(n3771), .B(n1960), .Z(n3774) );
  XOR U3414 ( .A(n3775), .B(n3776), .Z(n1960) );
  AND U3415 ( .A(n310), .B(n3777), .Z(n3776) );
  XOR U3416 ( .A(n3778), .B(n3775), .Z(n3777) );
  XNOR U3417 ( .A(n1957), .B(n3771), .Z(n3773) );
  XOR U3418 ( .A(n3779), .B(n3780), .Z(n1957) );
  AND U3419 ( .A(n307), .B(n3781), .Z(n3780) );
  XOR U3420 ( .A(n3782), .B(n3779), .Z(n3781) );
  XOR U3421 ( .A(n3783), .B(n3784), .Z(n3771) );
  AND U3422 ( .A(n3785), .B(n3786), .Z(n3784) );
  XOR U3423 ( .A(n3783), .B(n1972), .Z(n3786) );
  XOR U3424 ( .A(n3787), .B(n3788), .Z(n1972) );
  AND U3425 ( .A(n310), .B(n3789), .Z(n3788) );
  XOR U3426 ( .A(n3790), .B(n3787), .Z(n3789) );
  XNOR U3427 ( .A(n1969), .B(n3783), .Z(n3785) );
  XOR U3428 ( .A(n3791), .B(n3792), .Z(n1969) );
  AND U3429 ( .A(n307), .B(n3793), .Z(n3792) );
  XOR U3430 ( .A(n3794), .B(n3791), .Z(n3793) );
  XOR U3431 ( .A(n3795), .B(n3796), .Z(n3783) );
  AND U3432 ( .A(n3797), .B(n3798), .Z(n3796) );
  XOR U3433 ( .A(n3795), .B(n1984), .Z(n3798) );
  XOR U3434 ( .A(n3799), .B(n3800), .Z(n1984) );
  AND U3435 ( .A(n310), .B(n3801), .Z(n3800) );
  XOR U3436 ( .A(n3802), .B(n3799), .Z(n3801) );
  XNOR U3437 ( .A(n1981), .B(n3795), .Z(n3797) );
  XOR U3438 ( .A(n3803), .B(n3804), .Z(n1981) );
  AND U3439 ( .A(n307), .B(n3805), .Z(n3804) );
  XOR U3440 ( .A(n3806), .B(n3803), .Z(n3805) );
  XOR U3441 ( .A(n3807), .B(n3808), .Z(n3795) );
  AND U3442 ( .A(n3809), .B(n3810), .Z(n3808) );
  XOR U3443 ( .A(n3807), .B(n1996), .Z(n3810) );
  XOR U3444 ( .A(n3811), .B(n3812), .Z(n1996) );
  AND U3445 ( .A(n310), .B(n3813), .Z(n3812) );
  XOR U3446 ( .A(n3814), .B(n3811), .Z(n3813) );
  XNOR U3447 ( .A(n1993), .B(n3807), .Z(n3809) );
  XOR U3448 ( .A(n3815), .B(n3816), .Z(n1993) );
  AND U3449 ( .A(n307), .B(n3817), .Z(n3816) );
  XOR U3450 ( .A(n3818), .B(n3815), .Z(n3817) );
  XOR U3451 ( .A(n3819), .B(n3820), .Z(n3807) );
  AND U3452 ( .A(n3821), .B(n3822), .Z(n3820) );
  XOR U3453 ( .A(n3819), .B(n2008), .Z(n3822) );
  XOR U3454 ( .A(n3823), .B(n3824), .Z(n2008) );
  AND U3455 ( .A(n310), .B(n3825), .Z(n3824) );
  XOR U3456 ( .A(n3826), .B(n3823), .Z(n3825) );
  XNOR U3457 ( .A(n2005), .B(n3819), .Z(n3821) );
  XOR U3458 ( .A(n3827), .B(n3828), .Z(n2005) );
  AND U3459 ( .A(n307), .B(n3829), .Z(n3828) );
  XOR U3460 ( .A(n3830), .B(n3827), .Z(n3829) );
  XOR U3461 ( .A(n3831), .B(n3832), .Z(n3819) );
  AND U3462 ( .A(n3833), .B(n3834), .Z(n3832) );
  XOR U3463 ( .A(n3831), .B(n2020), .Z(n3834) );
  XOR U3464 ( .A(n3835), .B(n3836), .Z(n2020) );
  AND U3465 ( .A(n310), .B(n3837), .Z(n3836) );
  XOR U3466 ( .A(n3838), .B(n3835), .Z(n3837) );
  XNOR U3467 ( .A(n2017), .B(n3831), .Z(n3833) );
  XOR U3468 ( .A(n3839), .B(n3840), .Z(n2017) );
  AND U3469 ( .A(n307), .B(n3841), .Z(n3840) );
  XOR U3470 ( .A(n3842), .B(n3839), .Z(n3841) );
  XOR U3471 ( .A(n3843), .B(n3844), .Z(n3831) );
  AND U3472 ( .A(n3845), .B(n3846), .Z(n3844) );
  XOR U3473 ( .A(n3843), .B(n2032), .Z(n3846) );
  XOR U3474 ( .A(n3847), .B(n3848), .Z(n2032) );
  AND U3475 ( .A(n310), .B(n3849), .Z(n3848) );
  XOR U3476 ( .A(n3850), .B(n3847), .Z(n3849) );
  XNOR U3477 ( .A(n2029), .B(n3843), .Z(n3845) );
  XOR U3478 ( .A(n3851), .B(n3852), .Z(n2029) );
  AND U3479 ( .A(n307), .B(n3853), .Z(n3852) );
  XOR U3480 ( .A(n3854), .B(n3851), .Z(n3853) );
  XOR U3481 ( .A(n3855), .B(n3856), .Z(n3843) );
  AND U3482 ( .A(n3857), .B(n3858), .Z(n3856) );
  XOR U3483 ( .A(n3855), .B(n2044), .Z(n3858) );
  XOR U3484 ( .A(n3859), .B(n3860), .Z(n2044) );
  AND U3485 ( .A(n310), .B(n3861), .Z(n3860) );
  XOR U3486 ( .A(n3862), .B(n3859), .Z(n3861) );
  XNOR U3487 ( .A(n2041), .B(n3855), .Z(n3857) );
  XOR U3488 ( .A(n3863), .B(n3864), .Z(n2041) );
  AND U3489 ( .A(n307), .B(n3865), .Z(n3864) );
  XOR U3490 ( .A(n3866), .B(n3863), .Z(n3865) );
  XOR U3491 ( .A(n3867), .B(n3868), .Z(n3855) );
  AND U3492 ( .A(n3869), .B(n3870), .Z(n3868) );
  XOR U3493 ( .A(n3867), .B(n2056), .Z(n3870) );
  XOR U3494 ( .A(n3871), .B(n3872), .Z(n2056) );
  AND U3495 ( .A(n310), .B(n3873), .Z(n3872) );
  XOR U3496 ( .A(n3874), .B(n3871), .Z(n3873) );
  XNOR U3497 ( .A(n2053), .B(n3867), .Z(n3869) );
  XOR U3498 ( .A(n3875), .B(n3876), .Z(n2053) );
  AND U3499 ( .A(n307), .B(n3877), .Z(n3876) );
  XOR U3500 ( .A(n3878), .B(n3875), .Z(n3877) );
  XOR U3501 ( .A(n3879), .B(n3880), .Z(n3867) );
  AND U3502 ( .A(n3881), .B(n3882), .Z(n3880) );
  XOR U3503 ( .A(n3879), .B(n2068), .Z(n3882) );
  XOR U3504 ( .A(n3883), .B(n3884), .Z(n2068) );
  AND U3505 ( .A(n310), .B(n3885), .Z(n3884) );
  XOR U3506 ( .A(n3886), .B(n3883), .Z(n3885) );
  XNOR U3507 ( .A(n2065), .B(n3879), .Z(n3881) );
  XOR U3508 ( .A(n3887), .B(n3888), .Z(n2065) );
  AND U3509 ( .A(n307), .B(n3889), .Z(n3888) );
  XOR U3510 ( .A(n3890), .B(n3887), .Z(n3889) );
  XOR U3511 ( .A(n3891), .B(n3892), .Z(n3879) );
  AND U3512 ( .A(n3893), .B(n3894), .Z(n3892) );
  XOR U3513 ( .A(n3891), .B(n2080), .Z(n3894) );
  XOR U3514 ( .A(n3895), .B(n3896), .Z(n2080) );
  AND U3515 ( .A(n310), .B(n3897), .Z(n3896) );
  XOR U3516 ( .A(n3898), .B(n3895), .Z(n3897) );
  XNOR U3517 ( .A(n2077), .B(n3891), .Z(n3893) );
  XOR U3518 ( .A(n3899), .B(n3900), .Z(n2077) );
  AND U3519 ( .A(n307), .B(n3901), .Z(n3900) );
  XOR U3520 ( .A(n3902), .B(n3899), .Z(n3901) );
  XOR U3521 ( .A(n3903), .B(n3904), .Z(n3891) );
  AND U3522 ( .A(n3905), .B(n3906), .Z(n3904) );
  XOR U3523 ( .A(n3903), .B(n2092), .Z(n3906) );
  XOR U3524 ( .A(n3907), .B(n3908), .Z(n2092) );
  AND U3525 ( .A(n310), .B(n3909), .Z(n3908) );
  XOR U3526 ( .A(n3910), .B(n3907), .Z(n3909) );
  XNOR U3527 ( .A(n2089), .B(n3903), .Z(n3905) );
  XOR U3528 ( .A(n3911), .B(n3912), .Z(n2089) );
  AND U3529 ( .A(n307), .B(n3913), .Z(n3912) );
  XOR U3530 ( .A(n3914), .B(n3911), .Z(n3913) );
  XOR U3531 ( .A(n3915), .B(n3916), .Z(n3903) );
  AND U3532 ( .A(n3917), .B(n3918), .Z(n3916) );
  XOR U3533 ( .A(n3915), .B(n2104), .Z(n3918) );
  XOR U3534 ( .A(n3919), .B(n3920), .Z(n2104) );
  AND U3535 ( .A(n310), .B(n3921), .Z(n3920) );
  XOR U3536 ( .A(n3922), .B(n3919), .Z(n3921) );
  XNOR U3537 ( .A(n2101), .B(n3915), .Z(n3917) );
  XOR U3538 ( .A(n3923), .B(n3924), .Z(n2101) );
  AND U3539 ( .A(n307), .B(n3925), .Z(n3924) );
  XOR U3540 ( .A(n3926), .B(n3923), .Z(n3925) );
  XOR U3541 ( .A(n3927), .B(n3928), .Z(n3915) );
  AND U3542 ( .A(n3929), .B(n3930), .Z(n3928) );
  XOR U3543 ( .A(n3927), .B(n2116), .Z(n3930) );
  XOR U3544 ( .A(n3931), .B(n3932), .Z(n2116) );
  AND U3545 ( .A(n310), .B(n3933), .Z(n3932) );
  XOR U3546 ( .A(n3934), .B(n3931), .Z(n3933) );
  XNOR U3547 ( .A(n2113), .B(n3927), .Z(n3929) );
  XOR U3548 ( .A(n3935), .B(n3936), .Z(n2113) );
  AND U3549 ( .A(n307), .B(n3937), .Z(n3936) );
  XOR U3550 ( .A(n3938), .B(n3935), .Z(n3937) );
  XOR U3551 ( .A(n3939), .B(n3940), .Z(n3927) );
  AND U3552 ( .A(n3941), .B(n3942), .Z(n3940) );
  XOR U3553 ( .A(n2128), .B(n3939), .Z(n3942) );
  XOR U3554 ( .A(n3943), .B(n3944), .Z(n2128) );
  AND U3555 ( .A(n310), .B(n3945), .Z(n3944) );
  XOR U3556 ( .A(n3943), .B(n3946), .Z(n3945) );
  XNOR U3557 ( .A(n3939), .B(n2125), .Z(n3941) );
  XOR U3558 ( .A(n3947), .B(n3948), .Z(n2125) );
  AND U3559 ( .A(n307), .B(n3949), .Z(n3948) );
  XOR U3560 ( .A(n3947), .B(n3950), .Z(n3949) );
  XOR U3561 ( .A(n3951), .B(n3952), .Z(n3939) );
  AND U3562 ( .A(n3953), .B(n3954), .Z(n3952) );
  XNOR U3563 ( .A(n3955), .B(n2141), .Z(n3954) );
  XOR U3564 ( .A(n3956), .B(n3957), .Z(n2141) );
  AND U3565 ( .A(n310), .B(n3958), .Z(n3957) );
  XOR U3566 ( .A(n3959), .B(n3956), .Z(n3958) );
  XNOR U3567 ( .A(n2138), .B(n3951), .Z(n3953) );
  XOR U3568 ( .A(n3960), .B(n3961), .Z(n2138) );
  AND U3569 ( .A(n307), .B(n3962), .Z(n3961) );
  XOR U3570 ( .A(n3963), .B(n3960), .Z(n3962) );
  IV U3571 ( .A(n3955), .Z(n3951) );
  AND U3572 ( .A(n3587), .B(n3590), .Z(n3955) );
  XNOR U3573 ( .A(n3964), .B(n3965), .Z(n3590) );
  AND U3574 ( .A(n310), .B(n3966), .Z(n3965) );
  XNOR U3575 ( .A(n3967), .B(n3964), .Z(n3966) );
  XOR U3576 ( .A(n3968), .B(n3969), .Z(n310) );
  AND U3577 ( .A(n3970), .B(n3971), .Z(n3969) );
  XOR U3578 ( .A(n3598), .B(n3968), .Z(n3971) );
  IV U3579 ( .A(n3972), .Z(n3598) );
  AND U3580 ( .A(p_input[3839]), .B(p_input[3807]), .Z(n3972) );
  XOR U3581 ( .A(n3968), .B(n3595), .Z(n3970) );
  AND U3582 ( .A(p_input[3743]), .B(p_input[3775]), .Z(n3595) );
  XOR U3583 ( .A(n3973), .B(n3974), .Z(n3968) );
  AND U3584 ( .A(n3975), .B(n3976), .Z(n3974) );
  XOR U3585 ( .A(n3973), .B(n3610), .Z(n3976) );
  XNOR U3586 ( .A(p_input[3806]), .B(n3977), .Z(n3610) );
  AND U3587 ( .A(n194), .B(n3978), .Z(n3977) );
  XOR U3588 ( .A(p_input[3838]), .B(p_input[3806]), .Z(n3978) );
  XNOR U3589 ( .A(n3607), .B(n3973), .Z(n3975) );
  XOR U3590 ( .A(n3979), .B(n3980), .Z(n3607) );
  AND U3591 ( .A(n192), .B(n3981), .Z(n3980) );
  XOR U3592 ( .A(p_input[3774]), .B(p_input[3742]), .Z(n3981) );
  XOR U3593 ( .A(n3982), .B(n3983), .Z(n3973) );
  AND U3594 ( .A(n3984), .B(n3985), .Z(n3983) );
  XOR U3595 ( .A(n3982), .B(n3622), .Z(n3985) );
  XNOR U3596 ( .A(p_input[3805]), .B(n3986), .Z(n3622) );
  AND U3597 ( .A(n194), .B(n3987), .Z(n3986) );
  XOR U3598 ( .A(p_input[3837]), .B(p_input[3805]), .Z(n3987) );
  XNOR U3599 ( .A(n3619), .B(n3982), .Z(n3984) );
  XOR U3600 ( .A(n3988), .B(n3989), .Z(n3619) );
  AND U3601 ( .A(n192), .B(n3990), .Z(n3989) );
  XOR U3602 ( .A(p_input[3773]), .B(p_input[3741]), .Z(n3990) );
  XOR U3603 ( .A(n3991), .B(n3992), .Z(n3982) );
  AND U3604 ( .A(n3993), .B(n3994), .Z(n3992) );
  XOR U3605 ( .A(n3991), .B(n3634), .Z(n3994) );
  XNOR U3606 ( .A(p_input[3804]), .B(n3995), .Z(n3634) );
  AND U3607 ( .A(n194), .B(n3996), .Z(n3995) );
  XOR U3608 ( .A(p_input[3836]), .B(p_input[3804]), .Z(n3996) );
  XNOR U3609 ( .A(n3631), .B(n3991), .Z(n3993) );
  XOR U3610 ( .A(n3997), .B(n3998), .Z(n3631) );
  AND U3611 ( .A(n192), .B(n3999), .Z(n3998) );
  XOR U3612 ( .A(p_input[3772]), .B(p_input[3740]), .Z(n3999) );
  XOR U3613 ( .A(n4000), .B(n4001), .Z(n3991) );
  AND U3614 ( .A(n4002), .B(n4003), .Z(n4001) );
  XOR U3615 ( .A(n4000), .B(n3646), .Z(n4003) );
  XNOR U3616 ( .A(p_input[3803]), .B(n4004), .Z(n3646) );
  AND U3617 ( .A(n194), .B(n4005), .Z(n4004) );
  XOR U3618 ( .A(p_input[3835]), .B(p_input[3803]), .Z(n4005) );
  XNOR U3619 ( .A(n3643), .B(n4000), .Z(n4002) );
  XOR U3620 ( .A(n4006), .B(n4007), .Z(n3643) );
  AND U3621 ( .A(n192), .B(n4008), .Z(n4007) );
  XOR U3622 ( .A(p_input[3771]), .B(p_input[3739]), .Z(n4008) );
  XOR U3623 ( .A(n4009), .B(n4010), .Z(n4000) );
  AND U3624 ( .A(n4011), .B(n4012), .Z(n4010) );
  XOR U3625 ( .A(n4009), .B(n3658), .Z(n4012) );
  XNOR U3626 ( .A(p_input[3802]), .B(n4013), .Z(n3658) );
  AND U3627 ( .A(n194), .B(n4014), .Z(n4013) );
  XOR U3628 ( .A(p_input[3834]), .B(p_input[3802]), .Z(n4014) );
  XNOR U3629 ( .A(n3655), .B(n4009), .Z(n4011) );
  XOR U3630 ( .A(n4015), .B(n4016), .Z(n3655) );
  AND U3631 ( .A(n192), .B(n4017), .Z(n4016) );
  XOR U3632 ( .A(p_input[3770]), .B(p_input[3738]), .Z(n4017) );
  XOR U3633 ( .A(n4018), .B(n4019), .Z(n4009) );
  AND U3634 ( .A(n4020), .B(n4021), .Z(n4019) );
  XOR U3635 ( .A(n4018), .B(n3670), .Z(n4021) );
  XNOR U3636 ( .A(p_input[3801]), .B(n4022), .Z(n3670) );
  AND U3637 ( .A(n194), .B(n4023), .Z(n4022) );
  XOR U3638 ( .A(p_input[3833]), .B(p_input[3801]), .Z(n4023) );
  XNOR U3639 ( .A(n3667), .B(n4018), .Z(n4020) );
  XOR U3640 ( .A(n4024), .B(n4025), .Z(n3667) );
  AND U3641 ( .A(n192), .B(n4026), .Z(n4025) );
  XOR U3642 ( .A(p_input[3769]), .B(p_input[3737]), .Z(n4026) );
  XOR U3643 ( .A(n4027), .B(n4028), .Z(n4018) );
  AND U3644 ( .A(n4029), .B(n4030), .Z(n4028) );
  XOR U3645 ( .A(n4027), .B(n3682), .Z(n4030) );
  XNOR U3646 ( .A(p_input[3800]), .B(n4031), .Z(n3682) );
  AND U3647 ( .A(n194), .B(n4032), .Z(n4031) );
  XOR U3648 ( .A(p_input[3832]), .B(p_input[3800]), .Z(n4032) );
  XNOR U3649 ( .A(n3679), .B(n4027), .Z(n4029) );
  XOR U3650 ( .A(n4033), .B(n4034), .Z(n3679) );
  AND U3651 ( .A(n192), .B(n4035), .Z(n4034) );
  XOR U3652 ( .A(p_input[3768]), .B(p_input[3736]), .Z(n4035) );
  XOR U3653 ( .A(n4036), .B(n4037), .Z(n4027) );
  AND U3654 ( .A(n4038), .B(n4039), .Z(n4037) );
  XOR U3655 ( .A(n4036), .B(n3694), .Z(n4039) );
  XNOR U3656 ( .A(p_input[3799]), .B(n4040), .Z(n3694) );
  AND U3657 ( .A(n194), .B(n4041), .Z(n4040) );
  XOR U3658 ( .A(p_input[3831]), .B(p_input[3799]), .Z(n4041) );
  XNOR U3659 ( .A(n3691), .B(n4036), .Z(n4038) );
  XOR U3660 ( .A(n4042), .B(n4043), .Z(n3691) );
  AND U3661 ( .A(n192), .B(n4044), .Z(n4043) );
  XOR U3662 ( .A(p_input[3767]), .B(p_input[3735]), .Z(n4044) );
  XOR U3663 ( .A(n4045), .B(n4046), .Z(n4036) );
  AND U3664 ( .A(n4047), .B(n4048), .Z(n4046) );
  XOR U3665 ( .A(n4045), .B(n3706), .Z(n4048) );
  XNOR U3666 ( .A(p_input[3798]), .B(n4049), .Z(n3706) );
  AND U3667 ( .A(n194), .B(n4050), .Z(n4049) );
  XOR U3668 ( .A(p_input[3830]), .B(p_input[3798]), .Z(n4050) );
  XNOR U3669 ( .A(n3703), .B(n4045), .Z(n4047) );
  XOR U3670 ( .A(n4051), .B(n4052), .Z(n3703) );
  AND U3671 ( .A(n192), .B(n4053), .Z(n4052) );
  XOR U3672 ( .A(p_input[3766]), .B(p_input[3734]), .Z(n4053) );
  XOR U3673 ( .A(n4054), .B(n4055), .Z(n4045) );
  AND U3674 ( .A(n4056), .B(n4057), .Z(n4055) );
  XOR U3675 ( .A(n4054), .B(n3718), .Z(n4057) );
  XNOR U3676 ( .A(p_input[3797]), .B(n4058), .Z(n3718) );
  AND U3677 ( .A(n194), .B(n4059), .Z(n4058) );
  XOR U3678 ( .A(p_input[3829]), .B(p_input[3797]), .Z(n4059) );
  XNOR U3679 ( .A(n3715), .B(n4054), .Z(n4056) );
  XOR U3680 ( .A(n4060), .B(n4061), .Z(n3715) );
  AND U3681 ( .A(n192), .B(n4062), .Z(n4061) );
  XOR U3682 ( .A(p_input[3765]), .B(p_input[3733]), .Z(n4062) );
  XOR U3683 ( .A(n4063), .B(n4064), .Z(n4054) );
  AND U3684 ( .A(n4065), .B(n4066), .Z(n4064) );
  XOR U3685 ( .A(n4063), .B(n3730), .Z(n4066) );
  XNOR U3686 ( .A(p_input[3796]), .B(n4067), .Z(n3730) );
  AND U3687 ( .A(n194), .B(n4068), .Z(n4067) );
  XOR U3688 ( .A(p_input[3828]), .B(p_input[3796]), .Z(n4068) );
  XNOR U3689 ( .A(n3727), .B(n4063), .Z(n4065) );
  XOR U3690 ( .A(n4069), .B(n4070), .Z(n3727) );
  AND U3691 ( .A(n192), .B(n4071), .Z(n4070) );
  XOR U3692 ( .A(p_input[3764]), .B(p_input[3732]), .Z(n4071) );
  XOR U3693 ( .A(n4072), .B(n4073), .Z(n4063) );
  AND U3694 ( .A(n4074), .B(n4075), .Z(n4073) );
  XOR U3695 ( .A(n4072), .B(n3742), .Z(n4075) );
  XNOR U3696 ( .A(p_input[3795]), .B(n4076), .Z(n3742) );
  AND U3697 ( .A(n194), .B(n4077), .Z(n4076) );
  XOR U3698 ( .A(p_input[3827]), .B(p_input[3795]), .Z(n4077) );
  XNOR U3699 ( .A(n3739), .B(n4072), .Z(n4074) );
  XOR U3700 ( .A(n4078), .B(n4079), .Z(n3739) );
  AND U3701 ( .A(n192), .B(n4080), .Z(n4079) );
  XOR U3702 ( .A(p_input[3763]), .B(p_input[3731]), .Z(n4080) );
  XOR U3703 ( .A(n4081), .B(n4082), .Z(n4072) );
  AND U3704 ( .A(n4083), .B(n4084), .Z(n4082) );
  XOR U3705 ( .A(n4081), .B(n3754), .Z(n4084) );
  XNOR U3706 ( .A(p_input[3794]), .B(n4085), .Z(n3754) );
  AND U3707 ( .A(n194), .B(n4086), .Z(n4085) );
  XOR U3708 ( .A(p_input[3826]), .B(p_input[3794]), .Z(n4086) );
  XNOR U3709 ( .A(n3751), .B(n4081), .Z(n4083) );
  XOR U3710 ( .A(n4087), .B(n4088), .Z(n3751) );
  AND U3711 ( .A(n192), .B(n4089), .Z(n4088) );
  XOR U3712 ( .A(p_input[3762]), .B(p_input[3730]), .Z(n4089) );
  XOR U3713 ( .A(n4090), .B(n4091), .Z(n4081) );
  AND U3714 ( .A(n4092), .B(n4093), .Z(n4091) );
  XOR U3715 ( .A(n4090), .B(n3766), .Z(n4093) );
  XNOR U3716 ( .A(p_input[3793]), .B(n4094), .Z(n3766) );
  AND U3717 ( .A(n194), .B(n4095), .Z(n4094) );
  XOR U3718 ( .A(p_input[3825]), .B(p_input[3793]), .Z(n4095) );
  XNOR U3719 ( .A(n3763), .B(n4090), .Z(n4092) );
  XOR U3720 ( .A(n4096), .B(n4097), .Z(n3763) );
  AND U3721 ( .A(n192), .B(n4098), .Z(n4097) );
  XOR U3722 ( .A(p_input[3761]), .B(p_input[3729]), .Z(n4098) );
  XOR U3723 ( .A(n4099), .B(n4100), .Z(n4090) );
  AND U3724 ( .A(n4101), .B(n4102), .Z(n4100) );
  XOR U3725 ( .A(n4099), .B(n3778), .Z(n4102) );
  XNOR U3726 ( .A(p_input[3792]), .B(n4103), .Z(n3778) );
  AND U3727 ( .A(n194), .B(n4104), .Z(n4103) );
  XOR U3728 ( .A(p_input[3824]), .B(p_input[3792]), .Z(n4104) );
  XNOR U3729 ( .A(n3775), .B(n4099), .Z(n4101) );
  XOR U3730 ( .A(n4105), .B(n4106), .Z(n3775) );
  AND U3731 ( .A(n192), .B(n4107), .Z(n4106) );
  XOR U3732 ( .A(p_input[3760]), .B(p_input[3728]), .Z(n4107) );
  XOR U3733 ( .A(n4108), .B(n4109), .Z(n4099) );
  AND U3734 ( .A(n4110), .B(n4111), .Z(n4109) );
  XOR U3735 ( .A(n4108), .B(n3790), .Z(n4111) );
  XNOR U3736 ( .A(p_input[3791]), .B(n4112), .Z(n3790) );
  AND U3737 ( .A(n194), .B(n4113), .Z(n4112) );
  XOR U3738 ( .A(p_input[3823]), .B(p_input[3791]), .Z(n4113) );
  XNOR U3739 ( .A(n3787), .B(n4108), .Z(n4110) );
  XOR U3740 ( .A(n4114), .B(n4115), .Z(n3787) );
  AND U3741 ( .A(n192), .B(n4116), .Z(n4115) );
  XOR U3742 ( .A(p_input[3759]), .B(p_input[3727]), .Z(n4116) );
  XOR U3743 ( .A(n4117), .B(n4118), .Z(n4108) );
  AND U3744 ( .A(n4119), .B(n4120), .Z(n4118) );
  XOR U3745 ( .A(n4117), .B(n3802), .Z(n4120) );
  XNOR U3746 ( .A(p_input[3790]), .B(n4121), .Z(n3802) );
  AND U3747 ( .A(n194), .B(n4122), .Z(n4121) );
  XOR U3748 ( .A(p_input[3822]), .B(p_input[3790]), .Z(n4122) );
  XNOR U3749 ( .A(n3799), .B(n4117), .Z(n4119) );
  XOR U3750 ( .A(n4123), .B(n4124), .Z(n3799) );
  AND U3751 ( .A(n192), .B(n4125), .Z(n4124) );
  XOR U3752 ( .A(p_input[3758]), .B(p_input[3726]), .Z(n4125) );
  XOR U3753 ( .A(n4126), .B(n4127), .Z(n4117) );
  AND U3754 ( .A(n4128), .B(n4129), .Z(n4127) );
  XOR U3755 ( .A(n4126), .B(n3814), .Z(n4129) );
  XNOR U3756 ( .A(p_input[3789]), .B(n4130), .Z(n3814) );
  AND U3757 ( .A(n194), .B(n4131), .Z(n4130) );
  XOR U3758 ( .A(p_input[3821]), .B(p_input[3789]), .Z(n4131) );
  XNOR U3759 ( .A(n3811), .B(n4126), .Z(n4128) );
  XOR U3760 ( .A(n4132), .B(n4133), .Z(n3811) );
  AND U3761 ( .A(n192), .B(n4134), .Z(n4133) );
  XOR U3762 ( .A(p_input[3757]), .B(p_input[3725]), .Z(n4134) );
  XOR U3763 ( .A(n4135), .B(n4136), .Z(n4126) );
  AND U3764 ( .A(n4137), .B(n4138), .Z(n4136) );
  XOR U3765 ( .A(n4135), .B(n3826), .Z(n4138) );
  XNOR U3766 ( .A(p_input[3788]), .B(n4139), .Z(n3826) );
  AND U3767 ( .A(n194), .B(n4140), .Z(n4139) );
  XOR U3768 ( .A(p_input[3820]), .B(p_input[3788]), .Z(n4140) );
  XNOR U3769 ( .A(n3823), .B(n4135), .Z(n4137) );
  XOR U3770 ( .A(n4141), .B(n4142), .Z(n3823) );
  AND U3771 ( .A(n192), .B(n4143), .Z(n4142) );
  XOR U3772 ( .A(p_input[3756]), .B(p_input[3724]), .Z(n4143) );
  XOR U3773 ( .A(n4144), .B(n4145), .Z(n4135) );
  AND U3774 ( .A(n4146), .B(n4147), .Z(n4145) );
  XOR U3775 ( .A(n4144), .B(n3838), .Z(n4147) );
  XNOR U3776 ( .A(p_input[3787]), .B(n4148), .Z(n3838) );
  AND U3777 ( .A(n194), .B(n4149), .Z(n4148) );
  XOR U3778 ( .A(p_input[3819]), .B(p_input[3787]), .Z(n4149) );
  XNOR U3779 ( .A(n3835), .B(n4144), .Z(n4146) );
  XOR U3780 ( .A(n4150), .B(n4151), .Z(n3835) );
  AND U3781 ( .A(n192), .B(n4152), .Z(n4151) );
  XOR U3782 ( .A(p_input[3755]), .B(p_input[3723]), .Z(n4152) );
  XOR U3783 ( .A(n4153), .B(n4154), .Z(n4144) );
  AND U3784 ( .A(n4155), .B(n4156), .Z(n4154) );
  XOR U3785 ( .A(n4153), .B(n3850), .Z(n4156) );
  XNOR U3786 ( .A(p_input[3786]), .B(n4157), .Z(n3850) );
  AND U3787 ( .A(n194), .B(n4158), .Z(n4157) );
  XOR U3788 ( .A(p_input[3818]), .B(p_input[3786]), .Z(n4158) );
  XNOR U3789 ( .A(n3847), .B(n4153), .Z(n4155) );
  XOR U3790 ( .A(n4159), .B(n4160), .Z(n3847) );
  AND U3791 ( .A(n192), .B(n4161), .Z(n4160) );
  XOR U3792 ( .A(p_input[3754]), .B(p_input[3722]), .Z(n4161) );
  XOR U3793 ( .A(n4162), .B(n4163), .Z(n4153) );
  AND U3794 ( .A(n4164), .B(n4165), .Z(n4163) );
  XOR U3795 ( .A(n4162), .B(n3862), .Z(n4165) );
  XNOR U3796 ( .A(p_input[3785]), .B(n4166), .Z(n3862) );
  AND U3797 ( .A(n194), .B(n4167), .Z(n4166) );
  XOR U3798 ( .A(p_input[3817]), .B(p_input[3785]), .Z(n4167) );
  XNOR U3799 ( .A(n3859), .B(n4162), .Z(n4164) );
  XOR U3800 ( .A(n4168), .B(n4169), .Z(n3859) );
  AND U3801 ( .A(n192), .B(n4170), .Z(n4169) );
  XOR U3802 ( .A(p_input[3753]), .B(p_input[3721]), .Z(n4170) );
  XOR U3803 ( .A(n4171), .B(n4172), .Z(n4162) );
  AND U3804 ( .A(n4173), .B(n4174), .Z(n4172) );
  XOR U3805 ( .A(n4171), .B(n3874), .Z(n4174) );
  XNOR U3806 ( .A(p_input[3784]), .B(n4175), .Z(n3874) );
  AND U3807 ( .A(n194), .B(n4176), .Z(n4175) );
  XOR U3808 ( .A(p_input[3816]), .B(p_input[3784]), .Z(n4176) );
  XNOR U3809 ( .A(n3871), .B(n4171), .Z(n4173) );
  XOR U3810 ( .A(n4177), .B(n4178), .Z(n3871) );
  AND U3811 ( .A(n192), .B(n4179), .Z(n4178) );
  XOR U3812 ( .A(p_input[3752]), .B(p_input[3720]), .Z(n4179) );
  XOR U3813 ( .A(n4180), .B(n4181), .Z(n4171) );
  AND U3814 ( .A(n4182), .B(n4183), .Z(n4181) );
  XOR U3815 ( .A(n4180), .B(n3886), .Z(n4183) );
  XNOR U3816 ( .A(p_input[3783]), .B(n4184), .Z(n3886) );
  AND U3817 ( .A(n194), .B(n4185), .Z(n4184) );
  XOR U3818 ( .A(p_input[3815]), .B(p_input[3783]), .Z(n4185) );
  XNOR U3819 ( .A(n3883), .B(n4180), .Z(n4182) );
  XOR U3820 ( .A(n4186), .B(n4187), .Z(n3883) );
  AND U3821 ( .A(n192), .B(n4188), .Z(n4187) );
  XOR U3822 ( .A(p_input[3751]), .B(p_input[3719]), .Z(n4188) );
  XOR U3823 ( .A(n4189), .B(n4190), .Z(n4180) );
  AND U3824 ( .A(n4191), .B(n4192), .Z(n4190) );
  XOR U3825 ( .A(n4189), .B(n3898), .Z(n4192) );
  XNOR U3826 ( .A(p_input[3782]), .B(n4193), .Z(n3898) );
  AND U3827 ( .A(n194), .B(n4194), .Z(n4193) );
  XOR U3828 ( .A(p_input[3814]), .B(p_input[3782]), .Z(n4194) );
  XNOR U3829 ( .A(n3895), .B(n4189), .Z(n4191) );
  XOR U3830 ( .A(n4195), .B(n4196), .Z(n3895) );
  AND U3831 ( .A(n192), .B(n4197), .Z(n4196) );
  XOR U3832 ( .A(p_input[3750]), .B(p_input[3718]), .Z(n4197) );
  XOR U3833 ( .A(n4198), .B(n4199), .Z(n4189) );
  AND U3834 ( .A(n4200), .B(n4201), .Z(n4199) );
  XOR U3835 ( .A(n4198), .B(n3910), .Z(n4201) );
  XNOR U3836 ( .A(p_input[3781]), .B(n4202), .Z(n3910) );
  AND U3837 ( .A(n194), .B(n4203), .Z(n4202) );
  XOR U3838 ( .A(p_input[3813]), .B(p_input[3781]), .Z(n4203) );
  XNOR U3839 ( .A(n3907), .B(n4198), .Z(n4200) );
  XOR U3840 ( .A(n4204), .B(n4205), .Z(n3907) );
  AND U3841 ( .A(n192), .B(n4206), .Z(n4205) );
  XOR U3842 ( .A(p_input[3749]), .B(p_input[3717]), .Z(n4206) );
  XOR U3843 ( .A(n4207), .B(n4208), .Z(n4198) );
  AND U3844 ( .A(n4209), .B(n4210), .Z(n4208) );
  XOR U3845 ( .A(n4207), .B(n3922), .Z(n4210) );
  XNOR U3846 ( .A(p_input[3780]), .B(n4211), .Z(n3922) );
  AND U3847 ( .A(n194), .B(n4212), .Z(n4211) );
  XOR U3848 ( .A(p_input[3812]), .B(p_input[3780]), .Z(n4212) );
  XNOR U3849 ( .A(n3919), .B(n4207), .Z(n4209) );
  XOR U3850 ( .A(n4213), .B(n4214), .Z(n3919) );
  AND U3851 ( .A(n192), .B(n4215), .Z(n4214) );
  XOR U3852 ( .A(p_input[3748]), .B(p_input[3716]), .Z(n4215) );
  XOR U3853 ( .A(n4216), .B(n4217), .Z(n4207) );
  AND U3854 ( .A(n4218), .B(n4219), .Z(n4217) );
  XOR U3855 ( .A(n4216), .B(n3934), .Z(n4219) );
  XNOR U3856 ( .A(p_input[3779]), .B(n4220), .Z(n3934) );
  AND U3857 ( .A(n194), .B(n4221), .Z(n4220) );
  XOR U3858 ( .A(p_input[3811]), .B(p_input[3779]), .Z(n4221) );
  XNOR U3859 ( .A(n3931), .B(n4216), .Z(n4218) );
  XOR U3860 ( .A(n4222), .B(n4223), .Z(n3931) );
  AND U3861 ( .A(n192), .B(n4224), .Z(n4223) );
  XOR U3862 ( .A(p_input[3747]), .B(p_input[3715]), .Z(n4224) );
  XOR U3863 ( .A(n4225), .B(n4226), .Z(n4216) );
  AND U3864 ( .A(n4227), .B(n4228), .Z(n4226) );
  XOR U3865 ( .A(n3946), .B(n4225), .Z(n4228) );
  XNOR U3866 ( .A(p_input[3778]), .B(n4229), .Z(n3946) );
  AND U3867 ( .A(n194), .B(n4230), .Z(n4229) );
  XOR U3868 ( .A(p_input[3810]), .B(p_input[3778]), .Z(n4230) );
  XNOR U3869 ( .A(n4225), .B(n3943), .Z(n4227) );
  XOR U3870 ( .A(n4231), .B(n4232), .Z(n3943) );
  AND U3871 ( .A(n192), .B(n4233), .Z(n4232) );
  XOR U3872 ( .A(p_input[3746]), .B(p_input[3714]), .Z(n4233) );
  XOR U3873 ( .A(n4234), .B(n4235), .Z(n4225) );
  AND U3874 ( .A(n4236), .B(n4237), .Z(n4235) );
  XNOR U3875 ( .A(n4238), .B(n3959), .Z(n4237) );
  XNOR U3876 ( .A(p_input[3777]), .B(n4239), .Z(n3959) );
  AND U3877 ( .A(n194), .B(n4240), .Z(n4239) );
  XNOR U3878 ( .A(p_input[3809]), .B(n4241), .Z(n4240) );
  IV U3879 ( .A(p_input[3777]), .Z(n4241) );
  XNOR U3880 ( .A(n3956), .B(n4234), .Z(n4236) );
  XNOR U3881 ( .A(p_input[3713]), .B(n4242), .Z(n3956) );
  AND U3882 ( .A(n192), .B(n4243), .Z(n4242) );
  XOR U3883 ( .A(p_input[3745]), .B(p_input[3713]), .Z(n4243) );
  IV U3884 ( .A(n4238), .Z(n4234) );
  AND U3885 ( .A(n3964), .B(n3967), .Z(n4238) );
  XOR U3886 ( .A(p_input[3776]), .B(n4244), .Z(n3967) );
  AND U3887 ( .A(n194), .B(n4245), .Z(n4244) );
  XOR U3888 ( .A(p_input[3808]), .B(p_input[3776]), .Z(n4245) );
  XOR U3889 ( .A(n4246), .B(n4247), .Z(n194) );
  AND U3890 ( .A(n4248), .B(n4249), .Z(n4247) );
  XNOR U3891 ( .A(p_input[3839]), .B(n4246), .Z(n4249) );
  XOR U3892 ( .A(n4246), .B(p_input[3807]), .Z(n4248) );
  XOR U3893 ( .A(n4250), .B(n4251), .Z(n4246) );
  AND U3894 ( .A(n4252), .B(n4253), .Z(n4251) );
  XNOR U3895 ( .A(p_input[3838]), .B(n4250), .Z(n4253) );
  XOR U3896 ( .A(n4250), .B(p_input[3806]), .Z(n4252) );
  XOR U3897 ( .A(n4254), .B(n4255), .Z(n4250) );
  AND U3898 ( .A(n4256), .B(n4257), .Z(n4255) );
  XNOR U3899 ( .A(p_input[3837]), .B(n4254), .Z(n4257) );
  XOR U3900 ( .A(n4254), .B(p_input[3805]), .Z(n4256) );
  XOR U3901 ( .A(n4258), .B(n4259), .Z(n4254) );
  AND U3902 ( .A(n4260), .B(n4261), .Z(n4259) );
  XNOR U3903 ( .A(p_input[3836]), .B(n4258), .Z(n4261) );
  XOR U3904 ( .A(n4258), .B(p_input[3804]), .Z(n4260) );
  XOR U3905 ( .A(n4262), .B(n4263), .Z(n4258) );
  AND U3906 ( .A(n4264), .B(n4265), .Z(n4263) );
  XNOR U3907 ( .A(p_input[3835]), .B(n4262), .Z(n4265) );
  XOR U3908 ( .A(n4262), .B(p_input[3803]), .Z(n4264) );
  XOR U3909 ( .A(n4266), .B(n4267), .Z(n4262) );
  AND U3910 ( .A(n4268), .B(n4269), .Z(n4267) );
  XNOR U3911 ( .A(p_input[3834]), .B(n4266), .Z(n4269) );
  XOR U3912 ( .A(n4266), .B(p_input[3802]), .Z(n4268) );
  XOR U3913 ( .A(n4270), .B(n4271), .Z(n4266) );
  AND U3914 ( .A(n4272), .B(n4273), .Z(n4271) );
  XNOR U3915 ( .A(p_input[3833]), .B(n4270), .Z(n4273) );
  XOR U3916 ( .A(n4270), .B(p_input[3801]), .Z(n4272) );
  XOR U3917 ( .A(n4274), .B(n4275), .Z(n4270) );
  AND U3918 ( .A(n4276), .B(n4277), .Z(n4275) );
  XNOR U3919 ( .A(p_input[3832]), .B(n4274), .Z(n4277) );
  XOR U3920 ( .A(n4274), .B(p_input[3800]), .Z(n4276) );
  XOR U3921 ( .A(n4278), .B(n4279), .Z(n4274) );
  AND U3922 ( .A(n4280), .B(n4281), .Z(n4279) );
  XNOR U3923 ( .A(p_input[3831]), .B(n4278), .Z(n4281) );
  XOR U3924 ( .A(n4278), .B(p_input[3799]), .Z(n4280) );
  XOR U3925 ( .A(n4282), .B(n4283), .Z(n4278) );
  AND U3926 ( .A(n4284), .B(n4285), .Z(n4283) );
  XNOR U3927 ( .A(p_input[3830]), .B(n4282), .Z(n4285) );
  XOR U3928 ( .A(n4282), .B(p_input[3798]), .Z(n4284) );
  XOR U3929 ( .A(n4286), .B(n4287), .Z(n4282) );
  AND U3930 ( .A(n4288), .B(n4289), .Z(n4287) );
  XNOR U3931 ( .A(p_input[3829]), .B(n4286), .Z(n4289) );
  XOR U3932 ( .A(n4286), .B(p_input[3797]), .Z(n4288) );
  XOR U3933 ( .A(n4290), .B(n4291), .Z(n4286) );
  AND U3934 ( .A(n4292), .B(n4293), .Z(n4291) );
  XNOR U3935 ( .A(p_input[3828]), .B(n4290), .Z(n4293) );
  XOR U3936 ( .A(n4290), .B(p_input[3796]), .Z(n4292) );
  XOR U3937 ( .A(n4294), .B(n4295), .Z(n4290) );
  AND U3938 ( .A(n4296), .B(n4297), .Z(n4295) );
  XNOR U3939 ( .A(p_input[3827]), .B(n4294), .Z(n4297) );
  XOR U3940 ( .A(n4294), .B(p_input[3795]), .Z(n4296) );
  XOR U3941 ( .A(n4298), .B(n4299), .Z(n4294) );
  AND U3942 ( .A(n4300), .B(n4301), .Z(n4299) );
  XNOR U3943 ( .A(p_input[3826]), .B(n4298), .Z(n4301) );
  XOR U3944 ( .A(n4298), .B(p_input[3794]), .Z(n4300) );
  XOR U3945 ( .A(n4302), .B(n4303), .Z(n4298) );
  AND U3946 ( .A(n4304), .B(n4305), .Z(n4303) );
  XNOR U3947 ( .A(p_input[3825]), .B(n4302), .Z(n4305) );
  XOR U3948 ( .A(n4302), .B(p_input[3793]), .Z(n4304) );
  XOR U3949 ( .A(n4306), .B(n4307), .Z(n4302) );
  AND U3950 ( .A(n4308), .B(n4309), .Z(n4307) );
  XNOR U3951 ( .A(p_input[3824]), .B(n4306), .Z(n4309) );
  XOR U3952 ( .A(n4306), .B(p_input[3792]), .Z(n4308) );
  XOR U3953 ( .A(n4310), .B(n4311), .Z(n4306) );
  AND U3954 ( .A(n4312), .B(n4313), .Z(n4311) );
  XNOR U3955 ( .A(p_input[3823]), .B(n4310), .Z(n4313) );
  XOR U3956 ( .A(n4310), .B(p_input[3791]), .Z(n4312) );
  XOR U3957 ( .A(n4314), .B(n4315), .Z(n4310) );
  AND U3958 ( .A(n4316), .B(n4317), .Z(n4315) );
  XNOR U3959 ( .A(p_input[3822]), .B(n4314), .Z(n4317) );
  XOR U3960 ( .A(n4314), .B(p_input[3790]), .Z(n4316) );
  XOR U3961 ( .A(n4318), .B(n4319), .Z(n4314) );
  AND U3962 ( .A(n4320), .B(n4321), .Z(n4319) );
  XNOR U3963 ( .A(p_input[3821]), .B(n4318), .Z(n4321) );
  XOR U3964 ( .A(n4318), .B(p_input[3789]), .Z(n4320) );
  XOR U3965 ( .A(n4322), .B(n4323), .Z(n4318) );
  AND U3966 ( .A(n4324), .B(n4325), .Z(n4323) );
  XNOR U3967 ( .A(p_input[3820]), .B(n4322), .Z(n4325) );
  XOR U3968 ( .A(n4322), .B(p_input[3788]), .Z(n4324) );
  XOR U3969 ( .A(n4326), .B(n4327), .Z(n4322) );
  AND U3970 ( .A(n4328), .B(n4329), .Z(n4327) );
  XNOR U3971 ( .A(p_input[3819]), .B(n4326), .Z(n4329) );
  XOR U3972 ( .A(n4326), .B(p_input[3787]), .Z(n4328) );
  XOR U3973 ( .A(n4330), .B(n4331), .Z(n4326) );
  AND U3974 ( .A(n4332), .B(n4333), .Z(n4331) );
  XNOR U3975 ( .A(p_input[3818]), .B(n4330), .Z(n4333) );
  XOR U3976 ( .A(n4330), .B(p_input[3786]), .Z(n4332) );
  XOR U3977 ( .A(n4334), .B(n4335), .Z(n4330) );
  AND U3978 ( .A(n4336), .B(n4337), .Z(n4335) );
  XNOR U3979 ( .A(p_input[3817]), .B(n4334), .Z(n4337) );
  XOR U3980 ( .A(n4334), .B(p_input[3785]), .Z(n4336) );
  XOR U3981 ( .A(n4338), .B(n4339), .Z(n4334) );
  AND U3982 ( .A(n4340), .B(n4341), .Z(n4339) );
  XNOR U3983 ( .A(p_input[3816]), .B(n4338), .Z(n4341) );
  XOR U3984 ( .A(n4338), .B(p_input[3784]), .Z(n4340) );
  XOR U3985 ( .A(n4342), .B(n4343), .Z(n4338) );
  AND U3986 ( .A(n4344), .B(n4345), .Z(n4343) );
  XNOR U3987 ( .A(p_input[3815]), .B(n4342), .Z(n4345) );
  XOR U3988 ( .A(n4342), .B(p_input[3783]), .Z(n4344) );
  XOR U3989 ( .A(n4346), .B(n4347), .Z(n4342) );
  AND U3990 ( .A(n4348), .B(n4349), .Z(n4347) );
  XNOR U3991 ( .A(p_input[3814]), .B(n4346), .Z(n4349) );
  XOR U3992 ( .A(n4346), .B(p_input[3782]), .Z(n4348) );
  XOR U3993 ( .A(n4350), .B(n4351), .Z(n4346) );
  AND U3994 ( .A(n4352), .B(n4353), .Z(n4351) );
  XNOR U3995 ( .A(p_input[3813]), .B(n4350), .Z(n4353) );
  XOR U3996 ( .A(n4350), .B(p_input[3781]), .Z(n4352) );
  XOR U3997 ( .A(n4354), .B(n4355), .Z(n4350) );
  AND U3998 ( .A(n4356), .B(n4357), .Z(n4355) );
  XNOR U3999 ( .A(p_input[3812]), .B(n4354), .Z(n4357) );
  XOR U4000 ( .A(n4354), .B(p_input[3780]), .Z(n4356) );
  XOR U4001 ( .A(n4358), .B(n4359), .Z(n4354) );
  AND U4002 ( .A(n4360), .B(n4361), .Z(n4359) );
  XNOR U4003 ( .A(p_input[3811]), .B(n4358), .Z(n4361) );
  XOR U4004 ( .A(n4358), .B(p_input[3779]), .Z(n4360) );
  XOR U4005 ( .A(n4362), .B(n4363), .Z(n4358) );
  AND U4006 ( .A(n4364), .B(n4365), .Z(n4363) );
  XNOR U4007 ( .A(p_input[3810]), .B(n4362), .Z(n4365) );
  XOR U4008 ( .A(n4362), .B(p_input[3778]), .Z(n4364) );
  XNOR U4009 ( .A(n4366), .B(n4367), .Z(n4362) );
  AND U4010 ( .A(n4368), .B(n4369), .Z(n4367) );
  XOR U4011 ( .A(p_input[3809]), .B(n4366), .Z(n4369) );
  XNOR U4012 ( .A(p_input[3777]), .B(n4366), .Z(n4368) );
  AND U4013 ( .A(p_input[3808]), .B(n4370), .Z(n4366) );
  IV U4014 ( .A(p_input[3776]), .Z(n4370) );
  XNOR U4015 ( .A(p_input[3712]), .B(n4371), .Z(n3964) );
  AND U4016 ( .A(n192), .B(n4372), .Z(n4371) );
  XOR U4017 ( .A(p_input[3744]), .B(p_input[3712]), .Z(n4372) );
  XOR U4018 ( .A(n4373), .B(n4374), .Z(n192) );
  AND U4019 ( .A(n4375), .B(n4376), .Z(n4374) );
  XNOR U4020 ( .A(p_input[3775]), .B(n4373), .Z(n4376) );
  XOR U4021 ( .A(n4373), .B(p_input[3743]), .Z(n4375) );
  XOR U4022 ( .A(n4377), .B(n4378), .Z(n4373) );
  AND U4023 ( .A(n4379), .B(n4380), .Z(n4378) );
  XNOR U4024 ( .A(p_input[3774]), .B(n4377), .Z(n4380) );
  XNOR U4025 ( .A(n4377), .B(n3979), .Z(n4379) );
  IV U4026 ( .A(p_input[3742]), .Z(n3979) );
  XOR U4027 ( .A(n4381), .B(n4382), .Z(n4377) );
  AND U4028 ( .A(n4383), .B(n4384), .Z(n4382) );
  XNOR U4029 ( .A(p_input[3773]), .B(n4381), .Z(n4384) );
  XNOR U4030 ( .A(n4381), .B(n3988), .Z(n4383) );
  IV U4031 ( .A(p_input[3741]), .Z(n3988) );
  XOR U4032 ( .A(n4385), .B(n4386), .Z(n4381) );
  AND U4033 ( .A(n4387), .B(n4388), .Z(n4386) );
  XNOR U4034 ( .A(p_input[3772]), .B(n4385), .Z(n4388) );
  XNOR U4035 ( .A(n4385), .B(n3997), .Z(n4387) );
  IV U4036 ( .A(p_input[3740]), .Z(n3997) );
  XOR U4037 ( .A(n4389), .B(n4390), .Z(n4385) );
  AND U4038 ( .A(n4391), .B(n4392), .Z(n4390) );
  XNOR U4039 ( .A(p_input[3771]), .B(n4389), .Z(n4392) );
  XNOR U4040 ( .A(n4389), .B(n4006), .Z(n4391) );
  IV U4041 ( .A(p_input[3739]), .Z(n4006) );
  XOR U4042 ( .A(n4393), .B(n4394), .Z(n4389) );
  AND U4043 ( .A(n4395), .B(n4396), .Z(n4394) );
  XNOR U4044 ( .A(p_input[3770]), .B(n4393), .Z(n4396) );
  XNOR U4045 ( .A(n4393), .B(n4015), .Z(n4395) );
  IV U4046 ( .A(p_input[3738]), .Z(n4015) );
  XOR U4047 ( .A(n4397), .B(n4398), .Z(n4393) );
  AND U4048 ( .A(n4399), .B(n4400), .Z(n4398) );
  XNOR U4049 ( .A(p_input[3769]), .B(n4397), .Z(n4400) );
  XNOR U4050 ( .A(n4397), .B(n4024), .Z(n4399) );
  IV U4051 ( .A(p_input[3737]), .Z(n4024) );
  XOR U4052 ( .A(n4401), .B(n4402), .Z(n4397) );
  AND U4053 ( .A(n4403), .B(n4404), .Z(n4402) );
  XNOR U4054 ( .A(p_input[3768]), .B(n4401), .Z(n4404) );
  XNOR U4055 ( .A(n4401), .B(n4033), .Z(n4403) );
  IV U4056 ( .A(p_input[3736]), .Z(n4033) );
  XOR U4057 ( .A(n4405), .B(n4406), .Z(n4401) );
  AND U4058 ( .A(n4407), .B(n4408), .Z(n4406) );
  XNOR U4059 ( .A(p_input[3767]), .B(n4405), .Z(n4408) );
  XNOR U4060 ( .A(n4405), .B(n4042), .Z(n4407) );
  IV U4061 ( .A(p_input[3735]), .Z(n4042) );
  XOR U4062 ( .A(n4409), .B(n4410), .Z(n4405) );
  AND U4063 ( .A(n4411), .B(n4412), .Z(n4410) );
  XNOR U4064 ( .A(p_input[3766]), .B(n4409), .Z(n4412) );
  XNOR U4065 ( .A(n4409), .B(n4051), .Z(n4411) );
  IV U4066 ( .A(p_input[3734]), .Z(n4051) );
  XOR U4067 ( .A(n4413), .B(n4414), .Z(n4409) );
  AND U4068 ( .A(n4415), .B(n4416), .Z(n4414) );
  XNOR U4069 ( .A(p_input[3765]), .B(n4413), .Z(n4416) );
  XNOR U4070 ( .A(n4413), .B(n4060), .Z(n4415) );
  IV U4071 ( .A(p_input[3733]), .Z(n4060) );
  XOR U4072 ( .A(n4417), .B(n4418), .Z(n4413) );
  AND U4073 ( .A(n4419), .B(n4420), .Z(n4418) );
  XNOR U4074 ( .A(p_input[3764]), .B(n4417), .Z(n4420) );
  XNOR U4075 ( .A(n4417), .B(n4069), .Z(n4419) );
  IV U4076 ( .A(p_input[3732]), .Z(n4069) );
  XOR U4077 ( .A(n4421), .B(n4422), .Z(n4417) );
  AND U4078 ( .A(n4423), .B(n4424), .Z(n4422) );
  XNOR U4079 ( .A(p_input[3763]), .B(n4421), .Z(n4424) );
  XNOR U4080 ( .A(n4421), .B(n4078), .Z(n4423) );
  IV U4081 ( .A(p_input[3731]), .Z(n4078) );
  XOR U4082 ( .A(n4425), .B(n4426), .Z(n4421) );
  AND U4083 ( .A(n4427), .B(n4428), .Z(n4426) );
  XNOR U4084 ( .A(p_input[3762]), .B(n4425), .Z(n4428) );
  XNOR U4085 ( .A(n4425), .B(n4087), .Z(n4427) );
  IV U4086 ( .A(p_input[3730]), .Z(n4087) );
  XOR U4087 ( .A(n4429), .B(n4430), .Z(n4425) );
  AND U4088 ( .A(n4431), .B(n4432), .Z(n4430) );
  XNOR U4089 ( .A(p_input[3761]), .B(n4429), .Z(n4432) );
  XNOR U4090 ( .A(n4429), .B(n4096), .Z(n4431) );
  IV U4091 ( .A(p_input[3729]), .Z(n4096) );
  XOR U4092 ( .A(n4433), .B(n4434), .Z(n4429) );
  AND U4093 ( .A(n4435), .B(n4436), .Z(n4434) );
  XNOR U4094 ( .A(p_input[3760]), .B(n4433), .Z(n4436) );
  XNOR U4095 ( .A(n4433), .B(n4105), .Z(n4435) );
  IV U4096 ( .A(p_input[3728]), .Z(n4105) );
  XOR U4097 ( .A(n4437), .B(n4438), .Z(n4433) );
  AND U4098 ( .A(n4439), .B(n4440), .Z(n4438) );
  XNOR U4099 ( .A(p_input[3759]), .B(n4437), .Z(n4440) );
  XNOR U4100 ( .A(n4437), .B(n4114), .Z(n4439) );
  IV U4101 ( .A(p_input[3727]), .Z(n4114) );
  XOR U4102 ( .A(n4441), .B(n4442), .Z(n4437) );
  AND U4103 ( .A(n4443), .B(n4444), .Z(n4442) );
  XNOR U4104 ( .A(p_input[3758]), .B(n4441), .Z(n4444) );
  XNOR U4105 ( .A(n4441), .B(n4123), .Z(n4443) );
  IV U4106 ( .A(p_input[3726]), .Z(n4123) );
  XOR U4107 ( .A(n4445), .B(n4446), .Z(n4441) );
  AND U4108 ( .A(n4447), .B(n4448), .Z(n4446) );
  XNOR U4109 ( .A(p_input[3757]), .B(n4445), .Z(n4448) );
  XNOR U4110 ( .A(n4445), .B(n4132), .Z(n4447) );
  IV U4111 ( .A(p_input[3725]), .Z(n4132) );
  XOR U4112 ( .A(n4449), .B(n4450), .Z(n4445) );
  AND U4113 ( .A(n4451), .B(n4452), .Z(n4450) );
  XNOR U4114 ( .A(p_input[3756]), .B(n4449), .Z(n4452) );
  XNOR U4115 ( .A(n4449), .B(n4141), .Z(n4451) );
  IV U4116 ( .A(p_input[3724]), .Z(n4141) );
  XOR U4117 ( .A(n4453), .B(n4454), .Z(n4449) );
  AND U4118 ( .A(n4455), .B(n4456), .Z(n4454) );
  XNOR U4119 ( .A(p_input[3755]), .B(n4453), .Z(n4456) );
  XNOR U4120 ( .A(n4453), .B(n4150), .Z(n4455) );
  IV U4121 ( .A(p_input[3723]), .Z(n4150) );
  XOR U4122 ( .A(n4457), .B(n4458), .Z(n4453) );
  AND U4123 ( .A(n4459), .B(n4460), .Z(n4458) );
  XNOR U4124 ( .A(p_input[3754]), .B(n4457), .Z(n4460) );
  XNOR U4125 ( .A(n4457), .B(n4159), .Z(n4459) );
  IV U4126 ( .A(p_input[3722]), .Z(n4159) );
  XOR U4127 ( .A(n4461), .B(n4462), .Z(n4457) );
  AND U4128 ( .A(n4463), .B(n4464), .Z(n4462) );
  XNOR U4129 ( .A(p_input[3753]), .B(n4461), .Z(n4464) );
  XNOR U4130 ( .A(n4461), .B(n4168), .Z(n4463) );
  IV U4131 ( .A(p_input[3721]), .Z(n4168) );
  XOR U4132 ( .A(n4465), .B(n4466), .Z(n4461) );
  AND U4133 ( .A(n4467), .B(n4468), .Z(n4466) );
  XNOR U4134 ( .A(p_input[3752]), .B(n4465), .Z(n4468) );
  XNOR U4135 ( .A(n4465), .B(n4177), .Z(n4467) );
  IV U4136 ( .A(p_input[3720]), .Z(n4177) );
  XOR U4137 ( .A(n4469), .B(n4470), .Z(n4465) );
  AND U4138 ( .A(n4471), .B(n4472), .Z(n4470) );
  XNOR U4139 ( .A(p_input[3751]), .B(n4469), .Z(n4472) );
  XNOR U4140 ( .A(n4469), .B(n4186), .Z(n4471) );
  IV U4141 ( .A(p_input[3719]), .Z(n4186) );
  XOR U4142 ( .A(n4473), .B(n4474), .Z(n4469) );
  AND U4143 ( .A(n4475), .B(n4476), .Z(n4474) );
  XNOR U4144 ( .A(p_input[3750]), .B(n4473), .Z(n4476) );
  XNOR U4145 ( .A(n4473), .B(n4195), .Z(n4475) );
  IV U4146 ( .A(p_input[3718]), .Z(n4195) );
  XOR U4147 ( .A(n4477), .B(n4478), .Z(n4473) );
  AND U4148 ( .A(n4479), .B(n4480), .Z(n4478) );
  XNOR U4149 ( .A(p_input[3749]), .B(n4477), .Z(n4480) );
  XNOR U4150 ( .A(n4477), .B(n4204), .Z(n4479) );
  IV U4151 ( .A(p_input[3717]), .Z(n4204) );
  XOR U4152 ( .A(n4481), .B(n4482), .Z(n4477) );
  AND U4153 ( .A(n4483), .B(n4484), .Z(n4482) );
  XNOR U4154 ( .A(p_input[3748]), .B(n4481), .Z(n4484) );
  XNOR U4155 ( .A(n4481), .B(n4213), .Z(n4483) );
  IV U4156 ( .A(p_input[3716]), .Z(n4213) );
  XOR U4157 ( .A(n4485), .B(n4486), .Z(n4481) );
  AND U4158 ( .A(n4487), .B(n4488), .Z(n4486) );
  XNOR U4159 ( .A(p_input[3747]), .B(n4485), .Z(n4488) );
  XNOR U4160 ( .A(n4485), .B(n4222), .Z(n4487) );
  IV U4161 ( .A(p_input[3715]), .Z(n4222) );
  XOR U4162 ( .A(n4489), .B(n4490), .Z(n4485) );
  AND U4163 ( .A(n4491), .B(n4492), .Z(n4490) );
  XNOR U4164 ( .A(p_input[3746]), .B(n4489), .Z(n4492) );
  XNOR U4165 ( .A(n4489), .B(n4231), .Z(n4491) );
  IV U4166 ( .A(p_input[3714]), .Z(n4231) );
  XNOR U4167 ( .A(n4493), .B(n4494), .Z(n4489) );
  AND U4168 ( .A(n4495), .B(n4496), .Z(n4494) );
  XOR U4169 ( .A(p_input[3745]), .B(n4493), .Z(n4496) );
  XNOR U4170 ( .A(p_input[3713]), .B(n4493), .Z(n4495) );
  AND U4171 ( .A(p_input[3744]), .B(n4497), .Z(n4493) );
  IV U4172 ( .A(p_input[3712]), .Z(n4497) );
  XOR U4173 ( .A(n4498), .B(n4499), .Z(n3587) );
  AND U4174 ( .A(n307), .B(n4500), .Z(n4499) );
  XNOR U4175 ( .A(n4501), .B(n4498), .Z(n4500) );
  XOR U4176 ( .A(n4502), .B(n4503), .Z(n307) );
  AND U4177 ( .A(n4504), .B(n4505), .Z(n4503) );
  XNOR U4178 ( .A(n3602), .B(n4502), .Z(n4505) );
  AND U4179 ( .A(p_input[3711]), .B(p_input[3679]), .Z(n3602) );
  XNOR U4180 ( .A(n4502), .B(n3599), .Z(n4504) );
  IV U4181 ( .A(n4506), .Z(n3599) );
  AND U4182 ( .A(p_input[3615]), .B(p_input[3647]), .Z(n4506) );
  XOR U4183 ( .A(n4507), .B(n4508), .Z(n4502) );
  AND U4184 ( .A(n4509), .B(n4510), .Z(n4508) );
  XOR U4185 ( .A(n4507), .B(n3614), .Z(n4510) );
  XNOR U4186 ( .A(p_input[3678]), .B(n4511), .Z(n3614) );
  AND U4187 ( .A(n198), .B(n4512), .Z(n4511) );
  XOR U4188 ( .A(p_input[3710]), .B(p_input[3678]), .Z(n4512) );
  XNOR U4189 ( .A(n3611), .B(n4507), .Z(n4509) );
  XOR U4190 ( .A(n4513), .B(n4514), .Z(n3611) );
  AND U4191 ( .A(n195), .B(n4515), .Z(n4514) );
  XOR U4192 ( .A(p_input[3646]), .B(p_input[3614]), .Z(n4515) );
  XOR U4193 ( .A(n4516), .B(n4517), .Z(n4507) );
  AND U4194 ( .A(n4518), .B(n4519), .Z(n4517) );
  XOR U4195 ( .A(n4516), .B(n3626), .Z(n4519) );
  XNOR U4196 ( .A(p_input[3677]), .B(n4520), .Z(n3626) );
  AND U4197 ( .A(n198), .B(n4521), .Z(n4520) );
  XOR U4198 ( .A(p_input[3709]), .B(p_input[3677]), .Z(n4521) );
  XNOR U4199 ( .A(n3623), .B(n4516), .Z(n4518) );
  XOR U4200 ( .A(n4522), .B(n4523), .Z(n3623) );
  AND U4201 ( .A(n195), .B(n4524), .Z(n4523) );
  XOR U4202 ( .A(p_input[3645]), .B(p_input[3613]), .Z(n4524) );
  XOR U4203 ( .A(n4525), .B(n4526), .Z(n4516) );
  AND U4204 ( .A(n4527), .B(n4528), .Z(n4526) );
  XOR U4205 ( .A(n4525), .B(n3638), .Z(n4528) );
  XNOR U4206 ( .A(p_input[3676]), .B(n4529), .Z(n3638) );
  AND U4207 ( .A(n198), .B(n4530), .Z(n4529) );
  XOR U4208 ( .A(p_input[3708]), .B(p_input[3676]), .Z(n4530) );
  XNOR U4209 ( .A(n3635), .B(n4525), .Z(n4527) );
  XOR U4210 ( .A(n4531), .B(n4532), .Z(n3635) );
  AND U4211 ( .A(n195), .B(n4533), .Z(n4532) );
  XOR U4212 ( .A(p_input[3644]), .B(p_input[3612]), .Z(n4533) );
  XOR U4213 ( .A(n4534), .B(n4535), .Z(n4525) );
  AND U4214 ( .A(n4536), .B(n4537), .Z(n4535) );
  XOR U4215 ( .A(n4534), .B(n3650), .Z(n4537) );
  XNOR U4216 ( .A(p_input[3675]), .B(n4538), .Z(n3650) );
  AND U4217 ( .A(n198), .B(n4539), .Z(n4538) );
  XOR U4218 ( .A(p_input[3707]), .B(p_input[3675]), .Z(n4539) );
  XNOR U4219 ( .A(n3647), .B(n4534), .Z(n4536) );
  XOR U4220 ( .A(n4540), .B(n4541), .Z(n3647) );
  AND U4221 ( .A(n195), .B(n4542), .Z(n4541) );
  XOR U4222 ( .A(p_input[3643]), .B(p_input[3611]), .Z(n4542) );
  XOR U4223 ( .A(n4543), .B(n4544), .Z(n4534) );
  AND U4224 ( .A(n4545), .B(n4546), .Z(n4544) );
  XOR U4225 ( .A(n4543), .B(n3662), .Z(n4546) );
  XNOR U4226 ( .A(p_input[3674]), .B(n4547), .Z(n3662) );
  AND U4227 ( .A(n198), .B(n4548), .Z(n4547) );
  XOR U4228 ( .A(p_input[3706]), .B(p_input[3674]), .Z(n4548) );
  XNOR U4229 ( .A(n3659), .B(n4543), .Z(n4545) );
  XOR U4230 ( .A(n4549), .B(n4550), .Z(n3659) );
  AND U4231 ( .A(n195), .B(n4551), .Z(n4550) );
  XOR U4232 ( .A(p_input[3642]), .B(p_input[3610]), .Z(n4551) );
  XOR U4233 ( .A(n4552), .B(n4553), .Z(n4543) );
  AND U4234 ( .A(n4554), .B(n4555), .Z(n4553) );
  XOR U4235 ( .A(n4552), .B(n3674), .Z(n4555) );
  XNOR U4236 ( .A(p_input[3673]), .B(n4556), .Z(n3674) );
  AND U4237 ( .A(n198), .B(n4557), .Z(n4556) );
  XOR U4238 ( .A(p_input[3705]), .B(p_input[3673]), .Z(n4557) );
  XNOR U4239 ( .A(n3671), .B(n4552), .Z(n4554) );
  XOR U4240 ( .A(n4558), .B(n4559), .Z(n3671) );
  AND U4241 ( .A(n195), .B(n4560), .Z(n4559) );
  XOR U4242 ( .A(p_input[3641]), .B(p_input[3609]), .Z(n4560) );
  XOR U4243 ( .A(n4561), .B(n4562), .Z(n4552) );
  AND U4244 ( .A(n4563), .B(n4564), .Z(n4562) );
  XOR U4245 ( .A(n4561), .B(n3686), .Z(n4564) );
  XNOR U4246 ( .A(p_input[3672]), .B(n4565), .Z(n3686) );
  AND U4247 ( .A(n198), .B(n4566), .Z(n4565) );
  XOR U4248 ( .A(p_input[3704]), .B(p_input[3672]), .Z(n4566) );
  XNOR U4249 ( .A(n3683), .B(n4561), .Z(n4563) );
  XOR U4250 ( .A(n4567), .B(n4568), .Z(n3683) );
  AND U4251 ( .A(n195), .B(n4569), .Z(n4568) );
  XOR U4252 ( .A(p_input[3640]), .B(p_input[3608]), .Z(n4569) );
  XOR U4253 ( .A(n4570), .B(n4571), .Z(n4561) );
  AND U4254 ( .A(n4572), .B(n4573), .Z(n4571) );
  XOR U4255 ( .A(n4570), .B(n3698), .Z(n4573) );
  XNOR U4256 ( .A(p_input[3671]), .B(n4574), .Z(n3698) );
  AND U4257 ( .A(n198), .B(n4575), .Z(n4574) );
  XOR U4258 ( .A(p_input[3703]), .B(p_input[3671]), .Z(n4575) );
  XNOR U4259 ( .A(n3695), .B(n4570), .Z(n4572) );
  XOR U4260 ( .A(n4576), .B(n4577), .Z(n3695) );
  AND U4261 ( .A(n195), .B(n4578), .Z(n4577) );
  XOR U4262 ( .A(p_input[3639]), .B(p_input[3607]), .Z(n4578) );
  XOR U4263 ( .A(n4579), .B(n4580), .Z(n4570) );
  AND U4264 ( .A(n4581), .B(n4582), .Z(n4580) );
  XOR U4265 ( .A(n4579), .B(n3710), .Z(n4582) );
  XNOR U4266 ( .A(p_input[3670]), .B(n4583), .Z(n3710) );
  AND U4267 ( .A(n198), .B(n4584), .Z(n4583) );
  XOR U4268 ( .A(p_input[3702]), .B(p_input[3670]), .Z(n4584) );
  XNOR U4269 ( .A(n3707), .B(n4579), .Z(n4581) );
  XOR U4270 ( .A(n4585), .B(n4586), .Z(n3707) );
  AND U4271 ( .A(n195), .B(n4587), .Z(n4586) );
  XOR U4272 ( .A(p_input[3638]), .B(p_input[3606]), .Z(n4587) );
  XOR U4273 ( .A(n4588), .B(n4589), .Z(n4579) );
  AND U4274 ( .A(n4590), .B(n4591), .Z(n4589) );
  XOR U4275 ( .A(n4588), .B(n3722), .Z(n4591) );
  XNOR U4276 ( .A(p_input[3669]), .B(n4592), .Z(n3722) );
  AND U4277 ( .A(n198), .B(n4593), .Z(n4592) );
  XOR U4278 ( .A(p_input[3701]), .B(p_input[3669]), .Z(n4593) );
  XNOR U4279 ( .A(n3719), .B(n4588), .Z(n4590) );
  XOR U4280 ( .A(n4594), .B(n4595), .Z(n3719) );
  AND U4281 ( .A(n195), .B(n4596), .Z(n4595) );
  XOR U4282 ( .A(p_input[3637]), .B(p_input[3605]), .Z(n4596) );
  XOR U4283 ( .A(n4597), .B(n4598), .Z(n4588) );
  AND U4284 ( .A(n4599), .B(n4600), .Z(n4598) );
  XOR U4285 ( .A(n4597), .B(n3734), .Z(n4600) );
  XNOR U4286 ( .A(p_input[3668]), .B(n4601), .Z(n3734) );
  AND U4287 ( .A(n198), .B(n4602), .Z(n4601) );
  XOR U4288 ( .A(p_input[3700]), .B(p_input[3668]), .Z(n4602) );
  XNOR U4289 ( .A(n3731), .B(n4597), .Z(n4599) );
  XOR U4290 ( .A(n4603), .B(n4604), .Z(n3731) );
  AND U4291 ( .A(n195), .B(n4605), .Z(n4604) );
  XOR U4292 ( .A(p_input[3636]), .B(p_input[3604]), .Z(n4605) );
  XOR U4293 ( .A(n4606), .B(n4607), .Z(n4597) );
  AND U4294 ( .A(n4608), .B(n4609), .Z(n4607) );
  XOR U4295 ( .A(n4606), .B(n3746), .Z(n4609) );
  XNOR U4296 ( .A(p_input[3667]), .B(n4610), .Z(n3746) );
  AND U4297 ( .A(n198), .B(n4611), .Z(n4610) );
  XOR U4298 ( .A(p_input[3699]), .B(p_input[3667]), .Z(n4611) );
  XNOR U4299 ( .A(n3743), .B(n4606), .Z(n4608) );
  XOR U4300 ( .A(n4612), .B(n4613), .Z(n3743) );
  AND U4301 ( .A(n195), .B(n4614), .Z(n4613) );
  XOR U4302 ( .A(p_input[3635]), .B(p_input[3603]), .Z(n4614) );
  XOR U4303 ( .A(n4615), .B(n4616), .Z(n4606) );
  AND U4304 ( .A(n4617), .B(n4618), .Z(n4616) );
  XOR U4305 ( .A(n4615), .B(n3758), .Z(n4618) );
  XNOR U4306 ( .A(p_input[3666]), .B(n4619), .Z(n3758) );
  AND U4307 ( .A(n198), .B(n4620), .Z(n4619) );
  XOR U4308 ( .A(p_input[3698]), .B(p_input[3666]), .Z(n4620) );
  XNOR U4309 ( .A(n3755), .B(n4615), .Z(n4617) );
  XOR U4310 ( .A(n4621), .B(n4622), .Z(n3755) );
  AND U4311 ( .A(n195), .B(n4623), .Z(n4622) );
  XOR U4312 ( .A(p_input[3634]), .B(p_input[3602]), .Z(n4623) );
  XOR U4313 ( .A(n4624), .B(n4625), .Z(n4615) );
  AND U4314 ( .A(n4626), .B(n4627), .Z(n4625) );
  XOR U4315 ( .A(n4624), .B(n3770), .Z(n4627) );
  XNOR U4316 ( .A(p_input[3665]), .B(n4628), .Z(n3770) );
  AND U4317 ( .A(n198), .B(n4629), .Z(n4628) );
  XOR U4318 ( .A(p_input[3697]), .B(p_input[3665]), .Z(n4629) );
  XNOR U4319 ( .A(n3767), .B(n4624), .Z(n4626) );
  XOR U4320 ( .A(n4630), .B(n4631), .Z(n3767) );
  AND U4321 ( .A(n195), .B(n4632), .Z(n4631) );
  XOR U4322 ( .A(p_input[3633]), .B(p_input[3601]), .Z(n4632) );
  XOR U4323 ( .A(n4633), .B(n4634), .Z(n4624) );
  AND U4324 ( .A(n4635), .B(n4636), .Z(n4634) );
  XOR U4325 ( .A(n4633), .B(n3782), .Z(n4636) );
  XNOR U4326 ( .A(p_input[3664]), .B(n4637), .Z(n3782) );
  AND U4327 ( .A(n198), .B(n4638), .Z(n4637) );
  XOR U4328 ( .A(p_input[3696]), .B(p_input[3664]), .Z(n4638) );
  XNOR U4329 ( .A(n3779), .B(n4633), .Z(n4635) );
  XOR U4330 ( .A(n4639), .B(n4640), .Z(n3779) );
  AND U4331 ( .A(n195), .B(n4641), .Z(n4640) );
  XOR U4332 ( .A(p_input[3632]), .B(p_input[3600]), .Z(n4641) );
  XOR U4333 ( .A(n4642), .B(n4643), .Z(n4633) );
  AND U4334 ( .A(n4644), .B(n4645), .Z(n4643) );
  XOR U4335 ( .A(n4642), .B(n3794), .Z(n4645) );
  XNOR U4336 ( .A(p_input[3663]), .B(n4646), .Z(n3794) );
  AND U4337 ( .A(n198), .B(n4647), .Z(n4646) );
  XOR U4338 ( .A(p_input[3695]), .B(p_input[3663]), .Z(n4647) );
  XNOR U4339 ( .A(n3791), .B(n4642), .Z(n4644) );
  XOR U4340 ( .A(n4648), .B(n4649), .Z(n3791) );
  AND U4341 ( .A(n195), .B(n4650), .Z(n4649) );
  XOR U4342 ( .A(p_input[3631]), .B(p_input[3599]), .Z(n4650) );
  XOR U4343 ( .A(n4651), .B(n4652), .Z(n4642) );
  AND U4344 ( .A(n4653), .B(n4654), .Z(n4652) );
  XOR U4345 ( .A(n4651), .B(n3806), .Z(n4654) );
  XNOR U4346 ( .A(p_input[3662]), .B(n4655), .Z(n3806) );
  AND U4347 ( .A(n198), .B(n4656), .Z(n4655) );
  XOR U4348 ( .A(p_input[3694]), .B(p_input[3662]), .Z(n4656) );
  XNOR U4349 ( .A(n3803), .B(n4651), .Z(n4653) );
  XOR U4350 ( .A(n4657), .B(n4658), .Z(n3803) );
  AND U4351 ( .A(n195), .B(n4659), .Z(n4658) );
  XOR U4352 ( .A(p_input[3630]), .B(p_input[3598]), .Z(n4659) );
  XOR U4353 ( .A(n4660), .B(n4661), .Z(n4651) );
  AND U4354 ( .A(n4662), .B(n4663), .Z(n4661) );
  XOR U4355 ( .A(n4660), .B(n3818), .Z(n4663) );
  XNOR U4356 ( .A(p_input[3661]), .B(n4664), .Z(n3818) );
  AND U4357 ( .A(n198), .B(n4665), .Z(n4664) );
  XOR U4358 ( .A(p_input[3693]), .B(p_input[3661]), .Z(n4665) );
  XNOR U4359 ( .A(n3815), .B(n4660), .Z(n4662) );
  XOR U4360 ( .A(n4666), .B(n4667), .Z(n3815) );
  AND U4361 ( .A(n195), .B(n4668), .Z(n4667) );
  XOR U4362 ( .A(p_input[3629]), .B(p_input[3597]), .Z(n4668) );
  XOR U4363 ( .A(n4669), .B(n4670), .Z(n4660) );
  AND U4364 ( .A(n4671), .B(n4672), .Z(n4670) );
  XOR U4365 ( .A(n4669), .B(n3830), .Z(n4672) );
  XNOR U4366 ( .A(p_input[3660]), .B(n4673), .Z(n3830) );
  AND U4367 ( .A(n198), .B(n4674), .Z(n4673) );
  XOR U4368 ( .A(p_input[3692]), .B(p_input[3660]), .Z(n4674) );
  XNOR U4369 ( .A(n3827), .B(n4669), .Z(n4671) );
  XOR U4370 ( .A(n4675), .B(n4676), .Z(n3827) );
  AND U4371 ( .A(n195), .B(n4677), .Z(n4676) );
  XOR U4372 ( .A(p_input[3628]), .B(p_input[3596]), .Z(n4677) );
  XOR U4373 ( .A(n4678), .B(n4679), .Z(n4669) );
  AND U4374 ( .A(n4680), .B(n4681), .Z(n4679) );
  XOR U4375 ( .A(n4678), .B(n3842), .Z(n4681) );
  XNOR U4376 ( .A(p_input[3659]), .B(n4682), .Z(n3842) );
  AND U4377 ( .A(n198), .B(n4683), .Z(n4682) );
  XOR U4378 ( .A(p_input[3691]), .B(p_input[3659]), .Z(n4683) );
  XNOR U4379 ( .A(n3839), .B(n4678), .Z(n4680) );
  XOR U4380 ( .A(n4684), .B(n4685), .Z(n3839) );
  AND U4381 ( .A(n195), .B(n4686), .Z(n4685) );
  XOR U4382 ( .A(p_input[3627]), .B(p_input[3595]), .Z(n4686) );
  XOR U4383 ( .A(n4687), .B(n4688), .Z(n4678) );
  AND U4384 ( .A(n4689), .B(n4690), .Z(n4688) );
  XOR U4385 ( .A(n4687), .B(n3854), .Z(n4690) );
  XNOR U4386 ( .A(p_input[3658]), .B(n4691), .Z(n3854) );
  AND U4387 ( .A(n198), .B(n4692), .Z(n4691) );
  XOR U4388 ( .A(p_input[3690]), .B(p_input[3658]), .Z(n4692) );
  XNOR U4389 ( .A(n3851), .B(n4687), .Z(n4689) );
  XOR U4390 ( .A(n4693), .B(n4694), .Z(n3851) );
  AND U4391 ( .A(n195), .B(n4695), .Z(n4694) );
  XOR U4392 ( .A(p_input[3626]), .B(p_input[3594]), .Z(n4695) );
  XOR U4393 ( .A(n4696), .B(n4697), .Z(n4687) );
  AND U4394 ( .A(n4698), .B(n4699), .Z(n4697) );
  XOR U4395 ( .A(n4696), .B(n3866), .Z(n4699) );
  XNOR U4396 ( .A(p_input[3657]), .B(n4700), .Z(n3866) );
  AND U4397 ( .A(n198), .B(n4701), .Z(n4700) );
  XOR U4398 ( .A(p_input[3689]), .B(p_input[3657]), .Z(n4701) );
  XNOR U4399 ( .A(n3863), .B(n4696), .Z(n4698) );
  XOR U4400 ( .A(n4702), .B(n4703), .Z(n3863) );
  AND U4401 ( .A(n195), .B(n4704), .Z(n4703) );
  XOR U4402 ( .A(p_input[3625]), .B(p_input[3593]), .Z(n4704) );
  XOR U4403 ( .A(n4705), .B(n4706), .Z(n4696) );
  AND U4404 ( .A(n4707), .B(n4708), .Z(n4706) );
  XOR U4405 ( .A(n4705), .B(n3878), .Z(n4708) );
  XNOR U4406 ( .A(p_input[3656]), .B(n4709), .Z(n3878) );
  AND U4407 ( .A(n198), .B(n4710), .Z(n4709) );
  XOR U4408 ( .A(p_input[3688]), .B(p_input[3656]), .Z(n4710) );
  XNOR U4409 ( .A(n3875), .B(n4705), .Z(n4707) );
  XOR U4410 ( .A(n4711), .B(n4712), .Z(n3875) );
  AND U4411 ( .A(n195), .B(n4713), .Z(n4712) );
  XOR U4412 ( .A(p_input[3624]), .B(p_input[3592]), .Z(n4713) );
  XOR U4413 ( .A(n4714), .B(n4715), .Z(n4705) );
  AND U4414 ( .A(n4716), .B(n4717), .Z(n4715) );
  XOR U4415 ( .A(n4714), .B(n3890), .Z(n4717) );
  XNOR U4416 ( .A(p_input[3655]), .B(n4718), .Z(n3890) );
  AND U4417 ( .A(n198), .B(n4719), .Z(n4718) );
  XOR U4418 ( .A(p_input[3687]), .B(p_input[3655]), .Z(n4719) );
  XNOR U4419 ( .A(n3887), .B(n4714), .Z(n4716) );
  XOR U4420 ( .A(n4720), .B(n4721), .Z(n3887) );
  AND U4421 ( .A(n195), .B(n4722), .Z(n4721) );
  XOR U4422 ( .A(p_input[3623]), .B(p_input[3591]), .Z(n4722) );
  XOR U4423 ( .A(n4723), .B(n4724), .Z(n4714) );
  AND U4424 ( .A(n4725), .B(n4726), .Z(n4724) );
  XOR U4425 ( .A(n4723), .B(n3902), .Z(n4726) );
  XNOR U4426 ( .A(p_input[3654]), .B(n4727), .Z(n3902) );
  AND U4427 ( .A(n198), .B(n4728), .Z(n4727) );
  XOR U4428 ( .A(p_input[3686]), .B(p_input[3654]), .Z(n4728) );
  XNOR U4429 ( .A(n3899), .B(n4723), .Z(n4725) );
  XOR U4430 ( .A(n4729), .B(n4730), .Z(n3899) );
  AND U4431 ( .A(n195), .B(n4731), .Z(n4730) );
  XOR U4432 ( .A(p_input[3622]), .B(p_input[3590]), .Z(n4731) );
  XOR U4433 ( .A(n4732), .B(n4733), .Z(n4723) );
  AND U4434 ( .A(n4734), .B(n4735), .Z(n4733) );
  XOR U4435 ( .A(n4732), .B(n3914), .Z(n4735) );
  XNOR U4436 ( .A(p_input[3653]), .B(n4736), .Z(n3914) );
  AND U4437 ( .A(n198), .B(n4737), .Z(n4736) );
  XOR U4438 ( .A(p_input[3685]), .B(p_input[3653]), .Z(n4737) );
  XNOR U4439 ( .A(n3911), .B(n4732), .Z(n4734) );
  XOR U4440 ( .A(n4738), .B(n4739), .Z(n3911) );
  AND U4441 ( .A(n195), .B(n4740), .Z(n4739) );
  XOR U4442 ( .A(p_input[3621]), .B(p_input[3589]), .Z(n4740) );
  XOR U4443 ( .A(n4741), .B(n4742), .Z(n4732) );
  AND U4444 ( .A(n4743), .B(n4744), .Z(n4742) );
  XOR U4445 ( .A(n4741), .B(n3926), .Z(n4744) );
  XNOR U4446 ( .A(p_input[3652]), .B(n4745), .Z(n3926) );
  AND U4447 ( .A(n198), .B(n4746), .Z(n4745) );
  XOR U4448 ( .A(p_input[3684]), .B(p_input[3652]), .Z(n4746) );
  XNOR U4449 ( .A(n3923), .B(n4741), .Z(n4743) );
  XOR U4450 ( .A(n4747), .B(n4748), .Z(n3923) );
  AND U4451 ( .A(n195), .B(n4749), .Z(n4748) );
  XOR U4452 ( .A(p_input[3620]), .B(p_input[3588]), .Z(n4749) );
  XOR U4453 ( .A(n4750), .B(n4751), .Z(n4741) );
  AND U4454 ( .A(n4752), .B(n4753), .Z(n4751) );
  XOR U4455 ( .A(n4750), .B(n3938), .Z(n4753) );
  XNOR U4456 ( .A(p_input[3651]), .B(n4754), .Z(n3938) );
  AND U4457 ( .A(n198), .B(n4755), .Z(n4754) );
  XOR U4458 ( .A(p_input[3683]), .B(p_input[3651]), .Z(n4755) );
  XNOR U4459 ( .A(n3935), .B(n4750), .Z(n4752) );
  XOR U4460 ( .A(n4756), .B(n4757), .Z(n3935) );
  AND U4461 ( .A(n195), .B(n4758), .Z(n4757) );
  XOR U4462 ( .A(p_input[3619]), .B(p_input[3587]), .Z(n4758) );
  XOR U4463 ( .A(n4759), .B(n4760), .Z(n4750) );
  AND U4464 ( .A(n4761), .B(n4762), .Z(n4760) );
  XOR U4465 ( .A(n3950), .B(n4759), .Z(n4762) );
  XNOR U4466 ( .A(p_input[3650]), .B(n4763), .Z(n3950) );
  AND U4467 ( .A(n198), .B(n4764), .Z(n4763) );
  XOR U4468 ( .A(p_input[3682]), .B(p_input[3650]), .Z(n4764) );
  XNOR U4469 ( .A(n4759), .B(n3947), .Z(n4761) );
  XOR U4470 ( .A(n4765), .B(n4766), .Z(n3947) );
  AND U4471 ( .A(n195), .B(n4767), .Z(n4766) );
  XOR U4472 ( .A(p_input[3618]), .B(p_input[3586]), .Z(n4767) );
  XOR U4473 ( .A(n4768), .B(n4769), .Z(n4759) );
  AND U4474 ( .A(n4770), .B(n4771), .Z(n4769) );
  XNOR U4475 ( .A(n4772), .B(n3963), .Z(n4771) );
  XNOR U4476 ( .A(p_input[3649]), .B(n4773), .Z(n3963) );
  AND U4477 ( .A(n198), .B(n4774), .Z(n4773) );
  XNOR U4478 ( .A(p_input[3681]), .B(n4775), .Z(n4774) );
  IV U4479 ( .A(p_input[3649]), .Z(n4775) );
  XNOR U4480 ( .A(n3960), .B(n4768), .Z(n4770) );
  XNOR U4481 ( .A(p_input[3585]), .B(n4776), .Z(n3960) );
  AND U4482 ( .A(n195), .B(n4777), .Z(n4776) );
  XOR U4483 ( .A(p_input[3617]), .B(p_input[3585]), .Z(n4777) );
  IV U4484 ( .A(n4772), .Z(n4768) );
  AND U4485 ( .A(n4498), .B(n4501), .Z(n4772) );
  XOR U4486 ( .A(p_input[3648]), .B(n4778), .Z(n4501) );
  AND U4487 ( .A(n198), .B(n4779), .Z(n4778) );
  XOR U4488 ( .A(p_input[3680]), .B(p_input[3648]), .Z(n4779) );
  XOR U4489 ( .A(n4780), .B(n4781), .Z(n198) );
  AND U4490 ( .A(n4782), .B(n4783), .Z(n4781) );
  XNOR U4491 ( .A(p_input[3711]), .B(n4780), .Z(n4783) );
  XOR U4492 ( .A(n4780), .B(p_input[3679]), .Z(n4782) );
  XOR U4493 ( .A(n4784), .B(n4785), .Z(n4780) );
  AND U4494 ( .A(n4786), .B(n4787), .Z(n4785) );
  XNOR U4495 ( .A(p_input[3710]), .B(n4784), .Z(n4787) );
  XOR U4496 ( .A(n4784), .B(p_input[3678]), .Z(n4786) );
  XOR U4497 ( .A(n4788), .B(n4789), .Z(n4784) );
  AND U4498 ( .A(n4790), .B(n4791), .Z(n4789) );
  XNOR U4499 ( .A(p_input[3709]), .B(n4788), .Z(n4791) );
  XOR U4500 ( .A(n4788), .B(p_input[3677]), .Z(n4790) );
  XOR U4501 ( .A(n4792), .B(n4793), .Z(n4788) );
  AND U4502 ( .A(n4794), .B(n4795), .Z(n4793) );
  XNOR U4503 ( .A(p_input[3708]), .B(n4792), .Z(n4795) );
  XOR U4504 ( .A(n4792), .B(p_input[3676]), .Z(n4794) );
  XOR U4505 ( .A(n4796), .B(n4797), .Z(n4792) );
  AND U4506 ( .A(n4798), .B(n4799), .Z(n4797) );
  XNOR U4507 ( .A(p_input[3707]), .B(n4796), .Z(n4799) );
  XOR U4508 ( .A(n4796), .B(p_input[3675]), .Z(n4798) );
  XOR U4509 ( .A(n4800), .B(n4801), .Z(n4796) );
  AND U4510 ( .A(n4802), .B(n4803), .Z(n4801) );
  XNOR U4511 ( .A(p_input[3706]), .B(n4800), .Z(n4803) );
  XOR U4512 ( .A(n4800), .B(p_input[3674]), .Z(n4802) );
  XOR U4513 ( .A(n4804), .B(n4805), .Z(n4800) );
  AND U4514 ( .A(n4806), .B(n4807), .Z(n4805) );
  XNOR U4515 ( .A(p_input[3705]), .B(n4804), .Z(n4807) );
  XOR U4516 ( .A(n4804), .B(p_input[3673]), .Z(n4806) );
  XOR U4517 ( .A(n4808), .B(n4809), .Z(n4804) );
  AND U4518 ( .A(n4810), .B(n4811), .Z(n4809) );
  XNOR U4519 ( .A(p_input[3704]), .B(n4808), .Z(n4811) );
  XOR U4520 ( .A(n4808), .B(p_input[3672]), .Z(n4810) );
  XOR U4521 ( .A(n4812), .B(n4813), .Z(n4808) );
  AND U4522 ( .A(n4814), .B(n4815), .Z(n4813) );
  XNOR U4523 ( .A(p_input[3703]), .B(n4812), .Z(n4815) );
  XOR U4524 ( .A(n4812), .B(p_input[3671]), .Z(n4814) );
  XOR U4525 ( .A(n4816), .B(n4817), .Z(n4812) );
  AND U4526 ( .A(n4818), .B(n4819), .Z(n4817) );
  XNOR U4527 ( .A(p_input[3702]), .B(n4816), .Z(n4819) );
  XOR U4528 ( .A(n4816), .B(p_input[3670]), .Z(n4818) );
  XOR U4529 ( .A(n4820), .B(n4821), .Z(n4816) );
  AND U4530 ( .A(n4822), .B(n4823), .Z(n4821) );
  XNOR U4531 ( .A(p_input[3701]), .B(n4820), .Z(n4823) );
  XOR U4532 ( .A(n4820), .B(p_input[3669]), .Z(n4822) );
  XOR U4533 ( .A(n4824), .B(n4825), .Z(n4820) );
  AND U4534 ( .A(n4826), .B(n4827), .Z(n4825) );
  XNOR U4535 ( .A(p_input[3700]), .B(n4824), .Z(n4827) );
  XOR U4536 ( .A(n4824), .B(p_input[3668]), .Z(n4826) );
  XOR U4537 ( .A(n4828), .B(n4829), .Z(n4824) );
  AND U4538 ( .A(n4830), .B(n4831), .Z(n4829) );
  XNOR U4539 ( .A(p_input[3699]), .B(n4828), .Z(n4831) );
  XOR U4540 ( .A(n4828), .B(p_input[3667]), .Z(n4830) );
  XOR U4541 ( .A(n4832), .B(n4833), .Z(n4828) );
  AND U4542 ( .A(n4834), .B(n4835), .Z(n4833) );
  XNOR U4543 ( .A(p_input[3698]), .B(n4832), .Z(n4835) );
  XOR U4544 ( .A(n4832), .B(p_input[3666]), .Z(n4834) );
  XOR U4545 ( .A(n4836), .B(n4837), .Z(n4832) );
  AND U4546 ( .A(n4838), .B(n4839), .Z(n4837) );
  XNOR U4547 ( .A(p_input[3697]), .B(n4836), .Z(n4839) );
  XOR U4548 ( .A(n4836), .B(p_input[3665]), .Z(n4838) );
  XOR U4549 ( .A(n4840), .B(n4841), .Z(n4836) );
  AND U4550 ( .A(n4842), .B(n4843), .Z(n4841) );
  XNOR U4551 ( .A(p_input[3696]), .B(n4840), .Z(n4843) );
  XOR U4552 ( .A(n4840), .B(p_input[3664]), .Z(n4842) );
  XOR U4553 ( .A(n4844), .B(n4845), .Z(n4840) );
  AND U4554 ( .A(n4846), .B(n4847), .Z(n4845) );
  XNOR U4555 ( .A(p_input[3695]), .B(n4844), .Z(n4847) );
  XOR U4556 ( .A(n4844), .B(p_input[3663]), .Z(n4846) );
  XOR U4557 ( .A(n4848), .B(n4849), .Z(n4844) );
  AND U4558 ( .A(n4850), .B(n4851), .Z(n4849) );
  XNOR U4559 ( .A(p_input[3694]), .B(n4848), .Z(n4851) );
  XOR U4560 ( .A(n4848), .B(p_input[3662]), .Z(n4850) );
  XOR U4561 ( .A(n4852), .B(n4853), .Z(n4848) );
  AND U4562 ( .A(n4854), .B(n4855), .Z(n4853) );
  XNOR U4563 ( .A(p_input[3693]), .B(n4852), .Z(n4855) );
  XOR U4564 ( .A(n4852), .B(p_input[3661]), .Z(n4854) );
  XOR U4565 ( .A(n4856), .B(n4857), .Z(n4852) );
  AND U4566 ( .A(n4858), .B(n4859), .Z(n4857) );
  XNOR U4567 ( .A(p_input[3692]), .B(n4856), .Z(n4859) );
  XOR U4568 ( .A(n4856), .B(p_input[3660]), .Z(n4858) );
  XOR U4569 ( .A(n4860), .B(n4861), .Z(n4856) );
  AND U4570 ( .A(n4862), .B(n4863), .Z(n4861) );
  XNOR U4571 ( .A(p_input[3691]), .B(n4860), .Z(n4863) );
  XOR U4572 ( .A(n4860), .B(p_input[3659]), .Z(n4862) );
  XOR U4573 ( .A(n4864), .B(n4865), .Z(n4860) );
  AND U4574 ( .A(n4866), .B(n4867), .Z(n4865) );
  XNOR U4575 ( .A(p_input[3690]), .B(n4864), .Z(n4867) );
  XOR U4576 ( .A(n4864), .B(p_input[3658]), .Z(n4866) );
  XOR U4577 ( .A(n4868), .B(n4869), .Z(n4864) );
  AND U4578 ( .A(n4870), .B(n4871), .Z(n4869) );
  XNOR U4579 ( .A(p_input[3689]), .B(n4868), .Z(n4871) );
  XOR U4580 ( .A(n4868), .B(p_input[3657]), .Z(n4870) );
  XOR U4581 ( .A(n4872), .B(n4873), .Z(n4868) );
  AND U4582 ( .A(n4874), .B(n4875), .Z(n4873) );
  XNOR U4583 ( .A(p_input[3688]), .B(n4872), .Z(n4875) );
  XOR U4584 ( .A(n4872), .B(p_input[3656]), .Z(n4874) );
  XOR U4585 ( .A(n4876), .B(n4877), .Z(n4872) );
  AND U4586 ( .A(n4878), .B(n4879), .Z(n4877) );
  XNOR U4587 ( .A(p_input[3687]), .B(n4876), .Z(n4879) );
  XOR U4588 ( .A(n4876), .B(p_input[3655]), .Z(n4878) );
  XOR U4589 ( .A(n4880), .B(n4881), .Z(n4876) );
  AND U4590 ( .A(n4882), .B(n4883), .Z(n4881) );
  XNOR U4591 ( .A(p_input[3686]), .B(n4880), .Z(n4883) );
  XOR U4592 ( .A(n4880), .B(p_input[3654]), .Z(n4882) );
  XOR U4593 ( .A(n4884), .B(n4885), .Z(n4880) );
  AND U4594 ( .A(n4886), .B(n4887), .Z(n4885) );
  XNOR U4595 ( .A(p_input[3685]), .B(n4884), .Z(n4887) );
  XOR U4596 ( .A(n4884), .B(p_input[3653]), .Z(n4886) );
  XOR U4597 ( .A(n4888), .B(n4889), .Z(n4884) );
  AND U4598 ( .A(n4890), .B(n4891), .Z(n4889) );
  XNOR U4599 ( .A(p_input[3684]), .B(n4888), .Z(n4891) );
  XOR U4600 ( .A(n4888), .B(p_input[3652]), .Z(n4890) );
  XOR U4601 ( .A(n4892), .B(n4893), .Z(n4888) );
  AND U4602 ( .A(n4894), .B(n4895), .Z(n4893) );
  XNOR U4603 ( .A(p_input[3683]), .B(n4892), .Z(n4895) );
  XOR U4604 ( .A(n4892), .B(p_input[3651]), .Z(n4894) );
  XOR U4605 ( .A(n4896), .B(n4897), .Z(n4892) );
  AND U4606 ( .A(n4898), .B(n4899), .Z(n4897) );
  XNOR U4607 ( .A(p_input[3682]), .B(n4896), .Z(n4899) );
  XOR U4608 ( .A(n4896), .B(p_input[3650]), .Z(n4898) );
  XNOR U4609 ( .A(n4900), .B(n4901), .Z(n4896) );
  AND U4610 ( .A(n4902), .B(n4903), .Z(n4901) );
  XOR U4611 ( .A(p_input[3681]), .B(n4900), .Z(n4903) );
  XNOR U4612 ( .A(p_input[3649]), .B(n4900), .Z(n4902) );
  AND U4613 ( .A(p_input[3680]), .B(n4904), .Z(n4900) );
  IV U4614 ( .A(p_input[3648]), .Z(n4904) );
  XNOR U4615 ( .A(p_input[3584]), .B(n4905), .Z(n4498) );
  AND U4616 ( .A(n195), .B(n4906), .Z(n4905) );
  XOR U4617 ( .A(p_input[3616]), .B(p_input[3584]), .Z(n4906) );
  XOR U4618 ( .A(n4907), .B(n4908), .Z(n195) );
  AND U4619 ( .A(n4909), .B(n4910), .Z(n4908) );
  XNOR U4620 ( .A(p_input[3647]), .B(n4907), .Z(n4910) );
  XOR U4621 ( .A(n4907), .B(p_input[3615]), .Z(n4909) );
  XOR U4622 ( .A(n4911), .B(n4912), .Z(n4907) );
  AND U4623 ( .A(n4913), .B(n4914), .Z(n4912) );
  XNOR U4624 ( .A(p_input[3646]), .B(n4911), .Z(n4914) );
  XNOR U4625 ( .A(n4911), .B(n4513), .Z(n4913) );
  IV U4626 ( .A(p_input[3614]), .Z(n4513) );
  XOR U4627 ( .A(n4915), .B(n4916), .Z(n4911) );
  AND U4628 ( .A(n4917), .B(n4918), .Z(n4916) );
  XNOR U4629 ( .A(p_input[3645]), .B(n4915), .Z(n4918) );
  XNOR U4630 ( .A(n4915), .B(n4522), .Z(n4917) );
  IV U4631 ( .A(p_input[3613]), .Z(n4522) );
  XOR U4632 ( .A(n4919), .B(n4920), .Z(n4915) );
  AND U4633 ( .A(n4921), .B(n4922), .Z(n4920) );
  XNOR U4634 ( .A(p_input[3644]), .B(n4919), .Z(n4922) );
  XNOR U4635 ( .A(n4919), .B(n4531), .Z(n4921) );
  IV U4636 ( .A(p_input[3612]), .Z(n4531) );
  XOR U4637 ( .A(n4923), .B(n4924), .Z(n4919) );
  AND U4638 ( .A(n4925), .B(n4926), .Z(n4924) );
  XNOR U4639 ( .A(p_input[3643]), .B(n4923), .Z(n4926) );
  XNOR U4640 ( .A(n4923), .B(n4540), .Z(n4925) );
  IV U4641 ( .A(p_input[3611]), .Z(n4540) );
  XOR U4642 ( .A(n4927), .B(n4928), .Z(n4923) );
  AND U4643 ( .A(n4929), .B(n4930), .Z(n4928) );
  XNOR U4644 ( .A(p_input[3642]), .B(n4927), .Z(n4930) );
  XNOR U4645 ( .A(n4927), .B(n4549), .Z(n4929) );
  IV U4646 ( .A(p_input[3610]), .Z(n4549) );
  XOR U4647 ( .A(n4931), .B(n4932), .Z(n4927) );
  AND U4648 ( .A(n4933), .B(n4934), .Z(n4932) );
  XNOR U4649 ( .A(p_input[3641]), .B(n4931), .Z(n4934) );
  XNOR U4650 ( .A(n4931), .B(n4558), .Z(n4933) );
  IV U4651 ( .A(p_input[3609]), .Z(n4558) );
  XOR U4652 ( .A(n4935), .B(n4936), .Z(n4931) );
  AND U4653 ( .A(n4937), .B(n4938), .Z(n4936) );
  XNOR U4654 ( .A(p_input[3640]), .B(n4935), .Z(n4938) );
  XNOR U4655 ( .A(n4935), .B(n4567), .Z(n4937) );
  IV U4656 ( .A(p_input[3608]), .Z(n4567) );
  XOR U4657 ( .A(n4939), .B(n4940), .Z(n4935) );
  AND U4658 ( .A(n4941), .B(n4942), .Z(n4940) );
  XNOR U4659 ( .A(p_input[3639]), .B(n4939), .Z(n4942) );
  XNOR U4660 ( .A(n4939), .B(n4576), .Z(n4941) );
  IV U4661 ( .A(p_input[3607]), .Z(n4576) );
  XOR U4662 ( .A(n4943), .B(n4944), .Z(n4939) );
  AND U4663 ( .A(n4945), .B(n4946), .Z(n4944) );
  XNOR U4664 ( .A(p_input[3638]), .B(n4943), .Z(n4946) );
  XNOR U4665 ( .A(n4943), .B(n4585), .Z(n4945) );
  IV U4666 ( .A(p_input[3606]), .Z(n4585) );
  XOR U4667 ( .A(n4947), .B(n4948), .Z(n4943) );
  AND U4668 ( .A(n4949), .B(n4950), .Z(n4948) );
  XNOR U4669 ( .A(p_input[3637]), .B(n4947), .Z(n4950) );
  XNOR U4670 ( .A(n4947), .B(n4594), .Z(n4949) );
  IV U4671 ( .A(p_input[3605]), .Z(n4594) );
  XOR U4672 ( .A(n4951), .B(n4952), .Z(n4947) );
  AND U4673 ( .A(n4953), .B(n4954), .Z(n4952) );
  XNOR U4674 ( .A(p_input[3636]), .B(n4951), .Z(n4954) );
  XNOR U4675 ( .A(n4951), .B(n4603), .Z(n4953) );
  IV U4676 ( .A(p_input[3604]), .Z(n4603) );
  XOR U4677 ( .A(n4955), .B(n4956), .Z(n4951) );
  AND U4678 ( .A(n4957), .B(n4958), .Z(n4956) );
  XNOR U4679 ( .A(p_input[3635]), .B(n4955), .Z(n4958) );
  XNOR U4680 ( .A(n4955), .B(n4612), .Z(n4957) );
  IV U4681 ( .A(p_input[3603]), .Z(n4612) );
  XOR U4682 ( .A(n4959), .B(n4960), .Z(n4955) );
  AND U4683 ( .A(n4961), .B(n4962), .Z(n4960) );
  XNOR U4684 ( .A(p_input[3634]), .B(n4959), .Z(n4962) );
  XNOR U4685 ( .A(n4959), .B(n4621), .Z(n4961) );
  IV U4686 ( .A(p_input[3602]), .Z(n4621) );
  XOR U4687 ( .A(n4963), .B(n4964), .Z(n4959) );
  AND U4688 ( .A(n4965), .B(n4966), .Z(n4964) );
  XNOR U4689 ( .A(p_input[3633]), .B(n4963), .Z(n4966) );
  XNOR U4690 ( .A(n4963), .B(n4630), .Z(n4965) );
  IV U4691 ( .A(p_input[3601]), .Z(n4630) );
  XOR U4692 ( .A(n4967), .B(n4968), .Z(n4963) );
  AND U4693 ( .A(n4969), .B(n4970), .Z(n4968) );
  XNOR U4694 ( .A(p_input[3632]), .B(n4967), .Z(n4970) );
  XNOR U4695 ( .A(n4967), .B(n4639), .Z(n4969) );
  IV U4696 ( .A(p_input[3600]), .Z(n4639) );
  XOR U4697 ( .A(n4971), .B(n4972), .Z(n4967) );
  AND U4698 ( .A(n4973), .B(n4974), .Z(n4972) );
  XNOR U4699 ( .A(p_input[3631]), .B(n4971), .Z(n4974) );
  XNOR U4700 ( .A(n4971), .B(n4648), .Z(n4973) );
  IV U4701 ( .A(p_input[3599]), .Z(n4648) );
  XOR U4702 ( .A(n4975), .B(n4976), .Z(n4971) );
  AND U4703 ( .A(n4977), .B(n4978), .Z(n4976) );
  XNOR U4704 ( .A(p_input[3630]), .B(n4975), .Z(n4978) );
  XNOR U4705 ( .A(n4975), .B(n4657), .Z(n4977) );
  IV U4706 ( .A(p_input[3598]), .Z(n4657) );
  XOR U4707 ( .A(n4979), .B(n4980), .Z(n4975) );
  AND U4708 ( .A(n4981), .B(n4982), .Z(n4980) );
  XNOR U4709 ( .A(p_input[3629]), .B(n4979), .Z(n4982) );
  XNOR U4710 ( .A(n4979), .B(n4666), .Z(n4981) );
  IV U4711 ( .A(p_input[3597]), .Z(n4666) );
  XOR U4712 ( .A(n4983), .B(n4984), .Z(n4979) );
  AND U4713 ( .A(n4985), .B(n4986), .Z(n4984) );
  XNOR U4714 ( .A(p_input[3628]), .B(n4983), .Z(n4986) );
  XNOR U4715 ( .A(n4983), .B(n4675), .Z(n4985) );
  IV U4716 ( .A(p_input[3596]), .Z(n4675) );
  XOR U4717 ( .A(n4987), .B(n4988), .Z(n4983) );
  AND U4718 ( .A(n4989), .B(n4990), .Z(n4988) );
  XNOR U4719 ( .A(p_input[3627]), .B(n4987), .Z(n4990) );
  XNOR U4720 ( .A(n4987), .B(n4684), .Z(n4989) );
  IV U4721 ( .A(p_input[3595]), .Z(n4684) );
  XOR U4722 ( .A(n4991), .B(n4992), .Z(n4987) );
  AND U4723 ( .A(n4993), .B(n4994), .Z(n4992) );
  XNOR U4724 ( .A(p_input[3626]), .B(n4991), .Z(n4994) );
  XNOR U4725 ( .A(n4991), .B(n4693), .Z(n4993) );
  IV U4726 ( .A(p_input[3594]), .Z(n4693) );
  XOR U4727 ( .A(n4995), .B(n4996), .Z(n4991) );
  AND U4728 ( .A(n4997), .B(n4998), .Z(n4996) );
  XNOR U4729 ( .A(p_input[3625]), .B(n4995), .Z(n4998) );
  XNOR U4730 ( .A(n4995), .B(n4702), .Z(n4997) );
  IV U4731 ( .A(p_input[3593]), .Z(n4702) );
  XOR U4732 ( .A(n4999), .B(n5000), .Z(n4995) );
  AND U4733 ( .A(n5001), .B(n5002), .Z(n5000) );
  XNOR U4734 ( .A(p_input[3624]), .B(n4999), .Z(n5002) );
  XNOR U4735 ( .A(n4999), .B(n4711), .Z(n5001) );
  IV U4736 ( .A(p_input[3592]), .Z(n4711) );
  XOR U4737 ( .A(n5003), .B(n5004), .Z(n4999) );
  AND U4738 ( .A(n5005), .B(n5006), .Z(n5004) );
  XNOR U4739 ( .A(p_input[3623]), .B(n5003), .Z(n5006) );
  XNOR U4740 ( .A(n5003), .B(n4720), .Z(n5005) );
  IV U4741 ( .A(p_input[3591]), .Z(n4720) );
  XOR U4742 ( .A(n5007), .B(n5008), .Z(n5003) );
  AND U4743 ( .A(n5009), .B(n5010), .Z(n5008) );
  XNOR U4744 ( .A(p_input[3622]), .B(n5007), .Z(n5010) );
  XNOR U4745 ( .A(n5007), .B(n4729), .Z(n5009) );
  IV U4746 ( .A(p_input[3590]), .Z(n4729) );
  XOR U4747 ( .A(n5011), .B(n5012), .Z(n5007) );
  AND U4748 ( .A(n5013), .B(n5014), .Z(n5012) );
  XNOR U4749 ( .A(p_input[3621]), .B(n5011), .Z(n5014) );
  XNOR U4750 ( .A(n5011), .B(n4738), .Z(n5013) );
  IV U4751 ( .A(p_input[3589]), .Z(n4738) );
  XOR U4752 ( .A(n5015), .B(n5016), .Z(n5011) );
  AND U4753 ( .A(n5017), .B(n5018), .Z(n5016) );
  XNOR U4754 ( .A(p_input[3620]), .B(n5015), .Z(n5018) );
  XNOR U4755 ( .A(n5015), .B(n4747), .Z(n5017) );
  IV U4756 ( .A(p_input[3588]), .Z(n4747) );
  XOR U4757 ( .A(n5019), .B(n5020), .Z(n5015) );
  AND U4758 ( .A(n5021), .B(n5022), .Z(n5020) );
  XNOR U4759 ( .A(p_input[3619]), .B(n5019), .Z(n5022) );
  XNOR U4760 ( .A(n5019), .B(n4756), .Z(n5021) );
  IV U4761 ( .A(p_input[3587]), .Z(n4756) );
  XOR U4762 ( .A(n5023), .B(n5024), .Z(n5019) );
  AND U4763 ( .A(n5025), .B(n5026), .Z(n5024) );
  XNOR U4764 ( .A(p_input[3618]), .B(n5023), .Z(n5026) );
  XNOR U4765 ( .A(n5023), .B(n4765), .Z(n5025) );
  IV U4766 ( .A(p_input[3586]), .Z(n4765) );
  XNOR U4767 ( .A(n5027), .B(n5028), .Z(n5023) );
  AND U4768 ( .A(n5029), .B(n5030), .Z(n5028) );
  XOR U4769 ( .A(p_input[3617]), .B(n5027), .Z(n5030) );
  XNOR U4770 ( .A(p_input[3585]), .B(n5027), .Z(n5029) );
  AND U4771 ( .A(p_input[3616]), .B(n5031), .Z(n5027) );
  IV U4772 ( .A(p_input[3584]), .Z(n5031) );
  XOR U4773 ( .A(n5032), .B(n5033), .Z(n1388) );
  AND U4774 ( .A(n576), .B(n5034), .Z(n5033) );
  XNOR U4775 ( .A(n5035), .B(n5032), .Z(n5034) );
  XOR U4776 ( .A(n5036), .B(n5037), .Z(n576) );
  AND U4777 ( .A(n5038), .B(n5039), .Z(n5037) );
  XOR U4778 ( .A(n5036), .B(n1403), .Z(n5039) );
  XOR U4779 ( .A(n5040), .B(n5041), .Z(n1403) );
  AND U4780 ( .A(n494), .B(n5042), .Z(n5041) );
  XOR U4781 ( .A(n5043), .B(n5040), .Z(n5042) );
  XNOR U4782 ( .A(n1400), .B(n5036), .Z(n5038) );
  XOR U4783 ( .A(n5044), .B(n5045), .Z(n1400) );
  AND U4784 ( .A(n491), .B(n5046), .Z(n5045) );
  XOR U4785 ( .A(n5047), .B(n5044), .Z(n5046) );
  XOR U4786 ( .A(n5048), .B(n5049), .Z(n5036) );
  AND U4787 ( .A(n5050), .B(n5051), .Z(n5049) );
  XOR U4788 ( .A(n5048), .B(n1415), .Z(n5051) );
  XOR U4789 ( .A(n5052), .B(n5053), .Z(n1415) );
  AND U4790 ( .A(n494), .B(n5054), .Z(n5053) );
  XOR U4791 ( .A(n5055), .B(n5052), .Z(n5054) );
  XNOR U4792 ( .A(n1412), .B(n5048), .Z(n5050) );
  XOR U4793 ( .A(n5056), .B(n5057), .Z(n1412) );
  AND U4794 ( .A(n491), .B(n5058), .Z(n5057) );
  XOR U4795 ( .A(n5059), .B(n5056), .Z(n5058) );
  XOR U4796 ( .A(n5060), .B(n5061), .Z(n5048) );
  AND U4797 ( .A(n5062), .B(n5063), .Z(n5061) );
  XOR U4798 ( .A(n5060), .B(n1427), .Z(n5063) );
  XOR U4799 ( .A(n5064), .B(n5065), .Z(n1427) );
  AND U4800 ( .A(n494), .B(n5066), .Z(n5065) );
  XOR U4801 ( .A(n5067), .B(n5064), .Z(n5066) );
  XNOR U4802 ( .A(n1424), .B(n5060), .Z(n5062) );
  XOR U4803 ( .A(n5068), .B(n5069), .Z(n1424) );
  AND U4804 ( .A(n491), .B(n5070), .Z(n5069) );
  XOR U4805 ( .A(n5071), .B(n5068), .Z(n5070) );
  XOR U4806 ( .A(n5072), .B(n5073), .Z(n5060) );
  AND U4807 ( .A(n5074), .B(n5075), .Z(n5073) );
  XOR U4808 ( .A(n5072), .B(n1439), .Z(n5075) );
  XOR U4809 ( .A(n5076), .B(n5077), .Z(n1439) );
  AND U4810 ( .A(n494), .B(n5078), .Z(n5077) );
  XOR U4811 ( .A(n5079), .B(n5076), .Z(n5078) );
  XNOR U4812 ( .A(n1436), .B(n5072), .Z(n5074) );
  XOR U4813 ( .A(n5080), .B(n5081), .Z(n1436) );
  AND U4814 ( .A(n491), .B(n5082), .Z(n5081) );
  XOR U4815 ( .A(n5083), .B(n5080), .Z(n5082) );
  XOR U4816 ( .A(n5084), .B(n5085), .Z(n5072) );
  AND U4817 ( .A(n5086), .B(n5087), .Z(n5085) );
  XOR U4818 ( .A(n5084), .B(n1451), .Z(n5087) );
  XOR U4819 ( .A(n5088), .B(n5089), .Z(n1451) );
  AND U4820 ( .A(n494), .B(n5090), .Z(n5089) );
  XOR U4821 ( .A(n5091), .B(n5088), .Z(n5090) );
  XNOR U4822 ( .A(n1448), .B(n5084), .Z(n5086) );
  XOR U4823 ( .A(n5092), .B(n5093), .Z(n1448) );
  AND U4824 ( .A(n491), .B(n5094), .Z(n5093) );
  XOR U4825 ( .A(n5095), .B(n5092), .Z(n5094) );
  XOR U4826 ( .A(n5096), .B(n5097), .Z(n5084) );
  AND U4827 ( .A(n5098), .B(n5099), .Z(n5097) );
  XOR U4828 ( .A(n5096), .B(n1463), .Z(n5099) );
  XOR U4829 ( .A(n5100), .B(n5101), .Z(n1463) );
  AND U4830 ( .A(n494), .B(n5102), .Z(n5101) );
  XOR U4831 ( .A(n5103), .B(n5100), .Z(n5102) );
  XNOR U4832 ( .A(n1460), .B(n5096), .Z(n5098) );
  XOR U4833 ( .A(n5104), .B(n5105), .Z(n1460) );
  AND U4834 ( .A(n491), .B(n5106), .Z(n5105) );
  XOR U4835 ( .A(n5107), .B(n5104), .Z(n5106) );
  XOR U4836 ( .A(n5108), .B(n5109), .Z(n5096) );
  AND U4837 ( .A(n5110), .B(n5111), .Z(n5109) );
  XOR U4838 ( .A(n5108), .B(n1475), .Z(n5111) );
  XOR U4839 ( .A(n5112), .B(n5113), .Z(n1475) );
  AND U4840 ( .A(n494), .B(n5114), .Z(n5113) );
  XOR U4841 ( .A(n5115), .B(n5112), .Z(n5114) );
  XNOR U4842 ( .A(n1472), .B(n5108), .Z(n5110) );
  XOR U4843 ( .A(n5116), .B(n5117), .Z(n1472) );
  AND U4844 ( .A(n491), .B(n5118), .Z(n5117) );
  XOR U4845 ( .A(n5119), .B(n5116), .Z(n5118) );
  XOR U4846 ( .A(n5120), .B(n5121), .Z(n5108) );
  AND U4847 ( .A(n5122), .B(n5123), .Z(n5121) );
  XOR U4848 ( .A(n5120), .B(n1487), .Z(n5123) );
  XOR U4849 ( .A(n5124), .B(n5125), .Z(n1487) );
  AND U4850 ( .A(n494), .B(n5126), .Z(n5125) );
  XOR U4851 ( .A(n5127), .B(n5124), .Z(n5126) );
  XNOR U4852 ( .A(n1484), .B(n5120), .Z(n5122) );
  XOR U4853 ( .A(n5128), .B(n5129), .Z(n1484) );
  AND U4854 ( .A(n491), .B(n5130), .Z(n5129) );
  XOR U4855 ( .A(n5131), .B(n5128), .Z(n5130) );
  XOR U4856 ( .A(n5132), .B(n5133), .Z(n5120) );
  AND U4857 ( .A(n5134), .B(n5135), .Z(n5133) );
  XOR U4858 ( .A(n5132), .B(n1499), .Z(n5135) );
  XOR U4859 ( .A(n5136), .B(n5137), .Z(n1499) );
  AND U4860 ( .A(n494), .B(n5138), .Z(n5137) );
  XOR U4861 ( .A(n5139), .B(n5136), .Z(n5138) );
  XNOR U4862 ( .A(n1496), .B(n5132), .Z(n5134) );
  XOR U4863 ( .A(n5140), .B(n5141), .Z(n1496) );
  AND U4864 ( .A(n491), .B(n5142), .Z(n5141) );
  XOR U4865 ( .A(n5143), .B(n5140), .Z(n5142) );
  XOR U4866 ( .A(n5144), .B(n5145), .Z(n5132) );
  AND U4867 ( .A(n5146), .B(n5147), .Z(n5145) );
  XOR U4868 ( .A(n5144), .B(n1511), .Z(n5147) );
  XOR U4869 ( .A(n5148), .B(n5149), .Z(n1511) );
  AND U4870 ( .A(n494), .B(n5150), .Z(n5149) );
  XOR U4871 ( .A(n5151), .B(n5148), .Z(n5150) );
  XNOR U4872 ( .A(n1508), .B(n5144), .Z(n5146) );
  XOR U4873 ( .A(n5152), .B(n5153), .Z(n1508) );
  AND U4874 ( .A(n491), .B(n5154), .Z(n5153) );
  XOR U4875 ( .A(n5155), .B(n5152), .Z(n5154) );
  XOR U4876 ( .A(n5156), .B(n5157), .Z(n5144) );
  AND U4877 ( .A(n5158), .B(n5159), .Z(n5157) );
  XOR U4878 ( .A(n5156), .B(n1523), .Z(n5159) );
  XOR U4879 ( .A(n5160), .B(n5161), .Z(n1523) );
  AND U4880 ( .A(n494), .B(n5162), .Z(n5161) );
  XOR U4881 ( .A(n5163), .B(n5160), .Z(n5162) );
  XNOR U4882 ( .A(n1520), .B(n5156), .Z(n5158) );
  XOR U4883 ( .A(n5164), .B(n5165), .Z(n1520) );
  AND U4884 ( .A(n491), .B(n5166), .Z(n5165) );
  XOR U4885 ( .A(n5167), .B(n5164), .Z(n5166) );
  XOR U4886 ( .A(n5168), .B(n5169), .Z(n5156) );
  AND U4887 ( .A(n5170), .B(n5171), .Z(n5169) );
  XOR U4888 ( .A(n5168), .B(n1535), .Z(n5171) );
  XOR U4889 ( .A(n5172), .B(n5173), .Z(n1535) );
  AND U4890 ( .A(n494), .B(n5174), .Z(n5173) );
  XOR U4891 ( .A(n5175), .B(n5172), .Z(n5174) );
  XNOR U4892 ( .A(n1532), .B(n5168), .Z(n5170) );
  XOR U4893 ( .A(n5176), .B(n5177), .Z(n1532) );
  AND U4894 ( .A(n491), .B(n5178), .Z(n5177) );
  XOR U4895 ( .A(n5179), .B(n5176), .Z(n5178) );
  XOR U4896 ( .A(n5180), .B(n5181), .Z(n5168) );
  AND U4897 ( .A(n5182), .B(n5183), .Z(n5181) );
  XOR U4898 ( .A(n5180), .B(n1547), .Z(n5183) );
  XOR U4899 ( .A(n5184), .B(n5185), .Z(n1547) );
  AND U4900 ( .A(n494), .B(n5186), .Z(n5185) );
  XOR U4901 ( .A(n5187), .B(n5184), .Z(n5186) );
  XNOR U4902 ( .A(n1544), .B(n5180), .Z(n5182) );
  XOR U4903 ( .A(n5188), .B(n5189), .Z(n1544) );
  AND U4904 ( .A(n491), .B(n5190), .Z(n5189) );
  XOR U4905 ( .A(n5191), .B(n5188), .Z(n5190) );
  XOR U4906 ( .A(n5192), .B(n5193), .Z(n5180) );
  AND U4907 ( .A(n5194), .B(n5195), .Z(n5193) );
  XOR U4908 ( .A(n5192), .B(n1559), .Z(n5195) );
  XOR U4909 ( .A(n5196), .B(n5197), .Z(n1559) );
  AND U4910 ( .A(n494), .B(n5198), .Z(n5197) );
  XOR U4911 ( .A(n5199), .B(n5196), .Z(n5198) );
  XNOR U4912 ( .A(n1556), .B(n5192), .Z(n5194) );
  XOR U4913 ( .A(n5200), .B(n5201), .Z(n1556) );
  AND U4914 ( .A(n491), .B(n5202), .Z(n5201) );
  XOR U4915 ( .A(n5203), .B(n5200), .Z(n5202) );
  XOR U4916 ( .A(n5204), .B(n5205), .Z(n5192) );
  AND U4917 ( .A(n5206), .B(n5207), .Z(n5205) );
  XOR U4918 ( .A(n5204), .B(n1571), .Z(n5207) );
  XOR U4919 ( .A(n5208), .B(n5209), .Z(n1571) );
  AND U4920 ( .A(n494), .B(n5210), .Z(n5209) );
  XOR U4921 ( .A(n5211), .B(n5208), .Z(n5210) );
  XNOR U4922 ( .A(n1568), .B(n5204), .Z(n5206) );
  XOR U4923 ( .A(n5212), .B(n5213), .Z(n1568) );
  AND U4924 ( .A(n491), .B(n5214), .Z(n5213) );
  XOR U4925 ( .A(n5215), .B(n5212), .Z(n5214) );
  XOR U4926 ( .A(n5216), .B(n5217), .Z(n5204) );
  AND U4927 ( .A(n5218), .B(n5219), .Z(n5217) );
  XOR U4928 ( .A(n5216), .B(n1583), .Z(n5219) );
  XOR U4929 ( .A(n5220), .B(n5221), .Z(n1583) );
  AND U4930 ( .A(n494), .B(n5222), .Z(n5221) );
  XOR U4931 ( .A(n5223), .B(n5220), .Z(n5222) );
  XNOR U4932 ( .A(n1580), .B(n5216), .Z(n5218) );
  XOR U4933 ( .A(n5224), .B(n5225), .Z(n1580) );
  AND U4934 ( .A(n491), .B(n5226), .Z(n5225) );
  XOR U4935 ( .A(n5227), .B(n5224), .Z(n5226) );
  XOR U4936 ( .A(n5228), .B(n5229), .Z(n5216) );
  AND U4937 ( .A(n5230), .B(n5231), .Z(n5229) );
  XOR U4938 ( .A(n5228), .B(n1595), .Z(n5231) );
  XOR U4939 ( .A(n5232), .B(n5233), .Z(n1595) );
  AND U4940 ( .A(n494), .B(n5234), .Z(n5233) );
  XOR U4941 ( .A(n5235), .B(n5232), .Z(n5234) );
  XNOR U4942 ( .A(n1592), .B(n5228), .Z(n5230) );
  XOR U4943 ( .A(n5236), .B(n5237), .Z(n1592) );
  AND U4944 ( .A(n491), .B(n5238), .Z(n5237) );
  XOR U4945 ( .A(n5239), .B(n5236), .Z(n5238) );
  XOR U4946 ( .A(n5240), .B(n5241), .Z(n5228) );
  AND U4947 ( .A(n5242), .B(n5243), .Z(n5241) );
  XOR U4948 ( .A(n5240), .B(n1607), .Z(n5243) );
  XOR U4949 ( .A(n5244), .B(n5245), .Z(n1607) );
  AND U4950 ( .A(n494), .B(n5246), .Z(n5245) );
  XOR U4951 ( .A(n5247), .B(n5244), .Z(n5246) );
  XNOR U4952 ( .A(n1604), .B(n5240), .Z(n5242) );
  XOR U4953 ( .A(n5248), .B(n5249), .Z(n1604) );
  AND U4954 ( .A(n491), .B(n5250), .Z(n5249) );
  XOR U4955 ( .A(n5251), .B(n5248), .Z(n5250) );
  XOR U4956 ( .A(n5252), .B(n5253), .Z(n5240) );
  AND U4957 ( .A(n5254), .B(n5255), .Z(n5253) );
  XOR U4958 ( .A(n5252), .B(n1619), .Z(n5255) );
  XOR U4959 ( .A(n5256), .B(n5257), .Z(n1619) );
  AND U4960 ( .A(n494), .B(n5258), .Z(n5257) );
  XOR U4961 ( .A(n5259), .B(n5256), .Z(n5258) );
  XNOR U4962 ( .A(n1616), .B(n5252), .Z(n5254) );
  XOR U4963 ( .A(n5260), .B(n5261), .Z(n1616) );
  AND U4964 ( .A(n491), .B(n5262), .Z(n5261) );
  XOR U4965 ( .A(n5263), .B(n5260), .Z(n5262) );
  XOR U4966 ( .A(n5264), .B(n5265), .Z(n5252) );
  AND U4967 ( .A(n5266), .B(n5267), .Z(n5265) );
  XOR U4968 ( .A(n5264), .B(n1631), .Z(n5267) );
  XOR U4969 ( .A(n5268), .B(n5269), .Z(n1631) );
  AND U4970 ( .A(n494), .B(n5270), .Z(n5269) );
  XOR U4971 ( .A(n5271), .B(n5268), .Z(n5270) );
  XNOR U4972 ( .A(n1628), .B(n5264), .Z(n5266) );
  XOR U4973 ( .A(n5272), .B(n5273), .Z(n1628) );
  AND U4974 ( .A(n491), .B(n5274), .Z(n5273) );
  XOR U4975 ( .A(n5275), .B(n5272), .Z(n5274) );
  XOR U4976 ( .A(n5276), .B(n5277), .Z(n5264) );
  AND U4977 ( .A(n5278), .B(n5279), .Z(n5277) );
  XOR U4978 ( .A(n5276), .B(n1643), .Z(n5279) );
  XOR U4979 ( .A(n5280), .B(n5281), .Z(n1643) );
  AND U4980 ( .A(n494), .B(n5282), .Z(n5281) );
  XOR U4981 ( .A(n5283), .B(n5280), .Z(n5282) );
  XNOR U4982 ( .A(n1640), .B(n5276), .Z(n5278) );
  XOR U4983 ( .A(n5284), .B(n5285), .Z(n1640) );
  AND U4984 ( .A(n491), .B(n5286), .Z(n5285) );
  XOR U4985 ( .A(n5287), .B(n5284), .Z(n5286) );
  XOR U4986 ( .A(n5288), .B(n5289), .Z(n5276) );
  AND U4987 ( .A(n5290), .B(n5291), .Z(n5289) );
  XOR U4988 ( .A(n5288), .B(n1655), .Z(n5291) );
  XOR U4989 ( .A(n5292), .B(n5293), .Z(n1655) );
  AND U4990 ( .A(n494), .B(n5294), .Z(n5293) );
  XOR U4991 ( .A(n5295), .B(n5292), .Z(n5294) );
  XNOR U4992 ( .A(n1652), .B(n5288), .Z(n5290) );
  XOR U4993 ( .A(n5296), .B(n5297), .Z(n1652) );
  AND U4994 ( .A(n491), .B(n5298), .Z(n5297) );
  XOR U4995 ( .A(n5299), .B(n5296), .Z(n5298) );
  XOR U4996 ( .A(n5300), .B(n5301), .Z(n5288) );
  AND U4997 ( .A(n5302), .B(n5303), .Z(n5301) );
  XOR U4998 ( .A(n5300), .B(n1667), .Z(n5303) );
  XOR U4999 ( .A(n5304), .B(n5305), .Z(n1667) );
  AND U5000 ( .A(n494), .B(n5306), .Z(n5305) );
  XOR U5001 ( .A(n5307), .B(n5304), .Z(n5306) );
  XNOR U5002 ( .A(n1664), .B(n5300), .Z(n5302) );
  XOR U5003 ( .A(n5308), .B(n5309), .Z(n1664) );
  AND U5004 ( .A(n491), .B(n5310), .Z(n5309) );
  XOR U5005 ( .A(n5311), .B(n5308), .Z(n5310) );
  XOR U5006 ( .A(n5312), .B(n5313), .Z(n5300) );
  AND U5007 ( .A(n5314), .B(n5315), .Z(n5313) );
  XOR U5008 ( .A(n5312), .B(n1679), .Z(n5315) );
  XOR U5009 ( .A(n5316), .B(n5317), .Z(n1679) );
  AND U5010 ( .A(n494), .B(n5318), .Z(n5317) );
  XOR U5011 ( .A(n5319), .B(n5316), .Z(n5318) );
  XNOR U5012 ( .A(n1676), .B(n5312), .Z(n5314) );
  XOR U5013 ( .A(n5320), .B(n5321), .Z(n1676) );
  AND U5014 ( .A(n491), .B(n5322), .Z(n5321) );
  XOR U5015 ( .A(n5323), .B(n5320), .Z(n5322) );
  XOR U5016 ( .A(n5324), .B(n5325), .Z(n5312) );
  AND U5017 ( .A(n5326), .B(n5327), .Z(n5325) );
  XOR U5018 ( .A(n5324), .B(n1691), .Z(n5327) );
  XOR U5019 ( .A(n5328), .B(n5329), .Z(n1691) );
  AND U5020 ( .A(n494), .B(n5330), .Z(n5329) );
  XOR U5021 ( .A(n5331), .B(n5328), .Z(n5330) );
  XNOR U5022 ( .A(n1688), .B(n5324), .Z(n5326) );
  XOR U5023 ( .A(n5332), .B(n5333), .Z(n1688) );
  AND U5024 ( .A(n491), .B(n5334), .Z(n5333) );
  XOR U5025 ( .A(n5335), .B(n5332), .Z(n5334) );
  XOR U5026 ( .A(n5336), .B(n5337), .Z(n5324) );
  AND U5027 ( .A(n5338), .B(n5339), .Z(n5337) );
  XOR U5028 ( .A(n5336), .B(n1703), .Z(n5339) );
  XOR U5029 ( .A(n5340), .B(n5341), .Z(n1703) );
  AND U5030 ( .A(n494), .B(n5342), .Z(n5341) );
  XOR U5031 ( .A(n5343), .B(n5340), .Z(n5342) );
  XNOR U5032 ( .A(n1700), .B(n5336), .Z(n5338) );
  XOR U5033 ( .A(n5344), .B(n5345), .Z(n1700) );
  AND U5034 ( .A(n491), .B(n5346), .Z(n5345) );
  XOR U5035 ( .A(n5347), .B(n5344), .Z(n5346) );
  XOR U5036 ( .A(n5348), .B(n5349), .Z(n5336) );
  AND U5037 ( .A(n5350), .B(n5351), .Z(n5349) );
  XOR U5038 ( .A(n5348), .B(n1715), .Z(n5351) );
  XOR U5039 ( .A(n5352), .B(n5353), .Z(n1715) );
  AND U5040 ( .A(n494), .B(n5354), .Z(n5353) );
  XOR U5041 ( .A(n5355), .B(n5352), .Z(n5354) );
  XNOR U5042 ( .A(n1712), .B(n5348), .Z(n5350) );
  XOR U5043 ( .A(n5356), .B(n5357), .Z(n1712) );
  AND U5044 ( .A(n491), .B(n5358), .Z(n5357) );
  XOR U5045 ( .A(n5359), .B(n5356), .Z(n5358) );
  XOR U5046 ( .A(n5360), .B(n5361), .Z(n5348) );
  AND U5047 ( .A(n5362), .B(n5363), .Z(n5361) );
  XOR U5048 ( .A(n5360), .B(n1727), .Z(n5363) );
  XOR U5049 ( .A(n5364), .B(n5365), .Z(n1727) );
  AND U5050 ( .A(n494), .B(n5366), .Z(n5365) );
  XOR U5051 ( .A(n5367), .B(n5364), .Z(n5366) );
  XNOR U5052 ( .A(n1724), .B(n5360), .Z(n5362) );
  XOR U5053 ( .A(n5368), .B(n5369), .Z(n1724) );
  AND U5054 ( .A(n491), .B(n5370), .Z(n5369) );
  XOR U5055 ( .A(n5371), .B(n5368), .Z(n5370) );
  XOR U5056 ( .A(n5372), .B(n5373), .Z(n5360) );
  AND U5057 ( .A(n5374), .B(n5375), .Z(n5373) );
  XOR U5058 ( .A(n5372), .B(n1739), .Z(n5375) );
  XOR U5059 ( .A(n5376), .B(n5377), .Z(n1739) );
  AND U5060 ( .A(n494), .B(n5378), .Z(n5377) );
  XOR U5061 ( .A(n5379), .B(n5376), .Z(n5378) );
  XNOR U5062 ( .A(n1736), .B(n5372), .Z(n5374) );
  XOR U5063 ( .A(n5380), .B(n5381), .Z(n1736) );
  AND U5064 ( .A(n491), .B(n5382), .Z(n5381) );
  XOR U5065 ( .A(n5383), .B(n5380), .Z(n5382) );
  XOR U5066 ( .A(n5384), .B(n5385), .Z(n5372) );
  AND U5067 ( .A(n5386), .B(n5387), .Z(n5385) );
  XOR U5068 ( .A(n1751), .B(n5384), .Z(n5387) );
  XOR U5069 ( .A(n5388), .B(n5389), .Z(n1751) );
  AND U5070 ( .A(n494), .B(n5390), .Z(n5389) );
  XOR U5071 ( .A(n5388), .B(n5391), .Z(n5390) );
  XNOR U5072 ( .A(n5384), .B(n1748), .Z(n5386) );
  XOR U5073 ( .A(n5392), .B(n5393), .Z(n1748) );
  AND U5074 ( .A(n491), .B(n5394), .Z(n5393) );
  XOR U5075 ( .A(n5392), .B(n5395), .Z(n5394) );
  XOR U5076 ( .A(n5396), .B(n5397), .Z(n5384) );
  AND U5077 ( .A(n5398), .B(n5399), .Z(n5397) );
  XNOR U5078 ( .A(n5400), .B(n1764), .Z(n5399) );
  XOR U5079 ( .A(n5401), .B(n5402), .Z(n1764) );
  AND U5080 ( .A(n494), .B(n5403), .Z(n5402) );
  XOR U5081 ( .A(n5404), .B(n5401), .Z(n5403) );
  XNOR U5082 ( .A(n1761), .B(n5396), .Z(n5398) );
  XOR U5083 ( .A(n5405), .B(n5406), .Z(n1761) );
  AND U5084 ( .A(n491), .B(n5407), .Z(n5406) );
  XOR U5085 ( .A(n5408), .B(n5405), .Z(n5407) );
  IV U5086 ( .A(n5400), .Z(n5396) );
  AND U5087 ( .A(n5032), .B(n5035), .Z(n5400) );
  XNOR U5088 ( .A(n5409), .B(n5410), .Z(n5035) );
  AND U5089 ( .A(n494), .B(n5411), .Z(n5410) );
  XNOR U5090 ( .A(n5412), .B(n5409), .Z(n5411) );
  XOR U5091 ( .A(n5413), .B(n5414), .Z(n494) );
  AND U5092 ( .A(n5415), .B(n5416), .Z(n5414) );
  XOR U5093 ( .A(n5413), .B(n5043), .Z(n5416) );
  XNOR U5094 ( .A(n5417), .B(n5418), .Z(n5043) );
  AND U5095 ( .A(n5419), .B(n318), .Z(n5418) );
  AND U5096 ( .A(n5417), .B(n5420), .Z(n5419) );
  XNOR U5097 ( .A(n5040), .B(n5413), .Z(n5415) );
  XOR U5098 ( .A(n5421), .B(n5422), .Z(n5040) );
  AND U5099 ( .A(n5423), .B(n316), .Z(n5422) );
  NOR U5100 ( .A(n5421), .B(n5424), .Z(n5423) );
  XOR U5101 ( .A(n5425), .B(n5426), .Z(n5413) );
  AND U5102 ( .A(n5427), .B(n5428), .Z(n5426) );
  XOR U5103 ( .A(n5425), .B(n5055), .Z(n5428) );
  XOR U5104 ( .A(n5429), .B(n5430), .Z(n5055) );
  AND U5105 ( .A(n318), .B(n5431), .Z(n5430) );
  XOR U5106 ( .A(n5432), .B(n5429), .Z(n5431) );
  XNOR U5107 ( .A(n5052), .B(n5425), .Z(n5427) );
  XOR U5108 ( .A(n5433), .B(n5434), .Z(n5052) );
  AND U5109 ( .A(n316), .B(n5435), .Z(n5434) );
  XOR U5110 ( .A(n5436), .B(n5433), .Z(n5435) );
  XOR U5111 ( .A(n5437), .B(n5438), .Z(n5425) );
  AND U5112 ( .A(n5439), .B(n5440), .Z(n5438) );
  XOR U5113 ( .A(n5437), .B(n5067), .Z(n5440) );
  XOR U5114 ( .A(n5441), .B(n5442), .Z(n5067) );
  AND U5115 ( .A(n318), .B(n5443), .Z(n5442) );
  XOR U5116 ( .A(n5444), .B(n5441), .Z(n5443) );
  XNOR U5117 ( .A(n5064), .B(n5437), .Z(n5439) );
  XOR U5118 ( .A(n5445), .B(n5446), .Z(n5064) );
  AND U5119 ( .A(n316), .B(n5447), .Z(n5446) );
  XOR U5120 ( .A(n5448), .B(n5445), .Z(n5447) );
  XOR U5121 ( .A(n5449), .B(n5450), .Z(n5437) );
  AND U5122 ( .A(n5451), .B(n5452), .Z(n5450) );
  XOR U5123 ( .A(n5449), .B(n5079), .Z(n5452) );
  XOR U5124 ( .A(n5453), .B(n5454), .Z(n5079) );
  AND U5125 ( .A(n318), .B(n5455), .Z(n5454) );
  XOR U5126 ( .A(n5456), .B(n5453), .Z(n5455) );
  XNOR U5127 ( .A(n5076), .B(n5449), .Z(n5451) );
  XOR U5128 ( .A(n5457), .B(n5458), .Z(n5076) );
  AND U5129 ( .A(n316), .B(n5459), .Z(n5458) );
  XOR U5130 ( .A(n5460), .B(n5457), .Z(n5459) );
  XOR U5131 ( .A(n5461), .B(n5462), .Z(n5449) );
  AND U5132 ( .A(n5463), .B(n5464), .Z(n5462) );
  XOR U5133 ( .A(n5461), .B(n5091), .Z(n5464) );
  XOR U5134 ( .A(n5465), .B(n5466), .Z(n5091) );
  AND U5135 ( .A(n318), .B(n5467), .Z(n5466) );
  XOR U5136 ( .A(n5468), .B(n5465), .Z(n5467) );
  XNOR U5137 ( .A(n5088), .B(n5461), .Z(n5463) );
  XOR U5138 ( .A(n5469), .B(n5470), .Z(n5088) );
  AND U5139 ( .A(n316), .B(n5471), .Z(n5470) );
  XOR U5140 ( .A(n5472), .B(n5469), .Z(n5471) );
  XOR U5141 ( .A(n5473), .B(n5474), .Z(n5461) );
  AND U5142 ( .A(n5475), .B(n5476), .Z(n5474) );
  XOR U5143 ( .A(n5473), .B(n5103), .Z(n5476) );
  XOR U5144 ( .A(n5477), .B(n5478), .Z(n5103) );
  AND U5145 ( .A(n318), .B(n5479), .Z(n5478) );
  XOR U5146 ( .A(n5480), .B(n5477), .Z(n5479) );
  XNOR U5147 ( .A(n5100), .B(n5473), .Z(n5475) );
  XOR U5148 ( .A(n5481), .B(n5482), .Z(n5100) );
  AND U5149 ( .A(n316), .B(n5483), .Z(n5482) );
  XOR U5150 ( .A(n5484), .B(n5481), .Z(n5483) );
  XOR U5151 ( .A(n5485), .B(n5486), .Z(n5473) );
  AND U5152 ( .A(n5487), .B(n5488), .Z(n5486) );
  XOR U5153 ( .A(n5485), .B(n5115), .Z(n5488) );
  XOR U5154 ( .A(n5489), .B(n5490), .Z(n5115) );
  AND U5155 ( .A(n318), .B(n5491), .Z(n5490) );
  XOR U5156 ( .A(n5492), .B(n5489), .Z(n5491) );
  XNOR U5157 ( .A(n5112), .B(n5485), .Z(n5487) );
  XOR U5158 ( .A(n5493), .B(n5494), .Z(n5112) );
  AND U5159 ( .A(n316), .B(n5495), .Z(n5494) );
  XOR U5160 ( .A(n5496), .B(n5493), .Z(n5495) );
  XOR U5161 ( .A(n5497), .B(n5498), .Z(n5485) );
  AND U5162 ( .A(n5499), .B(n5500), .Z(n5498) );
  XOR U5163 ( .A(n5497), .B(n5127), .Z(n5500) );
  XOR U5164 ( .A(n5501), .B(n5502), .Z(n5127) );
  AND U5165 ( .A(n318), .B(n5503), .Z(n5502) );
  XOR U5166 ( .A(n5504), .B(n5501), .Z(n5503) );
  XNOR U5167 ( .A(n5124), .B(n5497), .Z(n5499) );
  XOR U5168 ( .A(n5505), .B(n5506), .Z(n5124) );
  AND U5169 ( .A(n316), .B(n5507), .Z(n5506) );
  XOR U5170 ( .A(n5508), .B(n5505), .Z(n5507) );
  XOR U5171 ( .A(n5509), .B(n5510), .Z(n5497) );
  AND U5172 ( .A(n5511), .B(n5512), .Z(n5510) );
  XOR U5173 ( .A(n5509), .B(n5139), .Z(n5512) );
  XOR U5174 ( .A(n5513), .B(n5514), .Z(n5139) );
  AND U5175 ( .A(n318), .B(n5515), .Z(n5514) );
  XOR U5176 ( .A(n5516), .B(n5513), .Z(n5515) );
  XNOR U5177 ( .A(n5136), .B(n5509), .Z(n5511) );
  XOR U5178 ( .A(n5517), .B(n5518), .Z(n5136) );
  AND U5179 ( .A(n316), .B(n5519), .Z(n5518) );
  XOR U5180 ( .A(n5520), .B(n5517), .Z(n5519) );
  XOR U5181 ( .A(n5521), .B(n5522), .Z(n5509) );
  AND U5182 ( .A(n5523), .B(n5524), .Z(n5522) );
  XOR U5183 ( .A(n5521), .B(n5151), .Z(n5524) );
  XOR U5184 ( .A(n5525), .B(n5526), .Z(n5151) );
  AND U5185 ( .A(n318), .B(n5527), .Z(n5526) );
  XOR U5186 ( .A(n5528), .B(n5525), .Z(n5527) );
  XNOR U5187 ( .A(n5148), .B(n5521), .Z(n5523) );
  XOR U5188 ( .A(n5529), .B(n5530), .Z(n5148) );
  AND U5189 ( .A(n316), .B(n5531), .Z(n5530) );
  XOR U5190 ( .A(n5532), .B(n5529), .Z(n5531) );
  XOR U5191 ( .A(n5533), .B(n5534), .Z(n5521) );
  AND U5192 ( .A(n5535), .B(n5536), .Z(n5534) );
  XOR U5193 ( .A(n5533), .B(n5163), .Z(n5536) );
  XOR U5194 ( .A(n5537), .B(n5538), .Z(n5163) );
  AND U5195 ( .A(n318), .B(n5539), .Z(n5538) );
  XOR U5196 ( .A(n5540), .B(n5537), .Z(n5539) );
  XNOR U5197 ( .A(n5160), .B(n5533), .Z(n5535) );
  XOR U5198 ( .A(n5541), .B(n5542), .Z(n5160) );
  AND U5199 ( .A(n316), .B(n5543), .Z(n5542) );
  XOR U5200 ( .A(n5544), .B(n5541), .Z(n5543) );
  XOR U5201 ( .A(n5545), .B(n5546), .Z(n5533) );
  AND U5202 ( .A(n5547), .B(n5548), .Z(n5546) );
  XOR U5203 ( .A(n5545), .B(n5175), .Z(n5548) );
  XOR U5204 ( .A(n5549), .B(n5550), .Z(n5175) );
  AND U5205 ( .A(n318), .B(n5551), .Z(n5550) );
  XOR U5206 ( .A(n5552), .B(n5549), .Z(n5551) );
  XNOR U5207 ( .A(n5172), .B(n5545), .Z(n5547) );
  XOR U5208 ( .A(n5553), .B(n5554), .Z(n5172) );
  AND U5209 ( .A(n316), .B(n5555), .Z(n5554) );
  XOR U5210 ( .A(n5556), .B(n5553), .Z(n5555) );
  XOR U5211 ( .A(n5557), .B(n5558), .Z(n5545) );
  AND U5212 ( .A(n5559), .B(n5560), .Z(n5558) );
  XOR U5213 ( .A(n5557), .B(n5187), .Z(n5560) );
  XOR U5214 ( .A(n5561), .B(n5562), .Z(n5187) );
  AND U5215 ( .A(n318), .B(n5563), .Z(n5562) );
  XOR U5216 ( .A(n5564), .B(n5561), .Z(n5563) );
  XNOR U5217 ( .A(n5184), .B(n5557), .Z(n5559) );
  XOR U5218 ( .A(n5565), .B(n5566), .Z(n5184) );
  AND U5219 ( .A(n316), .B(n5567), .Z(n5566) );
  XOR U5220 ( .A(n5568), .B(n5565), .Z(n5567) );
  XOR U5221 ( .A(n5569), .B(n5570), .Z(n5557) );
  AND U5222 ( .A(n5571), .B(n5572), .Z(n5570) );
  XOR U5223 ( .A(n5569), .B(n5199), .Z(n5572) );
  XOR U5224 ( .A(n5573), .B(n5574), .Z(n5199) );
  AND U5225 ( .A(n318), .B(n5575), .Z(n5574) );
  XOR U5226 ( .A(n5576), .B(n5573), .Z(n5575) );
  XNOR U5227 ( .A(n5196), .B(n5569), .Z(n5571) );
  XOR U5228 ( .A(n5577), .B(n5578), .Z(n5196) );
  AND U5229 ( .A(n316), .B(n5579), .Z(n5578) );
  XOR U5230 ( .A(n5580), .B(n5577), .Z(n5579) );
  XOR U5231 ( .A(n5581), .B(n5582), .Z(n5569) );
  AND U5232 ( .A(n5583), .B(n5584), .Z(n5582) );
  XOR U5233 ( .A(n5581), .B(n5211), .Z(n5584) );
  XOR U5234 ( .A(n5585), .B(n5586), .Z(n5211) );
  AND U5235 ( .A(n318), .B(n5587), .Z(n5586) );
  XOR U5236 ( .A(n5588), .B(n5585), .Z(n5587) );
  XNOR U5237 ( .A(n5208), .B(n5581), .Z(n5583) );
  XOR U5238 ( .A(n5589), .B(n5590), .Z(n5208) );
  AND U5239 ( .A(n316), .B(n5591), .Z(n5590) );
  XOR U5240 ( .A(n5592), .B(n5589), .Z(n5591) );
  XOR U5241 ( .A(n5593), .B(n5594), .Z(n5581) );
  AND U5242 ( .A(n5595), .B(n5596), .Z(n5594) );
  XOR U5243 ( .A(n5593), .B(n5223), .Z(n5596) );
  XOR U5244 ( .A(n5597), .B(n5598), .Z(n5223) );
  AND U5245 ( .A(n318), .B(n5599), .Z(n5598) );
  XOR U5246 ( .A(n5600), .B(n5597), .Z(n5599) );
  XNOR U5247 ( .A(n5220), .B(n5593), .Z(n5595) );
  XOR U5248 ( .A(n5601), .B(n5602), .Z(n5220) );
  AND U5249 ( .A(n316), .B(n5603), .Z(n5602) );
  XOR U5250 ( .A(n5604), .B(n5601), .Z(n5603) );
  XOR U5251 ( .A(n5605), .B(n5606), .Z(n5593) );
  AND U5252 ( .A(n5607), .B(n5608), .Z(n5606) );
  XOR U5253 ( .A(n5605), .B(n5235), .Z(n5608) );
  XOR U5254 ( .A(n5609), .B(n5610), .Z(n5235) );
  AND U5255 ( .A(n318), .B(n5611), .Z(n5610) );
  XOR U5256 ( .A(n5612), .B(n5609), .Z(n5611) );
  XNOR U5257 ( .A(n5232), .B(n5605), .Z(n5607) );
  XOR U5258 ( .A(n5613), .B(n5614), .Z(n5232) );
  AND U5259 ( .A(n316), .B(n5615), .Z(n5614) );
  XOR U5260 ( .A(n5616), .B(n5613), .Z(n5615) );
  XOR U5261 ( .A(n5617), .B(n5618), .Z(n5605) );
  AND U5262 ( .A(n5619), .B(n5620), .Z(n5618) );
  XOR U5263 ( .A(n5617), .B(n5247), .Z(n5620) );
  XOR U5264 ( .A(n5621), .B(n5622), .Z(n5247) );
  AND U5265 ( .A(n318), .B(n5623), .Z(n5622) );
  XOR U5266 ( .A(n5624), .B(n5621), .Z(n5623) );
  XNOR U5267 ( .A(n5244), .B(n5617), .Z(n5619) );
  XOR U5268 ( .A(n5625), .B(n5626), .Z(n5244) );
  AND U5269 ( .A(n316), .B(n5627), .Z(n5626) );
  XOR U5270 ( .A(n5628), .B(n5625), .Z(n5627) );
  XOR U5271 ( .A(n5629), .B(n5630), .Z(n5617) );
  AND U5272 ( .A(n5631), .B(n5632), .Z(n5630) );
  XOR U5273 ( .A(n5629), .B(n5259), .Z(n5632) );
  XOR U5274 ( .A(n5633), .B(n5634), .Z(n5259) );
  AND U5275 ( .A(n318), .B(n5635), .Z(n5634) );
  XOR U5276 ( .A(n5636), .B(n5633), .Z(n5635) );
  XNOR U5277 ( .A(n5256), .B(n5629), .Z(n5631) );
  XOR U5278 ( .A(n5637), .B(n5638), .Z(n5256) );
  AND U5279 ( .A(n316), .B(n5639), .Z(n5638) );
  XOR U5280 ( .A(n5640), .B(n5637), .Z(n5639) );
  XOR U5281 ( .A(n5641), .B(n5642), .Z(n5629) );
  AND U5282 ( .A(n5643), .B(n5644), .Z(n5642) );
  XOR U5283 ( .A(n5641), .B(n5271), .Z(n5644) );
  XOR U5284 ( .A(n5645), .B(n5646), .Z(n5271) );
  AND U5285 ( .A(n318), .B(n5647), .Z(n5646) );
  XOR U5286 ( .A(n5648), .B(n5645), .Z(n5647) );
  XNOR U5287 ( .A(n5268), .B(n5641), .Z(n5643) );
  XOR U5288 ( .A(n5649), .B(n5650), .Z(n5268) );
  AND U5289 ( .A(n316), .B(n5651), .Z(n5650) );
  XOR U5290 ( .A(n5652), .B(n5649), .Z(n5651) );
  XOR U5291 ( .A(n5653), .B(n5654), .Z(n5641) );
  AND U5292 ( .A(n5655), .B(n5656), .Z(n5654) );
  XOR U5293 ( .A(n5653), .B(n5283), .Z(n5656) );
  XOR U5294 ( .A(n5657), .B(n5658), .Z(n5283) );
  AND U5295 ( .A(n318), .B(n5659), .Z(n5658) );
  XOR U5296 ( .A(n5660), .B(n5657), .Z(n5659) );
  XNOR U5297 ( .A(n5280), .B(n5653), .Z(n5655) );
  XOR U5298 ( .A(n5661), .B(n5662), .Z(n5280) );
  AND U5299 ( .A(n316), .B(n5663), .Z(n5662) );
  XOR U5300 ( .A(n5664), .B(n5661), .Z(n5663) );
  XOR U5301 ( .A(n5665), .B(n5666), .Z(n5653) );
  AND U5302 ( .A(n5667), .B(n5668), .Z(n5666) );
  XOR U5303 ( .A(n5665), .B(n5295), .Z(n5668) );
  XOR U5304 ( .A(n5669), .B(n5670), .Z(n5295) );
  AND U5305 ( .A(n318), .B(n5671), .Z(n5670) );
  XOR U5306 ( .A(n5672), .B(n5669), .Z(n5671) );
  XNOR U5307 ( .A(n5292), .B(n5665), .Z(n5667) );
  XOR U5308 ( .A(n5673), .B(n5674), .Z(n5292) );
  AND U5309 ( .A(n316), .B(n5675), .Z(n5674) );
  XOR U5310 ( .A(n5676), .B(n5673), .Z(n5675) );
  XOR U5311 ( .A(n5677), .B(n5678), .Z(n5665) );
  AND U5312 ( .A(n5679), .B(n5680), .Z(n5678) );
  XOR U5313 ( .A(n5677), .B(n5307), .Z(n5680) );
  XOR U5314 ( .A(n5681), .B(n5682), .Z(n5307) );
  AND U5315 ( .A(n318), .B(n5683), .Z(n5682) );
  XOR U5316 ( .A(n5684), .B(n5681), .Z(n5683) );
  XNOR U5317 ( .A(n5304), .B(n5677), .Z(n5679) );
  XOR U5318 ( .A(n5685), .B(n5686), .Z(n5304) );
  AND U5319 ( .A(n316), .B(n5687), .Z(n5686) );
  XOR U5320 ( .A(n5688), .B(n5685), .Z(n5687) );
  XOR U5321 ( .A(n5689), .B(n5690), .Z(n5677) );
  AND U5322 ( .A(n5691), .B(n5692), .Z(n5690) );
  XOR U5323 ( .A(n5689), .B(n5319), .Z(n5692) );
  XOR U5324 ( .A(n5693), .B(n5694), .Z(n5319) );
  AND U5325 ( .A(n318), .B(n5695), .Z(n5694) );
  XOR U5326 ( .A(n5696), .B(n5693), .Z(n5695) );
  XNOR U5327 ( .A(n5316), .B(n5689), .Z(n5691) );
  XOR U5328 ( .A(n5697), .B(n5698), .Z(n5316) );
  AND U5329 ( .A(n316), .B(n5699), .Z(n5698) );
  XOR U5330 ( .A(n5700), .B(n5697), .Z(n5699) );
  XOR U5331 ( .A(n5701), .B(n5702), .Z(n5689) );
  AND U5332 ( .A(n5703), .B(n5704), .Z(n5702) );
  XOR U5333 ( .A(n5701), .B(n5331), .Z(n5704) );
  XOR U5334 ( .A(n5705), .B(n5706), .Z(n5331) );
  AND U5335 ( .A(n318), .B(n5707), .Z(n5706) );
  XOR U5336 ( .A(n5708), .B(n5705), .Z(n5707) );
  XNOR U5337 ( .A(n5328), .B(n5701), .Z(n5703) );
  XOR U5338 ( .A(n5709), .B(n5710), .Z(n5328) );
  AND U5339 ( .A(n316), .B(n5711), .Z(n5710) );
  XOR U5340 ( .A(n5712), .B(n5709), .Z(n5711) );
  XOR U5341 ( .A(n5713), .B(n5714), .Z(n5701) );
  AND U5342 ( .A(n5715), .B(n5716), .Z(n5714) );
  XOR U5343 ( .A(n5713), .B(n5343), .Z(n5716) );
  XOR U5344 ( .A(n5717), .B(n5718), .Z(n5343) );
  AND U5345 ( .A(n318), .B(n5719), .Z(n5718) );
  XOR U5346 ( .A(n5720), .B(n5717), .Z(n5719) );
  XNOR U5347 ( .A(n5340), .B(n5713), .Z(n5715) );
  XOR U5348 ( .A(n5721), .B(n5722), .Z(n5340) );
  AND U5349 ( .A(n316), .B(n5723), .Z(n5722) );
  XOR U5350 ( .A(n5724), .B(n5721), .Z(n5723) );
  XOR U5351 ( .A(n5725), .B(n5726), .Z(n5713) );
  AND U5352 ( .A(n5727), .B(n5728), .Z(n5726) );
  XOR U5353 ( .A(n5725), .B(n5355), .Z(n5728) );
  XOR U5354 ( .A(n5729), .B(n5730), .Z(n5355) );
  AND U5355 ( .A(n318), .B(n5731), .Z(n5730) );
  XOR U5356 ( .A(n5732), .B(n5729), .Z(n5731) );
  XNOR U5357 ( .A(n5352), .B(n5725), .Z(n5727) );
  XOR U5358 ( .A(n5733), .B(n5734), .Z(n5352) );
  AND U5359 ( .A(n316), .B(n5735), .Z(n5734) );
  XOR U5360 ( .A(n5736), .B(n5733), .Z(n5735) );
  XOR U5361 ( .A(n5737), .B(n5738), .Z(n5725) );
  AND U5362 ( .A(n5739), .B(n5740), .Z(n5738) );
  XOR U5363 ( .A(n5737), .B(n5367), .Z(n5740) );
  XOR U5364 ( .A(n5741), .B(n5742), .Z(n5367) );
  AND U5365 ( .A(n318), .B(n5743), .Z(n5742) );
  XOR U5366 ( .A(n5744), .B(n5741), .Z(n5743) );
  XNOR U5367 ( .A(n5364), .B(n5737), .Z(n5739) );
  XOR U5368 ( .A(n5745), .B(n5746), .Z(n5364) );
  AND U5369 ( .A(n316), .B(n5747), .Z(n5746) );
  XOR U5370 ( .A(n5748), .B(n5745), .Z(n5747) );
  XOR U5371 ( .A(n5749), .B(n5750), .Z(n5737) );
  AND U5372 ( .A(n5751), .B(n5752), .Z(n5750) );
  XOR U5373 ( .A(n5749), .B(n5379), .Z(n5752) );
  XOR U5374 ( .A(n5753), .B(n5754), .Z(n5379) );
  AND U5375 ( .A(n318), .B(n5755), .Z(n5754) );
  XOR U5376 ( .A(n5756), .B(n5753), .Z(n5755) );
  XNOR U5377 ( .A(n5376), .B(n5749), .Z(n5751) );
  XOR U5378 ( .A(n5757), .B(n5758), .Z(n5376) );
  AND U5379 ( .A(n316), .B(n5759), .Z(n5758) );
  XOR U5380 ( .A(n5760), .B(n5757), .Z(n5759) );
  XOR U5381 ( .A(n5761), .B(n5762), .Z(n5749) );
  AND U5382 ( .A(n5763), .B(n5764), .Z(n5762) );
  XOR U5383 ( .A(n5391), .B(n5761), .Z(n5764) );
  XOR U5384 ( .A(n5765), .B(n5766), .Z(n5391) );
  AND U5385 ( .A(n318), .B(n5767), .Z(n5766) );
  XOR U5386 ( .A(n5765), .B(n5768), .Z(n5767) );
  XNOR U5387 ( .A(n5761), .B(n5388), .Z(n5763) );
  XOR U5388 ( .A(n5769), .B(n5770), .Z(n5388) );
  AND U5389 ( .A(n316), .B(n5771), .Z(n5770) );
  XOR U5390 ( .A(n5769), .B(n5772), .Z(n5771) );
  XOR U5391 ( .A(n5773), .B(n5774), .Z(n5761) );
  AND U5392 ( .A(n5775), .B(n5776), .Z(n5774) );
  XNOR U5393 ( .A(n5777), .B(n5404), .Z(n5776) );
  XOR U5394 ( .A(n5778), .B(n5779), .Z(n5404) );
  AND U5395 ( .A(n318), .B(n5780), .Z(n5779) );
  XOR U5396 ( .A(n5781), .B(n5778), .Z(n5780) );
  XNOR U5397 ( .A(n5401), .B(n5773), .Z(n5775) );
  XOR U5398 ( .A(n5782), .B(n5783), .Z(n5401) );
  AND U5399 ( .A(n316), .B(n5784), .Z(n5783) );
  XOR U5400 ( .A(n5785), .B(n5782), .Z(n5784) );
  IV U5401 ( .A(n5777), .Z(n5773) );
  AND U5402 ( .A(n5409), .B(n5412), .Z(n5777) );
  XNOR U5403 ( .A(n5786), .B(n5787), .Z(n5412) );
  AND U5404 ( .A(n318), .B(n5788), .Z(n5787) );
  XNOR U5405 ( .A(n5789), .B(n5786), .Z(n5788) );
  XOR U5406 ( .A(n5790), .B(n5791), .Z(n318) );
  AND U5407 ( .A(n5792), .B(n5793), .Z(n5791) );
  XOR U5408 ( .A(n5420), .B(n5790), .Z(n5793) );
  IV U5409 ( .A(n5794), .Z(n5420) );
  AND U5410 ( .A(p_input[3583]), .B(p_input[3551]), .Z(n5794) );
  XOR U5411 ( .A(n5790), .B(n5417), .Z(n5792) );
  AND U5412 ( .A(p_input[3487]), .B(p_input[3519]), .Z(n5417) );
  XOR U5413 ( .A(n5795), .B(n5796), .Z(n5790) );
  AND U5414 ( .A(n5797), .B(n5798), .Z(n5796) );
  XOR U5415 ( .A(n5795), .B(n5432), .Z(n5798) );
  XNOR U5416 ( .A(p_input[3550]), .B(n5799), .Z(n5432) );
  AND U5417 ( .A(n210), .B(n5800), .Z(n5799) );
  XOR U5418 ( .A(p_input[3582]), .B(p_input[3550]), .Z(n5800) );
  XNOR U5419 ( .A(n5429), .B(n5795), .Z(n5797) );
  XOR U5420 ( .A(n5801), .B(n5802), .Z(n5429) );
  AND U5421 ( .A(n208), .B(n5803), .Z(n5802) );
  XOR U5422 ( .A(p_input[3518]), .B(p_input[3486]), .Z(n5803) );
  XOR U5423 ( .A(n5804), .B(n5805), .Z(n5795) );
  AND U5424 ( .A(n5806), .B(n5807), .Z(n5805) );
  XOR U5425 ( .A(n5804), .B(n5444), .Z(n5807) );
  XNOR U5426 ( .A(p_input[3549]), .B(n5808), .Z(n5444) );
  AND U5427 ( .A(n210), .B(n5809), .Z(n5808) );
  XOR U5428 ( .A(p_input[3581]), .B(p_input[3549]), .Z(n5809) );
  XNOR U5429 ( .A(n5441), .B(n5804), .Z(n5806) );
  XOR U5430 ( .A(n5810), .B(n5811), .Z(n5441) );
  AND U5431 ( .A(n208), .B(n5812), .Z(n5811) );
  XOR U5432 ( .A(p_input[3517]), .B(p_input[3485]), .Z(n5812) );
  XOR U5433 ( .A(n5813), .B(n5814), .Z(n5804) );
  AND U5434 ( .A(n5815), .B(n5816), .Z(n5814) );
  XOR U5435 ( .A(n5813), .B(n5456), .Z(n5816) );
  XNOR U5436 ( .A(p_input[3548]), .B(n5817), .Z(n5456) );
  AND U5437 ( .A(n210), .B(n5818), .Z(n5817) );
  XOR U5438 ( .A(p_input[3580]), .B(p_input[3548]), .Z(n5818) );
  XNOR U5439 ( .A(n5453), .B(n5813), .Z(n5815) );
  XOR U5440 ( .A(n5819), .B(n5820), .Z(n5453) );
  AND U5441 ( .A(n208), .B(n5821), .Z(n5820) );
  XOR U5442 ( .A(p_input[3516]), .B(p_input[3484]), .Z(n5821) );
  XOR U5443 ( .A(n5822), .B(n5823), .Z(n5813) );
  AND U5444 ( .A(n5824), .B(n5825), .Z(n5823) );
  XOR U5445 ( .A(n5822), .B(n5468), .Z(n5825) );
  XNOR U5446 ( .A(p_input[3547]), .B(n5826), .Z(n5468) );
  AND U5447 ( .A(n210), .B(n5827), .Z(n5826) );
  XOR U5448 ( .A(p_input[3579]), .B(p_input[3547]), .Z(n5827) );
  XNOR U5449 ( .A(n5465), .B(n5822), .Z(n5824) );
  XOR U5450 ( .A(n5828), .B(n5829), .Z(n5465) );
  AND U5451 ( .A(n208), .B(n5830), .Z(n5829) );
  XOR U5452 ( .A(p_input[3515]), .B(p_input[3483]), .Z(n5830) );
  XOR U5453 ( .A(n5831), .B(n5832), .Z(n5822) );
  AND U5454 ( .A(n5833), .B(n5834), .Z(n5832) );
  XOR U5455 ( .A(n5831), .B(n5480), .Z(n5834) );
  XNOR U5456 ( .A(p_input[3546]), .B(n5835), .Z(n5480) );
  AND U5457 ( .A(n210), .B(n5836), .Z(n5835) );
  XOR U5458 ( .A(p_input[3578]), .B(p_input[3546]), .Z(n5836) );
  XNOR U5459 ( .A(n5477), .B(n5831), .Z(n5833) );
  XOR U5460 ( .A(n5837), .B(n5838), .Z(n5477) );
  AND U5461 ( .A(n208), .B(n5839), .Z(n5838) );
  XOR U5462 ( .A(p_input[3514]), .B(p_input[3482]), .Z(n5839) );
  XOR U5463 ( .A(n5840), .B(n5841), .Z(n5831) );
  AND U5464 ( .A(n5842), .B(n5843), .Z(n5841) );
  XOR U5465 ( .A(n5840), .B(n5492), .Z(n5843) );
  XNOR U5466 ( .A(p_input[3545]), .B(n5844), .Z(n5492) );
  AND U5467 ( .A(n210), .B(n5845), .Z(n5844) );
  XOR U5468 ( .A(p_input[3577]), .B(p_input[3545]), .Z(n5845) );
  XNOR U5469 ( .A(n5489), .B(n5840), .Z(n5842) );
  XOR U5470 ( .A(n5846), .B(n5847), .Z(n5489) );
  AND U5471 ( .A(n208), .B(n5848), .Z(n5847) );
  XOR U5472 ( .A(p_input[3513]), .B(p_input[3481]), .Z(n5848) );
  XOR U5473 ( .A(n5849), .B(n5850), .Z(n5840) );
  AND U5474 ( .A(n5851), .B(n5852), .Z(n5850) );
  XOR U5475 ( .A(n5849), .B(n5504), .Z(n5852) );
  XNOR U5476 ( .A(p_input[3544]), .B(n5853), .Z(n5504) );
  AND U5477 ( .A(n210), .B(n5854), .Z(n5853) );
  XOR U5478 ( .A(p_input[3576]), .B(p_input[3544]), .Z(n5854) );
  XNOR U5479 ( .A(n5501), .B(n5849), .Z(n5851) );
  XOR U5480 ( .A(n5855), .B(n5856), .Z(n5501) );
  AND U5481 ( .A(n208), .B(n5857), .Z(n5856) );
  XOR U5482 ( .A(p_input[3512]), .B(p_input[3480]), .Z(n5857) );
  XOR U5483 ( .A(n5858), .B(n5859), .Z(n5849) );
  AND U5484 ( .A(n5860), .B(n5861), .Z(n5859) );
  XOR U5485 ( .A(n5858), .B(n5516), .Z(n5861) );
  XNOR U5486 ( .A(p_input[3543]), .B(n5862), .Z(n5516) );
  AND U5487 ( .A(n210), .B(n5863), .Z(n5862) );
  XOR U5488 ( .A(p_input[3575]), .B(p_input[3543]), .Z(n5863) );
  XNOR U5489 ( .A(n5513), .B(n5858), .Z(n5860) );
  XOR U5490 ( .A(n5864), .B(n5865), .Z(n5513) );
  AND U5491 ( .A(n208), .B(n5866), .Z(n5865) );
  XOR U5492 ( .A(p_input[3511]), .B(p_input[3479]), .Z(n5866) );
  XOR U5493 ( .A(n5867), .B(n5868), .Z(n5858) );
  AND U5494 ( .A(n5869), .B(n5870), .Z(n5868) );
  XOR U5495 ( .A(n5867), .B(n5528), .Z(n5870) );
  XNOR U5496 ( .A(p_input[3542]), .B(n5871), .Z(n5528) );
  AND U5497 ( .A(n210), .B(n5872), .Z(n5871) );
  XOR U5498 ( .A(p_input[3574]), .B(p_input[3542]), .Z(n5872) );
  XNOR U5499 ( .A(n5525), .B(n5867), .Z(n5869) );
  XOR U5500 ( .A(n5873), .B(n5874), .Z(n5525) );
  AND U5501 ( .A(n208), .B(n5875), .Z(n5874) );
  XOR U5502 ( .A(p_input[3510]), .B(p_input[3478]), .Z(n5875) );
  XOR U5503 ( .A(n5876), .B(n5877), .Z(n5867) );
  AND U5504 ( .A(n5878), .B(n5879), .Z(n5877) );
  XOR U5505 ( .A(n5876), .B(n5540), .Z(n5879) );
  XNOR U5506 ( .A(p_input[3541]), .B(n5880), .Z(n5540) );
  AND U5507 ( .A(n210), .B(n5881), .Z(n5880) );
  XOR U5508 ( .A(p_input[3573]), .B(p_input[3541]), .Z(n5881) );
  XNOR U5509 ( .A(n5537), .B(n5876), .Z(n5878) );
  XOR U5510 ( .A(n5882), .B(n5883), .Z(n5537) );
  AND U5511 ( .A(n208), .B(n5884), .Z(n5883) );
  XOR U5512 ( .A(p_input[3509]), .B(p_input[3477]), .Z(n5884) );
  XOR U5513 ( .A(n5885), .B(n5886), .Z(n5876) );
  AND U5514 ( .A(n5887), .B(n5888), .Z(n5886) );
  XOR U5515 ( .A(n5885), .B(n5552), .Z(n5888) );
  XNOR U5516 ( .A(p_input[3540]), .B(n5889), .Z(n5552) );
  AND U5517 ( .A(n210), .B(n5890), .Z(n5889) );
  XOR U5518 ( .A(p_input[3572]), .B(p_input[3540]), .Z(n5890) );
  XNOR U5519 ( .A(n5549), .B(n5885), .Z(n5887) );
  XOR U5520 ( .A(n5891), .B(n5892), .Z(n5549) );
  AND U5521 ( .A(n208), .B(n5893), .Z(n5892) );
  XOR U5522 ( .A(p_input[3508]), .B(p_input[3476]), .Z(n5893) );
  XOR U5523 ( .A(n5894), .B(n5895), .Z(n5885) );
  AND U5524 ( .A(n5896), .B(n5897), .Z(n5895) );
  XOR U5525 ( .A(n5894), .B(n5564), .Z(n5897) );
  XNOR U5526 ( .A(p_input[3539]), .B(n5898), .Z(n5564) );
  AND U5527 ( .A(n210), .B(n5899), .Z(n5898) );
  XOR U5528 ( .A(p_input[3571]), .B(p_input[3539]), .Z(n5899) );
  XNOR U5529 ( .A(n5561), .B(n5894), .Z(n5896) );
  XOR U5530 ( .A(n5900), .B(n5901), .Z(n5561) );
  AND U5531 ( .A(n208), .B(n5902), .Z(n5901) );
  XOR U5532 ( .A(p_input[3507]), .B(p_input[3475]), .Z(n5902) );
  XOR U5533 ( .A(n5903), .B(n5904), .Z(n5894) );
  AND U5534 ( .A(n5905), .B(n5906), .Z(n5904) );
  XOR U5535 ( .A(n5903), .B(n5576), .Z(n5906) );
  XNOR U5536 ( .A(p_input[3538]), .B(n5907), .Z(n5576) );
  AND U5537 ( .A(n210), .B(n5908), .Z(n5907) );
  XOR U5538 ( .A(p_input[3570]), .B(p_input[3538]), .Z(n5908) );
  XNOR U5539 ( .A(n5573), .B(n5903), .Z(n5905) );
  XOR U5540 ( .A(n5909), .B(n5910), .Z(n5573) );
  AND U5541 ( .A(n208), .B(n5911), .Z(n5910) );
  XOR U5542 ( .A(p_input[3506]), .B(p_input[3474]), .Z(n5911) );
  XOR U5543 ( .A(n5912), .B(n5913), .Z(n5903) );
  AND U5544 ( .A(n5914), .B(n5915), .Z(n5913) );
  XOR U5545 ( .A(n5912), .B(n5588), .Z(n5915) );
  XNOR U5546 ( .A(p_input[3537]), .B(n5916), .Z(n5588) );
  AND U5547 ( .A(n210), .B(n5917), .Z(n5916) );
  XOR U5548 ( .A(p_input[3569]), .B(p_input[3537]), .Z(n5917) );
  XNOR U5549 ( .A(n5585), .B(n5912), .Z(n5914) );
  XOR U5550 ( .A(n5918), .B(n5919), .Z(n5585) );
  AND U5551 ( .A(n208), .B(n5920), .Z(n5919) );
  XOR U5552 ( .A(p_input[3505]), .B(p_input[3473]), .Z(n5920) );
  XOR U5553 ( .A(n5921), .B(n5922), .Z(n5912) );
  AND U5554 ( .A(n5923), .B(n5924), .Z(n5922) );
  XOR U5555 ( .A(n5921), .B(n5600), .Z(n5924) );
  XNOR U5556 ( .A(p_input[3536]), .B(n5925), .Z(n5600) );
  AND U5557 ( .A(n210), .B(n5926), .Z(n5925) );
  XOR U5558 ( .A(p_input[3568]), .B(p_input[3536]), .Z(n5926) );
  XNOR U5559 ( .A(n5597), .B(n5921), .Z(n5923) );
  XOR U5560 ( .A(n5927), .B(n5928), .Z(n5597) );
  AND U5561 ( .A(n208), .B(n5929), .Z(n5928) );
  XOR U5562 ( .A(p_input[3504]), .B(p_input[3472]), .Z(n5929) );
  XOR U5563 ( .A(n5930), .B(n5931), .Z(n5921) );
  AND U5564 ( .A(n5932), .B(n5933), .Z(n5931) );
  XOR U5565 ( .A(n5930), .B(n5612), .Z(n5933) );
  XNOR U5566 ( .A(p_input[3535]), .B(n5934), .Z(n5612) );
  AND U5567 ( .A(n210), .B(n5935), .Z(n5934) );
  XOR U5568 ( .A(p_input[3567]), .B(p_input[3535]), .Z(n5935) );
  XNOR U5569 ( .A(n5609), .B(n5930), .Z(n5932) );
  XOR U5570 ( .A(n5936), .B(n5937), .Z(n5609) );
  AND U5571 ( .A(n208), .B(n5938), .Z(n5937) );
  XOR U5572 ( .A(p_input[3503]), .B(p_input[3471]), .Z(n5938) );
  XOR U5573 ( .A(n5939), .B(n5940), .Z(n5930) );
  AND U5574 ( .A(n5941), .B(n5942), .Z(n5940) );
  XOR U5575 ( .A(n5939), .B(n5624), .Z(n5942) );
  XNOR U5576 ( .A(p_input[3534]), .B(n5943), .Z(n5624) );
  AND U5577 ( .A(n210), .B(n5944), .Z(n5943) );
  XOR U5578 ( .A(p_input[3566]), .B(p_input[3534]), .Z(n5944) );
  XNOR U5579 ( .A(n5621), .B(n5939), .Z(n5941) );
  XOR U5580 ( .A(n5945), .B(n5946), .Z(n5621) );
  AND U5581 ( .A(n208), .B(n5947), .Z(n5946) );
  XOR U5582 ( .A(p_input[3502]), .B(p_input[3470]), .Z(n5947) );
  XOR U5583 ( .A(n5948), .B(n5949), .Z(n5939) );
  AND U5584 ( .A(n5950), .B(n5951), .Z(n5949) );
  XOR U5585 ( .A(n5948), .B(n5636), .Z(n5951) );
  XNOR U5586 ( .A(p_input[3533]), .B(n5952), .Z(n5636) );
  AND U5587 ( .A(n210), .B(n5953), .Z(n5952) );
  XOR U5588 ( .A(p_input[3565]), .B(p_input[3533]), .Z(n5953) );
  XNOR U5589 ( .A(n5633), .B(n5948), .Z(n5950) );
  XOR U5590 ( .A(n5954), .B(n5955), .Z(n5633) );
  AND U5591 ( .A(n208), .B(n5956), .Z(n5955) );
  XOR U5592 ( .A(p_input[3501]), .B(p_input[3469]), .Z(n5956) );
  XOR U5593 ( .A(n5957), .B(n5958), .Z(n5948) );
  AND U5594 ( .A(n5959), .B(n5960), .Z(n5958) );
  XOR U5595 ( .A(n5957), .B(n5648), .Z(n5960) );
  XNOR U5596 ( .A(p_input[3532]), .B(n5961), .Z(n5648) );
  AND U5597 ( .A(n210), .B(n5962), .Z(n5961) );
  XOR U5598 ( .A(p_input[3564]), .B(p_input[3532]), .Z(n5962) );
  XNOR U5599 ( .A(n5645), .B(n5957), .Z(n5959) );
  XOR U5600 ( .A(n5963), .B(n5964), .Z(n5645) );
  AND U5601 ( .A(n208), .B(n5965), .Z(n5964) );
  XOR U5602 ( .A(p_input[3500]), .B(p_input[3468]), .Z(n5965) );
  XOR U5603 ( .A(n5966), .B(n5967), .Z(n5957) );
  AND U5604 ( .A(n5968), .B(n5969), .Z(n5967) );
  XOR U5605 ( .A(n5966), .B(n5660), .Z(n5969) );
  XNOR U5606 ( .A(p_input[3531]), .B(n5970), .Z(n5660) );
  AND U5607 ( .A(n210), .B(n5971), .Z(n5970) );
  XOR U5608 ( .A(p_input[3563]), .B(p_input[3531]), .Z(n5971) );
  XNOR U5609 ( .A(n5657), .B(n5966), .Z(n5968) );
  XOR U5610 ( .A(n5972), .B(n5973), .Z(n5657) );
  AND U5611 ( .A(n208), .B(n5974), .Z(n5973) );
  XOR U5612 ( .A(p_input[3499]), .B(p_input[3467]), .Z(n5974) );
  XOR U5613 ( .A(n5975), .B(n5976), .Z(n5966) );
  AND U5614 ( .A(n5977), .B(n5978), .Z(n5976) );
  XOR U5615 ( .A(n5975), .B(n5672), .Z(n5978) );
  XNOR U5616 ( .A(p_input[3530]), .B(n5979), .Z(n5672) );
  AND U5617 ( .A(n210), .B(n5980), .Z(n5979) );
  XOR U5618 ( .A(p_input[3562]), .B(p_input[3530]), .Z(n5980) );
  XNOR U5619 ( .A(n5669), .B(n5975), .Z(n5977) );
  XOR U5620 ( .A(n5981), .B(n5982), .Z(n5669) );
  AND U5621 ( .A(n208), .B(n5983), .Z(n5982) );
  XOR U5622 ( .A(p_input[3498]), .B(p_input[3466]), .Z(n5983) );
  XOR U5623 ( .A(n5984), .B(n5985), .Z(n5975) );
  AND U5624 ( .A(n5986), .B(n5987), .Z(n5985) );
  XOR U5625 ( .A(n5984), .B(n5684), .Z(n5987) );
  XNOR U5626 ( .A(p_input[3529]), .B(n5988), .Z(n5684) );
  AND U5627 ( .A(n210), .B(n5989), .Z(n5988) );
  XOR U5628 ( .A(p_input[3561]), .B(p_input[3529]), .Z(n5989) );
  XNOR U5629 ( .A(n5681), .B(n5984), .Z(n5986) );
  XOR U5630 ( .A(n5990), .B(n5991), .Z(n5681) );
  AND U5631 ( .A(n208), .B(n5992), .Z(n5991) );
  XOR U5632 ( .A(p_input[3497]), .B(p_input[3465]), .Z(n5992) );
  XOR U5633 ( .A(n5993), .B(n5994), .Z(n5984) );
  AND U5634 ( .A(n5995), .B(n5996), .Z(n5994) );
  XOR U5635 ( .A(n5993), .B(n5696), .Z(n5996) );
  XNOR U5636 ( .A(p_input[3528]), .B(n5997), .Z(n5696) );
  AND U5637 ( .A(n210), .B(n5998), .Z(n5997) );
  XOR U5638 ( .A(p_input[3560]), .B(p_input[3528]), .Z(n5998) );
  XNOR U5639 ( .A(n5693), .B(n5993), .Z(n5995) );
  XOR U5640 ( .A(n5999), .B(n6000), .Z(n5693) );
  AND U5641 ( .A(n208), .B(n6001), .Z(n6000) );
  XOR U5642 ( .A(p_input[3496]), .B(p_input[3464]), .Z(n6001) );
  XOR U5643 ( .A(n6002), .B(n6003), .Z(n5993) );
  AND U5644 ( .A(n6004), .B(n6005), .Z(n6003) );
  XOR U5645 ( .A(n6002), .B(n5708), .Z(n6005) );
  XNOR U5646 ( .A(p_input[3527]), .B(n6006), .Z(n5708) );
  AND U5647 ( .A(n210), .B(n6007), .Z(n6006) );
  XOR U5648 ( .A(p_input[3559]), .B(p_input[3527]), .Z(n6007) );
  XNOR U5649 ( .A(n5705), .B(n6002), .Z(n6004) );
  XOR U5650 ( .A(n6008), .B(n6009), .Z(n5705) );
  AND U5651 ( .A(n208), .B(n6010), .Z(n6009) );
  XOR U5652 ( .A(p_input[3495]), .B(p_input[3463]), .Z(n6010) );
  XOR U5653 ( .A(n6011), .B(n6012), .Z(n6002) );
  AND U5654 ( .A(n6013), .B(n6014), .Z(n6012) );
  XOR U5655 ( .A(n6011), .B(n5720), .Z(n6014) );
  XNOR U5656 ( .A(p_input[3526]), .B(n6015), .Z(n5720) );
  AND U5657 ( .A(n210), .B(n6016), .Z(n6015) );
  XOR U5658 ( .A(p_input[3558]), .B(p_input[3526]), .Z(n6016) );
  XNOR U5659 ( .A(n5717), .B(n6011), .Z(n6013) );
  XOR U5660 ( .A(n6017), .B(n6018), .Z(n5717) );
  AND U5661 ( .A(n208), .B(n6019), .Z(n6018) );
  XOR U5662 ( .A(p_input[3494]), .B(p_input[3462]), .Z(n6019) );
  XOR U5663 ( .A(n6020), .B(n6021), .Z(n6011) );
  AND U5664 ( .A(n6022), .B(n6023), .Z(n6021) );
  XOR U5665 ( .A(n6020), .B(n5732), .Z(n6023) );
  XNOR U5666 ( .A(p_input[3525]), .B(n6024), .Z(n5732) );
  AND U5667 ( .A(n210), .B(n6025), .Z(n6024) );
  XOR U5668 ( .A(p_input[3557]), .B(p_input[3525]), .Z(n6025) );
  XNOR U5669 ( .A(n5729), .B(n6020), .Z(n6022) );
  XOR U5670 ( .A(n6026), .B(n6027), .Z(n5729) );
  AND U5671 ( .A(n208), .B(n6028), .Z(n6027) );
  XOR U5672 ( .A(p_input[3493]), .B(p_input[3461]), .Z(n6028) );
  XOR U5673 ( .A(n6029), .B(n6030), .Z(n6020) );
  AND U5674 ( .A(n6031), .B(n6032), .Z(n6030) );
  XOR U5675 ( .A(n6029), .B(n5744), .Z(n6032) );
  XNOR U5676 ( .A(p_input[3524]), .B(n6033), .Z(n5744) );
  AND U5677 ( .A(n210), .B(n6034), .Z(n6033) );
  XOR U5678 ( .A(p_input[3556]), .B(p_input[3524]), .Z(n6034) );
  XNOR U5679 ( .A(n5741), .B(n6029), .Z(n6031) );
  XOR U5680 ( .A(n6035), .B(n6036), .Z(n5741) );
  AND U5681 ( .A(n208), .B(n6037), .Z(n6036) );
  XOR U5682 ( .A(p_input[3492]), .B(p_input[3460]), .Z(n6037) );
  XOR U5683 ( .A(n6038), .B(n6039), .Z(n6029) );
  AND U5684 ( .A(n6040), .B(n6041), .Z(n6039) );
  XOR U5685 ( .A(n6038), .B(n5756), .Z(n6041) );
  XNOR U5686 ( .A(p_input[3523]), .B(n6042), .Z(n5756) );
  AND U5687 ( .A(n210), .B(n6043), .Z(n6042) );
  XOR U5688 ( .A(p_input[3555]), .B(p_input[3523]), .Z(n6043) );
  XNOR U5689 ( .A(n5753), .B(n6038), .Z(n6040) );
  XOR U5690 ( .A(n6044), .B(n6045), .Z(n5753) );
  AND U5691 ( .A(n208), .B(n6046), .Z(n6045) );
  XOR U5692 ( .A(p_input[3491]), .B(p_input[3459]), .Z(n6046) );
  XOR U5693 ( .A(n6047), .B(n6048), .Z(n6038) );
  AND U5694 ( .A(n6049), .B(n6050), .Z(n6048) );
  XOR U5695 ( .A(n5768), .B(n6047), .Z(n6050) );
  XNOR U5696 ( .A(p_input[3522]), .B(n6051), .Z(n5768) );
  AND U5697 ( .A(n210), .B(n6052), .Z(n6051) );
  XOR U5698 ( .A(p_input[3554]), .B(p_input[3522]), .Z(n6052) );
  XNOR U5699 ( .A(n6047), .B(n5765), .Z(n6049) );
  XOR U5700 ( .A(n6053), .B(n6054), .Z(n5765) );
  AND U5701 ( .A(n208), .B(n6055), .Z(n6054) );
  XOR U5702 ( .A(p_input[3490]), .B(p_input[3458]), .Z(n6055) );
  XOR U5703 ( .A(n6056), .B(n6057), .Z(n6047) );
  AND U5704 ( .A(n6058), .B(n6059), .Z(n6057) );
  XNOR U5705 ( .A(n6060), .B(n5781), .Z(n6059) );
  XNOR U5706 ( .A(p_input[3521]), .B(n6061), .Z(n5781) );
  AND U5707 ( .A(n210), .B(n6062), .Z(n6061) );
  XNOR U5708 ( .A(p_input[3553]), .B(n6063), .Z(n6062) );
  IV U5709 ( .A(p_input[3521]), .Z(n6063) );
  XNOR U5710 ( .A(n5778), .B(n6056), .Z(n6058) );
  XNOR U5711 ( .A(p_input[3457]), .B(n6064), .Z(n5778) );
  AND U5712 ( .A(n208), .B(n6065), .Z(n6064) );
  XOR U5713 ( .A(p_input[3489]), .B(p_input[3457]), .Z(n6065) );
  IV U5714 ( .A(n6060), .Z(n6056) );
  AND U5715 ( .A(n5786), .B(n5789), .Z(n6060) );
  XOR U5716 ( .A(p_input[3520]), .B(n6066), .Z(n5789) );
  AND U5717 ( .A(n210), .B(n6067), .Z(n6066) );
  XOR U5718 ( .A(p_input[3552]), .B(p_input[3520]), .Z(n6067) );
  XOR U5719 ( .A(n6068), .B(n6069), .Z(n210) );
  AND U5720 ( .A(n6070), .B(n6071), .Z(n6069) );
  XNOR U5721 ( .A(p_input[3583]), .B(n6068), .Z(n6071) );
  XOR U5722 ( .A(n6068), .B(p_input[3551]), .Z(n6070) );
  XOR U5723 ( .A(n6072), .B(n6073), .Z(n6068) );
  AND U5724 ( .A(n6074), .B(n6075), .Z(n6073) );
  XNOR U5725 ( .A(p_input[3582]), .B(n6072), .Z(n6075) );
  XOR U5726 ( .A(n6072), .B(p_input[3550]), .Z(n6074) );
  XOR U5727 ( .A(n6076), .B(n6077), .Z(n6072) );
  AND U5728 ( .A(n6078), .B(n6079), .Z(n6077) );
  XNOR U5729 ( .A(p_input[3581]), .B(n6076), .Z(n6079) );
  XOR U5730 ( .A(n6076), .B(p_input[3549]), .Z(n6078) );
  XOR U5731 ( .A(n6080), .B(n6081), .Z(n6076) );
  AND U5732 ( .A(n6082), .B(n6083), .Z(n6081) );
  XNOR U5733 ( .A(p_input[3580]), .B(n6080), .Z(n6083) );
  XOR U5734 ( .A(n6080), .B(p_input[3548]), .Z(n6082) );
  XOR U5735 ( .A(n6084), .B(n6085), .Z(n6080) );
  AND U5736 ( .A(n6086), .B(n6087), .Z(n6085) );
  XNOR U5737 ( .A(p_input[3579]), .B(n6084), .Z(n6087) );
  XOR U5738 ( .A(n6084), .B(p_input[3547]), .Z(n6086) );
  XOR U5739 ( .A(n6088), .B(n6089), .Z(n6084) );
  AND U5740 ( .A(n6090), .B(n6091), .Z(n6089) );
  XNOR U5741 ( .A(p_input[3578]), .B(n6088), .Z(n6091) );
  XOR U5742 ( .A(n6088), .B(p_input[3546]), .Z(n6090) );
  XOR U5743 ( .A(n6092), .B(n6093), .Z(n6088) );
  AND U5744 ( .A(n6094), .B(n6095), .Z(n6093) );
  XNOR U5745 ( .A(p_input[3577]), .B(n6092), .Z(n6095) );
  XOR U5746 ( .A(n6092), .B(p_input[3545]), .Z(n6094) );
  XOR U5747 ( .A(n6096), .B(n6097), .Z(n6092) );
  AND U5748 ( .A(n6098), .B(n6099), .Z(n6097) );
  XNOR U5749 ( .A(p_input[3576]), .B(n6096), .Z(n6099) );
  XOR U5750 ( .A(n6096), .B(p_input[3544]), .Z(n6098) );
  XOR U5751 ( .A(n6100), .B(n6101), .Z(n6096) );
  AND U5752 ( .A(n6102), .B(n6103), .Z(n6101) );
  XNOR U5753 ( .A(p_input[3575]), .B(n6100), .Z(n6103) );
  XOR U5754 ( .A(n6100), .B(p_input[3543]), .Z(n6102) );
  XOR U5755 ( .A(n6104), .B(n6105), .Z(n6100) );
  AND U5756 ( .A(n6106), .B(n6107), .Z(n6105) );
  XNOR U5757 ( .A(p_input[3574]), .B(n6104), .Z(n6107) );
  XOR U5758 ( .A(n6104), .B(p_input[3542]), .Z(n6106) );
  XOR U5759 ( .A(n6108), .B(n6109), .Z(n6104) );
  AND U5760 ( .A(n6110), .B(n6111), .Z(n6109) );
  XNOR U5761 ( .A(p_input[3573]), .B(n6108), .Z(n6111) );
  XOR U5762 ( .A(n6108), .B(p_input[3541]), .Z(n6110) );
  XOR U5763 ( .A(n6112), .B(n6113), .Z(n6108) );
  AND U5764 ( .A(n6114), .B(n6115), .Z(n6113) );
  XNOR U5765 ( .A(p_input[3572]), .B(n6112), .Z(n6115) );
  XOR U5766 ( .A(n6112), .B(p_input[3540]), .Z(n6114) );
  XOR U5767 ( .A(n6116), .B(n6117), .Z(n6112) );
  AND U5768 ( .A(n6118), .B(n6119), .Z(n6117) );
  XNOR U5769 ( .A(p_input[3571]), .B(n6116), .Z(n6119) );
  XOR U5770 ( .A(n6116), .B(p_input[3539]), .Z(n6118) );
  XOR U5771 ( .A(n6120), .B(n6121), .Z(n6116) );
  AND U5772 ( .A(n6122), .B(n6123), .Z(n6121) );
  XNOR U5773 ( .A(p_input[3570]), .B(n6120), .Z(n6123) );
  XOR U5774 ( .A(n6120), .B(p_input[3538]), .Z(n6122) );
  XOR U5775 ( .A(n6124), .B(n6125), .Z(n6120) );
  AND U5776 ( .A(n6126), .B(n6127), .Z(n6125) );
  XNOR U5777 ( .A(p_input[3569]), .B(n6124), .Z(n6127) );
  XOR U5778 ( .A(n6124), .B(p_input[3537]), .Z(n6126) );
  XOR U5779 ( .A(n6128), .B(n6129), .Z(n6124) );
  AND U5780 ( .A(n6130), .B(n6131), .Z(n6129) );
  XNOR U5781 ( .A(p_input[3568]), .B(n6128), .Z(n6131) );
  XOR U5782 ( .A(n6128), .B(p_input[3536]), .Z(n6130) );
  XOR U5783 ( .A(n6132), .B(n6133), .Z(n6128) );
  AND U5784 ( .A(n6134), .B(n6135), .Z(n6133) );
  XNOR U5785 ( .A(p_input[3567]), .B(n6132), .Z(n6135) );
  XOR U5786 ( .A(n6132), .B(p_input[3535]), .Z(n6134) );
  XOR U5787 ( .A(n6136), .B(n6137), .Z(n6132) );
  AND U5788 ( .A(n6138), .B(n6139), .Z(n6137) );
  XNOR U5789 ( .A(p_input[3566]), .B(n6136), .Z(n6139) );
  XOR U5790 ( .A(n6136), .B(p_input[3534]), .Z(n6138) );
  XOR U5791 ( .A(n6140), .B(n6141), .Z(n6136) );
  AND U5792 ( .A(n6142), .B(n6143), .Z(n6141) );
  XNOR U5793 ( .A(p_input[3565]), .B(n6140), .Z(n6143) );
  XOR U5794 ( .A(n6140), .B(p_input[3533]), .Z(n6142) );
  XOR U5795 ( .A(n6144), .B(n6145), .Z(n6140) );
  AND U5796 ( .A(n6146), .B(n6147), .Z(n6145) );
  XNOR U5797 ( .A(p_input[3564]), .B(n6144), .Z(n6147) );
  XOR U5798 ( .A(n6144), .B(p_input[3532]), .Z(n6146) );
  XOR U5799 ( .A(n6148), .B(n6149), .Z(n6144) );
  AND U5800 ( .A(n6150), .B(n6151), .Z(n6149) );
  XNOR U5801 ( .A(p_input[3563]), .B(n6148), .Z(n6151) );
  XOR U5802 ( .A(n6148), .B(p_input[3531]), .Z(n6150) );
  XOR U5803 ( .A(n6152), .B(n6153), .Z(n6148) );
  AND U5804 ( .A(n6154), .B(n6155), .Z(n6153) );
  XNOR U5805 ( .A(p_input[3562]), .B(n6152), .Z(n6155) );
  XOR U5806 ( .A(n6152), .B(p_input[3530]), .Z(n6154) );
  XOR U5807 ( .A(n6156), .B(n6157), .Z(n6152) );
  AND U5808 ( .A(n6158), .B(n6159), .Z(n6157) );
  XNOR U5809 ( .A(p_input[3561]), .B(n6156), .Z(n6159) );
  XOR U5810 ( .A(n6156), .B(p_input[3529]), .Z(n6158) );
  XOR U5811 ( .A(n6160), .B(n6161), .Z(n6156) );
  AND U5812 ( .A(n6162), .B(n6163), .Z(n6161) );
  XNOR U5813 ( .A(p_input[3560]), .B(n6160), .Z(n6163) );
  XOR U5814 ( .A(n6160), .B(p_input[3528]), .Z(n6162) );
  XOR U5815 ( .A(n6164), .B(n6165), .Z(n6160) );
  AND U5816 ( .A(n6166), .B(n6167), .Z(n6165) );
  XNOR U5817 ( .A(p_input[3559]), .B(n6164), .Z(n6167) );
  XOR U5818 ( .A(n6164), .B(p_input[3527]), .Z(n6166) );
  XOR U5819 ( .A(n6168), .B(n6169), .Z(n6164) );
  AND U5820 ( .A(n6170), .B(n6171), .Z(n6169) );
  XNOR U5821 ( .A(p_input[3558]), .B(n6168), .Z(n6171) );
  XOR U5822 ( .A(n6168), .B(p_input[3526]), .Z(n6170) );
  XOR U5823 ( .A(n6172), .B(n6173), .Z(n6168) );
  AND U5824 ( .A(n6174), .B(n6175), .Z(n6173) );
  XNOR U5825 ( .A(p_input[3557]), .B(n6172), .Z(n6175) );
  XOR U5826 ( .A(n6172), .B(p_input[3525]), .Z(n6174) );
  XOR U5827 ( .A(n6176), .B(n6177), .Z(n6172) );
  AND U5828 ( .A(n6178), .B(n6179), .Z(n6177) );
  XNOR U5829 ( .A(p_input[3556]), .B(n6176), .Z(n6179) );
  XOR U5830 ( .A(n6176), .B(p_input[3524]), .Z(n6178) );
  XOR U5831 ( .A(n6180), .B(n6181), .Z(n6176) );
  AND U5832 ( .A(n6182), .B(n6183), .Z(n6181) );
  XNOR U5833 ( .A(p_input[3555]), .B(n6180), .Z(n6183) );
  XOR U5834 ( .A(n6180), .B(p_input[3523]), .Z(n6182) );
  XOR U5835 ( .A(n6184), .B(n6185), .Z(n6180) );
  AND U5836 ( .A(n6186), .B(n6187), .Z(n6185) );
  XNOR U5837 ( .A(p_input[3554]), .B(n6184), .Z(n6187) );
  XOR U5838 ( .A(n6184), .B(p_input[3522]), .Z(n6186) );
  XNOR U5839 ( .A(n6188), .B(n6189), .Z(n6184) );
  AND U5840 ( .A(n6190), .B(n6191), .Z(n6189) );
  XOR U5841 ( .A(p_input[3553]), .B(n6188), .Z(n6191) );
  XNOR U5842 ( .A(p_input[3521]), .B(n6188), .Z(n6190) );
  AND U5843 ( .A(p_input[3552]), .B(n6192), .Z(n6188) );
  IV U5844 ( .A(p_input[3520]), .Z(n6192) );
  XNOR U5845 ( .A(p_input[3456]), .B(n6193), .Z(n5786) );
  AND U5846 ( .A(n208), .B(n6194), .Z(n6193) );
  XOR U5847 ( .A(p_input[3488]), .B(p_input[3456]), .Z(n6194) );
  XOR U5848 ( .A(n6195), .B(n6196), .Z(n208) );
  AND U5849 ( .A(n6197), .B(n6198), .Z(n6196) );
  XNOR U5850 ( .A(p_input[3519]), .B(n6195), .Z(n6198) );
  XOR U5851 ( .A(n6195), .B(p_input[3487]), .Z(n6197) );
  XOR U5852 ( .A(n6199), .B(n6200), .Z(n6195) );
  AND U5853 ( .A(n6201), .B(n6202), .Z(n6200) );
  XNOR U5854 ( .A(p_input[3518]), .B(n6199), .Z(n6202) );
  XNOR U5855 ( .A(n6199), .B(n5801), .Z(n6201) );
  IV U5856 ( .A(p_input[3486]), .Z(n5801) );
  XOR U5857 ( .A(n6203), .B(n6204), .Z(n6199) );
  AND U5858 ( .A(n6205), .B(n6206), .Z(n6204) );
  XNOR U5859 ( .A(p_input[3517]), .B(n6203), .Z(n6206) );
  XNOR U5860 ( .A(n6203), .B(n5810), .Z(n6205) );
  IV U5861 ( .A(p_input[3485]), .Z(n5810) );
  XOR U5862 ( .A(n6207), .B(n6208), .Z(n6203) );
  AND U5863 ( .A(n6209), .B(n6210), .Z(n6208) );
  XNOR U5864 ( .A(p_input[3516]), .B(n6207), .Z(n6210) );
  XNOR U5865 ( .A(n6207), .B(n5819), .Z(n6209) );
  IV U5866 ( .A(p_input[3484]), .Z(n5819) );
  XOR U5867 ( .A(n6211), .B(n6212), .Z(n6207) );
  AND U5868 ( .A(n6213), .B(n6214), .Z(n6212) );
  XNOR U5869 ( .A(p_input[3515]), .B(n6211), .Z(n6214) );
  XNOR U5870 ( .A(n6211), .B(n5828), .Z(n6213) );
  IV U5871 ( .A(p_input[3483]), .Z(n5828) );
  XOR U5872 ( .A(n6215), .B(n6216), .Z(n6211) );
  AND U5873 ( .A(n6217), .B(n6218), .Z(n6216) );
  XNOR U5874 ( .A(p_input[3514]), .B(n6215), .Z(n6218) );
  XNOR U5875 ( .A(n6215), .B(n5837), .Z(n6217) );
  IV U5876 ( .A(p_input[3482]), .Z(n5837) );
  XOR U5877 ( .A(n6219), .B(n6220), .Z(n6215) );
  AND U5878 ( .A(n6221), .B(n6222), .Z(n6220) );
  XNOR U5879 ( .A(p_input[3513]), .B(n6219), .Z(n6222) );
  XNOR U5880 ( .A(n6219), .B(n5846), .Z(n6221) );
  IV U5881 ( .A(p_input[3481]), .Z(n5846) );
  XOR U5882 ( .A(n6223), .B(n6224), .Z(n6219) );
  AND U5883 ( .A(n6225), .B(n6226), .Z(n6224) );
  XNOR U5884 ( .A(p_input[3512]), .B(n6223), .Z(n6226) );
  XNOR U5885 ( .A(n6223), .B(n5855), .Z(n6225) );
  IV U5886 ( .A(p_input[3480]), .Z(n5855) );
  XOR U5887 ( .A(n6227), .B(n6228), .Z(n6223) );
  AND U5888 ( .A(n6229), .B(n6230), .Z(n6228) );
  XNOR U5889 ( .A(p_input[3511]), .B(n6227), .Z(n6230) );
  XNOR U5890 ( .A(n6227), .B(n5864), .Z(n6229) );
  IV U5891 ( .A(p_input[3479]), .Z(n5864) );
  XOR U5892 ( .A(n6231), .B(n6232), .Z(n6227) );
  AND U5893 ( .A(n6233), .B(n6234), .Z(n6232) );
  XNOR U5894 ( .A(p_input[3510]), .B(n6231), .Z(n6234) );
  XNOR U5895 ( .A(n6231), .B(n5873), .Z(n6233) );
  IV U5896 ( .A(p_input[3478]), .Z(n5873) );
  XOR U5897 ( .A(n6235), .B(n6236), .Z(n6231) );
  AND U5898 ( .A(n6237), .B(n6238), .Z(n6236) );
  XNOR U5899 ( .A(p_input[3509]), .B(n6235), .Z(n6238) );
  XNOR U5900 ( .A(n6235), .B(n5882), .Z(n6237) );
  IV U5901 ( .A(p_input[3477]), .Z(n5882) );
  XOR U5902 ( .A(n6239), .B(n6240), .Z(n6235) );
  AND U5903 ( .A(n6241), .B(n6242), .Z(n6240) );
  XNOR U5904 ( .A(p_input[3508]), .B(n6239), .Z(n6242) );
  XNOR U5905 ( .A(n6239), .B(n5891), .Z(n6241) );
  IV U5906 ( .A(p_input[3476]), .Z(n5891) );
  XOR U5907 ( .A(n6243), .B(n6244), .Z(n6239) );
  AND U5908 ( .A(n6245), .B(n6246), .Z(n6244) );
  XNOR U5909 ( .A(p_input[3507]), .B(n6243), .Z(n6246) );
  XNOR U5910 ( .A(n6243), .B(n5900), .Z(n6245) );
  IV U5911 ( .A(p_input[3475]), .Z(n5900) );
  XOR U5912 ( .A(n6247), .B(n6248), .Z(n6243) );
  AND U5913 ( .A(n6249), .B(n6250), .Z(n6248) );
  XNOR U5914 ( .A(p_input[3506]), .B(n6247), .Z(n6250) );
  XNOR U5915 ( .A(n6247), .B(n5909), .Z(n6249) );
  IV U5916 ( .A(p_input[3474]), .Z(n5909) );
  XOR U5917 ( .A(n6251), .B(n6252), .Z(n6247) );
  AND U5918 ( .A(n6253), .B(n6254), .Z(n6252) );
  XNOR U5919 ( .A(p_input[3505]), .B(n6251), .Z(n6254) );
  XNOR U5920 ( .A(n6251), .B(n5918), .Z(n6253) );
  IV U5921 ( .A(p_input[3473]), .Z(n5918) );
  XOR U5922 ( .A(n6255), .B(n6256), .Z(n6251) );
  AND U5923 ( .A(n6257), .B(n6258), .Z(n6256) );
  XNOR U5924 ( .A(p_input[3504]), .B(n6255), .Z(n6258) );
  XNOR U5925 ( .A(n6255), .B(n5927), .Z(n6257) );
  IV U5926 ( .A(p_input[3472]), .Z(n5927) );
  XOR U5927 ( .A(n6259), .B(n6260), .Z(n6255) );
  AND U5928 ( .A(n6261), .B(n6262), .Z(n6260) );
  XNOR U5929 ( .A(p_input[3503]), .B(n6259), .Z(n6262) );
  XNOR U5930 ( .A(n6259), .B(n5936), .Z(n6261) );
  IV U5931 ( .A(p_input[3471]), .Z(n5936) );
  XOR U5932 ( .A(n6263), .B(n6264), .Z(n6259) );
  AND U5933 ( .A(n6265), .B(n6266), .Z(n6264) );
  XNOR U5934 ( .A(p_input[3502]), .B(n6263), .Z(n6266) );
  XNOR U5935 ( .A(n6263), .B(n5945), .Z(n6265) );
  IV U5936 ( .A(p_input[3470]), .Z(n5945) );
  XOR U5937 ( .A(n6267), .B(n6268), .Z(n6263) );
  AND U5938 ( .A(n6269), .B(n6270), .Z(n6268) );
  XNOR U5939 ( .A(p_input[3501]), .B(n6267), .Z(n6270) );
  XNOR U5940 ( .A(n6267), .B(n5954), .Z(n6269) );
  IV U5941 ( .A(p_input[3469]), .Z(n5954) );
  XOR U5942 ( .A(n6271), .B(n6272), .Z(n6267) );
  AND U5943 ( .A(n6273), .B(n6274), .Z(n6272) );
  XNOR U5944 ( .A(p_input[3500]), .B(n6271), .Z(n6274) );
  XNOR U5945 ( .A(n6271), .B(n5963), .Z(n6273) );
  IV U5946 ( .A(p_input[3468]), .Z(n5963) );
  XOR U5947 ( .A(n6275), .B(n6276), .Z(n6271) );
  AND U5948 ( .A(n6277), .B(n6278), .Z(n6276) );
  XNOR U5949 ( .A(p_input[3499]), .B(n6275), .Z(n6278) );
  XNOR U5950 ( .A(n6275), .B(n5972), .Z(n6277) );
  IV U5951 ( .A(p_input[3467]), .Z(n5972) );
  XOR U5952 ( .A(n6279), .B(n6280), .Z(n6275) );
  AND U5953 ( .A(n6281), .B(n6282), .Z(n6280) );
  XNOR U5954 ( .A(p_input[3498]), .B(n6279), .Z(n6282) );
  XNOR U5955 ( .A(n6279), .B(n5981), .Z(n6281) );
  IV U5956 ( .A(p_input[3466]), .Z(n5981) );
  XOR U5957 ( .A(n6283), .B(n6284), .Z(n6279) );
  AND U5958 ( .A(n6285), .B(n6286), .Z(n6284) );
  XNOR U5959 ( .A(p_input[3497]), .B(n6283), .Z(n6286) );
  XNOR U5960 ( .A(n6283), .B(n5990), .Z(n6285) );
  IV U5961 ( .A(p_input[3465]), .Z(n5990) );
  XOR U5962 ( .A(n6287), .B(n6288), .Z(n6283) );
  AND U5963 ( .A(n6289), .B(n6290), .Z(n6288) );
  XNOR U5964 ( .A(p_input[3496]), .B(n6287), .Z(n6290) );
  XNOR U5965 ( .A(n6287), .B(n5999), .Z(n6289) );
  IV U5966 ( .A(p_input[3464]), .Z(n5999) );
  XOR U5967 ( .A(n6291), .B(n6292), .Z(n6287) );
  AND U5968 ( .A(n6293), .B(n6294), .Z(n6292) );
  XNOR U5969 ( .A(p_input[3495]), .B(n6291), .Z(n6294) );
  XNOR U5970 ( .A(n6291), .B(n6008), .Z(n6293) );
  IV U5971 ( .A(p_input[3463]), .Z(n6008) );
  XOR U5972 ( .A(n6295), .B(n6296), .Z(n6291) );
  AND U5973 ( .A(n6297), .B(n6298), .Z(n6296) );
  XNOR U5974 ( .A(p_input[3494]), .B(n6295), .Z(n6298) );
  XNOR U5975 ( .A(n6295), .B(n6017), .Z(n6297) );
  IV U5976 ( .A(p_input[3462]), .Z(n6017) );
  XOR U5977 ( .A(n6299), .B(n6300), .Z(n6295) );
  AND U5978 ( .A(n6301), .B(n6302), .Z(n6300) );
  XNOR U5979 ( .A(p_input[3493]), .B(n6299), .Z(n6302) );
  XNOR U5980 ( .A(n6299), .B(n6026), .Z(n6301) );
  IV U5981 ( .A(p_input[3461]), .Z(n6026) );
  XOR U5982 ( .A(n6303), .B(n6304), .Z(n6299) );
  AND U5983 ( .A(n6305), .B(n6306), .Z(n6304) );
  XNOR U5984 ( .A(p_input[3492]), .B(n6303), .Z(n6306) );
  XNOR U5985 ( .A(n6303), .B(n6035), .Z(n6305) );
  IV U5986 ( .A(p_input[3460]), .Z(n6035) );
  XOR U5987 ( .A(n6307), .B(n6308), .Z(n6303) );
  AND U5988 ( .A(n6309), .B(n6310), .Z(n6308) );
  XNOR U5989 ( .A(p_input[3491]), .B(n6307), .Z(n6310) );
  XNOR U5990 ( .A(n6307), .B(n6044), .Z(n6309) );
  IV U5991 ( .A(p_input[3459]), .Z(n6044) );
  XOR U5992 ( .A(n6311), .B(n6312), .Z(n6307) );
  AND U5993 ( .A(n6313), .B(n6314), .Z(n6312) );
  XNOR U5994 ( .A(p_input[3490]), .B(n6311), .Z(n6314) );
  XNOR U5995 ( .A(n6311), .B(n6053), .Z(n6313) );
  IV U5996 ( .A(p_input[3458]), .Z(n6053) );
  XNOR U5997 ( .A(n6315), .B(n6316), .Z(n6311) );
  AND U5998 ( .A(n6317), .B(n6318), .Z(n6316) );
  XOR U5999 ( .A(p_input[3489]), .B(n6315), .Z(n6318) );
  XNOR U6000 ( .A(p_input[3457]), .B(n6315), .Z(n6317) );
  AND U6001 ( .A(p_input[3488]), .B(n6319), .Z(n6315) );
  IV U6002 ( .A(p_input[3456]), .Z(n6319) );
  XOR U6003 ( .A(n6320), .B(n6321), .Z(n5409) );
  AND U6004 ( .A(n316), .B(n6322), .Z(n6321) );
  XNOR U6005 ( .A(n6323), .B(n6320), .Z(n6322) );
  XOR U6006 ( .A(n6324), .B(n6325), .Z(n316) );
  AND U6007 ( .A(n6326), .B(n6327), .Z(n6325) );
  XNOR U6008 ( .A(n5424), .B(n6324), .Z(n6327) );
  AND U6009 ( .A(p_input[3455]), .B(p_input[3423]), .Z(n5424) );
  XNOR U6010 ( .A(n6324), .B(n5421), .Z(n6326) );
  IV U6011 ( .A(n6328), .Z(n5421) );
  AND U6012 ( .A(p_input[3359]), .B(p_input[3391]), .Z(n6328) );
  XOR U6013 ( .A(n6329), .B(n6330), .Z(n6324) );
  AND U6014 ( .A(n6331), .B(n6332), .Z(n6330) );
  XOR U6015 ( .A(n6329), .B(n5436), .Z(n6332) );
  XNOR U6016 ( .A(p_input[3422]), .B(n6333), .Z(n5436) );
  AND U6017 ( .A(n214), .B(n6334), .Z(n6333) );
  XOR U6018 ( .A(p_input[3454]), .B(p_input[3422]), .Z(n6334) );
  XNOR U6019 ( .A(n5433), .B(n6329), .Z(n6331) );
  XOR U6020 ( .A(n6335), .B(n6336), .Z(n5433) );
  AND U6021 ( .A(n211), .B(n6337), .Z(n6336) );
  XOR U6022 ( .A(p_input[3390]), .B(p_input[3358]), .Z(n6337) );
  XOR U6023 ( .A(n6338), .B(n6339), .Z(n6329) );
  AND U6024 ( .A(n6340), .B(n6341), .Z(n6339) );
  XOR U6025 ( .A(n6338), .B(n5448), .Z(n6341) );
  XNOR U6026 ( .A(p_input[3421]), .B(n6342), .Z(n5448) );
  AND U6027 ( .A(n214), .B(n6343), .Z(n6342) );
  XOR U6028 ( .A(p_input[3453]), .B(p_input[3421]), .Z(n6343) );
  XNOR U6029 ( .A(n5445), .B(n6338), .Z(n6340) );
  XOR U6030 ( .A(n6344), .B(n6345), .Z(n5445) );
  AND U6031 ( .A(n211), .B(n6346), .Z(n6345) );
  XOR U6032 ( .A(p_input[3389]), .B(p_input[3357]), .Z(n6346) );
  XOR U6033 ( .A(n6347), .B(n6348), .Z(n6338) );
  AND U6034 ( .A(n6349), .B(n6350), .Z(n6348) );
  XOR U6035 ( .A(n6347), .B(n5460), .Z(n6350) );
  XNOR U6036 ( .A(p_input[3420]), .B(n6351), .Z(n5460) );
  AND U6037 ( .A(n214), .B(n6352), .Z(n6351) );
  XOR U6038 ( .A(p_input[3452]), .B(p_input[3420]), .Z(n6352) );
  XNOR U6039 ( .A(n5457), .B(n6347), .Z(n6349) );
  XOR U6040 ( .A(n6353), .B(n6354), .Z(n5457) );
  AND U6041 ( .A(n211), .B(n6355), .Z(n6354) );
  XOR U6042 ( .A(p_input[3388]), .B(p_input[3356]), .Z(n6355) );
  XOR U6043 ( .A(n6356), .B(n6357), .Z(n6347) );
  AND U6044 ( .A(n6358), .B(n6359), .Z(n6357) );
  XOR U6045 ( .A(n6356), .B(n5472), .Z(n6359) );
  XNOR U6046 ( .A(p_input[3419]), .B(n6360), .Z(n5472) );
  AND U6047 ( .A(n214), .B(n6361), .Z(n6360) );
  XOR U6048 ( .A(p_input[3451]), .B(p_input[3419]), .Z(n6361) );
  XNOR U6049 ( .A(n5469), .B(n6356), .Z(n6358) );
  XOR U6050 ( .A(n6362), .B(n6363), .Z(n5469) );
  AND U6051 ( .A(n211), .B(n6364), .Z(n6363) );
  XOR U6052 ( .A(p_input[3387]), .B(p_input[3355]), .Z(n6364) );
  XOR U6053 ( .A(n6365), .B(n6366), .Z(n6356) );
  AND U6054 ( .A(n6367), .B(n6368), .Z(n6366) );
  XOR U6055 ( .A(n6365), .B(n5484), .Z(n6368) );
  XNOR U6056 ( .A(p_input[3418]), .B(n6369), .Z(n5484) );
  AND U6057 ( .A(n214), .B(n6370), .Z(n6369) );
  XOR U6058 ( .A(p_input[3450]), .B(p_input[3418]), .Z(n6370) );
  XNOR U6059 ( .A(n5481), .B(n6365), .Z(n6367) );
  XOR U6060 ( .A(n6371), .B(n6372), .Z(n5481) );
  AND U6061 ( .A(n211), .B(n6373), .Z(n6372) );
  XOR U6062 ( .A(p_input[3386]), .B(p_input[3354]), .Z(n6373) );
  XOR U6063 ( .A(n6374), .B(n6375), .Z(n6365) );
  AND U6064 ( .A(n6376), .B(n6377), .Z(n6375) );
  XOR U6065 ( .A(n6374), .B(n5496), .Z(n6377) );
  XNOR U6066 ( .A(p_input[3417]), .B(n6378), .Z(n5496) );
  AND U6067 ( .A(n214), .B(n6379), .Z(n6378) );
  XOR U6068 ( .A(p_input[3449]), .B(p_input[3417]), .Z(n6379) );
  XNOR U6069 ( .A(n5493), .B(n6374), .Z(n6376) );
  XOR U6070 ( .A(n6380), .B(n6381), .Z(n5493) );
  AND U6071 ( .A(n211), .B(n6382), .Z(n6381) );
  XOR U6072 ( .A(p_input[3385]), .B(p_input[3353]), .Z(n6382) );
  XOR U6073 ( .A(n6383), .B(n6384), .Z(n6374) );
  AND U6074 ( .A(n6385), .B(n6386), .Z(n6384) );
  XOR U6075 ( .A(n6383), .B(n5508), .Z(n6386) );
  XNOR U6076 ( .A(p_input[3416]), .B(n6387), .Z(n5508) );
  AND U6077 ( .A(n214), .B(n6388), .Z(n6387) );
  XOR U6078 ( .A(p_input[3448]), .B(p_input[3416]), .Z(n6388) );
  XNOR U6079 ( .A(n5505), .B(n6383), .Z(n6385) );
  XOR U6080 ( .A(n6389), .B(n6390), .Z(n5505) );
  AND U6081 ( .A(n211), .B(n6391), .Z(n6390) );
  XOR U6082 ( .A(p_input[3384]), .B(p_input[3352]), .Z(n6391) );
  XOR U6083 ( .A(n6392), .B(n6393), .Z(n6383) );
  AND U6084 ( .A(n6394), .B(n6395), .Z(n6393) );
  XOR U6085 ( .A(n6392), .B(n5520), .Z(n6395) );
  XNOR U6086 ( .A(p_input[3415]), .B(n6396), .Z(n5520) );
  AND U6087 ( .A(n214), .B(n6397), .Z(n6396) );
  XOR U6088 ( .A(p_input[3447]), .B(p_input[3415]), .Z(n6397) );
  XNOR U6089 ( .A(n5517), .B(n6392), .Z(n6394) );
  XOR U6090 ( .A(n6398), .B(n6399), .Z(n5517) );
  AND U6091 ( .A(n211), .B(n6400), .Z(n6399) );
  XOR U6092 ( .A(p_input[3383]), .B(p_input[3351]), .Z(n6400) );
  XOR U6093 ( .A(n6401), .B(n6402), .Z(n6392) );
  AND U6094 ( .A(n6403), .B(n6404), .Z(n6402) );
  XOR U6095 ( .A(n6401), .B(n5532), .Z(n6404) );
  XNOR U6096 ( .A(p_input[3414]), .B(n6405), .Z(n5532) );
  AND U6097 ( .A(n214), .B(n6406), .Z(n6405) );
  XOR U6098 ( .A(p_input[3446]), .B(p_input[3414]), .Z(n6406) );
  XNOR U6099 ( .A(n5529), .B(n6401), .Z(n6403) );
  XOR U6100 ( .A(n6407), .B(n6408), .Z(n5529) );
  AND U6101 ( .A(n211), .B(n6409), .Z(n6408) );
  XOR U6102 ( .A(p_input[3382]), .B(p_input[3350]), .Z(n6409) );
  XOR U6103 ( .A(n6410), .B(n6411), .Z(n6401) );
  AND U6104 ( .A(n6412), .B(n6413), .Z(n6411) );
  XOR U6105 ( .A(n6410), .B(n5544), .Z(n6413) );
  XNOR U6106 ( .A(p_input[3413]), .B(n6414), .Z(n5544) );
  AND U6107 ( .A(n214), .B(n6415), .Z(n6414) );
  XOR U6108 ( .A(p_input[3445]), .B(p_input[3413]), .Z(n6415) );
  XNOR U6109 ( .A(n5541), .B(n6410), .Z(n6412) );
  XOR U6110 ( .A(n6416), .B(n6417), .Z(n5541) );
  AND U6111 ( .A(n211), .B(n6418), .Z(n6417) );
  XOR U6112 ( .A(p_input[3381]), .B(p_input[3349]), .Z(n6418) );
  XOR U6113 ( .A(n6419), .B(n6420), .Z(n6410) );
  AND U6114 ( .A(n6421), .B(n6422), .Z(n6420) );
  XOR U6115 ( .A(n6419), .B(n5556), .Z(n6422) );
  XNOR U6116 ( .A(p_input[3412]), .B(n6423), .Z(n5556) );
  AND U6117 ( .A(n214), .B(n6424), .Z(n6423) );
  XOR U6118 ( .A(p_input[3444]), .B(p_input[3412]), .Z(n6424) );
  XNOR U6119 ( .A(n5553), .B(n6419), .Z(n6421) );
  XOR U6120 ( .A(n6425), .B(n6426), .Z(n5553) );
  AND U6121 ( .A(n211), .B(n6427), .Z(n6426) );
  XOR U6122 ( .A(p_input[3380]), .B(p_input[3348]), .Z(n6427) );
  XOR U6123 ( .A(n6428), .B(n6429), .Z(n6419) );
  AND U6124 ( .A(n6430), .B(n6431), .Z(n6429) );
  XOR U6125 ( .A(n6428), .B(n5568), .Z(n6431) );
  XNOR U6126 ( .A(p_input[3411]), .B(n6432), .Z(n5568) );
  AND U6127 ( .A(n214), .B(n6433), .Z(n6432) );
  XOR U6128 ( .A(p_input[3443]), .B(p_input[3411]), .Z(n6433) );
  XNOR U6129 ( .A(n5565), .B(n6428), .Z(n6430) );
  XOR U6130 ( .A(n6434), .B(n6435), .Z(n5565) );
  AND U6131 ( .A(n211), .B(n6436), .Z(n6435) );
  XOR U6132 ( .A(p_input[3379]), .B(p_input[3347]), .Z(n6436) );
  XOR U6133 ( .A(n6437), .B(n6438), .Z(n6428) );
  AND U6134 ( .A(n6439), .B(n6440), .Z(n6438) );
  XOR U6135 ( .A(n6437), .B(n5580), .Z(n6440) );
  XNOR U6136 ( .A(p_input[3410]), .B(n6441), .Z(n5580) );
  AND U6137 ( .A(n214), .B(n6442), .Z(n6441) );
  XOR U6138 ( .A(p_input[3442]), .B(p_input[3410]), .Z(n6442) );
  XNOR U6139 ( .A(n5577), .B(n6437), .Z(n6439) );
  XOR U6140 ( .A(n6443), .B(n6444), .Z(n5577) );
  AND U6141 ( .A(n211), .B(n6445), .Z(n6444) );
  XOR U6142 ( .A(p_input[3378]), .B(p_input[3346]), .Z(n6445) );
  XOR U6143 ( .A(n6446), .B(n6447), .Z(n6437) );
  AND U6144 ( .A(n6448), .B(n6449), .Z(n6447) );
  XOR U6145 ( .A(n6446), .B(n5592), .Z(n6449) );
  XNOR U6146 ( .A(p_input[3409]), .B(n6450), .Z(n5592) );
  AND U6147 ( .A(n214), .B(n6451), .Z(n6450) );
  XOR U6148 ( .A(p_input[3441]), .B(p_input[3409]), .Z(n6451) );
  XNOR U6149 ( .A(n5589), .B(n6446), .Z(n6448) );
  XOR U6150 ( .A(n6452), .B(n6453), .Z(n5589) );
  AND U6151 ( .A(n211), .B(n6454), .Z(n6453) );
  XOR U6152 ( .A(p_input[3377]), .B(p_input[3345]), .Z(n6454) );
  XOR U6153 ( .A(n6455), .B(n6456), .Z(n6446) );
  AND U6154 ( .A(n6457), .B(n6458), .Z(n6456) );
  XOR U6155 ( .A(n6455), .B(n5604), .Z(n6458) );
  XNOR U6156 ( .A(p_input[3408]), .B(n6459), .Z(n5604) );
  AND U6157 ( .A(n214), .B(n6460), .Z(n6459) );
  XOR U6158 ( .A(p_input[3440]), .B(p_input[3408]), .Z(n6460) );
  XNOR U6159 ( .A(n5601), .B(n6455), .Z(n6457) );
  XOR U6160 ( .A(n6461), .B(n6462), .Z(n5601) );
  AND U6161 ( .A(n211), .B(n6463), .Z(n6462) );
  XOR U6162 ( .A(p_input[3376]), .B(p_input[3344]), .Z(n6463) );
  XOR U6163 ( .A(n6464), .B(n6465), .Z(n6455) );
  AND U6164 ( .A(n6466), .B(n6467), .Z(n6465) );
  XOR U6165 ( .A(n6464), .B(n5616), .Z(n6467) );
  XNOR U6166 ( .A(p_input[3407]), .B(n6468), .Z(n5616) );
  AND U6167 ( .A(n214), .B(n6469), .Z(n6468) );
  XOR U6168 ( .A(p_input[3439]), .B(p_input[3407]), .Z(n6469) );
  XNOR U6169 ( .A(n5613), .B(n6464), .Z(n6466) );
  XOR U6170 ( .A(n6470), .B(n6471), .Z(n5613) );
  AND U6171 ( .A(n211), .B(n6472), .Z(n6471) );
  XOR U6172 ( .A(p_input[3375]), .B(p_input[3343]), .Z(n6472) );
  XOR U6173 ( .A(n6473), .B(n6474), .Z(n6464) );
  AND U6174 ( .A(n6475), .B(n6476), .Z(n6474) );
  XOR U6175 ( .A(n6473), .B(n5628), .Z(n6476) );
  XNOR U6176 ( .A(p_input[3406]), .B(n6477), .Z(n5628) );
  AND U6177 ( .A(n214), .B(n6478), .Z(n6477) );
  XOR U6178 ( .A(p_input[3438]), .B(p_input[3406]), .Z(n6478) );
  XNOR U6179 ( .A(n5625), .B(n6473), .Z(n6475) );
  XOR U6180 ( .A(n6479), .B(n6480), .Z(n5625) );
  AND U6181 ( .A(n211), .B(n6481), .Z(n6480) );
  XOR U6182 ( .A(p_input[3374]), .B(p_input[3342]), .Z(n6481) );
  XOR U6183 ( .A(n6482), .B(n6483), .Z(n6473) );
  AND U6184 ( .A(n6484), .B(n6485), .Z(n6483) );
  XOR U6185 ( .A(n6482), .B(n5640), .Z(n6485) );
  XNOR U6186 ( .A(p_input[3405]), .B(n6486), .Z(n5640) );
  AND U6187 ( .A(n214), .B(n6487), .Z(n6486) );
  XOR U6188 ( .A(p_input[3437]), .B(p_input[3405]), .Z(n6487) );
  XNOR U6189 ( .A(n5637), .B(n6482), .Z(n6484) );
  XOR U6190 ( .A(n6488), .B(n6489), .Z(n5637) );
  AND U6191 ( .A(n211), .B(n6490), .Z(n6489) );
  XOR U6192 ( .A(p_input[3373]), .B(p_input[3341]), .Z(n6490) );
  XOR U6193 ( .A(n6491), .B(n6492), .Z(n6482) );
  AND U6194 ( .A(n6493), .B(n6494), .Z(n6492) );
  XOR U6195 ( .A(n6491), .B(n5652), .Z(n6494) );
  XNOR U6196 ( .A(p_input[3404]), .B(n6495), .Z(n5652) );
  AND U6197 ( .A(n214), .B(n6496), .Z(n6495) );
  XOR U6198 ( .A(p_input[3436]), .B(p_input[3404]), .Z(n6496) );
  XNOR U6199 ( .A(n5649), .B(n6491), .Z(n6493) );
  XOR U6200 ( .A(n6497), .B(n6498), .Z(n5649) );
  AND U6201 ( .A(n211), .B(n6499), .Z(n6498) );
  XOR U6202 ( .A(p_input[3372]), .B(p_input[3340]), .Z(n6499) );
  XOR U6203 ( .A(n6500), .B(n6501), .Z(n6491) );
  AND U6204 ( .A(n6502), .B(n6503), .Z(n6501) );
  XOR U6205 ( .A(n6500), .B(n5664), .Z(n6503) );
  XNOR U6206 ( .A(p_input[3403]), .B(n6504), .Z(n5664) );
  AND U6207 ( .A(n214), .B(n6505), .Z(n6504) );
  XOR U6208 ( .A(p_input[3435]), .B(p_input[3403]), .Z(n6505) );
  XNOR U6209 ( .A(n5661), .B(n6500), .Z(n6502) );
  XOR U6210 ( .A(n6506), .B(n6507), .Z(n5661) );
  AND U6211 ( .A(n211), .B(n6508), .Z(n6507) );
  XOR U6212 ( .A(p_input[3371]), .B(p_input[3339]), .Z(n6508) );
  XOR U6213 ( .A(n6509), .B(n6510), .Z(n6500) );
  AND U6214 ( .A(n6511), .B(n6512), .Z(n6510) );
  XOR U6215 ( .A(n6509), .B(n5676), .Z(n6512) );
  XNOR U6216 ( .A(p_input[3402]), .B(n6513), .Z(n5676) );
  AND U6217 ( .A(n214), .B(n6514), .Z(n6513) );
  XOR U6218 ( .A(p_input[3434]), .B(p_input[3402]), .Z(n6514) );
  XNOR U6219 ( .A(n5673), .B(n6509), .Z(n6511) );
  XOR U6220 ( .A(n6515), .B(n6516), .Z(n5673) );
  AND U6221 ( .A(n211), .B(n6517), .Z(n6516) );
  XOR U6222 ( .A(p_input[3370]), .B(p_input[3338]), .Z(n6517) );
  XOR U6223 ( .A(n6518), .B(n6519), .Z(n6509) );
  AND U6224 ( .A(n6520), .B(n6521), .Z(n6519) );
  XOR U6225 ( .A(n6518), .B(n5688), .Z(n6521) );
  XNOR U6226 ( .A(p_input[3401]), .B(n6522), .Z(n5688) );
  AND U6227 ( .A(n214), .B(n6523), .Z(n6522) );
  XOR U6228 ( .A(p_input[3433]), .B(p_input[3401]), .Z(n6523) );
  XNOR U6229 ( .A(n5685), .B(n6518), .Z(n6520) );
  XOR U6230 ( .A(n6524), .B(n6525), .Z(n5685) );
  AND U6231 ( .A(n211), .B(n6526), .Z(n6525) );
  XOR U6232 ( .A(p_input[3369]), .B(p_input[3337]), .Z(n6526) );
  XOR U6233 ( .A(n6527), .B(n6528), .Z(n6518) );
  AND U6234 ( .A(n6529), .B(n6530), .Z(n6528) );
  XOR U6235 ( .A(n6527), .B(n5700), .Z(n6530) );
  XNOR U6236 ( .A(p_input[3400]), .B(n6531), .Z(n5700) );
  AND U6237 ( .A(n214), .B(n6532), .Z(n6531) );
  XOR U6238 ( .A(p_input[3432]), .B(p_input[3400]), .Z(n6532) );
  XNOR U6239 ( .A(n5697), .B(n6527), .Z(n6529) );
  XOR U6240 ( .A(n6533), .B(n6534), .Z(n5697) );
  AND U6241 ( .A(n211), .B(n6535), .Z(n6534) );
  XOR U6242 ( .A(p_input[3368]), .B(p_input[3336]), .Z(n6535) );
  XOR U6243 ( .A(n6536), .B(n6537), .Z(n6527) );
  AND U6244 ( .A(n6538), .B(n6539), .Z(n6537) );
  XOR U6245 ( .A(n6536), .B(n5712), .Z(n6539) );
  XNOR U6246 ( .A(p_input[3399]), .B(n6540), .Z(n5712) );
  AND U6247 ( .A(n214), .B(n6541), .Z(n6540) );
  XOR U6248 ( .A(p_input[3431]), .B(p_input[3399]), .Z(n6541) );
  XNOR U6249 ( .A(n5709), .B(n6536), .Z(n6538) );
  XOR U6250 ( .A(n6542), .B(n6543), .Z(n5709) );
  AND U6251 ( .A(n211), .B(n6544), .Z(n6543) );
  XOR U6252 ( .A(p_input[3367]), .B(p_input[3335]), .Z(n6544) );
  XOR U6253 ( .A(n6545), .B(n6546), .Z(n6536) );
  AND U6254 ( .A(n6547), .B(n6548), .Z(n6546) );
  XOR U6255 ( .A(n6545), .B(n5724), .Z(n6548) );
  XNOR U6256 ( .A(p_input[3398]), .B(n6549), .Z(n5724) );
  AND U6257 ( .A(n214), .B(n6550), .Z(n6549) );
  XOR U6258 ( .A(p_input[3430]), .B(p_input[3398]), .Z(n6550) );
  XNOR U6259 ( .A(n5721), .B(n6545), .Z(n6547) );
  XOR U6260 ( .A(n6551), .B(n6552), .Z(n5721) );
  AND U6261 ( .A(n211), .B(n6553), .Z(n6552) );
  XOR U6262 ( .A(p_input[3366]), .B(p_input[3334]), .Z(n6553) );
  XOR U6263 ( .A(n6554), .B(n6555), .Z(n6545) );
  AND U6264 ( .A(n6556), .B(n6557), .Z(n6555) );
  XOR U6265 ( .A(n6554), .B(n5736), .Z(n6557) );
  XNOR U6266 ( .A(p_input[3397]), .B(n6558), .Z(n5736) );
  AND U6267 ( .A(n214), .B(n6559), .Z(n6558) );
  XOR U6268 ( .A(p_input[3429]), .B(p_input[3397]), .Z(n6559) );
  XNOR U6269 ( .A(n5733), .B(n6554), .Z(n6556) );
  XOR U6270 ( .A(n6560), .B(n6561), .Z(n5733) );
  AND U6271 ( .A(n211), .B(n6562), .Z(n6561) );
  XOR U6272 ( .A(p_input[3365]), .B(p_input[3333]), .Z(n6562) );
  XOR U6273 ( .A(n6563), .B(n6564), .Z(n6554) );
  AND U6274 ( .A(n6565), .B(n6566), .Z(n6564) );
  XOR U6275 ( .A(n6563), .B(n5748), .Z(n6566) );
  XNOR U6276 ( .A(p_input[3396]), .B(n6567), .Z(n5748) );
  AND U6277 ( .A(n214), .B(n6568), .Z(n6567) );
  XOR U6278 ( .A(p_input[3428]), .B(p_input[3396]), .Z(n6568) );
  XNOR U6279 ( .A(n5745), .B(n6563), .Z(n6565) );
  XOR U6280 ( .A(n6569), .B(n6570), .Z(n5745) );
  AND U6281 ( .A(n211), .B(n6571), .Z(n6570) );
  XOR U6282 ( .A(p_input[3364]), .B(p_input[3332]), .Z(n6571) );
  XOR U6283 ( .A(n6572), .B(n6573), .Z(n6563) );
  AND U6284 ( .A(n6574), .B(n6575), .Z(n6573) );
  XOR U6285 ( .A(n6572), .B(n5760), .Z(n6575) );
  XNOR U6286 ( .A(p_input[3395]), .B(n6576), .Z(n5760) );
  AND U6287 ( .A(n214), .B(n6577), .Z(n6576) );
  XOR U6288 ( .A(p_input[3427]), .B(p_input[3395]), .Z(n6577) );
  XNOR U6289 ( .A(n5757), .B(n6572), .Z(n6574) );
  XOR U6290 ( .A(n6578), .B(n6579), .Z(n5757) );
  AND U6291 ( .A(n211), .B(n6580), .Z(n6579) );
  XOR U6292 ( .A(p_input[3363]), .B(p_input[3331]), .Z(n6580) );
  XOR U6293 ( .A(n6581), .B(n6582), .Z(n6572) );
  AND U6294 ( .A(n6583), .B(n6584), .Z(n6582) );
  XOR U6295 ( .A(n5772), .B(n6581), .Z(n6584) );
  XNOR U6296 ( .A(p_input[3394]), .B(n6585), .Z(n5772) );
  AND U6297 ( .A(n214), .B(n6586), .Z(n6585) );
  XOR U6298 ( .A(p_input[3426]), .B(p_input[3394]), .Z(n6586) );
  XNOR U6299 ( .A(n6581), .B(n5769), .Z(n6583) );
  XOR U6300 ( .A(n6587), .B(n6588), .Z(n5769) );
  AND U6301 ( .A(n211), .B(n6589), .Z(n6588) );
  XOR U6302 ( .A(p_input[3362]), .B(p_input[3330]), .Z(n6589) );
  XOR U6303 ( .A(n6590), .B(n6591), .Z(n6581) );
  AND U6304 ( .A(n6592), .B(n6593), .Z(n6591) );
  XNOR U6305 ( .A(n6594), .B(n5785), .Z(n6593) );
  XNOR U6306 ( .A(p_input[3393]), .B(n6595), .Z(n5785) );
  AND U6307 ( .A(n214), .B(n6596), .Z(n6595) );
  XNOR U6308 ( .A(p_input[3425]), .B(n6597), .Z(n6596) );
  IV U6309 ( .A(p_input[3393]), .Z(n6597) );
  XNOR U6310 ( .A(n5782), .B(n6590), .Z(n6592) );
  XNOR U6311 ( .A(p_input[3329]), .B(n6598), .Z(n5782) );
  AND U6312 ( .A(n211), .B(n6599), .Z(n6598) );
  XOR U6313 ( .A(p_input[3361]), .B(p_input[3329]), .Z(n6599) );
  IV U6314 ( .A(n6594), .Z(n6590) );
  AND U6315 ( .A(n6320), .B(n6323), .Z(n6594) );
  XOR U6316 ( .A(p_input[3392]), .B(n6600), .Z(n6323) );
  AND U6317 ( .A(n214), .B(n6601), .Z(n6600) );
  XOR U6318 ( .A(p_input[3424]), .B(p_input[3392]), .Z(n6601) );
  XOR U6319 ( .A(n6602), .B(n6603), .Z(n214) );
  AND U6320 ( .A(n6604), .B(n6605), .Z(n6603) );
  XNOR U6321 ( .A(p_input[3455]), .B(n6602), .Z(n6605) );
  XOR U6322 ( .A(n6602), .B(p_input[3423]), .Z(n6604) );
  XOR U6323 ( .A(n6606), .B(n6607), .Z(n6602) );
  AND U6324 ( .A(n6608), .B(n6609), .Z(n6607) );
  XNOR U6325 ( .A(p_input[3454]), .B(n6606), .Z(n6609) );
  XOR U6326 ( .A(n6606), .B(p_input[3422]), .Z(n6608) );
  XOR U6327 ( .A(n6610), .B(n6611), .Z(n6606) );
  AND U6328 ( .A(n6612), .B(n6613), .Z(n6611) );
  XNOR U6329 ( .A(p_input[3453]), .B(n6610), .Z(n6613) );
  XOR U6330 ( .A(n6610), .B(p_input[3421]), .Z(n6612) );
  XOR U6331 ( .A(n6614), .B(n6615), .Z(n6610) );
  AND U6332 ( .A(n6616), .B(n6617), .Z(n6615) );
  XNOR U6333 ( .A(p_input[3452]), .B(n6614), .Z(n6617) );
  XOR U6334 ( .A(n6614), .B(p_input[3420]), .Z(n6616) );
  XOR U6335 ( .A(n6618), .B(n6619), .Z(n6614) );
  AND U6336 ( .A(n6620), .B(n6621), .Z(n6619) );
  XNOR U6337 ( .A(p_input[3451]), .B(n6618), .Z(n6621) );
  XOR U6338 ( .A(n6618), .B(p_input[3419]), .Z(n6620) );
  XOR U6339 ( .A(n6622), .B(n6623), .Z(n6618) );
  AND U6340 ( .A(n6624), .B(n6625), .Z(n6623) );
  XNOR U6341 ( .A(p_input[3450]), .B(n6622), .Z(n6625) );
  XOR U6342 ( .A(n6622), .B(p_input[3418]), .Z(n6624) );
  XOR U6343 ( .A(n6626), .B(n6627), .Z(n6622) );
  AND U6344 ( .A(n6628), .B(n6629), .Z(n6627) );
  XNOR U6345 ( .A(p_input[3449]), .B(n6626), .Z(n6629) );
  XOR U6346 ( .A(n6626), .B(p_input[3417]), .Z(n6628) );
  XOR U6347 ( .A(n6630), .B(n6631), .Z(n6626) );
  AND U6348 ( .A(n6632), .B(n6633), .Z(n6631) );
  XNOR U6349 ( .A(p_input[3448]), .B(n6630), .Z(n6633) );
  XOR U6350 ( .A(n6630), .B(p_input[3416]), .Z(n6632) );
  XOR U6351 ( .A(n6634), .B(n6635), .Z(n6630) );
  AND U6352 ( .A(n6636), .B(n6637), .Z(n6635) );
  XNOR U6353 ( .A(p_input[3447]), .B(n6634), .Z(n6637) );
  XOR U6354 ( .A(n6634), .B(p_input[3415]), .Z(n6636) );
  XOR U6355 ( .A(n6638), .B(n6639), .Z(n6634) );
  AND U6356 ( .A(n6640), .B(n6641), .Z(n6639) );
  XNOR U6357 ( .A(p_input[3446]), .B(n6638), .Z(n6641) );
  XOR U6358 ( .A(n6638), .B(p_input[3414]), .Z(n6640) );
  XOR U6359 ( .A(n6642), .B(n6643), .Z(n6638) );
  AND U6360 ( .A(n6644), .B(n6645), .Z(n6643) );
  XNOR U6361 ( .A(p_input[3445]), .B(n6642), .Z(n6645) );
  XOR U6362 ( .A(n6642), .B(p_input[3413]), .Z(n6644) );
  XOR U6363 ( .A(n6646), .B(n6647), .Z(n6642) );
  AND U6364 ( .A(n6648), .B(n6649), .Z(n6647) );
  XNOR U6365 ( .A(p_input[3444]), .B(n6646), .Z(n6649) );
  XOR U6366 ( .A(n6646), .B(p_input[3412]), .Z(n6648) );
  XOR U6367 ( .A(n6650), .B(n6651), .Z(n6646) );
  AND U6368 ( .A(n6652), .B(n6653), .Z(n6651) );
  XNOR U6369 ( .A(p_input[3443]), .B(n6650), .Z(n6653) );
  XOR U6370 ( .A(n6650), .B(p_input[3411]), .Z(n6652) );
  XOR U6371 ( .A(n6654), .B(n6655), .Z(n6650) );
  AND U6372 ( .A(n6656), .B(n6657), .Z(n6655) );
  XNOR U6373 ( .A(p_input[3442]), .B(n6654), .Z(n6657) );
  XOR U6374 ( .A(n6654), .B(p_input[3410]), .Z(n6656) );
  XOR U6375 ( .A(n6658), .B(n6659), .Z(n6654) );
  AND U6376 ( .A(n6660), .B(n6661), .Z(n6659) );
  XNOR U6377 ( .A(p_input[3441]), .B(n6658), .Z(n6661) );
  XOR U6378 ( .A(n6658), .B(p_input[3409]), .Z(n6660) );
  XOR U6379 ( .A(n6662), .B(n6663), .Z(n6658) );
  AND U6380 ( .A(n6664), .B(n6665), .Z(n6663) );
  XNOR U6381 ( .A(p_input[3440]), .B(n6662), .Z(n6665) );
  XOR U6382 ( .A(n6662), .B(p_input[3408]), .Z(n6664) );
  XOR U6383 ( .A(n6666), .B(n6667), .Z(n6662) );
  AND U6384 ( .A(n6668), .B(n6669), .Z(n6667) );
  XNOR U6385 ( .A(p_input[3439]), .B(n6666), .Z(n6669) );
  XOR U6386 ( .A(n6666), .B(p_input[3407]), .Z(n6668) );
  XOR U6387 ( .A(n6670), .B(n6671), .Z(n6666) );
  AND U6388 ( .A(n6672), .B(n6673), .Z(n6671) );
  XNOR U6389 ( .A(p_input[3438]), .B(n6670), .Z(n6673) );
  XOR U6390 ( .A(n6670), .B(p_input[3406]), .Z(n6672) );
  XOR U6391 ( .A(n6674), .B(n6675), .Z(n6670) );
  AND U6392 ( .A(n6676), .B(n6677), .Z(n6675) );
  XNOR U6393 ( .A(p_input[3437]), .B(n6674), .Z(n6677) );
  XOR U6394 ( .A(n6674), .B(p_input[3405]), .Z(n6676) );
  XOR U6395 ( .A(n6678), .B(n6679), .Z(n6674) );
  AND U6396 ( .A(n6680), .B(n6681), .Z(n6679) );
  XNOR U6397 ( .A(p_input[3436]), .B(n6678), .Z(n6681) );
  XOR U6398 ( .A(n6678), .B(p_input[3404]), .Z(n6680) );
  XOR U6399 ( .A(n6682), .B(n6683), .Z(n6678) );
  AND U6400 ( .A(n6684), .B(n6685), .Z(n6683) );
  XNOR U6401 ( .A(p_input[3435]), .B(n6682), .Z(n6685) );
  XOR U6402 ( .A(n6682), .B(p_input[3403]), .Z(n6684) );
  XOR U6403 ( .A(n6686), .B(n6687), .Z(n6682) );
  AND U6404 ( .A(n6688), .B(n6689), .Z(n6687) );
  XNOR U6405 ( .A(p_input[3434]), .B(n6686), .Z(n6689) );
  XOR U6406 ( .A(n6686), .B(p_input[3402]), .Z(n6688) );
  XOR U6407 ( .A(n6690), .B(n6691), .Z(n6686) );
  AND U6408 ( .A(n6692), .B(n6693), .Z(n6691) );
  XNOR U6409 ( .A(p_input[3433]), .B(n6690), .Z(n6693) );
  XOR U6410 ( .A(n6690), .B(p_input[3401]), .Z(n6692) );
  XOR U6411 ( .A(n6694), .B(n6695), .Z(n6690) );
  AND U6412 ( .A(n6696), .B(n6697), .Z(n6695) );
  XNOR U6413 ( .A(p_input[3432]), .B(n6694), .Z(n6697) );
  XOR U6414 ( .A(n6694), .B(p_input[3400]), .Z(n6696) );
  XOR U6415 ( .A(n6698), .B(n6699), .Z(n6694) );
  AND U6416 ( .A(n6700), .B(n6701), .Z(n6699) );
  XNOR U6417 ( .A(p_input[3431]), .B(n6698), .Z(n6701) );
  XOR U6418 ( .A(n6698), .B(p_input[3399]), .Z(n6700) );
  XOR U6419 ( .A(n6702), .B(n6703), .Z(n6698) );
  AND U6420 ( .A(n6704), .B(n6705), .Z(n6703) );
  XNOR U6421 ( .A(p_input[3430]), .B(n6702), .Z(n6705) );
  XOR U6422 ( .A(n6702), .B(p_input[3398]), .Z(n6704) );
  XOR U6423 ( .A(n6706), .B(n6707), .Z(n6702) );
  AND U6424 ( .A(n6708), .B(n6709), .Z(n6707) );
  XNOR U6425 ( .A(p_input[3429]), .B(n6706), .Z(n6709) );
  XOR U6426 ( .A(n6706), .B(p_input[3397]), .Z(n6708) );
  XOR U6427 ( .A(n6710), .B(n6711), .Z(n6706) );
  AND U6428 ( .A(n6712), .B(n6713), .Z(n6711) );
  XNOR U6429 ( .A(p_input[3428]), .B(n6710), .Z(n6713) );
  XOR U6430 ( .A(n6710), .B(p_input[3396]), .Z(n6712) );
  XOR U6431 ( .A(n6714), .B(n6715), .Z(n6710) );
  AND U6432 ( .A(n6716), .B(n6717), .Z(n6715) );
  XNOR U6433 ( .A(p_input[3427]), .B(n6714), .Z(n6717) );
  XOR U6434 ( .A(n6714), .B(p_input[3395]), .Z(n6716) );
  XOR U6435 ( .A(n6718), .B(n6719), .Z(n6714) );
  AND U6436 ( .A(n6720), .B(n6721), .Z(n6719) );
  XNOR U6437 ( .A(p_input[3426]), .B(n6718), .Z(n6721) );
  XOR U6438 ( .A(n6718), .B(p_input[3394]), .Z(n6720) );
  XNOR U6439 ( .A(n6722), .B(n6723), .Z(n6718) );
  AND U6440 ( .A(n6724), .B(n6725), .Z(n6723) );
  XOR U6441 ( .A(p_input[3425]), .B(n6722), .Z(n6725) );
  XNOR U6442 ( .A(p_input[3393]), .B(n6722), .Z(n6724) );
  AND U6443 ( .A(p_input[3424]), .B(n6726), .Z(n6722) );
  IV U6444 ( .A(p_input[3392]), .Z(n6726) );
  XNOR U6445 ( .A(p_input[3328]), .B(n6727), .Z(n6320) );
  AND U6446 ( .A(n211), .B(n6728), .Z(n6727) );
  XOR U6447 ( .A(p_input[3360]), .B(p_input[3328]), .Z(n6728) );
  XOR U6448 ( .A(n6729), .B(n6730), .Z(n211) );
  AND U6449 ( .A(n6731), .B(n6732), .Z(n6730) );
  XNOR U6450 ( .A(p_input[3391]), .B(n6729), .Z(n6732) );
  XOR U6451 ( .A(n6729), .B(p_input[3359]), .Z(n6731) );
  XOR U6452 ( .A(n6733), .B(n6734), .Z(n6729) );
  AND U6453 ( .A(n6735), .B(n6736), .Z(n6734) );
  XNOR U6454 ( .A(p_input[3390]), .B(n6733), .Z(n6736) );
  XNOR U6455 ( .A(n6733), .B(n6335), .Z(n6735) );
  IV U6456 ( .A(p_input[3358]), .Z(n6335) );
  XOR U6457 ( .A(n6737), .B(n6738), .Z(n6733) );
  AND U6458 ( .A(n6739), .B(n6740), .Z(n6738) );
  XNOR U6459 ( .A(p_input[3389]), .B(n6737), .Z(n6740) );
  XNOR U6460 ( .A(n6737), .B(n6344), .Z(n6739) );
  IV U6461 ( .A(p_input[3357]), .Z(n6344) );
  XOR U6462 ( .A(n6741), .B(n6742), .Z(n6737) );
  AND U6463 ( .A(n6743), .B(n6744), .Z(n6742) );
  XNOR U6464 ( .A(p_input[3388]), .B(n6741), .Z(n6744) );
  XNOR U6465 ( .A(n6741), .B(n6353), .Z(n6743) );
  IV U6466 ( .A(p_input[3356]), .Z(n6353) );
  XOR U6467 ( .A(n6745), .B(n6746), .Z(n6741) );
  AND U6468 ( .A(n6747), .B(n6748), .Z(n6746) );
  XNOR U6469 ( .A(p_input[3387]), .B(n6745), .Z(n6748) );
  XNOR U6470 ( .A(n6745), .B(n6362), .Z(n6747) );
  IV U6471 ( .A(p_input[3355]), .Z(n6362) );
  XOR U6472 ( .A(n6749), .B(n6750), .Z(n6745) );
  AND U6473 ( .A(n6751), .B(n6752), .Z(n6750) );
  XNOR U6474 ( .A(p_input[3386]), .B(n6749), .Z(n6752) );
  XNOR U6475 ( .A(n6749), .B(n6371), .Z(n6751) );
  IV U6476 ( .A(p_input[3354]), .Z(n6371) );
  XOR U6477 ( .A(n6753), .B(n6754), .Z(n6749) );
  AND U6478 ( .A(n6755), .B(n6756), .Z(n6754) );
  XNOR U6479 ( .A(p_input[3385]), .B(n6753), .Z(n6756) );
  XNOR U6480 ( .A(n6753), .B(n6380), .Z(n6755) );
  IV U6481 ( .A(p_input[3353]), .Z(n6380) );
  XOR U6482 ( .A(n6757), .B(n6758), .Z(n6753) );
  AND U6483 ( .A(n6759), .B(n6760), .Z(n6758) );
  XNOR U6484 ( .A(p_input[3384]), .B(n6757), .Z(n6760) );
  XNOR U6485 ( .A(n6757), .B(n6389), .Z(n6759) );
  IV U6486 ( .A(p_input[3352]), .Z(n6389) );
  XOR U6487 ( .A(n6761), .B(n6762), .Z(n6757) );
  AND U6488 ( .A(n6763), .B(n6764), .Z(n6762) );
  XNOR U6489 ( .A(p_input[3383]), .B(n6761), .Z(n6764) );
  XNOR U6490 ( .A(n6761), .B(n6398), .Z(n6763) );
  IV U6491 ( .A(p_input[3351]), .Z(n6398) );
  XOR U6492 ( .A(n6765), .B(n6766), .Z(n6761) );
  AND U6493 ( .A(n6767), .B(n6768), .Z(n6766) );
  XNOR U6494 ( .A(p_input[3382]), .B(n6765), .Z(n6768) );
  XNOR U6495 ( .A(n6765), .B(n6407), .Z(n6767) );
  IV U6496 ( .A(p_input[3350]), .Z(n6407) );
  XOR U6497 ( .A(n6769), .B(n6770), .Z(n6765) );
  AND U6498 ( .A(n6771), .B(n6772), .Z(n6770) );
  XNOR U6499 ( .A(p_input[3381]), .B(n6769), .Z(n6772) );
  XNOR U6500 ( .A(n6769), .B(n6416), .Z(n6771) );
  IV U6501 ( .A(p_input[3349]), .Z(n6416) );
  XOR U6502 ( .A(n6773), .B(n6774), .Z(n6769) );
  AND U6503 ( .A(n6775), .B(n6776), .Z(n6774) );
  XNOR U6504 ( .A(p_input[3380]), .B(n6773), .Z(n6776) );
  XNOR U6505 ( .A(n6773), .B(n6425), .Z(n6775) );
  IV U6506 ( .A(p_input[3348]), .Z(n6425) );
  XOR U6507 ( .A(n6777), .B(n6778), .Z(n6773) );
  AND U6508 ( .A(n6779), .B(n6780), .Z(n6778) );
  XNOR U6509 ( .A(p_input[3379]), .B(n6777), .Z(n6780) );
  XNOR U6510 ( .A(n6777), .B(n6434), .Z(n6779) );
  IV U6511 ( .A(p_input[3347]), .Z(n6434) );
  XOR U6512 ( .A(n6781), .B(n6782), .Z(n6777) );
  AND U6513 ( .A(n6783), .B(n6784), .Z(n6782) );
  XNOR U6514 ( .A(p_input[3378]), .B(n6781), .Z(n6784) );
  XNOR U6515 ( .A(n6781), .B(n6443), .Z(n6783) );
  IV U6516 ( .A(p_input[3346]), .Z(n6443) );
  XOR U6517 ( .A(n6785), .B(n6786), .Z(n6781) );
  AND U6518 ( .A(n6787), .B(n6788), .Z(n6786) );
  XNOR U6519 ( .A(p_input[3377]), .B(n6785), .Z(n6788) );
  XNOR U6520 ( .A(n6785), .B(n6452), .Z(n6787) );
  IV U6521 ( .A(p_input[3345]), .Z(n6452) );
  XOR U6522 ( .A(n6789), .B(n6790), .Z(n6785) );
  AND U6523 ( .A(n6791), .B(n6792), .Z(n6790) );
  XNOR U6524 ( .A(p_input[3376]), .B(n6789), .Z(n6792) );
  XNOR U6525 ( .A(n6789), .B(n6461), .Z(n6791) );
  IV U6526 ( .A(p_input[3344]), .Z(n6461) );
  XOR U6527 ( .A(n6793), .B(n6794), .Z(n6789) );
  AND U6528 ( .A(n6795), .B(n6796), .Z(n6794) );
  XNOR U6529 ( .A(p_input[3375]), .B(n6793), .Z(n6796) );
  XNOR U6530 ( .A(n6793), .B(n6470), .Z(n6795) );
  IV U6531 ( .A(p_input[3343]), .Z(n6470) );
  XOR U6532 ( .A(n6797), .B(n6798), .Z(n6793) );
  AND U6533 ( .A(n6799), .B(n6800), .Z(n6798) );
  XNOR U6534 ( .A(p_input[3374]), .B(n6797), .Z(n6800) );
  XNOR U6535 ( .A(n6797), .B(n6479), .Z(n6799) );
  IV U6536 ( .A(p_input[3342]), .Z(n6479) );
  XOR U6537 ( .A(n6801), .B(n6802), .Z(n6797) );
  AND U6538 ( .A(n6803), .B(n6804), .Z(n6802) );
  XNOR U6539 ( .A(p_input[3373]), .B(n6801), .Z(n6804) );
  XNOR U6540 ( .A(n6801), .B(n6488), .Z(n6803) );
  IV U6541 ( .A(p_input[3341]), .Z(n6488) );
  XOR U6542 ( .A(n6805), .B(n6806), .Z(n6801) );
  AND U6543 ( .A(n6807), .B(n6808), .Z(n6806) );
  XNOR U6544 ( .A(p_input[3372]), .B(n6805), .Z(n6808) );
  XNOR U6545 ( .A(n6805), .B(n6497), .Z(n6807) );
  IV U6546 ( .A(p_input[3340]), .Z(n6497) );
  XOR U6547 ( .A(n6809), .B(n6810), .Z(n6805) );
  AND U6548 ( .A(n6811), .B(n6812), .Z(n6810) );
  XNOR U6549 ( .A(p_input[3371]), .B(n6809), .Z(n6812) );
  XNOR U6550 ( .A(n6809), .B(n6506), .Z(n6811) );
  IV U6551 ( .A(p_input[3339]), .Z(n6506) );
  XOR U6552 ( .A(n6813), .B(n6814), .Z(n6809) );
  AND U6553 ( .A(n6815), .B(n6816), .Z(n6814) );
  XNOR U6554 ( .A(p_input[3370]), .B(n6813), .Z(n6816) );
  XNOR U6555 ( .A(n6813), .B(n6515), .Z(n6815) );
  IV U6556 ( .A(p_input[3338]), .Z(n6515) );
  XOR U6557 ( .A(n6817), .B(n6818), .Z(n6813) );
  AND U6558 ( .A(n6819), .B(n6820), .Z(n6818) );
  XNOR U6559 ( .A(p_input[3369]), .B(n6817), .Z(n6820) );
  XNOR U6560 ( .A(n6817), .B(n6524), .Z(n6819) );
  IV U6561 ( .A(p_input[3337]), .Z(n6524) );
  XOR U6562 ( .A(n6821), .B(n6822), .Z(n6817) );
  AND U6563 ( .A(n6823), .B(n6824), .Z(n6822) );
  XNOR U6564 ( .A(p_input[3368]), .B(n6821), .Z(n6824) );
  XNOR U6565 ( .A(n6821), .B(n6533), .Z(n6823) );
  IV U6566 ( .A(p_input[3336]), .Z(n6533) );
  XOR U6567 ( .A(n6825), .B(n6826), .Z(n6821) );
  AND U6568 ( .A(n6827), .B(n6828), .Z(n6826) );
  XNOR U6569 ( .A(p_input[3367]), .B(n6825), .Z(n6828) );
  XNOR U6570 ( .A(n6825), .B(n6542), .Z(n6827) );
  IV U6571 ( .A(p_input[3335]), .Z(n6542) );
  XOR U6572 ( .A(n6829), .B(n6830), .Z(n6825) );
  AND U6573 ( .A(n6831), .B(n6832), .Z(n6830) );
  XNOR U6574 ( .A(p_input[3366]), .B(n6829), .Z(n6832) );
  XNOR U6575 ( .A(n6829), .B(n6551), .Z(n6831) );
  IV U6576 ( .A(p_input[3334]), .Z(n6551) );
  XOR U6577 ( .A(n6833), .B(n6834), .Z(n6829) );
  AND U6578 ( .A(n6835), .B(n6836), .Z(n6834) );
  XNOR U6579 ( .A(p_input[3365]), .B(n6833), .Z(n6836) );
  XNOR U6580 ( .A(n6833), .B(n6560), .Z(n6835) );
  IV U6581 ( .A(p_input[3333]), .Z(n6560) );
  XOR U6582 ( .A(n6837), .B(n6838), .Z(n6833) );
  AND U6583 ( .A(n6839), .B(n6840), .Z(n6838) );
  XNOR U6584 ( .A(p_input[3364]), .B(n6837), .Z(n6840) );
  XNOR U6585 ( .A(n6837), .B(n6569), .Z(n6839) );
  IV U6586 ( .A(p_input[3332]), .Z(n6569) );
  XOR U6587 ( .A(n6841), .B(n6842), .Z(n6837) );
  AND U6588 ( .A(n6843), .B(n6844), .Z(n6842) );
  XNOR U6589 ( .A(p_input[3363]), .B(n6841), .Z(n6844) );
  XNOR U6590 ( .A(n6841), .B(n6578), .Z(n6843) );
  IV U6591 ( .A(p_input[3331]), .Z(n6578) );
  XOR U6592 ( .A(n6845), .B(n6846), .Z(n6841) );
  AND U6593 ( .A(n6847), .B(n6848), .Z(n6846) );
  XNOR U6594 ( .A(p_input[3362]), .B(n6845), .Z(n6848) );
  XNOR U6595 ( .A(n6845), .B(n6587), .Z(n6847) );
  IV U6596 ( .A(p_input[3330]), .Z(n6587) );
  XNOR U6597 ( .A(n6849), .B(n6850), .Z(n6845) );
  AND U6598 ( .A(n6851), .B(n6852), .Z(n6850) );
  XOR U6599 ( .A(p_input[3361]), .B(n6849), .Z(n6852) );
  XNOR U6600 ( .A(p_input[3329]), .B(n6849), .Z(n6851) );
  AND U6601 ( .A(p_input[3360]), .B(n6853), .Z(n6849) );
  IV U6602 ( .A(p_input[3328]), .Z(n6853) );
  XOR U6603 ( .A(n6854), .B(n6855), .Z(n5032) );
  AND U6604 ( .A(n491), .B(n6856), .Z(n6855) );
  XNOR U6605 ( .A(n6857), .B(n6854), .Z(n6856) );
  XOR U6606 ( .A(n6858), .B(n6859), .Z(n491) );
  AND U6607 ( .A(n6860), .B(n6861), .Z(n6859) );
  XOR U6608 ( .A(n6858), .B(n5047), .Z(n6861) );
  XNOR U6609 ( .A(n6862), .B(n6863), .Z(n5047) );
  AND U6610 ( .A(n6864), .B(n322), .Z(n6863) );
  AND U6611 ( .A(n6862), .B(n6865), .Z(n6864) );
  XNOR U6612 ( .A(n5044), .B(n6858), .Z(n6860) );
  XOR U6613 ( .A(n6866), .B(n6867), .Z(n5044) );
  AND U6614 ( .A(n6868), .B(n319), .Z(n6867) );
  NOR U6615 ( .A(n6866), .B(n6869), .Z(n6868) );
  XOR U6616 ( .A(n6870), .B(n6871), .Z(n6858) );
  AND U6617 ( .A(n6872), .B(n6873), .Z(n6871) );
  XOR U6618 ( .A(n6870), .B(n5059), .Z(n6873) );
  XOR U6619 ( .A(n6874), .B(n6875), .Z(n5059) );
  AND U6620 ( .A(n322), .B(n6876), .Z(n6875) );
  XOR U6621 ( .A(n6877), .B(n6874), .Z(n6876) );
  XNOR U6622 ( .A(n5056), .B(n6870), .Z(n6872) );
  XOR U6623 ( .A(n6878), .B(n6879), .Z(n5056) );
  AND U6624 ( .A(n319), .B(n6880), .Z(n6879) );
  XOR U6625 ( .A(n6881), .B(n6878), .Z(n6880) );
  XOR U6626 ( .A(n6882), .B(n6883), .Z(n6870) );
  AND U6627 ( .A(n6884), .B(n6885), .Z(n6883) );
  XOR U6628 ( .A(n6882), .B(n5071), .Z(n6885) );
  XOR U6629 ( .A(n6886), .B(n6887), .Z(n5071) );
  AND U6630 ( .A(n322), .B(n6888), .Z(n6887) );
  XOR U6631 ( .A(n6889), .B(n6886), .Z(n6888) );
  XNOR U6632 ( .A(n5068), .B(n6882), .Z(n6884) );
  XOR U6633 ( .A(n6890), .B(n6891), .Z(n5068) );
  AND U6634 ( .A(n319), .B(n6892), .Z(n6891) );
  XOR U6635 ( .A(n6893), .B(n6890), .Z(n6892) );
  XOR U6636 ( .A(n6894), .B(n6895), .Z(n6882) );
  AND U6637 ( .A(n6896), .B(n6897), .Z(n6895) );
  XOR U6638 ( .A(n6894), .B(n5083), .Z(n6897) );
  XOR U6639 ( .A(n6898), .B(n6899), .Z(n5083) );
  AND U6640 ( .A(n322), .B(n6900), .Z(n6899) );
  XOR U6641 ( .A(n6901), .B(n6898), .Z(n6900) );
  XNOR U6642 ( .A(n5080), .B(n6894), .Z(n6896) );
  XOR U6643 ( .A(n6902), .B(n6903), .Z(n5080) );
  AND U6644 ( .A(n319), .B(n6904), .Z(n6903) );
  XOR U6645 ( .A(n6905), .B(n6902), .Z(n6904) );
  XOR U6646 ( .A(n6906), .B(n6907), .Z(n6894) );
  AND U6647 ( .A(n6908), .B(n6909), .Z(n6907) );
  XOR U6648 ( .A(n6906), .B(n5095), .Z(n6909) );
  XOR U6649 ( .A(n6910), .B(n6911), .Z(n5095) );
  AND U6650 ( .A(n322), .B(n6912), .Z(n6911) );
  XOR U6651 ( .A(n6913), .B(n6910), .Z(n6912) );
  XNOR U6652 ( .A(n5092), .B(n6906), .Z(n6908) );
  XOR U6653 ( .A(n6914), .B(n6915), .Z(n5092) );
  AND U6654 ( .A(n319), .B(n6916), .Z(n6915) );
  XOR U6655 ( .A(n6917), .B(n6914), .Z(n6916) );
  XOR U6656 ( .A(n6918), .B(n6919), .Z(n6906) );
  AND U6657 ( .A(n6920), .B(n6921), .Z(n6919) );
  XOR U6658 ( .A(n6918), .B(n5107), .Z(n6921) );
  XOR U6659 ( .A(n6922), .B(n6923), .Z(n5107) );
  AND U6660 ( .A(n322), .B(n6924), .Z(n6923) );
  XOR U6661 ( .A(n6925), .B(n6922), .Z(n6924) );
  XNOR U6662 ( .A(n5104), .B(n6918), .Z(n6920) );
  XOR U6663 ( .A(n6926), .B(n6927), .Z(n5104) );
  AND U6664 ( .A(n319), .B(n6928), .Z(n6927) );
  XOR U6665 ( .A(n6929), .B(n6926), .Z(n6928) );
  XOR U6666 ( .A(n6930), .B(n6931), .Z(n6918) );
  AND U6667 ( .A(n6932), .B(n6933), .Z(n6931) );
  XOR U6668 ( .A(n6930), .B(n5119), .Z(n6933) );
  XOR U6669 ( .A(n6934), .B(n6935), .Z(n5119) );
  AND U6670 ( .A(n322), .B(n6936), .Z(n6935) );
  XOR U6671 ( .A(n6937), .B(n6934), .Z(n6936) );
  XNOR U6672 ( .A(n5116), .B(n6930), .Z(n6932) );
  XOR U6673 ( .A(n6938), .B(n6939), .Z(n5116) );
  AND U6674 ( .A(n319), .B(n6940), .Z(n6939) );
  XOR U6675 ( .A(n6941), .B(n6938), .Z(n6940) );
  XOR U6676 ( .A(n6942), .B(n6943), .Z(n6930) );
  AND U6677 ( .A(n6944), .B(n6945), .Z(n6943) );
  XOR U6678 ( .A(n6942), .B(n5131), .Z(n6945) );
  XOR U6679 ( .A(n6946), .B(n6947), .Z(n5131) );
  AND U6680 ( .A(n322), .B(n6948), .Z(n6947) );
  XOR U6681 ( .A(n6949), .B(n6946), .Z(n6948) );
  XNOR U6682 ( .A(n5128), .B(n6942), .Z(n6944) );
  XOR U6683 ( .A(n6950), .B(n6951), .Z(n5128) );
  AND U6684 ( .A(n319), .B(n6952), .Z(n6951) );
  XOR U6685 ( .A(n6953), .B(n6950), .Z(n6952) );
  XOR U6686 ( .A(n6954), .B(n6955), .Z(n6942) );
  AND U6687 ( .A(n6956), .B(n6957), .Z(n6955) );
  XOR U6688 ( .A(n6954), .B(n5143), .Z(n6957) );
  XOR U6689 ( .A(n6958), .B(n6959), .Z(n5143) );
  AND U6690 ( .A(n322), .B(n6960), .Z(n6959) );
  XOR U6691 ( .A(n6961), .B(n6958), .Z(n6960) );
  XNOR U6692 ( .A(n5140), .B(n6954), .Z(n6956) );
  XOR U6693 ( .A(n6962), .B(n6963), .Z(n5140) );
  AND U6694 ( .A(n319), .B(n6964), .Z(n6963) );
  XOR U6695 ( .A(n6965), .B(n6962), .Z(n6964) );
  XOR U6696 ( .A(n6966), .B(n6967), .Z(n6954) );
  AND U6697 ( .A(n6968), .B(n6969), .Z(n6967) );
  XOR U6698 ( .A(n6966), .B(n5155), .Z(n6969) );
  XOR U6699 ( .A(n6970), .B(n6971), .Z(n5155) );
  AND U6700 ( .A(n322), .B(n6972), .Z(n6971) );
  XOR U6701 ( .A(n6973), .B(n6970), .Z(n6972) );
  XNOR U6702 ( .A(n5152), .B(n6966), .Z(n6968) );
  XOR U6703 ( .A(n6974), .B(n6975), .Z(n5152) );
  AND U6704 ( .A(n319), .B(n6976), .Z(n6975) );
  XOR U6705 ( .A(n6977), .B(n6974), .Z(n6976) );
  XOR U6706 ( .A(n6978), .B(n6979), .Z(n6966) );
  AND U6707 ( .A(n6980), .B(n6981), .Z(n6979) );
  XOR U6708 ( .A(n6978), .B(n5167), .Z(n6981) );
  XOR U6709 ( .A(n6982), .B(n6983), .Z(n5167) );
  AND U6710 ( .A(n322), .B(n6984), .Z(n6983) );
  XOR U6711 ( .A(n6985), .B(n6982), .Z(n6984) );
  XNOR U6712 ( .A(n5164), .B(n6978), .Z(n6980) );
  XOR U6713 ( .A(n6986), .B(n6987), .Z(n5164) );
  AND U6714 ( .A(n319), .B(n6988), .Z(n6987) );
  XOR U6715 ( .A(n6989), .B(n6986), .Z(n6988) );
  XOR U6716 ( .A(n6990), .B(n6991), .Z(n6978) );
  AND U6717 ( .A(n6992), .B(n6993), .Z(n6991) );
  XOR U6718 ( .A(n6990), .B(n5179), .Z(n6993) );
  XOR U6719 ( .A(n6994), .B(n6995), .Z(n5179) );
  AND U6720 ( .A(n322), .B(n6996), .Z(n6995) );
  XOR U6721 ( .A(n6997), .B(n6994), .Z(n6996) );
  XNOR U6722 ( .A(n5176), .B(n6990), .Z(n6992) );
  XOR U6723 ( .A(n6998), .B(n6999), .Z(n5176) );
  AND U6724 ( .A(n319), .B(n7000), .Z(n6999) );
  XOR U6725 ( .A(n7001), .B(n6998), .Z(n7000) );
  XOR U6726 ( .A(n7002), .B(n7003), .Z(n6990) );
  AND U6727 ( .A(n7004), .B(n7005), .Z(n7003) );
  XOR U6728 ( .A(n7002), .B(n5191), .Z(n7005) );
  XOR U6729 ( .A(n7006), .B(n7007), .Z(n5191) );
  AND U6730 ( .A(n322), .B(n7008), .Z(n7007) );
  XOR U6731 ( .A(n7009), .B(n7006), .Z(n7008) );
  XNOR U6732 ( .A(n5188), .B(n7002), .Z(n7004) );
  XOR U6733 ( .A(n7010), .B(n7011), .Z(n5188) );
  AND U6734 ( .A(n319), .B(n7012), .Z(n7011) );
  XOR U6735 ( .A(n7013), .B(n7010), .Z(n7012) );
  XOR U6736 ( .A(n7014), .B(n7015), .Z(n7002) );
  AND U6737 ( .A(n7016), .B(n7017), .Z(n7015) );
  XOR U6738 ( .A(n7014), .B(n5203), .Z(n7017) );
  XOR U6739 ( .A(n7018), .B(n7019), .Z(n5203) );
  AND U6740 ( .A(n322), .B(n7020), .Z(n7019) );
  XOR U6741 ( .A(n7021), .B(n7018), .Z(n7020) );
  XNOR U6742 ( .A(n5200), .B(n7014), .Z(n7016) );
  XOR U6743 ( .A(n7022), .B(n7023), .Z(n5200) );
  AND U6744 ( .A(n319), .B(n7024), .Z(n7023) );
  XOR U6745 ( .A(n7025), .B(n7022), .Z(n7024) );
  XOR U6746 ( .A(n7026), .B(n7027), .Z(n7014) );
  AND U6747 ( .A(n7028), .B(n7029), .Z(n7027) );
  XOR U6748 ( .A(n7026), .B(n5215), .Z(n7029) );
  XOR U6749 ( .A(n7030), .B(n7031), .Z(n5215) );
  AND U6750 ( .A(n322), .B(n7032), .Z(n7031) );
  XOR U6751 ( .A(n7033), .B(n7030), .Z(n7032) );
  XNOR U6752 ( .A(n5212), .B(n7026), .Z(n7028) );
  XOR U6753 ( .A(n7034), .B(n7035), .Z(n5212) );
  AND U6754 ( .A(n319), .B(n7036), .Z(n7035) );
  XOR U6755 ( .A(n7037), .B(n7034), .Z(n7036) );
  XOR U6756 ( .A(n7038), .B(n7039), .Z(n7026) );
  AND U6757 ( .A(n7040), .B(n7041), .Z(n7039) );
  XOR U6758 ( .A(n7038), .B(n5227), .Z(n7041) );
  XOR U6759 ( .A(n7042), .B(n7043), .Z(n5227) );
  AND U6760 ( .A(n322), .B(n7044), .Z(n7043) );
  XOR U6761 ( .A(n7045), .B(n7042), .Z(n7044) );
  XNOR U6762 ( .A(n5224), .B(n7038), .Z(n7040) );
  XOR U6763 ( .A(n7046), .B(n7047), .Z(n5224) );
  AND U6764 ( .A(n319), .B(n7048), .Z(n7047) );
  XOR U6765 ( .A(n7049), .B(n7046), .Z(n7048) );
  XOR U6766 ( .A(n7050), .B(n7051), .Z(n7038) );
  AND U6767 ( .A(n7052), .B(n7053), .Z(n7051) );
  XOR U6768 ( .A(n7050), .B(n5239), .Z(n7053) );
  XOR U6769 ( .A(n7054), .B(n7055), .Z(n5239) );
  AND U6770 ( .A(n322), .B(n7056), .Z(n7055) );
  XOR U6771 ( .A(n7057), .B(n7054), .Z(n7056) );
  XNOR U6772 ( .A(n5236), .B(n7050), .Z(n7052) );
  XOR U6773 ( .A(n7058), .B(n7059), .Z(n5236) );
  AND U6774 ( .A(n319), .B(n7060), .Z(n7059) );
  XOR U6775 ( .A(n7061), .B(n7058), .Z(n7060) );
  XOR U6776 ( .A(n7062), .B(n7063), .Z(n7050) );
  AND U6777 ( .A(n7064), .B(n7065), .Z(n7063) );
  XOR U6778 ( .A(n7062), .B(n5251), .Z(n7065) );
  XOR U6779 ( .A(n7066), .B(n7067), .Z(n5251) );
  AND U6780 ( .A(n322), .B(n7068), .Z(n7067) );
  XOR U6781 ( .A(n7069), .B(n7066), .Z(n7068) );
  XNOR U6782 ( .A(n5248), .B(n7062), .Z(n7064) );
  XOR U6783 ( .A(n7070), .B(n7071), .Z(n5248) );
  AND U6784 ( .A(n319), .B(n7072), .Z(n7071) );
  XOR U6785 ( .A(n7073), .B(n7070), .Z(n7072) );
  XOR U6786 ( .A(n7074), .B(n7075), .Z(n7062) );
  AND U6787 ( .A(n7076), .B(n7077), .Z(n7075) );
  XOR U6788 ( .A(n7074), .B(n5263), .Z(n7077) );
  XOR U6789 ( .A(n7078), .B(n7079), .Z(n5263) );
  AND U6790 ( .A(n322), .B(n7080), .Z(n7079) );
  XOR U6791 ( .A(n7081), .B(n7078), .Z(n7080) );
  XNOR U6792 ( .A(n5260), .B(n7074), .Z(n7076) );
  XOR U6793 ( .A(n7082), .B(n7083), .Z(n5260) );
  AND U6794 ( .A(n319), .B(n7084), .Z(n7083) );
  XOR U6795 ( .A(n7085), .B(n7082), .Z(n7084) );
  XOR U6796 ( .A(n7086), .B(n7087), .Z(n7074) );
  AND U6797 ( .A(n7088), .B(n7089), .Z(n7087) );
  XOR U6798 ( .A(n7086), .B(n5275), .Z(n7089) );
  XOR U6799 ( .A(n7090), .B(n7091), .Z(n5275) );
  AND U6800 ( .A(n322), .B(n7092), .Z(n7091) );
  XOR U6801 ( .A(n7093), .B(n7090), .Z(n7092) );
  XNOR U6802 ( .A(n5272), .B(n7086), .Z(n7088) );
  XOR U6803 ( .A(n7094), .B(n7095), .Z(n5272) );
  AND U6804 ( .A(n319), .B(n7096), .Z(n7095) );
  XOR U6805 ( .A(n7097), .B(n7094), .Z(n7096) );
  XOR U6806 ( .A(n7098), .B(n7099), .Z(n7086) );
  AND U6807 ( .A(n7100), .B(n7101), .Z(n7099) );
  XOR U6808 ( .A(n7098), .B(n5287), .Z(n7101) );
  XOR U6809 ( .A(n7102), .B(n7103), .Z(n5287) );
  AND U6810 ( .A(n322), .B(n7104), .Z(n7103) );
  XOR U6811 ( .A(n7105), .B(n7102), .Z(n7104) );
  XNOR U6812 ( .A(n5284), .B(n7098), .Z(n7100) );
  XOR U6813 ( .A(n7106), .B(n7107), .Z(n5284) );
  AND U6814 ( .A(n319), .B(n7108), .Z(n7107) );
  XOR U6815 ( .A(n7109), .B(n7106), .Z(n7108) );
  XOR U6816 ( .A(n7110), .B(n7111), .Z(n7098) );
  AND U6817 ( .A(n7112), .B(n7113), .Z(n7111) );
  XOR U6818 ( .A(n7110), .B(n5299), .Z(n7113) );
  XOR U6819 ( .A(n7114), .B(n7115), .Z(n5299) );
  AND U6820 ( .A(n322), .B(n7116), .Z(n7115) );
  XOR U6821 ( .A(n7117), .B(n7114), .Z(n7116) );
  XNOR U6822 ( .A(n5296), .B(n7110), .Z(n7112) );
  XOR U6823 ( .A(n7118), .B(n7119), .Z(n5296) );
  AND U6824 ( .A(n319), .B(n7120), .Z(n7119) );
  XOR U6825 ( .A(n7121), .B(n7118), .Z(n7120) );
  XOR U6826 ( .A(n7122), .B(n7123), .Z(n7110) );
  AND U6827 ( .A(n7124), .B(n7125), .Z(n7123) );
  XOR U6828 ( .A(n7122), .B(n5311), .Z(n7125) );
  XOR U6829 ( .A(n7126), .B(n7127), .Z(n5311) );
  AND U6830 ( .A(n322), .B(n7128), .Z(n7127) );
  XOR U6831 ( .A(n7129), .B(n7126), .Z(n7128) );
  XNOR U6832 ( .A(n5308), .B(n7122), .Z(n7124) );
  XOR U6833 ( .A(n7130), .B(n7131), .Z(n5308) );
  AND U6834 ( .A(n319), .B(n7132), .Z(n7131) );
  XOR U6835 ( .A(n7133), .B(n7130), .Z(n7132) );
  XOR U6836 ( .A(n7134), .B(n7135), .Z(n7122) );
  AND U6837 ( .A(n7136), .B(n7137), .Z(n7135) );
  XOR U6838 ( .A(n7134), .B(n5323), .Z(n7137) );
  XOR U6839 ( .A(n7138), .B(n7139), .Z(n5323) );
  AND U6840 ( .A(n322), .B(n7140), .Z(n7139) );
  XOR U6841 ( .A(n7141), .B(n7138), .Z(n7140) );
  XNOR U6842 ( .A(n5320), .B(n7134), .Z(n7136) );
  XOR U6843 ( .A(n7142), .B(n7143), .Z(n5320) );
  AND U6844 ( .A(n319), .B(n7144), .Z(n7143) );
  XOR U6845 ( .A(n7145), .B(n7142), .Z(n7144) );
  XOR U6846 ( .A(n7146), .B(n7147), .Z(n7134) );
  AND U6847 ( .A(n7148), .B(n7149), .Z(n7147) );
  XOR U6848 ( .A(n7146), .B(n5335), .Z(n7149) );
  XOR U6849 ( .A(n7150), .B(n7151), .Z(n5335) );
  AND U6850 ( .A(n322), .B(n7152), .Z(n7151) );
  XOR U6851 ( .A(n7153), .B(n7150), .Z(n7152) );
  XNOR U6852 ( .A(n5332), .B(n7146), .Z(n7148) );
  XOR U6853 ( .A(n7154), .B(n7155), .Z(n5332) );
  AND U6854 ( .A(n319), .B(n7156), .Z(n7155) );
  XOR U6855 ( .A(n7157), .B(n7154), .Z(n7156) );
  XOR U6856 ( .A(n7158), .B(n7159), .Z(n7146) );
  AND U6857 ( .A(n7160), .B(n7161), .Z(n7159) );
  XOR U6858 ( .A(n7158), .B(n5347), .Z(n7161) );
  XOR U6859 ( .A(n7162), .B(n7163), .Z(n5347) );
  AND U6860 ( .A(n322), .B(n7164), .Z(n7163) );
  XOR U6861 ( .A(n7165), .B(n7162), .Z(n7164) );
  XNOR U6862 ( .A(n5344), .B(n7158), .Z(n7160) );
  XOR U6863 ( .A(n7166), .B(n7167), .Z(n5344) );
  AND U6864 ( .A(n319), .B(n7168), .Z(n7167) );
  XOR U6865 ( .A(n7169), .B(n7166), .Z(n7168) );
  XOR U6866 ( .A(n7170), .B(n7171), .Z(n7158) );
  AND U6867 ( .A(n7172), .B(n7173), .Z(n7171) );
  XOR U6868 ( .A(n7170), .B(n5359), .Z(n7173) );
  XOR U6869 ( .A(n7174), .B(n7175), .Z(n5359) );
  AND U6870 ( .A(n322), .B(n7176), .Z(n7175) );
  XOR U6871 ( .A(n7177), .B(n7174), .Z(n7176) );
  XNOR U6872 ( .A(n5356), .B(n7170), .Z(n7172) );
  XOR U6873 ( .A(n7178), .B(n7179), .Z(n5356) );
  AND U6874 ( .A(n319), .B(n7180), .Z(n7179) );
  XOR U6875 ( .A(n7181), .B(n7178), .Z(n7180) );
  XOR U6876 ( .A(n7182), .B(n7183), .Z(n7170) );
  AND U6877 ( .A(n7184), .B(n7185), .Z(n7183) );
  XOR U6878 ( .A(n7182), .B(n5371), .Z(n7185) );
  XOR U6879 ( .A(n7186), .B(n7187), .Z(n5371) );
  AND U6880 ( .A(n322), .B(n7188), .Z(n7187) );
  XOR U6881 ( .A(n7189), .B(n7186), .Z(n7188) );
  XNOR U6882 ( .A(n5368), .B(n7182), .Z(n7184) );
  XOR U6883 ( .A(n7190), .B(n7191), .Z(n5368) );
  AND U6884 ( .A(n319), .B(n7192), .Z(n7191) );
  XOR U6885 ( .A(n7193), .B(n7190), .Z(n7192) );
  XOR U6886 ( .A(n7194), .B(n7195), .Z(n7182) );
  AND U6887 ( .A(n7196), .B(n7197), .Z(n7195) );
  XOR U6888 ( .A(n7194), .B(n5383), .Z(n7197) );
  XOR U6889 ( .A(n7198), .B(n7199), .Z(n5383) );
  AND U6890 ( .A(n322), .B(n7200), .Z(n7199) );
  XOR U6891 ( .A(n7201), .B(n7198), .Z(n7200) );
  XNOR U6892 ( .A(n5380), .B(n7194), .Z(n7196) );
  XOR U6893 ( .A(n7202), .B(n7203), .Z(n5380) );
  AND U6894 ( .A(n319), .B(n7204), .Z(n7203) );
  XOR U6895 ( .A(n7205), .B(n7202), .Z(n7204) );
  XOR U6896 ( .A(n7206), .B(n7207), .Z(n7194) );
  AND U6897 ( .A(n7208), .B(n7209), .Z(n7207) );
  XOR U6898 ( .A(n5395), .B(n7206), .Z(n7209) );
  XOR U6899 ( .A(n7210), .B(n7211), .Z(n5395) );
  AND U6900 ( .A(n322), .B(n7212), .Z(n7211) );
  XOR U6901 ( .A(n7210), .B(n7213), .Z(n7212) );
  XNOR U6902 ( .A(n7206), .B(n5392), .Z(n7208) );
  XOR U6903 ( .A(n7214), .B(n7215), .Z(n5392) );
  AND U6904 ( .A(n319), .B(n7216), .Z(n7215) );
  XOR U6905 ( .A(n7214), .B(n7217), .Z(n7216) );
  XOR U6906 ( .A(n7218), .B(n7219), .Z(n7206) );
  AND U6907 ( .A(n7220), .B(n7221), .Z(n7219) );
  XNOR U6908 ( .A(n7222), .B(n5408), .Z(n7221) );
  XOR U6909 ( .A(n7223), .B(n7224), .Z(n5408) );
  AND U6910 ( .A(n322), .B(n7225), .Z(n7224) );
  XOR U6911 ( .A(n7226), .B(n7223), .Z(n7225) );
  XNOR U6912 ( .A(n5405), .B(n7218), .Z(n7220) );
  XOR U6913 ( .A(n7227), .B(n7228), .Z(n5405) );
  AND U6914 ( .A(n319), .B(n7229), .Z(n7228) );
  XOR U6915 ( .A(n7230), .B(n7227), .Z(n7229) );
  IV U6916 ( .A(n7222), .Z(n7218) );
  AND U6917 ( .A(n6854), .B(n6857), .Z(n7222) );
  XNOR U6918 ( .A(n7231), .B(n7232), .Z(n6857) );
  AND U6919 ( .A(n322), .B(n7233), .Z(n7232) );
  XNOR U6920 ( .A(n7234), .B(n7231), .Z(n7233) );
  XOR U6921 ( .A(n7235), .B(n7236), .Z(n322) );
  AND U6922 ( .A(n7237), .B(n7238), .Z(n7236) );
  XOR U6923 ( .A(n6865), .B(n7235), .Z(n7238) );
  IV U6924 ( .A(n7239), .Z(n6865) );
  AND U6925 ( .A(p_input[3327]), .B(p_input[3295]), .Z(n7239) );
  XOR U6926 ( .A(n7235), .B(n6862), .Z(n7237) );
  AND U6927 ( .A(p_input[3231]), .B(p_input[3263]), .Z(n6862) );
  XOR U6928 ( .A(n7240), .B(n7241), .Z(n7235) );
  AND U6929 ( .A(n7242), .B(n7243), .Z(n7241) );
  XOR U6930 ( .A(n7240), .B(n6877), .Z(n7243) );
  XNOR U6931 ( .A(p_input[3294]), .B(n7244), .Z(n6877) );
  AND U6932 ( .A(n222), .B(n7245), .Z(n7244) );
  XOR U6933 ( .A(p_input[3326]), .B(p_input[3294]), .Z(n7245) );
  XNOR U6934 ( .A(n6874), .B(n7240), .Z(n7242) );
  XOR U6935 ( .A(n7246), .B(n7247), .Z(n6874) );
  AND U6936 ( .A(n220), .B(n7248), .Z(n7247) );
  XOR U6937 ( .A(p_input[3262]), .B(p_input[3230]), .Z(n7248) );
  XOR U6938 ( .A(n7249), .B(n7250), .Z(n7240) );
  AND U6939 ( .A(n7251), .B(n7252), .Z(n7250) );
  XOR U6940 ( .A(n7249), .B(n6889), .Z(n7252) );
  XNOR U6941 ( .A(p_input[3293]), .B(n7253), .Z(n6889) );
  AND U6942 ( .A(n222), .B(n7254), .Z(n7253) );
  XOR U6943 ( .A(p_input[3325]), .B(p_input[3293]), .Z(n7254) );
  XNOR U6944 ( .A(n6886), .B(n7249), .Z(n7251) );
  XOR U6945 ( .A(n7255), .B(n7256), .Z(n6886) );
  AND U6946 ( .A(n220), .B(n7257), .Z(n7256) );
  XOR U6947 ( .A(p_input[3261]), .B(p_input[3229]), .Z(n7257) );
  XOR U6948 ( .A(n7258), .B(n7259), .Z(n7249) );
  AND U6949 ( .A(n7260), .B(n7261), .Z(n7259) );
  XOR U6950 ( .A(n7258), .B(n6901), .Z(n7261) );
  XNOR U6951 ( .A(p_input[3292]), .B(n7262), .Z(n6901) );
  AND U6952 ( .A(n222), .B(n7263), .Z(n7262) );
  XOR U6953 ( .A(p_input[3324]), .B(p_input[3292]), .Z(n7263) );
  XNOR U6954 ( .A(n6898), .B(n7258), .Z(n7260) );
  XOR U6955 ( .A(n7264), .B(n7265), .Z(n6898) );
  AND U6956 ( .A(n220), .B(n7266), .Z(n7265) );
  XOR U6957 ( .A(p_input[3260]), .B(p_input[3228]), .Z(n7266) );
  XOR U6958 ( .A(n7267), .B(n7268), .Z(n7258) );
  AND U6959 ( .A(n7269), .B(n7270), .Z(n7268) );
  XOR U6960 ( .A(n7267), .B(n6913), .Z(n7270) );
  XNOR U6961 ( .A(p_input[3291]), .B(n7271), .Z(n6913) );
  AND U6962 ( .A(n222), .B(n7272), .Z(n7271) );
  XOR U6963 ( .A(p_input[3323]), .B(p_input[3291]), .Z(n7272) );
  XNOR U6964 ( .A(n6910), .B(n7267), .Z(n7269) );
  XOR U6965 ( .A(n7273), .B(n7274), .Z(n6910) );
  AND U6966 ( .A(n220), .B(n7275), .Z(n7274) );
  XOR U6967 ( .A(p_input[3259]), .B(p_input[3227]), .Z(n7275) );
  XOR U6968 ( .A(n7276), .B(n7277), .Z(n7267) );
  AND U6969 ( .A(n7278), .B(n7279), .Z(n7277) );
  XOR U6970 ( .A(n7276), .B(n6925), .Z(n7279) );
  XNOR U6971 ( .A(p_input[3290]), .B(n7280), .Z(n6925) );
  AND U6972 ( .A(n222), .B(n7281), .Z(n7280) );
  XOR U6973 ( .A(p_input[3322]), .B(p_input[3290]), .Z(n7281) );
  XNOR U6974 ( .A(n6922), .B(n7276), .Z(n7278) );
  XOR U6975 ( .A(n7282), .B(n7283), .Z(n6922) );
  AND U6976 ( .A(n220), .B(n7284), .Z(n7283) );
  XOR U6977 ( .A(p_input[3258]), .B(p_input[3226]), .Z(n7284) );
  XOR U6978 ( .A(n7285), .B(n7286), .Z(n7276) );
  AND U6979 ( .A(n7287), .B(n7288), .Z(n7286) );
  XOR U6980 ( .A(n7285), .B(n6937), .Z(n7288) );
  XNOR U6981 ( .A(p_input[3289]), .B(n7289), .Z(n6937) );
  AND U6982 ( .A(n222), .B(n7290), .Z(n7289) );
  XOR U6983 ( .A(p_input[3321]), .B(p_input[3289]), .Z(n7290) );
  XNOR U6984 ( .A(n6934), .B(n7285), .Z(n7287) );
  XOR U6985 ( .A(n7291), .B(n7292), .Z(n6934) );
  AND U6986 ( .A(n220), .B(n7293), .Z(n7292) );
  XOR U6987 ( .A(p_input[3257]), .B(p_input[3225]), .Z(n7293) );
  XOR U6988 ( .A(n7294), .B(n7295), .Z(n7285) );
  AND U6989 ( .A(n7296), .B(n7297), .Z(n7295) );
  XOR U6990 ( .A(n7294), .B(n6949), .Z(n7297) );
  XNOR U6991 ( .A(p_input[3288]), .B(n7298), .Z(n6949) );
  AND U6992 ( .A(n222), .B(n7299), .Z(n7298) );
  XOR U6993 ( .A(p_input[3320]), .B(p_input[3288]), .Z(n7299) );
  XNOR U6994 ( .A(n6946), .B(n7294), .Z(n7296) );
  XOR U6995 ( .A(n7300), .B(n7301), .Z(n6946) );
  AND U6996 ( .A(n220), .B(n7302), .Z(n7301) );
  XOR U6997 ( .A(p_input[3256]), .B(p_input[3224]), .Z(n7302) );
  XOR U6998 ( .A(n7303), .B(n7304), .Z(n7294) );
  AND U6999 ( .A(n7305), .B(n7306), .Z(n7304) );
  XOR U7000 ( .A(n7303), .B(n6961), .Z(n7306) );
  XNOR U7001 ( .A(p_input[3287]), .B(n7307), .Z(n6961) );
  AND U7002 ( .A(n222), .B(n7308), .Z(n7307) );
  XOR U7003 ( .A(p_input[3319]), .B(p_input[3287]), .Z(n7308) );
  XNOR U7004 ( .A(n6958), .B(n7303), .Z(n7305) );
  XOR U7005 ( .A(n7309), .B(n7310), .Z(n6958) );
  AND U7006 ( .A(n220), .B(n7311), .Z(n7310) );
  XOR U7007 ( .A(p_input[3255]), .B(p_input[3223]), .Z(n7311) );
  XOR U7008 ( .A(n7312), .B(n7313), .Z(n7303) );
  AND U7009 ( .A(n7314), .B(n7315), .Z(n7313) );
  XOR U7010 ( .A(n7312), .B(n6973), .Z(n7315) );
  XNOR U7011 ( .A(p_input[3286]), .B(n7316), .Z(n6973) );
  AND U7012 ( .A(n222), .B(n7317), .Z(n7316) );
  XOR U7013 ( .A(p_input[3318]), .B(p_input[3286]), .Z(n7317) );
  XNOR U7014 ( .A(n6970), .B(n7312), .Z(n7314) );
  XOR U7015 ( .A(n7318), .B(n7319), .Z(n6970) );
  AND U7016 ( .A(n220), .B(n7320), .Z(n7319) );
  XOR U7017 ( .A(p_input[3254]), .B(p_input[3222]), .Z(n7320) );
  XOR U7018 ( .A(n7321), .B(n7322), .Z(n7312) );
  AND U7019 ( .A(n7323), .B(n7324), .Z(n7322) );
  XOR U7020 ( .A(n7321), .B(n6985), .Z(n7324) );
  XNOR U7021 ( .A(p_input[3285]), .B(n7325), .Z(n6985) );
  AND U7022 ( .A(n222), .B(n7326), .Z(n7325) );
  XOR U7023 ( .A(p_input[3317]), .B(p_input[3285]), .Z(n7326) );
  XNOR U7024 ( .A(n6982), .B(n7321), .Z(n7323) );
  XOR U7025 ( .A(n7327), .B(n7328), .Z(n6982) );
  AND U7026 ( .A(n220), .B(n7329), .Z(n7328) );
  XOR U7027 ( .A(p_input[3253]), .B(p_input[3221]), .Z(n7329) );
  XOR U7028 ( .A(n7330), .B(n7331), .Z(n7321) );
  AND U7029 ( .A(n7332), .B(n7333), .Z(n7331) );
  XOR U7030 ( .A(n7330), .B(n6997), .Z(n7333) );
  XNOR U7031 ( .A(p_input[3284]), .B(n7334), .Z(n6997) );
  AND U7032 ( .A(n222), .B(n7335), .Z(n7334) );
  XOR U7033 ( .A(p_input[3316]), .B(p_input[3284]), .Z(n7335) );
  XNOR U7034 ( .A(n6994), .B(n7330), .Z(n7332) );
  XOR U7035 ( .A(n7336), .B(n7337), .Z(n6994) );
  AND U7036 ( .A(n220), .B(n7338), .Z(n7337) );
  XOR U7037 ( .A(p_input[3252]), .B(p_input[3220]), .Z(n7338) );
  XOR U7038 ( .A(n7339), .B(n7340), .Z(n7330) );
  AND U7039 ( .A(n7341), .B(n7342), .Z(n7340) );
  XOR U7040 ( .A(n7339), .B(n7009), .Z(n7342) );
  XNOR U7041 ( .A(p_input[3283]), .B(n7343), .Z(n7009) );
  AND U7042 ( .A(n222), .B(n7344), .Z(n7343) );
  XOR U7043 ( .A(p_input[3315]), .B(p_input[3283]), .Z(n7344) );
  XNOR U7044 ( .A(n7006), .B(n7339), .Z(n7341) );
  XOR U7045 ( .A(n7345), .B(n7346), .Z(n7006) );
  AND U7046 ( .A(n220), .B(n7347), .Z(n7346) );
  XOR U7047 ( .A(p_input[3251]), .B(p_input[3219]), .Z(n7347) );
  XOR U7048 ( .A(n7348), .B(n7349), .Z(n7339) );
  AND U7049 ( .A(n7350), .B(n7351), .Z(n7349) );
  XOR U7050 ( .A(n7348), .B(n7021), .Z(n7351) );
  XNOR U7051 ( .A(p_input[3282]), .B(n7352), .Z(n7021) );
  AND U7052 ( .A(n222), .B(n7353), .Z(n7352) );
  XOR U7053 ( .A(p_input[3314]), .B(p_input[3282]), .Z(n7353) );
  XNOR U7054 ( .A(n7018), .B(n7348), .Z(n7350) );
  XOR U7055 ( .A(n7354), .B(n7355), .Z(n7018) );
  AND U7056 ( .A(n220), .B(n7356), .Z(n7355) );
  XOR U7057 ( .A(p_input[3250]), .B(p_input[3218]), .Z(n7356) );
  XOR U7058 ( .A(n7357), .B(n7358), .Z(n7348) );
  AND U7059 ( .A(n7359), .B(n7360), .Z(n7358) );
  XOR U7060 ( .A(n7357), .B(n7033), .Z(n7360) );
  XNOR U7061 ( .A(p_input[3281]), .B(n7361), .Z(n7033) );
  AND U7062 ( .A(n222), .B(n7362), .Z(n7361) );
  XOR U7063 ( .A(p_input[3313]), .B(p_input[3281]), .Z(n7362) );
  XNOR U7064 ( .A(n7030), .B(n7357), .Z(n7359) );
  XOR U7065 ( .A(n7363), .B(n7364), .Z(n7030) );
  AND U7066 ( .A(n220), .B(n7365), .Z(n7364) );
  XOR U7067 ( .A(p_input[3249]), .B(p_input[3217]), .Z(n7365) );
  XOR U7068 ( .A(n7366), .B(n7367), .Z(n7357) );
  AND U7069 ( .A(n7368), .B(n7369), .Z(n7367) );
  XOR U7070 ( .A(n7366), .B(n7045), .Z(n7369) );
  XNOR U7071 ( .A(p_input[3280]), .B(n7370), .Z(n7045) );
  AND U7072 ( .A(n222), .B(n7371), .Z(n7370) );
  XOR U7073 ( .A(p_input[3312]), .B(p_input[3280]), .Z(n7371) );
  XNOR U7074 ( .A(n7042), .B(n7366), .Z(n7368) );
  XOR U7075 ( .A(n7372), .B(n7373), .Z(n7042) );
  AND U7076 ( .A(n220), .B(n7374), .Z(n7373) );
  XOR U7077 ( .A(p_input[3248]), .B(p_input[3216]), .Z(n7374) );
  XOR U7078 ( .A(n7375), .B(n7376), .Z(n7366) );
  AND U7079 ( .A(n7377), .B(n7378), .Z(n7376) );
  XOR U7080 ( .A(n7375), .B(n7057), .Z(n7378) );
  XNOR U7081 ( .A(p_input[3279]), .B(n7379), .Z(n7057) );
  AND U7082 ( .A(n222), .B(n7380), .Z(n7379) );
  XOR U7083 ( .A(p_input[3311]), .B(p_input[3279]), .Z(n7380) );
  XNOR U7084 ( .A(n7054), .B(n7375), .Z(n7377) );
  XOR U7085 ( .A(n7381), .B(n7382), .Z(n7054) );
  AND U7086 ( .A(n220), .B(n7383), .Z(n7382) );
  XOR U7087 ( .A(p_input[3247]), .B(p_input[3215]), .Z(n7383) );
  XOR U7088 ( .A(n7384), .B(n7385), .Z(n7375) );
  AND U7089 ( .A(n7386), .B(n7387), .Z(n7385) );
  XOR U7090 ( .A(n7384), .B(n7069), .Z(n7387) );
  XNOR U7091 ( .A(p_input[3278]), .B(n7388), .Z(n7069) );
  AND U7092 ( .A(n222), .B(n7389), .Z(n7388) );
  XOR U7093 ( .A(p_input[3310]), .B(p_input[3278]), .Z(n7389) );
  XNOR U7094 ( .A(n7066), .B(n7384), .Z(n7386) );
  XOR U7095 ( .A(n7390), .B(n7391), .Z(n7066) );
  AND U7096 ( .A(n220), .B(n7392), .Z(n7391) );
  XOR U7097 ( .A(p_input[3246]), .B(p_input[3214]), .Z(n7392) );
  XOR U7098 ( .A(n7393), .B(n7394), .Z(n7384) );
  AND U7099 ( .A(n7395), .B(n7396), .Z(n7394) );
  XOR U7100 ( .A(n7393), .B(n7081), .Z(n7396) );
  XNOR U7101 ( .A(p_input[3277]), .B(n7397), .Z(n7081) );
  AND U7102 ( .A(n222), .B(n7398), .Z(n7397) );
  XOR U7103 ( .A(p_input[3309]), .B(p_input[3277]), .Z(n7398) );
  XNOR U7104 ( .A(n7078), .B(n7393), .Z(n7395) );
  XOR U7105 ( .A(n7399), .B(n7400), .Z(n7078) );
  AND U7106 ( .A(n220), .B(n7401), .Z(n7400) );
  XOR U7107 ( .A(p_input[3245]), .B(p_input[3213]), .Z(n7401) );
  XOR U7108 ( .A(n7402), .B(n7403), .Z(n7393) );
  AND U7109 ( .A(n7404), .B(n7405), .Z(n7403) );
  XOR U7110 ( .A(n7402), .B(n7093), .Z(n7405) );
  XNOR U7111 ( .A(p_input[3276]), .B(n7406), .Z(n7093) );
  AND U7112 ( .A(n222), .B(n7407), .Z(n7406) );
  XOR U7113 ( .A(p_input[3308]), .B(p_input[3276]), .Z(n7407) );
  XNOR U7114 ( .A(n7090), .B(n7402), .Z(n7404) );
  XOR U7115 ( .A(n7408), .B(n7409), .Z(n7090) );
  AND U7116 ( .A(n220), .B(n7410), .Z(n7409) );
  XOR U7117 ( .A(p_input[3244]), .B(p_input[3212]), .Z(n7410) );
  XOR U7118 ( .A(n7411), .B(n7412), .Z(n7402) );
  AND U7119 ( .A(n7413), .B(n7414), .Z(n7412) );
  XOR U7120 ( .A(n7411), .B(n7105), .Z(n7414) );
  XNOR U7121 ( .A(p_input[3275]), .B(n7415), .Z(n7105) );
  AND U7122 ( .A(n222), .B(n7416), .Z(n7415) );
  XOR U7123 ( .A(p_input[3307]), .B(p_input[3275]), .Z(n7416) );
  XNOR U7124 ( .A(n7102), .B(n7411), .Z(n7413) );
  XOR U7125 ( .A(n7417), .B(n7418), .Z(n7102) );
  AND U7126 ( .A(n220), .B(n7419), .Z(n7418) );
  XOR U7127 ( .A(p_input[3243]), .B(p_input[3211]), .Z(n7419) );
  XOR U7128 ( .A(n7420), .B(n7421), .Z(n7411) );
  AND U7129 ( .A(n7422), .B(n7423), .Z(n7421) );
  XOR U7130 ( .A(n7420), .B(n7117), .Z(n7423) );
  XNOR U7131 ( .A(p_input[3274]), .B(n7424), .Z(n7117) );
  AND U7132 ( .A(n222), .B(n7425), .Z(n7424) );
  XOR U7133 ( .A(p_input[3306]), .B(p_input[3274]), .Z(n7425) );
  XNOR U7134 ( .A(n7114), .B(n7420), .Z(n7422) );
  XOR U7135 ( .A(n7426), .B(n7427), .Z(n7114) );
  AND U7136 ( .A(n220), .B(n7428), .Z(n7427) );
  XOR U7137 ( .A(p_input[3242]), .B(p_input[3210]), .Z(n7428) );
  XOR U7138 ( .A(n7429), .B(n7430), .Z(n7420) );
  AND U7139 ( .A(n7431), .B(n7432), .Z(n7430) );
  XOR U7140 ( .A(n7429), .B(n7129), .Z(n7432) );
  XNOR U7141 ( .A(p_input[3273]), .B(n7433), .Z(n7129) );
  AND U7142 ( .A(n222), .B(n7434), .Z(n7433) );
  XOR U7143 ( .A(p_input[3305]), .B(p_input[3273]), .Z(n7434) );
  XNOR U7144 ( .A(n7126), .B(n7429), .Z(n7431) );
  XOR U7145 ( .A(n7435), .B(n7436), .Z(n7126) );
  AND U7146 ( .A(n220), .B(n7437), .Z(n7436) );
  XOR U7147 ( .A(p_input[3241]), .B(p_input[3209]), .Z(n7437) );
  XOR U7148 ( .A(n7438), .B(n7439), .Z(n7429) );
  AND U7149 ( .A(n7440), .B(n7441), .Z(n7439) );
  XOR U7150 ( .A(n7438), .B(n7141), .Z(n7441) );
  XNOR U7151 ( .A(p_input[3272]), .B(n7442), .Z(n7141) );
  AND U7152 ( .A(n222), .B(n7443), .Z(n7442) );
  XOR U7153 ( .A(p_input[3304]), .B(p_input[3272]), .Z(n7443) );
  XNOR U7154 ( .A(n7138), .B(n7438), .Z(n7440) );
  XOR U7155 ( .A(n7444), .B(n7445), .Z(n7138) );
  AND U7156 ( .A(n220), .B(n7446), .Z(n7445) );
  XOR U7157 ( .A(p_input[3240]), .B(p_input[3208]), .Z(n7446) );
  XOR U7158 ( .A(n7447), .B(n7448), .Z(n7438) );
  AND U7159 ( .A(n7449), .B(n7450), .Z(n7448) );
  XOR U7160 ( .A(n7447), .B(n7153), .Z(n7450) );
  XNOR U7161 ( .A(p_input[3271]), .B(n7451), .Z(n7153) );
  AND U7162 ( .A(n222), .B(n7452), .Z(n7451) );
  XOR U7163 ( .A(p_input[3303]), .B(p_input[3271]), .Z(n7452) );
  XNOR U7164 ( .A(n7150), .B(n7447), .Z(n7449) );
  XOR U7165 ( .A(n7453), .B(n7454), .Z(n7150) );
  AND U7166 ( .A(n220), .B(n7455), .Z(n7454) );
  XOR U7167 ( .A(p_input[3239]), .B(p_input[3207]), .Z(n7455) );
  XOR U7168 ( .A(n7456), .B(n7457), .Z(n7447) );
  AND U7169 ( .A(n7458), .B(n7459), .Z(n7457) );
  XOR U7170 ( .A(n7456), .B(n7165), .Z(n7459) );
  XNOR U7171 ( .A(p_input[3270]), .B(n7460), .Z(n7165) );
  AND U7172 ( .A(n222), .B(n7461), .Z(n7460) );
  XOR U7173 ( .A(p_input[3302]), .B(p_input[3270]), .Z(n7461) );
  XNOR U7174 ( .A(n7162), .B(n7456), .Z(n7458) );
  XOR U7175 ( .A(n7462), .B(n7463), .Z(n7162) );
  AND U7176 ( .A(n220), .B(n7464), .Z(n7463) );
  XOR U7177 ( .A(p_input[3238]), .B(p_input[3206]), .Z(n7464) );
  XOR U7178 ( .A(n7465), .B(n7466), .Z(n7456) );
  AND U7179 ( .A(n7467), .B(n7468), .Z(n7466) );
  XOR U7180 ( .A(n7465), .B(n7177), .Z(n7468) );
  XNOR U7181 ( .A(p_input[3269]), .B(n7469), .Z(n7177) );
  AND U7182 ( .A(n222), .B(n7470), .Z(n7469) );
  XOR U7183 ( .A(p_input[3301]), .B(p_input[3269]), .Z(n7470) );
  XNOR U7184 ( .A(n7174), .B(n7465), .Z(n7467) );
  XOR U7185 ( .A(n7471), .B(n7472), .Z(n7174) );
  AND U7186 ( .A(n220), .B(n7473), .Z(n7472) );
  XOR U7187 ( .A(p_input[3237]), .B(p_input[3205]), .Z(n7473) );
  XOR U7188 ( .A(n7474), .B(n7475), .Z(n7465) );
  AND U7189 ( .A(n7476), .B(n7477), .Z(n7475) );
  XOR U7190 ( .A(n7474), .B(n7189), .Z(n7477) );
  XNOR U7191 ( .A(p_input[3268]), .B(n7478), .Z(n7189) );
  AND U7192 ( .A(n222), .B(n7479), .Z(n7478) );
  XOR U7193 ( .A(p_input[3300]), .B(p_input[3268]), .Z(n7479) );
  XNOR U7194 ( .A(n7186), .B(n7474), .Z(n7476) );
  XOR U7195 ( .A(n7480), .B(n7481), .Z(n7186) );
  AND U7196 ( .A(n220), .B(n7482), .Z(n7481) );
  XOR U7197 ( .A(p_input[3236]), .B(p_input[3204]), .Z(n7482) );
  XOR U7198 ( .A(n7483), .B(n7484), .Z(n7474) );
  AND U7199 ( .A(n7485), .B(n7486), .Z(n7484) );
  XOR U7200 ( .A(n7483), .B(n7201), .Z(n7486) );
  XNOR U7201 ( .A(p_input[3267]), .B(n7487), .Z(n7201) );
  AND U7202 ( .A(n222), .B(n7488), .Z(n7487) );
  XOR U7203 ( .A(p_input[3299]), .B(p_input[3267]), .Z(n7488) );
  XNOR U7204 ( .A(n7198), .B(n7483), .Z(n7485) );
  XOR U7205 ( .A(n7489), .B(n7490), .Z(n7198) );
  AND U7206 ( .A(n220), .B(n7491), .Z(n7490) );
  XOR U7207 ( .A(p_input[3235]), .B(p_input[3203]), .Z(n7491) );
  XOR U7208 ( .A(n7492), .B(n7493), .Z(n7483) );
  AND U7209 ( .A(n7494), .B(n7495), .Z(n7493) );
  XOR U7210 ( .A(n7213), .B(n7492), .Z(n7495) );
  XNOR U7211 ( .A(p_input[3266]), .B(n7496), .Z(n7213) );
  AND U7212 ( .A(n222), .B(n7497), .Z(n7496) );
  XOR U7213 ( .A(p_input[3298]), .B(p_input[3266]), .Z(n7497) );
  XNOR U7214 ( .A(n7492), .B(n7210), .Z(n7494) );
  XOR U7215 ( .A(n7498), .B(n7499), .Z(n7210) );
  AND U7216 ( .A(n220), .B(n7500), .Z(n7499) );
  XOR U7217 ( .A(p_input[3234]), .B(p_input[3202]), .Z(n7500) );
  XOR U7218 ( .A(n7501), .B(n7502), .Z(n7492) );
  AND U7219 ( .A(n7503), .B(n7504), .Z(n7502) );
  XNOR U7220 ( .A(n7505), .B(n7226), .Z(n7504) );
  XNOR U7221 ( .A(p_input[3265]), .B(n7506), .Z(n7226) );
  AND U7222 ( .A(n222), .B(n7507), .Z(n7506) );
  XNOR U7223 ( .A(p_input[3297]), .B(n7508), .Z(n7507) );
  IV U7224 ( .A(p_input[3265]), .Z(n7508) );
  XNOR U7225 ( .A(n7223), .B(n7501), .Z(n7503) );
  XNOR U7226 ( .A(p_input[3201]), .B(n7509), .Z(n7223) );
  AND U7227 ( .A(n220), .B(n7510), .Z(n7509) );
  XOR U7228 ( .A(p_input[3233]), .B(p_input[3201]), .Z(n7510) );
  IV U7229 ( .A(n7505), .Z(n7501) );
  AND U7230 ( .A(n7231), .B(n7234), .Z(n7505) );
  XOR U7231 ( .A(p_input[3264]), .B(n7511), .Z(n7234) );
  AND U7232 ( .A(n222), .B(n7512), .Z(n7511) );
  XOR U7233 ( .A(p_input[3296]), .B(p_input[3264]), .Z(n7512) );
  XOR U7234 ( .A(n7513), .B(n7514), .Z(n222) );
  AND U7235 ( .A(n7515), .B(n7516), .Z(n7514) );
  XNOR U7236 ( .A(p_input[3327]), .B(n7513), .Z(n7516) );
  XOR U7237 ( .A(n7513), .B(p_input[3295]), .Z(n7515) );
  XOR U7238 ( .A(n7517), .B(n7518), .Z(n7513) );
  AND U7239 ( .A(n7519), .B(n7520), .Z(n7518) );
  XNOR U7240 ( .A(p_input[3326]), .B(n7517), .Z(n7520) );
  XOR U7241 ( .A(n7517), .B(p_input[3294]), .Z(n7519) );
  XOR U7242 ( .A(n7521), .B(n7522), .Z(n7517) );
  AND U7243 ( .A(n7523), .B(n7524), .Z(n7522) );
  XNOR U7244 ( .A(p_input[3325]), .B(n7521), .Z(n7524) );
  XOR U7245 ( .A(n7521), .B(p_input[3293]), .Z(n7523) );
  XOR U7246 ( .A(n7525), .B(n7526), .Z(n7521) );
  AND U7247 ( .A(n7527), .B(n7528), .Z(n7526) );
  XNOR U7248 ( .A(p_input[3324]), .B(n7525), .Z(n7528) );
  XOR U7249 ( .A(n7525), .B(p_input[3292]), .Z(n7527) );
  XOR U7250 ( .A(n7529), .B(n7530), .Z(n7525) );
  AND U7251 ( .A(n7531), .B(n7532), .Z(n7530) );
  XNOR U7252 ( .A(p_input[3323]), .B(n7529), .Z(n7532) );
  XOR U7253 ( .A(n7529), .B(p_input[3291]), .Z(n7531) );
  XOR U7254 ( .A(n7533), .B(n7534), .Z(n7529) );
  AND U7255 ( .A(n7535), .B(n7536), .Z(n7534) );
  XNOR U7256 ( .A(p_input[3322]), .B(n7533), .Z(n7536) );
  XOR U7257 ( .A(n7533), .B(p_input[3290]), .Z(n7535) );
  XOR U7258 ( .A(n7537), .B(n7538), .Z(n7533) );
  AND U7259 ( .A(n7539), .B(n7540), .Z(n7538) );
  XNOR U7260 ( .A(p_input[3321]), .B(n7537), .Z(n7540) );
  XOR U7261 ( .A(n7537), .B(p_input[3289]), .Z(n7539) );
  XOR U7262 ( .A(n7541), .B(n7542), .Z(n7537) );
  AND U7263 ( .A(n7543), .B(n7544), .Z(n7542) );
  XNOR U7264 ( .A(p_input[3320]), .B(n7541), .Z(n7544) );
  XOR U7265 ( .A(n7541), .B(p_input[3288]), .Z(n7543) );
  XOR U7266 ( .A(n7545), .B(n7546), .Z(n7541) );
  AND U7267 ( .A(n7547), .B(n7548), .Z(n7546) );
  XNOR U7268 ( .A(p_input[3319]), .B(n7545), .Z(n7548) );
  XOR U7269 ( .A(n7545), .B(p_input[3287]), .Z(n7547) );
  XOR U7270 ( .A(n7549), .B(n7550), .Z(n7545) );
  AND U7271 ( .A(n7551), .B(n7552), .Z(n7550) );
  XNOR U7272 ( .A(p_input[3318]), .B(n7549), .Z(n7552) );
  XOR U7273 ( .A(n7549), .B(p_input[3286]), .Z(n7551) );
  XOR U7274 ( .A(n7553), .B(n7554), .Z(n7549) );
  AND U7275 ( .A(n7555), .B(n7556), .Z(n7554) );
  XNOR U7276 ( .A(p_input[3317]), .B(n7553), .Z(n7556) );
  XOR U7277 ( .A(n7553), .B(p_input[3285]), .Z(n7555) );
  XOR U7278 ( .A(n7557), .B(n7558), .Z(n7553) );
  AND U7279 ( .A(n7559), .B(n7560), .Z(n7558) );
  XNOR U7280 ( .A(p_input[3316]), .B(n7557), .Z(n7560) );
  XOR U7281 ( .A(n7557), .B(p_input[3284]), .Z(n7559) );
  XOR U7282 ( .A(n7561), .B(n7562), .Z(n7557) );
  AND U7283 ( .A(n7563), .B(n7564), .Z(n7562) );
  XNOR U7284 ( .A(p_input[3315]), .B(n7561), .Z(n7564) );
  XOR U7285 ( .A(n7561), .B(p_input[3283]), .Z(n7563) );
  XOR U7286 ( .A(n7565), .B(n7566), .Z(n7561) );
  AND U7287 ( .A(n7567), .B(n7568), .Z(n7566) );
  XNOR U7288 ( .A(p_input[3314]), .B(n7565), .Z(n7568) );
  XOR U7289 ( .A(n7565), .B(p_input[3282]), .Z(n7567) );
  XOR U7290 ( .A(n7569), .B(n7570), .Z(n7565) );
  AND U7291 ( .A(n7571), .B(n7572), .Z(n7570) );
  XNOR U7292 ( .A(p_input[3313]), .B(n7569), .Z(n7572) );
  XOR U7293 ( .A(n7569), .B(p_input[3281]), .Z(n7571) );
  XOR U7294 ( .A(n7573), .B(n7574), .Z(n7569) );
  AND U7295 ( .A(n7575), .B(n7576), .Z(n7574) );
  XNOR U7296 ( .A(p_input[3312]), .B(n7573), .Z(n7576) );
  XOR U7297 ( .A(n7573), .B(p_input[3280]), .Z(n7575) );
  XOR U7298 ( .A(n7577), .B(n7578), .Z(n7573) );
  AND U7299 ( .A(n7579), .B(n7580), .Z(n7578) );
  XNOR U7300 ( .A(p_input[3311]), .B(n7577), .Z(n7580) );
  XOR U7301 ( .A(n7577), .B(p_input[3279]), .Z(n7579) );
  XOR U7302 ( .A(n7581), .B(n7582), .Z(n7577) );
  AND U7303 ( .A(n7583), .B(n7584), .Z(n7582) );
  XNOR U7304 ( .A(p_input[3310]), .B(n7581), .Z(n7584) );
  XOR U7305 ( .A(n7581), .B(p_input[3278]), .Z(n7583) );
  XOR U7306 ( .A(n7585), .B(n7586), .Z(n7581) );
  AND U7307 ( .A(n7587), .B(n7588), .Z(n7586) );
  XNOR U7308 ( .A(p_input[3309]), .B(n7585), .Z(n7588) );
  XOR U7309 ( .A(n7585), .B(p_input[3277]), .Z(n7587) );
  XOR U7310 ( .A(n7589), .B(n7590), .Z(n7585) );
  AND U7311 ( .A(n7591), .B(n7592), .Z(n7590) );
  XNOR U7312 ( .A(p_input[3308]), .B(n7589), .Z(n7592) );
  XOR U7313 ( .A(n7589), .B(p_input[3276]), .Z(n7591) );
  XOR U7314 ( .A(n7593), .B(n7594), .Z(n7589) );
  AND U7315 ( .A(n7595), .B(n7596), .Z(n7594) );
  XNOR U7316 ( .A(p_input[3307]), .B(n7593), .Z(n7596) );
  XOR U7317 ( .A(n7593), .B(p_input[3275]), .Z(n7595) );
  XOR U7318 ( .A(n7597), .B(n7598), .Z(n7593) );
  AND U7319 ( .A(n7599), .B(n7600), .Z(n7598) );
  XNOR U7320 ( .A(p_input[3306]), .B(n7597), .Z(n7600) );
  XOR U7321 ( .A(n7597), .B(p_input[3274]), .Z(n7599) );
  XOR U7322 ( .A(n7601), .B(n7602), .Z(n7597) );
  AND U7323 ( .A(n7603), .B(n7604), .Z(n7602) );
  XNOR U7324 ( .A(p_input[3305]), .B(n7601), .Z(n7604) );
  XOR U7325 ( .A(n7601), .B(p_input[3273]), .Z(n7603) );
  XOR U7326 ( .A(n7605), .B(n7606), .Z(n7601) );
  AND U7327 ( .A(n7607), .B(n7608), .Z(n7606) );
  XNOR U7328 ( .A(p_input[3304]), .B(n7605), .Z(n7608) );
  XOR U7329 ( .A(n7605), .B(p_input[3272]), .Z(n7607) );
  XOR U7330 ( .A(n7609), .B(n7610), .Z(n7605) );
  AND U7331 ( .A(n7611), .B(n7612), .Z(n7610) );
  XNOR U7332 ( .A(p_input[3303]), .B(n7609), .Z(n7612) );
  XOR U7333 ( .A(n7609), .B(p_input[3271]), .Z(n7611) );
  XOR U7334 ( .A(n7613), .B(n7614), .Z(n7609) );
  AND U7335 ( .A(n7615), .B(n7616), .Z(n7614) );
  XNOR U7336 ( .A(p_input[3302]), .B(n7613), .Z(n7616) );
  XOR U7337 ( .A(n7613), .B(p_input[3270]), .Z(n7615) );
  XOR U7338 ( .A(n7617), .B(n7618), .Z(n7613) );
  AND U7339 ( .A(n7619), .B(n7620), .Z(n7618) );
  XNOR U7340 ( .A(p_input[3301]), .B(n7617), .Z(n7620) );
  XOR U7341 ( .A(n7617), .B(p_input[3269]), .Z(n7619) );
  XOR U7342 ( .A(n7621), .B(n7622), .Z(n7617) );
  AND U7343 ( .A(n7623), .B(n7624), .Z(n7622) );
  XNOR U7344 ( .A(p_input[3300]), .B(n7621), .Z(n7624) );
  XOR U7345 ( .A(n7621), .B(p_input[3268]), .Z(n7623) );
  XOR U7346 ( .A(n7625), .B(n7626), .Z(n7621) );
  AND U7347 ( .A(n7627), .B(n7628), .Z(n7626) );
  XNOR U7348 ( .A(p_input[3299]), .B(n7625), .Z(n7628) );
  XOR U7349 ( .A(n7625), .B(p_input[3267]), .Z(n7627) );
  XOR U7350 ( .A(n7629), .B(n7630), .Z(n7625) );
  AND U7351 ( .A(n7631), .B(n7632), .Z(n7630) );
  XNOR U7352 ( .A(p_input[3298]), .B(n7629), .Z(n7632) );
  XOR U7353 ( .A(n7629), .B(p_input[3266]), .Z(n7631) );
  XNOR U7354 ( .A(n7633), .B(n7634), .Z(n7629) );
  AND U7355 ( .A(n7635), .B(n7636), .Z(n7634) );
  XOR U7356 ( .A(p_input[3297]), .B(n7633), .Z(n7636) );
  XNOR U7357 ( .A(p_input[3265]), .B(n7633), .Z(n7635) );
  AND U7358 ( .A(p_input[3296]), .B(n7637), .Z(n7633) );
  IV U7359 ( .A(p_input[3264]), .Z(n7637) );
  XNOR U7360 ( .A(p_input[3200]), .B(n7638), .Z(n7231) );
  AND U7361 ( .A(n220), .B(n7639), .Z(n7638) );
  XOR U7362 ( .A(p_input[3232]), .B(p_input[3200]), .Z(n7639) );
  XOR U7363 ( .A(n7640), .B(n7641), .Z(n220) );
  AND U7364 ( .A(n7642), .B(n7643), .Z(n7641) );
  XNOR U7365 ( .A(p_input[3263]), .B(n7640), .Z(n7643) );
  XOR U7366 ( .A(n7640), .B(p_input[3231]), .Z(n7642) );
  XOR U7367 ( .A(n7644), .B(n7645), .Z(n7640) );
  AND U7368 ( .A(n7646), .B(n7647), .Z(n7645) );
  XNOR U7369 ( .A(p_input[3262]), .B(n7644), .Z(n7647) );
  XNOR U7370 ( .A(n7644), .B(n7246), .Z(n7646) );
  IV U7371 ( .A(p_input[3230]), .Z(n7246) );
  XOR U7372 ( .A(n7648), .B(n7649), .Z(n7644) );
  AND U7373 ( .A(n7650), .B(n7651), .Z(n7649) );
  XNOR U7374 ( .A(p_input[3261]), .B(n7648), .Z(n7651) );
  XNOR U7375 ( .A(n7648), .B(n7255), .Z(n7650) );
  IV U7376 ( .A(p_input[3229]), .Z(n7255) );
  XOR U7377 ( .A(n7652), .B(n7653), .Z(n7648) );
  AND U7378 ( .A(n7654), .B(n7655), .Z(n7653) );
  XNOR U7379 ( .A(p_input[3260]), .B(n7652), .Z(n7655) );
  XNOR U7380 ( .A(n7652), .B(n7264), .Z(n7654) );
  IV U7381 ( .A(p_input[3228]), .Z(n7264) );
  XOR U7382 ( .A(n7656), .B(n7657), .Z(n7652) );
  AND U7383 ( .A(n7658), .B(n7659), .Z(n7657) );
  XNOR U7384 ( .A(p_input[3259]), .B(n7656), .Z(n7659) );
  XNOR U7385 ( .A(n7656), .B(n7273), .Z(n7658) );
  IV U7386 ( .A(p_input[3227]), .Z(n7273) );
  XOR U7387 ( .A(n7660), .B(n7661), .Z(n7656) );
  AND U7388 ( .A(n7662), .B(n7663), .Z(n7661) );
  XNOR U7389 ( .A(p_input[3258]), .B(n7660), .Z(n7663) );
  XNOR U7390 ( .A(n7660), .B(n7282), .Z(n7662) );
  IV U7391 ( .A(p_input[3226]), .Z(n7282) );
  XOR U7392 ( .A(n7664), .B(n7665), .Z(n7660) );
  AND U7393 ( .A(n7666), .B(n7667), .Z(n7665) );
  XNOR U7394 ( .A(p_input[3257]), .B(n7664), .Z(n7667) );
  XNOR U7395 ( .A(n7664), .B(n7291), .Z(n7666) );
  IV U7396 ( .A(p_input[3225]), .Z(n7291) );
  XOR U7397 ( .A(n7668), .B(n7669), .Z(n7664) );
  AND U7398 ( .A(n7670), .B(n7671), .Z(n7669) );
  XNOR U7399 ( .A(p_input[3256]), .B(n7668), .Z(n7671) );
  XNOR U7400 ( .A(n7668), .B(n7300), .Z(n7670) );
  IV U7401 ( .A(p_input[3224]), .Z(n7300) );
  XOR U7402 ( .A(n7672), .B(n7673), .Z(n7668) );
  AND U7403 ( .A(n7674), .B(n7675), .Z(n7673) );
  XNOR U7404 ( .A(p_input[3255]), .B(n7672), .Z(n7675) );
  XNOR U7405 ( .A(n7672), .B(n7309), .Z(n7674) );
  IV U7406 ( .A(p_input[3223]), .Z(n7309) );
  XOR U7407 ( .A(n7676), .B(n7677), .Z(n7672) );
  AND U7408 ( .A(n7678), .B(n7679), .Z(n7677) );
  XNOR U7409 ( .A(p_input[3254]), .B(n7676), .Z(n7679) );
  XNOR U7410 ( .A(n7676), .B(n7318), .Z(n7678) );
  IV U7411 ( .A(p_input[3222]), .Z(n7318) );
  XOR U7412 ( .A(n7680), .B(n7681), .Z(n7676) );
  AND U7413 ( .A(n7682), .B(n7683), .Z(n7681) );
  XNOR U7414 ( .A(p_input[3253]), .B(n7680), .Z(n7683) );
  XNOR U7415 ( .A(n7680), .B(n7327), .Z(n7682) );
  IV U7416 ( .A(p_input[3221]), .Z(n7327) );
  XOR U7417 ( .A(n7684), .B(n7685), .Z(n7680) );
  AND U7418 ( .A(n7686), .B(n7687), .Z(n7685) );
  XNOR U7419 ( .A(p_input[3252]), .B(n7684), .Z(n7687) );
  XNOR U7420 ( .A(n7684), .B(n7336), .Z(n7686) );
  IV U7421 ( .A(p_input[3220]), .Z(n7336) );
  XOR U7422 ( .A(n7688), .B(n7689), .Z(n7684) );
  AND U7423 ( .A(n7690), .B(n7691), .Z(n7689) );
  XNOR U7424 ( .A(p_input[3251]), .B(n7688), .Z(n7691) );
  XNOR U7425 ( .A(n7688), .B(n7345), .Z(n7690) );
  IV U7426 ( .A(p_input[3219]), .Z(n7345) );
  XOR U7427 ( .A(n7692), .B(n7693), .Z(n7688) );
  AND U7428 ( .A(n7694), .B(n7695), .Z(n7693) );
  XNOR U7429 ( .A(p_input[3250]), .B(n7692), .Z(n7695) );
  XNOR U7430 ( .A(n7692), .B(n7354), .Z(n7694) );
  IV U7431 ( .A(p_input[3218]), .Z(n7354) );
  XOR U7432 ( .A(n7696), .B(n7697), .Z(n7692) );
  AND U7433 ( .A(n7698), .B(n7699), .Z(n7697) );
  XNOR U7434 ( .A(p_input[3249]), .B(n7696), .Z(n7699) );
  XNOR U7435 ( .A(n7696), .B(n7363), .Z(n7698) );
  IV U7436 ( .A(p_input[3217]), .Z(n7363) );
  XOR U7437 ( .A(n7700), .B(n7701), .Z(n7696) );
  AND U7438 ( .A(n7702), .B(n7703), .Z(n7701) );
  XNOR U7439 ( .A(p_input[3248]), .B(n7700), .Z(n7703) );
  XNOR U7440 ( .A(n7700), .B(n7372), .Z(n7702) );
  IV U7441 ( .A(p_input[3216]), .Z(n7372) );
  XOR U7442 ( .A(n7704), .B(n7705), .Z(n7700) );
  AND U7443 ( .A(n7706), .B(n7707), .Z(n7705) );
  XNOR U7444 ( .A(p_input[3247]), .B(n7704), .Z(n7707) );
  XNOR U7445 ( .A(n7704), .B(n7381), .Z(n7706) );
  IV U7446 ( .A(p_input[3215]), .Z(n7381) );
  XOR U7447 ( .A(n7708), .B(n7709), .Z(n7704) );
  AND U7448 ( .A(n7710), .B(n7711), .Z(n7709) );
  XNOR U7449 ( .A(p_input[3246]), .B(n7708), .Z(n7711) );
  XNOR U7450 ( .A(n7708), .B(n7390), .Z(n7710) );
  IV U7451 ( .A(p_input[3214]), .Z(n7390) );
  XOR U7452 ( .A(n7712), .B(n7713), .Z(n7708) );
  AND U7453 ( .A(n7714), .B(n7715), .Z(n7713) );
  XNOR U7454 ( .A(p_input[3245]), .B(n7712), .Z(n7715) );
  XNOR U7455 ( .A(n7712), .B(n7399), .Z(n7714) );
  IV U7456 ( .A(p_input[3213]), .Z(n7399) );
  XOR U7457 ( .A(n7716), .B(n7717), .Z(n7712) );
  AND U7458 ( .A(n7718), .B(n7719), .Z(n7717) );
  XNOR U7459 ( .A(p_input[3244]), .B(n7716), .Z(n7719) );
  XNOR U7460 ( .A(n7716), .B(n7408), .Z(n7718) );
  IV U7461 ( .A(p_input[3212]), .Z(n7408) );
  XOR U7462 ( .A(n7720), .B(n7721), .Z(n7716) );
  AND U7463 ( .A(n7722), .B(n7723), .Z(n7721) );
  XNOR U7464 ( .A(p_input[3243]), .B(n7720), .Z(n7723) );
  XNOR U7465 ( .A(n7720), .B(n7417), .Z(n7722) );
  IV U7466 ( .A(p_input[3211]), .Z(n7417) );
  XOR U7467 ( .A(n7724), .B(n7725), .Z(n7720) );
  AND U7468 ( .A(n7726), .B(n7727), .Z(n7725) );
  XNOR U7469 ( .A(p_input[3242]), .B(n7724), .Z(n7727) );
  XNOR U7470 ( .A(n7724), .B(n7426), .Z(n7726) );
  IV U7471 ( .A(p_input[3210]), .Z(n7426) );
  XOR U7472 ( .A(n7728), .B(n7729), .Z(n7724) );
  AND U7473 ( .A(n7730), .B(n7731), .Z(n7729) );
  XNOR U7474 ( .A(p_input[3241]), .B(n7728), .Z(n7731) );
  XNOR U7475 ( .A(n7728), .B(n7435), .Z(n7730) );
  IV U7476 ( .A(p_input[3209]), .Z(n7435) );
  XOR U7477 ( .A(n7732), .B(n7733), .Z(n7728) );
  AND U7478 ( .A(n7734), .B(n7735), .Z(n7733) );
  XNOR U7479 ( .A(p_input[3240]), .B(n7732), .Z(n7735) );
  XNOR U7480 ( .A(n7732), .B(n7444), .Z(n7734) );
  IV U7481 ( .A(p_input[3208]), .Z(n7444) );
  XOR U7482 ( .A(n7736), .B(n7737), .Z(n7732) );
  AND U7483 ( .A(n7738), .B(n7739), .Z(n7737) );
  XNOR U7484 ( .A(p_input[3239]), .B(n7736), .Z(n7739) );
  XNOR U7485 ( .A(n7736), .B(n7453), .Z(n7738) );
  IV U7486 ( .A(p_input[3207]), .Z(n7453) );
  XOR U7487 ( .A(n7740), .B(n7741), .Z(n7736) );
  AND U7488 ( .A(n7742), .B(n7743), .Z(n7741) );
  XNOR U7489 ( .A(p_input[3238]), .B(n7740), .Z(n7743) );
  XNOR U7490 ( .A(n7740), .B(n7462), .Z(n7742) );
  IV U7491 ( .A(p_input[3206]), .Z(n7462) );
  XOR U7492 ( .A(n7744), .B(n7745), .Z(n7740) );
  AND U7493 ( .A(n7746), .B(n7747), .Z(n7745) );
  XNOR U7494 ( .A(p_input[3237]), .B(n7744), .Z(n7747) );
  XNOR U7495 ( .A(n7744), .B(n7471), .Z(n7746) );
  IV U7496 ( .A(p_input[3205]), .Z(n7471) );
  XOR U7497 ( .A(n7748), .B(n7749), .Z(n7744) );
  AND U7498 ( .A(n7750), .B(n7751), .Z(n7749) );
  XNOR U7499 ( .A(p_input[3236]), .B(n7748), .Z(n7751) );
  XNOR U7500 ( .A(n7748), .B(n7480), .Z(n7750) );
  IV U7501 ( .A(p_input[3204]), .Z(n7480) );
  XOR U7502 ( .A(n7752), .B(n7753), .Z(n7748) );
  AND U7503 ( .A(n7754), .B(n7755), .Z(n7753) );
  XNOR U7504 ( .A(p_input[3235]), .B(n7752), .Z(n7755) );
  XNOR U7505 ( .A(n7752), .B(n7489), .Z(n7754) );
  IV U7506 ( .A(p_input[3203]), .Z(n7489) );
  XOR U7507 ( .A(n7756), .B(n7757), .Z(n7752) );
  AND U7508 ( .A(n7758), .B(n7759), .Z(n7757) );
  XNOR U7509 ( .A(p_input[3234]), .B(n7756), .Z(n7759) );
  XNOR U7510 ( .A(n7756), .B(n7498), .Z(n7758) );
  IV U7511 ( .A(p_input[3202]), .Z(n7498) );
  XNOR U7512 ( .A(n7760), .B(n7761), .Z(n7756) );
  AND U7513 ( .A(n7762), .B(n7763), .Z(n7761) );
  XOR U7514 ( .A(p_input[3233]), .B(n7760), .Z(n7763) );
  XNOR U7515 ( .A(p_input[3201]), .B(n7760), .Z(n7762) );
  AND U7516 ( .A(p_input[3232]), .B(n7764), .Z(n7760) );
  IV U7517 ( .A(p_input[3200]), .Z(n7764) );
  XOR U7518 ( .A(n7765), .B(n7766), .Z(n6854) );
  AND U7519 ( .A(n319), .B(n7767), .Z(n7766) );
  XNOR U7520 ( .A(n7768), .B(n7765), .Z(n7767) );
  XOR U7521 ( .A(n7769), .B(n7770), .Z(n319) );
  AND U7522 ( .A(n7771), .B(n7772), .Z(n7770) );
  XNOR U7523 ( .A(n6869), .B(n7769), .Z(n7772) );
  AND U7524 ( .A(p_input[3199]), .B(p_input[3167]), .Z(n6869) );
  XNOR U7525 ( .A(n7769), .B(n6866), .Z(n7771) );
  IV U7526 ( .A(n7773), .Z(n6866) );
  AND U7527 ( .A(p_input[3103]), .B(p_input[3135]), .Z(n7773) );
  XOR U7528 ( .A(n7774), .B(n7775), .Z(n7769) );
  AND U7529 ( .A(n7776), .B(n7777), .Z(n7775) );
  XOR U7530 ( .A(n7774), .B(n6881), .Z(n7777) );
  XNOR U7531 ( .A(p_input[3166]), .B(n7778), .Z(n6881) );
  AND U7532 ( .A(n226), .B(n7779), .Z(n7778) );
  XOR U7533 ( .A(p_input[3198]), .B(p_input[3166]), .Z(n7779) );
  XNOR U7534 ( .A(n6878), .B(n7774), .Z(n7776) );
  XOR U7535 ( .A(n7780), .B(n7781), .Z(n6878) );
  AND U7536 ( .A(n223), .B(n7782), .Z(n7781) );
  XOR U7537 ( .A(p_input[3134]), .B(p_input[3102]), .Z(n7782) );
  XOR U7538 ( .A(n7783), .B(n7784), .Z(n7774) );
  AND U7539 ( .A(n7785), .B(n7786), .Z(n7784) );
  XOR U7540 ( .A(n7783), .B(n6893), .Z(n7786) );
  XNOR U7541 ( .A(p_input[3165]), .B(n7787), .Z(n6893) );
  AND U7542 ( .A(n226), .B(n7788), .Z(n7787) );
  XOR U7543 ( .A(p_input[3197]), .B(p_input[3165]), .Z(n7788) );
  XNOR U7544 ( .A(n6890), .B(n7783), .Z(n7785) );
  XOR U7545 ( .A(n7789), .B(n7790), .Z(n6890) );
  AND U7546 ( .A(n223), .B(n7791), .Z(n7790) );
  XOR U7547 ( .A(p_input[3133]), .B(p_input[3101]), .Z(n7791) );
  XOR U7548 ( .A(n7792), .B(n7793), .Z(n7783) );
  AND U7549 ( .A(n7794), .B(n7795), .Z(n7793) );
  XOR U7550 ( .A(n7792), .B(n6905), .Z(n7795) );
  XNOR U7551 ( .A(p_input[3164]), .B(n7796), .Z(n6905) );
  AND U7552 ( .A(n226), .B(n7797), .Z(n7796) );
  XOR U7553 ( .A(p_input[3196]), .B(p_input[3164]), .Z(n7797) );
  XNOR U7554 ( .A(n6902), .B(n7792), .Z(n7794) );
  XOR U7555 ( .A(n7798), .B(n7799), .Z(n6902) );
  AND U7556 ( .A(n223), .B(n7800), .Z(n7799) );
  XOR U7557 ( .A(p_input[3132]), .B(p_input[3100]), .Z(n7800) );
  XOR U7558 ( .A(n7801), .B(n7802), .Z(n7792) );
  AND U7559 ( .A(n7803), .B(n7804), .Z(n7802) );
  XOR U7560 ( .A(n7801), .B(n6917), .Z(n7804) );
  XNOR U7561 ( .A(p_input[3163]), .B(n7805), .Z(n6917) );
  AND U7562 ( .A(n226), .B(n7806), .Z(n7805) );
  XOR U7563 ( .A(p_input[3195]), .B(p_input[3163]), .Z(n7806) );
  XNOR U7564 ( .A(n6914), .B(n7801), .Z(n7803) );
  XOR U7565 ( .A(n7807), .B(n7808), .Z(n6914) );
  AND U7566 ( .A(n223), .B(n7809), .Z(n7808) );
  XOR U7567 ( .A(p_input[3131]), .B(p_input[3099]), .Z(n7809) );
  XOR U7568 ( .A(n7810), .B(n7811), .Z(n7801) );
  AND U7569 ( .A(n7812), .B(n7813), .Z(n7811) );
  XOR U7570 ( .A(n7810), .B(n6929), .Z(n7813) );
  XNOR U7571 ( .A(p_input[3162]), .B(n7814), .Z(n6929) );
  AND U7572 ( .A(n226), .B(n7815), .Z(n7814) );
  XOR U7573 ( .A(p_input[3194]), .B(p_input[3162]), .Z(n7815) );
  XNOR U7574 ( .A(n6926), .B(n7810), .Z(n7812) );
  XOR U7575 ( .A(n7816), .B(n7817), .Z(n6926) );
  AND U7576 ( .A(n223), .B(n7818), .Z(n7817) );
  XOR U7577 ( .A(p_input[3130]), .B(p_input[3098]), .Z(n7818) );
  XOR U7578 ( .A(n7819), .B(n7820), .Z(n7810) );
  AND U7579 ( .A(n7821), .B(n7822), .Z(n7820) );
  XOR U7580 ( .A(n7819), .B(n6941), .Z(n7822) );
  XNOR U7581 ( .A(p_input[3161]), .B(n7823), .Z(n6941) );
  AND U7582 ( .A(n226), .B(n7824), .Z(n7823) );
  XOR U7583 ( .A(p_input[3193]), .B(p_input[3161]), .Z(n7824) );
  XNOR U7584 ( .A(n6938), .B(n7819), .Z(n7821) );
  XOR U7585 ( .A(n7825), .B(n7826), .Z(n6938) );
  AND U7586 ( .A(n223), .B(n7827), .Z(n7826) );
  XOR U7587 ( .A(p_input[3129]), .B(p_input[3097]), .Z(n7827) );
  XOR U7588 ( .A(n7828), .B(n7829), .Z(n7819) );
  AND U7589 ( .A(n7830), .B(n7831), .Z(n7829) );
  XOR U7590 ( .A(n7828), .B(n6953), .Z(n7831) );
  XNOR U7591 ( .A(p_input[3160]), .B(n7832), .Z(n6953) );
  AND U7592 ( .A(n226), .B(n7833), .Z(n7832) );
  XOR U7593 ( .A(p_input[3192]), .B(p_input[3160]), .Z(n7833) );
  XNOR U7594 ( .A(n6950), .B(n7828), .Z(n7830) );
  XOR U7595 ( .A(n7834), .B(n7835), .Z(n6950) );
  AND U7596 ( .A(n223), .B(n7836), .Z(n7835) );
  XOR U7597 ( .A(p_input[3128]), .B(p_input[3096]), .Z(n7836) );
  XOR U7598 ( .A(n7837), .B(n7838), .Z(n7828) );
  AND U7599 ( .A(n7839), .B(n7840), .Z(n7838) );
  XOR U7600 ( .A(n7837), .B(n6965), .Z(n7840) );
  XNOR U7601 ( .A(p_input[3159]), .B(n7841), .Z(n6965) );
  AND U7602 ( .A(n226), .B(n7842), .Z(n7841) );
  XOR U7603 ( .A(p_input[3191]), .B(p_input[3159]), .Z(n7842) );
  XNOR U7604 ( .A(n6962), .B(n7837), .Z(n7839) );
  XOR U7605 ( .A(n7843), .B(n7844), .Z(n6962) );
  AND U7606 ( .A(n223), .B(n7845), .Z(n7844) );
  XOR U7607 ( .A(p_input[3127]), .B(p_input[3095]), .Z(n7845) );
  XOR U7608 ( .A(n7846), .B(n7847), .Z(n7837) );
  AND U7609 ( .A(n7848), .B(n7849), .Z(n7847) );
  XOR U7610 ( .A(n7846), .B(n6977), .Z(n7849) );
  XNOR U7611 ( .A(p_input[3158]), .B(n7850), .Z(n6977) );
  AND U7612 ( .A(n226), .B(n7851), .Z(n7850) );
  XOR U7613 ( .A(p_input[3190]), .B(p_input[3158]), .Z(n7851) );
  XNOR U7614 ( .A(n6974), .B(n7846), .Z(n7848) );
  XOR U7615 ( .A(n7852), .B(n7853), .Z(n6974) );
  AND U7616 ( .A(n223), .B(n7854), .Z(n7853) );
  XOR U7617 ( .A(p_input[3126]), .B(p_input[3094]), .Z(n7854) );
  XOR U7618 ( .A(n7855), .B(n7856), .Z(n7846) );
  AND U7619 ( .A(n7857), .B(n7858), .Z(n7856) );
  XOR U7620 ( .A(n7855), .B(n6989), .Z(n7858) );
  XNOR U7621 ( .A(p_input[3157]), .B(n7859), .Z(n6989) );
  AND U7622 ( .A(n226), .B(n7860), .Z(n7859) );
  XOR U7623 ( .A(p_input[3189]), .B(p_input[3157]), .Z(n7860) );
  XNOR U7624 ( .A(n6986), .B(n7855), .Z(n7857) );
  XOR U7625 ( .A(n7861), .B(n7862), .Z(n6986) );
  AND U7626 ( .A(n223), .B(n7863), .Z(n7862) );
  XOR U7627 ( .A(p_input[3125]), .B(p_input[3093]), .Z(n7863) );
  XOR U7628 ( .A(n7864), .B(n7865), .Z(n7855) );
  AND U7629 ( .A(n7866), .B(n7867), .Z(n7865) );
  XOR U7630 ( .A(n7864), .B(n7001), .Z(n7867) );
  XNOR U7631 ( .A(p_input[3156]), .B(n7868), .Z(n7001) );
  AND U7632 ( .A(n226), .B(n7869), .Z(n7868) );
  XOR U7633 ( .A(p_input[3188]), .B(p_input[3156]), .Z(n7869) );
  XNOR U7634 ( .A(n6998), .B(n7864), .Z(n7866) );
  XOR U7635 ( .A(n7870), .B(n7871), .Z(n6998) );
  AND U7636 ( .A(n223), .B(n7872), .Z(n7871) );
  XOR U7637 ( .A(p_input[3124]), .B(p_input[3092]), .Z(n7872) );
  XOR U7638 ( .A(n7873), .B(n7874), .Z(n7864) );
  AND U7639 ( .A(n7875), .B(n7876), .Z(n7874) );
  XOR U7640 ( .A(n7873), .B(n7013), .Z(n7876) );
  XNOR U7641 ( .A(p_input[3155]), .B(n7877), .Z(n7013) );
  AND U7642 ( .A(n226), .B(n7878), .Z(n7877) );
  XOR U7643 ( .A(p_input[3187]), .B(p_input[3155]), .Z(n7878) );
  XNOR U7644 ( .A(n7010), .B(n7873), .Z(n7875) );
  XOR U7645 ( .A(n7879), .B(n7880), .Z(n7010) );
  AND U7646 ( .A(n223), .B(n7881), .Z(n7880) );
  XOR U7647 ( .A(p_input[3123]), .B(p_input[3091]), .Z(n7881) );
  XOR U7648 ( .A(n7882), .B(n7883), .Z(n7873) );
  AND U7649 ( .A(n7884), .B(n7885), .Z(n7883) );
  XOR U7650 ( .A(n7882), .B(n7025), .Z(n7885) );
  XNOR U7651 ( .A(p_input[3154]), .B(n7886), .Z(n7025) );
  AND U7652 ( .A(n226), .B(n7887), .Z(n7886) );
  XOR U7653 ( .A(p_input[3186]), .B(p_input[3154]), .Z(n7887) );
  XNOR U7654 ( .A(n7022), .B(n7882), .Z(n7884) );
  XOR U7655 ( .A(n7888), .B(n7889), .Z(n7022) );
  AND U7656 ( .A(n223), .B(n7890), .Z(n7889) );
  XOR U7657 ( .A(p_input[3122]), .B(p_input[3090]), .Z(n7890) );
  XOR U7658 ( .A(n7891), .B(n7892), .Z(n7882) );
  AND U7659 ( .A(n7893), .B(n7894), .Z(n7892) );
  XOR U7660 ( .A(n7891), .B(n7037), .Z(n7894) );
  XNOR U7661 ( .A(p_input[3153]), .B(n7895), .Z(n7037) );
  AND U7662 ( .A(n226), .B(n7896), .Z(n7895) );
  XOR U7663 ( .A(p_input[3185]), .B(p_input[3153]), .Z(n7896) );
  XNOR U7664 ( .A(n7034), .B(n7891), .Z(n7893) );
  XOR U7665 ( .A(n7897), .B(n7898), .Z(n7034) );
  AND U7666 ( .A(n223), .B(n7899), .Z(n7898) );
  XOR U7667 ( .A(p_input[3121]), .B(p_input[3089]), .Z(n7899) );
  XOR U7668 ( .A(n7900), .B(n7901), .Z(n7891) );
  AND U7669 ( .A(n7902), .B(n7903), .Z(n7901) );
  XOR U7670 ( .A(n7900), .B(n7049), .Z(n7903) );
  XNOR U7671 ( .A(p_input[3152]), .B(n7904), .Z(n7049) );
  AND U7672 ( .A(n226), .B(n7905), .Z(n7904) );
  XOR U7673 ( .A(p_input[3184]), .B(p_input[3152]), .Z(n7905) );
  XNOR U7674 ( .A(n7046), .B(n7900), .Z(n7902) );
  XOR U7675 ( .A(n7906), .B(n7907), .Z(n7046) );
  AND U7676 ( .A(n223), .B(n7908), .Z(n7907) );
  XOR U7677 ( .A(p_input[3120]), .B(p_input[3088]), .Z(n7908) );
  XOR U7678 ( .A(n7909), .B(n7910), .Z(n7900) );
  AND U7679 ( .A(n7911), .B(n7912), .Z(n7910) );
  XOR U7680 ( .A(n7909), .B(n7061), .Z(n7912) );
  XNOR U7681 ( .A(p_input[3151]), .B(n7913), .Z(n7061) );
  AND U7682 ( .A(n226), .B(n7914), .Z(n7913) );
  XOR U7683 ( .A(p_input[3183]), .B(p_input[3151]), .Z(n7914) );
  XNOR U7684 ( .A(n7058), .B(n7909), .Z(n7911) );
  XOR U7685 ( .A(n7915), .B(n7916), .Z(n7058) );
  AND U7686 ( .A(n223), .B(n7917), .Z(n7916) );
  XOR U7687 ( .A(p_input[3119]), .B(p_input[3087]), .Z(n7917) );
  XOR U7688 ( .A(n7918), .B(n7919), .Z(n7909) );
  AND U7689 ( .A(n7920), .B(n7921), .Z(n7919) );
  XOR U7690 ( .A(n7918), .B(n7073), .Z(n7921) );
  XNOR U7691 ( .A(p_input[3150]), .B(n7922), .Z(n7073) );
  AND U7692 ( .A(n226), .B(n7923), .Z(n7922) );
  XOR U7693 ( .A(p_input[3182]), .B(p_input[3150]), .Z(n7923) );
  XNOR U7694 ( .A(n7070), .B(n7918), .Z(n7920) );
  XOR U7695 ( .A(n7924), .B(n7925), .Z(n7070) );
  AND U7696 ( .A(n223), .B(n7926), .Z(n7925) );
  XOR U7697 ( .A(p_input[3118]), .B(p_input[3086]), .Z(n7926) );
  XOR U7698 ( .A(n7927), .B(n7928), .Z(n7918) );
  AND U7699 ( .A(n7929), .B(n7930), .Z(n7928) );
  XOR U7700 ( .A(n7927), .B(n7085), .Z(n7930) );
  XNOR U7701 ( .A(p_input[3149]), .B(n7931), .Z(n7085) );
  AND U7702 ( .A(n226), .B(n7932), .Z(n7931) );
  XOR U7703 ( .A(p_input[3181]), .B(p_input[3149]), .Z(n7932) );
  XNOR U7704 ( .A(n7082), .B(n7927), .Z(n7929) );
  XOR U7705 ( .A(n7933), .B(n7934), .Z(n7082) );
  AND U7706 ( .A(n223), .B(n7935), .Z(n7934) );
  XOR U7707 ( .A(p_input[3117]), .B(p_input[3085]), .Z(n7935) );
  XOR U7708 ( .A(n7936), .B(n7937), .Z(n7927) );
  AND U7709 ( .A(n7938), .B(n7939), .Z(n7937) );
  XOR U7710 ( .A(n7936), .B(n7097), .Z(n7939) );
  XNOR U7711 ( .A(p_input[3148]), .B(n7940), .Z(n7097) );
  AND U7712 ( .A(n226), .B(n7941), .Z(n7940) );
  XOR U7713 ( .A(p_input[3180]), .B(p_input[3148]), .Z(n7941) );
  XNOR U7714 ( .A(n7094), .B(n7936), .Z(n7938) );
  XOR U7715 ( .A(n7942), .B(n7943), .Z(n7094) );
  AND U7716 ( .A(n223), .B(n7944), .Z(n7943) );
  XOR U7717 ( .A(p_input[3116]), .B(p_input[3084]), .Z(n7944) );
  XOR U7718 ( .A(n7945), .B(n7946), .Z(n7936) );
  AND U7719 ( .A(n7947), .B(n7948), .Z(n7946) );
  XOR U7720 ( .A(n7945), .B(n7109), .Z(n7948) );
  XNOR U7721 ( .A(p_input[3147]), .B(n7949), .Z(n7109) );
  AND U7722 ( .A(n226), .B(n7950), .Z(n7949) );
  XOR U7723 ( .A(p_input[3179]), .B(p_input[3147]), .Z(n7950) );
  XNOR U7724 ( .A(n7106), .B(n7945), .Z(n7947) );
  XOR U7725 ( .A(n7951), .B(n7952), .Z(n7106) );
  AND U7726 ( .A(n223), .B(n7953), .Z(n7952) );
  XOR U7727 ( .A(p_input[3115]), .B(p_input[3083]), .Z(n7953) );
  XOR U7728 ( .A(n7954), .B(n7955), .Z(n7945) );
  AND U7729 ( .A(n7956), .B(n7957), .Z(n7955) );
  XOR U7730 ( .A(n7954), .B(n7121), .Z(n7957) );
  XNOR U7731 ( .A(p_input[3146]), .B(n7958), .Z(n7121) );
  AND U7732 ( .A(n226), .B(n7959), .Z(n7958) );
  XOR U7733 ( .A(p_input[3178]), .B(p_input[3146]), .Z(n7959) );
  XNOR U7734 ( .A(n7118), .B(n7954), .Z(n7956) );
  XOR U7735 ( .A(n7960), .B(n7961), .Z(n7118) );
  AND U7736 ( .A(n223), .B(n7962), .Z(n7961) );
  XOR U7737 ( .A(p_input[3114]), .B(p_input[3082]), .Z(n7962) );
  XOR U7738 ( .A(n7963), .B(n7964), .Z(n7954) );
  AND U7739 ( .A(n7965), .B(n7966), .Z(n7964) );
  XOR U7740 ( .A(n7963), .B(n7133), .Z(n7966) );
  XNOR U7741 ( .A(p_input[3145]), .B(n7967), .Z(n7133) );
  AND U7742 ( .A(n226), .B(n7968), .Z(n7967) );
  XOR U7743 ( .A(p_input[3177]), .B(p_input[3145]), .Z(n7968) );
  XNOR U7744 ( .A(n7130), .B(n7963), .Z(n7965) );
  XOR U7745 ( .A(n7969), .B(n7970), .Z(n7130) );
  AND U7746 ( .A(n223), .B(n7971), .Z(n7970) );
  XOR U7747 ( .A(p_input[3113]), .B(p_input[3081]), .Z(n7971) );
  XOR U7748 ( .A(n7972), .B(n7973), .Z(n7963) );
  AND U7749 ( .A(n7974), .B(n7975), .Z(n7973) );
  XOR U7750 ( .A(n7972), .B(n7145), .Z(n7975) );
  XNOR U7751 ( .A(p_input[3144]), .B(n7976), .Z(n7145) );
  AND U7752 ( .A(n226), .B(n7977), .Z(n7976) );
  XOR U7753 ( .A(p_input[3176]), .B(p_input[3144]), .Z(n7977) );
  XNOR U7754 ( .A(n7142), .B(n7972), .Z(n7974) );
  XOR U7755 ( .A(n7978), .B(n7979), .Z(n7142) );
  AND U7756 ( .A(n223), .B(n7980), .Z(n7979) );
  XOR U7757 ( .A(p_input[3112]), .B(p_input[3080]), .Z(n7980) );
  XOR U7758 ( .A(n7981), .B(n7982), .Z(n7972) );
  AND U7759 ( .A(n7983), .B(n7984), .Z(n7982) );
  XOR U7760 ( .A(n7981), .B(n7157), .Z(n7984) );
  XNOR U7761 ( .A(p_input[3143]), .B(n7985), .Z(n7157) );
  AND U7762 ( .A(n226), .B(n7986), .Z(n7985) );
  XOR U7763 ( .A(p_input[3175]), .B(p_input[3143]), .Z(n7986) );
  XNOR U7764 ( .A(n7154), .B(n7981), .Z(n7983) );
  XOR U7765 ( .A(n7987), .B(n7988), .Z(n7154) );
  AND U7766 ( .A(n223), .B(n7989), .Z(n7988) );
  XOR U7767 ( .A(p_input[3111]), .B(p_input[3079]), .Z(n7989) );
  XOR U7768 ( .A(n7990), .B(n7991), .Z(n7981) );
  AND U7769 ( .A(n7992), .B(n7993), .Z(n7991) );
  XOR U7770 ( .A(n7990), .B(n7169), .Z(n7993) );
  XNOR U7771 ( .A(p_input[3142]), .B(n7994), .Z(n7169) );
  AND U7772 ( .A(n226), .B(n7995), .Z(n7994) );
  XOR U7773 ( .A(p_input[3174]), .B(p_input[3142]), .Z(n7995) );
  XNOR U7774 ( .A(n7166), .B(n7990), .Z(n7992) );
  XOR U7775 ( .A(n7996), .B(n7997), .Z(n7166) );
  AND U7776 ( .A(n223), .B(n7998), .Z(n7997) );
  XOR U7777 ( .A(p_input[3110]), .B(p_input[3078]), .Z(n7998) );
  XOR U7778 ( .A(n7999), .B(n8000), .Z(n7990) );
  AND U7779 ( .A(n8001), .B(n8002), .Z(n8000) );
  XOR U7780 ( .A(n7999), .B(n7181), .Z(n8002) );
  XNOR U7781 ( .A(p_input[3141]), .B(n8003), .Z(n7181) );
  AND U7782 ( .A(n226), .B(n8004), .Z(n8003) );
  XOR U7783 ( .A(p_input[3173]), .B(p_input[3141]), .Z(n8004) );
  XNOR U7784 ( .A(n7178), .B(n7999), .Z(n8001) );
  XOR U7785 ( .A(n8005), .B(n8006), .Z(n7178) );
  AND U7786 ( .A(n223), .B(n8007), .Z(n8006) );
  XOR U7787 ( .A(p_input[3109]), .B(p_input[3077]), .Z(n8007) );
  XOR U7788 ( .A(n8008), .B(n8009), .Z(n7999) );
  AND U7789 ( .A(n8010), .B(n8011), .Z(n8009) );
  XOR U7790 ( .A(n8008), .B(n7193), .Z(n8011) );
  XNOR U7791 ( .A(p_input[3140]), .B(n8012), .Z(n7193) );
  AND U7792 ( .A(n226), .B(n8013), .Z(n8012) );
  XOR U7793 ( .A(p_input[3172]), .B(p_input[3140]), .Z(n8013) );
  XNOR U7794 ( .A(n7190), .B(n8008), .Z(n8010) );
  XOR U7795 ( .A(n8014), .B(n8015), .Z(n7190) );
  AND U7796 ( .A(n223), .B(n8016), .Z(n8015) );
  XOR U7797 ( .A(p_input[3108]), .B(p_input[3076]), .Z(n8016) );
  XOR U7798 ( .A(n8017), .B(n8018), .Z(n8008) );
  AND U7799 ( .A(n8019), .B(n8020), .Z(n8018) );
  XOR U7800 ( .A(n8017), .B(n7205), .Z(n8020) );
  XNOR U7801 ( .A(p_input[3139]), .B(n8021), .Z(n7205) );
  AND U7802 ( .A(n226), .B(n8022), .Z(n8021) );
  XOR U7803 ( .A(p_input[3171]), .B(p_input[3139]), .Z(n8022) );
  XNOR U7804 ( .A(n7202), .B(n8017), .Z(n8019) );
  XOR U7805 ( .A(n8023), .B(n8024), .Z(n7202) );
  AND U7806 ( .A(n223), .B(n8025), .Z(n8024) );
  XOR U7807 ( .A(p_input[3107]), .B(p_input[3075]), .Z(n8025) );
  XOR U7808 ( .A(n8026), .B(n8027), .Z(n8017) );
  AND U7809 ( .A(n8028), .B(n8029), .Z(n8027) );
  XOR U7810 ( .A(n7217), .B(n8026), .Z(n8029) );
  XNOR U7811 ( .A(p_input[3138]), .B(n8030), .Z(n7217) );
  AND U7812 ( .A(n226), .B(n8031), .Z(n8030) );
  XOR U7813 ( .A(p_input[3170]), .B(p_input[3138]), .Z(n8031) );
  XNOR U7814 ( .A(n8026), .B(n7214), .Z(n8028) );
  XOR U7815 ( .A(n8032), .B(n8033), .Z(n7214) );
  AND U7816 ( .A(n223), .B(n8034), .Z(n8033) );
  XOR U7817 ( .A(p_input[3106]), .B(p_input[3074]), .Z(n8034) );
  XOR U7818 ( .A(n8035), .B(n8036), .Z(n8026) );
  AND U7819 ( .A(n8037), .B(n8038), .Z(n8036) );
  XNOR U7820 ( .A(n8039), .B(n7230), .Z(n8038) );
  XNOR U7821 ( .A(p_input[3137]), .B(n8040), .Z(n7230) );
  AND U7822 ( .A(n226), .B(n8041), .Z(n8040) );
  XNOR U7823 ( .A(p_input[3169]), .B(n8042), .Z(n8041) );
  IV U7824 ( .A(p_input[3137]), .Z(n8042) );
  XNOR U7825 ( .A(n7227), .B(n8035), .Z(n8037) );
  XNOR U7826 ( .A(p_input[3073]), .B(n8043), .Z(n7227) );
  AND U7827 ( .A(n223), .B(n8044), .Z(n8043) );
  XOR U7828 ( .A(p_input[3105]), .B(p_input[3073]), .Z(n8044) );
  IV U7829 ( .A(n8039), .Z(n8035) );
  AND U7830 ( .A(n7765), .B(n7768), .Z(n8039) );
  XOR U7831 ( .A(p_input[3136]), .B(n8045), .Z(n7768) );
  AND U7832 ( .A(n226), .B(n8046), .Z(n8045) );
  XOR U7833 ( .A(p_input[3168]), .B(p_input[3136]), .Z(n8046) );
  XOR U7834 ( .A(n8047), .B(n8048), .Z(n226) );
  AND U7835 ( .A(n8049), .B(n8050), .Z(n8048) );
  XNOR U7836 ( .A(p_input[3199]), .B(n8047), .Z(n8050) );
  XOR U7837 ( .A(n8047), .B(p_input[3167]), .Z(n8049) );
  XOR U7838 ( .A(n8051), .B(n8052), .Z(n8047) );
  AND U7839 ( .A(n8053), .B(n8054), .Z(n8052) );
  XNOR U7840 ( .A(p_input[3198]), .B(n8051), .Z(n8054) );
  XOR U7841 ( .A(n8051), .B(p_input[3166]), .Z(n8053) );
  XOR U7842 ( .A(n8055), .B(n8056), .Z(n8051) );
  AND U7843 ( .A(n8057), .B(n8058), .Z(n8056) );
  XNOR U7844 ( .A(p_input[3197]), .B(n8055), .Z(n8058) );
  XOR U7845 ( .A(n8055), .B(p_input[3165]), .Z(n8057) );
  XOR U7846 ( .A(n8059), .B(n8060), .Z(n8055) );
  AND U7847 ( .A(n8061), .B(n8062), .Z(n8060) );
  XNOR U7848 ( .A(p_input[3196]), .B(n8059), .Z(n8062) );
  XOR U7849 ( .A(n8059), .B(p_input[3164]), .Z(n8061) );
  XOR U7850 ( .A(n8063), .B(n8064), .Z(n8059) );
  AND U7851 ( .A(n8065), .B(n8066), .Z(n8064) );
  XNOR U7852 ( .A(p_input[3195]), .B(n8063), .Z(n8066) );
  XOR U7853 ( .A(n8063), .B(p_input[3163]), .Z(n8065) );
  XOR U7854 ( .A(n8067), .B(n8068), .Z(n8063) );
  AND U7855 ( .A(n8069), .B(n8070), .Z(n8068) );
  XNOR U7856 ( .A(p_input[3194]), .B(n8067), .Z(n8070) );
  XOR U7857 ( .A(n8067), .B(p_input[3162]), .Z(n8069) );
  XOR U7858 ( .A(n8071), .B(n8072), .Z(n8067) );
  AND U7859 ( .A(n8073), .B(n8074), .Z(n8072) );
  XNOR U7860 ( .A(p_input[3193]), .B(n8071), .Z(n8074) );
  XOR U7861 ( .A(n8071), .B(p_input[3161]), .Z(n8073) );
  XOR U7862 ( .A(n8075), .B(n8076), .Z(n8071) );
  AND U7863 ( .A(n8077), .B(n8078), .Z(n8076) );
  XNOR U7864 ( .A(p_input[3192]), .B(n8075), .Z(n8078) );
  XOR U7865 ( .A(n8075), .B(p_input[3160]), .Z(n8077) );
  XOR U7866 ( .A(n8079), .B(n8080), .Z(n8075) );
  AND U7867 ( .A(n8081), .B(n8082), .Z(n8080) );
  XNOR U7868 ( .A(p_input[3191]), .B(n8079), .Z(n8082) );
  XOR U7869 ( .A(n8079), .B(p_input[3159]), .Z(n8081) );
  XOR U7870 ( .A(n8083), .B(n8084), .Z(n8079) );
  AND U7871 ( .A(n8085), .B(n8086), .Z(n8084) );
  XNOR U7872 ( .A(p_input[3190]), .B(n8083), .Z(n8086) );
  XOR U7873 ( .A(n8083), .B(p_input[3158]), .Z(n8085) );
  XOR U7874 ( .A(n8087), .B(n8088), .Z(n8083) );
  AND U7875 ( .A(n8089), .B(n8090), .Z(n8088) );
  XNOR U7876 ( .A(p_input[3189]), .B(n8087), .Z(n8090) );
  XOR U7877 ( .A(n8087), .B(p_input[3157]), .Z(n8089) );
  XOR U7878 ( .A(n8091), .B(n8092), .Z(n8087) );
  AND U7879 ( .A(n8093), .B(n8094), .Z(n8092) );
  XNOR U7880 ( .A(p_input[3188]), .B(n8091), .Z(n8094) );
  XOR U7881 ( .A(n8091), .B(p_input[3156]), .Z(n8093) );
  XOR U7882 ( .A(n8095), .B(n8096), .Z(n8091) );
  AND U7883 ( .A(n8097), .B(n8098), .Z(n8096) );
  XNOR U7884 ( .A(p_input[3187]), .B(n8095), .Z(n8098) );
  XOR U7885 ( .A(n8095), .B(p_input[3155]), .Z(n8097) );
  XOR U7886 ( .A(n8099), .B(n8100), .Z(n8095) );
  AND U7887 ( .A(n8101), .B(n8102), .Z(n8100) );
  XNOR U7888 ( .A(p_input[3186]), .B(n8099), .Z(n8102) );
  XOR U7889 ( .A(n8099), .B(p_input[3154]), .Z(n8101) );
  XOR U7890 ( .A(n8103), .B(n8104), .Z(n8099) );
  AND U7891 ( .A(n8105), .B(n8106), .Z(n8104) );
  XNOR U7892 ( .A(p_input[3185]), .B(n8103), .Z(n8106) );
  XOR U7893 ( .A(n8103), .B(p_input[3153]), .Z(n8105) );
  XOR U7894 ( .A(n8107), .B(n8108), .Z(n8103) );
  AND U7895 ( .A(n8109), .B(n8110), .Z(n8108) );
  XNOR U7896 ( .A(p_input[3184]), .B(n8107), .Z(n8110) );
  XOR U7897 ( .A(n8107), .B(p_input[3152]), .Z(n8109) );
  XOR U7898 ( .A(n8111), .B(n8112), .Z(n8107) );
  AND U7899 ( .A(n8113), .B(n8114), .Z(n8112) );
  XNOR U7900 ( .A(p_input[3183]), .B(n8111), .Z(n8114) );
  XOR U7901 ( .A(n8111), .B(p_input[3151]), .Z(n8113) );
  XOR U7902 ( .A(n8115), .B(n8116), .Z(n8111) );
  AND U7903 ( .A(n8117), .B(n8118), .Z(n8116) );
  XNOR U7904 ( .A(p_input[3182]), .B(n8115), .Z(n8118) );
  XOR U7905 ( .A(n8115), .B(p_input[3150]), .Z(n8117) );
  XOR U7906 ( .A(n8119), .B(n8120), .Z(n8115) );
  AND U7907 ( .A(n8121), .B(n8122), .Z(n8120) );
  XNOR U7908 ( .A(p_input[3181]), .B(n8119), .Z(n8122) );
  XOR U7909 ( .A(n8119), .B(p_input[3149]), .Z(n8121) );
  XOR U7910 ( .A(n8123), .B(n8124), .Z(n8119) );
  AND U7911 ( .A(n8125), .B(n8126), .Z(n8124) );
  XNOR U7912 ( .A(p_input[3180]), .B(n8123), .Z(n8126) );
  XOR U7913 ( .A(n8123), .B(p_input[3148]), .Z(n8125) );
  XOR U7914 ( .A(n8127), .B(n8128), .Z(n8123) );
  AND U7915 ( .A(n8129), .B(n8130), .Z(n8128) );
  XNOR U7916 ( .A(p_input[3179]), .B(n8127), .Z(n8130) );
  XOR U7917 ( .A(n8127), .B(p_input[3147]), .Z(n8129) );
  XOR U7918 ( .A(n8131), .B(n8132), .Z(n8127) );
  AND U7919 ( .A(n8133), .B(n8134), .Z(n8132) );
  XNOR U7920 ( .A(p_input[3178]), .B(n8131), .Z(n8134) );
  XOR U7921 ( .A(n8131), .B(p_input[3146]), .Z(n8133) );
  XOR U7922 ( .A(n8135), .B(n8136), .Z(n8131) );
  AND U7923 ( .A(n8137), .B(n8138), .Z(n8136) );
  XNOR U7924 ( .A(p_input[3177]), .B(n8135), .Z(n8138) );
  XOR U7925 ( .A(n8135), .B(p_input[3145]), .Z(n8137) );
  XOR U7926 ( .A(n8139), .B(n8140), .Z(n8135) );
  AND U7927 ( .A(n8141), .B(n8142), .Z(n8140) );
  XNOR U7928 ( .A(p_input[3176]), .B(n8139), .Z(n8142) );
  XOR U7929 ( .A(n8139), .B(p_input[3144]), .Z(n8141) );
  XOR U7930 ( .A(n8143), .B(n8144), .Z(n8139) );
  AND U7931 ( .A(n8145), .B(n8146), .Z(n8144) );
  XNOR U7932 ( .A(p_input[3175]), .B(n8143), .Z(n8146) );
  XOR U7933 ( .A(n8143), .B(p_input[3143]), .Z(n8145) );
  XOR U7934 ( .A(n8147), .B(n8148), .Z(n8143) );
  AND U7935 ( .A(n8149), .B(n8150), .Z(n8148) );
  XNOR U7936 ( .A(p_input[3174]), .B(n8147), .Z(n8150) );
  XOR U7937 ( .A(n8147), .B(p_input[3142]), .Z(n8149) );
  XOR U7938 ( .A(n8151), .B(n8152), .Z(n8147) );
  AND U7939 ( .A(n8153), .B(n8154), .Z(n8152) );
  XNOR U7940 ( .A(p_input[3173]), .B(n8151), .Z(n8154) );
  XOR U7941 ( .A(n8151), .B(p_input[3141]), .Z(n8153) );
  XOR U7942 ( .A(n8155), .B(n8156), .Z(n8151) );
  AND U7943 ( .A(n8157), .B(n8158), .Z(n8156) );
  XNOR U7944 ( .A(p_input[3172]), .B(n8155), .Z(n8158) );
  XOR U7945 ( .A(n8155), .B(p_input[3140]), .Z(n8157) );
  XOR U7946 ( .A(n8159), .B(n8160), .Z(n8155) );
  AND U7947 ( .A(n8161), .B(n8162), .Z(n8160) );
  XNOR U7948 ( .A(p_input[3171]), .B(n8159), .Z(n8162) );
  XOR U7949 ( .A(n8159), .B(p_input[3139]), .Z(n8161) );
  XOR U7950 ( .A(n8163), .B(n8164), .Z(n8159) );
  AND U7951 ( .A(n8165), .B(n8166), .Z(n8164) );
  XNOR U7952 ( .A(p_input[3170]), .B(n8163), .Z(n8166) );
  XOR U7953 ( .A(n8163), .B(p_input[3138]), .Z(n8165) );
  XNOR U7954 ( .A(n8167), .B(n8168), .Z(n8163) );
  AND U7955 ( .A(n8169), .B(n8170), .Z(n8168) );
  XOR U7956 ( .A(p_input[3169]), .B(n8167), .Z(n8170) );
  XNOR U7957 ( .A(p_input[3137]), .B(n8167), .Z(n8169) );
  AND U7958 ( .A(p_input[3168]), .B(n8171), .Z(n8167) );
  IV U7959 ( .A(p_input[3136]), .Z(n8171) );
  XNOR U7960 ( .A(p_input[3072]), .B(n8172), .Z(n7765) );
  AND U7961 ( .A(n223), .B(n8173), .Z(n8172) );
  XOR U7962 ( .A(p_input[3104]), .B(p_input[3072]), .Z(n8173) );
  XOR U7963 ( .A(n8174), .B(n8175), .Z(n223) );
  AND U7964 ( .A(n8176), .B(n8177), .Z(n8175) );
  XNOR U7965 ( .A(p_input[3135]), .B(n8174), .Z(n8177) );
  XOR U7966 ( .A(n8174), .B(p_input[3103]), .Z(n8176) );
  XOR U7967 ( .A(n8178), .B(n8179), .Z(n8174) );
  AND U7968 ( .A(n8180), .B(n8181), .Z(n8179) );
  XNOR U7969 ( .A(p_input[3134]), .B(n8178), .Z(n8181) );
  XNOR U7970 ( .A(n8178), .B(n7780), .Z(n8180) );
  IV U7971 ( .A(p_input[3102]), .Z(n7780) );
  XOR U7972 ( .A(n8182), .B(n8183), .Z(n8178) );
  AND U7973 ( .A(n8184), .B(n8185), .Z(n8183) );
  XNOR U7974 ( .A(p_input[3133]), .B(n8182), .Z(n8185) );
  XNOR U7975 ( .A(n8182), .B(n7789), .Z(n8184) );
  IV U7976 ( .A(p_input[3101]), .Z(n7789) );
  XOR U7977 ( .A(n8186), .B(n8187), .Z(n8182) );
  AND U7978 ( .A(n8188), .B(n8189), .Z(n8187) );
  XNOR U7979 ( .A(p_input[3132]), .B(n8186), .Z(n8189) );
  XNOR U7980 ( .A(n8186), .B(n7798), .Z(n8188) );
  IV U7981 ( .A(p_input[3100]), .Z(n7798) );
  XOR U7982 ( .A(n8190), .B(n8191), .Z(n8186) );
  AND U7983 ( .A(n8192), .B(n8193), .Z(n8191) );
  XNOR U7984 ( .A(p_input[3131]), .B(n8190), .Z(n8193) );
  XNOR U7985 ( .A(n8190), .B(n7807), .Z(n8192) );
  IV U7986 ( .A(p_input[3099]), .Z(n7807) );
  XOR U7987 ( .A(n8194), .B(n8195), .Z(n8190) );
  AND U7988 ( .A(n8196), .B(n8197), .Z(n8195) );
  XNOR U7989 ( .A(p_input[3130]), .B(n8194), .Z(n8197) );
  XNOR U7990 ( .A(n8194), .B(n7816), .Z(n8196) );
  IV U7991 ( .A(p_input[3098]), .Z(n7816) );
  XOR U7992 ( .A(n8198), .B(n8199), .Z(n8194) );
  AND U7993 ( .A(n8200), .B(n8201), .Z(n8199) );
  XNOR U7994 ( .A(p_input[3129]), .B(n8198), .Z(n8201) );
  XNOR U7995 ( .A(n8198), .B(n7825), .Z(n8200) );
  IV U7996 ( .A(p_input[3097]), .Z(n7825) );
  XOR U7997 ( .A(n8202), .B(n8203), .Z(n8198) );
  AND U7998 ( .A(n8204), .B(n8205), .Z(n8203) );
  XNOR U7999 ( .A(p_input[3128]), .B(n8202), .Z(n8205) );
  XNOR U8000 ( .A(n8202), .B(n7834), .Z(n8204) );
  IV U8001 ( .A(p_input[3096]), .Z(n7834) );
  XOR U8002 ( .A(n8206), .B(n8207), .Z(n8202) );
  AND U8003 ( .A(n8208), .B(n8209), .Z(n8207) );
  XNOR U8004 ( .A(p_input[3127]), .B(n8206), .Z(n8209) );
  XNOR U8005 ( .A(n8206), .B(n7843), .Z(n8208) );
  IV U8006 ( .A(p_input[3095]), .Z(n7843) );
  XOR U8007 ( .A(n8210), .B(n8211), .Z(n8206) );
  AND U8008 ( .A(n8212), .B(n8213), .Z(n8211) );
  XNOR U8009 ( .A(p_input[3126]), .B(n8210), .Z(n8213) );
  XNOR U8010 ( .A(n8210), .B(n7852), .Z(n8212) );
  IV U8011 ( .A(p_input[3094]), .Z(n7852) );
  XOR U8012 ( .A(n8214), .B(n8215), .Z(n8210) );
  AND U8013 ( .A(n8216), .B(n8217), .Z(n8215) );
  XNOR U8014 ( .A(p_input[3125]), .B(n8214), .Z(n8217) );
  XNOR U8015 ( .A(n8214), .B(n7861), .Z(n8216) );
  IV U8016 ( .A(p_input[3093]), .Z(n7861) );
  XOR U8017 ( .A(n8218), .B(n8219), .Z(n8214) );
  AND U8018 ( .A(n8220), .B(n8221), .Z(n8219) );
  XNOR U8019 ( .A(p_input[3124]), .B(n8218), .Z(n8221) );
  XNOR U8020 ( .A(n8218), .B(n7870), .Z(n8220) );
  IV U8021 ( .A(p_input[3092]), .Z(n7870) );
  XOR U8022 ( .A(n8222), .B(n8223), .Z(n8218) );
  AND U8023 ( .A(n8224), .B(n8225), .Z(n8223) );
  XNOR U8024 ( .A(p_input[3123]), .B(n8222), .Z(n8225) );
  XNOR U8025 ( .A(n8222), .B(n7879), .Z(n8224) );
  IV U8026 ( .A(p_input[3091]), .Z(n7879) );
  XOR U8027 ( .A(n8226), .B(n8227), .Z(n8222) );
  AND U8028 ( .A(n8228), .B(n8229), .Z(n8227) );
  XNOR U8029 ( .A(p_input[3122]), .B(n8226), .Z(n8229) );
  XNOR U8030 ( .A(n8226), .B(n7888), .Z(n8228) );
  IV U8031 ( .A(p_input[3090]), .Z(n7888) );
  XOR U8032 ( .A(n8230), .B(n8231), .Z(n8226) );
  AND U8033 ( .A(n8232), .B(n8233), .Z(n8231) );
  XNOR U8034 ( .A(p_input[3121]), .B(n8230), .Z(n8233) );
  XNOR U8035 ( .A(n8230), .B(n7897), .Z(n8232) );
  IV U8036 ( .A(p_input[3089]), .Z(n7897) );
  XOR U8037 ( .A(n8234), .B(n8235), .Z(n8230) );
  AND U8038 ( .A(n8236), .B(n8237), .Z(n8235) );
  XNOR U8039 ( .A(p_input[3120]), .B(n8234), .Z(n8237) );
  XNOR U8040 ( .A(n8234), .B(n7906), .Z(n8236) );
  IV U8041 ( .A(p_input[3088]), .Z(n7906) );
  XOR U8042 ( .A(n8238), .B(n8239), .Z(n8234) );
  AND U8043 ( .A(n8240), .B(n8241), .Z(n8239) );
  XNOR U8044 ( .A(p_input[3119]), .B(n8238), .Z(n8241) );
  XNOR U8045 ( .A(n8238), .B(n7915), .Z(n8240) );
  IV U8046 ( .A(p_input[3087]), .Z(n7915) );
  XOR U8047 ( .A(n8242), .B(n8243), .Z(n8238) );
  AND U8048 ( .A(n8244), .B(n8245), .Z(n8243) );
  XNOR U8049 ( .A(p_input[3118]), .B(n8242), .Z(n8245) );
  XNOR U8050 ( .A(n8242), .B(n7924), .Z(n8244) );
  IV U8051 ( .A(p_input[3086]), .Z(n7924) );
  XOR U8052 ( .A(n8246), .B(n8247), .Z(n8242) );
  AND U8053 ( .A(n8248), .B(n8249), .Z(n8247) );
  XNOR U8054 ( .A(p_input[3117]), .B(n8246), .Z(n8249) );
  XNOR U8055 ( .A(n8246), .B(n7933), .Z(n8248) );
  IV U8056 ( .A(p_input[3085]), .Z(n7933) );
  XOR U8057 ( .A(n8250), .B(n8251), .Z(n8246) );
  AND U8058 ( .A(n8252), .B(n8253), .Z(n8251) );
  XNOR U8059 ( .A(p_input[3116]), .B(n8250), .Z(n8253) );
  XNOR U8060 ( .A(n8250), .B(n7942), .Z(n8252) );
  IV U8061 ( .A(p_input[3084]), .Z(n7942) );
  XOR U8062 ( .A(n8254), .B(n8255), .Z(n8250) );
  AND U8063 ( .A(n8256), .B(n8257), .Z(n8255) );
  XNOR U8064 ( .A(p_input[3115]), .B(n8254), .Z(n8257) );
  XNOR U8065 ( .A(n8254), .B(n7951), .Z(n8256) );
  IV U8066 ( .A(p_input[3083]), .Z(n7951) );
  XOR U8067 ( .A(n8258), .B(n8259), .Z(n8254) );
  AND U8068 ( .A(n8260), .B(n8261), .Z(n8259) );
  XNOR U8069 ( .A(p_input[3114]), .B(n8258), .Z(n8261) );
  XNOR U8070 ( .A(n8258), .B(n7960), .Z(n8260) );
  IV U8071 ( .A(p_input[3082]), .Z(n7960) );
  XOR U8072 ( .A(n8262), .B(n8263), .Z(n8258) );
  AND U8073 ( .A(n8264), .B(n8265), .Z(n8263) );
  XNOR U8074 ( .A(p_input[3113]), .B(n8262), .Z(n8265) );
  XNOR U8075 ( .A(n8262), .B(n7969), .Z(n8264) );
  IV U8076 ( .A(p_input[3081]), .Z(n7969) );
  XOR U8077 ( .A(n8266), .B(n8267), .Z(n8262) );
  AND U8078 ( .A(n8268), .B(n8269), .Z(n8267) );
  XNOR U8079 ( .A(p_input[3112]), .B(n8266), .Z(n8269) );
  XNOR U8080 ( .A(n8266), .B(n7978), .Z(n8268) );
  IV U8081 ( .A(p_input[3080]), .Z(n7978) );
  XOR U8082 ( .A(n8270), .B(n8271), .Z(n8266) );
  AND U8083 ( .A(n8272), .B(n8273), .Z(n8271) );
  XNOR U8084 ( .A(p_input[3111]), .B(n8270), .Z(n8273) );
  XNOR U8085 ( .A(n8270), .B(n7987), .Z(n8272) );
  IV U8086 ( .A(p_input[3079]), .Z(n7987) );
  XOR U8087 ( .A(n8274), .B(n8275), .Z(n8270) );
  AND U8088 ( .A(n8276), .B(n8277), .Z(n8275) );
  XNOR U8089 ( .A(p_input[3110]), .B(n8274), .Z(n8277) );
  XNOR U8090 ( .A(n8274), .B(n7996), .Z(n8276) );
  IV U8091 ( .A(p_input[3078]), .Z(n7996) );
  XOR U8092 ( .A(n8278), .B(n8279), .Z(n8274) );
  AND U8093 ( .A(n8280), .B(n8281), .Z(n8279) );
  XNOR U8094 ( .A(p_input[3109]), .B(n8278), .Z(n8281) );
  XNOR U8095 ( .A(n8278), .B(n8005), .Z(n8280) );
  IV U8096 ( .A(p_input[3077]), .Z(n8005) );
  XOR U8097 ( .A(n8282), .B(n8283), .Z(n8278) );
  AND U8098 ( .A(n8284), .B(n8285), .Z(n8283) );
  XNOR U8099 ( .A(p_input[3108]), .B(n8282), .Z(n8285) );
  XNOR U8100 ( .A(n8282), .B(n8014), .Z(n8284) );
  IV U8101 ( .A(p_input[3076]), .Z(n8014) );
  XOR U8102 ( .A(n8286), .B(n8287), .Z(n8282) );
  AND U8103 ( .A(n8288), .B(n8289), .Z(n8287) );
  XNOR U8104 ( .A(p_input[3107]), .B(n8286), .Z(n8289) );
  XNOR U8105 ( .A(n8286), .B(n8023), .Z(n8288) );
  IV U8106 ( .A(p_input[3075]), .Z(n8023) );
  XOR U8107 ( .A(n8290), .B(n8291), .Z(n8286) );
  AND U8108 ( .A(n8292), .B(n8293), .Z(n8291) );
  XNOR U8109 ( .A(p_input[3106]), .B(n8290), .Z(n8293) );
  XNOR U8110 ( .A(n8290), .B(n8032), .Z(n8292) );
  IV U8111 ( .A(p_input[3074]), .Z(n8032) );
  XNOR U8112 ( .A(n8294), .B(n8295), .Z(n8290) );
  AND U8113 ( .A(n8296), .B(n8297), .Z(n8295) );
  XOR U8114 ( .A(p_input[3105]), .B(n8294), .Z(n8297) );
  XNOR U8115 ( .A(p_input[3073]), .B(n8294), .Z(n8296) );
  AND U8116 ( .A(p_input[3104]), .B(n8298), .Z(n8294) );
  IV U8117 ( .A(p_input[3072]), .Z(n8298) );
  XOR U8118 ( .A(n8299), .B(n8300), .Z(n1011) );
  AND U8119 ( .A(n616), .B(n8301), .Z(n8300) );
  XNOR U8120 ( .A(n8302), .B(n8299), .Z(n8301) );
  XOR U8121 ( .A(n8303), .B(n8304), .Z(n616) );
  AND U8122 ( .A(n8305), .B(n8306), .Z(n8304) );
  XOR U8123 ( .A(n8303), .B(n1026), .Z(n8306) );
  XOR U8124 ( .A(n8307), .B(n8308), .Z(n1026) );
  AND U8125 ( .A(n582), .B(n8309), .Z(n8308) );
  XOR U8126 ( .A(n8310), .B(n8307), .Z(n8309) );
  XNOR U8127 ( .A(n1023), .B(n8303), .Z(n8305) );
  XOR U8128 ( .A(n8311), .B(n8312), .Z(n1023) );
  AND U8129 ( .A(n579), .B(n8313), .Z(n8312) );
  XOR U8130 ( .A(n8314), .B(n8311), .Z(n8313) );
  XOR U8131 ( .A(n8315), .B(n8316), .Z(n8303) );
  AND U8132 ( .A(n8317), .B(n8318), .Z(n8316) );
  XOR U8133 ( .A(n8315), .B(n1038), .Z(n8318) );
  XOR U8134 ( .A(n8319), .B(n8320), .Z(n1038) );
  AND U8135 ( .A(n582), .B(n8321), .Z(n8320) );
  XOR U8136 ( .A(n8322), .B(n8319), .Z(n8321) );
  XNOR U8137 ( .A(n1035), .B(n8315), .Z(n8317) );
  XOR U8138 ( .A(n8323), .B(n8324), .Z(n1035) );
  AND U8139 ( .A(n579), .B(n8325), .Z(n8324) );
  XOR U8140 ( .A(n8326), .B(n8323), .Z(n8325) );
  XOR U8141 ( .A(n8327), .B(n8328), .Z(n8315) );
  AND U8142 ( .A(n8329), .B(n8330), .Z(n8328) );
  XOR U8143 ( .A(n8327), .B(n1050), .Z(n8330) );
  XOR U8144 ( .A(n8331), .B(n8332), .Z(n1050) );
  AND U8145 ( .A(n582), .B(n8333), .Z(n8332) );
  XOR U8146 ( .A(n8334), .B(n8331), .Z(n8333) );
  XNOR U8147 ( .A(n1047), .B(n8327), .Z(n8329) );
  XOR U8148 ( .A(n8335), .B(n8336), .Z(n1047) );
  AND U8149 ( .A(n579), .B(n8337), .Z(n8336) );
  XOR U8150 ( .A(n8338), .B(n8335), .Z(n8337) );
  XOR U8151 ( .A(n8339), .B(n8340), .Z(n8327) );
  AND U8152 ( .A(n8341), .B(n8342), .Z(n8340) );
  XOR U8153 ( .A(n8339), .B(n1062), .Z(n8342) );
  XOR U8154 ( .A(n8343), .B(n8344), .Z(n1062) );
  AND U8155 ( .A(n582), .B(n8345), .Z(n8344) );
  XOR U8156 ( .A(n8346), .B(n8343), .Z(n8345) );
  XNOR U8157 ( .A(n1059), .B(n8339), .Z(n8341) );
  XOR U8158 ( .A(n8347), .B(n8348), .Z(n1059) );
  AND U8159 ( .A(n579), .B(n8349), .Z(n8348) );
  XOR U8160 ( .A(n8350), .B(n8347), .Z(n8349) );
  XOR U8161 ( .A(n8351), .B(n8352), .Z(n8339) );
  AND U8162 ( .A(n8353), .B(n8354), .Z(n8352) );
  XOR U8163 ( .A(n8351), .B(n1074), .Z(n8354) );
  XOR U8164 ( .A(n8355), .B(n8356), .Z(n1074) );
  AND U8165 ( .A(n582), .B(n8357), .Z(n8356) );
  XOR U8166 ( .A(n8358), .B(n8355), .Z(n8357) );
  XNOR U8167 ( .A(n1071), .B(n8351), .Z(n8353) );
  XOR U8168 ( .A(n8359), .B(n8360), .Z(n1071) );
  AND U8169 ( .A(n579), .B(n8361), .Z(n8360) );
  XOR U8170 ( .A(n8362), .B(n8359), .Z(n8361) );
  XOR U8171 ( .A(n8363), .B(n8364), .Z(n8351) );
  AND U8172 ( .A(n8365), .B(n8366), .Z(n8364) );
  XOR U8173 ( .A(n8363), .B(n1086), .Z(n8366) );
  XOR U8174 ( .A(n8367), .B(n8368), .Z(n1086) );
  AND U8175 ( .A(n582), .B(n8369), .Z(n8368) );
  XOR U8176 ( .A(n8370), .B(n8367), .Z(n8369) );
  XNOR U8177 ( .A(n1083), .B(n8363), .Z(n8365) );
  XOR U8178 ( .A(n8371), .B(n8372), .Z(n1083) );
  AND U8179 ( .A(n579), .B(n8373), .Z(n8372) );
  XOR U8180 ( .A(n8374), .B(n8371), .Z(n8373) );
  XOR U8181 ( .A(n8375), .B(n8376), .Z(n8363) );
  AND U8182 ( .A(n8377), .B(n8378), .Z(n8376) );
  XOR U8183 ( .A(n8375), .B(n1098), .Z(n8378) );
  XOR U8184 ( .A(n8379), .B(n8380), .Z(n1098) );
  AND U8185 ( .A(n582), .B(n8381), .Z(n8380) );
  XOR U8186 ( .A(n8382), .B(n8379), .Z(n8381) );
  XNOR U8187 ( .A(n1095), .B(n8375), .Z(n8377) );
  XOR U8188 ( .A(n8383), .B(n8384), .Z(n1095) );
  AND U8189 ( .A(n579), .B(n8385), .Z(n8384) );
  XOR U8190 ( .A(n8386), .B(n8383), .Z(n8385) );
  XOR U8191 ( .A(n8387), .B(n8388), .Z(n8375) );
  AND U8192 ( .A(n8389), .B(n8390), .Z(n8388) );
  XOR U8193 ( .A(n8387), .B(n1110), .Z(n8390) );
  XOR U8194 ( .A(n8391), .B(n8392), .Z(n1110) );
  AND U8195 ( .A(n582), .B(n8393), .Z(n8392) );
  XOR U8196 ( .A(n8394), .B(n8391), .Z(n8393) );
  XNOR U8197 ( .A(n1107), .B(n8387), .Z(n8389) );
  XOR U8198 ( .A(n8395), .B(n8396), .Z(n1107) );
  AND U8199 ( .A(n579), .B(n8397), .Z(n8396) );
  XOR U8200 ( .A(n8398), .B(n8395), .Z(n8397) );
  XOR U8201 ( .A(n8399), .B(n8400), .Z(n8387) );
  AND U8202 ( .A(n8401), .B(n8402), .Z(n8400) );
  XOR U8203 ( .A(n8399), .B(n1122), .Z(n8402) );
  XOR U8204 ( .A(n8403), .B(n8404), .Z(n1122) );
  AND U8205 ( .A(n582), .B(n8405), .Z(n8404) );
  XOR U8206 ( .A(n8406), .B(n8403), .Z(n8405) );
  XNOR U8207 ( .A(n1119), .B(n8399), .Z(n8401) );
  XOR U8208 ( .A(n8407), .B(n8408), .Z(n1119) );
  AND U8209 ( .A(n579), .B(n8409), .Z(n8408) );
  XOR U8210 ( .A(n8410), .B(n8407), .Z(n8409) );
  XOR U8211 ( .A(n8411), .B(n8412), .Z(n8399) );
  AND U8212 ( .A(n8413), .B(n8414), .Z(n8412) );
  XOR U8213 ( .A(n8411), .B(n1134), .Z(n8414) );
  XOR U8214 ( .A(n8415), .B(n8416), .Z(n1134) );
  AND U8215 ( .A(n582), .B(n8417), .Z(n8416) );
  XOR U8216 ( .A(n8418), .B(n8415), .Z(n8417) );
  XNOR U8217 ( .A(n1131), .B(n8411), .Z(n8413) );
  XOR U8218 ( .A(n8419), .B(n8420), .Z(n1131) );
  AND U8219 ( .A(n579), .B(n8421), .Z(n8420) );
  XOR U8220 ( .A(n8422), .B(n8419), .Z(n8421) );
  XOR U8221 ( .A(n8423), .B(n8424), .Z(n8411) );
  AND U8222 ( .A(n8425), .B(n8426), .Z(n8424) );
  XOR U8223 ( .A(n8423), .B(n1146), .Z(n8426) );
  XOR U8224 ( .A(n8427), .B(n8428), .Z(n1146) );
  AND U8225 ( .A(n582), .B(n8429), .Z(n8428) );
  XOR U8226 ( .A(n8430), .B(n8427), .Z(n8429) );
  XNOR U8227 ( .A(n1143), .B(n8423), .Z(n8425) );
  XOR U8228 ( .A(n8431), .B(n8432), .Z(n1143) );
  AND U8229 ( .A(n579), .B(n8433), .Z(n8432) );
  XOR U8230 ( .A(n8434), .B(n8431), .Z(n8433) );
  XOR U8231 ( .A(n8435), .B(n8436), .Z(n8423) );
  AND U8232 ( .A(n8437), .B(n8438), .Z(n8436) );
  XOR U8233 ( .A(n8435), .B(n1158), .Z(n8438) );
  XOR U8234 ( .A(n8439), .B(n8440), .Z(n1158) );
  AND U8235 ( .A(n582), .B(n8441), .Z(n8440) );
  XOR U8236 ( .A(n8442), .B(n8439), .Z(n8441) );
  XNOR U8237 ( .A(n1155), .B(n8435), .Z(n8437) );
  XOR U8238 ( .A(n8443), .B(n8444), .Z(n1155) );
  AND U8239 ( .A(n579), .B(n8445), .Z(n8444) );
  XOR U8240 ( .A(n8446), .B(n8443), .Z(n8445) );
  XOR U8241 ( .A(n8447), .B(n8448), .Z(n8435) );
  AND U8242 ( .A(n8449), .B(n8450), .Z(n8448) );
  XOR U8243 ( .A(n8447), .B(n1170), .Z(n8450) );
  XOR U8244 ( .A(n8451), .B(n8452), .Z(n1170) );
  AND U8245 ( .A(n582), .B(n8453), .Z(n8452) );
  XOR U8246 ( .A(n8454), .B(n8451), .Z(n8453) );
  XNOR U8247 ( .A(n1167), .B(n8447), .Z(n8449) );
  XOR U8248 ( .A(n8455), .B(n8456), .Z(n1167) );
  AND U8249 ( .A(n579), .B(n8457), .Z(n8456) );
  XOR U8250 ( .A(n8458), .B(n8455), .Z(n8457) );
  XOR U8251 ( .A(n8459), .B(n8460), .Z(n8447) );
  AND U8252 ( .A(n8461), .B(n8462), .Z(n8460) );
  XOR U8253 ( .A(n8459), .B(n1182), .Z(n8462) );
  XOR U8254 ( .A(n8463), .B(n8464), .Z(n1182) );
  AND U8255 ( .A(n582), .B(n8465), .Z(n8464) );
  XOR U8256 ( .A(n8466), .B(n8463), .Z(n8465) );
  XNOR U8257 ( .A(n1179), .B(n8459), .Z(n8461) );
  XOR U8258 ( .A(n8467), .B(n8468), .Z(n1179) );
  AND U8259 ( .A(n579), .B(n8469), .Z(n8468) );
  XOR U8260 ( .A(n8470), .B(n8467), .Z(n8469) );
  XOR U8261 ( .A(n8471), .B(n8472), .Z(n8459) );
  AND U8262 ( .A(n8473), .B(n8474), .Z(n8472) );
  XOR U8263 ( .A(n8471), .B(n1194), .Z(n8474) );
  XOR U8264 ( .A(n8475), .B(n8476), .Z(n1194) );
  AND U8265 ( .A(n582), .B(n8477), .Z(n8476) );
  XOR U8266 ( .A(n8478), .B(n8475), .Z(n8477) );
  XNOR U8267 ( .A(n1191), .B(n8471), .Z(n8473) );
  XOR U8268 ( .A(n8479), .B(n8480), .Z(n1191) );
  AND U8269 ( .A(n579), .B(n8481), .Z(n8480) );
  XOR U8270 ( .A(n8482), .B(n8479), .Z(n8481) );
  XOR U8271 ( .A(n8483), .B(n8484), .Z(n8471) );
  AND U8272 ( .A(n8485), .B(n8486), .Z(n8484) );
  XOR U8273 ( .A(n8483), .B(n1206), .Z(n8486) );
  XOR U8274 ( .A(n8487), .B(n8488), .Z(n1206) );
  AND U8275 ( .A(n582), .B(n8489), .Z(n8488) );
  XOR U8276 ( .A(n8490), .B(n8487), .Z(n8489) );
  XNOR U8277 ( .A(n1203), .B(n8483), .Z(n8485) );
  XOR U8278 ( .A(n8491), .B(n8492), .Z(n1203) );
  AND U8279 ( .A(n579), .B(n8493), .Z(n8492) );
  XOR U8280 ( .A(n8494), .B(n8491), .Z(n8493) );
  XOR U8281 ( .A(n8495), .B(n8496), .Z(n8483) );
  AND U8282 ( .A(n8497), .B(n8498), .Z(n8496) );
  XOR U8283 ( .A(n8495), .B(n1218), .Z(n8498) );
  XOR U8284 ( .A(n8499), .B(n8500), .Z(n1218) );
  AND U8285 ( .A(n582), .B(n8501), .Z(n8500) );
  XOR U8286 ( .A(n8502), .B(n8499), .Z(n8501) );
  XNOR U8287 ( .A(n1215), .B(n8495), .Z(n8497) );
  XOR U8288 ( .A(n8503), .B(n8504), .Z(n1215) );
  AND U8289 ( .A(n579), .B(n8505), .Z(n8504) );
  XOR U8290 ( .A(n8506), .B(n8503), .Z(n8505) );
  XOR U8291 ( .A(n8507), .B(n8508), .Z(n8495) );
  AND U8292 ( .A(n8509), .B(n8510), .Z(n8508) );
  XOR U8293 ( .A(n8507), .B(n1230), .Z(n8510) );
  XOR U8294 ( .A(n8511), .B(n8512), .Z(n1230) );
  AND U8295 ( .A(n582), .B(n8513), .Z(n8512) );
  XOR U8296 ( .A(n8514), .B(n8511), .Z(n8513) );
  XNOR U8297 ( .A(n1227), .B(n8507), .Z(n8509) );
  XOR U8298 ( .A(n8515), .B(n8516), .Z(n1227) );
  AND U8299 ( .A(n579), .B(n8517), .Z(n8516) );
  XOR U8300 ( .A(n8518), .B(n8515), .Z(n8517) );
  XOR U8301 ( .A(n8519), .B(n8520), .Z(n8507) );
  AND U8302 ( .A(n8521), .B(n8522), .Z(n8520) );
  XOR U8303 ( .A(n8519), .B(n1242), .Z(n8522) );
  XOR U8304 ( .A(n8523), .B(n8524), .Z(n1242) );
  AND U8305 ( .A(n582), .B(n8525), .Z(n8524) );
  XOR U8306 ( .A(n8526), .B(n8523), .Z(n8525) );
  XNOR U8307 ( .A(n1239), .B(n8519), .Z(n8521) );
  XOR U8308 ( .A(n8527), .B(n8528), .Z(n1239) );
  AND U8309 ( .A(n579), .B(n8529), .Z(n8528) );
  XOR U8310 ( .A(n8530), .B(n8527), .Z(n8529) );
  XOR U8311 ( .A(n8531), .B(n8532), .Z(n8519) );
  AND U8312 ( .A(n8533), .B(n8534), .Z(n8532) );
  XOR U8313 ( .A(n8531), .B(n1254), .Z(n8534) );
  XOR U8314 ( .A(n8535), .B(n8536), .Z(n1254) );
  AND U8315 ( .A(n582), .B(n8537), .Z(n8536) );
  XOR U8316 ( .A(n8538), .B(n8535), .Z(n8537) );
  XNOR U8317 ( .A(n1251), .B(n8531), .Z(n8533) );
  XOR U8318 ( .A(n8539), .B(n8540), .Z(n1251) );
  AND U8319 ( .A(n579), .B(n8541), .Z(n8540) );
  XOR U8320 ( .A(n8542), .B(n8539), .Z(n8541) );
  XOR U8321 ( .A(n8543), .B(n8544), .Z(n8531) );
  AND U8322 ( .A(n8545), .B(n8546), .Z(n8544) );
  XOR U8323 ( .A(n8543), .B(n1266), .Z(n8546) );
  XOR U8324 ( .A(n8547), .B(n8548), .Z(n1266) );
  AND U8325 ( .A(n582), .B(n8549), .Z(n8548) );
  XOR U8326 ( .A(n8550), .B(n8547), .Z(n8549) );
  XNOR U8327 ( .A(n1263), .B(n8543), .Z(n8545) );
  XOR U8328 ( .A(n8551), .B(n8552), .Z(n1263) );
  AND U8329 ( .A(n579), .B(n8553), .Z(n8552) );
  XOR U8330 ( .A(n8554), .B(n8551), .Z(n8553) );
  XOR U8331 ( .A(n8555), .B(n8556), .Z(n8543) );
  AND U8332 ( .A(n8557), .B(n8558), .Z(n8556) );
  XOR U8333 ( .A(n8555), .B(n1278), .Z(n8558) );
  XOR U8334 ( .A(n8559), .B(n8560), .Z(n1278) );
  AND U8335 ( .A(n582), .B(n8561), .Z(n8560) );
  XOR U8336 ( .A(n8562), .B(n8559), .Z(n8561) );
  XNOR U8337 ( .A(n1275), .B(n8555), .Z(n8557) );
  XOR U8338 ( .A(n8563), .B(n8564), .Z(n1275) );
  AND U8339 ( .A(n579), .B(n8565), .Z(n8564) );
  XOR U8340 ( .A(n8566), .B(n8563), .Z(n8565) );
  XOR U8341 ( .A(n8567), .B(n8568), .Z(n8555) );
  AND U8342 ( .A(n8569), .B(n8570), .Z(n8568) );
  XOR U8343 ( .A(n8567), .B(n1290), .Z(n8570) );
  XOR U8344 ( .A(n8571), .B(n8572), .Z(n1290) );
  AND U8345 ( .A(n582), .B(n8573), .Z(n8572) );
  XOR U8346 ( .A(n8574), .B(n8571), .Z(n8573) );
  XNOR U8347 ( .A(n1287), .B(n8567), .Z(n8569) );
  XOR U8348 ( .A(n8575), .B(n8576), .Z(n1287) );
  AND U8349 ( .A(n579), .B(n8577), .Z(n8576) );
  XOR U8350 ( .A(n8578), .B(n8575), .Z(n8577) );
  XOR U8351 ( .A(n8579), .B(n8580), .Z(n8567) );
  AND U8352 ( .A(n8581), .B(n8582), .Z(n8580) );
  XOR U8353 ( .A(n8579), .B(n1302), .Z(n8582) );
  XOR U8354 ( .A(n8583), .B(n8584), .Z(n1302) );
  AND U8355 ( .A(n582), .B(n8585), .Z(n8584) );
  XOR U8356 ( .A(n8586), .B(n8583), .Z(n8585) );
  XNOR U8357 ( .A(n1299), .B(n8579), .Z(n8581) );
  XOR U8358 ( .A(n8587), .B(n8588), .Z(n1299) );
  AND U8359 ( .A(n579), .B(n8589), .Z(n8588) );
  XOR U8360 ( .A(n8590), .B(n8587), .Z(n8589) );
  XOR U8361 ( .A(n8591), .B(n8592), .Z(n8579) );
  AND U8362 ( .A(n8593), .B(n8594), .Z(n8592) );
  XOR U8363 ( .A(n8591), .B(n1314), .Z(n8594) );
  XOR U8364 ( .A(n8595), .B(n8596), .Z(n1314) );
  AND U8365 ( .A(n582), .B(n8597), .Z(n8596) );
  XOR U8366 ( .A(n8598), .B(n8595), .Z(n8597) );
  XNOR U8367 ( .A(n1311), .B(n8591), .Z(n8593) );
  XOR U8368 ( .A(n8599), .B(n8600), .Z(n1311) );
  AND U8369 ( .A(n579), .B(n8601), .Z(n8600) );
  XOR U8370 ( .A(n8602), .B(n8599), .Z(n8601) );
  XOR U8371 ( .A(n8603), .B(n8604), .Z(n8591) );
  AND U8372 ( .A(n8605), .B(n8606), .Z(n8604) );
  XOR U8373 ( .A(n8603), .B(n1326), .Z(n8606) );
  XOR U8374 ( .A(n8607), .B(n8608), .Z(n1326) );
  AND U8375 ( .A(n582), .B(n8609), .Z(n8608) );
  XOR U8376 ( .A(n8610), .B(n8607), .Z(n8609) );
  XNOR U8377 ( .A(n1323), .B(n8603), .Z(n8605) );
  XOR U8378 ( .A(n8611), .B(n8612), .Z(n1323) );
  AND U8379 ( .A(n579), .B(n8613), .Z(n8612) );
  XOR U8380 ( .A(n8614), .B(n8611), .Z(n8613) );
  XOR U8381 ( .A(n8615), .B(n8616), .Z(n8603) );
  AND U8382 ( .A(n8617), .B(n8618), .Z(n8616) );
  XOR U8383 ( .A(n8615), .B(n1338), .Z(n8618) );
  XOR U8384 ( .A(n8619), .B(n8620), .Z(n1338) );
  AND U8385 ( .A(n582), .B(n8621), .Z(n8620) );
  XOR U8386 ( .A(n8622), .B(n8619), .Z(n8621) );
  XNOR U8387 ( .A(n1335), .B(n8615), .Z(n8617) );
  XOR U8388 ( .A(n8623), .B(n8624), .Z(n1335) );
  AND U8389 ( .A(n579), .B(n8625), .Z(n8624) );
  XOR U8390 ( .A(n8626), .B(n8623), .Z(n8625) );
  XOR U8391 ( .A(n8627), .B(n8628), .Z(n8615) );
  AND U8392 ( .A(n8629), .B(n8630), .Z(n8628) );
  XOR U8393 ( .A(n8627), .B(n1350), .Z(n8630) );
  XOR U8394 ( .A(n8631), .B(n8632), .Z(n1350) );
  AND U8395 ( .A(n582), .B(n8633), .Z(n8632) );
  XOR U8396 ( .A(n8634), .B(n8631), .Z(n8633) );
  XNOR U8397 ( .A(n1347), .B(n8627), .Z(n8629) );
  XOR U8398 ( .A(n8635), .B(n8636), .Z(n1347) );
  AND U8399 ( .A(n579), .B(n8637), .Z(n8636) );
  XOR U8400 ( .A(n8638), .B(n8635), .Z(n8637) );
  XOR U8401 ( .A(n8639), .B(n8640), .Z(n8627) );
  AND U8402 ( .A(n8641), .B(n8642), .Z(n8640) );
  XOR U8403 ( .A(n8639), .B(n1362), .Z(n8642) );
  XOR U8404 ( .A(n8643), .B(n8644), .Z(n1362) );
  AND U8405 ( .A(n582), .B(n8645), .Z(n8644) );
  XOR U8406 ( .A(n8646), .B(n8643), .Z(n8645) );
  XNOR U8407 ( .A(n1359), .B(n8639), .Z(n8641) );
  XOR U8408 ( .A(n8647), .B(n8648), .Z(n1359) );
  AND U8409 ( .A(n579), .B(n8649), .Z(n8648) );
  XOR U8410 ( .A(n8650), .B(n8647), .Z(n8649) );
  XOR U8411 ( .A(n8651), .B(n8652), .Z(n8639) );
  AND U8412 ( .A(n8653), .B(n8654), .Z(n8652) );
  XOR U8413 ( .A(n1374), .B(n8651), .Z(n8654) );
  XOR U8414 ( .A(n8655), .B(n8656), .Z(n1374) );
  AND U8415 ( .A(n582), .B(n8657), .Z(n8656) );
  XOR U8416 ( .A(n8655), .B(n8658), .Z(n8657) );
  XNOR U8417 ( .A(n8651), .B(n1371), .Z(n8653) );
  XOR U8418 ( .A(n8659), .B(n8660), .Z(n1371) );
  AND U8419 ( .A(n579), .B(n8661), .Z(n8660) );
  XOR U8420 ( .A(n8659), .B(n8662), .Z(n8661) );
  XOR U8421 ( .A(n8663), .B(n8664), .Z(n8651) );
  AND U8422 ( .A(n8665), .B(n8666), .Z(n8664) );
  XNOR U8423 ( .A(n8667), .B(n1387), .Z(n8666) );
  XOR U8424 ( .A(n8668), .B(n8669), .Z(n1387) );
  AND U8425 ( .A(n582), .B(n8670), .Z(n8669) );
  XOR U8426 ( .A(n8671), .B(n8668), .Z(n8670) );
  XNOR U8427 ( .A(n1384), .B(n8663), .Z(n8665) );
  XOR U8428 ( .A(n8672), .B(n8673), .Z(n1384) );
  AND U8429 ( .A(n579), .B(n8674), .Z(n8673) );
  XOR U8430 ( .A(n8675), .B(n8672), .Z(n8674) );
  IV U8431 ( .A(n8667), .Z(n8663) );
  AND U8432 ( .A(n8299), .B(n8302), .Z(n8667) );
  XNOR U8433 ( .A(n8676), .B(n8677), .Z(n8302) );
  AND U8434 ( .A(n582), .B(n8678), .Z(n8677) );
  XNOR U8435 ( .A(n8679), .B(n8676), .Z(n8678) );
  XOR U8436 ( .A(n8680), .B(n8681), .Z(n582) );
  AND U8437 ( .A(n8682), .B(n8683), .Z(n8681) );
  XOR U8438 ( .A(n8680), .B(n8310), .Z(n8683) );
  XOR U8439 ( .A(n8684), .B(n8685), .Z(n8310) );
  AND U8440 ( .A(n502), .B(n8686), .Z(n8685) );
  XOR U8441 ( .A(n8687), .B(n8684), .Z(n8686) );
  XNOR U8442 ( .A(n8307), .B(n8680), .Z(n8682) );
  XOR U8443 ( .A(n8688), .B(n8689), .Z(n8307) );
  AND U8444 ( .A(n500), .B(n8690), .Z(n8689) );
  XOR U8445 ( .A(n8691), .B(n8688), .Z(n8690) );
  XOR U8446 ( .A(n8692), .B(n8693), .Z(n8680) );
  AND U8447 ( .A(n8694), .B(n8695), .Z(n8693) );
  XOR U8448 ( .A(n8692), .B(n8322), .Z(n8695) );
  XOR U8449 ( .A(n8696), .B(n8697), .Z(n8322) );
  AND U8450 ( .A(n502), .B(n8698), .Z(n8697) );
  XOR U8451 ( .A(n8699), .B(n8696), .Z(n8698) );
  XNOR U8452 ( .A(n8319), .B(n8692), .Z(n8694) );
  XOR U8453 ( .A(n8700), .B(n8701), .Z(n8319) );
  AND U8454 ( .A(n500), .B(n8702), .Z(n8701) );
  XOR U8455 ( .A(n8703), .B(n8700), .Z(n8702) );
  XOR U8456 ( .A(n8704), .B(n8705), .Z(n8692) );
  AND U8457 ( .A(n8706), .B(n8707), .Z(n8705) );
  XOR U8458 ( .A(n8704), .B(n8334), .Z(n8707) );
  XOR U8459 ( .A(n8708), .B(n8709), .Z(n8334) );
  AND U8460 ( .A(n502), .B(n8710), .Z(n8709) );
  XOR U8461 ( .A(n8711), .B(n8708), .Z(n8710) );
  XNOR U8462 ( .A(n8331), .B(n8704), .Z(n8706) );
  XOR U8463 ( .A(n8712), .B(n8713), .Z(n8331) );
  AND U8464 ( .A(n500), .B(n8714), .Z(n8713) );
  XOR U8465 ( .A(n8715), .B(n8712), .Z(n8714) );
  XOR U8466 ( .A(n8716), .B(n8717), .Z(n8704) );
  AND U8467 ( .A(n8718), .B(n8719), .Z(n8717) );
  XOR U8468 ( .A(n8716), .B(n8346), .Z(n8719) );
  XOR U8469 ( .A(n8720), .B(n8721), .Z(n8346) );
  AND U8470 ( .A(n502), .B(n8722), .Z(n8721) );
  XOR U8471 ( .A(n8723), .B(n8720), .Z(n8722) );
  XNOR U8472 ( .A(n8343), .B(n8716), .Z(n8718) );
  XOR U8473 ( .A(n8724), .B(n8725), .Z(n8343) );
  AND U8474 ( .A(n500), .B(n8726), .Z(n8725) );
  XOR U8475 ( .A(n8727), .B(n8724), .Z(n8726) );
  XOR U8476 ( .A(n8728), .B(n8729), .Z(n8716) );
  AND U8477 ( .A(n8730), .B(n8731), .Z(n8729) );
  XOR U8478 ( .A(n8728), .B(n8358), .Z(n8731) );
  XOR U8479 ( .A(n8732), .B(n8733), .Z(n8358) );
  AND U8480 ( .A(n502), .B(n8734), .Z(n8733) );
  XOR U8481 ( .A(n8735), .B(n8732), .Z(n8734) );
  XNOR U8482 ( .A(n8355), .B(n8728), .Z(n8730) );
  XOR U8483 ( .A(n8736), .B(n8737), .Z(n8355) );
  AND U8484 ( .A(n500), .B(n8738), .Z(n8737) );
  XOR U8485 ( .A(n8739), .B(n8736), .Z(n8738) );
  XOR U8486 ( .A(n8740), .B(n8741), .Z(n8728) );
  AND U8487 ( .A(n8742), .B(n8743), .Z(n8741) );
  XOR U8488 ( .A(n8740), .B(n8370), .Z(n8743) );
  XOR U8489 ( .A(n8744), .B(n8745), .Z(n8370) );
  AND U8490 ( .A(n502), .B(n8746), .Z(n8745) );
  XOR U8491 ( .A(n8747), .B(n8744), .Z(n8746) );
  XNOR U8492 ( .A(n8367), .B(n8740), .Z(n8742) );
  XOR U8493 ( .A(n8748), .B(n8749), .Z(n8367) );
  AND U8494 ( .A(n500), .B(n8750), .Z(n8749) );
  XOR U8495 ( .A(n8751), .B(n8748), .Z(n8750) );
  XOR U8496 ( .A(n8752), .B(n8753), .Z(n8740) );
  AND U8497 ( .A(n8754), .B(n8755), .Z(n8753) );
  XOR U8498 ( .A(n8752), .B(n8382), .Z(n8755) );
  XOR U8499 ( .A(n8756), .B(n8757), .Z(n8382) );
  AND U8500 ( .A(n502), .B(n8758), .Z(n8757) );
  XOR U8501 ( .A(n8759), .B(n8756), .Z(n8758) );
  XNOR U8502 ( .A(n8379), .B(n8752), .Z(n8754) );
  XOR U8503 ( .A(n8760), .B(n8761), .Z(n8379) );
  AND U8504 ( .A(n500), .B(n8762), .Z(n8761) );
  XOR U8505 ( .A(n8763), .B(n8760), .Z(n8762) );
  XOR U8506 ( .A(n8764), .B(n8765), .Z(n8752) );
  AND U8507 ( .A(n8766), .B(n8767), .Z(n8765) );
  XOR U8508 ( .A(n8764), .B(n8394), .Z(n8767) );
  XOR U8509 ( .A(n8768), .B(n8769), .Z(n8394) );
  AND U8510 ( .A(n502), .B(n8770), .Z(n8769) );
  XOR U8511 ( .A(n8771), .B(n8768), .Z(n8770) );
  XNOR U8512 ( .A(n8391), .B(n8764), .Z(n8766) );
  XOR U8513 ( .A(n8772), .B(n8773), .Z(n8391) );
  AND U8514 ( .A(n500), .B(n8774), .Z(n8773) );
  XOR U8515 ( .A(n8775), .B(n8772), .Z(n8774) );
  XOR U8516 ( .A(n8776), .B(n8777), .Z(n8764) );
  AND U8517 ( .A(n8778), .B(n8779), .Z(n8777) );
  XOR U8518 ( .A(n8776), .B(n8406), .Z(n8779) );
  XOR U8519 ( .A(n8780), .B(n8781), .Z(n8406) );
  AND U8520 ( .A(n502), .B(n8782), .Z(n8781) );
  XOR U8521 ( .A(n8783), .B(n8780), .Z(n8782) );
  XNOR U8522 ( .A(n8403), .B(n8776), .Z(n8778) );
  XOR U8523 ( .A(n8784), .B(n8785), .Z(n8403) );
  AND U8524 ( .A(n500), .B(n8786), .Z(n8785) );
  XOR U8525 ( .A(n8787), .B(n8784), .Z(n8786) );
  XOR U8526 ( .A(n8788), .B(n8789), .Z(n8776) );
  AND U8527 ( .A(n8790), .B(n8791), .Z(n8789) );
  XOR U8528 ( .A(n8788), .B(n8418), .Z(n8791) );
  XOR U8529 ( .A(n8792), .B(n8793), .Z(n8418) );
  AND U8530 ( .A(n502), .B(n8794), .Z(n8793) );
  XOR U8531 ( .A(n8795), .B(n8792), .Z(n8794) );
  XNOR U8532 ( .A(n8415), .B(n8788), .Z(n8790) );
  XOR U8533 ( .A(n8796), .B(n8797), .Z(n8415) );
  AND U8534 ( .A(n500), .B(n8798), .Z(n8797) );
  XOR U8535 ( .A(n8799), .B(n8796), .Z(n8798) );
  XOR U8536 ( .A(n8800), .B(n8801), .Z(n8788) );
  AND U8537 ( .A(n8802), .B(n8803), .Z(n8801) );
  XOR U8538 ( .A(n8800), .B(n8430), .Z(n8803) );
  XOR U8539 ( .A(n8804), .B(n8805), .Z(n8430) );
  AND U8540 ( .A(n502), .B(n8806), .Z(n8805) );
  XOR U8541 ( .A(n8807), .B(n8804), .Z(n8806) );
  XNOR U8542 ( .A(n8427), .B(n8800), .Z(n8802) );
  XOR U8543 ( .A(n8808), .B(n8809), .Z(n8427) );
  AND U8544 ( .A(n500), .B(n8810), .Z(n8809) );
  XOR U8545 ( .A(n8811), .B(n8808), .Z(n8810) );
  XOR U8546 ( .A(n8812), .B(n8813), .Z(n8800) );
  AND U8547 ( .A(n8814), .B(n8815), .Z(n8813) );
  XOR U8548 ( .A(n8812), .B(n8442), .Z(n8815) );
  XOR U8549 ( .A(n8816), .B(n8817), .Z(n8442) );
  AND U8550 ( .A(n502), .B(n8818), .Z(n8817) );
  XOR U8551 ( .A(n8819), .B(n8816), .Z(n8818) );
  XNOR U8552 ( .A(n8439), .B(n8812), .Z(n8814) );
  XOR U8553 ( .A(n8820), .B(n8821), .Z(n8439) );
  AND U8554 ( .A(n500), .B(n8822), .Z(n8821) );
  XOR U8555 ( .A(n8823), .B(n8820), .Z(n8822) );
  XOR U8556 ( .A(n8824), .B(n8825), .Z(n8812) );
  AND U8557 ( .A(n8826), .B(n8827), .Z(n8825) );
  XOR U8558 ( .A(n8824), .B(n8454), .Z(n8827) );
  XOR U8559 ( .A(n8828), .B(n8829), .Z(n8454) );
  AND U8560 ( .A(n502), .B(n8830), .Z(n8829) );
  XOR U8561 ( .A(n8831), .B(n8828), .Z(n8830) );
  XNOR U8562 ( .A(n8451), .B(n8824), .Z(n8826) );
  XOR U8563 ( .A(n8832), .B(n8833), .Z(n8451) );
  AND U8564 ( .A(n500), .B(n8834), .Z(n8833) );
  XOR U8565 ( .A(n8835), .B(n8832), .Z(n8834) );
  XOR U8566 ( .A(n8836), .B(n8837), .Z(n8824) );
  AND U8567 ( .A(n8838), .B(n8839), .Z(n8837) );
  XOR U8568 ( .A(n8836), .B(n8466), .Z(n8839) );
  XOR U8569 ( .A(n8840), .B(n8841), .Z(n8466) );
  AND U8570 ( .A(n502), .B(n8842), .Z(n8841) );
  XOR U8571 ( .A(n8843), .B(n8840), .Z(n8842) );
  XNOR U8572 ( .A(n8463), .B(n8836), .Z(n8838) );
  XOR U8573 ( .A(n8844), .B(n8845), .Z(n8463) );
  AND U8574 ( .A(n500), .B(n8846), .Z(n8845) );
  XOR U8575 ( .A(n8847), .B(n8844), .Z(n8846) );
  XOR U8576 ( .A(n8848), .B(n8849), .Z(n8836) );
  AND U8577 ( .A(n8850), .B(n8851), .Z(n8849) );
  XOR U8578 ( .A(n8848), .B(n8478), .Z(n8851) );
  XOR U8579 ( .A(n8852), .B(n8853), .Z(n8478) );
  AND U8580 ( .A(n502), .B(n8854), .Z(n8853) );
  XOR U8581 ( .A(n8855), .B(n8852), .Z(n8854) );
  XNOR U8582 ( .A(n8475), .B(n8848), .Z(n8850) );
  XOR U8583 ( .A(n8856), .B(n8857), .Z(n8475) );
  AND U8584 ( .A(n500), .B(n8858), .Z(n8857) );
  XOR U8585 ( .A(n8859), .B(n8856), .Z(n8858) );
  XOR U8586 ( .A(n8860), .B(n8861), .Z(n8848) );
  AND U8587 ( .A(n8862), .B(n8863), .Z(n8861) );
  XOR U8588 ( .A(n8860), .B(n8490), .Z(n8863) );
  XOR U8589 ( .A(n8864), .B(n8865), .Z(n8490) );
  AND U8590 ( .A(n502), .B(n8866), .Z(n8865) );
  XOR U8591 ( .A(n8867), .B(n8864), .Z(n8866) );
  XNOR U8592 ( .A(n8487), .B(n8860), .Z(n8862) );
  XOR U8593 ( .A(n8868), .B(n8869), .Z(n8487) );
  AND U8594 ( .A(n500), .B(n8870), .Z(n8869) );
  XOR U8595 ( .A(n8871), .B(n8868), .Z(n8870) );
  XOR U8596 ( .A(n8872), .B(n8873), .Z(n8860) );
  AND U8597 ( .A(n8874), .B(n8875), .Z(n8873) );
  XOR U8598 ( .A(n8872), .B(n8502), .Z(n8875) );
  XOR U8599 ( .A(n8876), .B(n8877), .Z(n8502) );
  AND U8600 ( .A(n502), .B(n8878), .Z(n8877) );
  XOR U8601 ( .A(n8879), .B(n8876), .Z(n8878) );
  XNOR U8602 ( .A(n8499), .B(n8872), .Z(n8874) );
  XOR U8603 ( .A(n8880), .B(n8881), .Z(n8499) );
  AND U8604 ( .A(n500), .B(n8882), .Z(n8881) );
  XOR U8605 ( .A(n8883), .B(n8880), .Z(n8882) );
  XOR U8606 ( .A(n8884), .B(n8885), .Z(n8872) );
  AND U8607 ( .A(n8886), .B(n8887), .Z(n8885) );
  XOR U8608 ( .A(n8884), .B(n8514), .Z(n8887) );
  XOR U8609 ( .A(n8888), .B(n8889), .Z(n8514) );
  AND U8610 ( .A(n502), .B(n8890), .Z(n8889) );
  XOR U8611 ( .A(n8891), .B(n8888), .Z(n8890) );
  XNOR U8612 ( .A(n8511), .B(n8884), .Z(n8886) );
  XOR U8613 ( .A(n8892), .B(n8893), .Z(n8511) );
  AND U8614 ( .A(n500), .B(n8894), .Z(n8893) );
  XOR U8615 ( .A(n8895), .B(n8892), .Z(n8894) );
  XOR U8616 ( .A(n8896), .B(n8897), .Z(n8884) );
  AND U8617 ( .A(n8898), .B(n8899), .Z(n8897) );
  XOR U8618 ( .A(n8896), .B(n8526), .Z(n8899) );
  XOR U8619 ( .A(n8900), .B(n8901), .Z(n8526) );
  AND U8620 ( .A(n502), .B(n8902), .Z(n8901) );
  XOR U8621 ( .A(n8903), .B(n8900), .Z(n8902) );
  XNOR U8622 ( .A(n8523), .B(n8896), .Z(n8898) );
  XOR U8623 ( .A(n8904), .B(n8905), .Z(n8523) );
  AND U8624 ( .A(n500), .B(n8906), .Z(n8905) );
  XOR U8625 ( .A(n8907), .B(n8904), .Z(n8906) );
  XOR U8626 ( .A(n8908), .B(n8909), .Z(n8896) );
  AND U8627 ( .A(n8910), .B(n8911), .Z(n8909) );
  XOR U8628 ( .A(n8908), .B(n8538), .Z(n8911) );
  XOR U8629 ( .A(n8912), .B(n8913), .Z(n8538) );
  AND U8630 ( .A(n502), .B(n8914), .Z(n8913) );
  XOR U8631 ( .A(n8915), .B(n8912), .Z(n8914) );
  XNOR U8632 ( .A(n8535), .B(n8908), .Z(n8910) );
  XOR U8633 ( .A(n8916), .B(n8917), .Z(n8535) );
  AND U8634 ( .A(n500), .B(n8918), .Z(n8917) );
  XOR U8635 ( .A(n8919), .B(n8916), .Z(n8918) );
  XOR U8636 ( .A(n8920), .B(n8921), .Z(n8908) );
  AND U8637 ( .A(n8922), .B(n8923), .Z(n8921) );
  XOR U8638 ( .A(n8920), .B(n8550), .Z(n8923) );
  XOR U8639 ( .A(n8924), .B(n8925), .Z(n8550) );
  AND U8640 ( .A(n502), .B(n8926), .Z(n8925) );
  XOR U8641 ( .A(n8927), .B(n8924), .Z(n8926) );
  XNOR U8642 ( .A(n8547), .B(n8920), .Z(n8922) );
  XOR U8643 ( .A(n8928), .B(n8929), .Z(n8547) );
  AND U8644 ( .A(n500), .B(n8930), .Z(n8929) );
  XOR U8645 ( .A(n8931), .B(n8928), .Z(n8930) );
  XOR U8646 ( .A(n8932), .B(n8933), .Z(n8920) );
  AND U8647 ( .A(n8934), .B(n8935), .Z(n8933) );
  XOR U8648 ( .A(n8932), .B(n8562), .Z(n8935) );
  XOR U8649 ( .A(n8936), .B(n8937), .Z(n8562) );
  AND U8650 ( .A(n502), .B(n8938), .Z(n8937) );
  XOR U8651 ( .A(n8939), .B(n8936), .Z(n8938) );
  XNOR U8652 ( .A(n8559), .B(n8932), .Z(n8934) );
  XOR U8653 ( .A(n8940), .B(n8941), .Z(n8559) );
  AND U8654 ( .A(n500), .B(n8942), .Z(n8941) );
  XOR U8655 ( .A(n8943), .B(n8940), .Z(n8942) );
  XOR U8656 ( .A(n8944), .B(n8945), .Z(n8932) );
  AND U8657 ( .A(n8946), .B(n8947), .Z(n8945) );
  XOR U8658 ( .A(n8944), .B(n8574), .Z(n8947) );
  XOR U8659 ( .A(n8948), .B(n8949), .Z(n8574) );
  AND U8660 ( .A(n502), .B(n8950), .Z(n8949) );
  XOR U8661 ( .A(n8951), .B(n8948), .Z(n8950) );
  XNOR U8662 ( .A(n8571), .B(n8944), .Z(n8946) );
  XOR U8663 ( .A(n8952), .B(n8953), .Z(n8571) );
  AND U8664 ( .A(n500), .B(n8954), .Z(n8953) );
  XOR U8665 ( .A(n8955), .B(n8952), .Z(n8954) );
  XOR U8666 ( .A(n8956), .B(n8957), .Z(n8944) );
  AND U8667 ( .A(n8958), .B(n8959), .Z(n8957) );
  XOR U8668 ( .A(n8956), .B(n8586), .Z(n8959) );
  XOR U8669 ( .A(n8960), .B(n8961), .Z(n8586) );
  AND U8670 ( .A(n502), .B(n8962), .Z(n8961) );
  XOR U8671 ( .A(n8963), .B(n8960), .Z(n8962) );
  XNOR U8672 ( .A(n8583), .B(n8956), .Z(n8958) );
  XOR U8673 ( .A(n8964), .B(n8965), .Z(n8583) );
  AND U8674 ( .A(n500), .B(n8966), .Z(n8965) );
  XOR U8675 ( .A(n8967), .B(n8964), .Z(n8966) );
  XOR U8676 ( .A(n8968), .B(n8969), .Z(n8956) );
  AND U8677 ( .A(n8970), .B(n8971), .Z(n8969) );
  XOR U8678 ( .A(n8968), .B(n8598), .Z(n8971) );
  XOR U8679 ( .A(n8972), .B(n8973), .Z(n8598) );
  AND U8680 ( .A(n502), .B(n8974), .Z(n8973) );
  XOR U8681 ( .A(n8975), .B(n8972), .Z(n8974) );
  XNOR U8682 ( .A(n8595), .B(n8968), .Z(n8970) );
  XOR U8683 ( .A(n8976), .B(n8977), .Z(n8595) );
  AND U8684 ( .A(n500), .B(n8978), .Z(n8977) );
  XOR U8685 ( .A(n8979), .B(n8976), .Z(n8978) );
  XOR U8686 ( .A(n8980), .B(n8981), .Z(n8968) );
  AND U8687 ( .A(n8982), .B(n8983), .Z(n8981) );
  XOR U8688 ( .A(n8980), .B(n8610), .Z(n8983) );
  XOR U8689 ( .A(n8984), .B(n8985), .Z(n8610) );
  AND U8690 ( .A(n502), .B(n8986), .Z(n8985) );
  XOR U8691 ( .A(n8987), .B(n8984), .Z(n8986) );
  XNOR U8692 ( .A(n8607), .B(n8980), .Z(n8982) );
  XOR U8693 ( .A(n8988), .B(n8989), .Z(n8607) );
  AND U8694 ( .A(n500), .B(n8990), .Z(n8989) );
  XOR U8695 ( .A(n8991), .B(n8988), .Z(n8990) );
  XOR U8696 ( .A(n8992), .B(n8993), .Z(n8980) );
  AND U8697 ( .A(n8994), .B(n8995), .Z(n8993) );
  XOR U8698 ( .A(n8992), .B(n8622), .Z(n8995) );
  XOR U8699 ( .A(n8996), .B(n8997), .Z(n8622) );
  AND U8700 ( .A(n502), .B(n8998), .Z(n8997) );
  XOR U8701 ( .A(n8999), .B(n8996), .Z(n8998) );
  XNOR U8702 ( .A(n8619), .B(n8992), .Z(n8994) );
  XOR U8703 ( .A(n9000), .B(n9001), .Z(n8619) );
  AND U8704 ( .A(n500), .B(n9002), .Z(n9001) );
  XOR U8705 ( .A(n9003), .B(n9000), .Z(n9002) );
  XOR U8706 ( .A(n9004), .B(n9005), .Z(n8992) );
  AND U8707 ( .A(n9006), .B(n9007), .Z(n9005) );
  XOR U8708 ( .A(n9004), .B(n8634), .Z(n9007) );
  XOR U8709 ( .A(n9008), .B(n9009), .Z(n8634) );
  AND U8710 ( .A(n502), .B(n9010), .Z(n9009) );
  XOR U8711 ( .A(n9011), .B(n9008), .Z(n9010) );
  XNOR U8712 ( .A(n8631), .B(n9004), .Z(n9006) );
  XOR U8713 ( .A(n9012), .B(n9013), .Z(n8631) );
  AND U8714 ( .A(n500), .B(n9014), .Z(n9013) );
  XOR U8715 ( .A(n9015), .B(n9012), .Z(n9014) );
  XOR U8716 ( .A(n9016), .B(n9017), .Z(n9004) );
  AND U8717 ( .A(n9018), .B(n9019), .Z(n9017) );
  XOR U8718 ( .A(n9016), .B(n8646), .Z(n9019) );
  XOR U8719 ( .A(n9020), .B(n9021), .Z(n8646) );
  AND U8720 ( .A(n502), .B(n9022), .Z(n9021) );
  XOR U8721 ( .A(n9023), .B(n9020), .Z(n9022) );
  XNOR U8722 ( .A(n8643), .B(n9016), .Z(n9018) );
  XOR U8723 ( .A(n9024), .B(n9025), .Z(n8643) );
  AND U8724 ( .A(n500), .B(n9026), .Z(n9025) );
  XOR U8725 ( .A(n9027), .B(n9024), .Z(n9026) );
  XOR U8726 ( .A(n9028), .B(n9029), .Z(n9016) );
  AND U8727 ( .A(n9030), .B(n9031), .Z(n9029) );
  XOR U8728 ( .A(n8658), .B(n9028), .Z(n9031) );
  XOR U8729 ( .A(n9032), .B(n9033), .Z(n8658) );
  AND U8730 ( .A(n502), .B(n9034), .Z(n9033) );
  XOR U8731 ( .A(n9032), .B(n9035), .Z(n9034) );
  XNOR U8732 ( .A(n9028), .B(n8655), .Z(n9030) );
  XOR U8733 ( .A(n9036), .B(n9037), .Z(n8655) );
  AND U8734 ( .A(n500), .B(n9038), .Z(n9037) );
  XOR U8735 ( .A(n9036), .B(n9039), .Z(n9038) );
  XOR U8736 ( .A(n9040), .B(n9041), .Z(n9028) );
  AND U8737 ( .A(n9042), .B(n9043), .Z(n9041) );
  XNOR U8738 ( .A(n9044), .B(n8671), .Z(n9043) );
  XOR U8739 ( .A(n9045), .B(n9046), .Z(n8671) );
  AND U8740 ( .A(n502), .B(n9047), .Z(n9046) );
  XOR U8741 ( .A(n9048), .B(n9045), .Z(n9047) );
  XNOR U8742 ( .A(n8668), .B(n9040), .Z(n9042) );
  XOR U8743 ( .A(n9049), .B(n9050), .Z(n8668) );
  AND U8744 ( .A(n500), .B(n9051), .Z(n9050) );
  XOR U8745 ( .A(n9052), .B(n9049), .Z(n9051) );
  IV U8746 ( .A(n9044), .Z(n9040) );
  AND U8747 ( .A(n8676), .B(n8679), .Z(n9044) );
  XNOR U8748 ( .A(n9053), .B(n9054), .Z(n8679) );
  AND U8749 ( .A(n502), .B(n9055), .Z(n9054) );
  XNOR U8750 ( .A(n9056), .B(n9053), .Z(n9055) );
  XOR U8751 ( .A(n9057), .B(n9058), .Z(n502) );
  AND U8752 ( .A(n9059), .B(n9060), .Z(n9058) );
  XOR U8753 ( .A(n9057), .B(n8687), .Z(n9060) );
  XNOR U8754 ( .A(n9061), .B(n9062), .Z(n8687) );
  AND U8755 ( .A(n9063), .B(n334), .Z(n9062) );
  AND U8756 ( .A(n9061), .B(n9064), .Z(n9063) );
  XNOR U8757 ( .A(n8684), .B(n9057), .Z(n9059) );
  XOR U8758 ( .A(n9065), .B(n9066), .Z(n8684) );
  AND U8759 ( .A(n9067), .B(n332), .Z(n9066) );
  NOR U8760 ( .A(n9065), .B(n9068), .Z(n9067) );
  XOR U8761 ( .A(n9069), .B(n9070), .Z(n9057) );
  AND U8762 ( .A(n9071), .B(n9072), .Z(n9070) );
  XOR U8763 ( .A(n9069), .B(n8699), .Z(n9072) );
  XOR U8764 ( .A(n9073), .B(n9074), .Z(n8699) );
  AND U8765 ( .A(n334), .B(n9075), .Z(n9074) );
  XOR U8766 ( .A(n9076), .B(n9073), .Z(n9075) );
  XNOR U8767 ( .A(n8696), .B(n9069), .Z(n9071) );
  XOR U8768 ( .A(n9077), .B(n9078), .Z(n8696) );
  AND U8769 ( .A(n332), .B(n9079), .Z(n9078) );
  XOR U8770 ( .A(n9080), .B(n9077), .Z(n9079) );
  XOR U8771 ( .A(n9081), .B(n9082), .Z(n9069) );
  AND U8772 ( .A(n9083), .B(n9084), .Z(n9082) );
  XOR U8773 ( .A(n9081), .B(n8711), .Z(n9084) );
  XOR U8774 ( .A(n9085), .B(n9086), .Z(n8711) );
  AND U8775 ( .A(n334), .B(n9087), .Z(n9086) );
  XOR U8776 ( .A(n9088), .B(n9085), .Z(n9087) );
  XNOR U8777 ( .A(n8708), .B(n9081), .Z(n9083) );
  XOR U8778 ( .A(n9089), .B(n9090), .Z(n8708) );
  AND U8779 ( .A(n332), .B(n9091), .Z(n9090) );
  XOR U8780 ( .A(n9092), .B(n9089), .Z(n9091) );
  XOR U8781 ( .A(n9093), .B(n9094), .Z(n9081) );
  AND U8782 ( .A(n9095), .B(n9096), .Z(n9094) );
  XOR U8783 ( .A(n9093), .B(n8723), .Z(n9096) );
  XOR U8784 ( .A(n9097), .B(n9098), .Z(n8723) );
  AND U8785 ( .A(n334), .B(n9099), .Z(n9098) );
  XOR U8786 ( .A(n9100), .B(n9097), .Z(n9099) );
  XNOR U8787 ( .A(n8720), .B(n9093), .Z(n9095) );
  XOR U8788 ( .A(n9101), .B(n9102), .Z(n8720) );
  AND U8789 ( .A(n332), .B(n9103), .Z(n9102) );
  XOR U8790 ( .A(n9104), .B(n9101), .Z(n9103) );
  XOR U8791 ( .A(n9105), .B(n9106), .Z(n9093) );
  AND U8792 ( .A(n9107), .B(n9108), .Z(n9106) );
  XOR U8793 ( .A(n9105), .B(n8735), .Z(n9108) );
  XOR U8794 ( .A(n9109), .B(n9110), .Z(n8735) );
  AND U8795 ( .A(n334), .B(n9111), .Z(n9110) );
  XOR U8796 ( .A(n9112), .B(n9109), .Z(n9111) );
  XNOR U8797 ( .A(n8732), .B(n9105), .Z(n9107) );
  XOR U8798 ( .A(n9113), .B(n9114), .Z(n8732) );
  AND U8799 ( .A(n332), .B(n9115), .Z(n9114) );
  XOR U8800 ( .A(n9116), .B(n9113), .Z(n9115) );
  XOR U8801 ( .A(n9117), .B(n9118), .Z(n9105) );
  AND U8802 ( .A(n9119), .B(n9120), .Z(n9118) );
  XOR U8803 ( .A(n9117), .B(n8747), .Z(n9120) );
  XOR U8804 ( .A(n9121), .B(n9122), .Z(n8747) );
  AND U8805 ( .A(n334), .B(n9123), .Z(n9122) );
  XOR U8806 ( .A(n9124), .B(n9121), .Z(n9123) );
  XNOR U8807 ( .A(n8744), .B(n9117), .Z(n9119) );
  XOR U8808 ( .A(n9125), .B(n9126), .Z(n8744) );
  AND U8809 ( .A(n332), .B(n9127), .Z(n9126) );
  XOR U8810 ( .A(n9128), .B(n9125), .Z(n9127) );
  XOR U8811 ( .A(n9129), .B(n9130), .Z(n9117) );
  AND U8812 ( .A(n9131), .B(n9132), .Z(n9130) );
  XOR U8813 ( .A(n9129), .B(n8759), .Z(n9132) );
  XOR U8814 ( .A(n9133), .B(n9134), .Z(n8759) );
  AND U8815 ( .A(n334), .B(n9135), .Z(n9134) );
  XOR U8816 ( .A(n9136), .B(n9133), .Z(n9135) );
  XNOR U8817 ( .A(n8756), .B(n9129), .Z(n9131) );
  XOR U8818 ( .A(n9137), .B(n9138), .Z(n8756) );
  AND U8819 ( .A(n332), .B(n9139), .Z(n9138) );
  XOR U8820 ( .A(n9140), .B(n9137), .Z(n9139) );
  XOR U8821 ( .A(n9141), .B(n9142), .Z(n9129) );
  AND U8822 ( .A(n9143), .B(n9144), .Z(n9142) );
  XOR U8823 ( .A(n9141), .B(n8771), .Z(n9144) );
  XOR U8824 ( .A(n9145), .B(n9146), .Z(n8771) );
  AND U8825 ( .A(n334), .B(n9147), .Z(n9146) );
  XOR U8826 ( .A(n9148), .B(n9145), .Z(n9147) );
  XNOR U8827 ( .A(n8768), .B(n9141), .Z(n9143) );
  XOR U8828 ( .A(n9149), .B(n9150), .Z(n8768) );
  AND U8829 ( .A(n332), .B(n9151), .Z(n9150) );
  XOR U8830 ( .A(n9152), .B(n9149), .Z(n9151) );
  XOR U8831 ( .A(n9153), .B(n9154), .Z(n9141) );
  AND U8832 ( .A(n9155), .B(n9156), .Z(n9154) );
  XOR U8833 ( .A(n9153), .B(n8783), .Z(n9156) );
  XOR U8834 ( .A(n9157), .B(n9158), .Z(n8783) );
  AND U8835 ( .A(n334), .B(n9159), .Z(n9158) );
  XOR U8836 ( .A(n9160), .B(n9157), .Z(n9159) );
  XNOR U8837 ( .A(n8780), .B(n9153), .Z(n9155) );
  XOR U8838 ( .A(n9161), .B(n9162), .Z(n8780) );
  AND U8839 ( .A(n332), .B(n9163), .Z(n9162) );
  XOR U8840 ( .A(n9164), .B(n9161), .Z(n9163) );
  XOR U8841 ( .A(n9165), .B(n9166), .Z(n9153) );
  AND U8842 ( .A(n9167), .B(n9168), .Z(n9166) );
  XOR U8843 ( .A(n9165), .B(n8795), .Z(n9168) );
  XOR U8844 ( .A(n9169), .B(n9170), .Z(n8795) );
  AND U8845 ( .A(n334), .B(n9171), .Z(n9170) );
  XOR U8846 ( .A(n9172), .B(n9169), .Z(n9171) );
  XNOR U8847 ( .A(n8792), .B(n9165), .Z(n9167) );
  XOR U8848 ( .A(n9173), .B(n9174), .Z(n8792) );
  AND U8849 ( .A(n332), .B(n9175), .Z(n9174) );
  XOR U8850 ( .A(n9176), .B(n9173), .Z(n9175) );
  XOR U8851 ( .A(n9177), .B(n9178), .Z(n9165) );
  AND U8852 ( .A(n9179), .B(n9180), .Z(n9178) );
  XOR U8853 ( .A(n9177), .B(n8807), .Z(n9180) );
  XOR U8854 ( .A(n9181), .B(n9182), .Z(n8807) );
  AND U8855 ( .A(n334), .B(n9183), .Z(n9182) );
  XOR U8856 ( .A(n9184), .B(n9181), .Z(n9183) );
  XNOR U8857 ( .A(n8804), .B(n9177), .Z(n9179) );
  XOR U8858 ( .A(n9185), .B(n9186), .Z(n8804) );
  AND U8859 ( .A(n332), .B(n9187), .Z(n9186) );
  XOR U8860 ( .A(n9188), .B(n9185), .Z(n9187) );
  XOR U8861 ( .A(n9189), .B(n9190), .Z(n9177) );
  AND U8862 ( .A(n9191), .B(n9192), .Z(n9190) );
  XOR U8863 ( .A(n9189), .B(n8819), .Z(n9192) );
  XOR U8864 ( .A(n9193), .B(n9194), .Z(n8819) );
  AND U8865 ( .A(n334), .B(n9195), .Z(n9194) );
  XOR U8866 ( .A(n9196), .B(n9193), .Z(n9195) );
  XNOR U8867 ( .A(n8816), .B(n9189), .Z(n9191) );
  XOR U8868 ( .A(n9197), .B(n9198), .Z(n8816) );
  AND U8869 ( .A(n332), .B(n9199), .Z(n9198) );
  XOR U8870 ( .A(n9200), .B(n9197), .Z(n9199) );
  XOR U8871 ( .A(n9201), .B(n9202), .Z(n9189) );
  AND U8872 ( .A(n9203), .B(n9204), .Z(n9202) );
  XOR U8873 ( .A(n9201), .B(n8831), .Z(n9204) );
  XOR U8874 ( .A(n9205), .B(n9206), .Z(n8831) );
  AND U8875 ( .A(n334), .B(n9207), .Z(n9206) );
  XOR U8876 ( .A(n9208), .B(n9205), .Z(n9207) );
  XNOR U8877 ( .A(n8828), .B(n9201), .Z(n9203) );
  XOR U8878 ( .A(n9209), .B(n9210), .Z(n8828) );
  AND U8879 ( .A(n332), .B(n9211), .Z(n9210) );
  XOR U8880 ( .A(n9212), .B(n9209), .Z(n9211) );
  XOR U8881 ( .A(n9213), .B(n9214), .Z(n9201) );
  AND U8882 ( .A(n9215), .B(n9216), .Z(n9214) );
  XOR U8883 ( .A(n9213), .B(n8843), .Z(n9216) );
  XOR U8884 ( .A(n9217), .B(n9218), .Z(n8843) );
  AND U8885 ( .A(n334), .B(n9219), .Z(n9218) );
  XOR U8886 ( .A(n9220), .B(n9217), .Z(n9219) );
  XNOR U8887 ( .A(n8840), .B(n9213), .Z(n9215) );
  XOR U8888 ( .A(n9221), .B(n9222), .Z(n8840) );
  AND U8889 ( .A(n332), .B(n9223), .Z(n9222) );
  XOR U8890 ( .A(n9224), .B(n9221), .Z(n9223) );
  XOR U8891 ( .A(n9225), .B(n9226), .Z(n9213) );
  AND U8892 ( .A(n9227), .B(n9228), .Z(n9226) );
  XOR U8893 ( .A(n9225), .B(n8855), .Z(n9228) );
  XOR U8894 ( .A(n9229), .B(n9230), .Z(n8855) );
  AND U8895 ( .A(n334), .B(n9231), .Z(n9230) );
  XOR U8896 ( .A(n9232), .B(n9229), .Z(n9231) );
  XNOR U8897 ( .A(n8852), .B(n9225), .Z(n9227) );
  XOR U8898 ( .A(n9233), .B(n9234), .Z(n8852) );
  AND U8899 ( .A(n332), .B(n9235), .Z(n9234) );
  XOR U8900 ( .A(n9236), .B(n9233), .Z(n9235) );
  XOR U8901 ( .A(n9237), .B(n9238), .Z(n9225) );
  AND U8902 ( .A(n9239), .B(n9240), .Z(n9238) );
  XOR U8903 ( .A(n9237), .B(n8867), .Z(n9240) );
  XOR U8904 ( .A(n9241), .B(n9242), .Z(n8867) );
  AND U8905 ( .A(n334), .B(n9243), .Z(n9242) );
  XOR U8906 ( .A(n9244), .B(n9241), .Z(n9243) );
  XNOR U8907 ( .A(n8864), .B(n9237), .Z(n9239) );
  XOR U8908 ( .A(n9245), .B(n9246), .Z(n8864) );
  AND U8909 ( .A(n332), .B(n9247), .Z(n9246) );
  XOR U8910 ( .A(n9248), .B(n9245), .Z(n9247) );
  XOR U8911 ( .A(n9249), .B(n9250), .Z(n9237) );
  AND U8912 ( .A(n9251), .B(n9252), .Z(n9250) );
  XOR U8913 ( .A(n9249), .B(n8879), .Z(n9252) );
  XOR U8914 ( .A(n9253), .B(n9254), .Z(n8879) );
  AND U8915 ( .A(n334), .B(n9255), .Z(n9254) );
  XOR U8916 ( .A(n9256), .B(n9253), .Z(n9255) );
  XNOR U8917 ( .A(n8876), .B(n9249), .Z(n9251) );
  XOR U8918 ( .A(n9257), .B(n9258), .Z(n8876) );
  AND U8919 ( .A(n332), .B(n9259), .Z(n9258) );
  XOR U8920 ( .A(n9260), .B(n9257), .Z(n9259) );
  XOR U8921 ( .A(n9261), .B(n9262), .Z(n9249) );
  AND U8922 ( .A(n9263), .B(n9264), .Z(n9262) );
  XOR U8923 ( .A(n9261), .B(n8891), .Z(n9264) );
  XOR U8924 ( .A(n9265), .B(n9266), .Z(n8891) );
  AND U8925 ( .A(n334), .B(n9267), .Z(n9266) );
  XOR U8926 ( .A(n9268), .B(n9265), .Z(n9267) );
  XNOR U8927 ( .A(n8888), .B(n9261), .Z(n9263) );
  XOR U8928 ( .A(n9269), .B(n9270), .Z(n8888) );
  AND U8929 ( .A(n332), .B(n9271), .Z(n9270) );
  XOR U8930 ( .A(n9272), .B(n9269), .Z(n9271) );
  XOR U8931 ( .A(n9273), .B(n9274), .Z(n9261) );
  AND U8932 ( .A(n9275), .B(n9276), .Z(n9274) );
  XOR U8933 ( .A(n9273), .B(n8903), .Z(n9276) );
  XOR U8934 ( .A(n9277), .B(n9278), .Z(n8903) );
  AND U8935 ( .A(n334), .B(n9279), .Z(n9278) );
  XOR U8936 ( .A(n9280), .B(n9277), .Z(n9279) );
  XNOR U8937 ( .A(n8900), .B(n9273), .Z(n9275) );
  XOR U8938 ( .A(n9281), .B(n9282), .Z(n8900) );
  AND U8939 ( .A(n332), .B(n9283), .Z(n9282) );
  XOR U8940 ( .A(n9284), .B(n9281), .Z(n9283) );
  XOR U8941 ( .A(n9285), .B(n9286), .Z(n9273) );
  AND U8942 ( .A(n9287), .B(n9288), .Z(n9286) );
  XOR U8943 ( .A(n9285), .B(n8915), .Z(n9288) );
  XOR U8944 ( .A(n9289), .B(n9290), .Z(n8915) );
  AND U8945 ( .A(n334), .B(n9291), .Z(n9290) );
  XOR U8946 ( .A(n9292), .B(n9289), .Z(n9291) );
  XNOR U8947 ( .A(n8912), .B(n9285), .Z(n9287) );
  XOR U8948 ( .A(n9293), .B(n9294), .Z(n8912) );
  AND U8949 ( .A(n332), .B(n9295), .Z(n9294) );
  XOR U8950 ( .A(n9296), .B(n9293), .Z(n9295) );
  XOR U8951 ( .A(n9297), .B(n9298), .Z(n9285) );
  AND U8952 ( .A(n9299), .B(n9300), .Z(n9298) );
  XOR U8953 ( .A(n9297), .B(n8927), .Z(n9300) );
  XOR U8954 ( .A(n9301), .B(n9302), .Z(n8927) );
  AND U8955 ( .A(n334), .B(n9303), .Z(n9302) );
  XOR U8956 ( .A(n9304), .B(n9301), .Z(n9303) );
  XNOR U8957 ( .A(n8924), .B(n9297), .Z(n9299) );
  XOR U8958 ( .A(n9305), .B(n9306), .Z(n8924) );
  AND U8959 ( .A(n332), .B(n9307), .Z(n9306) );
  XOR U8960 ( .A(n9308), .B(n9305), .Z(n9307) );
  XOR U8961 ( .A(n9309), .B(n9310), .Z(n9297) );
  AND U8962 ( .A(n9311), .B(n9312), .Z(n9310) );
  XOR U8963 ( .A(n9309), .B(n8939), .Z(n9312) );
  XOR U8964 ( .A(n9313), .B(n9314), .Z(n8939) );
  AND U8965 ( .A(n334), .B(n9315), .Z(n9314) );
  XOR U8966 ( .A(n9316), .B(n9313), .Z(n9315) );
  XNOR U8967 ( .A(n8936), .B(n9309), .Z(n9311) );
  XOR U8968 ( .A(n9317), .B(n9318), .Z(n8936) );
  AND U8969 ( .A(n332), .B(n9319), .Z(n9318) );
  XOR U8970 ( .A(n9320), .B(n9317), .Z(n9319) );
  XOR U8971 ( .A(n9321), .B(n9322), .Z(n9309) );
  AND U8972 ( .A(n9323), .B(n9324), .Z(n9322) );
  XOR U8973 ( .A(n9321), .B(n8951), .Z(n9324) );
  XOR U8974 ( .A(n9325), .B(n9326), .Z(n8951) );
  AND U8975 ( .A(n334), .B(n9327), .Z(n9326) );
  XOR U8976 ( .A(n9328), .B(n9325), .Z(n9327) );
  XNOR U8977 ( .A(n8948), .B(n9321), .Z(n9323) );
  XOR U8978 ( .A(n9329), .B(n9330), .Z(n8948) );
  AND U8979 ( .A(n332), .B(n9331), .Z(n9330) );
  XOR U8980 ( .A(n9332), .B(n9329), .Z(n9331) );
  XOR U8981 ( .A(n9333), .B(n9334), .Z(n9321) );
  AND U8982 ( .A(n9335), .B(n9336), .Z(n9334) );
  XOR U8983 ( .A(n9333), .B(n8963), .Z(n9336) );
  XOR U8984 ( .A(n9337), .B(n9338), .Z(n8963) );
  AND U8985 ( .A(n334), .B(n9339), .Z(n9338) );
  XOR U8986 ( .A(n9340), .B(n9337), .Z(n9339) );
  XNOR U8987 ( .A(n8960), .B(n9333), .Z(n9335) );
  XOR U8988 ( .A(n9341), .B(n9342), .Z(n8960) );
  AND U8989 ( .A(n332), .B(n9343), .Z(n9342) );
  XOR U8990 ( .A(n9344), .B(n9341), .Z(n9343) );
  XOR U8991 ( .A(n9345), .B(n9346), .Z(n9333) );
  AND U8992 ( .A(n9347), .B(n9348), .Z(n9346) );
  XOR U8993 ( .A(n9345), .B(n8975), .Z(n9348) );
  XOR U8994 ( .A(n9349), .B(n9350), .Z(n8975) );
  AND U8995 ( .A(n334), .B(n9351), .Z(n9350) );
  XOR U8996 ( .A(n9352), .B(n9349), .Z(n9351) );
  XNOR U8997 ( .A(n8972), .B(n9345), .Z(n9347) );
  XOR U8998 ( .A(n9353), .B(n9354), .Z(n8972) );
  AND U8999 ( .A(n332), .B(n9355), .Z(n9354) );
  XOR U9000 ( .A(n9356), .B(n9353), .Z(n9355) );
  XOR U9001 ( .A(n9357), .B(n9358), .Z(n9345) );
  AND U9002 ( .A(n9359), .B(n9360), .Z(n9358) );
  XOR U9003 ( .A(n9357), .B(n8987), .Z(n9360) );
  XOR U9004 ( .A(n9361), .B(n9362), .Z(n8987) );
  AND U9005 ( .A(n334), .B(n9363), .Z(n9362) );
  XOR U9006 ( .A(n9364), .B(n9361), .Z(n9363) );
  XNOR U9007 ( .A(n8984), .B(n9357), .Z(n9359) );
  XOR U9008 ( .A(n9365), .B(n9366), .Z(n8984) );
  AND U9009 ( .A(n332), .B(n9367), .Z(n9366) );
  XOR U9010 ( .A(n9368), .B(n9365), .Z(n9367) );
  XOR U9011 ( .A(n9369), .B(n9370), .Z(n9357) );
  AND U9012 ( .A(n9371), .B(n9372), .Z(n9370) );
  XOR U9013 ( .A(n9369), .B(n8999), .Z(n9372) );
  XOR U9014 ( .A(n9373), .B(n9374), .Z(n8999) );
  AND U9015 ( .A(n334), .B(n9375), .Z(n9374) );
  XOR U9016 ( .A(n9376), .B(n9373), .Z(n9375) );
  XNOR U9017 ( .A(n8996), .B(n9369), .Z(n9371) );
  XOR U9018 ( .A(n9377), .B(n9378), .Z(n8996) );
  AND U9019 ( .A(n332), .B(n9379), .Z(n9378) );
  XOR U9020 ( .A(n9380), .B(n9377), .Z(n9379) );
  XOR U9021 ( .A(n9381), .B(n9382), .Z(n9369) );
  AND U9022 ( .A(n9383), .B(n9384), .Z(n9382) );
  XOR U9023 ( .A(n9381), .B(n9011), .Z(n9384) );
  XOR U9024 ( .A(n9385), .B(n9386), .Z(n9011) );
  AND U9025 ( .A(n334), .B(n9387), .Z(n9386) );
  XOR U9026 ( .A(n9388), .B(n9385), .Z(n9387) );
  XNOR U9027 ( .A(n9008), .B(n9381), .Z(n9383) );
  XOR U9028 ( .A(n9389), .B(n9390), .Z(n9008) );
  AND U9029 ( .A(n332), .B(n9391), .Z(n9390) );
  XOR U9030 ( .A(n9392), .B(n9389), .Z(n9391) );
  XOR U9031 ( .A(n9393), .B(n9394), .Z(n9381) );
  AND U9032 ( .A(n9395), .B(n9396), .Z(n9394) );
  XOR U9033 ( .A(n9393), .B(n9023), .Z(n9396) );
  XOR U9034 ( .A(n9397), .B(n9398), .Z(n9023) );
  AND U9035 ( .A(n334), .B(n9399), .Z(n9398) );
  XOR U9036 ( .A(n9400), .B(n9397), .Z(n9399) );
  XNOR U9037 ( .A(n9020), .B(n9393), .Z(n9395) );
  XOR U9038 ( .A(n9401), .B(n9402), .Z(n9020) );
  AND U9039 ( .A(n332), .B(n9403), .Z(n9402) );
  XOR U9040 ( .A(n9404), .B(n9401), .Z(n9403) );
  XOR U9041 ( .A(n9405), .B(n9406), .Z(n9393) );
  AND U9042 ( .A(n9407), .B(n9408), .Z(n9406) );
  XOR U9043 ( .A(n9035), .B(n9405), .Z(n9408) );
  XOR U9044 ( .A(n9409), .B(n9410), .Z(n9035) );
  AND U9045 ( .A(n334), .B(n9411), .Z(n9410) );
  XOR U9046 ( .A(n9409), .B(n9412), .Z(n9411) );
  XNOR U9047 ( .A(n9405), .B(n9032), .Z(n9407) );
  XOR U9048 ( .A(n9413), .B(n9414), .Z(n9032) );
  AND U9049 ( .A(n332), .B(n9415), .Z(n9414) );
  XOR U9050 ( .A(n9413), .B(n9416), .Z(n9415) );
  XOR U9051 ( .A(n9417), .B(n9418), .Z(n9405) );
  AND U9052 ( .A(n9419), .B(n9420), .Z(n9418) );
  XNOR U9053 ( .A(n9421), .B(n9048), .Z(n9420) );
  XOR U9054 ( .A(n9422), .B(n9423), .Z(n9048) );
  AND U9055 ( .A(n334), .B(n9424), .Z(n9423) );
  XOR U9056 ( .A(n9425), .B(n9422), .Z(n9424) );
  XNOR U9057 ( .A(n9045), .B(n9417), .Z(n9419) );
  XOR U9058 ( .A(n9426), .B(n9427), .Z(n9045) );
  AND U9059 ( .A(n332), .B(n9428), .Z(n9427) );
  XOR U9060 ( .A(n9429), .B(n9426), .Z(n9428) );
  IV U9061 ( .A(n9421), .Z(n9417) );
  AND U9062 ( .A(n9053), .B(n9056), .Z(n9421) );
  XNOR U9063 ( .A(n9430), .B(n9431), .Z(n9056) );
  AND U9064 ( .A(n334), .B(n9432), .Z(n9431) );
  XNOR U9065 ( .A(n9433), .B(n9430), .Z(n9432) );
  XOR U9066 ( .A(n9434), .B(n9435), .Z(n334) );
  AND U9067 ( .A(n9436), .B(n9437), .Z(n9435) );
  XOR U9068 ( .A(n9064), .B(n9434), .Z(n9437) );
  IV U9069 ( .A(n9438), .Z(n9064) );
  AND U9070 ( .A(p_input[3071]), .B(p_input[3039]), .Z(n9438) );
  XOR U9071 ( .A(n9434), .B(n9061), .Z(n9436) );
  AND U9072 ( .A(p_input[2975]), .B(p_input[3007]), .Z(n9061) );
  XOR U9073 ( .A(n9439), .B(n9440), .Z(n9434) );
  AND U9074 ( .A(n9441), .B(n9442), .Z(n9440) );
  XOR U9075 ( .A(n9439), .B(n9076), .Z(n9442) );
  XNOR U9076 ( .A(p_input[3038]), .B(n9443), .Z(n9076) );
  AND U9077 ( .A(n242), .B(n9444), .Z(n9443) );
  XOR U9078 ( .A(p_input[3070]), .B(p_input[3038]), .Z(n9444) );
  XNOR U9079 ( .A(n9073), .B(n9439), .Z(n9441) );
  XOR U9080 ( .A(n9445), .B(n9446), .Z(n9073) );
  AND U9081 ( .A(n240), .B(n9447), .Z(n9446) );
  XOR U9082 ( .A(p_input[3006]), .B(p_input[2974]), .Z(n9447) );
  XOR U9083 ( .A(n9448), .B(n9449), .Z(n9439) );
  AND U9084 ( .A(n9450), .B(n9451), .Z(n9449) );
  XOR U9085 ( .A(n9448), .B(n9088), .Z(n9451) );
  XNOR U9086 ( .A(p_input[3037]), .B(n9452), .Z(n9088) );
  AND U9087 ( .A(n242), .B(n9453), .Z(n9452) );
  XOR U9088 ( .A(p_input[3069]), .B(p_input[3037]), .Z(n9453) );
  XNOR U9089 ( .A(n9085), .B(n9448), .Z(n9450) );
  XOR U9090 ( .A(n9454), .B(n9455), .Z(n9085) );
  AND U9091 ( .A(n240), .B(n9456), .Z(n9455) );
  XOR U9092 ( .A(p_input[3005]), .B(p_input[2973]), .Z(n9456) );
  XOR U9093 ( .A(n9457), .B(n9458), .Z(n9448) );
  AND U9094 ( .A(n9459), .B(n9460), .Z(n9458) );
  XOR U9095 ( .A(n9457), .B(n9100), .Z(n9460) );
  XNOR U9096 ( .A(p_input[3036]), .B(n9461), .Z(n9100) );
  AND U9097 ( .A(n242), .B(n9462), .Z(n9461) );
  XOR U9098 ( .A(p_input[3068]), .B(p_input[3036]), .Z(n9462) );
  XNOR U9099 ( .A(n9097), .B(n9457), .Z(n9459) );
  XOR U9100 ( .A(n9463), .B(n9464), .Z(n9097) );
  AND U9101 ( .A(n240), .B(n9465), .Z(n9464) );
  XOR U9102 ( .A(p_input[3004]), .B(p_input[2972]), .Z(n9465) );
  XOR U9103 ( .A(n9466), .B(n9467), .Z(n9457) );
  AND U9104 ( .A(n9468), .B(n9469), .Z(n9467) );
  XOR U9105 ( .A(n9466), .B(n9112), .Z(n9469) );
  XNOR U9106 ( .A(p_input[3035]), .B(n9470), .Z(n9112) );
  AND U9107 ( .A(n242), .B(n9471), .Z(n9470) );
  XOR U9108 ( .A(p_input[3067]), .B(p_input[3035]), .Z(n9471) );
  XNOR U9109 ( .A(n9109), .B(n9466), .Z(n9468) );
  XOR U9110 ( .A(n9472), .B(n9473), .Z(n9109) );
  AND U9111 ( .A(n240), .B(n9474), .Z(n9473) );
  XOR U9112 ( .A(p_input[3003]), .B(p_input[2971]), .Z(n9474) );
  XOR U9113 ( .A(n9475), .B(n9476), .Z(n9466) );
  AND U9114 ( .A(n9477), .B(n9478), .Z(n9476) );
  XOR U9115 ( .A(n9475), .B(n9124), .Z(n9478) );
  XNOR U9116 ( .A(p_input[3034]), .B(n9479), .Z(n9124) );
  AND U9117 ( .A(n242), .B(n9480), .Z(n9479) );
  XOR U9118 ( .A(p_input[3066]), .B(p_input[3034]), .Z(n9480) );
  XNOR U9119 ( .A(n9121), .B(n9475), .Z(n9477) );
  XOR U9120 ( .A(n9481), .B(n9482), .Z(n9121) );
  AND U9121 ( .A(n240), .B(n9483), .Z(n9482) );
  XOR U9122 ( .A(p_input[3002]), .B(p_input[2970]), .Z(n9483) );
  XOR U9123 ( .A(n9484), .B(n9485), .Z(n9475) );
  AND U9124 ( .A(n9486), .B(n9487), .Z(n9485) );
  XOR U9125 ( .A(n9484), .B(n9136), .Z(n9487) );
  XNOR U9126 ( .A(p_input[3033]), .B(n9488), .Z(n9136) );
  AND U9127 ( .A(n242), .B(n9489), .Z(n9488) );
  XOR U9128 ( .A(p_input[3065]), .B(p_input[3033]), .Z(n9489) );
  XNOR U9129 ( .A(n9133), .B(n9484), .Z(n9486) );
  XOR U9130 ( .A(n9490), .B(n9491), .Z(n9133) );
  AND U9131 ( .A(n240), .B(n9492), .Z(n9491) );
  XOR U9132 ( .A(p_input[3001]), .B(p_input[2969]), .Z(n9492) );
  XOR U9133 ( .A(n9493), .B(n9494), .Z(n9484) );
  AND U9134 ( .A(n9495), .B(n9496), .Z(n9494) );
  XOR U9135 ( .A(n9493), .B(n9148), .Z(n9496) );
  XNOR U9136 ( .A(p_input[3032]), .B(n9497), .Z(n9148) );
  AND U9137 ( .A(n242), .B(n9498), .Z(n9497) );
  XOR U9138 ( .A(p_input[3064]), .B(p_input[3032]), .Z(n9498) );
  XNOR U9139 ( .A(n9145), .B(n9493), .Z(n9495) );
  XOR U9140 ( .A(n9499), .B(n9500), .Z(n9145) );
  AND U9141 ( .A(n240), .B(n9501), .Z(n9500) );
  XOR U9142 ( .A(p_input[3000]), .B(p_input[2968]), .Z(n9501) );
  XOR U9143 ( .A(n9502), .B(n9503), .Z(n9493) );
  AND U9144 ( .A(n9504), .B(n9505), .Z(n9503) );
  XOR U9145 ( .A(n9502), .B(n9160), .Z(n9505) );
  XNOR U9146 ( .A(p_input[3031]), .B(n9506), .Z(n9160) );
  AND U9147 ( .A(n242), .B(n9507), .Z(n9506) );
  XOR U9148 ( .A(p_input[3063]), .B(p_input[3031]), .Z(n9507) );
  XNOR U9149 ( .A(n9157), .B(n9502), .Z(n9504) );
  XOR U9150 ( .A(n9508), .B(n9509), .Z(n9157) );
  AND U9151 ( .A(n240), .B(n9510), .Z(n9509) );
  XOR U9152 ( .A(p_input[2999]), .B(p_input[2967]), .Z(n9510) );
  XOR U9153 ( .A(n9511), .B(n9512), .Z(n9502) );
  AND U9154 ( .A(n9513), .B(n9514), .Z(n9512) );
  XOR U9155 ( .A(n9511), .B(n9172), .Z(n9514) );
  XNOR U9156 ( .A(p_input[3030]), .B(n9515), .Z(n9172) );
  AND U9157 ( .A(n242), .B(n9516), .Z(n9515) );
  XOR U9158 ( .A(p_input[3062]), .B(p_input[3030]), .Z(n9516) );
  XNOR U9159 ( .A(n9169), .B(n9511), .Z(n9513) );
  XOR U9160 ( .A(n9517), .B(n9518), .Z(n9169) );
  AND U9161 ( .A(n240), .B(n9519), .Z(n9518) );
  XOR U9162 ( .A(p_input[2998]), .B(p_input[2966]), .Z(n9519) );
  XOR U9163 ( .A(n9520), .B(n9521), .Z(n9511) );
  AND U9164 ( .A(n9522), .B(n9523), .Z(n9521) );
  XOR U9165 ( .A(n9520), .B(n9184), .Z(n9523) );
  XNOR U9166 ( .A(p_input[3029]), .B(n9524), .Z(n9184) );
  AND U9167 ( .A(n242), .B(n9525), .Z(n9524) );
  XOR U9168 ( .A(p_input[3061]), .B(p_input[3029]), .Z(n9525) );
  XNOR U9169 ( .A(n9181), .B(n9520), .Z(n9522) );
  XOR U9170 ( .A(n9526), .B(n9527), .Z(n9181) );
  AND U9171 ( .A(n240), .B(n9528), .Z(n9527) );
  XOR U9172 ( .A(p_input[2997]), .B(p_input[2965]), .Z(n9528) );
  XOR U9173 ( .A(n9529), .B(n9530), .Z(n9520) );
  AND U9174 ( .A(n9531), .B(n9532), .Z(n9530) );
  XOR U9175 ( .A(n9529), .B(n9196), .Z(n9532) );
  XNOR U9176 ( .A(p_input[3028]), .B(n9533), .Z(n9196) );
  AND U9177 ( .A(n242), .B(n9534), .Z(n9533) );
  XOR U9178 ( .A(p_input[3060]), .B(p_input[3028]), .Z(n9534) );
  XNOR U9179 ( .A(n9193), .B(n9529), .Z(n9531) );
  XOR U9180 ( .A(n9535), .B(n9536), .Z(n9193) );
  AND U9181 ( .A(n240), .B(n9537), .Z(n9536) );
  XOR U9182 ( .A(p_input[2996]), .B(p_input[2964]), .Z(n9537) );
  XOR U9183 ( .A(n9538), .B(n9539), .Z(n9529) );
  AND U9184 ( .A(n9540), .B(n9541), .Z(n9539) );
  XOR U9185 ( .A(n9538), .B(n9208), .Z(n9541) );
  XNOR U9186 ( .A(p_input[3027]), .B(n9542), .Z(n9208) );
  AND U9187 ( .A(n242), .B(n9543), .Z(n9542) );
  XOR U9188 ( .A(p_input[3059]), .B(p_input[3027]), .Z(n9543) );
  XNOR U9189 ( .A(n9205), .B(n9538), .Z(n9540) );
  XOR U9190 ( .A(n9544), .B(n9545), .Z(n9205) );
  AND U9191 ( .A(n240), .B(n9546), .Z(n9545) );
  XOR U9192 ( .A(p_input[2995]), .B(p_input[2963]), .Z(n9546) );
  XOR U9193 ( .A(n9547), .B(n9548), .Z(n9538) );
  AND U9194 ( .A(n9549), .B(n9550), .Z(n9548) );
  XOR U9195 ( .A(n9547), .B(n9220), .Z(n9550) );
  XNOR U9196 ( .A(p_input[3026]), .B(n9551), .Z(n9220) );
  AND U9197 ( .A(n242), .B(n9552), .Z(n9551) );
  XOR U9198 ( .A(p_input[3058]), .B(p_input[3026]), .Z(n9552) );
  XNOR U9199 ( .A(n9217), .B(n9547), .Z(n9549) );
  XOR U9200 ( .A(n9553), .B(n9554), .Z(n9217) );
  AND U9201 ( .A(n240), .B(n9555), .Z(n9554) );
  XOR U9202 ( .A(p_input[2994]), .B(p_input[2962]), .Z(n9555) );
  XOR U9203 ( .A(n9556), .B(n9557), .Z(n9547) );
  AND U9204 ( .A(n9558), .B(n9559), .Z(n9557) );
  XOR U9205 ( .A(n9556), .B(n9232), .Z(n9559) );
  XNOR U9206 ( .A(p_input[3025]), .B(n9560), .Z(n9232) );
  AND U9207 ( .A(n242), .B(n9561), .Z(n9560) );
  XOR U9208 ( .A(p_input[3057]), .B(p_input[3025]), .Z(n9561) );
  XNOR U9209 ( .A(n9229), .B(n9556), .Z(n9558) );
  XOR U9210 ( .A(n9562), .B(n9563), .Z(n9229) );
  AND U9211 ( .A(n240), .B(n9564), .Z(n9563) );
  XOR U9212 ( .A(p_input[2993]), .B(p_input[2961]), .Z(n9564) );
  XOR U9213 ( .A(n9565), .B(n9566), .Z(n9556) );
  AND U9214 ( .A(n9567), .B(n9568), .Z(n9566) );
  XOR U9215 ( .A(n9565), .B(n9244), .Z(n9568) );
  XNOR U9216 ( .A(p_input[3024]), .B(n9569), .Z(n9244) );
  AND U9217 ( .A(n242), .B(n9570), .Z(n9569) );
  XOR U9218 ( .A(p_input[3056]), .B(p_input[3024]), .Z(n9570) );
  XNOR U9219 ( .A(n9241), .B(n9565), .Z(n9567) );
  XOR U9220 ( .A(n9571), .B(n9572), .Z(n9241) );
  AND U9221 ( .A(n240), .B(n9573), .Z(n9572) );
  XOR U9222 ( .A(p_input[2992]), .B(p_input[2960]), .Z(n9573) );
  XOR U9223 ( .A(n9574), .B(n9575), .Z(n9565) );
  AND U9224 ( .A(n9576), .B(n9577), .Z(n9575) );
  XOR U9225 ( .A(n9574), .B(n9256), .Z(n9577) );
  XNOR U9226 ( .A(p_input[3023]), .B(n9578), .Z(n9256) );
  AND U9227 ( .A(n242), .B(n9579), .Z(n9578) );
  XOR U9228 ( .A(p_input[3055]), .B(p_input[3023]), .Z(n9579) );
  XNOR U9229 ( .A(n9253), .B(n9574), .Z(n9576) );
  XOR U9230 ( .A(n9580), .B(n9581), .Z(n9253) );
  AND U9231 ( .A(n240), .B(n9582), .Z(n9581) );
  XOR U9232 ( .A(p_input[2991]), .B(p_input[2959]), .Z(n9582) );
  XOR U9233 ( .A(n9583), .B(n9584), .Z(n9574) );
  AND U9234 ( .A(n9585), .B(n9586), .Z(n9584) );
  XOR U9235 ( .A(n9583), .B(n9268), .Z(n9586) );
  XNOR U9236 ( .A(p_input[3022]), .B(n9587), .Z(n9268) );
  AND U9237 ( .A(n242), .B(n9588), .Z(n9587) );
  XOR U9238 ( .A(p_input[3054]), .B(p_input[3022]), .Z(n9588) );
  XNOR U9239 ( .A(n9265), .B(n9583), .Z(n9585) );
  XOR U9240 ( .A(n9589), .B(n9590), .Z(n9265) );
  AND U9241 ( .A(n240), .B(n9591), .Z(n9590) );
  XOR U9242 ( .A(p_input[2990]), .B(p_input[2958]), .Z(n9591) );
  XOR U9243 ( .A(n9592), .B(n9593), .Z(n9583) );
  AND U9244 ( .A(n9594), .B(n9595), .Z(n9593) );
  XOR U9245 ( .A(n9592), .B(n9280), .Z(n9595) );
  XNOR U9246 ( .A(p_input[3021]), .B(n9596), .Z(n9280) );
  AND U9247 ( .A(n242), .B(n9597), .Z(n9596) );
  XOR U9248 ( .A(p_input[3053]), .B(p_input[3021]), .Z(n9597) );
  XNOR U9249 ( .A(n9277), .B(n9592), .Z(n9594) );
  XOR U9250 ( .A(n9598), .B(n9599), .Z(n9277) );
  AND U9251 ( .A(n240), .B(n9600), .Z(n9599) );
  XOR U9252 ( .A(p_input[2989]), .B(p_input[2957]), .Z(n9600) );
  XOR U9253 ( .A(n9601), .B(n9602), .Z(n9592) );
  AND U9254 ( .A(n9603), .B(n9604), .Z(n9602) );
  XOR U9255 ( .A(n9601), .B(n9292), .Z(n9604) );
  XNOR U9256 ( .A(p_input[3020]), .B(n9605), .Z(n9292) );
  AND U9257 ( .A(n242), .B(n9606), .Z(n9605) );
  XOR U9258 ( .A(p_input[3052]), .B(p_input[3020]), .Z(n9606) );
  XNOR U9259 ( .A(n9289), .B(n9601), .Z(n9603) );
  XOR U9260 ( .A(n9607), .B(n9608), .Z(n9289) );
  AND U9261 ( .A(n240), .B(n9609), .Z(n9608) );
  XOR U9262 ( .A(p_input[2988]), .B(p_input[2956]), .Z(n9609) );
  XOR U9263 ( .A(n9610), .B(n9611), .Z(n9601) );
  AND U9264 ( .A(n9612), .B(n9613), .Z(n9611) );
  XOR U9265 ( .A(n9610), .B(n9304), .Z(n9613) );
  XNOR U9266 ( .A(p_input[3019]), .B(n9614), .Z(n9304) );
  AND U9267 ( .A(n242), .B(n9615), .Z(n9614) );
  XOR U9268 ( .A(p_input[3051]), .B(p_input[3019]), .Z(n9615) );
  XNOR U9269 ( .A(n9301), .B(n9610), .Z(n9612) );
  XOR U9270 ( .A(n9616), .B(n9617), .Z(n9301) );
  AND U9271 ( .A(n240), .B(n9618), .Z(n9617) );
  XOR U9272 ( .A(p_input[2987]), .B(p_input[2955]), .Z(n9618) );
  XOR U9273 ( .A(n9619), .B(n9620), .Z(n9610) );
  AND U9274 ( .A(n9621), .B(n9622), .Z(n9620) );
  XOR U9275 ( .A(n9619), .B(n9316), .Z(n9622) );
  XNOR U9276 ( .A(p_input[3018]), .B(n9623), .Z(n9316) );
  AND U9277 ( .A(n242), .B(n9624), .Z(n9623) );
  XOR U9278 ( .A(p_input[3050]), .B(p_input[3018]), .Z(n9624) );
  XNOR U9279 ( .A(n9313), .B(n9619), .Z(n9621) );
  XOR U9280 ( .A(n9625), .B(n9626), .Z(n9313) );
  AND U9281 ( .A(n240), .B(n9627), .Z(n9626) );
  XOR U9282 ( .A(p_input[2986]), .B(p_input[2954]), .Z(n9627) );
  XOR U9283 ( .A(n9628), .B(n9629), .Z(n9619) );
  AND U9284 ( .A(n9630), .B(n9631), .Z(n9629) );
  XOR U9285 ( .A(n9628), .B(n9328), .Z(n9631) );
  XNOR U9286 ( .A(p_input[3017]), .B(n9632), .Z(n9328) );
  AND U9287 ( .A(n242), .B(n9633), .Z(n9632) );
  XOR U9288 ( .A(p_input[3049]), .B(p_input[3017]), .Z(n9633) );
  XNOR U9289 ( .A(n9325), .B(n9628), .Z(n9630) );
  XOR U9290 ( .A(n9634), .B(n9635), .Z(n9325) );
  AND U9291 ( .A(n240), .B(n9636), .Z(n9635) );
  XOR U9292 ( .A(p_input[2985]), .B(p_input[2953]), .Z(n9636) );
  XOR U9293 ( .A(n9637), .B(n9638), .Z(n9628) );
  AND U9294 ( .A(n9639), .B(n9640), .Z(n9638) );
  XOR U9295 ( .A(n9637), .B(n9340), .Z(n9640) );
  XNOR U9296 ( .A(p_input[3016]), .B(n9641), .Z(n9340) );
  AND U9297 ( .A(n242), .B(n9642), .Z(n9641) );
  XOR U9298 ( .A(p_input[3048]), .B(p_input[3016]), .Z(n9642) );
  XNOR U9299 ( .A(n9337), .B(n9637), .Z(n9639) );
  XOR U9300 ( .A(n9643), .B(n9644), .Z(n9337) );
  AND U9301 ( .A(n240), .B(n9645), .Z(n9644) );
  XOR U9302 ( .A(p_input[2984]), .B(p_input[2952]), .Z(n9645) );
  XOR U9303 ( .A(n9646), .B(n9647), .Z(n9637) );
  AND U9304 ( .A(n9648), .B(n9649), .Z(n9647) );
  XOR U9305 ( .A(n9646), .B(n9352), .Z(n9649) );
  XNOR U9306 ( .A(p_input[3015]), .B(n9650), .Z(n9352) );
  AND U9307 ( .A(n242), .B(n9651), .Z(n9650) );
  XOR U9308 ( .A(p_input[3047]), .B(p_input[3015]), .Z(n9651) );
  XNOR U9309 ( .A(n9349), .B(n9646), .Z(n9648) );
  XOR U9310 ( .A(n9652), .B(n9653), .Z(n9349) );
  AND U9311 ( .A(n240), .B(n9654), .Z(n9653) );
  XOR U9312 ( .A(p_input[2983]), .B(p_input[2951]), .Z(n9654) );
  XOR U9313 ( .A(n9655), .B(n9656), .Z(n9646) );
  AND U9314 ( .A(n9657), .B(n9658), .Z(n9656) );
  XOR U9315 ( .A(n9655), .B(n9364), .Z(n9658) );
  XNOR U9316 ( .A(p_input[3014]), .B(n9659), .Z(n9364) );
  AND U9317 ( .A(n242), .B(n9660), .Z(n9659) );
  XOR U9318 ( .A(p_input[3046]), .B(p_input[3014]), .Z(n9660) );
  XNOR U9319 ( .A(n9361), .B(n9655), .Z(n9657) );
  XOR U9320 ( .A(n9661), .B(n9662), .Z(n9361) );
  AND U9321 ( .A(n240), .B(n9663), .Z(n9662) );
  XOR U9322 ( .A(p_input[2982]), .B(p_input[2950]), .Z(n9663) );
  XOR U9323 ( .A(n9664), .B(n9665), .Z(n9655) );
  AND U9324 ( .A(n9666), .B(n9667), .Z(n9665) );
  XOR U9325 ( .A(n9664), .B(n9376), .Z(n9667) );
  XNOR U9326 ( .A(p_input[3013]), .B(n9668), .Z(n9376) );
  AND U9327 ( .A(n242), .B(n9669), .Z(n9668) );
  XOR U9328 ( .A(p_input[3045]), .B(p_input[3013]), .Z(n9669) );
  XNOR U9329 ( .A(n9373), .B(n9664), .Z(n9666) );
  XOR U9330 ( .A(n9670), .B(n9671), .Z(n9373) );
  AND U9331 ( .A(n240), .B(n9672), .Z(n9671) );
  XOR U9332 ( .A(p_input[2981]), .B(p_input[2949]), .Z(n9672) );
  XOR U9333 ( .A(n9673), .B(n9674), .Z(n9664) );
  AND U9334 ( .A(n9675), .B(n9676), .Z(n9674) );
  XOR U9335 ( .A(n9673), .B(n9388), .Z(n9676) );
  XNOR U9336 ( .A(p_input[3012]), .B(n9677), .Z(n9388) );
  AND U9337 ( .A(n242), .B(n9678), .Z(n9677) );
  XOR U9338 ( .A(p_input[3044]), .B(p_input[3012]), .Z(n9678) );
  XNOR U9339 ( .A(n9385), .B(n9673), .Z(n9675) );
  XOR U9340 ( .A(n9679), .B(n9680), .Z(n9385) );
  AND U9341 ( .A(n240), .B(n9681), .Z(n9680) );
  XOR U9342 ( .A(p_input[2980]), .B(p_input[2948]), .Z(n9681) );
  XOR U9343 ( .A(n9682), .B(n9683), .Z(n9673) );
  AND U9344 ( .A(n9684), .B(n9685), .Z(n9683) );
  XOR U9345 ( .A(n9682), .B(n9400), .Z(n9685) );
  XNOR U9346 ( .A(p_input[3011]), .B(n9686), .Z(n9400) );
  AND U9347 ( .A(n242), .B(n9687), .Z(n9686) );
  XOR U9348 ( .A(p_input[3043]), .B(p_input[3011]), .Z(n9687) );
  XNOR U9349 ( .A(n9397), .B(n9682), .Z(n9684) );
  XOR U9350 ( .A(n9688), .B(n9689), .Z(n9397) );
  AND U9351 ( .A(n240), .B(n9690), .Z(n9689) );
  XOR U9352 ( .A(p_input[2979]), .B(p_input[2947]), .Z(n9690) );
  XOR U9353 ( .A(n9691), .B(n9692), .Z(n9682) );
  AND U9354 ( .A(n9693), .B(n9694), .Z(n9692) );
  XOR U9355 ( .A(n9412), .B(n9691), .Z(n9694) );
  XNOR U9356 ( .A(p_input[3010]), .B(n9695), .Z(n9412) );
  AND U9357 ( .A(n242), .B(n9696), .Z(n9695) );
  XOR U9358 ( .A(p_input[3042]), .B(p_input[3010]), .Z(n9696) );
  XNOR U9359 ( .A(n9691), .B(n9409), .Z(n9693) );
  XOR U9360 ( .A(n9697), .B(n9698), .Z(n9409) );
  AND U9361 ( .A(n240), .B(n9699), .Z(n9698) );
  XOR U9362 ( .A(p_input[2978]), .B(p_input[2946]), .Z(n9699) );
  XOR U9363 ( .A(n9700), .B(n9701), .Z(n9691) );
  AND U9364 ( .A(n9702), .B(n9703), .Z(n9701) );
  XNOR U9365 ( .A(n9704), .B(n9425), .Z(n9703) );
  XNOR U9366 ( .A(p_input[3009]), .B(n9705), .Z(n9425) );
  AND U9367 ( .A(n242), .B(n9706), .Z(n9705) );
  XNOR U9368 ( .A(p_input[3041]), .B(n9707), .Z(n9706) );
  IV U9369 ( .A(p_input[3009]), .Z(n9707) );
  XNOR U9370 ( .A(n9422), .B(n9700), .Z(n9702) );
  XNOR U9371 ( .A(p_input[2945]), .B(n9708), .Z(n9422) );
  AND U9372 ( .A(n240), .B(n9709), .Z(n9708) );
  XOR U9373 ( .A(p_input[2977]), .B(p_input[2945]), .Z(n9709) );
  IV U9374 ( .A(n9704), .Z(n9700) );
  AND U9375 ( .A(n9430), .B(n9433), .Z(n9704) );
  XOR U9376 ( .A(p_input[3008]), .B(n9710), .Z(n9433) );
  AND U9377 ( .A(n242), .B(n9711), .Z(n9710) );
  XOR U9378 ( .A(p_input[3040]), .B(p_input[3008]), .Z(n9711) );
  XOR U9379 ( .A(n9712), .B(n9713), .Z(n242) );
  AND U9380 ( .A(n9714), .B(n9715), .Z(n9713) );
  XNOR U9381 ( .A(p_input[3071]), .B(n9712), .Z(n9715) );
  XOR U9382 ( .A(n9712), .B(p_input[3039]), .Z(n9714) );
  XOR U9383 ( .A(n9716), .B(n9717), .Z(n9712) );
  AND U9384 ( .A(n9718), .B(n9719), .Z(n9717) );
  XNOR U9385 ( .A(p_input[3070]), .B(n9716), .Z(n9719) );
  XOR U9386 ( .A(n9716), .B(p_input[3038]), .Z(n9718) );
  XOR U9387 ( .A(n9720), .B(n9721), .Z(n9716) );
  AND U9388 ( .A(n9722), .B(n9723), .Z(n9721) );
  XNOR U9389 ( .A(p_input[3069]), .B(n9720), .Z(n9723) );
  XOR U9390 ( .A(n9720), .B(p_input[3037]), .Z(n9722) );
  XOR U9391 ( .A(n9724), .B(n9725), .Z(n9720) );
  AND U9392 ( .A(n9726), .B(n9727), .Z(n9725) );
  XNOR U9393 ( .A(p_input[3068]), .B(n9724), .Z(n9727) );
  XOR U9394 ( .A(n9724), .B(p_input[3036]), .Z(n9726) );
  XOR U9395 ( .A(n9728), .B(n9729), .Z(n9724) );
  AND U9396 ( .A(n9730), .B(n9731), .Z(n9729) );
  XNOR U9397 ( .A(p_input[3067]), .B(n9728), .Z(n9731) );
  XOR U9398 ( .A(n9728), .B(p_input[3035]), .Z(n9730) );
  XOR U9399 ( .A(n9732), .B(n9733), .Z(n9728) );
  AND U9400 ( .A(n9734), .B(n9735), .Z(n9733) );
  XNOR U9401 ( .A(p_input[3066]), .B(n9732), .Z(n9735) );
  XOR U9402 ( .A(n9732), .B(p_input[3034]), .Z(n9734) );
  XOR U9403 ( .A(n9736), .B(n9737), .Z(n9732) );
  AND U9404 ( .A(n9738), .B(n9739), .Z(n9737) );
  XNOR U9405 ( .A(p_input[3065]), .B(n9736), .Z(n9739) );
  XOR U9406 ( .A(n9736), .B(p_input[3033]), .Z(n9738) );
  XOR U9407 ( .A(n9740), .B(n9741), .Z(n9736) );
  AND U9408 ( .A(n9742), .B(n9743), .Z(n9741) );
  XNOR U9409 ( .A(p_input[3064]), .B(n9740), .Z(n9743) );
  XOR U9410 ( .A(n9740), .B(p_input[3032]), .Z(n9742) );
  XOR U9411 ( .A(n9744), .B(n9745), .Z(n9740) );
  AND U9412 ( .A(n9746), .B(n9747), .Z(n9745) );
  XNOR U9413 ( .A(p_input[3063]), .B(n9744), .Z(n9747) );
  XOR U9414 ( .A(n9744), .B(p_input[3031]), .Z(n9746) );
  XOR U9415 ( .A(n9748), .B(n9749), .Z(n9744) );
  AND U9416 ( .A(n9750), .B(n9751), .Z(n9749) );
  XNOR U9417 ( .A(p_input[3062]), .B(n9748), .Z(n9751) );
  XOR U9418 ( .A(n9748), .B(p_input[3030]), .Z(n9750) );
  XOR U9419 ( .A(n9752), .B(n9753), .Z(n9748) );
  AND U9420 ( .A(n9754), .B(n9755), .Z(n9753) );
  XNOR U9421 ( .A(p_input[3061]), .B(n9752), .Z(n9755) );
  XOR U9422 ( .A(n9752), .B(p_input[3029]), .Z(n9754) );
  XOR U9423 ( .A(n9756), .B(n9757), .Z(n9752) );
  AND U9424 ( .A(n9758), .B(n9759), .Z(n9757) );
  XNOR U9425 ( .A(p_input[3060]), .B(n9756), .Z(n9759) );
  XOR U9426 ( .A(n9756), .B(p_input[3028]), .Z(n9758) );
  XOR U9427 ( .A(n9760), .B(n9761), .Z(n9756) );
  AND U9428 ( .A(n9762), .B(n9763), .Z(n9761) );
  XNOR U9429 ( .A(p_input[3059]), .B(n9760), .Z(n9763) );
  XOR U9430 ( .A(n9760), .B(p_input[3027]), .Z(n9762) );
  XOR U9431 ( .A(n9764), .B(n9765), .Z(n9760) );
  AND U9432 ( .A(n9766), .B(n9767), .Z(n9765) );
  XNOR U9433 ( .A(p_input[3058]), .B(n9764), .Z(n9767) );
  XOR U9434 ( .A(n9764), .B(p_input[3026]), .Z(n9766) );
  XOR U9435 ( .A(n9768), .B(n9769), .Z(n9764) );
  AND U9436 ( .A(n9770), .B(n9771), .Z(n9769) );
  XNOR U9437 ( .A(p_input[3057]), .B(n9768), .Z(n9771) );
  XOR U9438 ( .A(n9768), .B(p_input[3025]), .Z(n9770) );
  XOR U9439 ( .A(n9772), .B(n9773), .Z(n9768) );
  AND U9440 ( .A(n9774), .B(n9775), .Z(n9773) );
  XNOR U9441 ( .A(p_input[3056]), .B(n9772), .Z(n9775) );
  XOR U9442 ( .A(n9772), .B(p_input[3024]), .Z(n9774) );
  XOR U9443 ( .A(n9776), .B(n9777), .Z(n9772) );
  AND U9444 ( .A(n9778), .B(n9779), .Z(n9777) );
  XNOR U9445 ( .A(p_input[3055]), .B(n9776), .Z(n9779) );
  XOR U9446 ( .A(n9776), .B(p_input[3023]), .Z(n9778) );
  XOR U9447 ( .A(n9780), .B(n9781), .Z(n9776) );
  AND U9448 ( .A(n9782), .B(n9783), .Z(n9781) );
  XNOR U9449 ( .A(p_input[3054]), .B(n9780), .Z(n9783) );
  XOR U9450 ( .A(n9780), .B(p_input[3022]), .Z(n9782) );
  XOR U9451 ( .A(n9784), .B(n9785), .Z(n9780) );
  AND U9452 ( .A(n9786), .B(n9787), .Z(n9785) );
  XNOR U9453 ( .A(p_input[3053]), .B(n9784), .Z(n9787) );
  XOR U9454 ( .A(n9784), .B(p_input[3021]), .Z(n9786) );
  XOR U9455 ( .A(n9788), .B(n9789), .Z(n9784) );
  AND U9456 ( .A(n9790), .B(n9791), .Z(n9789) );
  XNOR U9457 ( .A(p_input[3052]), .B(n9788), .Z(n9791) );
  XOR U9458 ( .A(n9788), .B(p_input[3020]), .Z(n9790) );
  XOR U9459 ( .A(n9792), .B(n9793), .Z(n9788) );
  AND U9460 ( .A(n9794), .B(n9795), .Z(n9793) );
  XNOR U9461 ( .A(p_input[3051]), .B(n9792), .Z(n9795) );
  XOR U9462 ( .A(n9792), .B(p_input[3019]), .Z(n9794) );
  XOR U9463 ( .A(n9796), .B(n9797), .Z(n9792) );
  AND U9464 ( .A(n9798), .B(n9799), .Z(n9797) );
  XNOR U9465 ( .A(p_input[3050]), .B(n9796), .Z(n9799) );
  XOR U9466 ( .A(n9796), .B(p_input[3018]), .Z(n9798) );
  XOR U9467 ( .A(n9800), .B(n9801), .Z(n9796) );
  AND U9468 ( .A(n9802), .B(n9803), .Z(n9801) );
  XNOR U9469 ( .A(p_input[3049]), .B(n9800), .Z(n9803) );
  XOR U9470 ( .A(n9800), .B(p_input[3017]), .Z(n9802) );
  XOR U9471 ( .A(n9804), .B(n9805), .Z(n9800) );
  AND U9472 ( .A(n9806), .B(n9807), .Z(n9805) );
  XNOR U9473 ( .A(p_input[3048]), .B(n9804), .Z(n9807) );
  XOR U9474 ( .A(n9804), .B(p_input[3016]), .Z(n9806) );
  XOR U9475 ( .A(n9808), .B(n9809), .Z(n9804) );
  AND U9476 ( .A(n9810), .B(n9811), .Z(n9809) );
  XNOR U9477 ( .A(p_input[3047]), .B(n9808), .Z(n9811) );
  XOR U9478 ( .A(n9808), .B(p_input[3015]), .Z(n9810) );
  XOR U9479 ( .A(n9812), .B(n9813), .Z(n9808) );
  AND U9480 ( .A(n9814), .B(n9815), .Z(n9813) );
  XNOR U9481 ( .A(p_input[3046]), .B(n9812), .Z(n9815) );
  XOR U9482 ( .A(n9812), .B(p_input[3014]), .Z(n9814) );
  XOR U9483 ( .A(n9816), .B(n9817), .Z(n9812) );
  AND U9484 ( .A(n9818), .B(n9819), .Z(n9817) );
  XNOR U9485 ( .A(p_input[3045]), .B(n9816), .Z(n9819) );
  XOR U9486 ( .A(n9816), .B(p_input[3013]), .Z(n9818) );
  XOR U9487 ( .A(n9820), .B(n9821), .Z(n9816) );
  AND U9488 ( .A(n9822), .B(n9823), .Z(n9821) );
  XNOR U9489 ( .A(p_input[3044]), .B(n9820), .Z(n9823) );
  XOR U9490 ( .A(n9820), .B(p_input[3012]), .Z(n9822) );
  XOR U9491 ( .A(n9824), .B(n9825), .Z(n9820) );
  AND U9492 ( .A(n9826), .B(n9827), .Z(n9825) );
  XNOR U9493 ( .A(p_input[3043]), .B(n9824), .Z(n9827) );
  XOR U9494 ( .A(n9824), .B(p_input[3011]), .Z(n9826) );
  XOR U9495 ( .A(n9828), .B(n9829), .Z(n9824) );
  AND U9496 ( .A(n9830), .B(n9831), .Z(n9829) );
  XNOR U9497 ( .A(p_input[3042]), .B(n9828), .Z(n9831) );
  XOR U9498 ( .A(n9828), .B(p_input[3010]), .Z(n9830) );
  XNOR U9499 ( .A(n9832), .B(n9833), .Z(n9828) );
  AND U9500 ( .A(n9834), .B(n9835), .Z(n9833) );
  XOR U9501 ( .A(p_input[3041]), .B(n9832), .Z(n9835) );
  XNOR U9502 ( .A(p_input[3009]), .B(n9832), .Z(n9834) );
  AND U9503 ( .A(p_input[3040]), .B(n9836), .Z(n9832) );
  IV U9504 ( .A(p_input[3008]), .Z(n9836) );
  XNOR U9505 ( .A(p_input[2944]), .B(n9837), .Z(n9430) );
  AND U9506 ( .A(n240), .B(n9838), .Z(n9837) );
  XOR U9507 ( .A(p_input[2976]), .B(p_input[2944]), .Z(n9838) );
  XOR U9508 ( .A(n9839), .B(n9840), .Z(n240) );
  AND U9509 ( .A(n9841), .B(n9842), .Z(n9840) );
  XNOR U9510 ( .A(p_input[3007]), .B(n9839), .Z(n9842) );
  XOR U9511 ( .A(n9839), .B(p_input[2975]), .Z(n9841) );
  XOR U9512 ( .A(n9843), .B(n9844), .Z(n9839) );
  AND U9513 ( .A(n9845), .B(n9846), .Z(n9844) );
  XNOR U9514 ( .A(p_input[3006]), .B(n9843), .Z(n9846) );
  XNOR U9515 ( .A(n9843), .B(n9445), .Z(n9845) );
  IV U9516 ( .A(p_input[2974]), .Z(n9445) );
  XOR U9517 ( .A(n9847), .B(n9848), .Z(n9843) );
  AND U9518 ( .A(n9849), .B(n9850), .Z(n9848) );
  XNOR U9519 ( .A(p_input[3005]), .B(n9847), .Z(n9850) );
  XNOR U9520 ( .A(n9847), .B(n9454), .Z(n9849) );
  IV U9521 ( .A(p_input[2973]), .Z(n9454) );
  XOR U9522 ( .A(n9851), .B(n9852), .Z(n9847) );
  AND U9523 ( .A(n9853), .B(n9854), .Z(n9852) );
  XNOR U9524 ( .A(p_input[3004]), .B(n9851), .Z(n9854) );
  XNOR U9525 ( .A(n9851), .B(n9463), .Z(n9853) );
  IV U9526 ( .A(p_input[2972]), .Z(n9463) );
  XOR U9527 ( .A(n9855), .B(n9856), .Z(n9851) );
  AND U9528 ( .A(n9857), .B(n9858), .Z(n9856) );
  XNOR U9529 ( .A(p_input[3003]), .B(n9855), .Z(n9858) );
  XNOR U9530 ( .A(n9855), .B(n9472), .Z(n9857) );
  IV U9531 ( .A(p_input[2971]), .Z(n9472) );
  XOR U9532 ( .A(n9859), .B(n9860), .Z(n9855) );
  AND U9533 ( .A(n9861), .B(n9862), .Z(n9860) );
  XNOR U9534 ( .A(p_input[3002]), .B(n9859), .Z(n9862) );
  XNOR U9535 ( .A(n9859), .B(n9481), .Z(n9861) );
  IV U9536 ( .A(p_input[2970]), .Z(n9481) );
  XOR U9537 ( .A(n9863), .B(n9864), .Z(n9859) );
  AND U9538 ( .A(n9865), .B(n9866), .Z(n9864) );
  XNOR U9539 ( .A(p_input[3001]), .B(n9863), .Z(n9866) );
  XNOR U9540 ( .A(n9863), .B(n9490), .Z(n9865) );
  IV U9541 ( .A(p_input[2969]), .Z(n9490) );
  XOR U9542 ( .A(n9867), .B(n9868), .Z(n9863) );
  AND U9543 ( .A(n9869), .B(n9870), .Z(n9868) );
  XNOR U9544 ( .A(p_input[3000]), .B(n9867), .Z(n9870) );
  XNOR U9545 ( .A(n9867), .B(n9499), .Z(n9869) );
  IV U9546 ( .A(p_input[2968]), .Z(n9499) );
  XOR U9547 ( .A(n9871), .B(n9872), .Z(n9867) );
  AND U9548 ( .A(n9873), .B(n9874), .Z(n9872) );
  XNOR U9549 ( .A(p_input[2999]), .B(n9871), .Z(n9874) );
  XNOR U9550 ( .A(n9871), .B(n9508), .Z(n9873) );
  IV U9551 ( .A(p_input[2967]), .Z(n9508) );
  XOR U9552 ( .A(n9875), .B(n9876), .Z(n9871) );
  AND U9553 ( .A(n9877), .B(n9878), .Z(n9876) );
  XNOR U9554 ( .A(p_input[2998]), .B(n9875), .Z(n9878) );
  XNOR U9555 ( .A(n9875), .B(n9517), .Z(n9877) );
  IV U9556 ( .A(p_input[2966]), .Z(n9517) );
  XOR U9557 ( .A(n9879), .B(n9880), .Z(n9875) );
  AND U9558 ( .A(n9881), .B(n9882), .Z(n9880) );
  XNOR U9559 ( .A(p_input[2997]), .B(n9879), .Z(n9882) );
  XNOR U9560 ( .A(n9879), .B(n9526), .Z(n9881) );
  IV U9561 ( .A(p_input[2965]), .Z(n9526) );
  XOR U9562 ( .A(n9883), .B(n9884), .Z(n9879) );
  AND U9563 ( .A(n9885), .B(n9886), .Z(n9884) );
  XNOR U9564 ( .A(p_input[2996]), .B(n9883), .Z(n9886) );
  XNOR U9565 ( .A(n9883), .B(n9535), .Z(n9885) );
  IV U9566 ( .A(p_input[2964]), .Z(n9535) );
  XOR U9567 ( .A(n9887), .B(n9888), .Z(n9883) );
  AND U9568 ( .A(n9889), .B(n9890), .Z(n9888) );
  XNOR U9569 ( .A(p_input[2995]), .B(n9887), .Z(n9890) );
  XNOR U9570 ( .A(n9887), .B(n9544), .Z(n9889) );
  IV U9571 ( .A(p_input[2963]), .Z(n9544) );
  XOR U9572 ( .A(n9891), .B(n9892), .Z(n9887) );
  AND U9573 ( .A(n9893), .B(n9894), .Z(n9892) );
  XNOR U9574 ( .A(p_input[2994]), .B(n9891), .Z(n9894) );
  XNOR U9575 ( .A(n9891), .B(n9553), .Z(n9893) );
  IV U9576 ( .A(p_input[2962]), .Z(n9553) );
  XOR U9577 ( .A(n9895), .B(n9896), .Z(n9891) );
  AND U9578 ( .A(n9897), .B(n9898), .Z(n9896) );
  XNOR U9579 ( .A(p_input[2993]), .B(n9895), .Z(n9898) );
  XNOR U9580 ( .A(n9895), .B(n9562), .Z(n9897) );
  IV U9581 ( .A(p_input[2961]), .Z(n9562) );
  XOR U9582 ( .A(n9899), .B(n9900), .Z(n9895) );
  AND U9583 ( .A(n9901), .B(n9902), .Z(n9900) );
  XNOR U9584 ( .A(p_input[2992]), .B(n9899), .Z(n9902) );
  XNOR U9585 ( .A(n9899), .B(n9571), .Z(n9901) );
  IV U9586 ( .A(p_input[2960]), .Z(n9571) );
  XOR U9587 ( .A(n9903), .B(n9904), .Z(n9899) );
  AND U9588 ( .A(n9905), .B(n9906), .Z(n9904) );
  XNOR U9589 ( .A(p_input[2991]), .B(n9903), .Z(n9906) );
  XNOR U9590 ( .A(n9903), .B(n9580), .Z(n9905) );
  IV U9591 ( .A(p_input[2959]), .Z(n9580) );
  XOR U9592 ( .A(n9907), .B(n9908), .Z(n9903) );
  AND U9593 ( .A(n9909), .B(n9910), .Z(n9908) );
  XNOR U9594 ( .A(p_input[2990]), .B(n9907), .Z(n9910) );
  XNOR U9595 ( .A(n9907), .B(n9589), .Z(n9909) );
  IV U9596 ( .A(p_input[2958]), .Z(n9589) );
  XOR U9597 ( .A(n9911), .B(n9912), .Z(n9907) );
  AND U9598 ( .A(n9913), .B(n9914), .Z(n9912) );
  XNOR U9599 ( .A(p_input[2989]), .B(n9911), .Z(n9914) );
  XNOR U9600 ( .A(n9911), .B(n9598), .Z(n9913) );
  IV U9601 ( .A(p_input[2957]), .Z(n9598) );
  XOR U9602 ( .A(n9915), .B(n9916), .Z(n9911) );
  AND U9603 ( .A(n9917), .B(n9918), .Z(n9916) );
  XNOR U9604 ( .A(p_input[2988]), .B(n9915), .Z(n9918) );
  XNOR U9605 ( .A(n9915), .B(n9607), .Z(n9917) );
  IV U9606 ( .A(p_input[2956]), .Z(n9607) );
  XOR U9607 ( .A(n9919), .B(n9920), .Z(n9915) );
  AND U9608 ( .A(n9921), .B(n9922), .Z(n9920) );
  XNOR U9609 ( .A(p_input[2987]), .B(n9919), .Z(n9922) );
  XNOR U9610 ( .A(n9919), .B(n9616), .Z(n9921) );
  IV U9611 ( .A(p_input[2955]), .Z(n9616) );
  XOR U9612 ( .A(n9923), .B(n9924), .Z(n9919) );
  AND U9613 ( .A(n9925), .B(n9926), .Z(n9924) );
  XNOR U9614 ( .A(p_input[2986]), .B(n9923), .Z(n9926) );
  XNOR U9615 ( .A(n9923), .B(n9625), .Z(n9925) );
  IV U9616 ( .A(p_input[2954]), .Z(n9625) );
  XOR U9617 ( .A(n9927), .B(n9928), .Z(n9923) );
  AND U9618 ( .A(n9929), .B(n9930), .Z(n9928) );
  XNOR U9619 ( .A(p_input[2985]), .B(n9927), .Z(n9930) );
  XNOR U9620 ( .A(n9927), .B(n9634), .Z(n9929) );
  IV U9621 ( .A(p_input[2953]), .Z(n9634) );
  XOR U9622 ( .A(n9931), .B(n9932), .Z(n9927) );
  AND U9623 ( .A(n9933), .B(n9934), .Z(n9932) );
  XNOR U9624 ( .A(p_input[2984]), .B(n9931), .Z(n9934) );
  XNOR U9625 ( .A(n9931), .B(n9643), .Z(n9933) );
  IV U9626 ( .A(p_input[2952]), .Z(n9643) );
  XOR U9627 ( .A(n9935), .B(n9936), .Z(n9931) );
  AND U9628 ( .A(n9937), .B(n9938), .Z(n9936) );
  XNOR U9629 ( .A(p_input[2983]), .B(n9935), .Z(n9938) );
  XNOR U9630 ( .A(n9935), .B(n9652), .Z(n9937) );
  IV U9631 ( .A(p_input[2951]), .Z(n9652) );
  XOR U9632 ( .A(n9939), .B(n9940), .Z(n9935) );
  AND U9633 ( .A(n9941), .B(n9942), .Z(n9940) );
  XNOR U9634 ( .A(p_input[2982]), .B(n9939), .Z(n9942) );
  XNOR U9635 ( .A(n9939), .B(n9661), .Z(n9941) );
  IV U9636 ( .A(p_input[2950]), .Z(n9661) );
  XOR U9637 ( .A(n9943), .B(n9944), .Z(n9939) );
  AND U9638 ( .A(n9945), .B(n9946), .Z(n9944) );
  XNOR U9639 ( .A(p_input[2981]), .B(n9943), .Z(n9946) );
  XNOR U9640 ( .A(n9943), .B(n9670), .Z(n9945) );
  IV U9641 ( .A(p_input[2949]), .Z(n9670) );
  XOR U9642 ( .A(n9947), .B(n9948), .Z(n9943) );
  AND U9643 ( .A(n9949), .B(n9950), .Z(n9948) );
  XNOR U9644 ( .A(p_input[2980]), .B(n9947), .Z(n9950) );
  XNOR U9645 ( .A(n9947), .B(n9679), .Z(n9949) );
  IV U9646 ( .A(p_input[2948]), .Z(n9679) );
  XOR U9647 ( .A(n9951), .B(n9952), .Z(n9947) );
  AND U9648 ( .A(n9953), .B(n9954), .Z(n9952) );
  XNOR U9649 ( .A(p_input[2979]), .B(n9951), .Z(n9954) );
  XNOR U9650 ( .A(n9951), .B(n9688), .Z(n9953) );
  IV U9651 ( .A(p_input[2947]), .Z(n9688) );
  XOR U9652 ( .A(n9955), .B(n9956), .Z(n9951) );
  AND U9653 ( .A(n9957), .B(n9958), .Z(n9956) );
  XNOR U9654 ( .A(p_input[2978]), .B(n9955), .Z(n9958) );
  XNOR U9655 ( .A(n9955), .B(n9697), .Z(n9957) );
  IV U9656 ( .A(p_input[2946]), .Z(n9697) );
  XNOR U9657 ( .A(n9959), .B(n9960), .Z(n9955) );
  AND U9658 ( .A(n9961), .B(n9962), .Z(n9960) );
  XOR U9659 ( .A(p_input[2977]), .B(n9959), .Z(n9962) );
  XNOR U9660 ( .A(p_input[2945]), .B(n9959), .Z(n9961) );
  AND U9661 ( .A(p_input[2976]), .B(n9963), .Z(n9959) );
  IV U9662 ( .A(p_input[2944]), .Z(n9963) );
  XOR U9663 ( .A(n9964), .B(n9965), .Z(n9053) );
  AND U9664 ( .A(n332), .B(n9966), .Z(n9965) );
  XNOR U9665 ( .A(n9967), .B(n9964), .Z(n9966) );
  XOR U9666 ( .A(n9968), .B(n9969), .Z(n332) );
  AND U9667 ( .A(n9970), .B(n9971), .Z(n9969) );
  XNOR U9668 ( .A(n9068), .B(n9968), .Z(n9971) );
  AND U9669 ( .A(p_input[2943]), .B(p_input[2911]), .Z(n9068) );
  XNOR U9670 ( .A(n9968), .B(n9065), .Z(n9970) );
  IV U9671 ( .A(n9972), .Z(n9065) );
  AND U9672 ( .A(p_input[2847]), .B(p_input[2879]), .Z(n9972) );
  XOR U9673 ( .A(n9973), .B(n9974), .Z(n9968) );
  AND U9674 ( .A(n9975), .B(n9976), .Z(n9974) );
  XOR U9675 ( .A(n9973), .B(n9080), .Z(n9976) );
  XNOR U9676 ( .A(p_input[2910]), .B(n9977), .Z(n9080) );
  AND U9677 ( .A(n246), .B(n9978), .Z(n9977) );
  XOR U9678 ( .A(p_input[2942]), .B(p_input[2910]), .Z(n9978) );
  XNOR U9679 ( .A(n9077), .B(n9973), .Z(n9975) );
  XOR U9680 ( .A(n9979), .B(n9980), .Z(n9077) );
  AND U9681 ( .A(n243), .B(n9981), .Z(n9980) );
  XOR U9682 ( .A(p_input[2878]), .B(p_input[2846]), .Z(n9981) );
  XOR U9683 ( .A(n9982), .B(n9983), .Z(n9973) );
  AND U9684 ( .A(n9984), .B(n9985), .Z(n9983) );
  XOR U9685 ( .A(n9982), .B(n9092), .Z(n9985) );
  XNOR U9686 ( .A(p_input[2909]), .B(n9986), .Z(n9092) );
  AND U9687 ( .A(n246), .B(n9987), .Z(n9986) );
  XOR U9688 ( .A(p_input[2941]), .B(p_input[2909]), .Z(n9987) );
  XNOR U9689 ( .A(n9089), .B(n9982), .Z(n9984) );
  XOR U9690 ( .A(n9988), .B(n9989), .Z(n9089) );
  AND U9691 ( .A(n243), .B(n9990), .Z(n9989) );
  XOR U9692 ( .A(p_input[2877]), .B(p_input[2845]), .Z(n9990) );
  XOR U9693 ( .A(n9991), .B(n9992), .Z(n9982) );
  AND U9694 ( .A(n9993), .B(n9994), .Z(n9992) );
  XOR U9695 ( .A(n9991), .B(n9104), .Z(n9994) );
  XNOR U9696 ( .A(p_input[2908]), .B(n9995), .Z(n9104) );
  AND U9697 ( .A(n246), .B(n9996), .Z(n9995) );
  XOR U9698 ( .A(p_input[2940]), .B(p_input[2908]), .Z(n9996) );
  XNOR U9699 ( .A(n9101), .B(n9991), .Z(n9993) );
  XOR U9700 ( .A(n9997), .B(n9998), .Z(n9101) );
  AND U9701 ( .A(n243), .B(n9999), .Z(n9998) );
  XOR U9702 ( .A(p_input[2876]), .B(p_input[2844]), .Z(n9999) );
  XOR U9703 ( .A(n10000), .B(n10001), .Z(n9991) );
  AND U9704 ( .A(n10002), .B(n10003), .Z(n10001) );
  XOR U9705 ( .A(n10000), .B(n9116), .Z(n10003) );
  XNOR U9706 ( .A(p_input[2907]), .B(n10004), .Z(n9116) );
  AND U9707 ( .A(n246), .B(n10005), .Z(n10004) );
  XOR U9708 ( .A(p_input[2939]), .B(p_input[2907]), .Z(n10005) );
  XNOR U9709 ( .A(n9113), .B(n10000), .Z(n10002) );
  XOR U9710 ( .A(n10006), .B(n10007), .Z(n9113) );
  AND U9711 ( .A(n243), .B(n10008), .Z(n10007) );
  XOR U9712 ( .A(p_input[2875]), .B(p_input[2843]), .Z(n10008) );
  XOR U9713 ( .A(n10009), .B(n10010), .Z(n10000) );
  AND U9714 ( .A(n10011), .B(n10012), .Z(n10010) );
  XOR U9715 ( .A(n10009), .B(n9128), .Z(n10012) );
  XNOR U9716 ( .A(p_input[2906]), .B(n10013), .Z(n9128) );
  AND U9717 ( .A(n246), .B(n10014), .Z(n10013) );
  XOR U9718 ( .A(p_input[2938]), .B(p_input[2906]), .Z(n10014) );
  XNOR U9719 ( .A(n9125), .B(n10009), .Z(n10011) );
  XOR U9720 ( .A(n10015), .B(n10016), .Z(n9125) );
  AND U9721 ( .A(n243), .B(n10017), .Z(n10016) );
  XOR U9722 ( .A(p_input[2874]), .B(p_input[2842]), .Z(n10017) );
  XOR U9723 ( .A(n10018), .B(n10019), .Z(n10009) );
  AND U9724 ( .A(n10020), .B(n10021), .Z(n10019) );
  XOR U9725 ( .A(n10018), .B(n9140), .Z(n10021) );
  XNOR U9726 ( .A(p_input[2905]), .B(n10022), .Z(n9140) );
  AND U9727 ( .A(n246), .B(n10023), .Z(n10022) );
  XOR U9728 ( .A(p_input[2937]), .B(p_input[2905]), .Z(n10023) );
  XNOR U9729 ( .A(n9137), .B(n10018), .Z(n10020) );
  XOR U9730 ( .A(n10024), .B(n10025), .Z(n9137) );
  AND U9731 ( .A(n243), .B(n10026), .Z(n10025) );
  XOR U9732 ( .A(p_input[2873]), .B(p_input[2841]), .Z(n10026) );
  XOR U9733 ( .A(n10027), .B(n10028), .Z(n10018) );
  AND U9734 ( .A(n10029), .B(n10030), .Z(n10028) );
  XOR U9735 ( .A(n10027), .B(n9152), .Z(n10030) );
  XNOR U9736 ( .A(p_input[2904]), .B(n10031), .Z(n9152) );
  AND U9737 ( .A(n246), .B(n10032), .Z(n10031) );
  XOR U9738 ( .A(p_input[2936]), .B(p_input[2904]), .Z(n10032) );
  XNOR U9739 ( .A(n9149), .B(n10027), .Z(n10029) );
  XOR U9740 ( .A(n10033), .B(n10034), .Z(n9149) );
  AND U9741 ( .A(n243), .B(n10035), .Z(n10034) );
  XOR U9742 ( .A(p_input[2872]), .B(p_input[2840]), .Z(n10035) );
  XOR U9743 ( .A(n10036), .B(n10037), .Z(n10027) );
  AND U9744 ( .A(n10038), .B(n10039), .Z(n10037) );
  XOR U9745 ( .A(n10036), .B(n9164), .Z(n10039) );
  XNOR U9746 ( .A(p_input[2903]), .B(n10040), .Z(n9164) );
  AND U9747 ( .A(n246), .B(n10041), .Z(n10040) );
  XOR U9748 ( .A(p_input[2935]), .B(p_input[2903]), .Z(n10041) );
  XNOR U9749 ( .A(n9161), .B(n10036), .Z(n10038) );
  XOR U9750 ( .A(n10042), .B(n10043), .Z(n9161) );
  AND U9751 ( .A(n243), .B(n10044), .Z(n10043) );
  XOR U9752 ( .A(p_input[2871]), .B(p_input[2839]), .Z(n10044) );
  XOR U9753 ( .A(n10045), .B(n10046), .Z(n10036) );
  AND U9754 ( .A(n10047), .B(n10048), .Z(n10046) );
  XOR U9755 ( .A(n10045), .B(n9176), .Z(n10048) );
  XNOR U9756 ( .A(p_input[2902]), .B(n10049), .Z(n9176) );
  AND U9757 ( .A(n246), .B(n10050), .Z(n10049) );
  XOR U9758 ( .A(p_input[2934]), .B(p_input[2902]), .Z(n10050) );
  XNOR U9759 ( .A(n9173), .B(n10045), .Z(n10047) );
  XOR U9760 ( .A(n10051), .B(n10052), .Z(n9173) );
  AND U9761 ( .A(n243), .B(n10053), .Z(n10052) );
  XOR U9762 ( .A(p_input[2870]), .B(p_input[2838]), .Z(n10053) );
  XOR U9763 ( .A(n10054), .B(n10055), .Z(n10045) );
  AND U9764 ( .A(n10056), .B(n10057), .Z(n10055) );
  XOR U9765 ( .A(n10054), .B(n9188), .Z(n10057) );
  XNOR U9766 ( .A(p_input[2901]), .B(n10058), .Z(n9188) );
  AND U9767 ( .A(n246), .B(n10059), .Z(n10058) );
  XOR U9768 ( .A(p_input[2933]), .B(p_input[2901]), .Z(n10059) );
  XNOR U9769 ( .A(n9185), .B(n10054), .Z(n10056) );
  XOR U9770 ( .A(n10060), .B(n10061), .Z(n9185) );
  AND U9771 ( .A(n243), .B(n10062), .Z(n10061) );
  XOR U9772 ( .A(p_input[2869]), .B(p_input[2837]), .Z(n10062) );
  XOR U9773 ( .A(n10063), .B(n10064), .Z(n10054) );
  AND U9774 ( .A(n10065), .B(n10066), .Z(n10064) );
  XOR U9775 ( .A(n10063), .B(n9200), .Z(n10066) );
  XNOR U9776 ( .A(p_input[2900]), .B(n10067), .Z(n9200) );
  AND U9777 ( .A(n246), .B(n10068), .Z(n10067) );
  XOR U9778 ( .A(p_input[2932]), .B(p_input[2900]), .Z(n10068) );
  XNOR U9779 ( .A(n9197), .B(n10063), .Z(n10065) );
  XOR U9780 ( .A(n10069), .B(n10070), .Z(n9197) );
  AND U9781 ( .A(n243), .B(n10071), .Z(n10070) );
  XOR U9782 ( .A(p_input[2868]), .B(p_input[2836]), .Z(n10071) );
  XOR U9783 ( .A(n10072), .B(n10073), .Z(n10063) );
  AND U9784 ( .A(n10074), .B(n10075), .Z(n10073) );
  XOR U9785 ( .A(n10072), .B(n9212), .Z(n10075) );
  XNOR U9786 ( .A(p_input[2899]), .B(n10076), .Z(n9212) );
  AND U9787 ( .A(n246), .B(n10077), .Z(n10076) );
  XOR U9788 ( .A(p_input[2931]), .B(p_input[2899]), .Z(n10077) );
  XNOR U9789 ( .A(n9209), .B(n10072), .Z(n10074) );
  XOR U9790 ( .A(n10078), .B(n10079), .Z(n9209) );
  AND U9791 ( .A(n243), .B(n10080), .Z(n10079) );
  XOR U9792 ( .A(p_input[2867]), .B(p_input[2835]), .Z(n10080) );
  XOR U9793 ( .A(n10081), .B(n10082), .Z(n10072) );
  AND U9794 ( .A(n10083), .B(n10084), .Z(n10082) );
  XOR U9795 ( .A(n10081), .B(n9224), .Z(n10084) );
  XNOR U9796 ( .A(p_input[2898]), .B(n10085), .Z(n9224) );
  AND U9797 ( .A(n246), .B(n10086), .Z(n10085) );
  XOR U9798 ( .A(p_input[2930]), .B(p_input[2898]), .Z(n10086) );
  XNOR U9799 ( .A(n9221), .B(n10081), .Z(n10083) );
  XOR U9800 ( .A(n10087), .B(n10088), .Z(n9221) );
  AND U9801 ( .A(n243), .B(n10089), .Z(n10088) );
  XOR U9802 ( .A(p_input[2866]), .B(p_input[2834]), .Z(n10089) );
  XOR U9803 ( .A(n10090), .B(n10091), .Z(n10081) );
  AND U9804 ( .A(n10092), .B(n10093), .Z(n10091) );
  XOR U9805 ( .A(n10090), .B(n9236), .Z(n10093) );
  XNOR U9806 ( .A(p_input[2897]), .B(n10094), .Z(n9236) );
  AND U9807 ( .A(n246), .B(n10095), .Z(n10094) );
  XOR U9808 ( .A(p_input[2929]), .B(p_input[2897]), .Z(n10095) );
  XNOR U9809 ( .A(n9233), .B(n10090), .Z(n10092) );
  XOR U9810 ( .A(n10096), .B(n10097), .Z(n9233) );
  AND U9811 ( .A(n243), .B(n10098), .Z(n10097) );
  XOR U9812 ( .A(p_input[2865]), .B(p_input[2833]), .Z(n10098) );
  XOR U9813 ( .A(n10099), .B(n10100), .Z(n10090) );
  AND U9814 ( .A(n10101), .B(n10102), .Z(n10100) );
  XOR U9815 ( .A(n10099), .B(n9248), .Z(n10102) );
  XNOR U9816 ( .A(p_input[2896]), .B(n10103), .Z(n9248) );
  AND U9817 ( .A(n246), .B(n10104), .Z(n10103) );
  XOR U9818 ( .A(p_input[2928]), .B(p_input[2896]), .Z(n10104) );
  XNOR U9819 ( .A(n9245), .B(n10099), .Z(n10101) );
  XOR U9820 ( .A(n10105), .B(n10106), .Z(n9245) );
  AND U9821 ( .A(n243), .B(n10107), .Z(n10106) );
  XOR U9822 ( .A(p_input[2864]), .B(p_input[2832]), .Z(n10107) );
  XOR U9823 ( .A(n10108), .B(n10109), .Z(n10099) );
  AND U9824 ( .A(n10110), .B(n10111), .Z(n10109) );
  XOR U9825 ( .A(n10108), .B(n9260), .Z(n10111) );
  XNOR U9826 ( .A(p_input[2895]), .B(n10112), .Z(n9260) );
  AND U9827 ( .A(n246), .B(n10113), .Z(n10112) );
  XOR U9828 ( .A(p_input[2927]), .B(p_input[2895]), .Z(n10113) );
  XNOR U9829 ( .A(n9257), .B(n10108), .Z(n10110) );
  XOR U9830 ( .A(n10114), .B(n10115), .Z(n9257) );
  AND U9831 ( .A(n243), .B(n10116), .Z(n10115) );
  XOR U9832 ( .A(p_input[2863]), .B(p_input[2831]), .Z(n10116) );
  XOR U9833 ( .A(n10117), .B(n10118), .Z(n10108) );
  AND U9834 ( .A(n10119), .B(n10120), .Z(n10118) );
  XOR U9835 ( .A(n10117), .B(n9272), .Z(n10120) );
  XNOR U9836 ( .A(p_input[2894]), .B(n10121), .Z(n9272) );
  AND U9837 ( .A(n246), .B(n10122), .Z(n10121) );
  XOR U9838 ( .A(p_input[2926]), .B(p_input[2894]), .Z(n10122) );
  XNOR U9839 ( .A(n9269), .B(n10117), .Z(n10119) );
  XOR U9840 ( .A(n10123), .B(n10124), .Z(n9269) );
  AND U9841 ( .A(n243), .B(n10125), .Z(n10124) );
  XOR U9842 ( .A(p_input[2862]), .B(p_input[2830]), .Z(n10125) );
  XOR U9843 ( .A(n10126), .B(n10127), .Z(n10117) );
  AND U9844 ( .A(n10128), .B(n10129), .Z(n10127) );
  XOR U9845 ( .A(n10126), .B(n9284), .Z(n10129) );
  XNOR U9846 ( .A(p_input[2893]), .B(n10130), .Z(n9284) );
  AND U9847 ( .A(n246), .B(n10131), .Z(n10130) );
  XOR U9848 ( .A(p_input[2925]), .B(p_input[2893]), .Z(n10131) );
  XNOR U9849 ( .A(n9281), .B(n10126), .Z(n10128) );
  XOR U9850 ( .A(n10132), .B(n10133), .Z(n9281) );
  AND U9851 ( .A(n243), .B(n10134), .Z(n10133) );
  XOR U9852 ( .A(p_input[2861]), .B(p_input[2829]), .Z(n10134) );
  XOR U9853 ( .A(n10135), .B(n10136), .Z(n10126) );
  AND U9854 ( .A(n10137), .B(n10138), .Z(n10136) );
  XOR U9855 ( .A(n10135), .B(n9296), .Z(n10138) );
  XNOR U9856 ( .A(p_input[2892]), .B(n10139), .Z(n9296) );
  AND U9857 ( .A(n246), .B(n10140), .Z(n10139) );
  XOR U9858 ( .A(p_input[2924]), .B(p_input[2892]), .Z(n10140) );
  XNOR U9859 ( .A(n9293), .B(n10135), .Z(n10137) );
  XOR U9860 ( .A(n10141), .B(n10142), .Z(n9293) );
  AND U9861 ( .A(n243), .B(n10143), .Z(n10142) );
  XOR U9862 ( .A(p_input[2860]), .B(p_input[2828]), .Z(n10143) );
  XOR U9863 ( .A(n10144), .B(n10145), .Z(n10135) );
  AND U9864 ( .A(n10146), .B(n10147), .Z(n10145) );
  XOR U9865 ( .A(n10144), .B(n9308), .Z(n10147) );
  XNOR U9866 ( .A(p_input[2891]), .B(n10148), .Z(n9308) );
  AND U9867 ( .A(n246), .B(n10149), .Z(n10148) );
  XOR U9868 ( .A(p_input[2923]), .B(p_input[2891]), .Z(n10149) );
  XNOR U9869 ( .A(n9305), .B(n10144), .Z(n10146) );
  XOR U9870 ( .A(n10150), .B(n10151), .Z(n9305) );
  AND U9871 ( .A(n243), .B(n10152), .Z(n10151) );
  XOR U9872 ( .A(p_input[2859]), .B(p_input[2827]), .Z(n10152) );
  XOR U9873 ( .A(n10153), .B(n10154), .Z(n10144) );
  AND U9874 ( .A(n10155), .B(n10156), .Z(n10154) );
  XOR U9875 ( .A(n10153), .B(n9320), .Z(n10156) );
  XNOR U9876 ( .A(p_input[2890]), .B(n10157), .Z(n9320) );
  AND U9877 ( .A(n246), .B(n10158), .Z(n10157) );
  XOR U9878 ( .A(p_input[2922]), .B(p_input[2890]), .Z(n10158) );
  XNOR U9879 ( .A(n9317), .B(n10153), .Z(n10155) );
  XOR U9880 ( .A(n10159), .B(n10160), .Z(n9317) );
  AND U9881 ( .A(n243), .B(n10161), .Z(n10160) );
  XOR U9882 ( .A(p_input[2858]), .B(p_input[2826]), .Z(n10161) );
  XOR U9883 ( .A(n10162), .B(n10163), .Z(n10153) );
  AND U9884 ( .A(n10164), .B(n10165), .Z(n10163) );
  XOR U9885 ( .A(n10162), .B(n9332), .Z(n10165) );
  XNOR U9886 ( .A(p_input[2889]), .B(n10166), .Z(n9332) );
  AND U9887 ( .A(n246), .B(n10167), .Z(n10166) );
  XOR U9888 ( .A(p_input[2921]), .B(p_input[2889]), .Z(n10167) );
  XNOR U9889 ( .A(n9329), .B(n10162), .Z(n10164) );
  XOR U9890 ( .A(n10168), .B(n10169), .Z(n9329) );
  AND U9891 ( .A(n243), .B(n10170), .Z(n10169) );
  XOR U9892 ( .A(p_input[2857]), .B(p_input[2825]), .Z(n10170) );
  XOR U9893 ( .A(n10171), .B(n10172), .Z(n10162) );
  AND U9894 ( .A(n10173), .B(n10174), .Z(n10172) );
  XOR U9895 ( .A(n10171), .B(n9344), .Z(n10174) );
  XNOR U9896 ( .A(p_input[2888]), .B(n10175), .Z(n9344) );
  AND U9897 ( .A(n246), .B(n10176), .Z(n10175) );
  XOR U9898 ( .A(p_input[2920]), .B(p_input[2888]), .Z(n10176) );
  XNOR U9899 ( .A(n9341), .B(n10171), .Z(n10173) );
  XOR U9900 ( .A(n10177), .B(n10178), .Z(n9341) );
  AND U9901 ( .A(n243), .B(n10179), .Z(n10178) );
  XOR U9902 ( .A(p_input[2856]), .B(p_input[2824]), .Z(n10179) );
  XOR U9903 ( .A(n10180), .B(n10181), .Z(n10171) );
  AND U9904 ( .A(n10182), .B(n10183), .Z(n10181) );
  XOR U9905 ( .A(n10180), .B(n9356), .Z(n10183) );
  XNOR U9906 ( .A(p_input[2887]), .B(n10184), .Z(n9356) );
  AND U9907 ( .A(n246), .B(n10185), .Z(n10184) );
  XOR U9908 ( .A(p_input[2919]), .B(p_input[2887]), .Z(n10185) );
  XNOR U9909 ( .A(n9353), .B(n10180), .Z(n10182) );
  XOR U9910 ( .A(n10186), .B(n10187), .Z(n9353) );
  AND U9911 ( .A(n243), .B(n10188), .Z(n10187) );
  XOR U9912 ( .A(p_input[2855]), .B(p_input[2823]), .Z(n10188) );
  XOR U9913 ( .A(n10189), .B(n10190), .Z(n10180) );
  AND U9914 ( .A(n10191), .B(n10192), .Z(n10190) );
  XOR U9915 ( .A(n10189), .B(n9368), .Z(n10192) );
  XNOR U9916 ( .A(p_input[2886]), .B(n10193), .Z(n9368) );
  AND U9917 ( .A(n246), .B(n10194), .Z(n10193) );
  XOR U9918 ( .A(p_input[2918]), .B(p_input[2886]), .Z(n10194) );
  XNOR U9919 ( .A(n9365), .B(n10189), .Z(n10191) );
  XOR U9920 ( .A(n10195), .B(n10196), .Z(n9365) );
  AND U9921 ( .A(n243), .B(n10197), .Z(n10196) );
  XOR U9922 ( .A(p_input[2854]), .B(p_input[2822]), .Z(n10197) );
  XOR U9923 ( .A(n10198), .B(n10199), .Z(n10189) );
  AND U9924 ( .A(n10200), .B(n10201), .Z(n10199) );
  XOR U9925 ( .A(n10198), .B(n9380), .Z(n10201) );
  XNOR U9926 ( .A(p_input[2885]), .B(n10202), .Z(n9380) );
  AND U9927 ( .A(n246), .B(n10203), .Z(n10202) );
  XOR U9928 ( .A(p_input[2917]), .B(p_input[2885]), .Z(n10203) );
  XNOR U9929 ( .A(n9377), .B(n10198), .Z(n10200) );
  XOR U9930 ( .A(n10204), .B(n10205), .Z(n9377) );
  AND U9931 ( .A(n243), .B(n10206), .Z(n10205) );
  XOR U9932 ( .A(p_input[2853]), .B(p_input[2821]), .Z(n10206) );
  XOR U9933 ( .A(n10207), .B(n10208), .Z(n10198) );
  AND U9934 ( .A(n10209), .B(n10210), .Z(n10208) );
  XOR U9935 ( .A(n10207), .B(n9392), .Z(n10210) );
  XNOR U9936 ( .A(p_input[2884]), .B(n10211), .Z(n9392) );
  AND U9937 ( .A(n246), .B(n10212), .Z(n10211) );
  XOR U9938 ( .A(p_input[2916]), .B(p_input[2884]), .Z(n10212) );
  XNOR U9939 ( .A(n9389), .B(n10207), .Z(n10209) );
  XOR U9940 ( .A(n10213), .B(n10214), .Z(n9389) );
  AND U9941 ( .A(n243), .B(n10215), .Z(n10214) );
  XOR U9942 ( .A(p_input[2852]), .B(p_input[2820]), .Z(n10215) );
  XOR U9943 ( .A(n10216), .B(n10217), .Z(n10207) );
  AND U9944 ( .A(n10218), .B(n10219), .Z(n10217) );
  XOR U9945 ( .A(n10216), .B(n9404), .Z(n10219) );
  XNOR U9946 ( .A(p_input[2883]), .B(n10220), .Z(n9404) );
  AND U9947 ( .A(n246), .B(n10221), .Z(n10220) );
  XOR U9948 ( .A(p_input[2915]), .B(p_input[2883]), .Z(n10221) );
  XNOR U9949 ( .A(n9401), .B(n10216), .Z(n10218) );
  XOR U9950 ( .A(n10222), .B(n10223), .Z(n9401) );
  AND U9951 ( .A(n243), .B(n10224), .Z(n10223) );
  XOR U9952 ( .A(p_input[2851]), .B(p_input[2819]), .Z(n10224) );
  XOR U9953 ( .A(n10225), .B(n10226), .Z(n10216) );
  AND U9954 ( .A(n10227), .B(n10228), .Z(n10226) );
  XOR U9955 ( .A(n9416), .B(n10225), .Z(n10228) );
  XNOR U9956 ( .A(p_input[2882]), .B(n10229), .Z(n9416) );
  AND U9957 ( .A(n246), .B(n10230), .Z(n10229) );
  XOR U9958 ( .A(p_input[2914]), .B(p_input[2882]), .Z(n10230) );
  XNOR U9959 ( .A(n10225), .B(n9413), .Z(n10227) );
  XOR U9960 ( .A(n10231), .B(n10232), .Z(n9413) );
  AND U9961 ( .A(n243), .B(n10233), .Z(n10232) );
  XOR U9962 ( .A(p_input[2850]), .B(p_input[2818]), .Z(n10233) );
  XOR U9963 ( .A(n10234), .B(n10235), .Z(n10225) );
  AND U9964 ( .A(n10236), .B(n10237), .Z(n10235) );
  XNOR U9965 ( .A(n10238), .B(n9429), .Z(n10237) );
  XNOR U9966 ( .A(p_input[2881]), .B(n10239), .Z(n9429) );
  AND U9967 ( .A(n246), .B(n10240), .Z(n10239) );
  XNOR U9968 ( .A(p_input[2913]), .B(n10241), .Z(n10240) );
  IV U9969 ( .A(p_input[2881]), .Z(n10241) );
  XNOR U9970 ( .A(n9426), .B(n10234), .Z(n10236) );
  XNOR U9971 ( .A(p_input[2817]), .B(n10242), .Z(n9426) );
  AND U9972 ( .A(n243), .B(n10243), .Z(n10242) );
  XOR U9973 ( .A(p_input[2849]), .B(p_input[2817]), .Z(n10243) );
  IV U9974 ( .A(n10238), .Z(n10234) );
  AND U9975 ( .A(n9964), .B(n9967), .Z(n10238) );
  XOR U9976 ( .A(p_input[2880]), .B(n10244), .Z(n9967) );
  AND U9977 ( .A(n246), .B(n10245), .Z(n10244) );
  XOR U9978 ( .A(p_input[2912]), .B(p_input[2880]), .Z(n10245) );
  XOR U9979 ( .A(n10246), .B(n10247), .Z(n246) );
  AND U9980 ( .A(n10248), .B(n10249), .Z(n10247) );
  XNOR U9981 ( .A(p_input[2943]), .B(n10246), .Z(n10249) );
  XOR U9982 ( .A(n10246), .B(p_input[2911]), .Z(n10248) );
  XOR U9983 ( .A(n10250), .B(n10251), .Z(n10246) );
  AND U9984 ( .A(n10252), .B(n10253), .Z(n10251) );
  XNOR U9985 ( .A(p_input[2942]), .B(n10250), .Z(n10253) );
  XOR U9986 ( .A(n10250), .B(p_input[2910]), .Z(n10252) );
  XOR U9987 ( .A(n10254), .B(n10255), .Z(n10250) );
  AND U9988 ( .A(n10256), .B(n10257), .Z(n10255) );
  XNOR U9989 ( .A(p_input[2941]), .B(n10254), .Z(n10257) );
  XOR U9990 ( .A(n10254), .B(p_input[2909]), .Z(n10256) );
  XOR U9991 ( .A(n10258), .B(n10259), .Z(n10254) );
  AND U9992 ( .A(n10260), .B(n10261), .Z(n10259) );
  XNOR U9993 ( .A(p_input[2940]), .B(n10258), .Z(n10261) );
  XOR U9994 ( .A(n10258), .B(p_input[2908]), .Z(n10260) );
  XOR U9995 ( .A(n10262), .B(n10263), .Z(n10258) );
  AND U9996 ( .A(n10264), .B(n10265), .Z(n10263) );
  XNOR U9997 ( .A(p_input[2939]), .B(n10262), .Z(n10265) );
  XOR U9998 ( .A(n10262), .B(p_input[2907]), .Z(n10264) );
  XOR U9999 ( .A(n10266), .B(n10267), .Z(n10262) );
  AND U10000 ( .A(n10268), .B(n10269), .Z(n10267) );
  XNOR U10001 ( .A(p_input[2938]), .B(n10266), .Z(n10269) );
  XOR U10002 ( .A(n10266), .B(p_input[2906]), .Z(n10268) );
  XOR U10003 ( .A(n10270), .B(n10271), .Z(n10266) );
  AND U10004 ( .A(n10272), .B(n10273), .Z(n10271) );
  XNOR U10005 ( .A(p_input[2937]), .B(n10270), .Z(n10273) );
  XOR U10006 ( .A(n10270), .B(p_input[2905]), .Z(n10272) );
  XOR U10007 ( .A(n10274), .B(n10275), .Z(n10270) );
  AND U10008 ( .A(n10276), .B(n10277), .Z(n10275) );
  XNOR U10009 ( .A(p_input[2936]), .B(n10274), .Z(n10277) );
  XOR U10010 ( .A(n10274), .B(p_input[2904]), .Z(n10276) );
  XOR U10011 ( .A(n10278), .B(n10279), .Z(n10274) );
  AND U10012 ( .A(n10280), .B(n10281), .Z(n10279) );
  XNOR U10013 ( .A(p_input[2935]), .B(n10278), .Z(n10281) );
  XOR U10014 ( .A(n10278), .B(p_input[2903]), .Z(n10280) );
  XOR U10015 ( .A(n10282), .B(n10283), .Z(n10278) );
  AND U10016 ( .A(n10284), .B(n10285), .Z(n10283) );
  XNOR U10017 ( .A(p_input[2934]), .B(n10282), .Z(n10285) );
  XOR U10018 ( .A(n10282), .B(p_input[2902]), .Z(n10284) );
  XOR U10019 ( .A(n10286), .B(n10287), .Z(n10282) );
  AND U10020 ( .A(n10288), .B(n10289), .Z(n10287) );
  XNOR U10021 ( .A(p_input[2933]), .B(n10286), .Z(n10289) );
  XOR U10022 ( .A(n10286), .B(p_input[2901]), .Z(n10288) );
  XOR U10023 ( .A(n10290), .B(n10291), .Z(n10286) );
  AND U10024 ( .A(n10292), .B(n10293), .Z(n10291) );
  XNOR U10025 ( .A(p_input[2932]), .B(n10290), .Z(n10293) );
  XOR U10026 ( .A(n10290), .B(p_input[2900]), .Z(n10292) );
  XOR U10027 ( .A(n10294), .B(n10295), .Z(n10290) );
  AND U10028 ( .A(n10296), .B(n10297), .Z(n10295) );
  XNOR U10029 ( .A(p_input[2931]), .B(n10294), .Z(n10297) );
  XOR U10030 ( .A(n10294), .B(p_input[2899]), .Z(n10296) );
  XOR U10031 ( .A(n10298), .B(n10299), .Z(n10294) );
  AND U10032 ( .A(n10300), .B(n10301), .Z(n10299) );
  XNOR U10033 ( .A(p_input[2930]), .B(n10298), .Z(n10301) );
  XOR U10034 ( .A(n10298), .B(p_input[2898]), .Z(n10300) );
  XOR U10035 ( .A(n10302), .B(n10303), .Z(n10298) );
  AND U10036 ( .A(n10304), .B(n10305), .Z(n10303) );
  XNOR U10037 ( .A(p_input[2929]), .B(n10302), .Z(n10305) );
  XOR U10038 ( .A(n10302), .B(p_input[2897]), .Z(n10304) );
  XOR U10039 ( .A(n10306), .B(n10307), .Z(n10302) );
  AND U10040 ( .A(n10308), .B(n10309), .Z(n10307) );
  XNOR U10041 ( .A(p_input[2928]), .B(n10306), .Z(n10309) );
  XOR U10042 ( .A(n10306), .B(p_input[2896]), .Z(n10308) );
  XOR U10043 ( .A(n10310), .B(n10311), .Z(n10306) );
  AND U10044 ( .A(n10312), .B(n10313), .Z(n10311) );
  XNOR U10045 ( .A(p_input[2927]), .B(n10310), .Z(n10313) );
  XOR U10046 ( .A(n10310), .B(p_input[2895]), .Z(n10312) );
  XOR U10047 ( .A(n10314), .B(n10315), .Z(n10310) );
  AND U10048 ( .A(n10316), .B(n10317), .Z(n10315) );
  XNOR U10049 ( .A(p_input[2926]), .B(n10314), .Z(n10317) );
  XOR U10050 ( .A(n10314), .B(p_input[2894]), .Z(n10316) );
  XOR U10051 ( .A(n10318), .B(n10319), .Z(n10314) );
  AND U10052 ( .A(n10320), .B(n10321), .Z(n10319) );
  XNOR U10053 ( .A(p_input[2925]), .B(n10318), .Z(n10321) );
  XOR U10054 ( .A(n10318), .B(p_input[2893]), .Z(n10320) );
  XOR U10055 ( .A(n10322), .B(n10323), .Z(n10318) );
  AND U10056 ( .A(n10324), .B(n10325), .Z(n10323) );
  XNOR U10057 ( .A(p_input[2924]), .B(n10322), .Z(n10325) );
  XOR U10058 ( .A(n10322), .B(p_input[2892]), .Z(n10324) );
  XOR U10059 ( .A(n10326), .B(n10327), .Z(n10322) );
  AND U10060 ( .A(n10328), .B(n10329), .Z(n10327) );
  XNOR U10061 ( .A(p_input[2923]), .B(n10326), .Z(n10329) );
  XOR U10062 ( .A(n10326), .B(p_input[2891]), .Z(n10328) );
  XOR U10063 ( .A(n10330), .B(n10331), .Z(n10326) );
  AND U10064 ( .A(n10332), .B(n10333), .Z(n10331) );
  XNOR U10065 ( .A(p_input[2922]), .B(n10330), .Z(n10333) );
  XOR U10066 ( .A(n10330), .B(p_input[2890]), .Z(n10332) );
  XOR U10067 ( .A(n10334), .B(n10335), .Z(n10330) );
  AND U10068 ( .A(n10336), .B(n10337), .Z(n10335) );
  XNOR U10069 ( .A(p_input[2921]), .B(n10334), .Z(n10337) );
  XOR U10070 ( .A(n10334), .B(p_input[2889]), .Z(n10336) );
  XOR U10071 ( .A(n10338), .B(n10339), .Z(n10334) );
  AND U10072 ( .A(n10340), .B(n10341), .Z(n10339) );
  XNOR U10073 ( .A(p_input[2920]), .B(n10338), .Z(n10341) );
  XOR U10074 ( .A(n10338), .B(p_input[2888]), .Z(n10340) );
  XOR U10075 ( .A(n10342), .B(n10343), .Z(n10338) );
  AND U10076 ( .A(n10344), .B(n10345), .Z(n10343) );
  XNOR U10077 ( .A(p_input[2919]), .B(n10342), .Z(n10345) );
  XOR U10078 ( .A(n10342), .B(p_input[2887]), .Z(n10344) );
  XOR U10079 ( .A(n10346), .B(n10347), .Z(n10342) );
  AND U10080 ( .A(n10348), .B(n10349), .Z(n10347) );
  XNOR U10081 ( .A(p_input[2918]), .B(n10346), .Z(n10349) );
  XOR U10082 ( .A(n10346), .B(p_input[2886]), .Z(n10348) );
  XOR U10083 ( .A(n10350), .B(n10351), .Z(n10346) );
  AND U10084 ( .A(n10352), .B(n10353), .Z(n10351) );
  XNOR U10085 ( .A(p_input[2917]), .B(n10350), .Z(n10353) );
  XOR U10086 ( .A(n10350), .B(p_input[2885]), .Z(n10352) );
  XOR U10087 ( .A(n10354), .B(n10355), .Z(n10350) );
  AND U10088 ( .A(n10356), .B(n10357), .Z(n10355) );
  XNOR U10089 ( .A(p_input[2916]), .B(n10354), .Z(n10357) );
  XOR U10090 ( .A(n10354), .B(p_input[2884]), .Z(n10356) );
  XOR U10091 ( .A(n10358), .B(n10359), .Z(n10354) );
  AND U10092 ( .A(n10360), .B(n10361), .Z(n10359) );
  XNOR U10093 ( .A(p_input[2915]), .B(n10358), .Z(n10361) );
  XOR U10094 ( .A(n10358), .B(p_input[2883]), .Z(n10360) );
  XOR U10095 ( .A(n10362), .B(n10363), .Z(n10358) );
  AND U10096 ( .A(n10364), .B(n10365), .Z(n10363) );
  XNOR U10097 ( .A(p_input[2914]), .B(n10362), .Z(n10365) );
  XOR U10098 ( .A(n10362), .B(p_input[2882]), .Z(n10364) );
  XNOR U10099 ( .A(n10366), .B(n10367), .Z(n10362) );
  AND U10100 ( .A(n10368), .B(n10369), .Z(n10367) );
  XOR U10101 ( .A(p_input[2913]), .B(n10366), .Z(n10369) );
  XNOR U10102 ( .A(p_input[2881]), .B(n10366), .Z(n10368) );
  AND U10103 ( .A(p_input[2912]), .B(n10370), .Z(n10366) );
  IV U10104 ( .A(p_input[2880]), .Z(n10370) );
  XNOR U10105 ( .A(p_input[2816]), .B(n10371), .Z(n9964) );
  AND U10106 ( .A(n243), .B(n10372), .Z(n10371) );
  XOR U10107 ( .A(p_input[2848]), .B(p_input[2816]), .Z(n10372) );
  XOR U10108 ( .A(n10373), .B(n10374), .Z(n243) );
  AND U10109 ( .A(n10375), .B(n10376), .Z(n10374) );
  XNOR U10110 ( .A(p_input[2879]), .B(n10373), .Z(n10376) );
  XOR U10111 ( .A(n10373), .B(p_input[2847]), .Z(n10375) );
  XOR U10112 ( .A(n10377), .B(n10378), .Z(n10373) );
  AND U10113 ( .A(n10379), .B(n10380), .Z(n10378) );
  XNOR U10114 ( .A(p_input[2878]), .B(n10377), .Z(n10380) );
  XNOR U10115 ( .A(n10377), .B(n9979), .Z(n10379) );
  IV U10116 ( .A(p_input[2846]), .Z(n9979) );
  XOR U10117 ( .A(n10381), .B(n10382), .Z(n10377) );
  AND U10118 ( .A(n10383), .B(n10384), .Z(n10382) );
  XNOR U10119 ( .A(p_input[2877]), .B(n10381), .Z(n10384) );
  XNOR U10120 ( .A(n10381), .B(n9988), .Z(n10383) );
  IV U10121 ( .A(p_input[2845]), .Z(n9988) );
  XOR U10122 ( .A(n10385), .B(n10386), .Z(n10381) );
  AND U10123 ( .A(n10387), .B(n10388), .Z(n10386) );
  XNOR U10124 ( .A(p_input[2876]), .B(n10385), .Z(n10388) );
  XNOR U10125 ( .A(n10385), .B(n9997), .Z(n10387) );
  IV U10126 ( .A(p_input[2844]), .Z(n9997) );
  XOR U10127 ( .A(n10389), .B(n10390), .Z(n10385) );
  AND U10128 ( .A(n10391), .B(n10392), .Z(n10390) );
  XNOR U10129 ( .A(p_input[2875]), .B(n10389), .Z(n10392) );
  XNOR U10130 ( .A(n10389), .B(n10006), .Z(n10391) );
  IV U10131 ( .A(p_input[2843]), .Z(n10006) );
  XOR U10132 ( .A(n10393), .B(n10394), .Z(n10389) );
  AND U10133 ( .A(n10395), .B(n10396), .Z(n10394) );
  XNOR U10134 ( .A(p_input[2874]), .B(n10393), .Z(n10396) );
  XNOR U10135 ( .A(n10393), .B(n10015), .Z(n10395) );
  IV U10136 ( .A(p_input[2842]), .Z(n10015) );
  XOR U10137 ( .A(n10397), .B(n10398), .Z(n10393) );
  AND U10138 ( .A(n10399), .B(n10400), .Z(n10398) );
  XNOR U10139 ( .A(p_input[2873]), .B(n10397), .Z(n10400) );
  XNOR U10140 ( .A(n10397), .B(n10024), .Z(n10399) );
  IV U10141 ( .A(p_input[2841]), .Z(n10024) );
  XOR U10142 ( .A(n10401), .B(n10402), .Z(n10397) );
  AND U10143 ( .A(n10403), .B(n10404), .Z(n10402) );
  XNOR U10144 ( .A(p_input[2872]), .B(n10401), .Z(n10404) );
  XNOR U10145 ( .A(n10401), .B(n10033), .Z(n10403) );
  IV U10146 ( .A(p_input[2840]), .Z(n10033) );
  XOR U10147 ( .A(n10405), .B(n10406), .Z(n10401) );
  AND U10148 ( .A(n10407), .B(n10408), .Z(n10406) );
  XNOR U10149 ( .A(p_input[2871]), .B(n10405), .Z(n10408) );
  XNOR U10150 ( .A(n10405), .B(n10042), .Z(n10407) );
  IV U10151 ( .A(p_input[2839]), .Z(n10042) );
  XOR U10152 ( .A(n10409), .B(n10410), .Z(n10405) );
  AND U10153 ( .A(n10411), .B(n10412), .Z(n10410) );
  XNOR U10154 ( .A(p_input[2870]), .B(n10409), .Z(n10412) );
  XNOR U10155 ( .A(n10409), .B(n10051), .Z(n10411) );
  IV U10156 ( .A(p_input[2838]), .Z(n10051) );
  XOR U10157 ( .A(n10413), .B(n10414), .Z(n10409) );
  AND U10158 ( .A(n10415), .B(n10416), .Z(n10414) );
  XNOR U10159 ( .A(p_input[2869]), .B(n10413), .Z(n10416) );
  XNOR U10160 ( .A(n10413), .B(n10060), .Z(n10415) );
  IV U10161 ( .A(p_input[2837]), .Z(n10060) );
  XOR U10162 ( .A(n10417), .B(n10418), .Z(n10413) );
  AND U10163 ( .A(n10419), .B(n10420), .Z(n10418) );
  XNOR U10164 ( .A(p_input[2868]), .B(n10417), .Z(n10420) );
  XNOR U10165 ( .A(n10417), .B(n10069), .Z(n10419) );
  IV U10166 ( .A(p_input[2836]), .Z(n10069) );
  XOR U10167 ( .A(n10421), .B(n10422), .Z(n10417) );
  AND U10168 ( .A(n10423), .B(n10424), .Z(n10422) );
  XNOR U10169 ( .A(p_input[2867]), .B(n10421), .Z(n10424) );
  XNOR U10170 ( .A(n10421), .B(n10078), .Z(n10423) );
  IV U10171 ( .A(p_input[2835]), .Z(n10078) );
  XOR U10172 ( .A(n10425), .B(n10426), .Z(n10421) );
  AND U10173 ( .A(n10427), .B(n10428), .Z(n10426) );
  XNOR U10174 ( .A(p_input[2866]), .B(n10425), .Z(n10428) );
  XNOR U10175 ( .A(n10425), .B(n10087), .Z(n10427) );
  IV U10176 ( .A(p_input[2834]), .Z(n10087) );
  XOR U10177 ( .A(n10429), .B(n10430), .Z(n10425) );
  AND U10178 ( .A(n10431), .B(n10432), .Z(n10430) );
  XNOR U10179 ( .A(p_input[2865]), .B(n10429), .Z(n10432) );
  XNOR U10180 ( .A(n10429), .B(n10096), .Z(n10431) );
  IV U10181 ( .A(p_input[2833]), .Z(n10096) );
  XOR U10182 ( .A(n10433), .B(n10434), .Z(n10429) );
  AND U10183 ( .A(n10435), .B(n10436), .Z(n10434) );
  XNOR U10184 ( .A(p_input[2864]), .B(n10433), .Z(n10436) );
  XNOR U10185 ( .A(n10433), .B(n10105), .Z(n10435) );
  IV U10186 ( .A(p_input[2832]), .Z(n10105) );
  XOR U10187 ( .A(n10437), .B(n10438), .Z(n10433) );
  AND U10188 ( .A(n10439), .B(n10440), .Z(n10438) );
  XNOR U10189 ( .A(p_input[2863]), .B(n10437), .Z(n10440) );
  XNOR U10190 ( .A(n10437), .B(n10114), .Z(n10439) );
  IV U10191 ( .A(p_input[2831]), .Z(n10114) );
  XOR U10192 ( .A(n10441), .B(n10442), .Z(n10437) );
  AND U10193 ( .A(n10443), .B(n10444), .Z(n10442) );
  XNOR U10194 ( .A(p_input[2862]), .B(n10441), .Z(n10444) );
  XNOR U10195 ( .A(n10441), .B(n10123), .Z(n10443) );
  IV U10196 ( .A(p_input[2830]), .Z(n10123) );
  XOR U10197 ( .A(n10445), .B(n10446), .Z(n10441) );
  AND U10198 ( .A(n10447), .B(n10448), .Z(n10446) );
  XNOR U10199 ( .A(p_input[2861]), .B(n10445), .Z(n10448) );
  XNOR U10200 ( .A(n10445), .B(n10132), .Z(n10447) );
  IV U10201 ( .A(p_input[2829]), .Z(n10132) );
  XOR U10202 ( .A(n10449), .B(n10450), .Z(n10445) );
  AND U10203 ( .A(n10451), .B(n10452), .Z(n10450) );
  XNOR U10204 ( .A(p_input[2860]), .B(n10449), .Z(n10452) );
  XNOR U10205 ( .A(n10449), .B(n10141), .Z(n10451) );
  IV U10206 ( .A(p_input[2828]), .Z(n10141) );
  XOR U10207 ( .A(n10453), .B(n10454), .Z(n10449) );
  AND U10208 ( .A(n10455), .B(n10456), .Z(n10454) );
  XNOR U10209 ( .A(p_input[2859]), .B(n10453), .Z(n10456) );
  XNOR U10210 ( .A(n10453), .B(n10150), .Z(n10455) );
  IV U10211 ( .A(p_input[2827]), .Z(n10150) );
  XOR U10212 ( .A(n10457), .B(n10458), .Z(n10453) );
  AND U10213 ( .A(n10459), .B(n10460), .Z(n10458) );
  XNOR U10214 ( .A(p_input[2858]), .B(n10457), .Z(n10460) );
  XNOR U10215 ( .A(n10457), .B(n10159), .Z(n10459) );
  IV U10216 ( .A(p_input[2826]), .Z(n10159) );
  XOR U10217 ( .A(n10461), .B(n10462), .Z(n10457) );
  AND U10218 ( .A(n10463), .B(n10464), .Z(n10462) );
  XNOR U10219 ( .A(p_input[2857]), .B(n10461), .Z(n10464) );
  XNOR U10220 ( .A(n10461), .B(n10168), .Z(n10463) );
  IV U10221 ( .A(p_input[2825]), .Z(n10168) );
  XOR U10222 ( .A(n10465), .B(n10466), .Z(n10461) );
  AND U10223 ( .A(n10467), .B(n10468), .Z(n10466) );
  XNOR U10224 ( .A(p_input[2856]), .B(n10465), .Z(n10468) );
  XNOR U10225 ( .A(n10465), .B(n10177), .Z(n10467) );
  IV U10226 ( .A(p_input[2824]), .Z(n10177) );
  XOR U10227 ( .A(n10469), .B(n10470), .Z(n10465) );
  AND U10228 ( .A(n10471), .B(n10472), .Z(n10470) );
  XNOR U10229 ( .A(p_input[2855]), .B(n10469), .Z(n10472) );
  XNOR U10230 ( .A(n10469), .B(n10186), .Z(n10471) );
  IV U10231 ( .A(p_input[2823]), .Z(n10186) );
  XOR U10232 ( .A(n10473), .B(n10474), .Z(n10469) );
  AND U10233 ( .A(n10475), .B(n10476), .Z(n10474) );
  XNOR U10234 ( .A(p_input[2854]), .B(n10473), .Z(n10476) );
  XNOR U10235 ( .A(n10473), .B(n10195), .Z(n10475) );
  IV U10236 ( .A(p_input[2822]), .Z(n10195) );
  XOR U10237 ( .A(n10477), .B(n10478), .Z(n10473) );
  AND U10238 ( .A(n10479), .B(n10480), .Z(n10478) );
  XNOR U10239 ( .A(p_input[2853]), .B(n10477), .Z(n10480) );
  XNOR U10240 ( .A(n10477), .B(n10204), .Z(n10479) );
  IV U10241 ( .A(p_input[2821]), .Z(n10204) );
  XOR U10242 ( .A(n10481), .B(n10482), .Z(n10477) );
  AND U10243 ( .A(n10483), .B(n10484), .Z(n10482) );
  XNOR U10244 ( .A(p_input[2852]), .B(n10481), .Z(n10484) );
  XNOR U10245 ( .A(n10481), .B(n10213), .Z(n10483) );
  IV U10246 ( .A(p_input[2820]), .Z(n10213) );
  XOR U10247 ( .A(n10485), .B(n10486), .Z(n10481) );
  AND U10248 ( .A(n10487), .B(n10488), .Z(n10486) );
  XNOR U10249 ( .A(p_input[2851]), .B(n10485), .Z(n10488) );
  XNOR U10250 ( .A(n10485), .B(n10222), .Z(n10487) );
  IV U10251 ( .A(p_input[2819]), .Z(n10222) );
  XOR U10252 ( .A(n10489), .B(n10490), .Z(n10485) );
  AND U10253 ( .A(n10491), .B(n10492), .Z(n10490) );
  XNOR U10254 ( .A(p_input[2850]), .B(n10489), .Z(n10492) );
  XNOR U10255 ( .A(n10489), .B(n10231), .Z(n10491) );
  IV U10256 ( .A(p_input[2818]), .Z(n10231) );
  XNOR U10257 ( .A(n10493), .B(n10494), .Z(n10489) );
  AND U10258 ( .A(n10495), .B(n10496), .Z(n10494) );
  XOR U10259 ( .A(p_input[2849]), .B(n10493), .Z(n10496) );
  XNOR U10260 ( .A(p_input[2817]), .B(n10493), .Z(n10495) );
  AND U10261 ( .A(p_input[2848]), .B(n10497), .Z(n10493) );
  IV U10262 ( .A(p_input[2816]), .Z(n10497) );
  XOR U10263 ( .A(n10498), .B(n10499), .Z(n8676) );
  AND U10264 ( .A(n500), .B(n10500), .Z(n10499) );
  XNOR U10265 ( .A(n10501), .B(n10498), .Z(n10500) );
  XOR U10266 ( .A(n10502), .B(n10503), .Z(n500) );
  AND U10267 ( .A(n10504), .B(n10505), .Z(n10503) );
  XOR U10268 ( .A(n10502), .B(n8691), .Z(n10505) );
  XNOR U10269 ( .A(n10506), .B(n10507), .Z(n8691) );
  AND U10270 ( .A(n10508), .B(n338), .Z(n10507) );
  AND U10271 ( .A(n10506), .B(n10509), .Z(n10508) );
  XNOR U10272 ( .A(n8688), .B(n10502), .Z(n10504) );
  XOR U10273 ( .A(n10510), .B(n10511), .Z(n8688) );
  AND U10274 ( .A(n10512), .B(n335), .Z(n10511) );
  NOR U10275 ( .A(n10510), .B(n10513), .Z(n10512) );
  XOR U10276 ( .A(n10514), .B(n10515), .Z(n10502) );
  AND U10277 ( .A(n10516), .B(n10517), .Z(n10515) );
  XOR U10278 ( .A(n10514), .B(n8703), .Z(n10517) );
  XOR U10279 ( .A(n10518), .B(n10519), .Z(n8703) );
  AND U10280 ( .A(n338), .B(n10520), .Z(n10519) );
  XOR U10281 ( .A(n10521), .B(n10518), .Z(n10520) );
  XNOR U10282 ( .A(n8700), .B(n10514), .Z(n10516) );
  XOR U10283 ( .A(n10522), .B(n10523), .Z(n8700) );
  AND U10284 ( .A(n335), .B(n10524), .Z(n10523) );
  XOR U10285 ( .A(n10525), .B(n10522), .Z(n10524) );
  XOR U10286 ( .A(n10526), .B(n10527), .Z(n10514) );
  AND U10287 ( .A(n10528), .B(n10529), .Z(n10527) );
  XOR U10288 ( .A(n10526), .B(n8715), .Z(n10529) );
  XOR U10289 ( .A(n10530), .B(n10531), .Z(n8715) );
  AND U10290 ( .A(n338), .B(n10532), .Z(n10531) );
  XOR U10291 ( .A(n10533), .B(n10530), .Z(n10532) );
  XNOR U10292 ( .A(n8712), .B(n10526), .Z(n10528) );
  XOR U10293 ( .A(n10534), .B(n10535), .Z(n8712) );
  AND U10294 ( .A(n335), .B(n10536), .Z(n10535) );
  XOR U10295 ( .A(n10537), .B(n10534), .Z(n10536) );
  XOR U10296 ( .A(n10538), .B(n10539), .Z(n10526) );
  AND U10297 ( .A(n10540), .B(n10541), .Z(n10539) );
  XOR U10298 ( .A(n10538), .B(n8727), .Z(n10541) );
  XOR U10299 ( .A(n10542), .B(n10543), .Z(n8727) );
  AND U10300 ( .A(n338), .B(n10544), .Z(n10543) );
  XOR U10301 ( .A(n10545), .B(n10542), .Z(n10544) );
  XNOR U10302 ( .A(n8724), .B(n10538), .Z(n10540) );
  XOR U10303 ( .A(n10546), .B(n10547), .Z(n8724) );
  AND U10304 ( .A(n335), .B(n10548), .Z(n10547) );
  XOR U10305 ( .A(n10549), .B(n10546), .Z(n10548) );
  XOR U10306 ( .A(n10550), .B(n10551), .Z(n10538) );
  AND U10307 ( .A(n10552), .B(n10553), .Z(n10551) );
  XOR U10308 ( .A(n10550), .B(n8739), .Z(n10553) );
  XOR U10309 ( .A(n10554), .B(n10555), .Z(n8739) );
  AND U10310 ( .A(n338), .B(n10556), .Z(n10555) );
  XOR U10311 ( .A(n10557), .B(n10554), .Z(n10556) );
  XNOR U10312 ( .A(n8736), .B(n10550), .Z(n10552) );
  XOR U10313 ( .A(n10558), .B(n10559), .Z(n8736) );
  AND U10314 ( .A(n335), .B(n10560), .Z(n10559) );
  XOR U10315 ( .A(n10561), .B(n10558), .Z(n10560) );
  XOR U10316 ( .A(n10562), .B(n10563), .Z(n10550) );
  AND U10317 ( .A(n10564), .B(n10565), .Z(n10563) );
  XOR U10318 ( .A(n10562), .B(n8751), .Z(n10565) );
  XOR U10319 ( .A(n10566), .B(n10567), .Z(n8751) );
  AND U10320 ( .A(n338), .B(n10568), .Z(n10567) );
  XOR U10321 ( .A(n10569), .B(n10566), .Z(n10568) );
  XNOR U10322 ( .A(n8748), .B(n10562), .Z(n10564) );
  XOR U10323 ( .A(n10570), .B(n10571), .Z(n8748) );
  AND U10324 ( .A(n335), .B(n10572), .Z(n10571) );
  XOR U10325 ( .A(n10573), .B(n10570), .Z(n10572) );
  XOR U10326 ( .A(n10574), .B(n10575), .Z(n10562) );
  AND U10327 ( .A(n10576), .B(n10577), .Z(n10575) );
  XOR U10328 ( .A(n10574), .B(n8763), .Z(n10577) );
  XOR U10329 ( .A(n10578), .B(n10579), .Z(n8763) );
  AND U10330 ( .A(n338), .B(n10580), .Z(n10579) );
  XOR U10331 ( .A(n10581), .B(n10578), .Z(n10580) );
  XNOR U10332 ( .A(n8760), .B(n10574), .Z(n10576) );
  XOR U10333 ( .A(n10582), .B(n10583), .Z(n8760) );
  AND U10334 ( .A(n335), .B(n10584), .Z(n10583) );
  XOR U10335 ( .A(n10585), .B(n10582), .Z(n10584) );
  XOR U10336 ( .A(n10586), .B(n10587), .Z(n10574) );
  AND U10337 ( .A(n10588), .B(n10589), .Z(n10587) );
  XOR U10338 ( .A(n10586), .B(n8775), .Z(n10589) );
  XOR U10339 ( .A(n10590), .B(n10591), .Z(n8775) );
  AND U10340 ( .A(n338), .B(n10592), .Z(n10591) );
  XOR U10341 ( .A(n10593), .B(n10590), .Z(n10592) );
  XNOR U10342 ( .A(n8772), .B(n10586), .Z(n10588) );
  XOR U10343 ( .A(n10594), .B(n10595), .Z(n8772) );
  AND U10344 ( .A(n335), .B(n10596), .Z(n10595) );
  XOR U10345 ( .A(n10597), .B(n10594), .Z(n10596) );
  XOR U10346 ( .A(n10598), .B(n10599), .Z(n10586) );
  AND U10347 ( .A(n10600), .B(n10601), .Z(n10599) );
  XOR U10348 ( .A(n10598), .B(n8787), .Z(n10601) );
  XOR U10349 ( .A(n10602), .B(n10603), .Z(n8787) );
  AND U10350 ( .A(n338), .B(n10604), .Z(n10603) );
  XOR U10351 ( .A(n10605), .B(n10602), .Z(n10604) );
  XNOR U10352 ( .A(n8784), .B(n10598), .Z(n10600) );
  XOR U10353 ( .A(n10606), .B(n10607), .Z(n8784) );
  AND U10354 ( .A(n335), .B(n10608), .Z(n10607) );
  XOR U10355 ( .A(n10609), .B(n10606), .Z(n10608) );
  XOR U10356 ( .A(n10610), .B(n10611), .Z(n10598) );
  AND U10357 ( .A(n10612), .B(n10613), .Z(n10611) );
  XOR U10358 ( .A(n10610), .B(n8799), .Z(n10613) );
  XOR U10359 ( .A(n10614), .B(n10615), .Z(n8799) );
  AND U10360 ( .A(n338), .B(n10616), .Z(n10615) );
  XOR U10361 ( .A(n10617), .B(n10614), .Z(n10616) );
  XNOR U10362 ( .A(n8796), .B(n10610), .Z(n10612) );
  XOR U10363 ( .A(n10618), .B(n10619), .Z(n8796) );
  AND U10364 ( .A(n335), .B(n10620), .Z(n10619) );
  XOR U10365 ( .A(n10621), .B(n10618), .Z(n10620) );
  XOR U10366 ( .A(n10622), .B(n10623), .Z(n10610) );
  AND U10367 ( .A(n10624), .B(n10625), .Z(n10623) );
  XOR U10368 ( .A(n10622), .B(n8811), .Z(n10625) );
  XOR U10369 ( .A(n10626), .B(n10627), .Z(n8811) );
  AND U10370 ( .A(n338), .B(n10628), .Z(n10627) );
  XOR U10371 ( .A(n10629), .B(n10626), .Z(n10628) );
  XNOR U10372 ( .A(n8808), .B(n10622), .Z(n10624) );
  XOR U10373 ( .A(n10630), .B(n10631), .Z(n8808) );
  AND U10374 ( .A(n335), .B(n10632), .Z(n10631) );
  XOR U10375 ( .A(n10633), .B(n10630), .Z(n10632) );
  XOR U10376 ( .A(n10634), .B(n10635), .Z(n10622) );
  AND U10377 ( .A(n10636), .B(n10637), .Z(n10635) );
  XOR U10378 ( .A(n10634), .B(n8823), .Z(n10637) );
  XOR U10379 ( .A(n10638), .B(n10639), .Z(n8823) );
  AND U10380 ( .A(n338), .B(n10640), .Z(n10639) );
  XOR U10381 ( .A(n10641), .B(n10638), .Z(n10640) );
  XNOR U10382 ( .A(n8820), .B(n10634), .Z(n10636) );
  XOR U10383 ( .A(n10642), .B(n10643), .Z(n8820) );
  AND U10384 ( .A(n335), .B(n10644), .Z(n10643) );
  XOR U10385 ( .A(n10645), .B(n10642), .Z(n10644) );
  XOR U10386 ( .A(n10646), .B(n10647), .Z(n10634) );
  AND U10387 ( .A(n10648), .B(n10649), .Z(n10647) );
  XOR U10388 ( .A(n10646), .B(n8835), .Z(n10649) );
  XOR U10389 ( .A(n10650), .B(n10651), .Z(n8835) );
  AND U10390 ( .A(n338), .B(n10652), .Z(n10651) );
  XOR U10391 ( .A(n10653), .B(n10650), .Z(n10652) );
  XNOR U10392 ( .A(n8832), .B(n10646), .Z(n10648) );
  XOR U10393 ( .A(n10654), .B(n10655), .Z(n8832) );
  AND U10394 ( .A(n335), .B(n10656), .Z(n10655) );
  XOR U10395 ( .A(n10657), .B(n10654), .Z(n10656) );
  XOR U10396 ( .A(n10658), .B(n10659), .Z(n10646) );
  AND U10397 ( .A(n10660), .B(n10661), .Z(n10659) );
  XOR U10398 ( .A(n10658), .B(n8847), .Z(n10661) );
  XOR U10399 ( .A(n10662), .B(n10663), .Z(n8847) );
  AND U10400 ( .A(n338), .B(n10664), .Z(n10663) );
  XOR U10401 ( .A(n10665), .B(n10662), .Z(n10664) );
  XNOR U10402 ( .A(n8844), .B(n10658), .Z(n10660) );
  XOR U10403 ( .A(n10666), .B(n10667), .Z(n8844) );
  AND U10404 ( .A(n335), .B(n10668), .Z(n10667) );
  XOR U10405 ( .A(n10669), .B(n10666), .Z(n10668) );
  XOR U10406 ( .A(n10670), .B(n10671), .Z(n10658) );
  AND U10407 ( .A(n10672), .B(n10673), .Z(n10671) );
  XOR U10408 ( .A(n10670), .B(n8859), .Z(n10673) );
  XOR U10409 ( .A(n10674), .B(n10675), .Z(n8859) );
  AND U10410 ( .A(n338), .B(n10676), .Z(n10675) );
  XOR U10411 ( .A(n10677), .B(n10674), .Z(n10676) );
  XNOR U10412 ( .A(n8856), .B(n10670), .Z(n10672) );
  XOR U10413 ( .A(n10678), .B(n10679), .Z(n8856) );
  AND U10414 ( .A(n335), .B(n10680), .Z(n10679) );
  XOR U10415 ( .A(n10681), .B(n10678), .Z(n10680) );
  XOR U10416 ( .A(n10682), .B(n10683), .Z(n10670) );
  AND U10417 ( .A(n10684), .B(n10685), .Z(n10683) );
  XOR U10418 ( .A(n10682), .B(n8871), .Z(n10685) );
  XOR U10419 ( .A(n10686), .B(n10687), .Z(n8871) );
  AND U10420 ( .A(n338), .B(n10688), .Z(n10687) );
  XOR U10421 ( .A(n10689), .B(n10686), .Z(n10688) );
  XNOR U10422 ( .A(n8868), .B(n10682), .Z(n10684) );
  XOR U10423 ( .A(n10690), .B(n10691), .Z(n8868) );
  AND U10424 ( .A(n335), .B(n10692), .Z(n10691) );
  XOR U10425 ( .A(n10693), .B(n10690), .Z(n10692) );
  XOR U10426 ( .A(n10694), .B(n10695), .Z(n10682) );
  AND U10427 ( .A(n10696), .B(n10697), .Z(n10695) );
  XOR U10428 ( .A(n10694), .B(n8883), .Z(n10697) );
  XOR U10429 ( .A(n10698), .B(n10699), .Z(n8883) );
  AND U10430 ( .A(n338), .B(n10700), .Z(n10699) );
  XOR U10431 ( .A(n10701), .B(n10698), .Z(n10700) );
  XNOR U10432 ( .A(n8880), .B(n10694), .Z(n10696) );
  XOR U10433 ( .A(n10702), .B(n10703), .Z(n8880) );
  AND U10434 ( .A(n335), .B(n10704), .Z(n10703) );
  XOR U10435 ( .A(n10705), .B(n10702), .Z(n10704) );
  XOR U10436 ( .A(n10706), .B(n10707), .Z(n10694) );
  AND U10437 ( .A(n10708), .B(n10709), .Z(n10707) );
  XOR U10438 ( .A(n10706), .B(n8895), .Z(n10709) );
  XOR U10439 ( .A(n10710), .B(n10711), .Z(n8895) );
  AND U10440 ( .A(n338), .B(n10712), .Z(n10711) );
  XOR U10441 ( .A(n10713), .B(n10710), .Z(n10712) );
  XNOR U10442 ( .A(n8892), .B(n10706), .Z(n10708) );
  XOR U10443 ( .A(n10714), .B(n10715), .Z(n8892) );
  AND U10444 ( .A(n335), .B(n10716), .Z(n10715) );
  XOR U10445 ( .A(n10717), .B(n10714), .Z(n10716) );
  XOR U10446 ( .A(n10718), .B(n10719), .Z(n10706) );
  AND U10447 ( .A(n10720), .B(n10721), .Z(n10719) );
  XOR U10448 ( .A(n10718), .B(n8907), .Z(n10721) );
  XOR U10449 ( .A(n10722), .B(n10723), .Z(n8907) );
  AND U10450 ( .A(n338), .B(n10724), .Z(n10723) );
  XOR U10451 ( .A(n10725), .B(n10722), .Z(n10724) );
  XNOR U10452 ( .A(n8904), .B(n10718), .Z(n10720) );
  XOR U10453 ( .A(n10726), .B(n10727), .Z(n8904) );
  AND U10454 ( .A(n335), .B(n10728), .Z(n10727) );
  XOR U10455 ( .A(n10729), .B(n10726), .Z(n10728) );
  XOR U10456 ( .A(n10730), .B(n10731), .Z(n10718) );
  AND U10457 ( .A(n10732), .B(n10733), .Z(n10731) );
  XOR U10458 ( .A(n10730), .B(n8919), .Z(n10733) );
  XOR U10459 ( .A(n10734), .B(n10735), .Z(n8919) );
  AND U10460 ( .A(n338), .B(n10736), .Z(n10735) );
  XOR U10461 ( .A(n10737), .B(n10734), .Z(n10736) );
  XNOR U10462 ( .A(n8916), .B(n10730), .Z(n10732) );
  XOR U10463 ( .A(n10738), .B(n10739), .Z(n8916) );
  AND U10464 ( .A(n335), .B(n10740), .Z(n10739) );
  XOR U10465 ( .A(n10741), .B(n10738), .Z(n10740) );
  XOR U10466 ( .A(n10742), .B(n10743), .Z(n10730) );
  AND U10467 ( .A(n10744), .B(n10745), .Z(n10743) );
  XOR U10468 ( .A(n10742), .B(n8931), .Z(n10745) );
  XOR U10469 ( .A(n10746), .B(n10747), .Z(n8931) );
  AND U10470 ( .A(n338), .B(n10748), .Z(n10747) );
  XOR U10471 ( .A(n10749), .B(n10746), .Z(n10748) );
  XNOR U10472 ( .A(n8928), .B(n10742), .Z(n10744) );
  XOR U10473 ( .A(n10750), .B(n10751), .Z(n8928) );
  AND U10474 ( .A(n335), .B(n10752), .Z(n10751) );
  XOR U10475 ( .A(n10753), .B(n10750), .Z(n10752) );
  XOR U10476 ( .A(n10754), .B(n10755), .Z(n10742) );
  AND U10477 ( .A(n10756), .B(n10757), .Z(n10755) );
  XOR U10478 ( .A(n10754), .B(n8943), .Z(n10757) );
  XOR U10479 ( .A(n10758), .B(n10759), .Z(n8943) );
  AND U10480 ( .A(n338), .B(n10760), .Z(n10759) );
  XOR U10481 ( .A(n10761), .B(n10758), .Z(n10760) );
  XNOR U10482 ( .A(n8940), .B(n10754), .Z(n10756) );
  XOR U10483 ( .A(n10762), .B(n10763), .Z(n8940) );
  AND U10484 ( .A(n335), .B(n10764), .Z(n10763) );
  XOR U10485 ( .A(n10765), .B(n10762), .Z(n10764) );
  XOR U10486 ( .A(n10766), .B(n10767), .Z(n10754) );
  AND U10487 ( .A(n10768), .B(n10769), .Z(n10767) );
  XOR U10488 ( .A(n10766), .B(n8955), .Z(n10769) );
  XOR U10489 ( .A(n10770), .B(n10771), .Z(n8955) );
  AND U10490 ( .A(n338), .B(n10772), .Z(n10771) );
  XOR U10491 ( .A(n10773), .B(n10770), .Z(n10772) );
  XNOR U10492 ( .A(n8952), .B(n10766), .Z(n10768) );
  XOR U10493 ( .A(n10774), .B(n10775), .Z(n8952) );
  AND U10494 ( .A(n335), .B(n10776), .Z(n10775) );
  XOR U10495 ( .A(n10777), .B(n10774), .Z(n10776) );
  XOR U10496 ( .A(n10778), .B(n10779), .Z(n10766) );
  AND U10497 ( .A(n10780), .B(n10781), .Z(n10779) );
  XOR U10498 ( .A(n10778), .B(n8967), .Z(n10781) );
  XOR U10499 ( .A(n10782), .B(n10783), .Z(n8967) );
  AND U10500 ( .A(n338), .B(n10784), .Z(n10783) );
  XOR U10501 ( .A(n10785), .B(n10782), .Z(n10784) );
  XNOR U10502 ( .A(n8964), .B(n10778), .Z(n10780) );
  XOR U10503 ( .A(n10786), .B(n10787), .Z(n8964) );
  AND U10504 ( .A(n335), .B(n10788), .Z(n10787) );
  XOR U10505 ( .A(n10789), .B(n10786), .Z(n10788) );
  XOR U10506 ( .A(n10790), .B(n10791), .Z(n10778) );
  AND U10507 ( .A(n10792), .B(n10793), .Z(n10791) );
  XOR U10508 ( .A(n10790), .B(n8979), .Z(n10793) );
  XOR U10509 ( .A(n10794), .B(n10795), .Z(n8979) );
  AND U10510 ( .A(n338), .B(n10796), .Z(n10795) );
  XOR U10511 ( .A(n10797), .B(n10794), .Z(n10796) );
  XNOR U10512 ( .A(n8976), .B(n10790), .Z(n10792) );
  XOR U10513 ( .A(n10798), .B(n10799), .Z(n8976) );
  AND U10514 ( .A(n335), .B(n10800), .Z(n10799) );
  XOR U10515 ( .A(n10801), .B(n10798), .Z(n10800) );
  XOR U10516 ( .A(n10802), .B(n10803), .Z(n10790) );
  AND U10517 ( .A(n10804), .B(n10805), .Z(n10803) );
  XOR U10518 ( .A(n10802), .B(n8991), .Z(n10805) );
  XOR U10519 ( .A(n10806), .B(n10807), .Z(n8991) );
  AND U10520 ( .A(n338), .B(n10808), .Z(n10807) );
  XOR U10521 ( .A(n10809), .B(n10806), .Z(n10808) );
  XNOR U10522 ( .A(n8988), .B(n10802), .Z(n10804) );
  XOR U10523 ( .A(n10810), .B(n10811), .Z(n8988) );
  AND U10524 ( .A(n335), .B(n10812), .Z(n10811) );
  XOR U10525 ( .A(n10813), .B(n10810), .Z(n10812) );
  XOR U10526 ( .A(n10814), .B(n10815), .Z(n10802) );
  AND U10527 ( .A(n10816), .B(n10817), .Z(n10815) );
  XOR U10528 ( .A(n10814), .B(n9003), .Z(n10817) );
  XOR U10529 ( .A(n10818), .B(n10819), .Z(n9003) );
  AND U10530 ( .A(n338), .B(n10820), .Z(n10819) );
  XOR U10531 ( .A(n10821), .B(n10818), .Z(n10820) );
  XNOR U10532 ( .A(n9000), .B(n10814), .Z(n10816) );
  XOR U10533 ( .A(n10822), .B(n10823), .Z(n9000) );
  AND U10534 ( .A(n335), .B(n10824), .Z(n10823) );
  XOR U10535 ( .A(n10825), .B(n10822), .Z(n10824) );
  XOR U10536 ( .A(n10826), .B(n10827), .Z(n10814) );
  AND U10537 ( .A(n10828), .B(n10829), .Z(n10827) );
  XOR U10538 ( .A(n10826), .B(n9015), .Z(n10829) );
  XOR U10539 ( .A(n10830), .B(n10831), .Z(n9015) );
  AND U10540 ( .A(n338), .B(n10832), .Z(n10831) );
  XOR U10541 ( .A(n10833), .B(n10830), .Z(n10832) );
  XNOR U10542 ( .A(n9012), .B(n10826), .Z(n10828) );
  XOR U10543 ( .A(n10834), .B(n10835), .Z(n9012) );
  AND U10544 ( .A(n335), .B(n10836), .Z(n10835) );
  XOR U10545 ( .A(n10837), .B(n10834), .Z(n10836) );
  XOR U10546 ( .A(n10838), .B(n10839), .Z(n10826) );
  AND U10547 ( .A(n10840), .B(n10841), .Z(n10839) );
  XOR U10548 ( .A(n10838), .B(n9027), .Z(n10841) );
  XOR U10549 ( .A(n10842), .B(n10843), .Z(n9027) );
  AND U10550 ( .A(n338), .B(n10844), .Z(n10843) );
  XOR U10551 ( .A(n10845), .B(n10842), .Z(n10844) );
  XNOR U10552 ( .A(n9024), .B(n10838), .Z(n10840) );
  XOR U10553 ( .A(n10846), .B(n10847), .Z(n9024) );
  AND U10554 ( .A(n335), .B(n10848), .Z(n10847) );
  XOR U10555 ( .A(n10849), .B(n10846), .Z(n10848) );
  XOR U10556 ( .A(n10850), .B(n10851), .Z(n10838) );
  AND U10557 ( .A(n10852), .B(n10853), .Z(n10851) );
  XOR U10558 ( .A(n9039), .B(n10850), .Z(n10853) );
  XOR U10559 ( .A(n10854), .B(n10855), .Z(n9039) );
  AND U10560 ( .A(n338), .B(n10856), .Z(n10855) );
  XOR U10561 ( .A(n10854), .B(n10857), .Z(n10856) );
  XNOR U10562 ( .A(n10850), .B(n9036), .Z(n10852) );
  XOR U10563 ( .A(n10858), .B(n10859), .Z(n9036) );
  AND U10564 ( .A(n335), .B(n10860), .Z(n10859) );
  XOR U10565 ( .A(n10858), .B(n10861), .Z(n10860) );
  XOR U10566 ( .A(n10862), .B(n10863), .Z(n10850) );
  AND U10567 ( .A(n10864), .B(n10865), .Z(n10863) );
  XNOR U10568 ( .A(n10866), .B(n9052), .Z(n10865) );
  XOR U10569 ( .A(n10867), .B(n10868), .Z(n9052) );
  AND U10570 ( .A(n338), .B(n10869), .Z(n10868) );
  XOR U10571 ( .A(n10870), .B(n10867), .Z(n10869) );
  XNOR U10572 ( .A(n9049), .B(n10862), .Z(n10864) );
  XOR U10573 ( .A(n10871), .B(n10872), .Z(n9049) );
  AND U10574 ( .A(n335), .B(n10873), .Z(n10872) );
  XOR U10575 ( .A(n10874), .B(n10871), .Z(n10873) );
  IV U10576 ( .A(n10866), .Z(n10862) );
  AND U10577 ( .A(n10498), .B(n10501), .Z(n10866) );
  XNOR U10578 ( .A(n10875), .B(n10876), .Z(n10501) );
  AND U10579 ( .A(n338), .B(n10877), .Z(n10876) );
  XNOR U10580 ( .A(n10878), .B(n10875), .Z(n10877) );
  XOR U10581 ( .A(n10879), .B(n10880), .Z(n338) );
  AND U10582 ( .A(n10881), .B(n10882), .Z(n10880) );
  XOR U10583 ( .A(n10509), .B(n10879), .Z(n10882) );
  IV U10584 ( .A(n10883), .Z(n10509) );
  AND U10585 ( .A(p_input[2815]), .B(p_input[2783]), .Z(n10883) );
  XOR U10586 ( .A(n10879), .B(n10506), .Z(n10881) );
  AND U10587 ( .A(p_input[2719]), .B(p_input[2751]), .Z(n10506) );
  XOR U10588 ( .A(n10884), .B(n10885), .Z(n10879) );
  AND U10589 ( .A(n10886), .B(n10887), .Z(n10885) );
  XOR U10590 ( .A(n10884), .B(n10521), .Z(n10887) );
  XNOR U10591 ( .A(p_input[2782]), .B(n10888), .Z(n10521) );
  AND U10592 ( .A(n254), .B(n10889), .Z(n10888) );
  XOR U10593 ( .A(p_input[2814]), .B(p_input[2782]), .Z(n10889) );
  XNOR U10594 ( .A(n10518), .B(n10884), .Z(n10886) );
  XOR U10595 ( .A(n10890), .B(n10891), .Z(n10518) );
  AND U10596 ( .A(n252), .B(n10892), .Z(n10891) );
  XOR U10597 ( .A(p_input[2750]), .B(p_input[2718]), .Z(n10892) );
  XOR U10598 ( .A(n10893), .B(n10894), .Z(n10884) );
  AND U10599 ( .A(n10895), .B(n10896), .Z(n10894) );
  XOR U10600 ( .A(n10893), .B(n10533), .Z(n10896) );
  XNOR U10601 ( .A(p_input[2781]), .B(n10897), .Z(n10533) );
  AND U10602 ( .A(n254), .B(n10898), .Z(n10897) );
  XOR U10603 ( .A(p_input[2813]), .B(p_input[2781]), .Z(n10898) );
  XNOR U10604 ( .A(n10530), .B(n10893), .Z(n10895) );
  XOR U10605 ( .A(n10899), .B(n10900), .Z(n10530) );
  AND U10606 ( .A(n252), .B(n10901), .Z(n10900) );
  XOR U10607 ( .A(p_input[2749]), .B(p_input[2717]), .Z(n10901) );
  XOR U10608 ( .A(n10902), .B(n10903), .Z(n10893) );
  AND U10609 ( .A(n10904), .B(n10905), .Z(n10903) );
  XOR U10610 ( .A(n10902), .B(n10545), .Z(n10905) );
  XNOR U10611 ( .A(p_input[2780]), .B(n10906), .Z(n10545) );
  AND U10612 ( .A(n254), .B(n10907), .Z(n10906) );
  XOR U10613 ( .A(p_input[2812]), .B(p_input[2780]), .Z(n10907) );
  XNOR U10614 ( .A(n10542), .B(n10902), .Z(n10904) );
  XOR U10615 ( .A(n10908), .B(n10909), .Z(n10542) );
  AND U10616 ( .A(n252), .B(n10910), .Z(n10909) );
  XOR U10617 ( .A(p_input[2748]), .B(p_input[2716]), .Z(n10910) );
  XOR U10618 ( .A(n10911), .B(n10912), .Z(n10902) );
  AND U10619 ( .A(n10913), .B(n10914), .Z(n10912) );
  XOR U10620 ( .A(n10911), .B(n10557), .Z(n10914) );
  XNOR U10621 ( .A(p_input[2779]), .B(n10915), .Z(n10557) );
  AND U10622 ( .A(n254), .B(n10916), .Z(n10915) );
  XOR U10623 ( .A(p_input[2811]), .B(p_input[2779]), .Z(n10916) );
  XNOR U10624 ( .A(n10554), .B(n10911), .Z(n10913) );
  XOR U10625 ( .A(n10917), .B(n10918), .Z(n10554) );
  AND U10626 ( .A(n252), .B(n10919), .Z(n10918) );
  XOR U10627 ( .A(p_input[2747]), .B(p_input[2715]), .Z(n10919) );
  XOR U10628 ( .A(n10920), .B(n10921), .Z(n10911) );
  AND U10629 ( .A(n10922), .B(n10923), .Z(n10921) );
  XOR U10630 ( .A(n10920), .B(n10569), .Z(n10923) );
  XNOR U10631 ( .A(p_input[2778]), .B(n10924), .Z(n10569) );
  AND U10632 ( .A(n254), .B(n10925), .Z(n10924) );
  XOR U10633 ( .A(p_input[2810]), .B(p_input[2778]), .Z(n10925) );
  XNOR U10634 ( .A(n10566), .B(n10920), .Z(n10922) );
  XOR U10635 ( .A(n10926), .B(n10927), .Z(n10566) );
  AND U10636 ( .A(n252), .B(n10928), .Z(n10927) );
  XOR U10637 ( .A(p_input[2746]), .B(p_input[2714]), .Z(n10928) );
  XOR U10638 ( .A(n10929), .B(n10930), .Z(n10920) );
  AND U10639 ( .A(n10931), .B(n10932), .Z(n10930) );
  XOR U10640 ( .A(n10929), .B(n10581), .Z(n10932) );
  XNOR U10641 ( .A(p_input[2777]), .B(n10933), .Z(n10581) );
  AND U10642 ( .A(n254), .B(n10934), .Z(n10933) );
  XOR U10643 ( .A(p_input[2809]), .B(p_input[2777]), .Z(n10934) );
  XNOR U10644 ( .A(n10578), .B(n10929), .Z(n10931) );
  XOR U10645 ( .A(n10935), .B(n10936), .Z(n10578) );
  AND U10646 ( .A(n252), .B(n10937), .Z(n10936) );
  XOR U10647 ( .A(p_input[2745]), .B(p_input[2713]), .Z(n10937) );
  XOR U10648 ( .A(n10938), .B(n10939), .Z(n10929) );
  AND U10649 ( .A(n10940), .B(n10941), .Z(n10939) );
  XOR U10650 ( .A(n10938), .B(n10593), .Z(n10941) );
  XNOR U10651 ( .A(p_input[2776]), .B(n10942), .Z(n10593) );
  AND U10652 ( .A(n254), .B(n10943), .Z(n10942) );
  XOR U10653 ( .A(p_input[2808]), .B(p_input[2776]), .Z(n10943) );
  XNOR U10654 ( .A(n10590), .B(n10938), .Z(n10940) );
  XOR U10655 ( .A(n10944), .B(n10945), .Z(n10590) );
  AND U10656 ( .A(n252), .B(n10946), .Z(n10945) );
  XOR U10657 ( .A(p_input[2744]), .B(p_input[2712]), .Z(n10946) );
  XOR U10658 ( .A(n10947), .B(n10948), .Z(n10938) );
  AND U10659 ( .A(n10949), .B(n10950), .Z(n10948) );
  XOR U10660 ( .A(n10947), .B(n10605), .Z(n10950) );
  XNOR U10661 ( .A(p_input[2775]), .B(n10951), .Z(n10605) );
  AND U10662 ( .A(n254), .B(n10952), .Z(n10951) );
  XOR U10663 ( .A(p_input[2807]), .B(p_input[2775]), .Z(n10952) );
  XNOR U10664 ( .A(n10602), .B(n10947), .Z(n10949) );
  XOR U10665 ( .A(n10953), .B(n10954), .Z(n10602) );
  AND U10666 ( .A(n252), .B(n10955), .Z(n10954) );
  XOR U10667 ( .A(p_input[2743]), .B(p_input[2711]), .Z(n10955) );
  XOR U10668 ( .A(n10956), .B(n10957), .Z(n10947) );
  AND U10669 ( .A(n10958), .B(n10959), .Z(n10957) );
  XOR U10670 ( .A(n10956), .B(n10617), .Z(n10959) );
  XNOR U10671 ( .A(p_input[2774]), .B(n10960), .Z(n10617) );
  AND U10672 ( .A(n254), .B(n10961), .Z(n10960) );
  XOR U10673 ( .A(p_input[2806]), .B(p_input[2774]), .Z(n10961) );
  XNOR U10674 ( .A(n10614), .B(n10956), .Z(n10958) );
  XOR U10675 ( .A(n10962), .B(n10963), .Z(n10614) );
  AND U10676 ( .A(n252), .B(n10964), .Z(n10963) );
  XOR U10677 ( .A(p_input[2742]), .B(p_input[2710]), .Z(n10964) );
  XOR U10678 ( .A(n10965), .B(n10966), .Z(n10956) );
  AND U10679 ( .A(n10967), .B(n10968), .Z(n10966) );
  XOR U10680 ( .A(n10965), .B(n10629), .Z(n10968) );
  XNOR U10681 ( .A(p_input[2773]), .B(n10969), .Z(n10629) );
  AND U10682 ( .A(n254), .B(n10970), .Z(n10969) );
  XOR U10683 ( .A(p_input[2805]), .B(p_input[2773]), .Z(n10970) );
  XNOR U10684 ( .A(n10626), .B(n10965), .Z(n10967) );
  XOR U10685 ( .A(n10971), .B(n10972), .Z(n10626) );
  AND U10686 ( .A(n252), .B(n10973), .Z(n10972) );
  XOR U10687 ( .A(p_input[2741]), .B(p_input[2709]), .Z(n10973) );
  XOR U10688 ( .A(n10974), .B(n10975), .Z(n10965) );
  AND U10689 ( .A(n10976), .B(n10977), .Z(n10975) );
  XOR U10690 ( .A(n10974), .B(n10641), .Z(n10977) );
  XNOR U10691 ( .A(p_input[2772]), .B(n10978), .Z(n10641) );
  AND U10692 ( .A(n254), .B(n10979), .Z(n10978) );
  XOR U10693 ( .A(p_input[2804]), .B(p_input[2772]), .Z(n10979) );
  XNOR U10694 ( .A(n10638), .B(n10974), .Z(n10976) );
  XOR U10695 ( .A(n10980), .B(n10981), .Z(n10638) );
  AND U10696 ( .A(n252), .B(n10982), .Z(n10981) );
  XOR U10697 ( .A(p_input[2740]), .B(p_input[2708]), .Z(n10982) );
  XOR U10698 ( .A(n10983), .B(n10984), .Z(n10974) );
  AND U10699 ( .A(n10985), .B(n10986), .Z(n10984) );
  XOR U10700 ( .A(n10983), .B(n10653), .Z(n10986) );
  XNOR U10701 ( .A(p_input[2771]), .B(n10987), .Z(n10653) );
  AND U10702 ( .A(n254), .B(n10988), .Z(n10987) );
  XOR U10703 ( .A(p_input[2803]), .B(p_input[2771]), .Z(n10988) );
  XNOR U10704 ( .A(n10650), .B(n10983), .Z(n10985) );
  XOR U10705 ( .A(n10989), .B(n10990), .Z(n10650) );
  AND U10706 ( .A(n252), .B(n10991), .Z(n10990) );
  XOR U10707 ( .A(p_input[2739]), .B(p_input[2707]), .Z(n10991) );
  XOR U10708 ( .A(n10992), .B(n10993), .Z(n10983) );
  AND U10709 ( .A(n10994), .B(n10995), .Z(n10993) );
  XOR U10710 ( .A(n10992), .B(n10665), .Z(n10995) );
  XNOR U10711 ( .A(p_input[2770]), .B(n10996), .Z(n10665) );
  AND U10712 ( .A(n254), .B(n10997), .Z(n10996) );
  XOR U10713 ( .A(p_input[2802]), .B(p_input[2770]), .Z(n10997) );
  XNOR U10714 ( .A(n10662), .B(n10992), .Z(n10994) );
  XOR U10715 ( .A(n10998), .B(n10999), .Z(n10662) );
  AND U10716 ( .A(n252), .B(n11000), .Z(n10999) );
  XOR U10717 ( .A(p_input[2738]), .B(p_input[2706]), .Z(n11000) );
  XOR U10718 ( .A(n11001), .B(n11002), .Z(n10992) );
  AND U10719 ( .A(n11003), .B(n11004), .Z(n11002) );
  XOR U10720 ( .A(n11001), .B(n10677), .Z(n11004) );
  XNOR U10721 ( .A(p_input[2769]), .B(n11005), .Z(n10677) );
  AND U10722 ( .A(n254), .B(n11006), .Z(n11005) );
  XOR U10723 ( .A(p_input[2801]), .B(p_input[2769]), .Z(n11006) );
  XNOR U10724 ( .A(n10674), .B(n11001), .Z(n11003) );
  XOR U10725 ( .A(n11007), .B(n11008), .Z(n10674) );
  AND U10726 ( .A(n252), .B(n11009), .Z(n11008) );
  XOR U10727 ( .A(p_input[2737]), .B(p_input[2705]), .Z(n11009) );
  XOR U10728 ( .A(n11010), .B(n11011), .Z(n11001) );
  AND U10729 ( .A(n11012), .B(n11013), .Z(n11011) );
  XOR U10730 ( .A(n11010), .B(n10689), .Z(n11013) );
  XNOR U10731 ( .A(p_input[2768]), .B(n11014), .Z(n10689) );
  AND U10732 ( .A(n254), .B(n11015), .Z(n11014) );
  XOR U10733 ( .A(p_input[2800]), .B(p_input[2768]), .Z(n11015) );
  XNOR U10734 ( .A(n10686), .B(n11010), .Z(n11012) );
  XOR U10735 ( .A(n11016), .B(n11017), .Z(n10686) );
  AND U10736 ( .A(n252), .B(n11018), .Z(n11017) );
  XOR U10737 ( .A(p_input[2736]), .B(p_input[2704]), .Z(n11018) );
  XOR U10738 ( .A(n11019), .B(n11020), .Z(n11010) );
  AND U10739 ( .A(n11021), .B(n11022), .Z(n11020) );
  XOR U10740 ( .A(n11019), .B(n10701), .Z(n11022) );
  XNOR U10741 ( .A(p_input[2767]), .B(n11023), .Z(n10701) );
  AND U10742 ( .A(n254), .B(n11024), .Z(n11023) );
  XOR U10743 ( .A(p_input[2799]), .B(p_input[2767]), .Z(n11024) );
  XNOR U10744 ( .A(n10698), .B(n11019), .Z(n11021) );
  XOR U10745 ( .A(n11025), .B(n11026), .Z(n10698) );
  AND U10746 ( .A(n252), .B(n11027), .Z(n11026) );
  XOR U10747 ( .A(p_input[2735]), .B(p_input[2703]), .Z(n11027) );
  XOR U10748 ( .A(n11028), .B(n11029), .Z(n11019) );
  AND U10749 ( .A(n11030), .B(n11031), .Z(n11029) );
  XOR U10750 ( .A(n11028), .B(n10713), .Z(n11031) );
  XNOR U10751 ( .A(p_input[2766]), .B(n11032), .Z(n10713) );
  AND U10752 ( .A(n254), .B(n11033), .Z(n11032) );
  XOR U10753 ( .A(p_input[2798]), .B(p_input[2766]), .Z(n11033) );
  XNOR U10754 ( .A(n10710), .B(n11028), .Z(n11030) );
  XOR U10755 ( .A(n11034), .B(n11035), .Z(n10710) );
  AND U10756 ( .A(n252), .B(n11036), .Z(n11035) );
  XOR U10757 ( .A(p_input[2734]), .B(p_input[2702]), .Z(n11036) );
  XOR U10758 ( .A(n11037), .B(n11038), .Z(n11028) );
  AND U10759 ( .A(n11039), .B(n11040), .Z(n11038) );
  XOR U10760 ( .A(n11037), .B(n10725), .Z(n11040) );
  XNOR U10761 ( .A(p_input[2765]), .B(n11041), .Z(n10725) );
  AND U10762 ( .A(n254), .B(n11042), .Z(n11041) );
  XOR U10763 ( .A(p_input[2797]), .B(p_input[2765]), .Z(n11042) );
  XNOR U10764 ( .A(n10722), .B(n11037), .Z(n11039) );
  XOR U10765 ( .A(n11043), .B(n11044), .Z(n10722) );
  AND U10766 ( .A(n252), .B(n11045), .Z(n11044) );
  XOR U10767 ( .A(p_input[2733]), .B(p_input[2701]), .Z(n11045) );
  XOR U10768 ( .A(n11046), .B(n11047), .Z(n11037) );
  AND U10769 ( .A(n11048), .B(n11049), .Z(n11047) );
  XOR U10770 ( .A(n11046), .B(n10737), .Z(n11049) );
  XNOR U10771 ( .A(p_input[2764]), .B(n11050), .Z(n10737) );
  AND U10772 ( .A(n254), .B(n11051), .Z(n11050) );
  XOR U10773 ( .A(p_input[2796]), .B(p_input[2764]), .Z(n11051) );
  XNOR U10774 ( .A(n10734), .B(n11046), .Z(n11048) );
  XOR U10775 ( .A(n11052), .B(n11053), .Z(n10734) );
  AND U10776 ( .A(n252), .B(n11054), .Z(n11053) );
  XOR U10777 ( .A(p_input[2732]), .B(p_input[2700]), .Z(n11054) );
  XOR U10778 ( .A(n11055), .B(n11056), .Z(n11046) );
  AND U10779 ( .A(n11057), .B(n11058), .Z(n11056) );
  XOR U10780 ( .A(n11055), .B(n10749), .Z(n11058) );
  XNOR U10781 ( .A(p_input[2763]), .B(n11059), .Z(n10749) );
  AND U10782 ( .A(n254), .B(n11060), .Z(n11059) );
  XOR U10783 ( .A(p_input[2795]), .B(p_input[2763]), .Z(n11060) );
  XNOR U10784 ( .A(n10746), .B(n11055), .Z(n11057) );
  XOR U10785 ( .A(n11061), .B(n11062), .Z(n10746) );
  AND U10786 ( .A(n252), .B(n11063), .Z(n11062) );
  XOR U10787 ( .A(p_input[2731]), .B(p_input[2699]), .Z(n11063) );
  XOR U10788 ( .A(n11064), .B(n11065), .Z(n11055) );
  AND U10789 ( .A(n11066), .B(n11067), .Z(n11065) );
  XOR U10790 ( .A(n11064), .B(n10761), .Z(n11067) );
  XNOR U10791 ( .A(p_input[2762]), .B(n11068), .Z(n10761) );
  AND U10792 ( .A(n254), .B(n11069), .Z(n11068) );
  XOR U10793 ( .A(p_input[2794]), .B(p_input[2762]), .Z(n11069) );
  XNOR U10794 ( .A(n10758), .B(n11064), .Z(n11066) );
  XOR U10795 ( .A(n11070), .B(n11071), .Z(n10758) );
  AND U10796 ( .A(n252), .B(n11072), .Z(n11071) );
  XOR U10797 ( .A(p_input[2730]), .B(p_input[2698]), .Z(n11072) );
  XOR U10798 ( .A(n11073), .B(n11074), .Z(n11064) );
  AND U10799 ( .A(n11075), .B(n11076), .Z(n11074) );
  XOR U10800 ( .A(n11073), .B(n10773), .Z(n11076) );
  XNOR U10801 ( .A(p_input[2761]), .B(n11077), .Z(n10773) );
  AND U10802 ( .A(n254), .B(n11078), .Z(n11077) );
  XOR U10803 ( .A(p_input[2793]), .B(p_input[2761]), .Z(n11078) );
  XNOR U10804 ( .A(n10770), .B(n11073), .Z(n11075) );
  XOR U10805 ( .A(n11079), .B(n11080), .Z(n10770) );
  AND U10806 ( .A(n252), .B(n11081), .Z(n11080) );
  XOR U10807 ( .A(p_input[2729]), .B(p_input[2697]), .Z(n11081) );
  XOR U10808 ( .A(n11082), .B(n11083), .Z(n11073) );
  AND U10809 ( .A(n11084), .B(n11085), .Z(n11083) );
  XOR U10810 ( .A(n11082), .B(n10785), .Z(n11085) );
  XNOR U10811 ( .A(p_input[2760]), .B(n11086), .Z(n10785) );
  AND U10812 ( .A(n254), .B(n11087), .Z(n11086) );
  XOR U10813 ( .A(p_input[2792]), .B(p_input[2760]), .Z(n11087) );
  XNOR U10814 ( .A(n10782), .B(n11082), .Z(n11084) );
  XOR U10815 ( .A(n11088), .B(n11089), .Z(n10782) );
  AND U10816 ( .A(n252), .B(n11090), .Z(n11089) );
  XOR U10817 ( .A(p_input[2728]), .B(p_input[2696]), .Z(n11090) );
  XOR U10818 ( .A(n11091), .B(n11092), .Z(n11082) );
  AND U10819 ( .A(n11093), .B(n11094), .Z(n11092) );
  XOR U10820 ( .A(n11091), .B(n10797), .Z(n11094) );
  XNOR U10821 ( .A(p_input[2759]), .B(n11095), .Z(n10797) );
  AND U10822 ( .A(n254), .B(n11096), .Z(n11095) );
  XOR U10823 ( .A(p_input[2791]), .B(p_input[2759]), .Z(n11096) );
  XNOR U10824 ( .A(n10794), .B(n11091), .Z(n11093) );
  XOR U10825 ( .A(n11097), .B(n11098), .Z(n10794) );
  AND U10826 ( .A(n252), .B(n11099), .Z(n11098) );
  XOR U10827 ( .A(p_input[2727]), .B(p_input[2695]), .Z(n11099) );
  XOR U10828 ( .A(n11100), .B(n11101), .Z(n11091) );
  AND U10829 ( .A(n11102), .B(n11103), .Z(n11101) );
  XOR U10830 ( .A(n11100), .B(n10809), .Z(n11103) );
  XNOR U10831 ( .A(p_input[2758]), .B(n11104), .Z(n10809) );
  AND U10832 ( .A(n254), .B(n11105), .Z(n11104) );
  XOR U10833 ( .A(p_input[2790]), .B(p_input[2758]), .Z(n11105) );
  XNOR U10834 ( .A(n10806), .B(n11100), .Z(n11102) );
  XOR U10835 ( .A(n11106), .B(n11107), .Z(n10806) );
  AND U10836 ( .A(n252), .B(n11108), .Z(n11107) );
  XOR U10837 ( .A(p_input[2726]), .B(p_input[2694]), .Z(n11108) );
  XOR U10838 ( .A(n11109), .B(n11110), .Z(n11100) );
  AND U10839 ( .A(n11111), .B(n11112), .Z(n11110) );
  XOR U10840 ( .A(n11109), .B(n10821), .Z(n11112) );
  XNOR U10841 ( .A(p_input[2757]), .B(n11113), .Z(n10821) );
  AND U10842 ( .A(n254), .B(n11114), .Z(n11113) );
  XOR U10843 ( .A(p_input[2789]), .B(p_input[2757]), .Z(n11114) );
  XNOR U10844 ( .A(n10818), .B(n11109), .Z(n11111) );
  XOR U10845 ( .A(n11115), .B(n11116), .Z(n10818) );
  AND U10846 ( .A(n252), .B(n11117), .Z(n11116) );
  XOR U10847 ( .A(p_input[2725]), .B(p_input[2693]), .Z(n11117) );
  XOR U10848 ( .A(n11118), .B(n11119), .Z(n11109) );
  AND U10849 ( .A(n11120), .B(n11121), .Z(n11119) );
  XOR U10850 ( .A(n11118), .B(n10833), .Z(n11121) );
  XNOR U10851 ( .A(p_input[2756]), .B(n11122), .Z(n10833) );
  AND U10852 ( .A(n254), .B(n11123), .Z(n11122) );
  XOR U10853 ( .A(p_input[2788]), .B(p_input[2756]), .Z(n11123) );
  XNOR U10854 ( .A(n10830), .B(n11118), .Z(n11120) );
  XOR U10855 ( .A(n11124), .B(n11125), .Z(n10830) );
  AND U10856 ( .A(n252), .B(n11126), .Z(n11125) );
  XOR U10857 ( .A(p_input[2724]), .B(p_input[2692]), .Z(n11126) );
  XOR U10858 ( .A(n11127), .B(n11128), .Z(n11118) );
  AND U10859 ( .A(n11129), .B(n11130), .Z(n11128) );
  XOR U10860 ( .A(n11127), .B(n10845), .Z(n11130) );
  XNOR U10861 ( .A(p_input[2755]), .B(n11131), .Z(n10845) );
  AND U10862 ( .A(n254), .B(n11132), .Z(n11131) );
  XOR U10863 ( .A(p_input[2787]), .B(p_input[2755]), .Z(n11132) );
  XNOR U10864 ( .A(n10842), .B(n11127), .Z(n11129) );
  XOR U10865 ( .A(n11133), .B(n11134), .Z(n10842) );
  AND U10866 ( .A(n252), .B(n11135), .Z(n11134) );
  XOR U10867 ( .A(p_input[2723]), .B(p_input[2691]), .Z(n11135) );
  XOR U10868 ( .A(n11136), .B(n11137), .Z(n11127) );
  AND U10869 ( .A(n11138), .B(n11139), .Z(n11137) );
  XOR U10870 ( .A(n10857), .B(n11136), .Z(n11139) );
  XNOR U10871 ( .A(p_input[2754]), .B(n11140), .Z(n10857) );
  AND U10872 ( .A(n254), .B(n11141), .Z(n11140) );
  XOR U10873 ( .A(p_input[2786]), .B(p_input[2754]), .Z(n11141) );
  XNOR U10874 ( .A(n11136), .B(n10854), .Z(n11138) );
  XOR U10875 ( .A(n11142), .B(n11143), .Z(n10854) );
  AND U10876 ( .A(n252), .B(n11144), .Z(n11143) );
  XOR U10877 ( .A(p_input[2722]), .B(p_input[2690]), .Z(n11144) );
  XOR U10878 ( .A(n11145), .B(n11146), .Z(n11136) );
  AND U10879 ( .A(n11147), .B(n11148), .Z(n11146) );
  XNOR U10880 ( .A(n11149), .B(n10870), .Z(n11148) );
  XNOR U10881 ( .A(p_input[2753]), .B(n11150), .Z(n10870) );
  AND U10882 ( .A(n254), .B(n11151), .Z(n11150) );
  XNOR U10883 ( .A(p_input[2785]), .B(n11152), .Z(n11151) );
  IV U10884 ( .A(p_input[2753]), .Z(n11152) );
  XNOR U10885 ( .A(n10867), .B(n11145), .Z(n11147) );
  XNOR U10886 ( .A(p_input[2689]), .B(n11153), .Z(n10867) );
  AND U10887 ( .A(n252), .B(n11154), .Z(n11153) );
  XOR U10888 ( .A(p_input[2721]), .B(p_input[2689]), .Z(n11154) );
  IV U10889 ( .A(n11149), .Z(n11145) );
  AND U10890 ( .A(n10875), .B(n10878), .Z(n11149) );
  XOR U10891 ( .A(p_input[2752]), .B(n11155), .Z(n10878) );
  AND U10892 ( .A(n254), .B(n11156), .Z(n11155) );
  XOR U10893 ( .A(p_input[2784]), .B(p_input[2752]), .Z(n11156) );
  XOR U10894 ( .A(n11157), .B(n11158), .Z(n254) );
  AND U10895 ( .A(n11159), .B(n11160), .Z(n11158) );
  XNOR U10896 ( .A(p_input[2815]), .B(n11157), .Z(n11160) );
  XOR U10897 ( .A(n11157), .B(p_input[2783]), .Z(n11159) );
  XOR U10898 ( .A(n11161), .B(n11162), .Z(n11157) );
  AND U10899 ( .A(n11163), .B(n11164), .Z(n11162) );
  XNOR U10900 ( .A(p_input[2814]), .B(n11161), .Z(n11164) );
  XOR U10901 ( .A(n11161), .B(p_input[2782]), .Z(n11163) );
  XOR U10902 ( .A(n11165), .B(n11166), .Z(n11161) );
  AND U10903 ( .A(n11167), .B(n11168), .Z(n11166) );
  XNOR U10904 ( .A(p_input[2813]), .B(n11165), .Z(n11168) );
  XOR U10905 ( .A(n11165), .B(p_input[2781]), .Z(n11167) );
  XOR U10906 ( .A(n11169), .B(n11170), .Z(n11165) );
  AND U10907 ( .A(n11171), .B(n11172), .Z(n11170) );
  XNOR U10908 ( .A(p_input[2812]), .B(n11169), .Z(n11172) );
  XOR U10909 ( .A(n11169), .B(p_input[2780]), .Z(n11171) );
  XOR U10910 ( .A(n11173), .B(n11174), .Z(n11169) );
  AND U10911 ( .A(n11175), .B(n11176), .Z(n11174) );
  XNOR U10912 ( .A(p_input[2811]), .B(n11173), .Z(n11176) );
  XOR U10913 ( .A(n11173), .B(p_input[2779]), .Z(n11175) );
  XOR U10914 ( .A(n11177), .B(n11178), .Z(n11173) );
  AND U10915 ( .A(n11179), .B(n11180), .Z(n11178) );
  XNOR U10916 ( .A(p_input[2810]), .B(n11177), .Z(n11180) );
  XOR U10917 ( .A(n11177), .B(p_input[2778]), .Z(n11179) );
  XOR U10918 ( .A(n11181), .B(n11182), .Z(n11177) );
  AND U10919 ( .A(n11183), .B(n11184), .Z(n11182) );
  XNOR U10920 ( .A(p_input[2809]), .B(n11181), .Z(n11184) );
  XOR U10921 ( .A(n11181), .B(p_input[2777]), .Z(n11183) );
  XOR U10922 ( .A(n11185), .B(n11186), .Z(n11181) );
  AND U10923 ( .A(n11187), .B(n11188), .Z(n11186) );
  XNOR U10924 ( .A(p_input[2808]), .B(n11185), .Z(n11188) );
  XOR U10925 ( .A(n11185), .B(p_input[2776]), .Z(n11187) );
  XOR U10926 ( .A(n11189), .B(n11190), .Z(n11185) );
  AND U10927 ( .A(n11191), .B(n11192), .Z(n11190) );
  XNOR U10928 ( .A(p_input[2807]), .B(n11189), .Z(n11192) );
  XOR U10929 ( .A(n11189), .B(p_input[2775]), .Z(n11191) );
  XOR U10930 ( .A(n11193), .B(n11194), .Z(n11189) );
  AND U10931 ( .A(n11195), .B(n11196), .Z(n11194) );
  XNOR U10932 ( .A(p_input[2806]), .B(n11193), .Z(n11196) );
  XOR U10933 ( .A(n11193), .B(p_input[2774]), .Z(n11195) );
  XOR U10934 ( .A(n11197), .B(n11198), .Z(n11193) );
  AND U10935 ( .A(n11199), .B(n11200), .Z(n11198) );
  XNOR U10936 ( .A(p_input[2805]), .B(n11197), .Z(n11200) );
  XOR U10937 ( .A(n11197), .B(p_input[2773]), .Z(n11199) );
  XOR U10938 ( .A(n11201), .B(n11202), .Z(n11197) );
  AND U10939 ( .A(n11203), .B(n11204), .Z(n11202) );
  XNOR U10940 ( .A(p_input[2804]), .B(n11201), .Z(n11204) );
  XOR U10941 ( .A(n11201), .B(p_input[2772]), .Z(n11203) );
  XOR U10942 ( .A(n11205), .B(n11206), .Z(n11201) );
  AND U10943 ( .A(n11207), .B(n11208), .Z(n11206) );
  XNOR U10944 ( .A(p_input[2803]), .B(n11205), .Z(n11208) );
  XOR U10945 ( .A(n11205), .B(p_input[2771]), .Z(n11207) );
  XOR U10946 ( .A(n11209), .B(n11210), .Z(n11205) );
  AND U10947 ( .A(n11211), .B(n11212), .Z(n11210) );
  XNOR U10948 ( .A(p_input[2802]), .B(n11209), .Z(n11212) );
  XOR U10949 ( .A(n11209), .B(p_input[2770]), .Z(n11211) );
  XOR U10950 ( .A(n11213), .B(n11214), .Z(n11209) );
  AND U10951 ( .A(n11215), .B(n11216), .Z(n11214) );
  XNOR U10952 ( .A(p_input[2801]), .B(n11213), .Z(n11216) );
  XOR U10953 ( .A(n11213), .B(p_input[2769]), .Z(n11215) );
  XOR U10954 ( .A(n11217), .B(n11218), .Z(n11213) );
  AND U10955 ( .A(n11219), .B(n11220), .Z(n11218) );
  XNOR U10956 ( .A(p_input[2800]), .B(n11217), .Z(n11220) );
  XOR U10957 ( .A(n11217), .B(p_input[2768]), .Z(n11219) );
  XOR U10958 ( .A(n11221), .B(n11222), .Z(n11217) );
  AND U10959 ( .A(n11223), .B(n11224), .Z(n11222) );
  XNOR U10960 ( .A(p_input[2799]), .B(n11221), .Z(n11224) );
  XOR U10961 ( .A(n11221), .B(p_input[2767]), .Z(n11223) );
  XOR U10962 ( .A(n11225), .B(n11226), .Z(n11221) );
  AND U10963 ( .A(n11227), .B(n11228), .Z(n11226) );
  XNOR U10964 ( .A(p_input[2798]), .B(n11225), .Z(n11228) );
  XOR U10965 ( .A(n11225), .B(p_input[2766]), .Z(n11227) );
  XOR U10966 ( .A(n11229), .B(n11230), .Z(n11225) );
  AND U10967 ( .A(n11231), .B(n11232), .Z(n11230) );
  XNOR U10968 ( .A(p_input[2797]), .B(n11229), .Z(n11232) );
  XOR U10969 ( .A(n11229), .B(p_input[2765]), .Z(n11231) );
  XOR U10970 ( .A(n11233), .B(n11234), .Z(n11229) );
  AND U10971 ( .A(n11235), .B(n11236), .Z(n11234) );
  XNOR U10972 ( .A(p_input[2796]), .B(n11233), .Z(n11236) );
  XOR U10973 ( .A(n11233), .B(p_input[2764]), .Z(n11235) );
  XOR U10974 ( .A(n11237), .B(n11238), .Z(n11233) );
  AND U10975 ( .A(n11239), .B(n11240), .Z(n11238) );
  XNOR U10976 ( .A(p_input[2795]), .B(n11237), .Z(n11240) );
  XOR U10977 ( .A(n11237), .B(p_input[2763]), .Z(n11239) );
  XOR U10978 ( .A(n11241), .B(n11242), .Z(n11237) );
  AND U10979 ( .A(n11243), .B(n11244), .Z(n11242) );
  XNOR U10980 ( .A(p_input[2794]), .B(n11241), .Z(n11244) );
  XOR U10981 ( .A(n11241), .B(p_input[2762]), .Z(n11243) );
  XOR U10982 ( .A(n11245), .B(n11246), .Z(n11241) );
  AND U10983 ( .A(n11247), .B(n11248), .Z(n11246) );
  XNOR U10984 ( .A(p_input[2793]), .B(n11245), .Z(n11248) );
  XOR U10985 ( .A(n11245), .B(p_input[2761]), .Z(n11247) );
  XOR U10986 ( .A(n11249), .B(n11250), .Z(n11245) );
  AND U10987 ( .A(n11251), .B(n11252), .Z(n11250) );
  XNOR U10988 ( .A(p_input[2792]), .B(n11249), .Z(n11252) );
  XOR U10989 ( .A(n11249), .B(p_input[2760]), .Z(n11251) );
  XOR U10990 ( .A(n11253), .B(n11254), .Z(n11249) );
  AND U10991 ( .A(n11255), .B(n11256), .Z(n11254) );
  XNOR U10992 ( .A(p_input[2791]), .B(n11253), .Z(n11256) );
  XOR U10993 ( .A(n11253), .B(p_input[2759]), .Z(n11255) );
  XOR U10994 ( .A(n11257), .B(n11258), .Z(n11253) );
  AND U10995 ( .A(n11259), .B(n11260), .Z(n11258) );
  XNOR U10996 ( .A(p_input[2790]), .B(n11257), .Z(n11260) );
  XOR U10997 ( .A(n11257), .B(p_input[2758]), .Z(n11259) );
  XOR U10998 ( .A(n11261), .B(n11262), .Z(n11257) );
  AND U10999 ( .A(n11263), .B(n11264), .Z(n11262) );
  XNOR U11000 ( .A(p_input[2789]), .B(n11261), .Z(n11264) );
  XOR U11001 ( .A(n11261), .B(p_input[2757]), .Z(n11263) );
  XOR U11002 ( .A(n11265), .B(n11266), .Z(n11261) );
  AND U11003 ( .A(n11267), .B(n11268), .Z(n11266) );
  XNOR U11004 ( .A(p_input[2788]), .B(n11265), .Z(n11268) );
  XOR U11005 ( .A(n11265), .B(p_input[2756]), .Z(n11267) );
  XOR U11006 ( .A(n11269), .B(n11270), .Z(n11265) );
  AND U11007 ( .A(n11271), .B(n11272), .Z(n11270) );
  XNOR U11008 ( .A(p_input[2787]), .B(n11269), .Z(n11272) );
  XOR U11009 ( .A(n11269), .B(p_input[2755]), .Z(n11271) );
  XOR U11010 ( .A(n11273), .B(n11274), .Z(n11269) );
  AND U11011 ( .A(n11275), .B(n11276), .Z(n11274) );
  XNOR U11012 ( .A(p_input[2786]), .B(n11273), .Z(n11276) );
  XOR U11013 ( .A(n11273), .B(p_input[2754]), .Z(n11275) );
  XNOR U11014 ( .A(n11277), .B(n11278), .Z(n11273) );
  AND U11015 ( .A(n11279), .B(n11280), .Z(n11278) );
  XOR U11016 ( .A(p_input[2785]), .B(n11277), .Z(n11280) );
  XNOR U11017 ( .A(p_input[2753]), .B(n11277), .Z(n11279) );
  AND U11018 ( .A(p_input[2784]), .B(n11281), .Z(n11277) );
  IV U11019 ( .A(p_input[2752]), .Z(n11281) );
  XNOR U11020 ( .A(p_input[2688]), .B(n11282), .Z(n10875) );
  AND U11021 ( .A(n252), .B(n11283), .Z(n11282) );
  XOR U11022 ( .A(p_input[2720]), .B(p_input[2688]), .Z(n11283) );
  XOR U11023 ( .A(n11284), .B(n11285), .Z(n252) );
  AND U11024 ( .A(n11286), .B(n11287), .Z(n11285) );
  XNOR U11025 ( .A(p_input[2751]), .B(n11284), .Z(n11287) );
  XOR U11026 ( .A(n11284), .B(p_input[2719]), .Z(n11286) );
  XOR U11027 ( .A(n11288), .B(n11289), .Z(n11284) );
  AND U11028 ( .A(n11290), .B(n11291), .Z(n11289) );
  XNOR U11029 ( .A(p_input[2750]), .B(n11288), .Z(n11291) );
  XNOR U11030 ( .A(n11288), .B(n10890), .Z(n11290) );
  IV U11031 ( .A(p_input[2718]), .Z(n10890) );
  XOR U11032 ( .A(n11292), .B(n11293), .Z(n11288) );
  AND U11033 ( .A(n11294), .B(n11295), .Z(n11293) );
  XNOR U11034 ( .A(p_input[2749]), .B(n11292), .Z(n11295) );
  XNOR U11035 ( .A(n11292), .B(n10899), .Z(n11294) );
  IV U11036 ( .A(p_input[2717]), .Z(n10899) );
  XOR U11037 ( .A(n11296), .B(n11297), .Z(n11292) );
  AND U11038 ( .A(n11298), .B(n11299), .Z(n11297) );
  XNOR U11039 ( .A(p_input[2748]), .B(n11296), .Z(n11299) );
  XNOR U11040 ( .A(n11296), .B(n10908), .Z(n11298) );
  IV U11041 ( .A(p_input[2716]), .Z(n10908) );
  XOR U11042 ( .A(n11300), .B(n11301), .Z(n11296) );
  AND U11043 ( .A(n11302), .B(n11303), .Z(n11301) );
  XNOR U11044 ( .A(p_input[2747]), .B(n11300), .Z(n11303) );
  XNOR U11045 ( .A(n11300), .B(n10917), .Z(n11302) );
  IV U11046 ( .A(p_input[2715]), .Z(n10917) );
  XOR U11047 ( .A(n11304), .B(n11305), .Z(n11300) );
  AND U11048 ( .A(n11306), .B(n11307), .Z(n11305) );
  XNOR U11049 ( .A(p_input[2746]), .B(n11304), .Z(n11307) );
  XNOR U11050 ( .A(n11304), .B(n10926), .Z(n11306) );
  IV U11051 ( .A(p_input[2714]), .Z(n10926) );
  XOR U11052 ( .A(n11308), .B(n11309), .Z(n11304) );
  AND U11053 ( .A(n11310), .B(n11311), .Z(n11309) );
  XNOR U11054 ( .A(p_input[2745]), .B(n11308), .Z(n11311) );
  XNOR U11055 ( .A(n11308), .B(n10935), .Z(n11310) );
  IV U11056 ( .A(p_input[2713]), .Z(n10935) );
  XOR U11057 ( .A(n11312), .B(n11313), .Z(n11308) );
  AND U11058 ( .A(n11314), .B(n11315), .Z(n11313) );
  XNOR U11059 ( .A(p_input[2744]), .B(n11312), .Z(n11315) );
  XNOR U11060 ( .A(n11312), .B(n10944), .Z(n11314) );
  IV U11061 ( .A(p_input[2712]), .Z(n10944) );
  XOR U11062 ( .A(n11316), .B(n11317), .Z(n11312) );
  AND U11063 ( .A(n11318), .B(n11319), .Z(n11317) );
  XNOR U11064 ( .A(p_input[2743]), .B(n11316), .Z(n11319) );
  XNOR U11065 ( .A(n11316), .B(n10953), .Z(n11318) );
  IV U11066 ( .A(p_input[2711]), .Z(n10953) );
  XOR U11067 ( .A(n11320), .B(n11321), .Z(n11316) );
  AND U11068 ( .A(n11322), .B(n11323), .Z(n11321) );
  XNOR U11069 ( .A(p_input[2742]), .B(n11320), .Z(n11323) );
  XNOR U11070 ( .A(n11320), .B(n10962), .Z(n11322) );
  IV U11071 ( .A(p_input[2710]), .Z(n10962) );
  XOR U11072 ( .A(n11324), .B(n11325), .Z(n11320) );
  AND U11073 ( .A(n11326), .B(n11327), .Z(n11325) );
  XNOR U11074 ( .A(p_input[2741]), .B(n11324), .Z(n11327) );
  XNOR U11075 ( .A(n11324), .B(n10971), .Z(n11326) );
  IV U11076 ( .A(p_input[2709]), .Z(n10971) );
  XOR U11077 ( .A(n11328), .B(n11329), .Z(n11324) );
  AND U11078 ( .A(n11330), .B(n11331), .Z(n11329) );
  XNOR U11079 ( .A(p_input[2740]), .B(n11328), .Z(n11331) );
  XNOR U11080 ( .A(n11328), .B(n10980), .Z(n11330) );
  IV U11081 ( .A(p_input[2708]), .Z(n10980) );
  XOR U11082 ( .A(n11332), .B(n11333), .Z(n11328) );
  AND U11083 ( .A(n11334), .B(n11335), .Z(n11333) );
  XNOR U11084 ( .A(p_input[2739]), .B(n11332), .Z(n11335) );
  XNOR U11085 ( .A(n11332), .B(n10989), .Z(n11334) );
  IV U11086 ( .A(p_input[2707]), .Z(n10989) );
  XOR U11087 ( .A(n11336), .B(n11337), .Z(n11332) );
  AND U11088 ( .A(n11338), .B(n11339), .Z(n11337) );
  XNOR U11089 ( .A(p_input[2738]), .B(n11336), .Z(n11339) );
  XNOR U11090 ( .A(n11336), .B(n10998), .Z(n11338) );
  IV U11091 ( .A(p_input[2706]), .Z(n10998) );
  XOR U11092 ( .A(n11340), .B(n11341), .Z(n11336) );
  AND U11093 ( .A(n11342), .B(n11343), .Z(n11341) );
  XNOR U11094 ( .A(p_input[2737]), .B(n11340), .Z(n11343) );
  XNOR U11095 ( .A(n11340), .B(n11007), .Z(n11342) );
  IV U11096 ( .A(p_input[2705]), .Z(n11007) );
  XOR U11097 ( .A(n11344), .B(n11345), .Z(n11340) );
  AND U11098 ( .A(n11346), .B(n11347), .Z(n11345) );
  XNOR U11099 ( .A(p_input[2736]), .B(n11344), .Z(n11347) );
  XNOR U11100 ( .A(n11344), .B(n11016), .Z(n11346) );
  IV U11101 ( .A(p_input[2704]), .Z(n11016) );
  XOR U11102 ( .A(n11348), .B(n11349), .Z(n11344) );
  AND U11103 ( .A(n11350), .B(n11351), .Z(n11349) );
  XNOR U11104 ( .A(p_input[2735]), .B(n11348), .Z(n11351) );
  XNOR U11105 ( .A(n11348), .B(n11025), .Z(n11350) );
  IV U11106 ( .A(p_input[2703]), .Z(n11025) );
  XOR U11107 ( .A(n11352), .B(n11353), .Z(n11348) );
  AND U11108 ( .A(n11354), .B(n11355), .Z(n11353) );
  XNOR U11109 ( .A(p_input[2734]), .B(n11352), .Z(n11355) );
  XNOR U11110 ( .A(n11352), .B(n11034), .Z(n11354) );
  IV U11111 ( .A(p_input[2702]), .Z(n11034) );
  XOR U11112 ( .A(n11356), .B(n11357), .Z(n11352) );
  AND U11113 ( .A(n11358), .B(n11359), .Z(n11357) );
  XNOR U11114 ( .A(p_input[2733]), .B(n11356), .Z(n11359) );
  XNOR U11115 ( .A(n11356), .B(n11043), .Z(n11358) );
  IV U11116 ( .A(p_input[2701]), .Z(n11043) );
  XOR U11117 ( .A(n11360), .B(n11361), .Z(n11356) );
  AND U11118 ( .A(n11362), .B(n11363), .Z(n11361) );
  XNOR U11119 ( .A(p_input[2732]), .B(n11360), .Z(n11363) );
  XNOR U11120 ( .A(n11360), .B(n11052), .Z(n11362) );
  IV U11121 ( .A(p_input[2700]), .Z(n11052) );
  XOR U11122 ( .A(n11364), .B(n11365), .Z(n11360) );
  AND U11123 ( .A(n11366), .B(n11367), .Z(n11365) );
  XNOR U11124 ( .A(p_input[2731]), .B(n11364), .Z(n11367) );
  XNOR U11125 ( .A(n11364), .B(n11061), .Z(n11366) );
  IV U11126 ( .A(p_input[2699]), .Z(n11061) );
  XOR U11127 ( .A(n11368), .B(n11369), .Z(n11364) );
  AND U11128 ( .A(n11370), .B(n11371), .Z(n11369) );
  XNOR U11129 ( .A(p_input[2730]), .B(n11368), .Z(n11371) );
  XNOR U11130 ( .A(n11368), .B(n11070), .Z(n11370) );
  IV U11131 ( .A(p_input[2698]), .Z(n11070) );
  XOR U11132 ( .A(n11372), .B(n11373), .Z(n11368) );
  AND U11133 ( .A(n11374), .B(n11375), .Z(n11373) );
  XNOR U11134 ( .A(p_input[2729]), .B(n11372), .Z(n11375) );
  XNOR U11135 ( .A(n11372), .B(n11079), .Z(n11374) );
  IV U11136 ( .A(p_input[2697]), .Z(n11079) );
  XOR U11137 ( .A(n11376), .B(n11377), .Z(n11372) );
  AND U11138 ( .A(n11378), .B(n11379), .Z(n11377) );
  XNOR U11139 ( .A(p_input[2728]), .B(n11376), .Z(n11379) );
  XNOR U11140 ( .A(n11376), .B(n11088), .Z(n11378) );
  IV U11141 ( .A(p_input[2696]), .Z(n11088) );
  XOR U11142 ( .A(n11380), .B(n11381), .Z(n11376) );
  AND U11143 ( .A(n11382), .B(n11383), .Z(n11381) );
  XNOR U11144 ( .A(p_input[2727]), .B(n11380), .Z(n11383) );
  XNOR U11145 ( .A(n11380), .B(n11097), .Z(n11382) );
  IV U11146 ( .A(p_input[2695]), .Z(n11097) );
  XOR U11147 ( .A(n11384), .B(n11385), .Z(n11380) );
  AND U11148 ( .A(n11386), .B(n11387), .Z(n11385) );
  XNOR U11149 ( .A(p_input[2726]), .B(n11384), .Z(n11387) );
  XNOR U11150 ( .A(n11384), .B(n11106), .Z(n11386) );
  IV U11151 ( .A(p_input[2694]), .Z(n11106) );
  XOR U11152 ( .A(n11388), .B(n11389), .Z(n11384) );
  AND U11153 ( .A(n11390), .B(n11391), .Z(n11389) );
  XNOR U11154 ( .A(p_input[2725]), .B(n11388), .Z(n11391) );
  XNOR U11155 ( .A(n11388), .B(n11115), .Z(n11390) );
  IV U11156 ( .A(p_input[2693]), .Z(n11115) );
  XOR U11157 ( .A(n11392), .B(n11393), .Z(n11388) );
  AND U11158 ( .A(n11394), .B(n11395), .Z(n11393) );
  XNOR U11159 ( .A(p_input[2724]), .B(n11392), .Z(n11395) );
  XNOR U11160 ( .A(n11392), .B(n11124), .Z(n11394) );
  IV U11161 ( .A(p_input[2692]), .Z(n11124) );
  XOR U11162 ( .A(n11396), .B(n11397), .Z(n11392) );
  AND U11163 ( .A(n11398), .B(n11399), .Z(n11397) );
  XNOR U11164 ( .A(p_input[2723]), .B(n11396), .Z(n11399) );
  XNOR U11165 ( .A(n11396), .B(n11133), .Z(n11398) );
  IV U11166 ( .A(p_input[2691]), .Z(n11133) );
  XOR U11167 ( .A(n11400), .B(n11401), .Z(n11396) );
  AND U11168 ( .A(n11402), .B(n11403), .Z(n11401) );
  XNOR U11169 ( .A(p_input[2722]), .B(n11400), .Z(n11403) );
  XNOR U11170 ( .A(n11400), .B(n11142), .Z(n11402) );
  IV U11171 ( .A(p_input[2690]), .Z(n11142) );
  XNOR U11172 ( .A(n11404), .B(n11405), .Z(n11400) );
  AND U11173 ( .A(n11406), .B(n11407), .Z(n11405) );
  XOR U11174 ( .A(p_input[2721]), .B(n11404), .Z(n11407) );
  XNOR U11175 ( .A(p_input[2689]), .B(n11404), .Z(n11406) );
  AND U11176 ( .A(p_input[2720]), .B(n11408), .Z(n11404) );
  IV U11177 ( .A(p_input[2688]), .Z(n11408) );
  XOR U11178 ( .A(n11409), .B(n11410), .Z(n10498) );
  AND U11179 ( .A(n335), .B(n11411), .Z(n11410) );
  XNOR U11180 ( .A(n11412), .B(n11409), .Z(n11411) );
  XOR U11181 ( .A(n11413), .B(n11414), .Z(n335) );
  AND U11182 ( .A(n11415), .B(n11416), .Z(n11414) );
  XNOR U11183 ( .A(n10513), .B(n11413), .Z(n11416) );
  AND U11184 ( .A(p_input[2687]), .B(p_input[2655]), .Z(n10513) );
  XNOR U11185 ( .A(n11413), .B(n10510), .Z(n11415) );
  IV U11186 ( .A(n11417), .Z(n10510) );
  AND U11187 ( .A(p_input[2591]), .B(p_input[2623]), .Z(n11417) );
  XOR U11188 ( .A(n11418), .B(n11419), .Z(n11413) );
  AND U11189 ( .A(n11420), .B(n11421), .Z(n11419) );
  XOR U11190 ( .A(n11418), .B(n10525), .Z(n11421) );
  XNOR U11191 ( .A(p_input[2654]), .B(n11422), .Z(n10525) );
  AND U11192 ( .A(n258), .B(n11423), .Z(n11422) );
  XOR U11193 ( .A(p_input[2686]), .B(p_input[2654]), .Z(n11423) );
  XNOR U11194 ( .A(n10522), .B(n11418), .Z(n11420) );
  XOR U11195 ( .A(n11424), .B(n11425), .Z(n10522) );
  AND U11196 ( .A(n255), .B(n11426), .Z(n11425) );
  XOR U11197 ( .A(p_input[2622]), .B(p_input[2590]), .Z(n11426) );
  XOR U11198 ( .A(n11427), .B(n11428), .Z(n11418) );
  AND U11199 ( .A(n11429), .B(n11430), .Z(n11428) );
  XOR U11200 ( .A(n11427), .B(n10537), .Z(n11430) );
  XNOR U11201 ( .A(p_input[2653]), .B(n11431), .Z(n10537) );
  AND U11202 ( .A(n258), .B(n11432), .Z(n11431) );
  XOR U11203 ( .A(p_input[2685]), .B(p_input[2653]), .Z(n11432) );
  XNOR U11204 ( .A(n10534), .B(n11427), .Z(n11429) );
  XOR U11205 ( .A(n11433), .B(n11434), .Z(n10534) );
  AND U11206 ( .A(n255), .B(n11435), .Z(n11434) );
  XOR U11207 ( .A(p_input[2621]), .B(p_input[2589]), .Z(n11435) );
  XOR U11208 ( .A(n11436), .B(n11437), .Z(n11427) );
  AND U11209 ( .A(n11438), .B(n11439), .Z(n11437) );
  XOR U11210 ( .A(n11436), .B(n10549), .Z(n11439) );
  XNOR U11211 ( .A(p_input[2652]), .B(n11440), .Z(n10549) );
  AND U11212 ( .A(n258), .B(n11441), .Z(n11440) );
  XOR U11213 ( .A(p_input[2684]), .B(p_input[2652]), .Z(n11441) );
  XNOR U11214 ( .A(n10546), .B(n11436), .Z(n11438) );
  XOR U11215 ( .A(n11442), .B(n11443), .Z(n10546) );
  AND U11216 ( .A(n255), .B(n11444), .Z(n11443) );
  XOR U11217 ( .A(p_input[2620]), .B(p_input[2588]), .Z(n11444) );
  XOR U11218 ( .A(n11445), .B(n11446), .Z(n11436) );
  AND U11219 ( .A(n11447), .B(n11448), .Z(n11446) );
  XOR U11220 ( .A(n11445), .B(n10561), .Z(n11448) );
  XNOR U11221 ( .A(p_input[2651]), .B(n11449), .Z(n10561) );
  AND U11222 ( .A(n258), .B(n11450), .Z(n11449) );
  XOR U11223 ( .A(p_input[2683]), .B(p_input[2651]), .Z(n11450) );
  XNOR U11224 ( .A(n10558), .B(n11445), .Z(n11447) );
  XOR U11225 ( .A(n11451), .B(n11452), .Z(n10558) );
  AND U11226 ( .A(n255), .B(n11453), .Z(n11452) );
  XOR U11227 ( .A(p_input[2619]), .B(p_input[2587]), .Z(n11453) );
  XOR U11228 ( .A(n11454), .B(n11455), .Z(n11445) );
  AND U11229 ( .A(n11456), .B(n11457), .Z(n11455) );
  XOR U11230 ( .A(n11454), .B(n10573), .Z(n11457) );
  XNOR U11231 ( .A(p_input[2650]), .B(n11458), .Z(n10573) );
  AND U11232 ( .A(n258), .B(n11459), .Z(n11458) );
  XOR U11233 ( .A(p_input[2682]), .B(p_input[2650]), .Z(n11459) );
  XNOR U11234 ( .A(n10570), .B(n11454), .Z(n11456) );
  XOR U11235 ( .A(n11460), .B(n11461), .Z(n10570) );
  AND U11236 ( .A(n255), .B(n11462), .Z(n11461) );
  XOR U11237 ( .A(p_input[2618]), .B(p_input[2586]), .Z(n11462) );
  XOR U11238 ( .A(n11463), .B(n11464), .Z(n11454) );
  AND U11239 ( .A(n11465), .B(n11466), .Z(n11464) );
  XOR U11240 ( .A(n11463), .B(n10585), .Z(n11466) );
  XNOR U11241 ( .A(p_input[2649]), .B(n11467), .Z(n10585) );
  AND U11242 ( .A(n258), .B(n11468), .Z(n11467) );
  XOR U11243 ( .A(p_input[2681]), .B(p_input[2649]), .Z(n11468) );
  XNOR U11244 ( .A(n10582), .B(n11463), .Z(n11465) );
  XOR U11245 ( .A(n11469), .B(n11470), .Z(n10582) );
  AND U11246 ( .A(n255), .B(n11471), .Z(n11470) );
  XOR U11247 ( .A(p_input[2617]), .B(p_input[2585]), .Z(n11471) );
  XOR U11248 ( .A(n11472), .B(n11473), .Z(n11463) );
  AND U11249 ( .A(n11474), .B(n11475), .Z(n11473) );
  XOR U11250 ( .A(n11472), .B(n10597), .Z(n11475) );
  XNOR U11251 ( .A(p_input[2648]), .B(n11476), .Z(n10597) );
  AND U11252 ( .A(n258), .B(n11477), .Z(n11476) );
  XOR U11253 ( .A(p_input[2680]), .B(p_input[2648]), .Z(n11477) );
  XNOR U11254 ( .A(n10594), .B(n11472), .Z(n11474) );
  XOR U11255 ( .A(n11478), .B(n11479), .Z(n10594) );
  AND U11256 ( .A(n255), .B(n11480), .Z(n11479) );
  XOR U11257 ( .A(p_input[2616]), .B(p_input[2584]), .Z(n11480) );
  XOR U11258 ( .A(n11481), .B(n11482), .Z(n11472) );
  AND U11259 ( .A(n11483), .B(n11484), .Z(n11482) );
  XOR U11260 ( .A(n11481), .B(n10609), .Z(n11484) );
  XNOR U11261 ( .A(p_input[2647]), .B(n11485), .Z(n10609) );
  AND U11262 ( .A(n258), .B(n11486), .Z(n11485) );
  XOR U11263 ( .A(p_input[2679]), .B(p_input[2647]), .Z(n11486) );
  XNOR U11264 ( .A(n10606), .B(n11481), .Z(n11483) );
  XOR U11265 ( .A(n11487), .B(n11488), .Z(n10606) );
  AND U11266 ( .A(n255), .B(n11489), .Z(n11488) );
  XOR U11267 ( .A(p_input[2615]), .B(p_input[2583]), .Z(n11489) );
  XOR U11268 ( .A(n11490), .B(n11491), .Z(n11481) );
  AND U11269 ( .A(n11492), .B(n11493), .Z(n11491) );
  XOR U11270 ( .A(n11490), .B(n10621), .Z(n11493) );
  XNOR U11271 ( .A(p_input[2646]), .B(n11494), .Z(n10621) );
  AND U11272 ( .A(n258), .B(n11495), .Z(n11494) );
  XOR U11273 ( .A(p_input[2678]), .B(p_input[2646]), .Z(n11495) );
  XNOR U11274 ( .A(n10618), .B(n11490), .Z(n11492) );
  XOR U11275 ( .A(n11496), .B(n11497), .Z(n10618) );
  AND U11276 ( .A(n255), .B(n11498), .Z(n11497) );
  XOR U11277 ( .A(p_input[2614]), .B(p_input[2582]), .Z(n11498) );
  XOR U11278 ( .A(n11499), .B(n11500), .Z(n11490) );
  AND U11279 ( .A(n11501), .B(n11502), .Z(n11500) );
  XOR U11280 ( .A(n11499), .B(n10633), .Z(n11502) );
  XNOR U11281 ( .A(p_input[2645]), .B(n11503), .Z(n10633) );
  AND U11282 ( .A(n258), .B(n11504), .Z(n11503) );
  XOR U11283 ( .A(p_input[2677]), .B(p_input[2645]), .Z(n11504) );
  XNOR U11284 ( .A(n10630), .B(n11499), .Z(n11501) );
  XOR U11285 ( .A(n11505), .B(n11506), .Z(n10630) );
  AND U11286 ( .A(n255), .B(n11507), .Z(n11506) );
  XOR U11287 ( .A(p_input[2613]), .B(p_input[2581]), .Z(n11507) );
  XOR U11288 ( .A(n11508), .B(n11509), .Z(n11499) );
  AND U11289 ( .A(n11510), .B(n11511), .Z(n11509) );
  XOR U11290 ( .A(n11508), .B(n10645), .Z(n11511) );
  XNOR U11291 ( .A(p_input[2644]), .B(n11512), .Z(n10645) );
  AND U11292 ( .A(n258), .B(n11513), .Z(n11512) );
  XOR U11293 ( .A(p_input[2676]), .B(p_input[2644]), .Z(n11513) );
  XNOR U11294 ( .A(n10642), .B(n11508), .Z(n11510) );
  XOR U11295 ( .A(n11514), .B(n11515), .Z(n10642) );
  AND U11296 ( .A(n255), .B(n11516), .Z(n11515) );
  XOR U11297 ( .A(p_input[2612]), .B(p_input[2580]), .Z(n11516) );
  XOR U11298 ( .A(n11517), .B(n11518), .Z(n11508) );
  AND U11299 ( .A(n11519), .B(n11520), .Z(n11518) );
  XOR U11300 ( .A(n11517), .B(n10657), .Z(n11520) );
  XNOR U11301 ( .A(p_input[2643]), .B(n11521), .Z(n10657) );
  AND U11302 ( .A(n258), .B(n11522), .Z(n11521) );
  XOR U11303 ( .A(p_input[2675]), .B(p_input[2643]), .Z(n11522) );
  XNOR U11304 ( .A(n10654), .B(n11517), .Z(n11519) );
  XOR U11305 ( .A(n11523), .B(n11524), .Z(n10654) );
  AND U11306 ( .A(n255), .B(n11525), .Z(n11524) );
  XOR U11307 ( .A(p_input[2611]), .B(p_input[2579]), .Z(n11525) );
  XOR U11308 ( .A(n11526), .B(n11527), .Z(n11517) );
  AND U11309 ( .A(n11528), .B(n11529), .Z(n11527) );
  XOR U11310 ( .A(n11526), .B(n10669), .Z(n11529) );
  XNOR U11311 ( .A(p_input[2642]), .B(n11530), .Z(n10669) );
  AND U11312 ( .A(n258), .B(n11531), .Z(n11530) );
  XOR U11313 ( .A(p_input[2674]), .B(p_input[2642]), .Z(n11531) );
  XNOR U11314 ( .A(n10666), .B(n11526), .Z(n11528) );
  XOR U11315 ( .A(n11532), .B(n11533), .Z(n10666) );
  AND U11316 ( .A(n255), .B(n11534), .Z(n11533) );
  XOR U11317 ( .A(p_input[2610]), .B(p_input[2578]), .Z(n11534) );
  XOR U11318 ( .A(n11535), .B(n11536), .Z(n11526) );
  AND U11319 ( .A(n11537), .B(n11538), .Z(n11536) );
  XOR U11320 ( .A(n11535), .B(n10681), .Z(n11538) );
  XNOR U11321 ( .A(p_input[2641]), .B(n11539), .Z(n10681) );
  AND U11322 ( .A(n258), .B(n11540), .Z(n11539) );
  XOR U11323 ( .A(p_input[2673]), .B(p_input[2641]), .Z(n11540) );
  XNOR U11324 ( .A(n10678), .B(n11535), .Z(n11537) );
  XOR U11325 ( .A(n11541), .B(n11542), .Z(n10678) );
  AND U11326 ( .A(n255), .B(n11543), .Z(n11542) );
  XOR U11327 ( .A(p_input[2609]), .B(p_input[2577]), .Z(n11543) );
  XOR U11328 ( .A(n11544), .B(n11545), .Z(n11535) );
  AND U11329 ( .A(n11546), .B(n11547), .Z(n11545) );
  XOR U11330 ( .A(n11544), .B(n10693), .Z(n11547) );
  XNOR U11331 ( .A(p_input[2640]), .B(n11548), .Z(n10693) );
  AND U11332 ( .A(n258), .B(n11549), .Z(n11548) );
  XOR U11333 ( .A(p_input[2672]), .B(p_input[2640]), .Z(n11549) );
  XNOR U11334 ( .A(n10690), .B(n11544), .Z(n11546) );
  XOR U11335 ( .A(n11550), .B(n11551), .Z(n10690) );
  AND U11336 ( .A(n255), .B(n11552), .Z(n11551) );
  XOR U11337 ( .A(p_input[2608]), .B(p_input[2576]), .Z(n11552) );
  XOR U11338 ( .A(n11553), .B(n11554), .Z(n11544) );
  AND U11339 ( .A(n11555), .B(n11556), .Z(n11554) );
  XOR U11340 ( .A(n11553), .B(n10705), .Z(n11556) );
  XNOR U11341 ( .A(p_input[2639]), .B(n11557), .Z(n10705) );
  AND U11342 ( .A(n258), .B(n11558), .Z(n11557) );
  XOR U11343 ( .A(p_input[2671]), .B(p_input[2639]), .Z(n11558) );
  XNOR U11344 ( .A(n10702), .B(n11553), .Z(n11555) );
  XOR U11345 ( .A(n11559), .B(n11560), .Z(n10702) );
  AND U11346 ( .A(n255), .B(n11561), .Z(n11560) );
  XOR U11347 ( .A(p_input[2607]), .B(p_input[2575]), .Z(n11561) );
  XOR U11348 ( .A(n11562), .B(n11563), .Z(n11553) );
  AND U11349 ( .A(n11564), .B(n11565), .Z(n11563) );
  XOR U11350 ( .A(n11562), .B(n10717), .Z(n11565) );
  XNOR U11351 ( .A(p_input[2638]), .B(n11566), .Z(n10717) );
  AND U11352 ( .A(n258), .B(n11567), .Z(n11566) );
  XOR U11353 ( .A(p_input[2670]), .B(p_input[2638]), .Z(n11567) );
  XNOR U11354 ( .A(n10714), .B(n11562), .Z(n11564) );
  XOR U11355 ( .A(n11568), .B(n11569), .Z(n10714) );
  AND U11356 ( .A(n255), .B(n11570), .Z(n11569) );
  XOR U11357 ( .A(p_input[2606]), .B(p_input[2574]), .Z(n11570) );
  XOR U11358 ( .A(n11571), .B(n11572), .Z(n11562) );
  AND U11359 ( .A(n11573), .B(n11574), .Z(n11572) );
  XOR U11360 ( .A(n11571), .B(n10729), .Z(n11574) );
  XNOR U11361 ( .A(p_input[2637]), .B(n11575), .Z(n10729) );
  AND U11362 ( .A(n258), .B(n11576), .Z(n11575) );
  XOR U11363 ( .A(p_input[2669]), .B(p_input[2637]), .Z(n11576) );
  XNOR U11364 ( .A(n10726), .B(n11571), .Z(n11573) );
  XOR U11365 ( .A(n11577), .B(n11578), .Z(n10726) );
  AND U11366 ( .A(n255), .B(n11579), .Z(n11578) );
  XOR U11367 ( .A(p_input[2605]), .B(p_input[2573]), .Z(n11579) );
  XOR U11368 ( .A(n11580), .B(n11581), .Z(n11571) );
  AND U11369 ( .A(n11582), .B(n11583), .Z(n11581) );
  XOR U11370 ( .A(n11580), .B(n10741), .Z(n11583) );
  XNOR U11371 ( .A(p_input[2636]), .B(n11584), .Z(n10741) );
  AND U11372 ( .A(n258), .B(n11585), .Z(n11584) );
  XOR U11373 ( .A(p_input[2668]), .B(p_input[2636]), .Z(n11585) );
  XNOR U11374 ( .A(n10738), .B(n11580), .Z(n11582) );
  XOR U11375 ( .A(n11586), .B(n11587), .Z(n10738) );
  AND U11376 ( .A(n255), .B(n11588), .Z(n11587) );
  XOR U11377 ( .A(p_input[2604]), .B(p_input[2572]), .Z(n11588) );
  XOR U11378 ( .A(n11589), .B(n11590), .Z(n11580) );
  AND U11379 ( .A(n11591), .B(n11592), .Z(n11590) );
  XOR U11380 ( .A(n11589), .B(n10753), .Z(n11592) );
  XNOR U11381 ( .A(p_input[2635]), .B(n11593), .Z(n10753) );
  AND U11382 ( .A(n258), .B(n11594), .Z(n11593) );
  XOR U11383 ( .A(p_input[2667]), .B(p_input[2635]), .Z(n11594) );
  XNOR U11384 ( .A(n10750), .B(n11589), .Z(n11591) );
  XOR U11385 ( .A(n11595), .B(n11596), .Z(n10750) );
  AND U11386 ( .A(n255), .B(n11597), .Z(n11596) );
  XOR U11387 ( .A(p_input[2603]), .B(p_input[2571]), .Z(n11597) );
  XOR U11388 ( .A(n11598), .B(n11599), .Z(n11589) );
  AND U11389 ( .A(n11600), .B(n11601), .Z(n11599) );
  XOR U11390 ( .A(n11598), .B(n10765), .Z(n11601) );
  XNOR U11391 ( .A(p_input[2634]), .B(n11602), .Z(n10765) );
  AND U11392 ( .A(n258), .B(n11603), .Z(n11602) );
  XOR U11393 ( .A(p_input[2666]), .B(p_input[2634]), .Z(n11603) );
  XNOR U11394 ( .A(n10762), .B(n11598), .Z(n11600) );
  XOR U11395 ( .A(n11604), .B(n11605), .Z(n10762) );
  AND U11396 ( .A(n255), .B(n11606), .Z(n11605) );
  XOR U11397 ( .A(p_input[2602]), .B(p_input[2570]), .Z(n11606) );
  XOR U11398 ( .A(n11607), .B(n11608), .Z(n11598) );
  AND U11399 ( .A(n11609), .B(n11610), .Z(n11608) );
  XOR U11400 ( .A(n11607), .B(n10777), .Z(n11610) );
  XNOR U11401 ( .A(p_input[2633]), .B(n11611), .Z(n10777) );
  AND U11402 ( .A(n258), .B(n11612), .Z(n11611) );
  XOR U11403 ( .A(p_input[2665]), .B(p_input[2633]), .Z(n11612) );
  XNOR U11404 ( .A(n10774), .B(n11607), .Z(n11609) );
  XOR U11405 ( .A(n11613), .B(n11614), .Z(n10774) );
  AND U11406 ( .A(n255), .B(n11615), .Z(n11614) );
  XOR U11407 ( .A(p_input[2601]), .B(p_input[2569]), .Z(n11615) );
  XOR U11408 ( .A(n11616), .B(n11617), .Z(n11607) );
  AND U11409 ( .A(n11618), .B(n11619), .Z(n11617) );
  XOR U11410 ( .A(n11616), .B(n10789), .Z(n11619) );
  XNOR U11411 ( .A(p_input[2632]), .B(n11620), .Z(n10789) );
  AND U11412 ( .A(n258), .B(n11621), .Z(n11620) );
  XOR U11413 ( .A(p_input[2664]), .B(p_input[2632]), .Z(n11621) );
  XNOR U11414 ( .A(n10786), .B(n11616), .Z(n11618) );
  XOR U11415 ( .A(n11622), .B(n11623), .Z(n10786) );
  AND U11416 ( .A(n255), .B(n11624), .Z(n11623) );
  XOR U11417 ( .A(p_input[2600]), .B(p_input[2568]), .Z(n11624) );
  XOR U11418 ( .A(n11625), .B(n11626), .Z(n11616) );
  AND U11419 ( .A(n11627), .B(n11628), .Z(n11626) );
  XOR U11420 ( .A(n11625), .B(n10801), .Z(n11628) );
  XNOR U11421 ( .A(p_input[2631]), .B(n11629), .Z(n10801) );
  AND U11422 ( .A(n258), .B(n11630), .Z(n11629) );
  XOR U11423 ( .A(p_input[2663]), .B(p_input[2631]), .Z(n11630) );
  XNOR U11424 ( .A(n10798), .B(n11625), .Z(n11627) );
  XOR U11425 ( .A(n11631), .B(n11632), .Z(n10798) );
  AND U11426 ( .A(n255), .B(n11633), .Z(n11632) );
  XOR U11427 ( .A(p_input[2599]), .B(p_input[2567]), .Z(n11633) );
  XOR U11428 ( .A(n11634), .B(n11635), .Z(n11625) );
  AND U11429 ( .A(n11636), .B(n11637), .Z(n11635) );
  XOR U11430 ( .A(n11634), .B(n10813), .Z(n11637) );
  XNOR U11431 ( .A(p_input[2630]), .B(n11638), .Z(n10813) );
  AND U11432 ( .A(n258), .B(n11639), .Z(n11638) );
  XOR U11433 ( .A(p_input[2662]), .B(p_input[2630]), .Z(n11639) );
  XNOR U11434 ( .A(n10810), .B(n11634), .Z(n11636) );
  XOR U11435 ( .A(n11640), .B(n11641), .Z(n10810) );
  AND U11436 ( .A(n255), .B(n11642), .Z(n11641) );
  XOR U11437 ( .A(p_input[2598]), .B(p_input[2566]), .Z(n11642) );
  XOR U11438 ( .A(n11643), .B(n11644), .Z(n11634) );
  AND U11439 ( .A(n11645), .B(n11646), .Z(n11644) );
  XOR U11440 ( .A(n11643), .B(n10825), .Z(n11646) );
  XNOR U11441 ( .A(p_input[2629]), .B(n11647), .Z(n10825) );
  AND U11442 ( .A(n258), .B(n11648), .Z(n11647) );
  XOR U11443 ( .A(p_input[2661]), .B(p_input[2629]), .Z(n11648) );
  XNOR U11444 ( .A(n10822), .B(n11643), .Z(n11645) );
  XOR U11445 ( .A(n11649), .B(n11650), .Z(n10822) );
  AND U11446 ( .A(n255), .B(n11651), .Z(n11650) );
  XOR U11447 ( .A(p_input[2597]), .B(p_input[2565]), .Z(n11651) );
  XOR U11448 ( .A(n11652), .B(n11653), .Z(n11643) );
  AND U11449 ( .A(n11654), .B(n11655), .Z(n11653) );
  XOR U11450 ( .A(n11652), .B(n10837), .Z(n11655) );
  XNOR U11451 ( .A(p_input[2628]), .B(n11656), .Z(n10837) );
  AND U11452 ( .A(n258), .B(n11657), .Z(n11656) );
  XOR U11453 ( .A(p_input[2660]), .B(p_input[2628]), .Z(n11657) );
  XNOR U11454 ( .A(n10834), .B(n11652), .Z(n11654) );
  XOR U11455 ( .A(n11658), .B(n11659), .Z(n10834) );
  AND U11456 ( .A(n255), .B(n11660), .Z(n11659) );
  XOR U11457 ( .A(p_input[2596]), .B(p_input[2564]), .Z(n11660) );
  XOR U11458 ( .A(n11661), .B(n11662), .Z(n11652) );
  AND U11459 ( .A(n11663), .B(n11664), .Z(n11662) );
  XOR U11460 ( .A(n11661), .B(n10849), .Z(n11664) );
  XNOR U11461 ( .A(p_input[2627]), .B(n11665), .Z(n10849) );
  AND U11462 ( .A(n258), .B(n11666), .Z(n11665) );
  XOR U11463 ( .A(p_input[2659]), .B(p_input[2627]), .Z(n11666) );
  XNOR U11464 ( .A(n10846), .B(n11661), .Z(n11663) );
  XOR U11465 ( .A(n11667), .B(n11668), .Z(n10846) );
  AND U11466 ( .A(n255), .B(n11669), .Z(n11668) );
  XOR U11467 ( .A(p_input[2595]), .B(p_input[2563]), .Z(n11669) );
  XOR U11468 ( .A(n11670), .B(n11671), .Z(n11661) );
  AND U11469 ( .A(n11672), .B(n11673), .Z(n11671) );
  XOR U11470 ( .A(n10861), .B(n11670), .Z(n11673) );
  XNOR U11471 ( .A(p_input[2626]), .B(n11674), .Z(n10861) );
  AND U11472 ( .A(n258), .B(n11675), .Z(n11674) );
  XOR U11473 ( .A(p_input[2658]), .B(p_input[2626]), .Z(n11675) );
  XNOR U11474 ( .A(n11670), .B(n10858), .Z(n11672) );
  XOR U11475 ( .A(n11676), .B(n11677), .Z(n10858) );
  AND U11476 ( .A(n255), .B(n11678), .Z(n11677) );
  XOR U11477 ( .A(p_input[2594]), .B(p_input[2562]), .Z(n11678) );
  XOR U11478 ( .A(n11679), .B(n11680), .Z(n11670) );
  AND U11479 ( .A(n11681), .B(n11682), .Z(n11680) );
  XNOR U11480 ( .A(n11683), .B(n10874), .Z(n11682) );
  XNOR U11481 ( .A(p_input[2625]), .B(n11684), .Z(n10874) );
  AND U11482 ( .A(n258), .B(n11685), .Z(n11684) );
  XNOR U11483 ( .A(p_input[2657]), .B(n11686), .Z(n11685) );
  IV U11484 ( .A(p_input[2625]), .Z(n11686) );
  XNOR U11485 ( .A(n10871), .B(n11679), .Z(n11681) );
  XNOR U11486 ( .A(p_input[2561]), .B(n11687), .Z(n10871) );
  AND U11487 ( .A(n255), .B(n11688), .Z(n11687) );
  XOR U11488 ( .A(p_input[2593]), .B(p_input[2561]), .Z(n11688) );
  IV U11489 ( .A(n11683), .Z(n11679) );
  AND U11490 ( .A(n11409), .B(n11412), .Z(n11683) );
  XOR U11491 ( .A(p_input[2624]), .B(n11689), .Z(n11412) );
  AND U11492 ( .A(n258), .B(n11690), .Z(n11689) );
  XOR U11493 ( .A(p_input[2656]), .B(p_input[2624]), .Z(n11690) );
  XOR U11494 ( .A(n11691), .B(n11692), .Z(n258) );
  AND U11495 ( .A(n11693), .B(n11694), .Z(n11692) );
  XNOR U11496 ( .A(p_input[2687]), .B(n11691), .Z(n11694) );
  XOR U11497 ( .A(n11691), .B(p_input[2655]), .Z(n11693) );
  XOR U11498 ( .A(n11695), .B(n11696), .Z(n11691) );
  AND U11499 ( .A(n11697), .B(n11698), .Z(n11696) );
  XNOR U11500 ( .A(p_input[2686]), .B(n11695), .Z(n11698) );
  XOR U11501 ( .A(n11695), .B(p_input[2654]), .Z(n11697) );
  XOR U11502 ( .A(n11699), .B(n11700), .Z(n11695) );
  AND U11503 ( .A(n11701), .B(n11702), .Z(n11700) );
  XNOR U11504 ( .A(p_input[2685]), .B(n11699), .Z(n11702) );
  XOR U11505 ( .A(n11699), .B(p_input[2653]), .Z(n11701) );
  XOR U11506 ( .A(n11703), .B(n11704), .Z(n11699) );
  AND U11507 ( .A(n11705), .B(n11706), .Z(n11704) );
  XNOR U11508 ( .A(p_input[2684]), .B(n11703), .Z(n11706) );
  XOR U11509 ( .A(n11703), .B(p_input[2652]), .Z(n11705) );
  XOR U11510 ( .A(n11707), .B(n11708), .Z(n11703) );
  AND U11511 ( .A(n11709), .B(n11710), .Z(n11708) );
  XNOR U11512 ( .A(p_input[2683]), .B(n11707), .Z(n11710) );
  XOR U11513 ( .A(n11707), .B(p_input[2651]), .Z(n11709) );
  XOR U11514 ( .A(n11711), .B(n11712), .Z(n11707) );
  AND U11515 ( .A(n11713), .B(n11714), .Z(n11712) );
  XNOR U11516 ( .A(p_input[2682]), .B(n11711), .Z(n11714) );
  XOR U11517 ( .A(n11711), .B(p_input[2650]), .Z(n11713) );
  XOR U11518 ( .A(n11715), .B(n11716), .Z(n11711) );
  AND U11519 ( .A(n11717), .B(n11718), .Z(n11716) );
  XNOR U11520 ( .A(p_input[2681]), .B(n11715), .Z(n11718) );
  XOR U11521 ( .A(n11715), .B(p_input[2649]), .Z(n11717) );
  XOR U11522 ( .A(n11719), .B(n11720), .Z(n11715) );
  AND U11523 ( .A(n11721), .B(n11722), .Z(n11720) );
  XNOR U11524 ( .A(p_input[2680]), .B(n11719), .Z(n11722) );
  XOR U11525 ( .A(n11719), .B(p_input[2648]), .Z(n11721) );
  XOR U11526 ( .A(n11723), .B(n11724), .Z(n11719) );
  AND U11527 ( .A(n11725), .B(n11726), .Z(n11724) );
  XNOR U11528 ( .A(p_input[2679]), .B(n11723), .Z(n11726) );
  XOR U11529 ( .A(n11723), .B(p_input[2647]), .Z(n11725) );
  XOR U11530 ( .A(n11727), .B(n11728), .Z(n11723) );
  AND U11531 ( .A(n11729), .B(n11730), .Z(n11728) );
  XNOR U11532 ( .A(p_input[2678]), .B(n11727), .Z(n11730) );
  XOR U11533 ( .A(n11727), .B(p_input[2646]), .Z(n11729) );
  XOR U11534 ( .A(n11731), .B(n11732), .Z(n11727) );
  AND U11535 ( .A(n11733), .B(n11734), .Z(n11732) );
  XNOR U11536 ( .A(p_input[2677]), .B(n11731), .Z(n11734) );
  XOR U11537 ( .A(n11731), .B(p_input[2645]), .Z(n11733) );
  XOR U11538 ( .A(n11735), .B(n11736), .Z(n11731) );
  AND U11539 ( .A(n11737), .B(n11738), .Z(n11736) );
  XNOR U11540 ( .A(p_input[2676]), .B(n11735), .Z(n11738) );
  XOR U11541 ( .A(n11735), .B(p_input[2644]), .Z(n11737) );
  XOR U11542 ( .A(n11739), .B(n11740), .Z(n11735) );
  AND U11543 ( .A(n11741), .B(n11742), .Z(n11740) );
  XNOR U11544 ( .A(p_input[2675]), .B(n11739), .Z(n11742) );
  XOR U11545 ( .A(n11739), .B(p_input[2643]), .Z(n11741) );
  XOR U11546 ( .A(n11743), .B(n11744), .Z(n11739) );
  AND U11547 ( .A(n11745), .B(n11746), .Z(n11744) );
  XNOR U11548 ( .A(p_input[2674]), .B(n11743), .Z(n11746) );
  XOR U11549 ( .A(n11743), .B(p_input[2642]), .Z(n11745) );
  XOR U11550 ( .A(n11747), .B(n11748), .Z(n11743) );
  AND U11551 ( .A(n11749), .B(n11750), .Z(n11748) );
  XNOR U11552 ( .A(p_input[2673]), .B(n11747), .Z(n11750) );
  XOR U11553 ( .A(n11747), .B(p_input[2641]), .Z(n11749) );
  XOR U11554 ( .A(n11751), .B(n11752), .Z(n11747) );
  AND U11555 ( .A(n11753), .B(n11754), .Z(n11752) );
  XNOR U11556 ( .A(p_input[2672]), .B(n11751), .Z(n11754) );
  XOR U11557 ( .A(n11751), .B(p_input[2640]), .Z(n11753) );
  XOR U11558 ( .A(n11755), .B(n11756), .Z(n11751) );
  AND U11559 ( .A(n11757), .B(n11758), .Z(n11756) );
  XNOR U11560 ( .A(p_input[2671]), .B(n11755), .Z(n11758) );
  XOR U11561 ( .A(n11755), .B(p_input[2639]), .Z(n11757) );
  XOR U11562 ( .A(n11759), .B(n11760), .Z(n11755) );
  AND U11563 ( .A(n11761), .B(n11762), .Z(n11760) );
  XNOR U11564 ( .A(p_input[2670]), .B(n11759), .Z(n11762) );
  XOR U11565 ( .A(n11759), .B(p_input[2638]), .Z(n11761) );
  XOR U11566 ( .A(n11763), .B(n11764), .Z(n11759) );
  AND U11567 ( .A(n11765), .B(n11766), .Z(n11764) );
  XNOR U11568 ( .A(p_input[2669]), .B(n11763), .Z(n11766) );
  XOR U11569 ( .A(n11763), .B(p_input[2637]), .Z(n11765) );
  XOR U11570 ( .A(n11767), .B(n11768), .Z(n11763) );
  AND U11571 ( .A(n11769), .B(n11770), .Z(n11768) );
  XNOR U11572 ( .A(p_input[2668]), .B(n11767), .Z(n11770) );
  XOR U11573 ( .A(n11767), .B(p_input[2636]), .Z(n11769) );
  XOR U11574 ( .A(n11771), .B(n11772), .Z(n11767) );
  AND U11575 ( .A(n11773), .B(n11774), .Z(n11772) );
  XNOR U11576 ( .A(p_input[2667]), .B(n11771), .Z(n11774) );
  XOR U11577 ( .A(n11771), .B(p_input[2635]), .Z(n11773) );
  XOR U11578 ( .A(n11775), .B(n11776), .Z(n11771) );
  AND U11579 ( .A(n11777), .B(n11778), .Z(n11776) );
  XNOR U11580 ( .A(p_input[2666]), .B(n11775), .Z(n11778) );
  XOR U11581 ( .A(n11775), .B(p_input[2634]), .Z(n11777) );
  XOR U11582 ( .A(n11779), .B(n11780), .Z(n11775) );
  AND U11583 ( .A(n11781), .B(n11782), .Z(n11780) );
  XNOR U11584 ( .A(p_input[2665]), .B(n11779), .Z(n11782) );
  XOR U11585 ( .A(n11779), .B(p_input[2633]), .Z(n11781) );
  XOR U11586 ( .A(n11783), .B(n11784), .Z(n11779) );
  AND U11587 ( .A(n11785), .B(n11786), .Z(n11784) );
  XNOR U11588 ( .A(p_input[2664]), .B(n11783), .Z(n11786) );
  XOR U11589 ( .A(n11783), .B(p_input[2632]), .Z(n11785) );
  XOR U11590 ( .A(n11787), .B(n11788), .Z(n11783) );
  AND U11591 ( .A(n11789), .B(n11790), .Z(n11788) );
  XNOR U11592 ( .A(p_input[2663]), .B(n11787), .Z(n11790) );
  XOR U11593 ( .A(n11787), .B(p_input[2631]), .Z(n11789) );
  XOR U11594 ( .A(n11791), .B(n11792), .Z(n11787) );
  AND U11595 ( .A(n11793), .B(n11794), .Z(n11792) );
  XNOR U11596 ( .A(p_input[2662]), .B(n11791), .Z(n11794) );
  XOR U11597 ( .A(n11791), .B(p_input[2630]), .Z(n11793) );
  XOR U11598 ( .A(n11795), .B(n11796), .Z(n11791) );
  AND U11599 ( .A(n11797), .B(n11798), .Z(n11796) );
  XNOR U11600 ( .A(p_input[2661]), .B(n11795), .Z(n11798) );
  XOR U11601 ( .A(n11795), .B(p_input[2629]), .Z(n11797) );
  XOR U11602 ( .A(n11799), .B(n11800), .Z(n11795) );
  AND U11603 ( .A(n11801), .B(n11802), .Z(n11800) );
  XNOR U11604 ( .A(p_input[2660]), .B(n11799), .Z(n11802) );
  XOR U11605 ( .A(n11799), .B(p_input[2628]), .Z(n11801) );
  XOR U11606 ( .A(n11803), .B(n11804), .Z(n11799) );
  AND U11607 ( .A(n11805), .B(n11806), .Z(n11804) );
  XNOR U11608 ( .A(p_input[2659]), .B(n11803), .Z(n11806) );
  XOR U11609 ( .A(n11803), .B(p_input[2627]), .Z(n11805) );
  XOR U11610 ( .A(n11807), .B(n11808), .Z(n11803) );
  AND U11611 ( .A(n11809), .B(n11810), .Z(n11808) );
  XNOR U11612 ( .A(p_input[2658]), .B(n11807), .Z(n11810) );
  XOR U11613 ( .A(n11807), .B(p_input[2626]), .Z(n11809) );
  XNOR U11614 ( .A(n11811), .B(n11812), .Z(n11807) );
  AND U11615 ( .A(n11813), .B(n11814), .Z(n11812) );
  XOR U11616 ( .A(p_input[2657]), .B(n11811), .Z(n11814) );
  XNOR U11617 ( .A(p_input[2625]), .B(n11811), .Z(n11813) );
  AND U11618 ( .A(p_input[2656]), .B(n11815), .Z(n11811) );
  IV U11619 ( .A(p_input[2624]), .Z(n11815) );
  XNOR U11620 ( .A(p_input[2560]), .B(n11816), .Z(n11409) );
  AND U11621 ( .A(n255), .B(n11817), .Z(n11816) );
  XOR U11622 ( .A(p_input[2592]), .B(p_input[2560]), .Z(n11817) );
  XOR U11623 ( .A(n11818), .B(n11819), .Z(n255) );
  AND U11624 ( .A(n11820), .B(n11821), .Z(n11819) );
  XNOR U11625 ( .A(p_input[2623]), .B(n11818), .Z(n11821) );
  XOR U11626 ( .A(n11818), .B(p_input[2591]), .Z(n11820) );
  XOR U11627 ( .A(n11822), .B(n11823), .Z(n11818) );
  AND U11628 ( .A(n11824), .B(n11825), .Z(n11823) );
  XNOR U11629 ( .A(p_input[2622]), .B(n11822), .Z(n11825) );
  XNOR U11630 ( .A(n11822), .B(n11424), .Z(n11824) );
  IV U11631 ( .A(p_input[2590]), .Z(n11424) );
  XOR U11632 ( .A(n11826), .B(n11827), .Z(n11822) );
  AND U11633 ( .A(n11828), .B(n11829), .Z(n11827) );
  XNOR U11634 ( .A(p_input[2621]), .B(n11826), .Z(n11829) );
  XNOR U11635 ( .A(n11826), .B(n11433), .Z(n11828) );
  IV U11636 ( .A(p_input[2589]), .Z(n11433) );
  XOR U11637 ( .A(n11830), .B(n11831), .Z(n11826) );
  AND U11638 ( .A(n11832), .B(n11833), .Z(n11831) );
  XNOR U11639 ( .A(p_input[2620]), .B(n11830), .Z(n11833) );
  XNOR U11640 ( .A(n11830), .B(n11442), .Z(n11832) );
  IV U11641 ( .A(p_input[2588]), .Z(n11442) );
  XOR U11642 ( .A(n11834), .B(n11835), .Z(n11830) );
  AND U11643 ( .A(n11836), .B(n11837), .Z(n11835) );
  XNOR U11644 ( .A(p_input[2619]), .B(n11834), .Z(n11837) );
  XNOR U11645 ( .A(n11834), .B(n11451), .Z(n11836) );
  IV U11646 ( .A(p_input[2587]), .Z(n11451) );
  XOR U11647 ( .A(n11838), .B(n11839), .Z(n11834) );
  AND U11648 ( .A(n11840), .B(n11841), .Z(n11839) );
  XNOR U11649 ( .A(p_input[2618]), .B(n11838), .Z(n11841) );
  XNOR U11650 ( .A(n11838), .B(n11460), .Z(n11840) );
  IV U11651 ( .A(p_input[2586]), .Z(n11460) );
  XOR U11652 ( .A(n11842), .B(n11843), .Z(n11838) );
  AND U11653 ( .A(n11844), .B(n11845), .Z(n11843) );
  XNOR U11654 ( .A(p_input[2617]), .B(n11842), .Z(n11845) );
  XNOR U11655 ( .A(n11842), .B(n11469), .Z(n11844) );
  IV U11656 ( .A(p_input[2585]), .Z(n11469) );
  XOR U11657 ( .A(n11846), .B(n11847), .Z(n11842) );
  AND U11658 ( .A(n11848), .B(n11849), .Z(n11847) );
  XNOR U11659 ( .A(p_input[2616]), .B(n11846), .Z(n11849) );
  XNOR U11660 ( .A(n11846), .B(n11478), .Z(n11848) );
  IV U11661 ( .A(p_input[2584]), .Z(n11478) );
  XOR U11662 ( .A(n11850), .B(n11851), .Z(n11846) );
  AND U11663 ( .A(n11852), .B(n11853), .Z(n11851) );
  XNOR U11664 ( .A(p_input[2615]), .B(n11850), .Z(n11853) );
  XNOR U11665 ( .A(n11850), .B(n11487), .Z(n11852) );
  IV U11666 ( .A(p_input[2583]), .Z(n11487) );
  XOR U11667 ( .A(n11854), .B(n11855), .Z(n11850) );
  AND U11668 ( .A(n11856), .B(n11857), .Z(n11855) );
  XNOR U11669 ( .A(p_input[2614]), .B(n11854), .Z(n11857) );
  XNOR U11670 ( .A(n11854), .B(n11496), .Z(n11856) );
  IV U11671 ( .A(p_input[2582]), .Z(n11496) );
  XOR U11672 ( .A(n11858), .B(n11859), .Z(n11854) );
  AND U11673 ( .A(n11860), .B(n11861), .Z(n11859) );
  XNOR U11674 ( .A(p_input[2613]), .B(n11858), .Z(n11861) );
  XNOR U11675 ( .A(n11858), .B(n11505), .Z(n11860) );
  IV U11676 ( .A(p_input[2581]), .Z(n11505) );
  XOR U11677 ( .A(n11862), .B(n11863), .Z(n11858) );
  AND U11678 ( .A(n11864), .B(n11865), .Z(n11863) );
  XNOR U11679 ( .A(p_input[2612]), .B(n11862), .Z(n11865) );
  XNOR U11680 ( .A(n11862), .B(n11514), .Z(n11864) );
  IV U11681 ( .A(p_input[2580]), .Z(n11514) );
  XOR U11682 ( .A(n11866), .B(n11867), .Z(n11862) );
  AND U11683 ( .A(n11868), .B(n11869), .Z(n11867) );
  XNOR U11684 ( .A(p_input[2611]), .B(n11866), .Z(n11869) );
  XNOR U11685 ( .A(n11866), .B(n11523), .Z(n11868) );
  IV U11686 ( .A(p_input[2579]), .Z(n11523) );
  XOR U11687 ( .A(n11870), .B(n11871), .Z(n11866) );
  AND U11688 ( .A(n11872), .B(n11873), .Z(n11871) );
  XNOR U11689 ( .A(p_input[2610]), .B(n11870), .Z(n11873) );
  XNOR U11690 ( .A(n11870), .B(n11532), .Z(n11872) );
  IV U11691 ( .A(p_input[2578]), .Z(n11532) );
  XOR U11692 ( .A(n11874), .B(n11875), .Z(n11870) );
  AND U11693 ( .A(n11876), .B(n11877), .Z(n11875) );
  XNOR U11694 ( .A(p_input[2609]), .B(n11874), .Z(n11877) );
  XNOR U11695 ( .A(n11874), .B(n11541), .Z(n11876) );
  IV U11696 ( .A(p_input[2577]), .Z(n11541) );
  XOR U11697 ( .A(n11878), .B(n11879), .Z(n11874) );
  AND U11698 ( .A(n11880), .B(n11881), .Z(n11879) );
  XNOR U11699 ( .A(p_input[2608]), .B(n11878), .Z(n11881) );
  XNOR U11700 ( .A(n11878), .B(n11550), .Z(n11880) );
  IV U11701 ( .A(p_input[2576]), .Z(n11550) );
  XOR U11702 ( .A(n11882), .B(n11883), .Z(n11878) );
  AND U11703 ( .A(n11884), .B(n11885), .Z(n11883) );
  XNOR U11704 ( .A(p_input[2607]), .B(n11882), .Z(n11885) );
  XNOR U11705 ( .A(n11882), .B(n11559), .Z(n11884) );
  IV U11706 ( .A(p_input[2575]), .Z(n11559) );
  XOR U11707 ( .A(n11886), .B(n11887), .Z(n11882) );
  AND U11708 ( .A(n11888), .B(n11889), .Z(n11887) );
  XNOR U11709 ( .A(p_input[2606]), .B(n11886), .Z(n11889) );
  XNOR U11710 ( .A(n11886), .B(n11568), .Z(n11888) );
  IV U11711 ( .A(p_input[2574]), .Z(n11568) );
  XOR U11712 ( .A(n11890), .B(n11891), .Z(n11886) );
  AND U11713 ( .A(n11892), .B(n11893), .Z(n11891) );
  XNOR U11714 ( .A(p_input[2605]), .B(n11890), .Z(n11893) );
  XNOR U11715 ( .A(n11890), .B(n11577), .Z(n11892) );
  IV U11716 ( .A(p_input[2573]), .Z(n11577) );
  XOR U11717 ( .A(n11894), .B(n11895), .Z(n11890) );
  AND U11718 ( .A(n11896), .B(n11897), .Z(n11895) );
  XNOR U11719 ( .A(p_input[2604]), .B(n11894), .Z(n11897) );
  XNOR U11720 ( .A(n11894), .B(n11586), .Z(n11896) );
  IV U11721 ( .A(p_input[2572]), .Z(n11586) );
  XOR U11722 ( .A(n11898), .B(n11899), .Z(n11894) );
  AND U11723 ( .A(n11900), .B(n11901), .Z(n11899) );
  XNOR U11724 ( .A(p_input[2603]), .B(n11898), .Z(n11901) );
  XNOR U11725 ( .A(n11898), .B(n11595), .Z(n11900) );
  IV U11726 ( .A(p_input[2571]), .Z(n11595) );
  XOR U11727 ( .A(n11902), .B(n11903), .Z(n11898) );
  AND U11728 ( .A(n11904), .B(n11905), .Z(n11903) );
  XNOR U11729 ( .A(p_input[2602]), .B(n11902), .Z(n11905) );
  XNOR U11730 ( .A(n11902), .B(n11604), .Z(n11904) );
  IV U11731 ( .A(p_input[2570]), .Z(n11604) );
  XOR U11732 ( .A(n11906), .B(n11907), .Z(n11902) );
  AND U11733 ( .A(n11908), .B(n11909), .Z(n11907) );
  XNOR U11734 ( .A(p_input[2601]), .B(n11906), .Z(n11909) );
  XNOR U11735 ( .A(n11906), .B(n11613), .Z(n11908) );
  IV U11736 ( .A(p_input[2569]), .Z(n11613) );
  XOR U11737 ( .A(n11910), .B(n11911), .Z(n11906) );
  AND U11738 ( .A(n11912), .B(n11913), .Z(n11911) );
  XNOR U11739 ( .A(p_input[2600]), .B(n11910), .Z(n11913) );
  XNOR U11740 ( .A(n11910), .B(n11622), .Z(n11912) );
  IV U11741 ( .A(p_input[2568]), .Z(n11622) );
  XOR U11742 ( .A(n11914), .B(n11915), .Z(n11910) );
  AND U11743 ( .A(n11916), .B(n11917), .Z(n11915) );
  XNOR U11744 ( .A(p_input[2599]), .B(n11914), .Z(n11917) );
  XNOR U11745 ( .A(n11914), .B(n11631), .Z(n11916) );
  IV U11746 ( .A(p_input[2567]), .Z(n11631) );
  XOR U11747 ( .A(n11918), .B(n11919), .Z(n11914) );
  AND U11748 ( .A(n11920), .B(n11921), .Z(n11919) );
  XNOR U11749 ( .A(p_input[2598]), .B(n11918), .Z(n11921) );
  XNOR U11750 ( .A(n11918), .B(n11640), .Z(n11920) );
  IV U11751 ( .A(p_input[2566]), .Z(n11640) );
  XOR U11752 ( .A(n11922), .B(n11923), .Z(n11918) );
  AND U11753 ( .A(n11924), .B(n11925), .Z(n11923) );
  XNOR U11754 ( .A(p_input[2597]), .B(n11922), .Z(n11925) );
  XNOR U11755 ( .A(n11922), .B(n11649), .Z(n11924) );
  IV U11756 ( .A(p_input[2565]), .Z(n11649) );
  XOR U11757 ( .A(n11926), .B(n11927), .Z(n11922) );
  AND U11758 ( .A(n11928), .B(n11929), .Z(n11927) );
  XNOR U11759 ( .A(p_input[2596]), .B(n11926), .Z(n11929) );
  XNOR U11760 ( .A(n11926), .B(n11658), .Z(n11928) );
  IV U11761 ( .A(p_input[2564]), .Z(n11658) );
  XOR U11762 ( .A(n11930), .B(n11931), .Z(n11926) );
  AND U11763 ( .A(n11932), .B(n11933), .Z(n11931) );
  XNOR U11764 ( .A(p_input[2595]), .B(n11930), .Z(n11933) );
  XNOR U11765 ( .A(n11930), .B(n11667), .Z(n11932) );
  IV U11766 ( .A(p_input[2563]), .Z(n11667) );
  XOR U11767 ( .A(n11934), .B(n11935), .Z(n11930) );
  AND U11768 ( .A(n11936), .B(n11937), .Z(n11935) );
  XNOR U11769 ( .A(p_input[2594]), .B(n11934), .Z(n11937) );
  XNOR U11770 ( .A(n11934), .B(n11676), .Z(n11936) );
  IV U11771 ( .A(p_input[2562]), .Z(n11676) );
  XNOR U11772 ( .A(n11938), .B(n11939), .Z(n11934) );
  AND U11773 ( .A(n11940), .B(n11941), .Z(n11939) );
  XOR U11774 ( .A(p_input[2593]), .B(n11938), .Z(n11941) );
  XNOR U11775 ( .A(p_input[2561]), .B(n11938), .Z(n11940) );
  AND U11776 ( .A(p_input[2592]), .B(n11942), .Z(n11938) );
  IV U11777 ( .A(p_input[2560]), .Z(n11942) );
  XOR U11778 ( .A(n11943), .B(n11944), .Z(n8299) );
  AND U11779 ( .A(n579), .B(n11945), .Z(n11944) );
  XNOR U11780 ( .A(n11946), .B(n11943), .Z(n11945) );
  XOR U11781 ( .A(n11947), .B(n11948), .Z(n579) );
  AND U11782 ( .A(n11949), .B(n11950), .Z(n11948) );
  XOR U11783 ( .A(n11947), .B(n8314), .Z(n11950) );
  XOR U11784 ( .A(n11951), .B(n11952), .Z(n8314) );
  AND U11785 ( .A(n506), .B(n11953), .Z(n11952) );
  XOR U11786 ( .A(n11954), .B(n11951), .Z(n11953) );
  XNOR U11787 ( .A(n8311), .B(n11947), .Z(n11949) );
  XOR U11788 ( .A(n11955), .B(n11956), .Z(n8311) );
  AND U11789 ( .A(n503), .B(n11957), .Z(n11956) );
  XOR U11790 ( .A(n11958), .B(n11955), .Z(n11957) );
  XOR U11791 ( .A(n11959), .B(n11960), .Z(n11947) );
  AND U11792 ( .A(n11961), .B(n11962), .Z(n11960) );
  XOR U11793 ( .A(n11959), .B(n8326), .Z(n11962) );
  XOR U11794 ( .A(n11963), .B(n11964), .Z(n8326) );
  AND U11795 ( .A(n506), .B(n11965), .Z(n11964) );
  XOR U11796 ( .A(n11966), .B(n11963), .Z(n11965) );
  XNOR U11797 ( .A(n8323), .B(n11959), .Z(n11961) );
  XOR U11798 ( .A(n11967), .B(n11968), .Z(n8323) );
  AND U11799 ( .A(n503), .B(n11969), .Z(n11968) );
  XOR U11800 ( .A(n11970), .B(n11967), .Z(n11969) );
  XOR U11801 ( .A(n11971), .B(n11972), .Z(n11959) );
  AND U11802 ( .A(n11973), .B(n11974), .Z(n11972) );
  XOR U11803 ( .A(n11971), .B(n8338), .Z(n11974) );
  XOR U11804 ( .A(n11975), .B(n11976), .Z(n8338) );
  AND U11805 ( .A(n506), .B(n11977), .Z(n11976) );
  XOR U11806 ( .A(n11978), .B(n11975), .Z(n11977) );
  XNOR U11807 ( .A(n8335), .B(n11971), .Z(n11973) );
  XOR U11808 ( .A(n11979), .B(n11980), .Z(n8335) );
  AND U11809 ( .A(n503), .B(n11981), .Z(n11980) );
  XOR U11810 ( .A(n11982), .B(n11979), .Z(n11981) );
  XOR U11811 ( .A(n11983), .B(n11984), .Z(n11971) );
  AND U11812 ( .A(n11985), .B(n11986), .Z(n11984) );
  XOR U11813 ( .A(n11983), .B(n8350), .Z(n11986) );
  XOR U11814 ( .A(n11987), .B(n11988), .Z(n8350) );
  AND U11815 ( .A(n506), .B(n11989), .Z(n11988) );
  XOR U11816 ( .A(n11990), .B(n11987), .Z(n11989) );
  XNOR U11817 ( .A(n8347), .B(n11983), .Z(n11985) );
  XOR U11818 ( .A(n11991), .B(n11992), .Z(n8347) );
  AND U11819 ( .A(n503), .B(n11993), .Z(n11992) );
  XOR U11820 ( .A(n11994), .B(n11991), .Z(n11993) );
  XOR U11821 ( .A(n11995), .B(n11996), .Z(n11983) );
  AND U11822 ( .A(n11997), .B(n11998), .Z(n11996) );
  XOR U11823 ( .A(n11995), .B(n8362), .Z(n11998) );
  XOR U11824 ( .A(n11999), .B(n12000), .Z(n8362) );
  AND U11825 ( .A(n506), .B(n12001), .Z(n12000) );
  XOR U11826 ( .A(n12002), .B(n11999), .Z(n12001) );
  XNOR U11827 ( .A(n8359), .B(n11995), .Z(n11997) );
  XOR U11828 ( .A(n12003), .B(n12004), .Z(n8359) );
  AND U11829 ( .A(n503), .B(n12005), .Z(n12004) );
  XOR U11830 ( .A(n12006), .B(n12003), .Z(n12005) );
  XOR U11831 ( .A(n12007), .B(n12008), .Z(n11995) );
  AND U11832 ( .A(n12009), .B(n12010), .Z(n12008) );
  XOR U11833 ( .A(n12007), .B(n8374), .Z(n12010) );
  XOR U11834 ( .A(n12011), .B(n12012), .Z(n8374) );
  AND U11835 ( .A(n506), .B(n12013), .Z(n12012) );
  XOR U11836 ( .A(n12014), .B(n12011), .Z(n12013) );
  XNOR U11837 ( .A(n8371), .B(n12007), .Z(n12009) );
  XOR U11838 ( .A(n12015), .B(n12016), .Z(n8371) );
  AND U11839 ( .A(n503), .B(n12017), .Z(n12016) );
  XOR U11840 ( .A(n12018), .B(n12015), .Z(n12017) );
  XOR U11841 ( .A(n12019), .B(n12020), .Z(n12007) );
  AND U11842 ( .A(n12021), .B(n12022), .Z(n12020) );
  XOR U11843 ( .A(n12019), .B(n8386), .Z(n12022) );
  XOR U11844 ( .A(n12023), .B(n12024), .Z(n8386) );
  AND U11845 ( .A(n506), .B(n12025), .Z(n12024) );
  XOR U11846 ( .A(n12026), .B(n12023), .Z(n12025) );
  XNOR U11847 ( .A(n8383), .B(n12019), .Z(n12021) );
  XOR U11848 ( .A(n12027), .B(n12028), .Z(n8383) );
  AND U11849 ( .A(n503), .B(n12029), .Z(n12028) );
  XOR U11850 ( .A(n12030), .B(n12027), .Z(n12029) );
  XOR U11851 ( .A(n12031), .B(n12032), .Z(n12019) );
  AND U11852 ( .A(n12033), .B(n12034), .Z(n12032) );
  XOR U11853 ( .A(n12031), .B(n8398), .Z(n12034) );
  XOR U11854 ( .A(n12035), .B(n12036), .Z(n8398) );
  AND U11855 ( .A(n506), .B(n12037), .Z(n12036) );
  XOR U11856 ( .A(n12038), .B(n12035), .Z(n12037) );
  XNOR U11857 ( .A(n8395), .B(n12031), .Z(n12033) );
  XOR U11858 ( .A(n12039), .B(n12040), .Z(n8395) );
  AND U11859 ( .A(n503), .B(n12041), .Z(n12040) );
  XOR U11860 ( .A(n12042), .B(n12039), .Z(n12041) );
  XOR U11861 ( .A(n12043), .B(n12044), .Z(n12031) );
  AND U11862 ( .A(n12045), .B(n12046), .Z(n12044) );
  XOR U11863 ( .A(n12043), .B(n8410), .Z(n12046) );
  XOR U11864 ( .A(n12047), .B(n12048), .Z(n8410) );
  AND U11865 ( .A(n506), .B(n12049), .Z(n12048) );
  XOR U11866 ( .A(n12050), .B(n12047), .Z(n12049) );
  XNOR U11867 ( .A(n8407), .B(n12043), .Z(n12045) );
  XOR U11868 ( .A(n12051), .B(n12052), .Z(n8407) );
  AND U11869 ( .A(n503), .B(n12053), .Z(n12052) );
  XOR U11870 ( .A(n12054), .B(n12051), .Z(n12053) );
  XOR U11871 ( .A(n12055), .B(n12056), .Z(n12043) );
  AND U11872 ( .A(n12057), .B(n12058), .Z(n12056) );
  XOR U11873 ( .A(n12055), .B(n8422), .Z(n12058) );
  XOR U11874 ( .A(n12059), .B(n12060), .Z(n8422) );
  AND U11875 ( .A(n506), .B(n12061), .Z(n12060) );
  XOR U11876 ( .A(n12062), .B(n12059), .Z(n12061) );
  XNOR U11877 ( .A(n8419), .B(n12055), .Z(n12057) );
  XOR U11878 ( .A(n12063), .B(n12064), .Z(n8419) );
  AND U11879 ( .A(n503), .B(n12065), .Z(n12064) );
  XOR U11880 ( .A(n12066), .B(n12063), .Z(n12065) );
  XOR U11881 ( .A(n12067), .B(n12068), .Z(n12055) );
  AND U11882 ( .A(n12069), .B(n12070), .Z(n12068) );
  XOR U11883 ( .A(n12067), .B(n8434), .Z(n12070) );
  XOR U11884 ( .A(n12071), .B(n12072), .Z(n8434) );
  AND U11885 ( .A(n506), .B(n12073), .Z(n12072) );
  XOR U11886 ( .A(n12074), .B(n12071), .Z(n12073) );
  XNOR U11887 ( .A(n8431), .B(n12067), .Z(n12069) );
  XOR U11888 ( .A(n12075), .B(n12076), .Z(n8431) );
  AND U11889 ( .A(n503), .B(n12077), .Z(n12076) );
  XOR U11890 ( .A(n12078), .B(n12075), .Z(n12077) );
  XOR U11891 ( .A(n12079), .B(n12080), .Z(n12067) );
  AND U11892 ( .A(n12081), .B(n12082), .Z(n12080) );
  XOR U11893 ( .A(n12079), .B(n8446), .Z(n12082) );
  XOR U11894 ( .A(n12083), .B(n12084), .Z(n8446) );
  AND U11895 ( .A(n506), .B(n12085), .Z(n12084) );
  XOR U11896 ( .A(n12086), .B(n12083), .Z(n12085) );
  XNOR U11897 ( .A(n8443), .B(n12079), .Z(n12081) );
  XOR U11898 ( .A(n12087), .B(n12088), .Z(n8443) );
  AND U11899 ( .A(n503), .B(n12089), .Z(n12088) );
  XOR U11900 ( .A(n12090), .B(n12087), .Z(n12089) );
  XOR U11901 ( .A(n12091), .B(n12092), .Z(n12079) );
  AND U11902 ( .A(n12093), .B(n12094), .Z(n12092) );
  XOR U11903 ( .A(n12091), .B(n8458), .Z(n12094) );
  XOR U11904 ( .A(n12095), .B(n12096), .Z(n8458) );
  AND U11905 ( .A(n506), .B(n12097), .Z(n12096) );
  XOR U11906 ( .A(n12098), .B(n12095), .Z(n12097) );
  XNOR U11907 ( .A(n8455), .B(n12091), .Z(n12093) );
  XOR U11908 ( .A(n12099), .B(n12100), .Z(n8455) );
  AND U11909 ( .A(n503), .B(n12101), .Z(n12100) );
  XOR U11910 ( .A(n12102), .B(n12099), .Z(n12101) );
  XOR U11911 ( .A(n12103), .B(n12104), .Z(n12091) );
  AND U11912 ( .A(n12105), .B(n12106), .Z(n12104) );
  XOR U11913 ( .A(n12103), .B(n8470), .Z(n12106) );
  XOR U11914 ( .A(n12107), .B(n12108), .Z(n8470) );
  AND U11915 ( .A(n506), .B(n12109), .Z(n12108) );
  XOR U11916 ( .A(n12110), .B(n12107), .Z(n12109) );
  XNOR U11917 ( .A(n8467), .B(n12103), .Z(n12105) );
  XOR U11918 ( .A(n12111), .B(n12112), .Z(n8467) );
  AND U11919 ( .A(n503), .B(n12113), .Z(n12112) );
  XOR U11920 ( .A(n12114), .B(n12111), .Z(n12113) );
  XOR U11921 ( .A(n12115), .B(n12116), .Z(n12103) );
  AND U11922 ( .A(n12117), .B(n12118), .Z(n12116) );
  XOR U11923 ( .A(n12115), .B(n8482), .Z(n12118) );
  XOR U11924 ( .A(n12119), .B(n12120), .Z(n8482) );
  AND U11925 ( .A(n506), .B(n12121), .Z(n12120) );
  XOR U11926 ( .A(n12122), .B(n12119), .Z(n12121) );
  XNOR U11927 ( .A(n8479), .B(n12115), .Z(n12117) );
  XOR U11928 ( .A(n12123), .B(n12124), .Z(n8479) );
  AND U11929 ( .A(n503), .B(n12125), .Z(n12124) );
  XOR U11930 ( .A(n12126), .B(n12123), .Z(n12125) );
  XOR U11931 ( .A(n12127), .B(n12128), .Z(n12115) );
  AND U11932 ( .A(n12129), .B(n12130), .Z(n12128) );
  XOR U11933 ( .A(n12127), .B(n8494), .Z(n12130) );
  XOR U11934 ( .A(n12131), .B(n12132), .Z(n8494) );
  AND U11935 ( .A(n506), .B(n12133), .Z(n12132) );
  XOR U11936 ( .A(n12134), .B(n12131), .Z(n12133) );
  XNOR U11937 ( .A(n8491), .B(n12127), .Z(n12129) );
  XOR U11938 ( .A(n12135), .B(n12136), .Z(n8491) );
  AND U11939 ( .A(n503), .B(n12137), .Z(n12136) );
  XOR U11940 ( .A(n12138), .B(n12135), .Z(n12137) );
  XOR U11941 ( .A(n12139), .B(n12140), .Z(n12127) );
  AND U11942 ( .A(n12141), .B(n12142), .Z(n12140) );
  XOR U11943 ( .A(n12139), .B(n8506), .Z(n12142) );
  XOR U11944 ( .A(n12143), .B(n12144), .Z(n8506) );
  AND U11945 ( .A(n506), .B(n12145), .Z(n12144) );
  XOR U11946 ( .A(n12146), .B(n12143), .Z(n12145) );
  XNOR U11947 ( .A(n8503), .B(n12139), .Z(n12141) );
  XOR U11948 ( .A(n12147), .B(n12148), .Z(n8503) );
  AND U11949 ( .A(n503), .B(n12149), .Z(n12148) );
  XOR U11950 ( .A(n12150), .B(n12147), .Z(n12149) );
  XOR U11951 ( .A(n12151), .B(n12152), .Z(n12139) );
  AND U11952 ( .A(n12153), .B(n12154), .Z(n12152) );
  XOR U11953 ( .A(n12151), .B(n8518), .Z(n12154) );
  XOR U11954 ( .A(n12155), .B(n12156), .Z(n8518) );
  AND U11955 ( .A(n506), .B(n12157), .Z(n12156) );
  XOR U11956 ( .A(n12158), .B(n12155), .Z(n12157) );
  XNOR U11957 ( .A(n8515), .B(n12151), .Z(n12153) );
  XOR U11958 ( .A(n12159), .B(n12160), .Z(n8515) );
  AND U11959 ( .A(n503), .B(n12161), .Z(n12160) );
  XOR U11960 ( .A(n12162), .B(n12159), .Z(n12161) );
  XOR U11961 ( .A(n12163), .B(n12164), .Z(n12151) );
  AND U11962 ( .A(n12165), .B(n12166), .Z(n12164) );
  XOR U11963 ( .A(n12163), .B(n8530), .Z(n12166) );
  XOR U11964 ( .A(n12167), .B(n12168), .Z(n8530) );
  AND U11965 ( .A(n506), .B(n12169), .Z(n12168) );
  XOR U11966 ( .A(n12170), .B(n12167), .Z(n12169) );
  XNOR U11967 ( .A(n8527), .B(n12163), .Z(n12165) );
  XOR U11968 ( .A(n12171), .B(n12172), .Z(n8527) );
  AND U11969 ( .A(n503), .B(n12173), .Z(n12172) );
  XOR U11970 ( .A(n12174), .B(n12171), .Z(n12173) );
  XOR U11971 ( .A(n12175), .B(n12176), .Z(n12163) );
  AND U11972 ( .A(n12177), .B(n12178), .Z(n12176) );
  XOR U11973 ( .A(n12175), .B(n8542), .Z(n12178) );
  XOR U11974 ( .A(n12179), .B(n12180), .Z(n8542) );
  AND U11975 ( .A(n506), .B(n12181), .Z(n12180) );
  XOR U11976 ( .A(n12182), .B(n12179), .Z(n12181) );
  XNOR U11977 ( .A(n8539), .B(n12175), .Z(n12177) );
  XOR U11978 ( .A(n12183), .B(n12184), .Z(n8539) );
  AND U11979 ( .A(n503), .B(n12185), .Z(n12184) );
  XOR U11980 ( .A(n12186), .B(n12183), .Z(n12185) );
  XOR U11981 ( .A(n12187), .B(n12188), .Z(n12175) );
  AND U11982 ( .A(n12189), .B(n12190), .Z(n12188) );
  XOR U11983 ( .A(n12187), .B(n8554), .Z(n12190) );
  XOR U11984 ( .A(n12191), .B(n12192), .Z(n8554) );
  AND U11985 ( .A(n506), .B(n12193), .Z(n12192) );
  XOR U11986 ( .A(n12194), .B(n12191), .Z(n12193) );
  XNOR U11987 ( .A(n8551), .B(n12187), .Z(n12189) );
  XOR U11988 ( .A(n12195), .B(n12196), .Z(n8551) );
  AND U11989 ( .A(n503), .B(n12197), .Z(n12196) );
  XOR U11990 ( .A(n12198), .B(n12195), .Z(n12197) );
  XOR U11991 ( .A(n12199), .B(n12200), .Z(n12187) );
  AND U11992 ( .A(n12201), .B(n12202), .Z(n12200) );
  XOR U11993 ( .A(n12199), .B(n8566), .Z(n12202) );
  XOR U11994 ( .A(n12203), .B(n12204), .Z(n8566) );
  AND U11995 ( .A(n506), .B(n12205), .Z(n12204) );
  XOR U11996 ( .A(n12206), .B(n12203), .Z(n12205) );
  XNOR U11997 ( .A(n8563), .B(n12199), .Z(n12201) );
  XOR U11998 ( .A(n12207), .B(n12208), .Z(n8563) );
  AND U11999 ( .A(n503), .B(n12209), .Z(n12208) );
  XOR U12000 ( .A(n12210), .B(n12207), .Z(n12209) );
  XOR U12001 ( .A(n12211), .B(n12212), .Z(n12199) );
  AND U12002 ( .A(n12213), .B(n12214), .Z(n12212) );
  XOR U12003 ( .A(n12211), .B(n8578), .Z(n12214) );
  XOR U12004 ( .A(n12215), .B(n12216), .Z(n8578) );
  AND U12005 ( .A(n506), .B(n12217), .Z(n12216) );
  XOR U12006 ( .A(n12218), .B(n12215), .Z(n12217) );
  XNOR U12007 ( .A(n8575), .B(n12211), .Z(n12213) );
  XOR U12008 ( .A(n12219), .B(n12220), .Z(n8575) );
  AND U12009 ( .A(n503), .B(n12221), .Z(n12220) );
  XOR U12010 ( .A(n12222), .B(n12219), .Z(n12221) );
  XOR U12011 ( .A(n12223), .B(n12224), .Z(n12211) );
  AND U12012 ( .A(n12225), .B(n12226), .Z(n12224) );
  XOR U12013 ( .A(n12223), .B(n8590), .Z(n12226) );
  XOR U12014 ( .A(n12227), .B(n12228), .Z(n8590) );
  AND U12015 ( .A(n506), .B(n12229), .Z(n12228) );
  XOR U12016 ( .A(n12230), .B(n12227), .Z(n12229) );
  XNOR U12017 ( .A(n8587), .B(n12223), .Z(n12225) );
  XOR U12018 ( .A(n12231), .B(n12232), .Z(n8587) );
  AND U12019 ( .A(n503), .B(n12233), .Z(n12232) );
  XOR U12020 ( .A(n12234), .B(n12231), .Z(n12233) );
  XOR U12021 ( .A(n12235), .B(n12236), .Z(n12223) );
  AND U12022 ( .A(n12237), .B(n12238), .Z(n12236) );
  XOR U12023 ( .A(n12235), .B(n8602), .Z(n12238) );
  XOR U12024 ( .A(n12239), .B(n12240), .Z(n8602) );
  AND U12025 ( .A(n506), .B(n12241), .Z(n12240) );
  XOR U12026 ( .A(n12242), .B(n12239), .Z(n12241) );
  XNOR U12027 ( .A(n8599), .B(n12235), .Z(n12237) );
  XOR U12028 ( .A(n12243), .B(n12244), .Z(n8599) );
  AND U12029 ( .A(n503), .B(n12245), .Z(n12244) );
  XOR U12030 ( .A(n12246), .B(n12243), .Z(n12245) );
  XOR U12031 ( .A(n12247), .B(n12248), .Z(n12235) );
  AND U12032 ( .A(n12249), .B(n12250), .Z(n12248) );
  XOR U12033 ( .A(n12247), .B(n8614), .Z(n12250) );
  XOR U12034 ( .A(n12251), .B(n12252), .Z(n8614) );
  AND U12035 ( .A(n506), .B(n12253), .Z(n12252) );
  XOR U12036 ( .A(n12254), .B(n12251), .Z(n12253) );
  XNOR U12037 ( .A(n8611), .B(n12247), .Z(n12249) );
  XOR U12038 ( .A(n12255), .B(n12256), .Z(n8611) );
  AND U12039 ( .A(n503), .B(n12257), .Z(n12256) );
  XOR U12040 ( .A(n12258), .B(n12255), .Z(n12257) );
  XOR U12041 ( .A(n12259), .B(n12260), .Z(n12247) );
  AND U12042 ( .A(n12261), .B(n12262), .Z(n12260) );
  XOR U12043 ( .A(n12259), .B(n8626), .Z(n12262) );
  XOR U12044 ( .A(n12263), .B(n12264), .Z(n8626) );
  AND U12045 ( .A(n506), .B(n12265), .Z(n12264) );
  XOR U12046 ( .A(n12266), .B(n12263), .Z(n12265) );
  XNOR U12047 ( .A(n8623), .B(n12259), .Z(n12261) );
  XOR U12048 ( .A(n12267), .B(n12268), .Z(n8623) );
  AND U12049 ( .A(n503), .B(n12269), .Z(n12268) );
  XOR U12050 ( .A(n12270), .B(n12267), .Z(n12269) );
  XOR U12051 ( .A(n12271), .B(n12272), .Z(n12259) );
  AND U12052 ( .A(n12273), .B(n12274), .Z(n12272) );
  XOR U12053 ( .A(n12271), .B(n8638), .Z(n12274) );
  XOR U12054 ( .A(n12275), .B(n12276), .Z(n8638) );
  AND U12055 ( .A(n506), .B(n12277), .Z(n12276) );
  XOR U12056 ( .A(n12278), .B(n12275), .Z(n12277) );
  XNOR U12057 ( .A(n8635), .B(n12271), .Z(n12273) );
  XOR U12058 ( .A(n12279), .B(n12280), .Z(n8635) );
  AND U12059 ( .A(n503), .B(n12281), .Z(n12280) );
  XOR U12060 ( .A(n12282), .B(n12279), .Z(n12281) );
  XOR U12061 ( .A(n12283), .B(n12284), .Z(n12271) );
  AND U12062 ( .A(n12285), .B(n12286), .Z(n12284) );
  XOR U12063 ( .A(n12283), .B(n8650), .Z(n12286) );
  XOR U12064 ( .A(n12287), .B(n12288), .Z(n8650) );
  AND U12065 ( .A(n506), .B(n12289), .Z(n12288) );
  XOR U12066 ( .A(n12290), .B(n12287), .Z(n12289) );
  XNOR U12067 ( .A(n8647), .B(n12283), .Z(n12285) );
  XOR U12068 ( .A(n12291), .B(n12292), .Z(n8647) );
  AND U12069 ( .A(n503), .B(n12293), .Z(n12292) );
  XOR U12070 ( .A(n12294), .B(n12291), .Z(n12293) );
  XOR U12071 ( .A(n12295), .B(n12296), .Z(n12283) );
  AND U12072 ( .A(n12297), .B(n12298), .Z(n12296) );
  XOR U12073 ( .A(n8662), .B(n12295), .Z(n12298) );
  XOR U12074 ( .A(n12299), .B(n12300), .Z(n8662) );
  AND U12075 ( .A(n506), .B(n12301), .Z(n12300) );
  XOR U12076 ( .A(n12299), .B(n12302), .Z(n12301) );
  XNOR U12077 ( .A(n12295), .B(n8659), .Z(n12297) );
  XOR U12078 ( .A(n12303), .B(n12304), .Z(n8659) );
  AND U12079 ( .A(n503), .B(n12305), .Z(n12304) );
  XOR U12080 ( .A(n12303), .B(n12306), .Z(n12305) );
  XOR U12081 ( .A(n12307), .B(n12308), .Z(n12295) );
  AND U12082 ( .A(n12309), .B(n12310), .Z(n12308) );
  XNOR U12083 ( .A(n12311), .B(n8675), .Z(n12310) );
  XOR U12084 ( .A(n12312), .B(n12313), .Z(n8675) );
  AND U12085 ( .A(n506), .B(n12314), .Z(n12313) );
  XOR U12086 ( .A(n12315), .B(n12312), .Z(n12314) );
  XNOR U12087 ( .A(n8672), .B(n12307), .Z(n12309) );
  XOR U12088 ( .A(n12316), .B(n12317), .Z(n8672) );
  AND U12089 ( .A(n503), .B(n12318), .Z(n12317) );
  XOR U12090 ( .A(n12319), .B(n12316), .Z(n12318) );
  IV U12091 ( .A(n12311), .Z(n12307) );
  AND U12092 ( .A(n11943), .B(n11946), .Z(n12311) );
  XNOR U12093 ( .A(n12320), .B(n12321), .Z(n11946) );
  AND U12094 ( .A(n506), .B(n12322), .Z(n12321) );
  XNOR U12095 ( .A(n12323), .B(n12320), .Z(n12322) );
  XOR U12096 ( .A(n12324), .B(n12325), .Z(n506) );
  AND U12097 ( .A(n12326), .B(n12327), .Z(n12325) );
  XOR U12098 ( .A(n12324), .B(n11954), .Z(n12327) );
  XNOR U12099 ( .A(n12328), .B(n12329), .Z(n11954) );
  AND U12100 ( .A(n12330), .B(n346), .Z(n12329) );
  AND U12101 ( .A(n12328), .B(n12331), .Z(n12330) );
  XNOR U12102 ( .A(n11951), .B(n12324), .Z(n12326) );
  XOR U12103 ( .A(n12332), .B(n12333), .Z(n11951) );
  AND U12104 ( .A(n12334), .B(n344), .Z(n12333) );
  NOR U12105 ( .A(n12332), .B(n12335), .Z(n12334) );
  XOR U12106 ( .A(n12336), .B(n12337), .Z(n12324) );
  AND U12107 ( .A(n12338), .B(n12339), .Z(n12337) );
  XOR U12108 ( .A(n12336), .B(n11966), .Z(n12339) );
  XOR U12109 ( .A(n12340), .B(n12341), .Z(n11966) );
  AND U12110 ( .A(n346), .B(n12342), .Z(n12341) );
  XOR U12111 ( .A(n12343), .B(n12340), .Z(n12342) );
  XNOR U12112 ( .A(n11963), .B(n12336), .Z(n12338) );
  XOR U12113 ( .A(n12344), .B(n12345), .Z(n11963) );
  AND U12114 ( .A(n344), .B(n12346), .Z(n12345) );
  XOR U12115 ( .A(n12347), .B(n12344), .Z(n12346) );
  XOR U12116 ( .A(n12348), .B(n12349), .Z(n12336) );
  AND U12117 ( .A(n12350), .B(n12351), .Z(n12349) );
  XOR U12118 ( .A(n12348), .B(n11978), .Z(n12351) );
  XOR U12119 ( .A(n12352), .B(n12353), .Z(n11978) );
  AND U12120 ( .A(n346), .B(n12354), .Z(n12353) );
  XOR U12121 ( .A(n12355), .B(n12352), .Z(n12354) );
  XNOR U12122 ( .A(n11975), .B(n12348), .Z(n12350) );
  XOR U12123 ( .A(n12356), .B(n12357), .Z(n11975) );
  AND U12124 ( .A(n344), .B(n12358), .Z(n12357) );
  XOR U12125 ( .A(n12359), .B(n12356), .Z(n12358) );
  XOR U12126 ( .A(n12360), .B(n12361), .Z(n12348) );
  AND U12127 ( .A(n12362), .B(n12363), .Z(n12361) );
  XOR U12128 ( .A(n12360), .B(n11990), .Z(n12363) );
  XOR U12129 ( .A(n12364), .B(n12365), .Z(n11990) );
  AND U12130 ( .A(n346), .B(n12366), .Z(n12365) );
  XOR U12131 ( .A(n12367), .B(n12364), .Z(n12366) );
  XNOR U12132 ( .A(n11987), .B(n12360), .Z(n12362) );
  XOR U12133 ( .A(n12368), .B(n12369), .Z(n11987) );
  AND U12134 ( .A(n344), .B(n12370), .Z(n12369) );
  XOR U12135 ( .A(n12371), .B(n12368), .Z(n12370) );
  XOR U12136 ( .A(n12372), .B(n12373), .Z(n12360) );
  AND U12137 ( .A(n12374), .B(n12375), .Z(n12373) );
  XOR U12138 ( .A(n12372), .B(n12002), .Z(n12375) );
  XOR U12139 ( .A(n12376), .B(n12377), .Z(n12002) );
  AND U12140 ( .A(n346), .B(n12378), .Z(n12377) );
  XOR U12141 ( .A(n12379), .B(n12376), .Z(n12378) );
  XNOR U12142 ( .A(n11999), .B(n12372), .Z(n12374) );
  XOR U12143 ( .A(n12380), .B(n12381), .Z(n11999) );
  AND U12144 ( .A(n344), .B(n12382), .Z(n12381) );
  XOR U12145 ( .A(n12383), .B(n12380), .Z(n12382) );
  XOR U12146 ( .A(n12384), .B(n12385), .Z(n12372) );
  AND U12147 ( .A(n12386), .B(n12387), .Z(n12385) );
  XOR U12148 ( .A(n12384), .B(n12014), .Z(n12387) );
  XOR U12149 ( .A(n12388), .B(n12389), .Z(n12014) );
  AND U12150 ( .A(n346), .B(n12390), .Z(n12389) );
  XOR U12151 ( .A(n12391), .B(n12388), .Z(n12390) );
  XNOR U12152 ( .A(n12011), .B(n12384), .Z(n12386) );
  XOR U12153 ( .A(n12392), .B(n12393), .Z(n12011) );
  AND U12154 ( .A(n344), .B(n12394), .Z(n12393) );
  XOR U12155 ( .A(n12395), .B(n12392), .Z(n12394) );
  XOR U12156 ( .A(n12396), .B(n12397), .Z(n12384) );
  AND U12157 ( .A(n12398), .B(n12399), .Z(n12397) );
  XOR U12158 ( .A(n12396), .B(n12026), .Z(n12399) );
  XOR U12159 ( .A(n12400), .B(n12401), .Z(n12026) );
  AND U12160 ( .A(n346), .B(n12402), .Z(n12401) );
  XOR U12161 ( .A(n12403), .B(n12400), .Z(n12402) );
  XNOR U12162 ( .A(n12023), .B(n12396), .Z(n12398) );
  XOR U12163 ( .A(n12404), .B(n12405), .Z(n12023) );
  AND U12164 ( .A(n344), .B(n12406), .Z(n12405) );
  XOR U12165 ( .A(n12407), .B(n12404), .Z(n12406) );
  XOR U12166 ( .A(n12408), .B(n12409), .Z(n12396) );
  AND U12167 ( .A(n12410), .B(n12411), .Z(n12409) );
  XOR U12168 ( .A(n12408), .B(n12038), .Z(n12411) );
  XOR U12169 ( .A(n12412), .B(n12413), .Z(n12038) );
  AND U12170 ( .A(n346), .B(n12414), .Z(n12413) );
  XOR U12171 ( .A(n12415), .B(n12412), .Z(n12414) );
  XNOR U12172 ( .A(n12035), .B(n12408), .Z(n12410) );
  XOR U12173 ( .A(n12416), .B(n12417), .Z(n12035) );
  AND U12174 ( .A(n344), .B(n12418), .Z(n12417) );
  XOR U12175 ( .A(n12419), .B(n12416), .Z(n12418) );
  XOR U12176 ( .A(n12420), .B(n12421), .Z(n12408) );
  AND U12177 ( .A(n12422), .B(n12423), .Z(n12421) );
  XOR U12178 ( .A(n12420), .B(n12050), .Z(n12423) );
  XOR U12179 ( .A(n12424), .B(n12425), .Z(n12050) );
  AND U12180 ( .A(n346), .B(n12426), .Z(n12425) );
  XOR U12181 ( .A(n12427), .B(n12424), .Z(n12426) );
  XNOR U12182 ( .A(n12047), .B(n12420), .Z(n12422) );
  XOR U12183 ( .A(n12428), .B(n12429), .Z(n12047) );
  AND U12184 ( .A(n344), .B(n12430), .Z(n12429) );
  XOR U12185 ( .A(n12431), .B(n12428), .Z(n12430) );
  XOR U12186 ( .A(n12432), .B(n12433), .Z(n12420) );
  AND U12187 ( .A(n12434), .B(n12435), .Z(n12433) );
  XOR U12188 ( .A(n12432), .B(n12062), .Z(n12435) );
  XOR U12189 ( .A(n12436), .B(n12437), .Z(n12062) );
  AND U12190 ( .A(n346), .B(n12438), .Z(n12437) );
  XOR U12191 ( .A(n12439), .B(n12436), .Z(n12438) );
  XNOR U12192 ( .A(n12059), .B(n12432), .Z(n12434) );
  XOR U12193 ( .A(n12440), .B(n12441), .Z(n12059) );
  AND U12194 ( .A(n344), .B(n12442), .Z(n12441) );
  XOR U12195 ( .A(n12443), .B(n12440), .Z(n12442) );
  XOR U12196 ( .A(n12444), .B(n12445), .Z(n12432) );
  AND U12197 ( .A(n12446), .B(n12447), .Z(n12445) );
  XOR U12198 ( .A(n12444), .B(n12074), .Z(n12447) );
  XOR U12199 ( .A(n12448), .B(n12449), .Z(n12074) );
  AND U12200 ( .A(n346), .B(n12450), .Z(n12449) );
  XOR U12201 ( .A(n12451), .B(n12448), .Z(n12450) );
  XNOR U12202 ( .A(n12071), .B(n12444), .Z(n12446) );
  XOR U12203 ( .A(n12452), .B(n12453), .Z(n12071) );
  AND U12204 ( .A(n344), .B(n12454), .Z(n12453) );
  XOR U12205 ( .A(n12455), .B(n12452), .Z(n12454) );
  XOR U12206 ( .A(n12456), .B(n12457), .Z(n12444) );
  AND U12207 ( .A(n12458), .B(n12459), .Z(n12457) );
  XOR U12208 ( .A(n12456), .B(n12086), .Z(n12459) );
  XOR U12209 ( .A(n12460), .B(n12461), .Z(n12086) );
  AND U12210 ( .A(n346), .B(n12462), .Z(n12461) );
  XOR U12211 ( .A(n12463), .B(n12460), .Z(n12462) );
  XNOR U12212 ( .A(n12083), .B(n12456), .Z(n12458) );
  XOR U12213 ( .A(n12464), .B(n12465), .Z(n12083) );
  AND U12214 ( .A(n344), .B(n12466), .Z(n12465) );
  XOR U12215 ( .A(n12467), .B(n12464), .Z(n12466) );
  XOR U12216 ( .A(n12468), .B(n12469), .Z(n12456) );
  AND U12217 ( .A(n12470), .B(n12471), .Z(n12469) );
  XOR U12218 ( .A(n12468), .B(n12098), .Z(n12471) );
  XOR U12219 ( .A(n12472), .B(n12473), .Z(n12098) );
  AND U12220 ( .A(n346), .B(n12474), .Z(n12473) );
  XOR U12221 ( .A(n12475), .B(n12472), .Z(n12474) );
  XNOR U12222 ( .A(n12095), .B(n12468), .Z(n12470) );
  XOR U12223 ( .A(n12476), .B(n12477), .Z(n12095) );
  AND U12224 ( .A(n344), .B(n12478), .Z(n12477) );
  XOR U12225 ( .A(n12479), .B(n12476), .Z(n12478) );
  XOR U12226 ( .A(n12480), .B(n12481), .Z(n12468) );
  AND U12227 ( .A(n12482), .B(n12483), .Z(n12481) );
  XOR U12228 ( .A(n12480), .B(n12110), .Z(n12483) );
  XOR U12229 ( .A(n12484), .B(n12485), .Z(n12110) );
  AND U12230 ( .A(n346), .B(n12486), .Z(n12485) );
  XOR U12231 ( .A(n12487), .B(n12484), .Z(n12486) );
  XNOR U12232 ( .A(n12107), .B(n12480), .Z(n12482) );
  XOR U12233 ( .A(n12488), .B(n12489), .Z(n12107) );
  AND U12234 ( .A(n344), .B(n12490), .Z(n12489) );
  XOR U12235 ( .A(n12491), .B(n12488), .Z(n12490) );
  XOR U12236 ( .A(n12492), .B(n12493), .Z(n12480) );
  AND U12237 ( .A(n12494), .B(n12495), .Z(n12493) );
  XOR U12238 ( .A(n12492), .B(n12122), .Z(n12495) );
  XOR U12239 ( .A(n12496), .B(n12497), .Z(n12122) );
  AND U12240 ( .A(n346), .B(n12498), .Z(n12497) );
  XOR U12241 ( .A(n12499), .B(n12496), .Z(n12498) );
  XNOR U12242 ( .A(n12119), .B(n12492), .Z(n12494) );
  XOR U12243 ( .A(n12500), .B(n12501), .Z(n12119) );
  AND U12244 ( .A(n344), .B(n12502), .Z(n12501) );
  XOR U12245 ( .A(n12503), .B(n12500), .Z(n12502) );
  XOR U12246 ( .A(n12504), .B(n12505), .Z(n12492) );
  AND U12247 ( .A(n12506), .B(n12507), .Z(n12505) );
  XOR U12248 ( .A(n12504), .B(n12134), .Z(n12507) );
  XOR U12249 ( .A(n12508), .B(n12509), .Z(n12134) );
  AND U12250 ( .A(n346), .B(n12510), .Z(n12509) );
  XOR U12251 ( .A(n12511), .B(n12508), .Z(n12510) );
  XNOR U12252 ( .A(n12131), .B(n12504), .Z(n12506) );
  XOR U12253 ( .A(n12512), .B(n12513), .Z(n12131) );
  AND U12254 ( .A(n344), .B(n12514), .Z(n12513) );
  XOR U12255 ( .A(n12515), .B(n12512), .Z(n12514) );
  XOR U12256 ( .A(n12516), .B(n12517), .Z(n12504) );
  AND U12257 ( .A(n12518), .B(n12519), .Z(n12517) );
  XOR U12258 ( .A(n12516), .B(n12146), .Z(n12519) );
  XOR U12259 ( .A(n12520), .B(n12521), .Z(n12146) );
  AND U12260 ( .A(n346), .B(n12522), .Z(n12521) );
  XOR U12261 ( .A(n12523), .B(n12520), .Z(n12522) );
  XNOR U12262 ( .A(n12143), .B(n12516), .Z(n12518) );
  XOR U12263 ( .A(n12524), .B(n12525), .Z(n12143) );
  AND U12264 ( .A(n344), .B(n12526), .Z(n12525) );
  XOR U12265 ( .A(n12527), .B(n12524), .Z(n12526) );
  XOR U12266 ( .A(n12528), .B(n12529), .Z(n12516) );
  AND U12267 ( .A(n12530), .B(n12531), .Z(n12529) );
  XOR U12268 ( .A(n12528), .B(n12158), .Z(n12531) );
  XOR U12269 ( .A(n12532), .B(n12533), .Z(n12158) );
  AND U12270 ( .A(n346), .B(n12534), .Z(n12533) );
  XOR U12271 ( .A(n12535), .B(n12532), .Z(n12534) );
  XNOR U12272 ( .A(n12155), .B(n12528), .Z(n12530) );
  XOR U12273 ( .A(n12536), .B(n12537), .Z(n12155) );
  AND U12274 ( .A(n344), .B(n12538), .Z(n12537) );
  XOR U12275 ( .A(n12539), .B(n12536), .Z(n12538) );
  XOR U12276 ( .A(n12540), .B(n12541), .Z(n12528) );
  AND U12277 ( .A(n12542), .B(n12543), .Z(n12541) );
  XOR U12278 ( .A(n12540), .B(n12170), .Z(n12543) );
  XOR U12279 ( .A(n12544), .B(n12545), .Z(n12170) );
  AND U12280 ( .A(n346), .B(n12546), .Z(n12545) );
  XOR U12281 ( .A(n12547), .B(n12544), .Z(n12546) );
  XNOR U12282 ( .A(n12167), .B(n12540), .Z(n12542) );
  XOR U12283 ( .A(n12548), .B(n12549), .Z(n12167) );
  AND U12284 ( .A(n344), .B(n12550), .Z(n12549) );
  XOR U12285 ( .A(n12551), .B(n12548), .Z(n12550) );
  XOR U12286 ( .A(n12552), .B(n12553), .Z(n12540) );
  AND U12287 ( .A(n12554), .B(n12555), .Z(n12553) );
  XOR U12288 ( .A(n12552), .B(n12182), .Z(n12555) );
  XOR U12289 ( .A(n12556), .B(n12557), .Z(n12182) );
  AND U12290 ( .A(n346), .B(n12558), .Z(n12557) );
  XOR U12291 ( .A(n12559), .B(n12556), .Z(n12558) );
  XNOR U12292 ( .A(n12179), .B(n12552), .Z(n12554) );
  XOR U12293 ( .A(n12560), .B(n12561), .Z(n12179) );
  AND U12294 ( .A(n344), .B(n12562), .Z(n12561) );
  XOR U12295 ( .A(n12563), .B(n12560), .Z(n12562) );
  XOR U12296 ( .A(n12564), .B(n12565), .Z(n12552) );
  AND U12297 ( .A(n12566), .B(n12567), .Z(n12565) );
  XOR U12298 ( .A(n12564), .B(n12194), .Z(n12567) );
  XOR U12299 ( .A(n12568), .B(n12569), .Z(n12194) );
  AND U12300 ( .A(n346), .B(n12570), .Z(n12569) );
  XOR U12301 ( .A(n12571), .B(n12568), .Z(n12570) );
  XNOR U12302 ( .A(n12191), .B(n12564), .Z(n12566) );
  XOR U12303 ( .A(n12572), .B(n12573), .Z(n12191) );
  AND U12304 ( .A(n344), .B(n12574), .Z(n12573) );
  XOR U12305 ( .A(n12575), .B(n12572), .Z(n12574) );
  XOR U12306 ( .A(n12576), .B(n12577), .Z(n12564) );
  AND U12307 ( .A(n12578), .B(n12579), .Z(n12577) );
  XOR U12308 ( .A(n12576), .B(n12206), .Z(n12579) );
  XOR U12309 ( .A(n12580), .B(n12581), .Z(n12206) );
  AND U12310 ( .A(n346), .B(n12582), .Z(n12581) );
  XOR U12311 ( .A(n12583), .B(n12580), .Z(n12582) );
  XNOR U12312 ( .A(n12203), .B(n12576), .Z(n12578) );
  XOR U12313 ( .A(n12584), .B(n12585), .Z(n12203) );
  AND U12314 ( .A(n344), .B(n12586), .Z(n12585) );
  XOR U12315 ( .A(n12587), .B(n12584), .Z(n12586) );
  XOR U12316 ( .A(n12588), .B(n12589), .Z(n12576) );
  AND U12317 ( .A(n12590), .B(n12591), .Z(n12589) );
  XOR U12318 ( .A(n12588), .B(n12218), .Z(n12591) );
  XOR U12319 ( .A(n12592), .B(n12593), .Z(n12218) );
  AND U12320 ( .A(n346), .B(n12594), .Z(n12593) );
  XOR U12321 ( .A(n12595), .B(n12592), .Z(n12594) );
  XNOR U12322 ( .A(n12215), .B(n12588), .Z(n12590) );
  XOR U12323 ( .A(n12596), .B(n12597), .Z(n12215) );
  AND U12324 ( .A(n344), .B(n12598), .Z(n12597) );
  XOR U12325 ( .A(n12599), .B(n12596), .Z(n12598) );
  XOR U12326 ( .A(n12600), .B(n12601), .Z(n12588) );
  AND U12327 ( .A(n12602), .B(n12603), .Z(n12601) );
  XOR U12328 ( .A(n12600), .B(n12230), .Z(n12603) );
  XOR U12329 ( .A(n12604), .B(n12605), .Z(n12230) );
  AND U12330 ( .A(n346), .B(n12606), .Z(n12605) );
  XOR U12331 ( .A(n12607), .B(n12604), .Z(n12606) );
  XNOR U12332 ( .A(n12227), .B(n12600), .Z(n12602) );
  XOR U12333 ( .A(n12608), .B(n12609), .Z(n12227) );
  AND U12334 ( .A(n344), .B(n12610), .Z(n12609) );
  XOR U12335 ( .A(n12611), .B(n12608), .Z(n12610) );
  XOR U12336 ( .A(n12612), .B(n12613), .Z(n12600) );
  AND U12337 ( .A(n12614), .B(n12615), .Z(n12613) );
  XOR U12338 ( .A(n12612), .B(n12242), .Z(n12615) );
  XOR U12339 ( .A(n12616), .B(n12617), .Z(n12242) );
  AND U12340 ( .A(n346), .B(n12618), .Z(n12617) );
  XOR U12341 ( .A(n12619), .B(n12616), .Z(n12618) );
  XNOR U12342 ( .A(n12239), .B(n12612), .Z(n12614) );
  XOR U12343 ( .A(n12620), .B(n12621), .Z(n12239) );
  AND U12344 ( .A(n344), .B(n12622), .Z(n12621) );
  XOR U12345 ( .A(n12623), .B(n12620), .Z(n12622) );
  XOR U12346 ( .A(n12624), .B(n12625), .Z(n12612) );
  AND U12347 ( .A(n12626), .B(n12627), .Z(n12625) );
  XOR U12348 ( .A(n12624), .B(n12254), .Z(n12627) );
  XOR U12349 ( .A(n12628), .B(n12629), .Z(n12254) );
  AND U12350 ( .A(n346), .B(n12630), .Z(n12629) );
  XOR U12351 ( .A(n12631), .B(n12628), .Z(n12630) );
  XNOR U12352 ( .A(n12251), .B(n12624), .Z(n12626) );
  XOR U12353 ( .A(n12632), .B(n12633), .Z(n12251) );
  AND U12354 ( .A(n344), .B(n12634), .Z(n12633) );
  XOR U12355 ( .A(n12635), .B(n12632), .Z(n12634) );
  XOR U12356 ( .A(n12636), .B(n12637), .Z(n12624) );
  AND U12357 ( .A(n12638), .B(n12639), .Z(n12637) );
  XOR U12358 ( .A(n12636), .B(n12266), .Z(n12639) );
  XOR U12359 ( .A(n12640), .B(n12641), .Z(n12266) );
  AND U12360 ( .A(n346), .B(n12642), .Z(n12641) );
  XOR U12361 ( .A(n12643), .B(n12640), .Z(n12642) );
  XNOR U12362 ( .A(n12263), .B(n12636), .Z(n12638) );
  XOR U12363 ( .A(n12644), .B(n12645), .Z(n12263) );
  AND U12364 ( .A(n344), .B(n12646), .Z(n12645) );
  XOR U12365 ( .A(n12647), .B(n12644), .Z(n12646) );
  XOR U12366 ( .A(n12648), .B(n12649), .Z(n12636) );
  AND U12367 ( .A(n12650), .B(n12651), .Z(n12649) );
  XOR U12368 ( .A(n12648), .B(n12278), .Z(n12651) );
  XOR U12369 ( .A(n12652), .B(n12653), .Z(n12278) );
  AND U12370 ( .A(n346), .B(n12654), .Z(n12653) );
  XOR U12371 ( .A(n12655), .B(n12652), .Z(n12654) );
  XNOR U12372 ( .A(n12275), .B(n12648), .Z(n12650) );
  XOR U12373 ( .A(n12656), .B(n12657), .Z(n12275) );
  AND U12374 ( .A(n344), .B(n12658), .Z(n12657) );
  XOR U12375 ( .A(n12659), .B(n12656), .Z(n12658) );
  XOR U12376 ( .A(n12660), .B(n12661), .Z(n12648) );
  AND U12377 ( .A(n12662), .B(n12663), .Z(n12661) );
  XOR U12378 ( .A(n12660), .B(n12290), .Z(n12663) );
  XOR U12379 ( .A(n12664), .B(n12665), .Z(n12290) );
  AND U12380 ( .A(n346), .B(n12666), .Z(n12665) );
  XOR U12381 ( .A(n12667), .B(n12664), .Z(n12666) );
  XNOR U12382 ( .A(n12287), .B(n12660), .Z(n12662) );
  XOR U12383 ( .A(n12668), .B(n12669), .Z(n12287) );
  AND U12384 ( .A(n344), .B(n12670), .Z(n12669) );
  XOR U12385 ( .A(n12671), .B(n12668), .Z(n12670) );
  XOR U12386 ( .A(n12672), .B(n12673), .Z(n12660) );
  AND U12387 ( .A(n12674), .B(n12675), .Z(n12673) );
  XOR U12388 ( .A(n12302), .B(n12672), .Z(n12675) );
  XOR U12389 ( .A(n12676), .B(n12677), .Z(n12302) );
  AND U12390 ( .A(n346), .B(n12678), .Z(n12677) );
  XOR U12391 ( .A(n12676), .B(n12679), .Z(n12678) );
  XNOR U12392 ( .A(n12672), .B(n12299), .Z(n12674) );
  XOR U12393 ( .A(n12680), .B(n12681), .Z(n12299) );
  AND U12394 ( .A(n344), .B(n12682), .Z(n12681) );
  XOR U12395 ( .A(n12680), .B(n12683), .Z(n12682) );
  XOR U12396 ( .A(n12684), .B(n12685), .Z(n12672) );
  AND U12397 ( .A(n12686), .B(n12687), .Z(n12685) );
  XNOR U12398 ( .A(n12688), .B(n12315), .Z(n12687) );
  XOR U12399 ( .A(n12689), .B(n12690), .Z(n12315) );
  AND U12400 ( .A(n346), .B(n12691), .Z(n12690) );
  XOR U12401 ( .A(n12692), .B(n12689), .Z(n12691) );
  XNOR U12402 ( .A(n12312), .B(n12684), .Z(n12686) );
  XOR U12403 ( .A(n12693), .B(n12694), .Z(n12312) );
  AND U12404 ( .A(n344), .B(n12695), .Z(n12694) );
  XOR U12405 ( .A(n12696), .B(n12693), .Z(n12695) );
  IV U12406 ( .A(n12688), .Z(n12684) );
  AND U12407 ( .A(n12320), .B(n12323), .Z(n12688) );
  XNOR U12408 ( .A(n12697), .B(n12698), .Z(n12323) );
  AND U12409 ( .A(n346), .B(n12699), .Z(n12698) );
  XNOR U12410 ( .A(n12700), .B(n12697), .Z(n12699) );
  XOR U12411 ( .A(n12701), .B(n12702), .Z(n346) );
  AND U12412 ( .A(n12703), .B(n12704), .Z(n12702) );
  XOR U12413 ( .A(n12331), .B(n12701), .Z(n12704) );
  IV U12414 ( .A(n12705), .Z(n12331) );
  AND U12415 ( .A(p_input[2559]), .B(p_input[2527]), .Z(n12705) );
  XOR U12416 ( .A(n12701), .B(n12328), .Z(n12703) );
  AND U12417 ( .A(p_input[2463]), .B(p_input[2495]), .Z(n12328) );
  XOR U12418 ( .A(n12706), .B(n12707), .Z(n12701) );
  AND U12419 ( .A(n12708), .B(n12709), .Z(n12707) );
  XOR U12420 ( .A(n12706), .B(n12343), .Z(n12709) );
  XNOR U12421 ( .A(p_input[2526]), .B(n12710), .Z(n12343) );
  AND U12422 ( .A(n270), .B(n12711), .Z(n12710) );
  XOR U12423 ( .A(p_input[2558]), .B(p_input[2526]), .Z(n12711) );
  XNOR U12424 ( .A(n12340), .B(n12706), .Z(n12708) );
  XOR U12425 ( .A(n12712), .B(n12713), .Z(n12340) );
  AND U12426 ( .A(n268), .B(n12714), .Z(n12713) );
  XOR U12427 ( .A(p_input[2494]), .B(p_input[2462]), .Z(n12714) );
  XOR U12428 ( .A(n12715), .B(n12716), .Z(n12706) );
  AND U12429 ( .A(n12717), .B(n12718), .Z(n12716) );
  XOR U12430 ( .A(n12715), .B(n12355), .Z(n12718) );
  XNOR U12431 ( .A(p_input[2525]), .B(n12719), .Z(n12355) );
  AND U12432 ( .A(n270), .B(n12720), .Z(n12719) );
  XOR U12433 ( .A(p_input[2557]), .B(p_input[2525]), .Z(n12720) );
  XNOR U12434 ( .A(n12352), .B(n12715), .Z(n12717) );
  XOR U12435 ( .A(n12721), .B(n12722), .Z(n12352) );
  AND U12436 ( .A(n268), .B(n12723), .Z(n12722) );
  XOR U12437 ( .A(p_input[2493]), .B(p_input[2461]), .Z(n12723) );
  XOR U12438 ( .A(n12724), .B(n12725), .Z(n12715) );
  AND U12439 ( .A(n12726), .B(n12727), .Z(n12725) );
  XOR U12440 ( .A(n12724), .B(n12367), .Z(n12727) );
  XNOR U12441 ( .A(p_input[2524]), .B(n12728), .Z(n12367) );
  AND U12442 ( .A(n270), .B(n12729), .Z(n12728) );
  XOR U12443 ( .A(p_input[2556]), .B(p_input[2524]), .Z(n12729) );
  XNOR U12444 ( .A(n12364), .B(n12724), .Z(n12726) );
  XOR U12445 ( .A(n12730), .B(n12731), .Z(n12364) );
  AND U12446 ( .A(n268), .B(n12732), .Z(n12731) );
  XOR U12447 ( .A(p_input[2492]), .B(p_input[2460]), .Z(n12732) );
  XOR U12448 ( .A(n12733), .B(n12734), .Z(n12724) );
  AND U12449 ( .A(n12735), .B(n12736), .Z(n12734) );
  XOR U12450 ( .A(n12733), .B(n12379), .Z(n12736) );
  XNOR U12451 ( .A(p_input[2523]), .B(n12737), .Z(n12379) );
  AND U12452 ( .A(n270), .B(n12738), .Z(n12737) );
  XOR U12453 ( .A(p_input[2555]), .B(p_input[2523]), .Z(n12738) );
  XNOR U12454 ( .A(n12376), .B(n12733), .Z(n12735) );
  XOR U12455 ( .A(n12739), .B(n12740), .Z(n12376) );
  AND U12456 ( .A(n268), .B(n12741), .Z(n12740) );
  XOR U12457 ( .A(p_input[2491]), .B(p_input[2459]), .Z(n12741) );
  XOR U12458 ( .A(n12742), .B(n12743), .Z(n12733) );
  AND U12459 ( .A(n12744), .B(n12745), .Z(n12743) );
  XOR U12460 ( .A(n12742), .B(n12391), .Z(n12745) );
  XNOR U12461 ( .A(p_input[2522]), .B(n12746), .Z(n12391) );
  AND U12462 ( .A(n270), .B(n12747), .Z(n12746) );
  XOR U12463 ( .A(p_input[2554]), .B(p_input[2522]), .Z(n12747) );
  XNOR U12464 ( .A(n12388), .B(n12742), .Z(n12744) );
  XOR U12465 ( .A(n12748), .B(n12749), .Z(n12388) );
  AND U12466 ( .A(n268), .B(n12750), .Z(n12749) );
  XOR U12467 ( .A(p_input[2490]), .B(p_input[2458]), .Z(n12750) );
  XOR U12468 ( .A(n12751), .B(n12752), .Z(n12742) );
  AND U12469 ( .A(n12753), .B(n12754), .Z(n12752) );
  XOR U12470 ( .A(n12751), .B(n12403), .Z(n12754) );
  XNOR U12471 ( .A(p_input[2521]), .B(n12755), .Z(n12403) );
  AND U12472 ( .A(n270), .B(n12756), .Z(n12755) );
  XOR U12473 ( .A(p_input[2553]), .B(p_input[2521]), .Z(n12756) );
  XNOR U12474 ( .A(n12400), .B(n12751), .Z(n12753) );
  XOR U12475 ( .A(n12757), .B(n12758), .Z(n12400) );
  AND U12476 ( .A(n268), .B(n12759), .Z(n12758) );
  XOR U12477 ( .A(p_input[2489]), .B(p_input[2457]), .Z(n12759) );
  XOR U12478 ( .A(n12760), .B(n12761), .Z(n12751) );
  AND U12479 ( .A(n12762), .B(n12763), .Z(n12761) );
  XOR U12480 ( .A(n12760), .B(n12415), .Z(n12763) );
  XNOR U12481 ( .A(p_input[2520]), .B(n12764), .Z(n12415) );
  AND U12482 ( .A(n270), .B(n12765), .Z(n12764) );
  XOR U12483 ( .A(p_input[2552]), .B(p_input[2520]), .Z(n12765) );
  XNOR U12484 ( .A(n12412), .B(n12760), .Z(n12762) );
  XOR U12485 ( .A(n12766), .B(n12767), .Z(n12412) );
  AND U12486 ( .A(n268), .B(n12768), .Z(n12767) );
  XOR U12487 ( .A(p_input[2488]), .B(p_input[2456]), .Z(n12768) );
  XOR U12488 ( .A(n12769), .B(n12770), .Z(n12760) );
  AND U12489 ( .A(n12771), .B(n12772), .Z(n12770) );
  XOR U12490 ( .A(n12769), .B(n12427), .Z(n12772) );
  XNOR U12491 ( .A(p_input[2519]), .B(n12773), .Z(n12427) );
  AND U12492 ( .A(n270), .B(n12774), .Z(n12773) );
  XOR U12493 ( .A(p_input[2551]), .B(p_input[2519]), .Z(n12774) );
  XNOR U12494 ( .A(n12424), .B(n12769), .Z(n12771) );
  XOR U12495 ( .A(n12775), .B(n12776), .Z(n12424) );
  AND U12496 ( .A(n268), .B(n12777), .Z(n12776) );
  XOR U12497 ( .A(p_input[2487]), .B(p_input[2455]), .Z(n12777) );
  XOR U12498 ( .A(n12778), .B(n12779), .Z(n12769) );
  AND U12499 ( .A(n12780), .B(n12781), .Z(n12779) );
  XOR U12500 ( .A(n12778), .B(n12439), .Z(n12781) );
  XNOR U12501 ( .A(p_input[2518]), .B(n12782), .Z(n12439) );
  AND U12502 ( .A(n270), .B(n12783), .Z(n12782) );
  XOR U12503 ( .A(p_input[2550]), .B(p_input[2518]), .Z(n12783) );
  XNOR U12504 ( .A(n12436), .B(n12778), .Z(n12780) );
  XOR U12505 ( .A(n12784), .B(n12785), .Z(n12436) );
  AND U12506 ( .A(n268), .B(n12786), .Z(n12785) );
  XOR U12507 ( .A(p_input[2486]), .B(p_input[2454]), .Z(n12786) );
  XOR U12508 ( .A(n12787), .B(n12788), .Z(n12778) );
  AND U12509 ( .A(n12789), .B(n12790), .Z(n12788) );
  XOR U12510 ( .A(n12787), .B(n12451), .Z(n12790) );
  XNOR U12511 ( .A(p_input[2517]), .B(n12791), .Z(n12451) );
  AND U12512 ( .A(n270), .B(n12792), .Z(n12791) );
  XOR U12513 ( .A(p_input[2549]), .B(p_input[2517]), .Z(n12792) );
  XNOR U12514 ( .A(n12448), .B(n12787), .Z(n12789) );
  XOR U12515 ( .A(n12793), .B(n12794), .Z(n12448) );
  AND U12516 ( .A(n268), .B(n12795), .Z(n12794) );
  XOR U12517 ( .A(p_input[2485]), .B(p_input[2453]), .Z(n12795) );
  XOR U12518 ( .A(n12796), .B(n12797), .Z(n12787) );
  AND U12519 ( .A(n12798), .B(n12799), .Z(n12797) );
  XOR U12520 ( .A(n12796), .B(n12463), .Z(n12799) );
  XNOR U12521 ( .A(p_input[2516]), .B(n12800), .Z(n12463) );
  AND U12522 ( .A(n270), .B(n12801), .Z(n12800) );
  XOR U12523 ( .A(p_input[2548]), .B(p_input[2516]), .Z(n12801) );
  XNOR U12524 ( .A(n12460), .B(n12796), .Z(n12798) );
  XOR U12525 ( .A(n12802), .B(n12803), .Z(n12460) );
  AND U12526 ( .A(n268), .B(n12804), .Z(n12803) );
  XOR U12527 ( .A(p_input[2484]), .B(p_input[2452]), .Z(n12804) );
  XOR U12528 ( .A(n12805), .B(n12806), .Z(n12796) );
  AND U12529 ( .A(n12807), .B(n12808), .Z(n12806) );
  XOR U12530 ( .A(n12805), .B(n12475), .Z(n12808) );
  XNOR U12531 ( .A(p_input[2515]), .B(n12809), .Z(n12475) );
  AND U12532 ( .A(n270), .B(n12810), .Z(n12809) );
  XOR U12533 ( .A(p_input[2547]), .B(p_input[2515]), .Z(n12810) );
  XNOR U12534 ( .A(n12472), .B(n12805), .Z(n12807) );
  XOR U12535 ( .A(n12811), .B(n12812), .Z(n12472) );
  AND U12536 ( .A(n268), .B(n12813), .Z(n12812) );
  XOR U12537 ( .A(p_input[2483]), .B(p_input[2451]), .Z(n12813) );
  XOR U12538 ( .A(n12814), .B(n12815), .Z(n12805) );
  AND U12539 ( .A(n12816), .B(n12817), .Z(n12815) );
  XOR U12540 ( .A(n12814), .B(n12487), .Z(n12817) );
  XNOR U12541 ( .A(p_input[2514]), .B(n12818), .Z(n12487) );
  AND U12542 ( .A(n270), .B(n12819), .Z(n12818) );
  XOR U12543 ( .A(p_input[2546]), .B(p_input[2514]), .Z(n12819) );
  XNOR U12544 ( .A(n12484), .B(n12814), .Z(n12816) );
  XOR U12545 ( .A(n12820), .B(n12821), .Z(n12484) );
  AND U12546 ( .A(n268), .B(n12822), .Z(n12821) );
  XOR U12547 ( .A(p_input[2482]), .B(p_input[2450]), .Z(n12822) );
  XOR U12548 ( .A(n12823), .B(n12824), .Z(n12814) );
  AND U12549 ( .A(n12825), .B(n12826), .Z(n12824) );
  XOR U12550 ( .A(n12823), .B(n12499), .Z(n12826) );
  XNOR U12551 ( .A(p_input[2513]), .B(n12827), .Z(n12499) );
  AND U12552 ( .A(n270), .B(n12828), .Z(n12827) );
  XOR U12553 ( .A(p_input[2545]), .B(p_input[2513]), .Z(n12828) );
  XNOR U12554 ( .A(n12496), .B(n12823), .Z(n12825) );
  XOR U12555 ( .A(n12829), .B(n12830), .Z(n12496) );
  AND U12556 ( .A(n268), .B(n12831), .Z(n12830) );
  XOR U12557 ( .A(p_input[2481]), .B(p_input[2449]), .Z(n12831) );
  XOR U12558 ( .A(n12832), .B(n12833), .Z(n12823) );
  AND U12559 ( .A(n12834), .B(n12835), .Z(n12833) );
  XOR U12560 ( .A(n12832), .B(n12511), .Z(n12835) );
  XNOR U12561 ( .A(p_input[2512]), .B(n12836), .Z(n12511) );
  AND U12562 ( .A(n270), .B(n12837), .Z(n12836) );
  XOR U12563 ( .A(p_input[2544]), .B(p_input[2512]), .Z(n12837) );
  XNOR U12564 ( .A(n12508), .B(n12832), .Z(n12834) );
  XOR U12565 ( .A(n12838), .B(n12839), .Z(n12508) );
  AND U12566 ( .A(n268), .B(n12840), .Z(n12839) );
  XOR U12567 ( .A(p_input[2480]), .B(p_input[2448]), .Z(n12840) );
  XOR U12568 ( .A(n12841), .B(n12842), .Z(n12832) );
  AND U12569 ( .A(n12843), .B(n12844), .Z(n12842) );
  XOR U12570 ( .A(n12841), .B(n12523), .Z(n12844) );
  XNOR U12571 ( .A(p_input[2511]), .B(n12845), .Z(n12523) );
  AND U12572 ( .A(n270), .B(n12846), .Z(n12845) );
  XOR U12573 ( .A(p_input[2543]), .B(p_input[2511]), .Z(n12846) );
  XNOR U12574 ( .A(n12520), .B(n12841), .Z(n12843) );
  XOR U12575 ( .A(n12847), .B(n12848), .Z(n12520) );
  AND U12576 ( .A(n268), .B(n12849), .Z(n12848) );
  XOR U12577 ( .A(p_input[2479]), .B(p_input[2447]), .Z(n12849) );
  XOR U12578 ( .A(n12850), .B(n12851), .Z(n12841) );
  AND U12579 ( .A(n12852), .B(n12853), .Z(n12851) );
  XOR U12580 ( .A(n12850), .B(n12535), .Z(n12853) );
  XNOR U12581 ( .A(p_input[2510]), .B(n12854), .Z(n12535) );
  AND U12582 ( .A(n270), .B(n12855), .Z(n12854) );
  XOR U12583 ( .A(p_input[2542]), .B(p_input[2510]), .Z(n12855) );
  XNOR U12584 ( .A(n12532), .B(n12850), .Z(n12852) );
  XOR U12585 ( .A(n12856), .B(n12857), .Z(n12532) );
  AND U12586 ( .A(n268), .B(n12858), .Z(n12857) );
  XOR U12587 ( .A(p_input[2478]), .B(p_input[2446]), .Z(n12858) );
  XOR U12588 ( .A(n12859), .B(n12860), .Z(n12850) );
  AND U12589 ( .A(n12861), .B(n12862), .Z(n12860) );
  XOR U12590 ( .A(n12859), .B(n12547), .Z(n12862) );
  XNOR U12591 ( .A(p_input[2509]), .B(n12863), .Z(n12547) );
  AND U12592 ( .A(n270), .B(n12864), .Z(n12863) );
  XOR U12593 ( .A(p_input[2541]), .B(p_input[2509]), .Z(n12864) );
  XNOR U12594 ( .A(n12544), .B(n12859), .Z(n12861) );
  XOR U12595 ( .A(n12865), .B(n12866), .Z(n12544) );
  AND U12596 ( .A(n268), .B(n12867), .Z(n12866) );
  XOR U12597 ( .A(p_input[2477]), .B(p_input[2445]), .Z(n12867) );
  XOR U12598 ( .A(n12868), .B(n12869), .Z(n12859) );
  AND U12599 ( .A(n12870), .B(n12871), .Z(n12869) );
  XOR U12600 ( .A(n12868), .B(n12559), .Z(n12871) );
  XNOR U12601 ( .A(p_input[2508]), .B(n12872), .Z(n12559) );
  AND U12602 ( .A(n270), .B(n12873), .Z(n12872) );
  XOR U12603 ( .A(p_input[2540]), .B(p_input[2508]), .Z(n12873) );
  XNOR U12604 ( .A(n12556), .B(n12868), .Z(n12870) );
  XOR U12605 ( .A(n12874), .B(n12875), .Z(n12556) );
  AND U12606 ( .A(n268), .B(n12876), .Z(n12875) );
  XOR U12607 ( .A(p_input[2476]), .B(p_input[2444]), .Z(n12876) );
  XOR U12608 ( .A(n12877), .B(n12878), .Z(n12868) );
  AND U12609 ( .A(n12879), .B(n12880), .Z(n12878) );
  XOR U12610 ( .A(n12877), .B(n12571), .Z(n12880) );
  XNOR U12611 ( .A(p_input[2507]), .B(n12881), .Z(n12571) );
  AND U12612 ( .A(n270), .B(n12882), .Z(n12881) );
  XOR U12613 ( .A(p_input[2539]), .B(p_input[2507]), .Z(n12882) );
  XNOR U12614 ( .A(n12568), .B(n12877), .Z(n12879) );
  XOR U12615 ( .A(n12883), .B(n12884), .Z(n12568) );
  AND U12616 ( .A(n268), .B(n12885), .Z(n12884) );
  XOR U12617 ( .A(p_input[2475]), .B(p_input[2443]), .Z(n12885) );
  XOR U12618 ( .A(n12886), .B(n12887), .Z(n12877) );
  AND U12619 ( .A(n12888), .B(n12889), .Z(n12887) );
  XOR U12620 ( .A(n12886), .B(n12583), .Z(n12889) );
  XNOR U12621 ( .A(p_input[2506]), .B(n12890), .Z(n12583) );
  AND U12622 ( .A(n270), .B(n12891), .Z(n12890) );
  XOR U12623 ( .A(p_input[2538]), .B(p_input[2506]), .Z(n12891) );
  XNOR U12624 ( .A(n12580), .B(n12886), .Z(n12888) );
  XOR U12625 ( .A(n12892), .B(n12893), .Z(n12580) );
  AND U12626 ( .A(n268), .B(n12894), .Z(n12893) );
  XOR U12627 ( .A(p_input[2474]), .B(p_input[2442]), .Z(n12894) );
  XOR U12628 ( .A(n12895), .B(n12896), .Z(n12886) );
  AND U12629 ( .A(n12897), .B(n12898), .Z(n12896) );
  XOR U12630 ( .A(n12895), .B(n12595), .Z(n12898) );
  XNOR U12631 ( .A(p_input[2505]), .B(n12899), .Z(n12595) );
  AND U12632 ( .A(n270), .B(n12900), .Z(n12899) );
  XOR U12633 ( .A(p_input[2537]), .B(p_input[2505]), .Z(n12900) );
  XNOR U12634 ( .A(n12592), .B(n12895), .Z(n12897) );
  XOR U12635 ( .A(n12901), .B(n12902), .Z(n12592) );
  AND U12636 ( .A(n268), .B(n12903), .Z(n12902) );
  XOR U12637 ( .A(p_input[2473]), .B(p_input[2441]), .Z(n12903) );
  XOR U12638 ( .A(n12904), .B(n12905), .Z(n12895) );
  AND U12639 ( .A(n12906), .B(n12907), .Z(n12905) );
  XOR U12640 ( .A(n12904), .B(n12607), .Z(n12907) );
  XNOR U12641 ( .A(p_input[2504]), .B(n12908), .Z(n12607) );
  AND U12642 ( .A(n270), .B(n12909), .Z(n12908) );
  XOR U12643 ( .A(p_input[2536]), .B(p_input[2504]), .Z(n12909) );
  XNOR U12644 ( .A(n12604), .B(n12904), .Z(n12906) );
  XOR U12645 ( .A(n12910), .B(n12911), .Z(n12604) );
  AND U12646 ( .A(n268), .B(n12912), .Z(n12911) );
  XOR U12647 ( .A(p_input[2472]), .B(p_input[2440]), .Z(n12912) );
  XOR U12648 ( .A(n12913), .B(n12914), .Z(n12904) );
  AND U12649 ( .A(n12915), .B(n12916), .Z(n12914) );
  XOR U12650 ( .A(n12913), .B(n12619), .Z(n12916) );
  XNOR U12651 ( .A(p_input[2503]), .B(n12917), .Z(n12619) );
  AND U12652 ( .A(n270), .B(n12918), .Z(n12917) );
  XOR U12653 ( .A(p_input[2535]), .B(p_input[2503]), .Z(n12918) );
  XNOR U12654 ( .A(n12616), .B(n12913), .Z(n12915) );
  XOR U12655 ( .A(n12919), .B(n12920), .Z(n12616) );
  AND U12656 ( .A(n268), .B(n12921), .Z(n12920) );
  XOR U12657 ( .A(p_input[2471]), .B(p_input[2439]), .Z(n12921) );
  XOR U12658 ( .A(n12922), .B(n12923), .Z(n12913) );
  AND U12659 ( .A(n12924), .B(n12925), .Z(n12923) );
  XOR U12660 ( .A(n12922), .B(n12631), .Z(n12925) );
  XNOR U12661 ( .A(p_input[2502]), .B(n12926), .Z(n12631) );
  AND U12662 ( .A(n270), .B(n12927), .Z(n12926) );
  XOR U12663 ( .A(p_input[2534]), .B(p_input[2502]), .Z(n12927) );
  XNOR U12664 ( .A(n12628), .B(n12922), .Z(n12924) );
  XOR U12665 ( .A(n12928), .B(n12929), .Z(n12628) );
  AND U12666 ( .A(n268), .B(n12930), .Z(n12929) );
  XOR U12667 ( .A(p_input[2470]), .B(p_input[2438]), .Z(n12930) );
  XOR U12668 ( .A(n12931), .B(n12932), .Z(n12922) );
  AND U12669 ( .A(n12933), .B(n12934), .Z(n12932) );
  XOR U12670 ( .A(n12931), .B(n12643), .Z(n12934) );
  XNOR U12671 ( .A(p_input[2501]), .B(n12935), .Z(n12643) );
  AND U12672 ( .A(n270), .B(n12936), .Z(n12935) );
  XOR U12673 ( .A(p_input[2533]), .B(p_input[2501]), .Z(n12936) );
  XNOR U12674 ( .A(n12640), .B(n12931), .Z(n12933) );
  XOR U12675 ( .A(n12937), .B(n12938), .Z(n12640) );
  AND U12676 ( .A(n268), .B(n12939), .Z(n12938) );
  XOR U12677 ( .A(p_input[2469]), .B(p_input[2437]), .Z(n12939) );
  XOR U12678 ( .A(n12940), .B(n12941), .Z(n12931) );
  AND U12679 ( .A(n12942), .B(n12943), .Z(n12941) );
  XOR U12680 ( .A(n12940), .B(n12655), .Z(n12943) );
  XNOR U12681 ( .A(p_input[2500]), .B(n12944), .Z(n12655) );
  AND U12682 ( .A(n270), .B(n12945), .Z(n12944) );
  XOR U12683 ( .A(p_input[2532]), .B(p_input[2500]), .Z(n12945) );
  XNOR U12684 ( .A(n12652), .B(n12940), .Z(n12942) );
  XOR U12685 ( .A(n12946), .B(n12947), .Z(n12652) );
  AND U12686 ( .A(n268), .B(n12948), .Z(n12947) );
  XOR U12687 ( .A(p_input[2468]), .B(p_input[2436]), .Z(n12948) );
  XOR U12688 ( .A(n12949), .B(n12950), .Z(n12940) );
  AND U12689 ( .A(n12951), .B(n12952), .Z(n12950) );
  XOR U12690 ( .A(n12949), .B(n12667), .Z(n12952) );
  XNOR U12691 ( .A(p_input[2499]), .B(n12953), .Z(n12667) );
  AND U12692 ( .A(n270), .B(n12954), .Z(n12953) );
  XOR U12693 ( .A(p_input[2531]), .B(p_input[2499]), .Z(n12954) );
  XNOR U12694 ( .A(n12664), .B(n12949), .Z(n12951) );
  XOR U12695 ( .A(n12955), .B(n12956), .Z(n12664) );
  AND U12696 ( .A(n268), .B(n12957), .Z(n12956) );
  XOR U12697 ( .A(p_input[2467]), .B(p_input[2435]), .Z(n12957) );
  XOR U12698 ( .A(n12958), .B(n12959), .Z(n12949) );
  AND U12699 ( .A(n12960), .B(n12961), .Z(n12959) );
  XOR U12700 ( .A(n12679), .B(n12958), .Z(n12961) );
  XNOR U12701 ( .A(p_input[2498]), .B(n12962), .Z(n12679) );
  AND U12702 ( .A(n270), .B(n12963), .Z(n12962) );
  XOR U12703 ( .A(p_input[2530]), .B(p_input[2498]), .Z(n12963) );
  XNOR U12704 ( .A(n12958), .B(n12676), .Z(n12960) );
  XOR U12705 ( .A(n12964), .B(n12965), .Z(n12676) );
  AND U12706 ( .A(n268), .B(n12966), .Z(n12965) );
  XOR U12707 ( .A(p_input[2466]), .B(p_input[2434]), .Z(n12966) );
  XOR U12708 ( .A(n12967), .B(n12968), .Z(n12958) );
  AND U12709 ( .A(n12969), .B(n12970), .Z(n12968) );
  XNOR U12710 ( .A(n12971), .B(n12692), .Z(n12970) );
  XNOR U12711 ( .A(p_input[2497]), .B(n12972), .Z(n12692) );
  AND U12712 ( .A(n270), .B(n12973), .Z(n12972) );
  XNOR U12713 ( .A(p_input[2529]), .B(n12974), .Z(n12973) );
  IV U12714 ( .A(p_input[2497]), .Z(n12974) );
  XNOR U12715 ( .A(n12689), .B(n12967), .Z(n12969) );
  XNOR U12716 ( .A(p_input[2433]), .B(n12975), .Z(n12689) );
  AND U12717 ( .A(n268), .B(n12976), .Z(n12975) );
  XOR U12718 ( .A(p_input[2465]), .B(p_input[2433]), .Z(n12976) );
  IV U12719 ( .A(n12971), .Z(n12967) );
  AND U12720 ( .A(n12697), .B(n12700), .Z(n12971) );
  XOR U12721 ( .A(p_input[2496]), .B(n12977), .Z(n12700) );
  AND U12722 ( .A(n270), .B(n12978), .Z(n12977) );
  XOR U12723 ( .A(p_input[2528]), .B(p_input[2496]), .Z(n12978) );
  XOR U12724 ( .A(n12979), .B(n12980), .Z(n270) );
  AND U12725 ( .A(n12981), .B(n12982), .Z(n12980) );
  XNOR U12726 ( .A(p_input[2559]), .B(n12979), .Z(n12982) );
  XOR U12727 ( .A(n12979), .B(p_input[2527]), .Z(n12981) );
  XOR U12728 ( .A(n12983), .B(n12984), .Z(n12979) );
  AND U12729 ( .A(n12985), .B(n12986), .Z(n12984) );
  XNOR U12730 ( .A(p_input[2558]), .B(n12983), .Z(n12986) );
  XOR U12731 ( .A(n12983), .B(p_input[2526]), .Z(n12985) );
  XOR U12732 ( .A(n12987), .B(n12988), .Z(n12983) );
  AND U12733 ( .A(n12989), .B(n12990), .Z(n12988) );
  XNOR U12734 ( .A(p_input[2557]), .B(n12987), .Z(n12990) );
  XOR U12735 ( .A(n12987), .B(p_input[2525]), .Z(n12989) );
  XOR U12736 ( .A(n12991), .B(n12992), .Z(n12987) );
  AND U12737 ( .A(n12993), .B(n12994), .Z(n12992) );
  XNOR U12738 ( .A(p_input[2556]), .B(n12991), .Z(n12994) );
  XOR U12739 ( .A(n12991), .B(p_input[2524]), .Z(n12993) );
  XOR U12740 ( .A(n12995), .B(n12996), .Z(n12991) );
  AND U12741 ( .A(n12997), .B(n12998), .Z(n12996) );
  XNOR U12742 ( .A(p_input[2555]), .B(n12995), .Z(n12998) );
  XOR U12743 ( .A(n12995), .B(p_input[2523]), .Z(n12997) );
  XOR U12744 ( .A(n12999), .B(n13000), .Z(n12995) );
  AND U12745 ( .A(n13001), .B(n13002), .Z(n13000) );
  XNOR U12746 ( .A(p_input[2554]), .B(n12999), .Z(n13002) );
  XOR U12747 ( .A(n12999), .B(p_input[2522]), .Z(n13001) );
  XOR U12748 ( .A(n13003), .B(n13004), .Z(n12999) );
  AND U12749 ( .A(n13005), .B(n13006), .Z(n13004) );
  XNOR U12750 ( .A(p_input[2553]), .B(n13003), .Z(n13006) );
  XOR U12751 ( .A(n13003), .B(p_input[2521]), .Z(n13005) );
  XOR U12752 ( .A(n13007), .B(n13008), .Z(n13003) );
  AND U12753 ( .A(n13009), .B(n13010), .Z(n13008) );
  XNOR U12754 ( .A(p_input[2552]), .B(n13007), .Z(n13010) );
  XOR U12755 ( .A(n13007), .B(p_input[2520]), .Z(n13009) );
  XOR U12756 ( .A(n13011), .B(n13012), .Z(n13007) );
  AND U12757 ( .A(n13013), .B(n13014), .Z(n13012) );
  XNOR U12758 ( .A(p_input[2551]), .B(n13011), .Z(n13014) );
  XOR U12759 ( .A(n13011), .B(p_input[2519]), .Z(n13013) );
  XOR U12760 ( .A(n13015), .B(n13016), .Z(n13011) );
  AND U12761 ( .A(n13017), .B(n13018), .Z(n13016) );
  XNOR U12762 ( .A(p_input[2550]), .B(n13015), .Z(n13018) );
  XOR U12763 ( .A(n13015), .B(p_input[2518]), .Z(n13017) );
  XOR U12764 ( .A(n13019), .B(n13020), .Z(n13015) );
  AND U12765 ( .A(n13021), .B(n13022), .Z(n13020) );
  XNOR U12766 ( .A(p_input[2549]), .B(n13019), .Z(n13022) );
  XOR U12767 ( .A(n13019), .B(p_input[2517]), .Z(n13021) );
  XOR U12768 ( .A(n13023), .B(n13024), .Z(n13019) );
  AND U12769 ( .A(n13025), .B(n13026), .Z(n13024) );
  XNOR U12770 ( .A(p_input[2548]), .B(n13023), .Z(n13026) );
  XOR U12771 ( .A(n13023), .B(p_input[2516]), .Z(n13025) );
  XOR U12772 ( .A(n13027), .B(n13028), .Z(n13023) );
  AND U12773 ( .A(n13029), .B(n13030), .Z(n13028) );
  XNOR U12774 ( .A(p_input[2547]), .B(n13027), .Z(n13030) );
  XOR U12775 ( .A(n13027), .B(p_input[2515]), .Z(n13029) );
  XOR U12776 ( .A(n13031), .B(n13032), .Z(n13027) );
  AND U12777 ( .A(n13033), .B(n13034), .Z(n13032) );
  XNOR U12778 ( .A(p_input[2546]), .B(n13031), .Z(n13034) );
  XOR U12779 ( .A(n13031), .B(p_input[2514]), .Z(n13033) );
  XOR U12780 ( .A(n13035), .B(n13036), .Z(n13031) );
  AND U12781 ( .A(n13037), .B(n13038), .Z(n13036) );
  XNOR U12782 ( .A(p_input[2545]), .B(n13035), .Z(n13038) );
  XOR U12783 ( .A(n13035), .B(p_input[2513]), .Z(n13037) );
  XOR U12784 ( .A(n13039), .B(n13040), .Z(n13035) );
  AND U12785 ( .A(n13041), .B(n13042), .Z(n13040) );
  XNOR U12786 ( .A(p_input[2544]), .B(n13039), .Z(n13042) );
  XOR U12787 ( .A(n13039), .B(p_input[2512]), .Z(n13041) );
  XOR U12788 ( .A(n13043), .B(n13044), .Z(n13039) );
  AND U12789 ( .A(n13045), .B(n13046), .Z(n13044) );
  XNOR U12790 ( .A(p_input[2543]), .B(n13043), .Z(n13046) );
  XOR U12791 ( .A(n13043), .B(p_input[2511]), .Z(n13045) );
  XOR U12792 ( .A(n13047), .B(n13048), .Z(n13043) );
  AND U12793 ( .A(n13049), .B(n13050), .Z(n13048) );
  XNOR U12794 ( .A(p_input[2542]), .B(n13047), .Z(n13050) );
  XOR U12795 ( .A(n13047), .B(p_input[2510]), .Z(n13049) );
  XOR U12796 ( .A(n13051), .B(n13052), .Z(n13047) );
  AND U12797 ( .A(n13053), .B(n13054), .Z(n13052) );
  XNOR U12798 ( .A(p_input[2541]), .B(n13051), .Z(n13054) );
  XOR U12799 ( .A(n13051), .B(p_input[2509]), .Z(n13053) );
  XOR U12800 ( .A(n13055), .B(n13056), .Z(n13051) );
  AND U12801 ( .A(n13057), .B(n13058), .Z(n13056) );
  XNOR U12802 ( .A(p_input[2540]), .B(n13055), .Z(n13058) );
  XOR U12803 ( .A(n13055), .B(p_input[2508]), .Z(n13057) );
  XOR U12804 ( .A(n13059), .B(n13060), .Z(n13055) );
  AND U12805 ( .A(n13061), .B(n13062), .Z(n13060) );
  XNOR U12806 ( .A(p_input[2539]), .B(n13059), .Z(n13062) );
  XOR U12807 ( .A(n13059), .B(p_input[2507]), .Z(n13061) );
  XOR U12808 ( .A(n13063), .B(n13064), .Z(n13059) );
  AND U12809 ( .A(n13065), .B(n13066), .Z(n13064) );
  XNOR U12810 ( .A(p_input[2538]), .B(n13063), .Z(n13066) );
  XOR U12811 ( .A(n13063), .B(p_input[2506]), .Z(n13065) );
  XOR U12812 ( .A(n13067), .B(n13068), .Z(n13063) );
  AND U12813 ( .A(n13069), .B(n13070), .Z(n13068) );
  XNOR U12814 ( .A(p_input[2537]), .B(n13067), .Z(n13070) );
  XOR U12815 ( .A(n13067), .B(p_input[2505]), .Z(n13069) );
  XOR U12816 ( .A(n13071), .B(n13072), .Z(n13067) );
  AND U12817 ( .A(n13073), .B(n13074), .Z(n13072) );
  XNOR U12818 ( .A(p_input[2536]), .B(n13071), .Z(n13074) );
  XOR U12819 ( .A(n13071), .B(p_input[2504]), .Z(n13073) );
  XOR U12820 ( .A(n13075), .B(n13076), .Z(n13071) );
  AND U12821 ( .A(n13077), .B(n13078), .Z(n13076) );
  XNOR U12822 ( .A(p_input[2535]), .B(n13075), .Z(n13078) );
  XOR U12823 ( .A(n13075), .B(p_input[2503]), .Z(n13077) );
  XOR U12824 ( .A(n13079), .B(n13080), .Z(n13075) );
  AND U12825 ( .A(n13081), .B(n13082), .Z(n13080) );
  XNOR U12826 ( .A(p_input[2534]), .B(n13079), .Z(n13082) );
  XOR U12827 ( .A(n13079), .B(p_input[2502]), .Z(n13081) );
  XOR U12828 ( .A(n13083), .B(n13084), .Z(n13079) );
  AND U12829 ( .A(n13085), .B(n13086), .Z(n13084) );
  XNOR U12830 ( .A(p_input[2533]), .B(n13083), .Z(n13086) );
  XOR U12831 ( .A(n13083), .B(p_input[2501]), .Z(n13085) );
  XOR U12832 ( .A(n13087), .B(n13088), .Z(n13083) );
  AND U12833 ( .A(n13089), .B(n13090), .Z(n13088) );
  XNOR U12834 ( .A(p_input[2532]), .B(n13087), .Z(n13090) );
  XOR U12835 ( .A(n13087), .B(p_input[2500]), .Z(n13089) );
  XOR U12836 ( .A(n13091), .B(n13092), .Z(n13087) );
  AND U12837 ( .A(n13093), .B(n13094), .Z(n13092) );
  XNOR U12838 ( .A(p_input[2531]), .B(n13091), .Z(n13094) );
  XOR U12839 ( .A(n13091), .B(p_input[2499]), .Z(n13093) );
  XOR U12840 ( .A(n13095), .B(n13096), .Z(n13091) );
  AND U12841 ( .A(n13097), .B(n13098), .Z(n13096) );
  XNOR U12842 ( .A(p_input[2530]), .B(n13095), .Z(n13098) );
  XOR U12843 ( .A(n13095), .B(p_input[2498]), .Z(n13097) );
  XNOR U12844 ( .A(n13099), .B(n13100), .Z(n13095) );
  AND U12845 ( .A(n13101), .B(n13102), .Z(n13100) );
  XOR U12846 ( .A(p_input[2529]), .B(n13099), .Z(n13102) );
  XNOR U12847 ( .A(p_input[2497]), .B(n13099), .Z(n13101) );
  AND U12848 ( .A(p_input[2528]), .B(n13103), .Z(n13099) );
  IV U12849 ( .A(p_input[2496]), .Z(n13103) );
  XNOR U12850 ( .A(p_input[2432]), .B(n13104), .Z(n12697) );
  AND U12851 ( .A(n268), .B(n13105), .Z(n13104) );
  XOR U12852 ( .A(p_input[2464]), .B(p_input[2432]), .Z(n13105) );
  XOR U12853 ( .A(n13106), .B(n13107), .Z(n268) );
  AND U12854 ( .A(n13108), .B(n13109), .Z(n13107) );
  XNOR U12855 ( .A(p_input[2495]), .B(n13106), .Z(n13109) );
  XOR U12856 ( .A(n13106), .B(p_input[2463]), .Z(n13108) );
  XOR U12857 ( .A(n13110), .B(n13111), .Z(n13106) );
  AND U12858 ( .A(n13112), .B(n13113), .Z(n13111) );
  XNOR U12859 ( .A(p_input[2494]), .B(n13110), .Z(n13113) );
  XNOR U12860 ( .A(n13110), .B(n12712), .Z(n13112) );
  IV U12861 ( .A(p_input[2462]), .Z(n12712) );
  XOR U12862 ( .A(n13114), .B(n13115), .Z(n13110) );
  AND U12863 ( .A(n13116), .B(n13117), .Z(n13115) );
  XNOR U12864 ( .A(p_input[2493]), .B(n13114), .Z(n13117) );
  XNOR U12865 ( .A(n13114), .B(n12721), .Z(n13116) );
  IV U12866 ( .A(p_input[2461]), .Z(n12721) );
  XOR U12867 ( .A(n13118), .B(n13119), .Z(n13114) );
  AND U12868 ( .A(n13120), .B(n13121), .Z(n13119) );
  XNOR U12869 ( .A(p_input[2492]), .B(n13118), .Z(n13121) );
  XNOR U12870 ( .A(n13118), .B(n12730), .Z(n13120) );
  IV U12871 ( .A(p_input[2460]), .Z(n12730) );
  XOR U12872 ( .A(n13122), .B(n13123), .Z(n13118) );
  AND U12873 ( .A(n13124), .B(n13125), .Z(n13123) );
  XNOR U12874 ( .A(p_input[2491]), .B(n13122), .Z(n13125) );
  XNOR U12875 ( .A(n13122), .B(n12739), .Z(n13124) );
  IV U12876 ( .A(p_input[2459]), .Z(n12739) );
  XOR U12877 ( .A(n13126), .B(n13127), .Z(n13122) );
  AND U12878 ( .A(n13128), .B(n13129), .Z(n13127) );
  XNOR U12879 ( .A(p_input[2490]), .B(n13126), .Z(n13129) );
  XNOR U12880 ( .A(n13126), .B(n12748), .Z(n13128) );
  IV U12881 ( .A(p_input[2458]), .Z(n12748) );
  XOR U12882 ( .A(n13130), .B(n13131), .Z(n13126) );
  AND U12883 ( .A(n13132), .B(n13133), .Z(n13131) );
  XNOR U12884 ( .A(p_input[2489]), .B(n13130), .Z(n13133) );
  XNOR U12885 ( .A(n13130), .B(n12757), .Z(n13132) );
  IV U12886 ( .A(p_input[2457]), .Z(n12757) );
  XOR U12887 ( .A(n13134), .B(n13135), .Z(n13130) );
  AND U12888 ( .A(n13136), .B(n13137), .Z(n13135) );
  XNOR U12889 ( .A(p_input[2488]), .B(n13134), .Z(n13137) );
  XNOR U12890 ( .A(n13134), .B(n12766), .Z(n13136) );
  IV U12891 ( .A(p_input[2456]), .Z(n12766) );
  XOR U12892 ( .A(n13138), .B(n13139), .Z(n13134) );
  AND U12893 ( .A(n13140), .B(n13141), .Z(n13139) );
  XNOR U12894 ( .A(p_input[2487]), .B(n13138), .Z(n13141) );
  XNOR U12895 ( .A(n13138), .B(n12775), .Z(n13140) );
  IV U12896 ( .A(p_input[2455]), .Z(n12775) );
  XOR U12897 ( .A(n13142), .B(n13143), .Z(n13138) );
  AND U12898 ( .A(n13144), .B(n13145), .Z(n13143) );
  XNOR U12899 ( .A(p_input[2486]), .B(n13142), .Z(n13145) );
  XNOR U12900 ( .A(n13142), .B(n12784), .Z(n13144) );
  IV U12901 ( .A(p_input[2454]), .Z(n12784) );
  XOR U12902 ( .A(n13146), .B(n13147), .Z(n13142) );
  AND U12903 ( .A(n13148), .B(n13149), .Z(n13147) );
  XNOR U12904 ( .A(p_input[2485]), .B(n13146), .Z(n13149) );
  XNOR U12905 ( .A(n13146), .B(n12793), .Z(n13148) );
  IV U12906 ( .A(p_input[2453]), .Z(n12793) );
  XOR U12907 ( .A(n13150), .B(n13151), .Z(n13146) );
  AND U12908 ( .A(n13152), .B(n13153), .Z(n13151) );
  XNOR U12909 ( .A(p_input[2484]), .B(n13150), .Z(n13153) );
  XNOR U12910 ( .A(n13150), .B(n12802), .Z(n13152) );
  IV U12911 ( .A(p_input[2452]), .Z(n12802) );
  XOR U12912 ( .A(n13154), .B(n13155), .Z(n13150) );
  AND U12913 ( .A(n13156), .B(n13157), .Z(n13155) );
  XNOR U12914 ( .A(p_input[2483]), .B(n13154), .Z(n13157) );
  XNOR U12915 ( .A(n13154), .B(n12811), .Z(n13156) );
  IV U12916 ( .A(p_input[2451]), .Z(n12811) );
  XOR U12917 ( .A(n13158), .B(n13159), .Z(n13154) );
  AND U12918 ( .A(n13160), .B(n13161), .Z(n13159) );
  XNOR U12919 ( .A(p_input[2482]), .B(n13158), .Z(n13161) );
  XNOR U12920 ( .A(n13158), .B(n12820), .Z(n13160) );
  IV U12921 ( .A(p_input[2450]), .Z(n12820) );
  XOR U12922 ( .A(n13162), .B(n13163), .Z(n13158) );
  AND U12923 ( .A(n13164), .B(n13165), .Z(n13163) );
  XNOR U12924 ( .A(p_input[2481]), .B(n13162), .Z(n13165) );
  XNOR U12925 ( .A(n13162), .B(n12829), .Z(n13164) );
  IV U12926 ( .A(p_input[2449]), .Z(n12829) );
  XOR U12927 ( .A(n13166), .B(n13167), .Z(n13162) );
  AND U12928 ( .A(n13168), .B(n13169), .Z(n13167) );
  XNOR U12929 ( .A(p_input[2480]), .B(n13166), .Z(n13169) );
  XNOR U12930 ( .A(n13166), .B(n12838), .Z(n13168) );
  IV U12931 ( .A(p_input[2448]), .Z(n12838) );
  XOR U12932 ( .A(n13170), .B(n13171), .Z(n13166) );
  AND U12933 ( .A(n13172), .B(n13173), .Z(n13171) );
  XNOR U12934 ( .A(p_input[2479]), .B(n13170), .Z(n13173) );
  XNOR U12935 ( .A(n13170), .B(n12847), .Z(n13172) );
  IV U12936 ( .A(p_input[2447]), .Z(n12847) );
  XOR U12937 ( .A(n13174), .B(n13175), .Z(n13170) );
  AND U12938 ( .A(n13176), .B(n13177), .Z(n13175) );
  XNOR U12939 ( .A(p_input[2478]), .B(n13174), .Z(n13177) );
  XNOR U12940 ( .A(n13174), .B(n12856), .Z(n13176) );
  IV U12941 ( .A(p_input[2446]), .Z(n12856) );
  XOR U12942 ( .A(n13178), .B(n13179), .Z(n13174) );
  AND U12943 ( .A(n13180), .B(n13181), .Z(n13179) );
  XNOR U12944 ( .A(p_input[2477]), .B(n13178), .Z(n13181) );
  XNOR U12945 ( .A(n13178), .B(n12865), .Z(n13180) );
  IV U12946 ( .A(p_input[2445]), .Z(n12865) );
  XOR U12947 ( .A(n13182), .B(n13183), .Z(n13178) );
  AND U12948 ( .A(n13184), .B(n13185), .Z(n13183) );
  XNOR U12949 ( .A(p_input[2476]), .B(n13182), .Z(n13185) );
  XNOR U12950 ( .A(n13182), .B(n12874), .Z(n13184) );
  IV U12951 ( .A(p_input[2444]), .Z(n12874) );
  XOR U12952 ( .A(n13186), .B(n13187), .Z(n13182) );
  AND U12953 ( .A(n13188), .B(n13189), .Z(n13187) );
  XNOR U12954 ( .A(p_input[2475]), .B(n13186), .Z(n13189) );
  XNOR U12955 ( .A(n13186), .B(n12883), .Z(n13188) );
  IV U12956 ( .A(p_input[2443]), .Z(n12883) );
  XOR U12957 ( .A(n13190), .B(n13191), .Z(n13186) );
  AND U12958 ( .A(n13192), .B(n13193), .Z(n13191) );
  XNOR U12959 ( .A(p_input[2474]), .B(n13190), .Z(n13193) );
  XNOR U12960 ( .A(n13190), .B(n12892), .Z(n13192) );
  IV U12961 ( .A(p_input[2442]), .Z(n12892) );
  XOR U12962 ( .A(n13194), .B(n13195), .Z(n13190) );
  AND U12963 ( .A(n13196), .B(n13197), .Z(n13195) );
  XNOR U12964 ( .A(p_input[2473]), .B(n13194), .Z(n13197) );
  XNOR U12965 ( .A(n13194), .B(n12901), .Z(n13196) );
  IV U12966 ( .A(p_input[2441]), .Z(n12901) );
  XOR U12967 ( .A(n13198), .B(n13199), .Z(n13194) );
  AND U12968 ( .A(n13200), .B(n13201), .Z(n13199) );
  XNOR U12969 ( .A(p_input[2472]), .B(n13198), .Z(n13201) );
  XNOR U12970 ( .A(n13198), .B(n12910), .Z(n13200) );
  IV U12971 ( .A(p_input[2440]), .Z(n12910) );
  XOR U12972 ( .A(n13202), .B(n13203), .Z(n13198) );
  AND U12973 ( .A(n13204), .B(n13205), .Z(n13203) );
  XNOR U12974 ( .A(p_input[2471]), .B(n13202), .Z(n13205) );
  XNOR U12975 ( .A(n13202), .B(n12919), .Z(n13204) );
  IV U12976 ( .A(p_input[2439]), .Z(n12919) );
  XOR U12977 ( .A(n13206), .B(n13207), .Z(n13202) );
  AND U12978 ( .A(n13208), .B(n13209), .Z(n13207) );
  XNOR U12979 ( .A(p_input[2470]), .B(n13206), .Z(n13209) );
  XNOR U12980 ( .A(n13206), .B(n12928), .Z(n13208) );
  IV U12981 ( .A(p_input[2438]), .Z(n12928) );
  XOR U12982 ( .A(n13210), .B(n13211), .Z(n13206) );
  AND U12983 ( .A(n13212), .B(n13213), .Z(n13211) );
  XNOR U12984 ( .A(p_input[2469]), .B(n13210), .Z(n13213) );
  XNOR U12985 ( .A(n13210), .B(n12937), .Z(n13212) );
  IV U12986 ( .A(p_input[2437]), .Z(n12937) );
  XOR U12987 ( .A(n13214), .B(n13215), .Z(n13210) );
  AND U12988 ( .A(n13216), .B(n13217), .Z(n13215) );
  XNOR U12989 ( .A(p_input[2468]), .B(n13214), .Z(n13217) );
  XNOR U12990 ( .A(n13214), .B(n12946), .Z(n13216) );
  IV U12991 ( .A(p_input[2436]), .Z(n12946) );
  XOR U12992 ( .A(n13218), .B(n13219), .Z(n13214) );
  AND U12993 ( .A(n13220), .B(n13221), .Z(n13219) );
  XNOR U12994 ( .A(p_input[2467]), .B(n13218), .Z(n13221) );
  XNOR U12995 ( .A(n13218), .B(n12955), .Z(n13220) );
  IV U12996 ( .A(p_input[2435]), .Z(n12955) );
  XOR U12997 ( .A(n13222), .B(n13223), .Z(n13218) );
  AND U12998 ( .A(n13224), .B(n13225), .Z(n13223) );
  XNOR U12999 ( .A(p_input[2466]), .B(n13222), .Z(n13225) );
  XNOR U13000 ( .A(n13222), .B(n12964), .Z(n13224) );
  IV U13001 ( .A(p_input[2434]), .Z(n12964) );
  XNOR U13002 ( .A(n13226), .B(n13227), .Z(n13222) );
  AND U13003 ( .A(n13228), .B(n13229), .Z(n13227) );
  XOR U13004 ( .A(p_input[2465]), .B(n13226), .Z(n13229) );
  XNOR U13005 ( .A(p_input[2433]), .B(n13226), .Z(n13228) );
  AND U13006 ( .A(p_input[2464]), .B(n13230), .Z(n13226) );
  IV U13007 ( .A(p_input[2432]), .Z(n13230) );
  XOR U13008 ( .A(n13231), .B(n13232), .Z(n12320) );
  AND U13009 ( .A(n344), .B(n13233), .Z(n13232) );
  XNOR U13010 ( .A(n13234), .B(n13231), .Z(n13233) );
  XOR U13011 ( .A(n13235), .B(n13236), .Z(n344) );
  AND U13012 ( .A(n13237), .B(n13238), .Z(n13236) );
  XNOR U13013 ( .A(n12335), .B(n13235), .Z(n13238) );
  AND U13014 ( .A(p_input[2431]), .B(p_input[2399]), .Z(n12335) );
  XNOR U13015 ( .A(n13235), .B(n12332), .Z(n13237) );
  IV U13016 ( .A(n13239), .Z(n12332) );
  AND U13017 ( .A(p_input[2335]), .B(p_input[2367]), .Z(n13239) );
  XOR U13018 ( .A(n13240), .B(n13241), .Z(n13235) );
  AND U13019 ( .A(n13242), .B(n13243), .Z(n13241) );
  XOR U13020 ( .A(n13240), .B(n12347), .Z(n13243) );
  XNOR U13021 ( .A(p_input[2398]), .B(n13244), .Z(n12347) );
  AND U13022 ( .A(n274), .B(n13245), .Z(n13244) );
  XOR U13023 ( .A(p_input[2430]), .B(p_input[2398]), .Z(n13245) );
  XNOR U13024 ( .A(n12344), .B(n13240), .Z(n13242) );
  XOR U13025 ( .A(n13246), .B(n13247), .Z(n12344) );
  AND U13026 ( .A(n271), .B(n13248), .Z(n13247) );
  XOR U13027 ( .A(p_input[2366]), .B(p_input[2334]), .Z(n13248) );
  XOR U13028 ( .A(n13249), .B(n13250), .Z(n13240) );
  AND U13029 ( .A(n13251), .B(n13252), .Z(n13250) );
  XOR U13030 ( .A(n13249), .B(n12359), .Z(n13252) );
  XNOR U13031 ( .A(p_input[2397]), .B(n13253), .Z(n12359) );
  AND U13032 ( .A(n274), .B(n13254), .Z(n13253) );
  XOR U13033 ( .A(p_input[2429]), .B(p_input[2397]), .Z(n13254) );
  XNOR U13034 ( .A(n12356), .B(n13249), .Z(n13251) );
  XOR U13035 ( .A(n13255), .B(n13256), .Z(n12356) );
  AND U13036 ( .A(n271), .B(n13257), .Z(n13256) );
  XOR U13037 ( .A(p_input[2365]), .B(p_input[2333]), .Z(n13257) );
  XOR U13038 ( .A(n13258), .B(n13259), .Z(n13249) );
  AND U13039 ( .A(n13260), .B(n13261), .Z(n13259) );
  XOR U13040 ( .A(n13258), .B(n12371), .Z(n13261) );
  XNOR U13041 ( .A(p_input[2396]), .B(n13262), .Z(n12371) );
  AND U13042 ( .A(n274), .B(n13263), .Z(n13262) );
  XOR U13043 ( .A(p_input[2428]), .B(p_input[2396]), .Z(n13263) );
  XNOR U13044 ( .A(n12368), .B(n13258), .Z(n13260) );
  XOR U13045 ( .A(n13264), .B(n13265), .Z(n12368) );
  AND U13046 ( .A(n271), .B(n13266), .Z(n13265) );
  XOR U13047 ( .A(p_input[2364]), .B(p_input[2332]), .Z(n13266) );
  XOR U13048 ( .A(n13267), .B(n13268), .Z(n13258) );
  AND U13049 ( .A(n13269), .B(n13270), .Z(n13268) );
  XOR U13050 ( .A(n13267), .B(n12383), .Z(n13270) );
  XNOR U13051 ( .A(p_input[2395]), .B(n13271), .Z(n12383) );
  AND U13052 ( .A(n274), .B(n13272), .Z(n13271) );
  XOR U13053 ( .A(p_input[2427]), .B(p_input[2395]), .Z(n13272) );
  XNOR U13054 ( .A(n12380), .B(n13267), .Z(n13269) );
  XOR U13055 ( .A(n13273), .B(n13274), .Z(n12380) );
  AND U13056 ( .A(n271), .B(n13275), .Z(n13274) );
  XOR U13057 ( .A(p_input[2363]), .B(p_input[2331]), .Z(n13275) );
  XOR U13058 ( .A(n13276), .B(n13277), .Z(n13267) );
  AND U13059 ( .A(n13278), .B(n13279), .Z(n13277) );
  XOR U13060 ( .A(n13276), .B(n12395), .Z(n13279) );
  XNOR U13061 ( .A(p_input[2394]), .B(n13280), .Z(n12395) );
  AND U13062 ( .A(n274), .B(n13281), .Z(n13280) );
  XOR U13063 ( .A(p_input[2426]), .B(p_input[2394]), .Z(n13281) );
  XNOR U13064 ( .A(n12392), .B(n13276), .Z(n13278) );
  XOR U13065 ( .A(n13282), .B(n13283), .Z(n12392) );
  AND U13066 ( .A(n271), .B(n13284), .Z(n13283) );
  XOR U13067 ( .A(p_input[2362]), .B(p_input[2330]), .Z(n13284) );
  XOR U13068 ( .A(n13285), .B(n13286), .Z(n13276) );
  AND U13069 ( .A(n13287), .B(n13288), .Z(n13286) );
  XOR U13070 ( .A(n13285), .B(n12407), .Z(n13288) );
  XNOR U13071 ( .A(p_input[2393]), .B(n13289), .Z(n12407) );
  AND U13072 ( .A(n274), .B(n13290), .Z(n13289) );
  XOR U13073 ( .A(p_input[2425]), .B(p_input[2393]), .Z(n13290) );
  XNOR U13074 ( .A(n12404), .B(n13285), .Z(n13287) );
  XOR U13075 ( .A(n13291), .B(n13292), .Z(n12404) );
  AND U13076 ( .A(n271), .B(n13293), .Z(n13292) );
  XOR U13077 ( .A(p_input[2361]), .B(p_input[2329]), .Z(n13293) );
  XOR U13078 ( .A(n13294), .B(n13295), .Z(n13285) );
  AND U13079 ( .A(n13296), .B(n13297), .Z(n13295) );
  XOR U13080 ( .A(n13294), .B(n12419), .Z(n13297) );
  XNOR U13081 ( .A(p_input[2392]), .B(n13298), .Z(n12419) );
  AND U13082 ( .A(n274), .B(n13299), .Z(n13298) );
  XOR U13083 ( .A(p_input[2424]), .B(p_input[2392]), .Z(n13299) );
  XNOR U13084 ( .A(n12416), .B(n13294), .Z(n13296) );
  XOR U13085 ( .A(n13300), .B(n13301), .Z(n12416) );
  AND U13086 ( .A(n271), .B(n13302), .Z(n13301) );
  XOR U13087 ( .A(p_input[2360]), .B(p_input[2328]), .Z(n13302) );
  XOR U13088 ( .A(n13303), .B(n13304), .Z(n13294) );
  AND U13089 ( .A(n13305), .B(n13306), .Z(n13304) );
  XOR U13090 ( .A(n13303), .B(n12431), .Z(n13306) );
  XNOR U13091 ( .A(p_input[2391]), .B(n13307), .Z(n12431) );
  AND U13092 ( .A(n274), .B(n13308), .Z(n13307) );
  XOR U13093 ( .A(p_input[2423]), .B(p_input[2391]), .Z(n13308) );
  XNOR U13094 ( .A(n12428), .B(n13303), .Z(n13305) );
  XOR U13095 ( .A(n13309), .B(n13310), .Z(n12428) );
  AND U13096 ( .A(n271), .B(n13311), .Z(n13310) );
  XOR U13097 ( .A(p_input[2359]), .B(p_input[2327]), .Z(n13311) );
  XOR U13098 ( .A(n13312), .B(n13313), .Z(n13303) );
  AND U13099 ( .A(n13314), .B(n13315), .Z(n13313) );
  XOR U13100 ( .A(n13312), .B(n12443), .Z(n13315) );
  XNOR U13101 ( .A(p_input[2390]), .B(n13316), .Z(n12443) );
  AND U13102 ( .A(n274), .B(n13317), .Z(n13316) );
  XOR U13103 ( .A(p_input[2422]), .B(p_input[2390]), .Z(n13317) );
  XNOR U13104 ( .A(n12440), .B(n13312), .Z(n13314) );
  XOR U13105 ( .A(n13318), .B(n13319), .Z(n12440) );
  AND U13106 ( .A(n271), .B(n13320), .Z(n13319) );
  XOR U13107 ( .A(p_input[2358]), .B(p_input[2326]), .Z(n13320) );
  XOR U13108 ( .A(n13321), .B(n13322), .Z(n13312) );
  AND U13109 ( .A(n13323), .B(n13324), .Z(n13322) );
  XOR U13110 ( .A(n13321), .B(n12455), .Z(n13324) );
  XNOR U13111 ( .A(p_input[2389]), .B(n13325), .Z(n12455) );
  AND U13112 ( .A(n274), .B(n13326), .Z(n13325) );
  XOR U13113 ( .A(p_input[2421]), .B(p_input[2389]), .Z(n13326) );
  XNOR U13114 ( .A(n12452), .B(n13321), .Z(n13323) );
  XOR U13115 ( .A(n13327), .B(n13328), .Z(n12452) );
  AND U13116 ( .A(n271), .B(n13329), .Z(n13328) );
  XOR U13117 ( .A(p_input[2357]), .B(p_input[2325]), .Z(n13329) );
  XOR U13118 ( .A(n13330), .B(n13331), .Z(n13321) );
  AND U13119 ( .A(n13332), .B(n13333), .Z(n13331) );
  XOR U13120 ( .A(n13330), .B(n12467), .Z(n13333) );
  XNOR U13121 ( .A(p_input[2388]), .B(n13334), .Z(n12467) );
  AND U13122 ( .A(n274), .B(n13335), .Z(n13334) );
  XOR U13123 ( .A(p_input[2420]), .B(p_input[2388]), .Z(n13335) );
  XNOR U13124 ( .A(n12464), .B(n13330), .Z(n13332) );
  XOR U13125 ( .A(n13336), .B(n13337), .Z(n12464) );
  AND U13126 ( .A(n271), .B(n13338), .Z(n13337) );
  XOR U13127 ( .A(p_input[2356]), .B(p_input[2324]), .Z(n13338) );
  XOR U13128 ( .A(n13339), .B(n13340), .Z(n13330) );
  AND U13129 ( .A(n13341), .B(n13342), .Z(n13340) );
  XOR U13130 ( .A(n13339), .B(n12479), .Z(n13342) );
  XNOR U13131 ( .A(p_input[2387]), .B(n13343), .Z(n12479) );
  AND U13132 ( .A(n274), .B(n13344), .Z(n13343) );
  XOR U13133 ( .A(p_input[2419]), .B(p_input[2387]), .Z(n13344) );
  XNOR U13134 ( .A(n12476), .B(n13339), .Z(n13341) );
  XOR U13135 ( .A(n13345), .B(n13346), .Z(n12476) );
  AND U13136 ( .A(n271), .B(n13347), .Z(n13346) );
  XOR U13137 ( .A(p_input[2355]), .B(p_input[2323]), .Z(n13347) );
  XOR U13138 ( .A(n13348), .B(n13349), .Z(n13339) );
  AND U13139 ( .A(n13350), .B(n13351), .Z(n13349) );
  XOR U13140 ( .A(n13348), .B(n12491), .Z(n13351) );
  XNOR U13141 ( .A(p_input[2386]), .B(n13352), .Z(n12491) );
  AND U13142 ( .A(n274), .B(n13353), .Z(n13352) );
  XOR U13143 ( .A(p_input[2418]), .B(p_input[2386]), .Z(n13353) );
  XNOR U13144 ( .A(n12488), .B(n13348), .Z(n13350) );
  XOR U13145 ( .A(n13354), .B(n13355), .Z(n12488) );
  AND U13146 ( .A(n271), .B(n13356), .Z(n13355) );
  XOR U13147 ( .A(p_input[2354]), .B(p_input[2322]), .Z(n13356) );
  XOR U13148 ( .A(n13357), .B(n13358), .Z(n13348) );
  AND U13149 ( .A(n13359), .B(n13360), .Z(n13358) );
  XOR U13150 ( .A(n13357), .B(n12503), .Z(n13360) );
  XNOR U13151 ( .A(p_input[2385]), .B(n13361), .Z(n12503) );
  AND U13152 ( .A(n274), .B(n13362), .Z(n13361) );
  XOR U13153 ( .A(p_input[2417]), .B(p_input[2385]), .Z(n13362) );
  XNOR U13154 ( .A(n12500), .B(n13357), .Z(n13359) );
  XOR U13155 ( .A(n13363), .B(n13364), .Z(n12500) );
  AND U13156 ( .A(n271), .B(n13365), .Z(n13364) );
  XOR U13157 ( .A(p_input[2353]), .B(p_input[2321]), .Z(n13365) );
  XOR U13158 ( .A(n13366), .B(n13367), .Z(n13357) );
  AND U13159 ( .A(n13368), .B(n13369), .Z(n13367) );
  XOR U13160 ( .A(n13366), .B(n12515), .Z(n13369) );
  XNOR U13161 ( .A(p_input[2384]), .B(n13370), .Z(n12515) );
  AND U13162 ( .A(n274), .B(n13371), .Z(n13370) );
  XOR U13163 ( .A(p_input[2416]), .B(p_input[2384]), .Z(n13371) );
  XNOR U13164 ( .A(n12512), .B(n13366), .Z(n13368) );
  XOR U13165 ( .A(n13372), .B(n13373), .Z(n12512) );
  AND U13166 ( .A(n271), .B(n13374), .Z(n13373) );
  XOR U13167 ( .A(p_input[2352]), .B(p_input[2320]), .Z(n13374) );
  XOR U13168 ( .A(n13375), .B(n13376), .Z(n13366) );
  AND U13169 ( .A(n13377), .B(n13378), .Z(n13376) );
  XOR U13170 ( .A(n13375), .B(n12527), .Z(n13378) );
  XNOR U13171 ( .A(p_input[2383]), .B(n13379), .Z(n12527) );
  AND U13172 ( .A(n274), .B(n13380), .Z(n13379) );
  XOR U13173 ( .A(p_input[2415]), .B(p_input[2383]), .Z(n13380) );
  XNOR U13174 ( .A(n12524), .B(n13375), .Z(n13377) );
  XOR U13175 ( .A(n13381), .B(n13382), .Z(n12524) );
  AND U13176 ( .A(n271), .B(n13383), .Z(n13382) );
  XOR U13177 ( .A(p_input[2351]), .B(p_input[2319]), .Z(n13383) );
  XOR U13178 ( .A(n13384), .B(n13385), .Z(n13375) );
  AND U13179 ( .A(n13386), .B(n13387), .Z(n13385) );
  XOR U13180 ( .A(n13384), .B(n12539), .Z(n13387) );
  XNOR U13181 ( .A(p_input[2382]), .B(n13388), .Z(n12539) );
  AND U13182 ( .A(n274), .B(n13389), .Z(n13388) );
  XOR U13183 ( .A(p_input[2414]), .B(p_input[2382]), .Z(n13389) );
  XNOR U13184 ( .A(n12536), .B(n13384), .Z(n13386) );
  XOR U13185 ( .A(n13390), .B(n13391), .Z(n12536) );
  AND U13186 ( .A(n271), .B(n13392), .Z(n13391) );
  XOR U13187 ( .A(p_input[2350]), .B(p_input[2318]), .Z(n13392) );
  XOR U13188 ( .A(n13393), .B(n13394), .Z(n13384) );
  AND U13189 ( .A(n13395), .B(n13396), .Z(n13394) );
  XOR U13190 ( .A(n13393), .B(n12551), .Z(n13396) );
  XNOR U13191 ( .A(p_input[2381]), .B(n13397), .Z(n12551) );
  AND U13192 ( .A(n274), .B(n13398), .Z(n13397) );
  XOR U13193 ( .A(p_input[2413]), .B(p_input[2381]), .Z(n13398) );
  XNOR U13194 ( .A(n12548), .B(n13393), .Z(n13395) );
  XOR U13195 ( .A(n13399), .B(n13400), .Z(n12548) );
  AND U13196 ( .A(n271), .B(n13401), .Z(n13400) );
  XOR U13197 ( .A(p_input[2349]), .B(p_input[2317]), .Z(n13401) );
  XOR U13198 ( .A(n13402), .B(n13403), .Z(n13393) );
  AND U13199 ( .A(n13404), .B(n13405), .Z(n13403) );
  XOR U13200 ( .A(n13402), .B(n12563), .Z(n13405) );
  XNOR U13201 ( .A(p_input[2380]), .B(n13406), .Z(n12563) );
  AND U13202 ( .A(n274), .B(n13407), .Z(n13406) );
  XOR U13203 ( .A(p_input[2412]), .B(p_input[2380]), .Z(n13407) );
  XNOR U13204 ( .A(n12560), .B(n13402), .Z(n13404) );
  XOR U13205 ( .A(n13408), .B(n13409), .Z(n12560) );
  AND U13206 ( .A(n271), .B(n13410), .Z(n13409) );
  XOR U13207 ( .A(p_input[2348]), .B(p_input[2316]), .Z(n13410) );
  XOR U13208 ( .A(n13411), .B(n13412), .Z(n13402) );
  AND U13209 ( .A(n13413), .B(n13414), .Z(n13412) );
  XOR U13210 ( .A(n13411), .B(n12575), .Z(n13414) );
  XNOR U13211 ( .A(p_input[2379]), .B(n13415), .Z(n12575) );
  AND U13212 ( .A(n274), .B(n13416), .Z(n13415) );
  XOR U13213 ( .A(p_input[2411]), .B(p_input[2379]), .Z(n13416) );
  XNOR U13214 ( .A(n12572), .B(n13411), .Z(n13413) );
  XOR U13215 ( .A(n13417), .B(n13418), .Z(n12572) );
  AND U13216 ( .A(n271), .B(n13419), .Z(n13418) );
  XOR U13217 ( .A(p_input[2347]), .B(p_input[2315]), .Z(n13419) );
  XOR U13218 ( .A(n13420), .B(n13421), .Z(n13411) );
  AND U13219 ( .A(n13422), .B(n13423), .Z(n13421) );
  XOR U13220 ( .A(n13420), .B(n12587), .Z(n13423) );
  XNOR U13221 ( .A(p_input[2378]), .B(n13424), .Z(n12587) );
  AND U13222 ( .A(n274), .B(n13425), .Z(n13424) );
  XOR U13223 ( .A(p_input[2410]), .B(p_input[2378]), .Z(n13425) );
  XNOR U13224 ( .A(n12584), .B(n13420), .Z(n13422) );
  XOR U13225 ( .A(n13426), .B(n13427), .Z(n12584) );
  AND U13226 ( .A(n271), .B(n13428), .Z(n13427) );
  XOR U13227 ( .A(p_input[2346]), .B(p_input[2314]), .Z(n13428) );
  XOR U13228 ( .A(n13429), .B(n13430), .Z(n13420) );
  AND U13229 ( .A(n13431), .B(n13432), .Z(n13430) );
  XOR U13230 ( .A(n13429), .B(n12599), .Z(n13432) );
  XNOR U13231 ( .A(p_input[2377]), .B(n13433), .Z(n12599) );
  AND U13232 ( .A(n274), .B(n13434), .Z(n13433) );
  XOR U13233 ( .A(p_input[2409]), .B(p_input[2377]), .Z(n13434) );
  XNOR U13234 ( .A(n12596), .B(n13429), .Z(n13431) );
  XOR U13235 ( .A(n13435), .B(n13436), .Z(n12596) );
  AND U13236 ( .A(n271), .B(n13437), .Z(n13436) );
  XOR U13237 ( .A(p_input[2345]), .B(p_input[2313]), .Z(n13437) );
  XOR U13238 ( .A(n13438), .B(n13439), .Z(n13429) );
  AND U13239 ( .A(n13440), .B(n13441), .Z(n13439) );
  XOR U13240 ( .A(n13438), .B(n12611), .Z(n13441) );
  XNOR U13241 ( .A(p_input[2376]), .B(n13442), .Z(n12611) );
  AND U13242 ( .A(n274), .B(n13443), .Z(n13442) );
  XOR U13243 ( .A(p_input[2408]), .B(p_input[2376]), .Z(n13443) );
  XNOR U13244 ( .A(n12608), .B(n13438), .Z(n13440) );
  XOR U13245 ( .A(n13444), .B(n13445), .Z(n12608) );
  AND U13246 ( .A(n271), .B(n13446), .Z(n13445) );
  XOR U13247 ( .A(p_input[2344]), .B(p_input[2312]), .Z(n13446) );
  XOR U13248 ( .A(n13447), .B(n13448), .Z(n13438) );
  AND U13249 ( .A(n13449), .B(n13450), .Z(n13448) );
  XOR U13250 ( .A(n13447), .B(n12623), .Z(n13450) );
  XNOR U13251 ( .A(p_input[2375]), .B(n13451), .Z(n12623) );
  AND U13252 ( .A(n274), .B(n13452), .Z(n13451) );
  XOR U13253 ( .A(p_input[2407]), .B(p_input[2375]), .Z(n13452) );
  XNOR U13254 ( .A(n12620), .B(n13447), .Z(n13449) );
  XOR U13255 ( .A(n13453), .B(n13454), .Z(n12620) );
  AND U13256 ( .A(n271), .B(n13455), .Z(n13454) );
  XOR U13257 ( .A(p_input[2343]), .B(p_input[2311]), .Z(n13455) );
  XOR U13258 ( .A(n13456), .B(n13457), .Z(n13447) );
  AND U13259 ( .A(n13458), .B(n13459), .Z(n13457) );
  XOR U13260 ( .A(n13456), .B(n12635), .Z(n13459) );
  XNOR U13261 ( .A(p_input[2374]), .B(n13460), .Z(n12635) );
  AND U13262 ( .A(n274), .B(n13461), .Z(n13460) );
  XOR U13263 ( .A(p_input[2406]), .B(p_input[2374]), .Z(n13461) );
  XNOR U13264 ( .A(n12632), .B(n13456), .Z(n13458) );
  XOR U13265 ( .A(n13462), .B(n13463), .Z(n12632) );
  AND U13266 ( .A(n271), .B(n13464), .Z(n13463) );
  XOR U13267 ( .A(p_input[2342]), .B(p_input[2310]), .Z(n13464) );
  XOR U13268 ( .A(n13465), .B(n13466), .Z(n13456) );
  AND U13269 ( .A(n13467), .B(n13468), .Z(n13466) );
  XOR U13270 ( .A(n13465), .B(n12647), .Z(n13468) );
  XNOR U13271 ( .A(p_input[2373]), .B(n13469), .Z(n12647) );
  AND U13272 ( .A(n274), .B(n13470), .Z(n13469) );
  XOR U13273 ( .A(p_input[2405]), .B(p_input[2373]), .Z(n13470) );
  XNOR U13274 ( .A(n12644), .B(n13465), .Z(n13467) );
  XOR U13275 ( .A(n13471), .B(n13472), .Z(n12644) );
  AND U13276 ( .A(n271), .B(n13473), .Z(n13472) );
  XOR U13277 ( .A(p_input[2341]), .B(p_input[2309]), .Z(n13473) );
  XOR U13278 ( .A(n13474), .B(n13475), .Z(n13465) );
  AND U13279 ( .A(n13476), .B(n13477), .Z(n13475) );
  XOR U13280 ( .A(n13474), .B(n12659), .Z(n13477) );
  XNOR U13281 ( .A(p_input[2372]), .B(n13478), .Z(n12659) );
  AND U13282 ( .A(n274), .B(n13479), .Z(n13478) );
  XOR U13283 ( .A(p_input[2404]), .B(p_input[2372]), .Z(n13479) );
  XNOR U13284 ( .A(n12656), .B(n13474), .Z(n13476) );
  XOR U13285 ( .A(n13480), .B(n13481), .Z(n12656) );
  AND U13286 ( .A(n271), .B(n13482), .Z(n13481) );
  XOR U13287 ( .A(p_input[2340]), .B(p_input[2308]), .Z(n13482) );
  XOR U13288 ( .A(n13483), .B(n13484), .Z(n13474) );
  AND U13289 ( .A(n13485), .B(n13486), .Z(n13484) );
  XOR U13290 ( .A(n13483), .B(n12671), .Z(n13486) );
  XNOR U13291 ( .A(p_input[2371]), .B(n13487), .Z(n12671) );
  AND U13292 ( .A(n274), .B(n13488), .Z(n13487) );
  XOR U13293 ( .A(p_input[2403]), .B(p_input[2371]), .Z(n13488) );
  XNOR U13294 ( .A(n12668), .B(n13483), .Z(n13485) );
  XOR U13295 ( .A(n13489), .B(n13490), .Z(n12668) );
  AND U13296 ( .A(n271), .B(n13491), .Z(n13490) );
  XOR U13297 ( .A(p_input[2339]), .B(p_input[2307]), .Z(n13491) );
  XOR U13298 ( .A(n13492), .B(n13493), .Z(n13483) );
  AND U13299 ( .A(n13494), .B(n13495), .Z(n13493) );
  XOR U13300 ( .A(n12683), .B(n13492), .Z(n13495) );
  XNOR U13301 ( .A(p_input[2370]), .B(n13496), .Z(n12683) );
  AND U13302 ( .A(n274), .B(n13497), .Z(n13496) );
  XOR U13303 ( .A(p_input[2402]), .B(p_input[2370]), .Z(n13497) );
  XNOR U13304 ( .A(n13492), .B(n12680), .Z(n13494) );
  XOR U13305 ( .A(n13498), .B(n13499), .Z(n12680) );
  AND U13306 ( .A(n271), .B(n13500), .Z(n13499) );
  XOR U13307 ( .A(p_input[2338]), .B(p_input[2306]), .Z(n13500) );
  XOR U13308 ( .A(n13501), .B(n13502), .Z(n13492) );
  AND U13309 ( .A(n13503), .B(n13504), .Z(n13502) );
  XNOR U13310 ( .A(n13505), .B(n12696), .Z(n13504) );
  XNOR U13311 ( .A(p_input[2369]), .B(n13506), .Z(n12696) );
  AND U13312 ( .A(n274), .B(n13507), .Z(n13506) );
  XNOR U13313 ( .A(p_input[2401]), .B(n13508), .Z(n13507) );
  IV U13314 ( .A(p_input[2369]), .Z(n13508) );
  XNOR U13315 ( .A(n12693), .B(n13501), .Z(n13503) );
  XNOR U13316 ( .A(p_input[2305]), .B(n13509), .Z(n12693) );
  AND U13317 ( .A(n271), .B(n13510), .Z(n13509) );
  XOR U13318 ( .A(p_input[2337]), .B(p_input[2305]), .Z(n13510) );
  IV U13319 ( .A(n13505), .Z(n13501) );
  AND U13320 ( .A(n13231), .B(n13234), .Z(n13505) );
  XOR U13321 ( .A(p_input[2368]), .B(n13511), .Z(n13234) );
  AND U13322 ( .A(n274), .B(n13512), .Z(n13511) );
  XOR U13323 ( .A(p_input[2400]), .B(p_input[2368]), .Z(n13512) );
  XOR U13324 ( .A(n13513), .B(n13514), .Z(n274) );
  AND U13325 ( .A(n13515), .B(n13516), .Z(n13514) );
  XNOR U13326 ( .A(p_input[2431]), .B(n13513), .Z(n13516) );
  XOR U13327 ( .A(n13513), .B(p_input[2399]), .Z(n13515) );
  XOR U13328 ( .A(n13517), .B(n13518), .Z(n13513) );
  AND U13329 ( .A(n13519), .B(n13520), .Z(n13518) );
  XNOR U13330 ( .A(p_input[2430]), .B(n13517), .Z(n13520) );
  XOR U13331 ( .A(n13517), .B(p_input[2398]), .Z(n13519) );
  XOR U13332 ( .A(n13521), .B(n13522), .Z(n13517) );
  AND U13333 ( .A(n13523), .B(n13524), .Z(n13522) );
  XNOR U13334 ( .A(p_input[2429]), .B(n13521), .Z(n13524) );
  XOR U13335 ( .A(n13521), .B(p_input[2397]), .Z(n13523) );
  XOR U13336 ( .A(n13525), .B(n13526), .Z(n13521) );
  AND U13337 ( .A(n13527), .B(n13528), .Z(n13526) );
  XNOR U13338 ( .A(p_input[2428]), .B(n13525), .Z(n13528) );
  XOR U13339 ( .A(n13525), .B(p_input[2396]), .Z(n13527) );
  XOR U13340 ( .A(n13529), .B(n13530), .Z(n13525) );
  AND U13341 ( .A(n13531), .B(n13532), .Z(n13530) );
  XNOR U13342 ( .A(p_input[2427]), .B(n13529), .Z(n13532) );
  XOR U13343 ( .A(n13529), .B(p_input[2395]), .Z(n13531) );
  XOR U13344 ( .A(n13533), .B(n13534), .Z(n13529) );
  AND U13345 ( .A(n13535), .B(n13536), .Z(n13534) );
  XNOR U13346 ( .A(p_input[2426]), .B(n13533), .Z(n13536) );
  XOR U13347 ( .A(n13533), .B(p_input[2394]), .Z(n13535) );
  XOR U13348 ( .A(n13537), .B(n13538), .Z(n13533) );
  AND U13349 ( .A(n13539), .B(n13540), .Z(n13538) );
  XNOR U13350 ( .A(p_input[2425]), .B(n13537), .Z(n13540) );
  XOR U13351 ( .A(n13537), .B(p_input[2393]), .Z(n13539) );
  XOR U13352 ( .A(n13541), .B(n13542), .Z(n13537) );
  AND U13353 ( .A(n13543), .B(n13544), .Z(n13542) );
  XNOR U13354 ( .A(p_input[2424]), .B(n13541), .Z(n13544) );
  XOR U13355 ( .A(n13541), .B(p_input[2392]), .Z(n13543) );
  XOR U13356 ( .A(n13545), .B(n13546), .Z(n13541) );
  AND U13357 ( .A(n13547), .B(n13548), .Z(n13546) );
  XNOR U13358 ( .A(p_input[2423]), .B(n13545), .Z(n13548) );
  XOR U13359 ( .A(n13545), .B(p_input[2391]), .Z(n13547) );
  XOR U13360 ( .A(n13549), .B(n13550), .Z(n13545) );
  AND U13361 ( .A(n13551), .B(n13552), .Z(n13550) );
  XNOR U13362 ( .A(p_input[2422]), .B(n13549), .Z(n13552) );
  XOR U13363 ( .A(n13549), .B(p_input[2390]), .Z(n13551) );
  XOR U13364 ( .A(n13553), .B(n13554), .Z(n13549) );
  AND U13365 ( .A(n13555), .B(n13556), .Z(n13554) );
  XNOR U13366 ( .A(p_input[2421]), .B(n13553), .Z(n13556) );
  XOR U13367 ( .A(n13553), .B(p_input[2389]), .Z(n13555) );
  XOR U13368 ( .A(n13557), .B(n13558), .Z(n13553) );
  AND U13369 ( .A(n13559), .B(n13560), .Z(n13558) );
  XNOR U13370 ( .A(p_input[2420]), .B(n13557), .Z(n13560) );
  XOR U13371 ( .A(n13557), .B(p_input[2388]), .Z(n13559) );
  XOR U13372 ( .A(n13561), .B(n13562), .Z(n13557) );
  AND U13373 ( .A(n13563), .B(n13564), .Z(n13562) );
  XNOR U13374 ( .A(p_input[2419]), .B(n13561), .Z(n13564) );
  XOR U13375 ( .A(n13561), .B(p_input[2387]), .Z(n13563) );
  XOR U13376 ( .A(n13565), .B(n13566), .Z(n13561) );
  AND U13377 ( .A(n13567), .B(n13568), .Z(n13566) );
  XNOR U13378 ( .A(p_input[2418]), .B(n13565), .Z(n13568) );
  XOR U13379 ( .A(n13565), .B(p_input[2386]), .Z(n13567) );
  XOR U13380 ( .A(n13569), .B(n13570), .Z(n13565) );
  AND U13381 ( .A(n13571), .B(n13572), .Z(n13570) );
  XNOR U13382 ( .A(p_input[2417]), .B(n13569), .Z(n13572) );
  XOR U13383 ( .A(n13569), .B(p_input[2385]), .Z(n13571) );
  XOR U13384 ( .A(n13573), .B(n13574), .Z(n13569) );
  AND U13385 ( .A(n13575), .B(n13576), .Z(n13574) );
  XNOR U13386 ( .A(p_input[2416]), .B(n13573), .Z(n13576) );
  XOR U13387 ( .A(n13573), .B(p_input[2384]), .Z(n13575) );
  XOR U13388 ( .A(n13577), .B(n13578), .Z(n13573) );
  AND U13389 ( .A(n13579), .B(n13580), .Z(n13578) );
  XNOR U13390 ( .A(p_input[2415]), .B(n13577), .Z(n13580) );
  XOR U13391 ( .A(n13577), .B(p_input[2383]), .Z(n13579) );
  XOR U13392 ( .A(n13581), .B(n13582), .Z(n13577) );
  AND U13393 ( .A(n13583), .B(n13584), .Z(n13582) );
  XNOR U13394 ( .A(p_input[2414]), .B(n13581), .Z(n13584) );
  XOR U13395 ( .A(n13581), .B(p_input[2382]), .Z(n13583) );
  XOR U13396 ( .A(n13585), .B(n13586), .Z(n13581) );
  AND U13397 ( .A(n13587), .B(n13588), .Z(n13586) );
  XNOR U13398 ( .A(p_input[2413]), .B(n13585), .Z(n13588) );
  XOR U13399 ( .A(n13585), .B(p_input[2381]), .Z(n13587) );
  XOR U13400 ( .A(n13589), .B(n13590), .Z(n13585) );
  AND U13401 ( .A(n13591), .B(n13592), .Z(n13590) );
  XNOR U13402 ( .A(p_input[2412]), .B(n13589), .Z(n13592) );
  XOR U13403 ( .A(n13589), .B(p_input[2380]), .Z(n13591) );
  XOR U13404 ( .A(n13593), .B(n13594), .Z(n13589) );
  AND U13405 ( .A(n13595), .B(n13596), .Z(n13594) );
  XNOR U13406 ( .A(p_input[2411]), .B(n13593), .Z(n13596) );
  XOR U13407 ( .A(n13593), .B(p_input[2379]), .Z(n13595) );
  XOR U13408 ( .A(n13597), .B(n13598), .Z(n13593) );
  AND U13409 ( .A(n13599), .B(n13600), .Z(n13598) );
  XNOR U13410 ( .A(p_input[2410]), .B(n13597), .Z(n13600) );
  XOR U13411 ( .A(n13597), .B(p_input[2378]), .Z(n13599) );
  XOR U13412 ( .A(n13601), .B(n13602), .Z(n13597) );
  AND U13413 ( .A(n13603), .B(n13604), .Z(n13602) );
  XNOR U13414 ( .A(p_input[2409]), .B(n13601), .Z(n13604) );
  XOR U13415 ( .A(n13601), .B(p_input[2377]), .Z(n13603) );
  XOR U13416 ( .A(n13605), .B(n13606), .Z(n13601) );
  AND U13417 ( .A(n13607), .B(n13608), .Z(n13606) );
  XNOR U13418 ( .A(p_input[2408]), .B(n13605), .Z(n13608) );
  XOR U13419 ( .A(n13605), .B(p_input[2376]), .Z(n13607) );
  XOR U13420 ( .A(n13609), .B(n13610), .Z(n13605) );
  AND U13421 ( .A(n13611), .B(n13612), .Z(n13610) );
  XNOR U13422 ( .A(p_input[2407]), .B(n13609), .Z(n13612) );
  XOR U13423 ( .A(n13609), .B(p_input[2375]), .Z(n13611) );
  XOR U13424 ( .A(n13613), .B(n13614), .Z(n13609) );
  AND U13425 ( .A(n13615), .B(n13616), .Z(n13614) );
  XNOR U13426 ( .A(p_input[2406]), .B(n13613), .Z(n13616) );
  XOR U13427 ( .A(n13613), .B(p_input[2374]), .Z(n13615) );
  XOR U13428 ( .A(n13617), .B(n13618), .Z(n13613) );
  AND U13429 ( .A(n13619), .B(n13620), .Z(n13618) );
  XNOR U13430 ( .A(p_input[2405]), .B(n13617), .Z(n13620) );
  XOR U13431 ( .A(n13617), .B(p_input[2373]), .Z(n13619) );
  XOR U13432 ( .A(n13621), .B(n13622), .Z(n13617) );
  AND U13433 ( .A(n13623), .B(n13624), .Z(n13622) );
  XNOR U13434 ( .A(p_input[2404]), .B(n13621), .Z(n13624) );
  XOR U13435 ( .A(n13621), .B(p_input[2372]), .Z(n13623) );
  XOR U13436 ( .A(n13625), .B(n13626), .Z(n13621) );
  AND U13437 ( .A(n13627), .B(n13628), .Z(n13626) );
  XNOR U13438 ( .A(p_input[2403]), .B(n13625), .Z(n13628) );
  XOR U13439 ( .A(n13625), .B(p_input[2371]), .Z(n13627) );
  XOR U13440 ( .A(n13629), .B(n13630), .Z(n13625) );
  AND U13441 ( .A(n13631), .B(n13632), .Z(n13630) );
  XNOR U13442 ( .A(p_input[2402]), .B(n13629), .Z(n13632) );
  XOR U13443 ( .A(n13629), .B(p_input[2370]), .Z(n13631) );
  XNOR U13444 ( .A(n13633), .B(n13634), .Z(n13629) );
  AND U13445 ( .A(n13635), .B(n13636), .Z(n13634) );
  XOR U13446 ( .A(p_input[2401]), .B(n13633), .Z(n13636) );
  XNOR U13447 ( .A(p_input[2369]), .B(n13633), .Z(n13635) );
  AND U13448 ( .A(p_input[2400]), .B(n13637), .Z(n13633) );
  IV U13449 ( .A(p_input[2368]), .Z(n13637) );
  XNOR U13450 ( .A(p_input[2304]), .B(n13638), .Z(n13231) );
  AND U13451 ( .A(n271), .B(n13639), .Z(n13638) );
  XOR U13452 ( .A(p_input[2336]), .B(p_input[2304]), .Z(n13639) );
  XOR U13453 ( .A(n13640), .B(n13641), .Z(n271) );
  AND U13454 ( .A(n13642), .B(n13643), .Z(n13641) );
  XNOR U13455 ( .A(p_input[2367]), .B(n13640), .Z(n13643) );
  XOR U13456 ( .A(n13640), .B(p_input[2335]), .Z(n13642) );
  XOR U13457 ( .A(n13644), .B(n13645), .Z(n13640) );
  AND U13458 ( .A(n13646), .B(n13647), .Z(n13645) );
  XNOR U13459 ( .A(p_input[2366]), .B(n13644), .Z(n13647) );
  XNOR U13460 ( .A(n13644), .B(n13246), .Z(n13646) );
  IV U13461 ( .A(p_input[2334]), .Z(n13246) );
  XOR U13462 ( .A(n13648), .B(n13649), .Z(n13644) );
  AND U13463 ( .A(n13650), .B(n13651), .Z(n13649) );
  XNOR U13464 ( .A(p_input[2365]), .B(n13648), .Z(n13651) );
  XNOR U13465 ( .A(n13648), .B(n13255), .Z(n13650) );
  IV U13466 ( .A(p_input[2333]), .Z(n13255) );
  XOR U13467 ( .A(n13652), .B(n13653), .Z(n13648) );
  AND U13468 ( .A(n13654), .B(n13655), .Z(n13653) );
  XNOR U13469 ( .A(p_input[2364]), .B(n13652), .Z(n13655) );
  XNOR U13470 ( .A(n13652), .B(n13264), .Z(n13654) );
  IV U13471 ( .A(p_input[2332]), .Z(n13264) );
  XOR U13472 ( .A(n13656), .B(n13657), .Z(n13652) );
  AND U13473 ( .A(n13658), .B(n13659), .Z(n13657) );
  XNOR U13474 ( .A(p_input[2363]), .B(n13656), .Z(n13659) );
  XNOR U13475 ( .A(n13656), .B(n13273), .Z(n13658) );
  IV U13476 ( .A(p_input[2331]), .Z(n13273) );
  XOR U13477 ( .A(n13660), .B(n13661), .Z(n13656) );
  AND U13478 ( .A(n13662), .B(n13663), .Z(n13661) );
  XNOR U13479 ( .A(p_input[2362]), .B(n13660), .Z(n13663) );
  XNOR U13480 ( .A(n13660), .B(n13282), .Z(n13662) );
  IV U13481 ( .A(p_input[2330]), .Z(n13282) );
  XOR U13482 ( .A(n13664), .B(n13665), .Z(n13660) );
  AND U13483 ( .A(n13666), .B(n13667), .Z(n13665) );
  XNOR U13484 ( .A(p_input[2361]), .B(n13664), .Z(n13667) );
  XNOR U13485 ( .A(n13664), .B(n13291), .Z(n13666) );
  IV U13486 ( .A(p_input[2329]), .Z(n13291) );
  XOR U13487 ( .A(n13668), .B(n13669), .Z(n13664) );
  AND U13488 ( .A(n13670), .B(n13671), .Z(n13669) );
  XNOR U13489 ( .A(p_input[2360]), .B(n13668), .Z(n13671) );
  XNOR U13490 ( .A(n13668), .B(n13300), .Z(n13670) );
  IV U13491 ( .A(p_input[2328]), .Z(n13300) );
  XOR U13492 ( .A(n13672), .B(n13673), .Z(n13668) );
  AND U13493 ( .A(n13674), .B(n13675), .Z(n13673) );
  XNOR U13494 ( .A(p_input[2359]), .B(n13672), .Z(n13675) );
  XNOR U13495 ( .A(n13672), .B(n13309), .Z(n13674) );
  IV U13496 ( .A(p_input[2327]), .Z(n13309) );
  XOR U13497 ( .A(n13676), .B(n13677), .Z(n13672) );
  AND U13498 ( .A(n13678), .B(n13679), .Z(n13677) );
  XNOR U13499 ( .A(p_input[2358]), .B(n13676), .Z(n13679) );
  XNOR U13500 ( .A(n13676), .B(n13318), .Z(n13678) );
  IV U13501 ( .A(p_input[2326]), .Z(n13318) );
  XOR U13502 ( .A(n13680), .B(n13681), .Z(n13676) );
  AND U13503 ( .A(n13682), .B(n13683), .Z(n13681) );
  XNOR U13504 ( .A(p_input[2357]), .B(n13680), .Z(n13683) );
  XNOR U13505 ( .A(n13680), .B(n13327), .Z(n13682) );
  IV U13506 ( .A(p_input[2325]), .Z(n13327) );
  XOR U13507 ( .A(n13684), .B(n13685), .Z(n13680) );
  AND U13508 ( .A(n13686), .B(n13687), .Z(n13685) );
  XNOR U13509 ( .A(p_input[2356]), .B(n13684), .Z(n13687) );
  XNOR U13510 ( .A(n13684), .B(n13336), .Z(n13686) );
  IV U13511 ( .A(p_input[2324]), .Z(n13336) );
  XOR U13512 ( .A(n13688), .B(n13689), .Z(n13684) );
  AND U13513 ( .A(n13690), .B(n13691), .Z(n13689) );
  XNOR U13514 ( .A(p_input[2355]), .B(n13688), .Z(n13691) );
  XNOR U13515 ( .A(n13688), .B(n13345), .Z(n13690) );
  IV U13516 ( .A(p_input[2323]), .Z(n13345) );
  XOR U13517 ( .A(n13692), .B(n13693), .Z(n13688) );
  AND U13518 ( .A(n13694), .B(n13695), .Z(n13693) );
  XNOR U13519 ( .A(p_input[2354]), .B(n13692), .Z(n13695) );
  XNOR U13520 ( .A(n13692), .B(n13354), .Z(n13694) );
  IV U13521 ( .A(p_input[2322]), .Z(n13354) );
  XOR U13522 ( .A(n13696), .B(n13697), .Z(n13692) );
  AND U13523 ( .A(n13698), .B(n13699), .Z(n13697) );
  XNOR U13524 ( .A(p_input[2353]), .B(n13696), .Z(n13699) );
  XNOR U13525 ( .A(n13696), .B(n13363), .Z(n13698) );
  IV U13526 ( .A(p_input[2321]), .Z(n13363) );
  XOR U13527 ( .A(n13700), .B(n13701), .Z(n13696) );
  AND U13528 ( .A(n13702), .B(n13703), .Z(n13701) );
  XNOR U13529 ( .A(p_input[2352]), .B(n13700), .Z(n13703) );
  XNOR U13530 ( .A(n13700), .B(n13372), .Z(n13702) );
  IV U13531 ( .A(p_input[2320]), .Z(n13372) );
  XOR U13532 ( .A(n13704), .B(n13705), .Z(n13700) );
  AND U13533 ( .A(n13706), .B(n13707), .Z(n13705) );
  XNOR U13534 ( .A(p_input[2351]), .B(n13704), .Z(n13707) );
  XNOR U13535 ( .A(n13704), .B(n13381), .Z(n13706) );
  IV U13536 ( .A(p_input[2319]), .Z(n13381) );
  XOR U13537 ( .A(n13708), .B(n13709), .Z(n13704) );
  AND U13538 ( .A(n13710), .B(n13711), .Z(n13709) );
  XNOR U13539 ( .A(p_input[2350]), .B(n13708), .Z(n13711) );
  XNOR U13540 ( .A(n13708), .B(n13390), .Z(n13710) );
  IV U13541 ( .A(p_input[2318]), .Z(n13390) );
  XOR U13542 ( .A(n13712), .B(n13713), .Z(n13708) );
  AND U13543 ( .A(n13714), .B(n13715), .Z(n13713) );
  XNOR U13544 ( .A(p_input[2349]), .B(n13712), .Z(n13715) );
  XNOR U13545 ( .A(n13712), .B(n13399), .Z(n13714) );
  IV U13546 ( .A(p_input[2317]), .Z(n13399) );
  XOR U13547 ( .A(n13716), .B(n13717), .Z(n13712) );
  AND U13548 ( .A(n13718), .B(n13719), .Z(n13717) );
  XNOR U13549 ( .A(p_input[2348]), .B(n13716), .Z(n13719) );
  XNOR U13550 ( .A(n13716), .B(n13408), .Z(n13718) );
  IV U13551 ( .A(p_input[2316]), .Z(n13408) );
  XOR U13552 ( .A(n13720), .B(n13721), .Z(n13716) );
  AND U13553 ( .A(n13722), .B(n13723), .Z(n13721) );
  XNOR U13554 ( .A(p_input[2347]), .B(n13720), .Z(n13723) );
  XNOR U13555 ( .A(n13720), .B(n13417), .Z(n13722) );
  IV U13556 ( .A(p_input[2315]), .Z(n13417) );
  XOR U13557 ( .A(n13724), .B(n13725), .Z(n13720) );
  AND U13558 ( .A(n13726), .B(n13727), .Z(n13725) );
  XNOR U13559 ( .A(p_input[2346]), .B(n13724), .Z(n13727) );
  XNOR U13560 ( .A(n13724), .B(n13426), .Z(n13726) );
  IV U13561 ( .A(p_input[2314]), .Z(n13426) );
  XOR U13562 ( .A(n13728), .B(n13729), .Z(n13724) );
  AND U13563 ( .A(n13730), .B(n13731), .Z(n13729) );
  XNOR U13564 ( .A(p_input[2345]), .B(n13728), .Z(n13731) );
  XNOR U13565 ( .A(n13728), .B(n13435), .Z(n13730) );
  IV U13566 ( .A(p_input[2313]), .Z(n13435) );
  XOR U13567 ( .A(n13732), .B(n13733), .Z(n13728) );
  AND U13568 ( .A(n13734), .B(n13735), .Z(n13733) );
  XNOR U13569 ( .A(p_input[2344]), .B(n13732), .Z(n13735) );
  XNOR U13570 ( .A(n13732), .B(n13444), .Z(n13734) );
  IV U13571 ( .A(p_input[2312]), .Z(n13444) );
  XOR U13572 ( .A(n13736), .B(n13737), .Z(n13732) );
  AND U13573 ( .A(n13738), .B(n13739), .Z(n13737) );
  XNOR U13574 ( .A(p_input[2343]), .B(n13736), .Z(n13739) );
  XNOR U13575 ( .A(n13736), .B(n13453), .Z(n13738) );
  IV U13576 ( .A(p_input[2311]), .Z(n13453) );
  XOR U13577 ( .A(n13740), .B(n13741), .Z(n13736) );
  AND U13578 ( .A(n13742), .B(n13743), .Z(n13741) );
  XNOR U13579 ( .A(p_input[2342]), .B(n13740), .Z(n13743) );
  XNOR U13580 ( .A(n13740), .B(n13462), .Z(n13742) );
  IV U13581 ( .A(p_input[2310]), .Z(n13462) );
  XOR U13582 ( .A(n13744), .B(n13745), .Z(n13740) );
  AND U13583 ( .A(n13746), .B(n13747), .Z(n13745) );
  XNOR U13584 ( .A(p_input[2341]), .B(n13744), .Z(n13747) );
  XNOR U13585 ( .A(n13744), .B(n13471), .Z(n13746) );
  IV U13586 ( .A(p_input[2309]), .Z(n13471) );
  XOR U13587 ( .A(n13748), .B(n13749), .Z(n13744) );
  AND U13588 ( .A(n13750), .B(n13751), .Z(n13749) );
  XNOR U13589 ( .A(p_input[2340]), .B(n13748), .Z(n13751) );
  XNOR U13590 ( .A(n13748), .B(n13480), .Z(n13750) );
  IV U13591 ( .A(p_input[2308]), .Z(n13480) );
  XOR U13592 ( .A(n13752), .B(n13753), .Z(n13748) );
  AND U13593 ( .A(n13754), .B(n13755), .Z(n13753) );
  XNOR U13594 ( .A(p_input[2339]), .B(n13752), .Z(n13755) );
  XNOR U13595 ( .A(n13752), .B(n13489), .Z(n13754) );
  IV U13596 ( .A(p_input[2307]), .Z(n13489) );
  XOR U13597 ( .A(n13756), .B(n13757), .Z(n13752) );
  AND U13598 ( .A(n13758), .B(n13759), .Z(n13757) );
  XNOR U13599 ( .A(p_input[2338]), .B(n13756), .Z(n13759) );
  XNOR U13600 ( .A(n13756), .B(n13498), .Z(n13758) );
  IV U13601 ( .A(p_input[2306]), .Z(n13498) );
  XNOR U13602 ( .A(n13760), .B(n13761), .Z(n13756) );
  AND U13603 ( .A(n13762), .B(n13763), .Z(n13761) );
  XOR U13604 ( .A(p_input[2337]), .B(n13760), .Z(n13763) );
  XNOR U13605 ( .A(p_input[2305]), .B(n13760), .Z(n13762) );
  AND U13606 ( .A(p_input[2336]), .B(n13764), .Z(n13760) );
  IV U13607 ( .A(p_input[2304]), .Z(n13764) );
  XOR U13608 ( .A(n13765), .B(n13766), .Z(n11943) );
  AND U13609 ( .A(n503), .B(n13767), .Z(n13766) );
  XNOR U13610 ( .A(n13768), .B(n13765), .Z(n13767) );
  XOR U13611 ( .A(n13769), .B(n13770), .Z(n503) );
  AND U13612 ( .A(n13771), .B(n13772), .Z(n13770) );
  XOR U13613 ( .A(n13769), .B(n11958), .Z(n13772) );
  XNOR U13614 ( .A(n13773), .B(n13774), .Z(n11958) );
  AND U13615 ( .A(n13775), .B(n350), .Z(n13774) );
  AND U13616 ( .A(n13773), .B(n13776), .Z(n13775) );
  XNOR U13617 ( .A(n11955), .B(n13769), .Z(n13771) );
  XOR U13618 ( .A(n13777), .B(n13778), .Z(n11955) );
  AND U13619 ( .A(n13779), .B(n347), .Z(n13778) );
  NOR U13620 ( .A(n13777), .B(n13780), .Z(n13779) );
  XOR U13621 ( .A(n13781), .B(n13782), .Z(n13769) );
  AND U13622 ( .A(n13783), .B(n13784), .Z(n13782) );
  XOR U13623 ( .A(n13781), .B(n11970), .Z(n13784) );
  XOR U13624 ( .A(n13785), .B(n13786), .Z(n11970) );
  AND U13625 ( .A(n350), .B(n13787), .Z(n13786) );
  XOR U13626 ( .A(n13788), .B(n13785), .Z(n13787) );
  XNOR U13627 ( .A(n11967), .B(n13781), .Z(n13783) );
  XOR U13628 ( .A(n13789), .B(n13790), .Z(n11967) );
  AND U13629 ( .A(n347), .B(n13791), .Z(n13790) );
  XOR U13630 ( .A(n13792), .B(n13789), .Z(n13791) );
  XOR U13631 ( .A(n13793), .B(n13794), .Z(n13781) );
  AND U13632 ( .A(n13795), .B(n13796), .Z(n13794) );
  XOR U13633 ( .A(n13793), .B(n11982), .Z(n13796) );
  XOR U13634 ( .A(n13797), .B(n13798), .Z(n11982) );
  AND U13635 ( .A(n350), .B(n13799), .Z(n13798) );
  XOR U13636 ( .A(n13800), .B(n13797), .Z(n13799) );
  XNOR U13637 ( .A(n11979), .B(n13793), .Z(n13795) );
  XOR U13638 ( .A(n13801), .B(n13802), .Z(n11979) );
  AND U13639 ( .A(n347), .B(n13803), .Z(n13802) );
  XOR U13640 ( .A(n13804), .B(n13801), .Z(n13803) );
  XOR U13641 ( .A(n13805), .B(n13806), .Z(n13793) );
  AND U13642 ( .A(n13807), .B(n13808), .Z(n13806) );
  XOR U13643 ( .A(n13805), .B(n11994), .Z(n13808) );
  XOR U13644 ( .A(n13809), .B(n13810), .Z(n11994) );
  AND U13645 ( .A(n350), .B(n13811), .Z(n13810) );
  XOR U13646 ( .A(n13812), .B(n13809), .Z(n13811) );
  XNOR U13647 ( .A(n11991), .B(n13805), .Z(n13807) );
  XOR U13648 ( .A(n13813), .B(n13814), .Z(n11991) );
  AND U13649 ( .A(n347), .B(n13815), .Z(n13814) );
  XOR U13650 ( .A(n13816), .B(n13813), .Z(n13815) );
  XOR U13651 ( .A(n13817), .B(n13818), .Z(n13805) );
  AND U13652 ( .A(n13819), .B(n13820), .Z(n13818) );
  XOR U13653 ( .A(n13817), .B(n12006), .Z(n13820) );
  XOR U13654 ( .A(n13821), .B(n13822), .Z(n12006) );
  AND U13655 ( .A(n350), .B(n13823), .Z(n13822) );
  XOR U13656 ( .A(n13824), .B(n13821), .Z(n13823) );
  XNOR U13657 ( .A(n12003), .B(n13817), .Z(n13819) );
  XOR U13658 ( .A(n13825), .B(n13826), .Z(n12003) );
  AND U13659 ( .A(n347), .B(n13827), .Z(n13826) );
  XOR U13660 ( .A(n13828), .B(n13825), .Z(n13827) );
  XOR U13661 ( .A(n13829), .B(n13830), .Z(n13817) );
  AND U13662 ( .A(n13831), .B(n13832), .Z(n13830) );
  XOR U13663 ( .A(n13829), .B(n12018), .Z(n13832) );
  XOR U13664 ( .A(n13833), .B(n13834), .Z(n12018) );
  AND U13665 ( .A(n350), .B(n13835), .Z(n13834) );
  XOR U13666 ( .A(n13836), .B(n13833), .Z(n13835) );
  XNOR U13667 ( .A(n12015), .B(n13829), .Z(n13831) );
  XOR U13668 ( .A(n13837), .B(n13838), .Z(n12015) );
  AND U13669 ( .A(n347), .B(n13839), .Z(n13838) );
  XOR U13670 ( .A(n13840), .B(n13837), .Z(n13839) );
  XOR U13671 ( .A(n13841), .B(n13842), .Z(n13829) );
  AND U13672 ( .A(n13843), .B(n13844), .Z(n13842) );
  XOR U13673 ( .A(n13841), .B(n12030), .Z(n13844) );
  XOR U13674 ( .A(n13845), .B(n13846), .Z(n12030) );
  AND U13675 ( .A(n350), .B(n13847), .Z(n13846) );
  XOR U13676 ( .A(n13848), .B(n13845), .Z(n13847) );
  XNOR U13677 ( .A(n12027), .B(n13841), .Z(n13843) );
  XOR U13678 ( .A(n13849), .B(n13850), .Z(n12027) );
  AND U13679 ( .A(n347), .B(n13851), .Z(n13850) );
  XOR U13680 ( .A(n13852), .B(n13849), .Z(n13851) );
  XOR U13681 ( .A(n13853), .B(n13854), .Z(n13841) );
  AND U13682 ( .A(n13855), .B(n13856), .Z(n13854) );
  XOR U13683 ( .A(n13853), .B(n12042), .Z(n13856) );
  XOR U13684 ( .A(n13857), .B(n13858), .Z(n12042) );
  AND U13685 ( .A(n350), .B(n13859), .Z(n13858) );
  XOR U13686 ( .A(n13860), .B(n13857), .Z(n13859) );
  XNOR U13687 ( .A(n12039), .B(n13853), .Z(n13855) );
  XOR U13688 ( .A(n13861), .B(n13862), .Z(n12039) );
  AND U13689 ( .A(n347), .B(n13863), .Z(n13862) );
  XOR U13690 ( .A(n13864), .B(n13861), .Z(n13863) );
  XOR U13691 ( .A(n13865), .B(n13866), .Z(n13853) );
  AND U13692 ( .A(n13867), .B(n13868), .Z(n13866) );
  XOR U13693 ( .A(n13865), .B(n12054), .Z(n13868) );
  XOR U13694 ( .A(n13869), .B(n13870), .Z(n12054) );
  AND U13695 ( .A(n350), .B(n13871), .Z(n13870) );
  XOR U13696 ( .A(n13872), .B(n13869), .Z(n13871) );
  XNOR U13697 ( .A(n12051), .B(n13865), .Z(n13867) );
  XOR U13698 ( .A(n13873), .B(n13874), .Z(n12051) );
  AND U13699 ( .A(n347), .B(n13875), .Z(n13874) );
  XOR U13700 ( .A(n13876), .B(n13873), .Z(n13875) );
  XOR U13701 ( .A(n13877), .B(n13878), .Z(n13865) );
  AND U13702 ( .A(n13879), .B(n13880), .Z(n13878) );
  XOR U13703 ( .A(n13877), .B(n12066), .Z(n13880) );
  XOR U13704 ( .A(n13881), .B(n13882), .Z(n12066) );
  AND U13705 ( .A(n350), .B(n13883), .Z(n13882) );
  XOR U13706 ( .A(n13884), .B(n13881), .Z(n13883) );
  XNOR U13707 ( .A(n12063), .B(n13877), .Z(n13879) );
  XOR U13708 ( .A(n13885), .B(n13886), .Z(n12063) );
  AND U13709 ( .A(n347), .B(n13887), .Z(n13886) );
  XOR U13710 ( .A(n13888), .B(n13885), .Z(n13887) );
  XOR U13711 ( .A(n13889), .B(n13890), .Z(n13877) );
  AND U13712 ( .A(n13891), .B(n13892), .Z(n13890) );
  XOR U13713 ( .A(n13889), .B(n12078), .Z(n13892) );
  XOR U13714 ( .A(n13893), .B(n13894), .Z(n12078) );
  AND U13715 ( .A(n350), .B(n13895), .Z(n13894) );
  XOR U13716 ( .A(n13896), .B(n13893), .Z(n13895) );
  XNOR U13717 ( .A(n12075), .B(n13889), .Z(n13891) );
  XOR U13718 ( .A(n13897), .B(n13898), .Z(n12075) );
  AND U13719 ( .A(n347), .B(n13899), .Z(n13898) );
  XOR U13720 ( .A(n13900), .B(n13897), .Z(n13899) );
  XOR U13721 ( .A(n13901), .B(n13902), .Z(n13889) );
  AND U13722 ( .A(n13903), .B(n13904), .Z(n13902) );
  XOR U13723 ( .A(n13901), .B(n12090), .Z(n13904) );
  XOR U13724 ( .A(n13905), .B(n13906), .Z(n12090) );
  AND U13725 ( .A(n350), .B(n13907), .Z(n13906) );
  XOR U13726 ( .A(n13908), .B(n13905), .Z(n13907) );
  XNOR U13727 ( .A(n12087), .B(n13901), .Z(n13903) );
  XOR U13728 ( .A(n13909), .B(n13910), .Z(n12087) );
  AND U13729 ( .A(n347), .B(n13911), .Z(n13910) );
  XOR U13730 ( .A(n13912), .B(n13909), .Z(n13911) );
  XOR U13731 ( .A(n13913), .B(n13914), .Z(n13901) );
  AND U13732 ( .A(n13915), .B(n13916), .Z(n13914) );
  XOR U13733 ( .A(n13913), .B(n12102), .Z(n13916) );
  XOR U13734 ( .A(n13917), .B(n13918), .Z(n12102) );
  AND U13735 ( .A(n350), .B(n13919), .Z(n13918) );
  XOR U13736 ( .A(n13920), .B(n13917), .Z(n13919) );
  XNOR U13737 ( .A(n12099), .B(n13913), .Z(n13915) );
  XOR U13738 ( .A(n13921), .B(n13922), .Z(n12099) );
  AND U13739 ( .A(n347), .B(n13923), .Z(n13922) );
  XOR U13740 ( .A(n13924), .B(n13921), .Z(n13923) );
  XOR U13741 ( .A(n13925), .B(n13926), .Z(n13913) );
  AND U13742 ( .A(n13927), .B(n13928), .Z(n13926) );
  XOR U13743 ( .A(n13925), .B(n12114), .Z(n13928) );
  XOR U13744 ( .A(n13929), .B(n13930), .Z(n12114) );
  AND U13745 ( .A(n350), .B(n13931), .Z(n13930) );
  XOR U13746 ( .A(n13932), .B(n13929), .Z(n13931) );
  XNOR U13747 ( .A(n12111), .B(n13925), .Z(n13927) );
  XOR U13748 ( .A(n13933), .B(n13934), .Z(n12111) );
  AND U13749 ( .A(n347), .B(n13935), .Z(n13934) );
  XOR U13750 ( .A(n13936), .B(n13933), .Z(n13935) );
  XOR U13751 ( .A(n13937), .B(n13938), .Z(n13925) );
  AND U13752 ( .A(n13939), .B(n13940), .Z(n13938) );
  XOR U13753 ( .A(n13937), .B(n12126), .Z(n13940) );
  XOR U13754 ( .A(n13941), .B(n13942), .Z(n12126) );
  AND U13755 ( .A(n350), .B(n13943), .Z(n13942) );
  XOR U13756 ( .A(n13944), .B(n13941), .Z(n13943) );
  XNOR U13757 ( .A(n12123), .B(n13937), .Z(n13939) );
  XOR U13758 ( .A(n13945), .B(n13946), .Z(n12123) );
  AND U13759 ( .A(n347), .B(n13947), .Z(n13946) );
  XOR U13760 ( .A(n13948), .B(n13945), .Z(n13947) );
  XOR U13761 ( .A(n13949), .B(n13950), .Z(n13937) );
  AND U13762 ( .A(n13951), .B(n13952), .Z(n13950) );
  XOR U13763 ( .A(n13949), .B(n12138), .Z(n13952) );
  XOR U13764 ( .A(n13953), .B(n13954), .Z(n12138) );
  AND U13765 ( .A(n350), .B(n13955), .Z(n13954) );
  XOR U13766 ( .A(n13956), .B(n13953), .Z(n13955) );
  XNOR U13767 ( .A(n12135), .B(n13949), .Z(n13951) );
  XOR U13768 ( .A(n13957), .B(n13958), .Z(n12135) );
  AND U13769 ( .A(n347), .B(n13959), .Z(n13958) );
  XOR U13770 ( .A(n13960), .B(n13957), .Z(n13959) );
  XOR U13771 ( .A(n13961), .B(n13962), .Z(n13949) );
  AND U13772 ( .A(n13963), .B(n13964), .Z(n13962) );
  XOR U13773 ( .A(n13961), .B(n12150), .Z(n13964) );
  XOR U13774 ( .A(n13965), .B(n13966), .Z(n12150) );
  AND U13775 ( .A(n350), .B(n13967), .Z(n13966) );
  XOR U13776 ( .A(n13968), .B(n13965), .Z(n13967) );
  XNOR U13777 ( .A(n12147), .B(n13961), .Z(n13963) );
  XOR U13778 ( .A(n13969), .B(n13970), .Z(n12147) );
  AND U13779 ( .A(n347), .B(n13971), .Z(n13970) );
  XOR U13780 ( .A(n13972), .B(n13969), .Z(n13971) );
  XOR U13781 ( .A(n13973), .B(n13974), .Z(n13961) );
  AND U13782 ( .A(n13975), .B(n13976), .Z(n13974) );
  XOR U13783 ( .A(n13973), .B(n12162), .Z(n13976) );
  XOR U13784 ( .A(n13977), .B(n13978), .Z(n12162) );
  AND U13785 ( .A(n350), .B(n13979), .Z(n13978) );
  XOR U13786 ( .A(n13980), .B(n13977), .Z(n13979) );
  XNOR U13787 ( .A(n12159), .B(n13973), .Z(n13975) );
  XOR U13788 ( .A(n13981), .B(n13982), .Z(n12159) );
  AND U13789 ( .A(n347), .B(n13983), .Z(n13982) );
  XOR U13790 ( .A(n13984), .B(n13981), .Z(n13983) );
  XOR U13791 ( .A(n13985), .B(n13986), .Z(n13973) );
  AND U13792 ( .A(n13987), .B(n13988), .Z(n13986) );
  XOR U13793 ( .A(n13985), .B(n12174), .Z(n13988) );
  XOR U13794 ( .A(n13989), .B(n13990), .Z(n12174) );
  AND U13795 ( .A(n350), .B(n13991), .Z(n13990) );
  XOR U13796 ( .A(n13992), .B(n13989), .Z(n13991) );
  XNOR U13797 ( .A(n12171), .B(n13985), .Z(n13987) );
  XOR U13798 ( .A(n13993), .B(n13994), .Z(n12171) );
  AND U13799 ( .A(n347), .B(n13995), .Z(n13994) );
  XOR U13800 ( .A(n13996), .B(n13993), .Z(n13995) );
  XOR U13801 ( .A(n13997), .B(n13998), .Z(n13985) );
  AND U13802 ( .A(n13999), .B(n14000), .Z(n13998) );
  XOR U13803 ( .A(n13997), .B(n12186), .Z(n14000) );
  XOR U13804 ( .A(n14001), .B(n14002), .Z(n12186) );
  AND U13805 ( .A(n350), .B(n14003), .Z(n14002) );
  XOR U13806 ( .A(n14004), .B(n14001), .Z(n14003) );
  XNOR U13807 ( .A(n12183), .B(n13997), .Z(n13999) );
  XOR U13808 ( .A(n14005), .B(n14006), .Z(n12183) );
  AND U13809 ( .A(n347), .B(n14007), .Z(n14006) );
  XOR U13810 ( .A(n14008), .B(n14005), .Z(n14007) );
  XOR U13811 ( .A(n14009), .B(n14010), .Z(n13997) );
  AND U13812 ( .A(n14011), .B(n14012), .Z(n14010) );
  XOR U13813 ( .A(n14009), .B(n12198), .Z(n14012) );
  XOR U13814 ( .A(n14013), .B(n14014), .Z(n12198) );
  AND U13815 ( .A(n350), .B(n14015), .Z(n14014) );
  XOR U13816 ( .A(n14016), .B(n14013), .Z(n14015) );
  XNOR U13817 ( .A(n12195), .B(n14009), .Z(n14011) );
  XOR U13818 ( .A(n14017), .B(n14018), .Z(n12195) );
  AND U13819 ( .A(n347), .B(n14019), .Z(n14018) );
  XOR U13820 ( .A(n14020), .B(n14017), .Z(n14019) );
  XOR U13821 ( .A(n14021), .B(n14022), .Z(n14009) );
  AND U13822 ( .A(n14023), .B(n14024), .Z(n14022) );
  XOR U13823 ( .A(n14021), .B(n12210), .Z(n14024) );
  XOR U13824 ( .A(n14025), .B(n14026), .Z(n12210) );
  AND U13825 ( .A(n350), .B(n14027), .Z(n14026) );
  XOR U13826 ( .A(n14028), .B(n14025), .Z(n14027) );
  XNOR U13827 ( .A(n12207), .B(n14021), .Z(n14023) );
  XOR U13828 ( .A(n14029), .B(n14030), .Z(n12207) );
  AND U13829 ( .A(n347), .B(n14031), .Z(n14030) );
  XOR U13830 ( .A(n14032), .B(n14029), .Z(n14031) );
  XOR U13831 ( .A(n14033), .B(n14034), .Z(n14021) );
  AND U13832 ( .A(n14035), .B(n14036), .Z(n14034) );
  XOR U13833 ( .A(n14033), .B(n12222), .Z(n14036) );
  XOR U13834 ( .A(n14037), .B(n14038), .Z(n12222) );
  AND U13835 ( .A(n350), .B(n14039), .Z(n14038) );
  XOR U13836 ( .A(n14040), .B(n14037), .Z(n14039) );
  XNOR U13837 ( .A(n12219), .B(n14033), .Z(n14035) );
  XOR U13838 ( .A(n14041), .B(n14042), .Z(n12219) );
  AND U13839 ( .A(n347), .B(n14043), .Z(n14042) );
  XOR U13840 ( .A(n14044), .B(n14041), .Z(n14043) );
  XOR U13841 ( .A(n14045), .B(n14046), .Z(n14033) );
  AND U13842 ( .A(n14047), .B(n14048), .Z(n14046) );
  XOR U13843 ( .A(n14045), .B(n12234), .Z(n14048) );
  XOR U13844 ( .A(n14049), .B(n14050), .Z(n12234) );
  AND U13845 ( .A(n350), .B(n14051), .Z(n14050) );
  XOR U13846 ( .A(n14052), .B(n14049), .Z(n14051) );
  XNOR U13847 ( .A(n12231), .B(n14045), .Z(n14047) );
  XOR U13848 ( .A(n14053), .B(n14054), .Z(n12231) );
  AND U13849 ( .A(n347), .B(n14055), .Z(n14054) );
  XOR U13850 ( .A(n14056), .B(n14053), .Z(n14055) );
  XOR U13851 ( .A(n14057), .B(n14058), .Z(n14045) );
  AND U13852 ( .A(n14059), .B(n14060), .Z(n14058) );
  XOR U13853 ( .A(n14057), .B(n12246), .Z(n14060) );
  XOR U13854 ( .A(n14061), .B(n14062), .Z(n12246) );
  AND U13855 ( .A(n350), .B(n14063), .Z(n14062) );
  XOR U13856 ( .A(n14064), .B(n14061), .Z(n14063) );
  XNOR U13857 ( .A(n12243), .B(n14057), .Z(n14059) );
  XOR U13858 ( .A(n14065), .B(n14066), .Z(n12243) );
  AND U13859 ( .A(n347), .B(n14067), .Z(n14066) );
  XOR U13860 ( .A(n14068), .B(n14065), .Z(n14067) );
  XOR U13861 ( .A(n14069), .B(n14070), .Z(n14057) );
  AND U13862 ( .A(n14071), .B(n14072), .Z(n14070) );
  XOR U13863 ( .A(n14069), .B(n12258), .Z(n14072) );
  XOR U13864 ( .A(n14073), .B(n14074), .Z(n12258) );
  AND U13865 ( .A(n350), .B(n14075), .Z(n14074) );
  XOR U13866 ( .A(n14076), .B(n14073), .Z(n14075) );
  XNOR U13867 ( .A(n12255), .B(n14069), .Z(n14071) );
  XOR U13868 ( .A(n14077), .B(n14078), .Z(n12255) );
  AND U13869 ( .A(n347), .B(n14079), .Z(n14078) );
  XOR U13870 ( .A(n14080), .B(n14077), .Z(n14079) );
  XOR U13871 ( .A(n14081), .B(n14082), .Z(n14069) );
  AND U13872 ( .A(n14083), .B(n14084), .Z(n14082) );
  XOR U13873 ( .A(n14081), .B(n12270), .Z(n14084) );
  XOR U13874 ( .A(n14085), .B(n14086), .Z(n12270) );
  AND U13875 ( .A(n350), .B(n14087), .Z(n14086) );
  XOR U13876 ( .A(n14088), .B(n14085), .Z(n14087) );
  XNOR U13877 ( .A(n12267), .B(n14081), .Z(n14083) );
  XOR U13878 ( .A(n14089), .B(n14090), .Z(n12267) );
  AND U13879 ( .A(n347), .B(n14091), .Z(n14090) );
  XOR U13880 ( .A(n14092), .B(n14089), .Z(n14091) );
  XOR U13881 ( .A(n14093), .B(n14094), .Z(n14081) );
  AND U13882 ( .A(n14095), .B(n14096), .Z(n14094) );
  XOR U13883 ( .A(n14093), .B(n12282), .Z(n14096) );
  XOR U13884 ( .A(n14097), .B(n14098), .Z(n12282) );
  AND U13885 ( .A(n350), .B(n14099), .Z(n14098) );
  XOR U13886 ( .A(n14100), .B(n14097), .Z(n14099) );
  XNOR U13887 ( .A(n12279), .B(n14093), .Z(n14095) );
  XOR U13888 ( .A(n14101), .B(n14102), .Z(n12279) );
  AND U13889 ( .A(n347), .B(n14103), .Z(n14102) );
  XOR U13890 ( .A(n14104), .B(n14101), .Z(n14103) );
  XOR U13891 ( .A(n14105), .B(n14106), .Z(n14093) );
  AND U13892 ( .A(n14107), .B(n14108), .Z(n14106) );
  XOR U13893 ( .A(n14105), .B(n12294), .Z(n14108) );
  XOR U13894 ( .A(n14109), .B(n14110), .Z(n12294) );
  AND U13895 ( .A(n350), .B(n14111), .Z(n14110) );
  XOR U13896 ( .A(n14112), .B(n14109), .Z(n14111) );
  XNOR U13897 ( .A(n12291), .B(n14105), .Z(n14107) );
  XOR U13898 ( .A(n14113), .B(n14114), .Z(n12291) );
  AND U13899 ( .A(n347), .B(n14115), .Z(n14114) );
  XOR U13900 ( .A(n14116), .B(n14113), .Z(n14115) );
  XOR U13901 ( .A(n14117), .B(n14118), .Z(n14105) );
  AND U13902 ( .A(n14119), .B(n14120), .Z(n14118) );
  XOR U13903 ( .A(n12306), .B(n14117), .Z(n14120) );
  XOR U13904 ( .A(n14121), .B(n14122), .Z(n12306) );
  AND U13905 ( .A(n350), .B(n14123), .Z(n14122) );
  XOR U13906 ( .A(n14121), .B(n14124), .Z(n14123) );
  XNOR U13907 ( .A(n14117), .B(n12303), .Z(n14119) );
  XOR U13908 ( .A(n14125), .B(n14126), .Z(n12303) );
  AND U13909 ( .A(n347), .B(n14127), .Z(n14126) );
  XOR U13910 ( .A(n14125), .B(n14128), .Z(n14127) );
  XOR U13911 ( .A(n14129), .B(n14130), .Z(n14117) );
  AND U13912 ( .A(n14131), .B(n14132), .Z(n14130) );
  XNOR U13913 ( .A(n14133), .B(n12319), .Z(n14132) );
  XOR U13914 ( .A(n14134), .B(n14135), .Z(n12319) );
  AND U13915 ( .A(n350), .B(n14136), .Z(n14135) );
  XOR U13916 ( .A(n14137), .B(n14134), .Z(n14136) );
  XNOR U13917 ( .A(n12316), .B(n14129), .Z(n14131) );
  XOR U13918 ( .A(n14138), .B(n14139), .Z(n12316) );
  AND U13919 ( .A(n347), .B(n14140), .Z(n14139) );
  XOR U13920 ( .A(n14141), .B(n14138), .Z(n14140) );
  IV U13921 ( .A(n14133), .Z(n14129) );
  AND U13922 ( .A(n13765), .B(n13768), .Z(n14133) );
  XNOR U13923 ( .A(n14142), .B(n14143), .Z(n13768) );
  AND U13924 ( .A(n350), .B(n14144), .Z(n14143) );
  XNOR U13925 ( .A(n14145), .B(n14142), .Z(n14144) );
  XOR U13926 ( .A(n14146), .B(n14147), .Z(n350) );
  AND U13927 ( .A(n14148), .B(n14149), .Z(n14147) );
  XOR U13928 ( .A(n13776), .B(n14146), .Z(n14149) );
  IV U13929 ( .A(n14150), .Z(n13776) );
  AND U13930 ( .A(p_input[2303]), .B(p_input[2271]), .Z(n14150) );
  XOR U13931 ( .A(n14146), .B(n13773), .Z(n14148) );
  AND U13932 ( .A(p_input[2207]), .B(p_input[2239]), .Z(n13773) );
  XOR U13933 ( .A(n14151), .B(n14152), .Z(n14146) );
  AND U13934 ( .A(n14153), .B(n14154), .Z(n14152) );
  XOR U13935 ( .A(n14151), .B(n13788), .Z(n14154) );
  XNOR U13936 ( .A(p_input[2270]), .B(n14155), .Z(n13788) );
  AND U13937 ( .A(n282), .B(n14156), .Z(n14155) );
  XOR U13938 ( .A(p_input[2302]), .B(p_input[2270]), .Z(n14156) );
  XNOR U13939 ( .A(n13785), .B(n14151), .Z(n14153) );
  XOR U13940 ( .A(n14157), .B(n14158), .Z(n13785) );
  AND U13941 ( .A(n280), .B(n14159), .Z(n14158) );
  XOR U13942 ( .A(p_input[2238]), .B(p_input[2206]), .Z(n14159) );
  XOR U13943 ( .A(n14160), .B(n14161), .Z(n14151) );
  AND U13944 ( .A(n14162), .B(n14163), .Z(n14161) );
  XOR U13945 ( .A(n14160), .B(n13800), .Z(n14163) );
  XNOR U13946 ( .A(p_input[2269]), .B(n14164), .Z(n13800) );
  AND U13947 ( .A(n282), .B(n14165), .Z(n14164) );
  XOR U13948 ( .A(p_input[2301]), .B(p_input[2269]), .Z(n14165) );
  XNOR U13949 ( .A(n13797), .B(n14160), .Z(n14162) );
  XOR U13950 ( .A(n14166), .B(n14167), .Z(n13797) );
  AND U13951 ( .A(n280), .B(n14168), .Z(n14167) );
  XOR U13952 ( .A(p_input[2237]), .B(p_input[2205]), .Z(n14168) );
  XOR U13953 ( .A(n14169), .B(n14170), .Z(n14160) );
  AND U13954 ( .A(n14171), .B(n14172), .Z(n14170) );
  XOR U13955 ( .A(n14169), .B(n13812), .Z(n14172) );
  XNOR U13956 ( .A(p_input[2268]), .B(n14173), .Z(n13812) );
  AND U13957 ( .A(n282), .B(n14174), .Z(n14173) );
  XOR U13958 ( .A(p_input[2300]), .B(p_input[2268]), .Z(n14174) );
  XNOR U13959 ( .A(n13809), .B(n14169), .Z(n14171) );
  XOR U13960 ( .A(n14175), .B(n14176), .Z(n13809) );
  AND U13961 ( .A(n280), .B(n14177), .Z(n14176) );
  XOR U13962 ( .A(p_input[2236]), .B(p_input[2204]), .Z(n14177) );
  XOR U13963 ( .A(n14178), .B(n14179), .Z(n14169) );
  AND U13964 ( .A(n14180), .B(n14181), .Z(n14179) );
  XOR U13965 ( .A(n14178), .B(n13824), .Z(n14181) );
  XNOR U13966 ( .A(p_input[2267]), .B(n14182), .Z(n13824) );
  AND U13967 ( .A(n282), .B(n14183), .Z(n14182) );
  XOR U13968 ( .A(p_input[2299]), .B(p_input[2267]), .Z(n14183) );
  XNOR U13969 ( .A(n13821), .B(n14178), .Z(n14180) );
  XOR U13970 ( .A(n14184), .B(n14185), .Z(n13821) );
  AND U13971 ( .A(n280), .B(n14186), .Z(n14185) );
  XOR U13972 ( .A(p_input[2235]), .B(p_input[2203]), .Z(n14186) );
  XOR U13973 ( .A(n14187), .B(n14188), .Z(n14178) );
  AND U13974 ( .A(n14189), .B(n14190), .Z(n14188) );
  XOR U13975 ( .A(n14187), .B(n13836), .Z(n14190) );
  XNOR U13976 ( .A(p_input[2266]), .B(n14191), .Z(n13836) );
  AND U13977 ( .A(n282), .B(n14192), .Z(n14191) );
  XOR U13978 ( .A(p_input[2298]), .B(p_input[2266]), .Z(n14192) );
  XNOR U13979 ( .A(n13833), .B(n14187), .Z(n14189) );
  XOR U13980 ( .A(n14193), .B(n14194), .Z(n13833) );
  AND U13981 ( .A(n280), .B(n14195), .Z(n14194) );
  XOR U13982 ( .A(p_input[2234]), .B(p_input[2202]), .Z(n14195) );
  XOR U13983 ( .A(n14196), .B(n14197), .Z(n14187) );
  AND U13984 ( .A(n14198), .B(n14199), .Z(n14197) );
  XOR U13985 ( .A(n14196), .B(n13848), .Z(n14199) );
  XNOR U13986 ( .A(p_input[2265]), .B(n14200), .Z(n13848) );
  AND U13987 ( .A(n282), .B(n14201), .Z(n14200) );
  XOR U13988 ( .A(p_input[2297]), .B(p_input[2265]), .Z(n14201) );
  XNOR U13989 ( .A(n13845), .B(n14196), .Z(n14198) );
  XOR U13990 ( .A(n14202), .B(n14203), .Z(n13845) );
  AND U13991 ( .A(n280), .B(n14204), .Z(n14203) );
  XOR U13992 ( .A(p_input[2233]), .B(p_input[2201]), .Z(n14204) );
  XOR U13993 ( .A(n14205), .B(n14206), .Z(n14196) );
  AND U13994 ( .A(n14207), .B(n14208), .Z(n14206) );
  XOR U13995 ( .A(n14205), .B(n13860), .Z(n14208) );
  XNOR U13996 ( .A(p_input[2264]), .B(n14209), .Z(n13860) );
  AND U13997 ( .A(n282), .B(n14210), .Z(n14209) );
  XOR U13998 ( .A(p_input[2296]), .B(p_input[2264]), .Z(n14210) );
  XNOR U13999 ( .A(n13857), .B(n14205), .Z(n14207) );
  XOR U14000 ( .A(n14211), .B(n14212), .Z(n13857) );
  AND U14001 ( .A(n280), .B(n14213), .Z(n14212) );
  XOR U14002 ( .A(p_input[2232]), .B(p_input[2200]), .Z(n14213) );
  XOR U14003 ( .A(n14214), .B(n14215), .Z(n14205) );
  AND U14004 ( .A(n14216), .B(n14217), .Z(n14215) );
  XOR U14005 ( .A(n14214), .B(n13872), .Z(n14217) );
  XNOR U14006 ( .A(p_input[2263]), .B(n14218), .Z(n13872) );
  AND U14007 ( .A(n282), .B(n14219), .Z(n14218) );
  XOR U14008 ( .A(p_input[2295]), .B(p_input[2263]), .Z(n14219) );
  XNOR U14009 ( .A(n13869), .B(n14214), .Z(n14216) );
  XOR U14010 ( .A(n14220), .B(n14221), .Z(n13869) );
  AND U14011 ( .A(n280), .B(n14222), .Z(n14221) );
  XOR U14012 ( .A(p_input[2231]), .B(p_input[2199]), .Z(n14222) );
  XOR U14013 ( .A(n14223), .B(n14224), .Z(n14214) );
  AND U14014 ( .A(n14225), .B(n14226), .Z(n14224) );
  XOR U14015 ( .A(n14223), .B(n13884), .Z(n14226) );
  XNOR U14016 ( .A(p_input[2262]), .B(n14227), .Z(n13884) );
  AND U14017 ( .A(n282), .B(n14228), .Z(n14227) );
  XOR U14018 ( .A(p_input[2294]), .B(p_input[2262]), .Z(n14228) );
  XNOR U14019 ( .A(n13881), .B(n14223), .Z(n14225) );
  XOR U14020 ( .A(n14229), .B(n14230), .Z(n13881) );
  AND U14021 ( .A(n280), .B(n14231), .Z(n14230) );
  XOR U14022 ( .A(p_input[2230]), .B(p_input[2198]), .Z(n14231) );
  XOR U14023 ( .A(n14232), .B(n14233), .Z(n14223) );
  AND U14024 ( .A(n14234), .B(n14235), .Z(n14233) );
  XOR U14025 ( .A(n14232), .B(n13896), .Z(n14235) );
  XNOR U14026 ( .A(p_input[2261]), .B(n14236), .Z(n13896) );
  AND U14027 ( .A(n282), .B(n14237), .Z(n14236) );
  XOR U14028 ( .A(p_input[2293]), .B(p_input[2261]), .Z(n14237) );
  XNOR U14029 ( .A(n13893), .B(n14232), .Z(n14234) );
  XOR U14030 ( .A(n14238), .B(n14239), .Z(n13893) );
  AND U14031 ( .A(n280), .B(n14240), .Z(n14239) );
  XOR U14032 ( .A(p_input[2229]), .B(p_input[2197]), .Z(n14240) );
  XOR U14033 ( .A(n14241), .B(n14242), .Z(n14232) );
  AND U14034 ( .A(n14243), .B(n14244), .Z(n14242) );
  XOR U14035 ( .A(n14241), .B(n13908), .Z(n14244) );
  XNOR U14036 ( .A(p_input[2260]), .B(n14245), .Z(n13908) );
  AND U14037 ( .A(n282), .B(n14246), .Z(n14245) );
  XOR U14038 ( .A(p_input[2292]), .B(p_input[2260]), .Z(n14246) );
  XNOR U14039 ( .A(n13905), .B(n14241), .Z(n14243) );
  XOR U14040 ( .A(n14247), .B(n14248), .Z(n13905) );
  AND U14041 ( .A(n280), .B(n14249), .Z(n14248) );
  XOR U14042 ( .A(p_input[2228]), .B(p_input[2196]), .Z(n14249) );
  XOR U14043 ( .A(n14250), .B(n14251), .Z(n14241) );
  AND U14044 ( .A(n14252), .B(n14253), .Z(n14251) );
  XOR U14045 ( .A(n14250), .B(n13920), .Z(n14253) );
  XNOR U14046 ( .A(p_input[2259]), .B(n14254), .Z(n13920) );
  AND U14047 ( .A(n282), .B(n14255), .Z(n14254) );
  XOR U14048 ( .A(p_input[2291]), .B(p_input[2259]), .Z(n14255) );
  XNOR U14049 ( .A(n13917), .B(n14250), .Z(n14252) );
  XOR U14050 ( .A(n14256), .B(n14257), .Z(n13917) );
  AND U14051 ( .A(n280), .B(n14258), .Z(n14257) );
  XOR U14052 ( .A(p_input[2227]), .B(p_input[2195]), .Z(n14258) );
  XOR U14053 ( .A(n14259), .B(n14260), .Z(n14250) );
  AND U14054 ( .A(n14261), .B(n14262), .Z(n14260) );
  XOR U14055 ( .A(n14259), .B(n13932), .Z(n14262) );
  XNOR U14056 ( .A(p_input[2258]), .B(n14263), .Z(n13932) );
  AND U14057 ( .A(n282), .B(n14264), .Z(n14263) );
  XOR U14058 ( .A(p_input[2290]), .B(p_input[2258]), .Z(n14264) );
  XNOR U14059 ( .A(n13929), .B(n14259), .Z(n14261) );
  XOR U14060 ( .A(n14265), .B(n14266), .Z(n13929) );
  AND U14061 ( .A(n280), .B(n14267), .Z(n14266) );
  XOR U14062 ( .A(p_input[2226]), .B(p_input[2194]), .Z(n14267) );
  XOR U14063 ( .A(n14268), .B(n14269), .Z(n14259) );
  AND U14064 ( .A(n14270), .B(n14271), .Z(n14269) );
  XOR U14065 ( .A(n14268), .B(n13944), .Z(n14271) );
  XNOR U14066 ( .A(p_input[2257]), .B(n14272), .Z(n13944) );
  AND U14067 ( .A(n282), .B(n14273), .Z(n14272) );
  XOR U14068 ( .A(p_input[2289]), .B(p_input[2257]), .Z(n14273) );
  XNOR U14069 ( .A(n13941), .B(n14268), .Z(n14270) );
  XOR U14070 ( .A(n14274), .B(n14275), .Z(n13941) );
  AND U14071 ( .A(n280), .B(n14276), .Z(n14275) );
  XOR U14072 ( .A(p_input[2225]), .B(p_input[2193]), .Z(n14276) );
  XOR U14073 ( .A(n14277), .B(n14278), .Z(n14268) );
  AND U14074 ( .A(n14279), .B(n14280), .Z(n14278) );
  XOR U14075 ( .A(n14277), .B(n13956), .Z(n14280) );
  XNOR U14076 ( .A(p_input[2256]), .B(n14281), .Z(n13956) );
  AND U14077 ( .A(n282), .B(n14282), .Z(n14281) );
  XOR U14078 ( .A(p_input[2288]), .B(p_input[2256]), .Z(n14282) );
  XNOR U14079 ( .A(n13953), .B(n14277), .Z(n14279) );
  XOR U14080 ( .A(n14283), .B(n14284), .Z(n13953) );
  AND U14081 ( .A(n280), .B(n14285), .Z(n14284) );
  XOR U14082 ( .A(p_input[2224]), .B(p_input[2192]), .Z(n14285) );
  XOR U14083 ( .A(n14286), .B(n14287), .Z(n14277) );
  AND U14084 ( .A(n14288), .B(n14289), .Z(n14287) );
  XOR U14085 ( .A(n14286), .B(n13968), .Z(n14289) );
  XNOR U14086 ( .A(p_input[2255]), .B(n14290), .Z(n13968) );
  AND U14087 ( .A(n282), .B(n14291), .Z(n14290) );
  XOR U14088 ( .A(p_input[2287]), .B(p_input[2255]), .Z(n14291) );
  XNOR U14089 ( .A(n13965), .B(n14286), .Z(n14288) );
  XOR U14090 ( .A(n14292), .B(n14293), .Z(n13965) );
  AND U14091 ( .A(n280), .B(n14294), .Z(n14293) );
  XOR U14092 ( .A(p_input[2223]), .B(p_input[2191]), .Z(n14294) );
  XOR U14093 ( .A(n14295), .B(n14296), .Z(n14286) );
  AND U14094 ( .A(n14297), .B(n14298), .Z(n14296) );
  XOR U14095 ( .A(n14295), .B(n13980), .Z(n14298) );
  XNOR U14096 ( .A(p_input[2254]), .B(n14299), .Z(n13980) );
  AND U14097 ( .A(n282), .B(n14300), .Z(n14299) );
  XOR U14098 ( .A(p_input[2286]), .B(p_input[2254]), .Z(n14300) );
  XNOR U14099 ( .A(n13977), .B(n14295), .Z(n14297) );
  XOR U14100 ( .A(n14301), .B(n14302), .Z(n13977) );
  AND U14101 ( .A(n280), .B(n14303), .Z(n14302) );
  XOR U14102 ( .A(p_input[2222]), .B(p_input[2190]), .Z(n14303) );
  XOR U14103 ( .A(n14304), .B(n14305), .Z(n14295) );
  AND U14104 ( .A(n14306), .B(n14307), .Z(n14305) );
  XOR U14105 ( .A(n14304), .B(n13992), .Z(n14307) );
  XNOR U14106 ( .A(p_input[2253]), .B(n14308), .Z(n13992) );
  AND U14107 ( .A(n282), .B(n14309), .Z(n14308) );
  XOR U14108 ( .A(p_input[2285]), .B(p_input[2253]), .Z(n14309) );
  XNOR U14109 ( .A(n13989), .B(n14304), .Z(n14306) );
  XOR U14110 ( .A(n14310), .B(n14311), .Z(n13989) );
  AND U14111 ( .A(n280), .B(n14312), .Z(n14311) );
  XOR U14112 ( .A(p_input[2221]), .B(p_input[2189]), .Z(n14312) );
  XOR U14113 ( .A(n14313), .B(n14314), .Z(n14304) );
  AND U14114 ( .A(n14315), .B(n14316), .Z(n14314) );
  XOR U14115 ( .A(n14313), .B(n14004), .Z(n14316) );
  XNOR U14116 ( .A(p_input[2252]), .B(n14317), .Z(n14004) );
  AND U14117 ( .A(n282), .B(n14318), .Z(n14317) );
  XOR U14118 ( .A(p_input[2284]), .B(p_input[2252]), .Z(n14318) );
  XNOR U14119 ( .A(n14001), .B(n14313), .Z(n14315) );
  XOR U14120 ( .A(n14319), .B(n14320), .Z(n14001) );
  AND U14121 ( .A(n280), .B(n14321), .Z(n14320) );
  XOR U14122 ( .A(p_input[2220]), .B(p_input[2188]), .Z(n14321) );
  XOR U14123 ( .A(n14322), .B(n14323), .Z(n14313) );
  AND U14124 ( .A(n14324), .B(n14325), .Z(n14323) );
  XOR U14125 ( .A(n14322), .B(n14016), .Z(n14325) );
  XNOR U14126 ( .A(p_input[2251]), .B(n14326), .Z(n14016) );
  AND U14127 ( .A(n282), .B(n14327), .Z(n14326) );
  XOR U14128 ( .A(p_input[2283]), .B(p_input[2251]), .Z(n14327) );
  XNOR U14129 ( .A(n14013), .B(n14322), .Z(n14324) );
  XOR U14130 ( .A(n14328), .B(n14329), .Z(n14013) );
  AND U14131 ( .A(n280), .B(n14330), .Z(n14329) );
  XOR U14132 ( .A(p_input[2219]), .B(p_input[2187]), .Z(n14330) );
  XOR U14133 ( .A(n14331), .B(n14332), .Z(n14322) );
  AND U14134 ( .A(n14333), .B(n14334), .Z(n14332) );
  XOR U14135 ( .A(n14331), .B(n14028), .Z(n14334) );
  XNOR U14136 ( .A(p_input[2250]), .B(n14335), .Z(n14028) );
  AND U14137 ( .A(n282), .B(n14336), .Z(n14335) );
  XOR U14138 ( .A(p_input[2282]), .B(p_input[2250]), .Z(n14336) );
  XNOR U14139 ( .A(n14025), .B(n14331), .Z(n14333) );
  XOR U14140 ( .A(n14337), .B(n14338), .Z(n14025) );
  AND U14141 ( .A(n280), .B(n14339), .Z(n14338) );
  XOR U14142 ( .A(p_input[2218]), .B(p_input[2186]), .Z(n14339) );
  XOR U14143 ( .A(n14340), .B(n14341), .Z(n14331) );
  AND U14144 ( .A(n14342), .B(n14343), .Z(n14341) );
  XOR U14145 ( .A(n14340), .B(n14040), .Z(n14343) );
  XNOR U14146 ( .A(p_input[2249]), .B(n14344), .Z(n14040) );
  AND U14147 ( .A(n282), .B(n14345), .Z(n14344) );
  XOR U14148 ( .A(p_input[2281]), .B(p_input[2249]), .Z(n14345) );
  XNOR U14149 ( .A(n14037), .B(n14340), .Z(n14342) );
  XOR U14150 ( .A(n14346), .B(n14347), .Z(n14037) );
  AND U14151 ( .A(n280), .B(n14348), .Z(n14347) );
  XOR U14152 ( .A(p_input[2217]), .B(p_input[2185]), .Z(n14348) );
  XOR U14153 ( .A(n14349), .B(n14350), .Z(n14340) );
  AND U14154 ( .A(n14351), .B(n14352), .Z(n14350) );
  XOR U14155 ( .A(n14349), .B(n14052), .Z(n14352) );
  XNOR U14156 ( .A(p_input[2248]), .B(n14353), .Z(n14052) );
  AND U14157 ( .A(n282), .B(n14354), .Z(n14353) );
  XOR U14158 ( .A(p_input[2280]), .B(p_input[2248]), .Z(n14354) );
  XNOR U14159 ( .A(n14049), .B(n14349), .Z(n14351) );
  XOR U14160 ( .A(n14355), .B(n14356), .Z(n14049) );
  AND U14161 ( .A(n280), .B(n14357), .Z(n14356) );
  XOR U14162 ( .A(p_input[2216]), .B(p_input[2184]), .Z(n14357) );
  XOR U14163 ( .A(n14358), .B(n14359), .Z(n14349) );
  AND U14164 ( .A(n14360), .B(n14361), .Z(n14359) );
  XOR U14165 ( .A(n14358), .B(n14064), .Z(n14361) );
  XNOR U14166 ( .A(p_input[2247]), .B(n14362), .Z(n14064) );
  AND U14167 ( .A(n282), .B(n14363), .Z(n14362) );
  XOR U14168 ( .A(p_input[2279]), .B(p_input[2247]), .Z(n14363) );
  XNOR U14169 ( .A(n14061), .B(n14358), .Z(n14360) );
  XOR U14170 ( .A(n14364), .B(n14365), .Z(n14061) );
  AND U14171 ( .A(n280), .B(n14366), .Z(n14365) );
  XOR U14172 ( .A(p_input[2215]), .B(p_input[2183]), .Z(n14366) );
  XOR U14173 ( .A(n14367), .B(n14368), .Z(n14358) );
  AND U14174 ( .A(n14369), .B(n14370), .Z(n14368) );
  XOR U14175 ( .A(n14367), .B(n14076), .Z(n14370) );
  XNOR U14176 ( .A(p_input[2246]), .B(n14371), .Z(n14076) );
  AND U14177 ( .A(n282), .B(n14372), .Z(n14371) );
  XOR U14178 ( .A(p_input[2278]), .B(p_input[2246]), .Z(n14372) );
  XNOR U14179 ( .A(n14073), .B(n14367), .Z(n14369) );
  XOR U14180 ( .A(n14373), .B(n14374), .Z(n14073) );
  AND U14181 ( .A(n280), .B(n14375), .Z(n14374) );
  XOR U14182 ( .A(p_input[2214]), .B(p_input[2182]), .Z(n14375) );
  XOR U14183 ( .A(n14376), .B(n14377), .Z(n14367) );
  AND U14184 ( .A(n14378), .B(n14379), .Z(n14377) );
  XOR U14185 ( .A(n14376), .B(n14088), .Z(n14379) );
  XNOR U14186 ( .A(p_input[2245]), .B(n14380), .Z(n14088) );
  AND U14187 ( .A(n282), .B(n14381), .Z(n14380) );
  XOR U14188 ( .A(p_input[2277]), .B(p_input[2245]), .Z(n14381) );
  XNOR U14189 ( .A(n14085), .B(n14376), .Z(n14378) );
  XOR U14190 ( .A(n14382), .B(n14383), .Z(n14085) );
  AND U14191 ( .A(n280), .B(n14384), .Z(n14383) );
  XOR U14192 ( .A(p_input[2213]), .B(p_input[2181]), .Z(n14384) );
  XOR U14193 ( .A(n14385), .B(n14386), .Z(n14376) );
  AND U14194 ( .A(n14387), .B(n14388), .Z(n14386) );
  XOR U14195 ( .A(n14385), .B(n14100), .Z(n14388) );
  XNOR U14196 ( .A(p_input[2244]), .B(n14389), .Z(n14100) );
  AND U14197 ( .A(n282), .B(n14390), .Z(n14389) );
  XOR U14198 ( .A(p_input[2276]), .B(p_input[2244]), .Z(n14390) );
  XNOR U14199 ( .A(n14097), .B(n14385), .Z(n14387) );
  XOR U14200 ( .A(n14391), .B(n14392), .Z(n14097) );
  AND U14201 ( .A(n280), .B(n14393), .Z(n14392) );
  XOR U14202 ( .A(p_input[2212]), .B(p_input[2180]), .Z(n14393) );
  XOR U14203 ( .A(n14394), .B(n14395), .Z(n14385) );
  AND U14204 ( .A(n14396), .B(n14397), .Z(n14395) );
  XOR U14205 ( .A(n14394), .B(n14112), .Z(n14397) );
  XNOR U14206 ( .A(p_input[2243]), .B(n14398), .Z(n14112) );
  AND U14207 ( .A(n282), .B(n14399), .Z(n14398) );
  XOR U14208 ( .A(p_input[2275]), .B(p_input[2243]), .Z(n14399) );
  XNOR U14209 ( .A(n14109), .B(n14394), .Z(n14396) );
  XOR U14210 ( .A(n14400), .B(n14401), .Z(n14109) );
  AND U14211 ( .A(n280), .B(n14402), .Z(n14401) );
  XOR U14212 ( .A(p_input[2211]), .B(p_input[2179]), .Z(n14402) );
  XOR U14213 ( .A(n14403), .B(n14404), .Z(n14394) );
  AND U14214 ( .A(n14405), .B(n14406), .Z(n14404) );
  XOR U14215 ( .A(n14124), .B(n14403), .Z(n14406) );
  XNOR U14216 ( .A(p_input[2242]), .B(n14407), .Z(n14124) );
  AND U14217 ( .A(n282), .B(n14408), .Z(n14407) );
  XOR U14218 ( .A(p_input[2274]), .B(p_input[2242]), .Z(n14408) );
  XNOR U14219 ( .A(n14403), .B(n14121), .Z(n14405) );
  XOR U14220 ( .A(n14409), .B(n14410), .Z(n14121) );
  AND U14221 ( .A(n280), .B(n14411), .Z(n14410) );
  XOR U14222 ( .A(p_input[2210]), .B(p_input[2178]), .Z(n14411) );
  XOR U14223 ( .A(n14412), .B(n14413), .Z(n14403) );
  AND U14224 ( .A(n14414), .B(n14415), .Z(n14413) );
  XNOR U14225 ( .A(n14416), .B(n14137), .Z(n14415) );
  XNOR U14226 ( .A(p_input[2241]), .B(n14417), .Z(n14137) );
  AND U14227 ( .A(n282), .B(n14418), .Z(n14417) );
  XNOR U14228 ( .A(p_input[2273]), .B(n14419), .Z(n14418) );
  IV U14229 ( .A(p_input[2241]), .Z(n14419) );
  XNOR U14230 ( .A(n14134), .B(n14412), .Z(n14414) );
  XNOR U14231 ( .A(p_input[2177]), .B(n14420), .Z(n14134) );
  AND U14232 ( .A(n280), .B(n14421), .Z(n14420) );
  XOR U14233 ( .A(p_input[2209]), .B(p_input[2177]), .Z(n14421) );
  IV U14234 ( .A(n14416), .Z(n14412) );
  AND U14235 ( .A(n14142), .B(n14145), .Z(n14416) );
  XOR U14236 ( .A(p_input[2240]), .B(n14422), .Z(n14145) );
  AND U14237 ( .A(n282), .B(n14423), .Z(n14422) );
  XOR U14238 ( .A(p_input[2272]), .B(p_input[2240]), .Z(n14423) );
  XOR U14239 ( .A(n14424), .B(n14425), .Z(n282) );
  AND U14240 ( .A(n14426), .B(n14427), .Z(n14425) );
  XNOR U14241 ( .A(p_input[2303]), .B(n14424), .Z(n14427) );
  XOR U14242 ( .A(n14424), .B(p_input[2271]), .Z(n14426) );
  XOR U14243 ( .A(n14428), .B(n14429), .Z(n14424) );
  AND U14244 ( .A(n14430), .B(n14431), .Z(n14429) );
  XNOR U14245 ( .A(p_input[2302]), .B(n14428), .Z(n14431) );
  XOR U14246 ( .A(n14428), .B(p_input[2270]), .Z(n14430) );
  XOR U14247 ( .A(n14432), .B(n14433), .Z(n14428) );
  AND U14248 ( .A(n14434), .B(n14435), .Z(n14433) );
  XNOR U14249 ( .A(p_input[2301]), .B(n14432), .Z(n14435) );
  XOR U14250 ( .A(n14432), .B(p_input[2269]), .Z(n14434) );
  XOR U14251 ( .A(n14436), .B(n14437), .Z(n14432) );
  AND U14252 ( .A(n14438), .B(n14439), .Z(n14437) );
  XNOR U14253 ( .A(p_input[2300]), .B(n14436), .Z(n14439) );
  XOR U14254 ( .A(n14436), .B(p_input[2268]), .Z(n14438) );
  XOR U14255 ( .A(n14440), .B(n14441), .Z(n14436) );
  AND U14256 ( .A(n14442), .B(n14443), .Z(n14441) );
  XNOR U14257 ( .A(p_input[2299]), .B(n14440), .Z(n14443) );
  XOR U14258 ( .A(n14440), .B(p_input[2267]), .Z(n14442) );
  XOR U14259 ( .A(n14444), .B(n14445), .Z(n14440) );
  AND U14260 ( .A(n14446), .B(n14447), .Z(n14445) );
  XNOR U14261 ( .A(p_input[2298]), .B(n14444), .Z(n14447) );
  XOR U14262 ( .A(n14444), .B(p_input[2266]), .Z(n14446) );
  XOR U14263 ( .A(n14448), .B(n14449), .Z(n14444) );
  AND U14264 ( .A(n14450), .B(n14451), .Z(n14449) );
  XNOR U14265 ( .A(p_input[2297]), .B(n14448), .Z(n14451) );
  XOR U14266 ( .A(n14448), .B(p_input[2265]), .Z(n14450) );
  XOR U14267 ( .A(n14452), .B(n14453), .Z(n14448) );
  AND U14268 ( .A(n14454), .B(n14455), .Z(n14453) );
  XNOR U14269 ( .A(p_input[2296]), .B(n14452), .Z(n14455) );
  XOR U14270 ( .A(n14452), .B(p_input[2264]), .Z(n14454) );
  XOR U14271 ( .A(n14456), .B(n14457), .Z(n14452) );
  AND U14272 ( .A(n14458), .B(n14459), .Z(n14457) );
  XNOR U14273 ( .A(p_input[2295]), .B(n14456), .Z(n14459) );
  XOR U14274 ( .A(n14456), .B(p_input[2263]), .Z(n14458) );
  XOR U14275 ( .A(n14460), .B(n14461), .Z(n14456) );
  AND U14276 ( .A(n14462), .B(n14463), .Z(n14461) );
  XNOR U14277 ( .A(p_input[2294]), .B(n14460), .Z(n14463) );
  XOR U14278 ( .A(n14460), .B(p_input[2262]), .Z(n14462) );
  XOR U14279 ( .A(n14464), .B(n14465), .Z(n14460) );
  AND U14280 ( .A(n14466), .B(n14467), .Z(n14465) );
  XNOR U14281 ( .A(p_input[2293]), .B(n14464), .Z(n14467) );
  XOR U14282 ( .A(n14464), .B(p_input[2261]), .Z(n14466) );
  XOR U14283 ( .A(n14468), .B(n14469), .Z(n14464) );
  AND U14284 ( .A(n14470), .B(n14471), .Z(n14469) );
  XNOR U14285 ( .A(p_input[2292]), .B(n14468), .Z(n14471) );
  XOR U14286 ( .A(n14468), .B(p_input[2260]), .Z(n14470) );
  XOR U14287 ( .A(n14472), .B(n14473), .Z(n14468) );
  AND U14288 ( .A(n14474), .B(n14475), .Z(n14473) );
  XNOR U14289 ( .A(p_input[2291]), .B(n14472), .Z(n14475) );
  XOR U14290 ( .A(n14472), .B(p_input[2259]), .Z(n14474) );
  XOR U14291 ( .A(n14476), .B(n14477), .Z(n14472) );
  AND U14292 ( .A(n14478), .B(n14479), .Z(n14477) );
  XNOR U14293 ( .A(p_input[2290]), .B(n14476), .Z(n14479) );
  XOR U14294 ( .A(n14476), .B(p_input[2258]), .Z(n14478) );
  XOR U14295 ( .A(n14480), .B(n14481), .Z(n14476) );
  AND U14296 ( .A(n14482), .B(n14483), .Z(n14481) );
  XNOR U14297 ( .A(p_input[2289]), .B(n14480), .Z(n14483) );
  XOR U14298 ( .A(n14480), .B(p_input[2257]), .Z(n14482) );
  XOR U14299 ( .A(n14484), .B(n14485), .Z(n14480) );
  AND U14300 ( .A(n14486), .B(n14487), .Z(n14485) );
  XNOR U14301 ( .A(p_input[2288]), .B(n14484), .Z(n14487) );
  XOR U14302 ( .A(n14484), .B(p_input[2256]), .Z(n14486) );
  XOR U14303 ( .A(n14488), .B(n14489), .Z(n14484) );
  AND U14304 ( .A(n14490), .B(n14491), .Z(n14489) );
  XNOR U14305 ( .A(p_input[2287]), .B(n14488), .Z(n14491) );
  XOR U14306 ( .A(n14488), .B(p_input[2255]), .Z(n14490) );
  XOR U14307 ( .A(n14492), .B(n14493), .Z(n14488) );
  AND U14308 ( .A(n14494), .B(n14495), .Z(n14493) );
  XNOR U14309 ( .A(p_input[2286]), .B(n14492), .Z(n14495) );
  XOR U14310 ( .A(n14492), .B(p_input[2254]), .Z(n14494) );
  XOR U14311 ( .A(n14496), .B(n14497), .Z(n14492) );
  AND U14312 ( .A(n14498), .B(n14499), .Z(n14497) );
  XNOR U14313 ( .A(p_input[2285]), .B(n14496), .Z(n14499) );
  XOR U14314 ( .A(n14496), .B(p_input[2253]), .Z(n14498) );
  XOR U14315 ( .A(n14500), .B(n14501), .Z(n14496) );
  AND U14316 ( .A(n14502), .B(n14503), .Z(n14501) );
  XNOR U14317 ( .A(p_input[2284]), .B(n14500), .Z(n14503) );
  XOR U14318 ( .A(n14500), .B(p_input[2252]), .Z(n14502) );
  XOR U14319 ( .A(n14504), .B(n14505), .Z(n14500) );
  AND U14320 ( .A(n14506), .B(n14507), .Z(n14505) );
  XNOR U14321 ( .A(p_input[2283]), .B(n14504), .Z(n14507) );
  XOR U14322 ( .A(n14504), .B(p_input[2251]), .Z(n14506) );
  XOR U14323 ( .A(n14508), .B(n14509), .Z(n14504) );
  AND U14324 ( .A(n14510), .B(n14511), .Z(n14509) );
  XNOR U14325 ( .A(p_input[2282]), .B(n14508), .Z(n14511) );
  XOR U14326 ( .A(n14508), .B(p_input[2250]), .Z(n14510) );
  XOR U14327 ( .A(n14512), .B(n14513), .Z(n14508) );
  AND U14328 ( .A(n14514), .B(n14515), .Z(n14513) );
  XNOR U14329 ( .A(p_input[2281]), .B(n14512), .Z(n14515) );
  XOR U14330 ( .A(n14512), .B(p_input[2249]), .Z(n14514) );
  XOR U14331 ( .A(n14516), .B(n14517), .Z(n14512) );
  AND U14332 ( .A(n14518), .B(n14519), .Z(n14517) );
  XNOR U14333 ( .A(p_input[2280]), .B(n14516), .Z(n14519) );
  XOR U14334 ( .A(n14516), .B(p_input[2248]), .Z(n14518) );
  XOR U14335 ( .A(n14520), .B(n14521), .Z(n14516) );
  AND U14336 ( .A(n14522), .B(n14523), .Z(n14521) );
  XNOR U14337 ( .A(p_input[2279]), .B(n14520), .Z(n14523) );
  XOR U14338 ( .A(n14520), .B(p_input[2247]), .Z(n14522) );
  XOR U14339 ( .A(n14524), .B(n14525), .Z(n14520) );
  AND U14340 ( .A(n14526), .B(n14527), .Z(n14525) );
  XNOR U14341 ( .A(p_input[2278]), .B(n14524), .Z(n14527) );
  XOR U14342 ( .A(n14524), .B(p_input[2246]), .Z(n14526) );
  XOR U14343 ( .A(n14528), .B(n14529), .Z(n14524) );
  AND U14344 ( .A(n14530), .B(n14531), .Z(n14529) );
  XNOR U14345 ( .A(p_input[2277]), .B(n14528), .Z(n14531) );
  XOR U14346 ( .A(n14528), .B(p_input[2245]), .Z(n14530) );
  XOR U14347 ( .A(n14532), .B(n14533), .Z(n14528) );
  AND U14348 ( .A(n14534), .B(n14535), .Z(n14533) );
  XNOR U14349 ( .A(p_input[2276]), .B(n14532), .Z(n14535) );
  XOR U14350 ( .A(n14532), .B(p_input[2244]), .Z(n14534) );
  XOR U14351 ( .A(n14536), .B(n14537), .Z(n14532) );
  AND U14352 ( .A(n14538), .B(n14539), .Z(n14537) );
  XNOR U14353 ( .A(p_input[2275]), .B(n14536), .Z(n14539) );
  XOR U14354 ( .A(n14536), .B(p_input[2243]), .Z(n14538) );
  XOR U14355 ( .A(n14540), .B(n14541), .Z(n14536) );
  AND U14356 ( .A(n14542), .B(n14543), .Z(n14541) );
  XNOR U14357 ( .A(p_input[2274]), .B(n14540), .Z(n14543) );
  XOR U14358 ( .A(n14540), .B(p_input[2242]), .Z(n14542) );
  XNOR U14359 ( .A(n14544), .B(n14545), .Z(n14540) );
  AND U14360 ( .A(n14546), .B(n14547), .Z(n14545) );
  XOR U14361 ( .A(p_input[2273]), .B(n14544), .Z(n14547) );
  XNOR U14362 ( .A(p_input[2241]), .B(n14544), .Z(n14546) );
  AND U14363 ( .A(p_input[2272]), .B(n14548), .Z(n14544) );
  IV U14364 ( .A(p_input[2240]), .Z(n14548) );
  XNOR U14365 ( .A(p_input[2176]), .B(n14549), .Z(n14142) );
  AND U14366 ( .A(n280), .B(n14550), .Z(n14549) );
  XOR U14367 ( .A(p_input[2208]), .B(p_input[2176]), .Z(n14550) );
  XOR U14368 ( .A(n14551), .B(n14552), .Z(n280) );
  AND U14369 ( .A(n14553), .B(n14554), .Z(n14552) );
  XNOR U14370 ( .A(p_input[2239]), .B(n14551), .Z(n14554) );
  XOR U14371 ( .A(n14551), .B(p_input[2207]), .Z(n14553) );
  XOR U14372 ( .A(n14555), .B(n14556), .Z(n14551) );
  AND U14373 ( .A(n14557), .B(n14558), .Z(n14556) );
  XNOR U14374 ( .A(p_input[2238]), .B(n14555), .Z(n14558) );
  XNOR U14375 ( .A(n14555), .B(n14157), .Z(n14557) );
  IV U14376 ( .A(p_input[2206]), .Z(n14157) );
  XOR U14377 ( .A(n14559), .B(n14560), .Z(n14555) );
  AND U14378 ( .A(n14561), .B(n14562), .Z(n14560) );
  XNOR U14379 ( .A(p_input[2237]), .B(n14559), .Z(n14562) );
  XNOR U14380 ( .A(n14559), .B(n14166), .Z(n14561) );
  IV U14381 ( .A(p_input[2205]), .Z(n14166) );
  XOR U14382 ( .A(n14563), .B(n14564), .Z(n14559) );
  AND U14383 ( .A(n14565), .B(n14566), .Z(n14564) );
  XNOR U14384 ( .A(p_input[2236]), .B(n14563), .Z(n14566) );
  XNOR U14385 ( .A(n14563), .B(n14175), .Z(n14565) );
  IV U14386 ( .A(p_input[2204]), .Z(n14175) );
  XOR U14387 ( .A(n14567), .B(n14568), .Z(n14563) );
  AND U14388 ( .A(n14569), .B(n14570), .Z(n14568) );
  XNOR U14389 ( .A(p_input[2235]), .B(n14567), .Z(n14570) );
  XNOR U14390 ( .A(n14567), .B(n14184), .Z(n14569) );
  IV U14391 ( .A(p_input[2203]), .Z(n14184) );
  XOR U14392 ( .A(n14571), .B(n14572), .Z(n14567) );
  AND U14393 ( .A(n14573), .B(n14574), .Z(n14572) );
  XNOR U14394 ( .A(p_input[2234]), .B(n14571), .Z(n14574) );
  XNOR U14395 ( .A(n14571), .B(n14193), .Z(n14573) );
  IV U14396 ( .A(p_input[2202]), .Z(n14193) );
  XOR U14397 ( .A(n14575), .B(n14576), .Z(n14571) );
  AND U14398 ( .A(n14577), .B(n14578), .Z(n14576) );
  XNOR U14399 ( .A(p_input[2233]), .B(n14575), .Z(n14578) );
  XNOR U14400 ( .A(n14575), .B(n14202), .Z(n14577) );
  IV U14401 ( .A(p_input[2201]), .Z(n14202) );
  XOR U14402 ( .A(n14579), .B(n14580), .Z(n14575) );
  AND U14403 ( .A(n14581), .B(n14582), .Z(n14580) );
  XNOR U14404 ( .A(p_input[2232]), .B(n14579), .Z(n14582) );
  XNOR U14405 ( .A(n14579), .B(n14211), .Z(n14581) );
  IV U14406 ( .A(p_input[2200]), .Z(n14211) );
  XOR U14407 ( .A(n14583), .B(n14584), .Z(n14579) );
  AND U14408 ( .A(n14585), .B(n14586), .Z(n14584) );
  XNOR U14409 ( .A(p_input[2231]), .B(n14583), .Z(n14586) );
  XNOR U14410 ( .A(n14583), .B(n14220), .Z(n14585) );
  IV U14411 ( .A(p_input[2199]), .Z(n14220) );
  XOR U14412 ( .A(n14587), .B(n14588), .Z(n14583) );
  AND U14413 ( .A(n14589), .B(n14590), .Z(n14588) );
  XNOR U14414 ( .A(p_input[2230]), .B(n14587), .Z(n14590) );
  XNOR U14415 ( .A(n14587), .B(n14229), .Z(n14589) );
  IV U14416 ( .A(p_input[2198]), .Z(n14229) );
  XOR U14417 ( .A(n14591), .B(n14592), .Z(n14587) );
  AND U14418 ( .A(n14593), .B(n14594), .Z(n14592) );
  XNOR U14419 ( .A(p_input[2229]), .B(n14591), .Z(n14594) );
  XNOR U14420 ( .A(n14591), .B(n14238), .Z(n14593) );
  IV U14421 ( .A(p_input[2197]), .Z(n14238) );
  XOR U14422 ( .A(n14595), .B(n14596), .Z(n14591) );
  AND U14423 ( .A(n14597), .B(n14598), .Z(n14596) );
  XNOR U14424 ( .A(p_input[2228]), .B(n14595), .Z(n14598) );
  XNOR U14425 ( .A(n14595), .B(n14247), .Z(n14597) );
  IV U14426 ( .A(p_input[2196]), .Z(n14247) );
  XOR U14427 ( .A(n14599), .B(n14600), .Z(n14595) );
  AND U14428 ( .A(n14601), .B(n14602), .Z(n14600) );
  XNOR U14429 ( .A(p_input[2227]), .B(n14599), .Z(n14602) );
  XNOR U14430 ( .A(n14599), .B(n14256), .Z(n14601) );
  IV U14431 ( .A(p_input[2195]), .Z(n14256) );
  XOR U14432 ( .A(n14603), .B(n14604), .Z(n14599) );
  AND U14433 ( .A(n14605), .B(n14606), .Z(n14604) );
  XNOR U14434 ( .A(p_input[2226]), .B(n14603), .Z(n14606) );
  XNOR U14435 ( .A(n14603), .B(n14265), .Z(n14605) );
  IV U14436 ( .A(p_input[2194]), .Z(n14265) );
  XOR U14437 ( .A(n14607), .B(n14608), .Z(n14603) );
  AND U14438 ( .A(n14609), .B(n14610), .Z(n14608) );
  XNOR U14439 ( .A(p_input[2225]), .B(n14607), .Z(n14610) );
  XNOR U14440 ( .A(n14607), .B(n14274), .Z(n14609) );
  IV U14441 ( .A(p_input[2193]), .Z(n14274) );
  XOR U14442 ( .A(n14611), .B(n14612), .Z(n14607) );
  AND U14443 ( .A(n14613), .B(n14614), .Z(n14612) );
  XNOR U14444 ( .A(p_input[2224]), .B(n14611), .Z(n14614) );
  XNOR U14445 ( .A(n14611), .B(n14283), .Z(n14613) );
  IV U14446 ( .A(p_input[2192]), .Z(n14283) );
  XOR U14447 ( .A(n14615), .B(n14616), .Z(n14611) );
  AND U14448 ( .A(n14617), .B(n14618), .Z(n14616) );
  XNOR U14449 ( .A(p_input[2223]), .B(n14615), .Z(n14618) );
  XNOR U14450 ( .A(n14615), .B(n14292), .Z(n14617) );
  IV U14451 ( .A(p_input[2191]), .Z(n14292) );
  XOR U14452 ( .A(n14619), .B(n14620), .Z(n14615) );
  AND U14453 ( .A(n14621), .B(n14622), .Z(n14620) );
  XNOR U14454 ( .A(p_input[2222]), .B(n14619), .Z(n14622) );
  XNOR U14455 ( .A(n14619), .B(n14301), .Z(n14621) );
  IV U14456 ( .A(p_input[2190]), .Z(n14301) );
  XOR U14457 ( .A(n14623), .B(n14624), .Z(n14619) );
  AND U14458 ( .A(n14625), .B(n14626), .Z(n14624) );
  XNOR U14459 ( .A(p_input[2221]), .B(n14623), .Z(n14626) );
  XNOR U14460 ( .A(n14623), .B(n14310), .Z(n14625) );
  IV U14461 ( .A(p_input[2189]), .Z(n14310) );
  XOR U14462 ( .A(n14627), .B(n14628), .Z(n14623) );
  AND U14463 ( .A(n14629), .B(n14630), .Z(n14628) );
  XNOR U14464 ( .A(p_input[2220]), .B(n14627), .Z(n14630) );
  XNOR U14465 ( .A(n14627), .B(n14319), .Z(n14629) );
  IV U14466 ( .A(p_input[2188]), .Z(n14319) );
  XOR U14467 ( .A(n14631), .B(n14632), .Z(n14627) );
  AND U14468 ( .A(n14633), .B(n14634), .Z(n14632) );
  XNOR U14469 ( .A(p_input[2219]), .B(n14631), .Z(n14634) );
  XNOR U14470 ( .A(n14631), .B(n14328), .Z(n14633) );
  IV U14471 ( .A(p_input[2187]), .Z(n14328) );
  XOR U14472 ( .A(n14635), .B(n14636), .Z(n14631) );
  AND U14473 ( .A(n14637), .B(n14638), .Z(n14636) );
  XNOR U14474 ( .A(p_input[2218]), .B(n14635), .Z(n14638) );
  XNOR U14475 ( .A(n14635), .B(n14337), .Z(n14637) );
  IV U14476 ( .A(p_input[2186]), .Z(n14337) );
  XOR U14477 ( .A(n14639), .B(n14640), .Z(n14635) );
  AND U14478 ( .A(n14641), .B(n14642), .Z(n14640) );
  XNOR U14479 ( .A(p_input[2217]), .B(n14639), .Z(n14642) );
  XNOR U14480 ( .A(n14639), .B(n14346), .Z(n14641) );
  IV U14481 ( .A(p_input[2185]), .Z(n14346) );
  XOR U14482 ( .A(n14643), .B(n14644), .Z(n14639) );
  AND U14483 ( .A(n14645), .B(n14646), .Z(n14644) );
  XNOR U14484 ( .A(p_input[2216]), .B(n14643), .Z(n14646) );
  XNOR U14485 ( .A(n14643), .B(n14355), .Z(n14645) );
  IV U14486 ( .A(p_input[2184]), .Z(n14355) );
  XOR U14487 ( .A(n14647), .B(n14648), .Z(n14643) );
  AND U14488 ( .A(n14649), .B(n14650), .Z(n14648) );
  XNOR U14489 ( .A(p_input[2215]), .B(n14647), .Z(n14650) );
  XNOR U14490 ( .A(n14647), .B(n14364), .Z(n14649) );
  IV U14491 ( .A(p_input[2183]), .Z(n14364) );
  XOR U14492 ( .A(n14651), .B(n14652), .Z(n14647) );
  AND U14493 ( .A(n14653), .B(n14654), .Z(n14652) );
  XNOR U14494 ( .A(p_input[2214]), .B(n14651), .Z(n14654) );
  XNOR U14495 ( .A(n14651), .B(n14373), .Z(n14653) );
  IV U14496 ( .A(p_input[2182]), .Z(n14373) );
  XOR U14497 ( .A(n14655), .B(n14656), .Z(n14651) );
  AND U14498 ( .A(n14657), .B(n14658), .Z(n14656) );
  XNOR U14499 ( .A(p_input[2213]), .B(n14655), .Z(n14658) );
  XNOR U14500 ( .A(n14655), .B(n14382), .Z(n14657) );
  IV U14501 ( .A(p_input[2181]), .Z(n14382) );
  XOR U14502 ( .A(n14659), .B(n14660), .Z(n14655) );
  AND U14503 ( .A(n14661), .B(n14662), .Z(n14660) );
  XNOR U14504 ( .A(p_input[2212]), .B(n14659), .Z(n14662) );
  XNOR U14505 ( .A(n14659), .B(n14391), .Z(n14661) );
  IV U14506 ( .A(p_input[2180]), .Z(n14391) );
  XOR U14507 ( .A(n14663), .B(n14664), .Z(n14659) );
  AND U14508 ( .A(n14665), .B(n14666), .Z(n14664) );
  XNOR U14509 ( .A(p_input[2211]), .B(n14663), .Z(n14666) );
  XNOR U14510 ( .A(n14663), .B(n14400), .Z(n14665) );
  IV U14511 ( .A(p_input[2179]), .Z(n14400) );
  XOR U14512 ( .A(n14667), .B(n14668), .Z(n14663) );
  AND U14513 ( .A(n14669), .B(n14670), .Z(n14668) );
  XNOR U14514 ( .A(p_input[2210]), .B(n14667), .Z(n14670) );
  XNOR U14515 ( .A(n14667), .B(n14409), .Z(n14669) );
  IV U14516 ( .A(p_input[2178]), .Z(n14409) );
  XNOR U14517 ( .A(n14671), .B(n14672), .Z(n14667) );
  AND U14518 ( .A(n14673), .B(n14674), .Z(n14672) );
  XOR U14519 ( .A(p_input[2209]), .B(n14671), .Z(n14674) );
  XNOR U14520 ( .A(p_input[2177]), .B(n14671), .Z(n14673) );
  AND U14521 ( .A(p_input[2208]), .B(n14675), .Z(n14671) );
  IV U14522 ( .A(p_input[2176]), .Z(n14675) );
  XOR U14523 ( .A(n14676), .B(n14677), .Z(n13765) );
  AND U14524 ( .A(n347), .B(n14678), .Z(n14677) );
  XNOR U14525 ( .A(n14679), .B(n14676), .Z(n14678) );
  XOR U14526 ( .A(n14680), .B(n14681), .Z(n347) );
  AND U14527 ( .A(n14682), .B(n14683), .Z(n14681) );
  XNOR U14528 ( .A(n13780), .B(n14680), .Z(n14683) );
  AND U14529 ( .A(p_input[2175]), .B(p_input[2143]), .Z(n13780) );
  XNOR U14530 ( .A(n14680), .B(n13777), .Z(n14682) );
  IV U14531 ( .A(n14684), .Z(n13777) );
  AND U14532 ( .A(p_input[2079]), .B(p_input[2111]), .Z(n14684) );
  XOR U14533 ( .A(n14685), .B(n14686), .Z(n14680) );
  AND U14534 ( .A(n14687), .B(n14688), .Z(n14686) );
  XOR U14535 ( .A(n14685), .B(n13792), .Z(n14688) );
  XNOR U14536 ( .A(p_input[2142]), .B(n14689), .Z(n13792) );
  AND U14537 ( .A(n286), .B(n14690), .Z(n14689) );
  XOR U14538 ( .A(p_input[2174]), .B(p_input[2142]), .Z(n14690) );
  XNOR U14539 ( .A(n13789), .B(n14685), .Z(n14687) );
  XOR U14540 ( .A(n14691), .B(n14692), .Z(n13789) );
  AND U14541 ( .A(n283), .B(n14693), .Z(n14692) );
  XOR U14542 ( .A(p_input[2110]), .B(p_input[2078]), .Z(n14693) );
  XOR U14543 ( .A(n14694), .B(n14695), .Z(n14685) );
  AND U14544 ( .A(n14696), .B(n14697), .Z(n14695) );
  XOR U14545 ( .A(n14694), .B(n13804), .Z(n14697) );
  XNOR U14546 ( .A(p_input[2141]), .B(n14698), .Z(n13804) );
  AND U14547 ( .A(n286), .B(n14699), .Z(n14698) );
  XOR U14548 ( .A(p_input[2173]), .B(p_input[2141]), .Z(n14699) );
  XNOR U14549 ( .A(n13801), .B(n14694), .Z(n14696) );
  XOR U14550 ( .A(n14700), .B(n14701), .Z(n13801) );
  AND U14551 ( .A(n283), .B(n14702), .Z(n14701) );
  XOR U14552 ( .A(p_input[2109]), .B(p_input[2077]), .Z(n14702) );
  XOR U14553 ( .A(n14703), .B(n14704), .Z(n14694) );
  AND U14554 ( .A(n14705), .B(n14706), .Z(n14704) );
  XOR U14555 ( .A(n14703), .B(n13816), .Z(n14706) );
  XNOR U14556 ( .A(p_input[2140]), .B(n14707), .Z(n13816) );
  AND U14557 ( .A(n286), .B(n14708), .Z(n14707) );
  XOR U14558 ( .A(p_input[2172]), .B(p_input[2140]), .Z(n14708) );
  XNOR U14559 ( .A(n13813), .B(n14703), .Z(n14705) );
  XOR U14560 ( .A(n14709), .B(n14710), .Z(n13813) );
  AND U14561 ( .A(n283), .B(n14711), .Z(n14710) );
  XOR U14562 ( .A(p_input[2108]), .B(p_input[2076]), .Z(n14711) );
  XOR U14563 ( .A(n14712), .B(n14713), .Z(n14703) );
  AND U14564 ( .A(n14714), .B(n14715), .Z(n14713) );
  XOR U14565 ( .A(n14712), .B(n13828), .Z(n14715) );
  XNOR U14566 ( .A(p_input[2139]), .B(n14716), .Z(n13828) );
  AND U14567 ( .A(n286), .B(n14717), .Z(n14716) );
  XOR U14568 ( .A(p_input[2171]), .B(p_input[2139]), .Z(n14717) );
  XNOR U14569 ( .A(n13825), .B(n14712), .Z(n14714) );
  XOR U14570 ( .A(n14718), .B(n14719), .Z(n13825) );
  AND U14571 ( .A(n283), .B(n14720), .Z(n14719) );
  XOR U14572 ( .A(p_input[2107]), .B(p_input[2075]), .Z(n14720) );
  XOR U14573 ( .A(n14721), .B(n14722), .Z(n14712) );
  AND U14574 ( .A(n14723), .B(n14724), .Z(n14722) );
  XOR U14575 ( .A(n14721), .B(n13840), .Z(n14724) );
  XNOR U14576 ( .A(p_input[2138]), .B(n14725), .Z(n13840) );
  AND U14577 ( .A(n286), .B(n14726), .Z(n14725) );
  XOR U14578 ( .A(p_input[2170]), .B(p_input[2138]), .Z(n14726) );
  XNOR U14579 ( .A(n13837), .B(n14721), .Z(n14723) );
  XOR U14580 ( .A(n14727), .B(n14728), .Z(n13837) );
  AND U14581 ( .A(n283), .B(n14729), .Z(n14728) );
  XOR U14582 ( .A(p_input[2106]), .B(p_input[2074]), .Z(n14729) );
  XOR U14583 ( .A(n14730), .B(n14731), .Z(n14721) );
  AND U14584 ( .A(n14732), .B(n14733), .Z(n14731) );
  XOR U14585 ( .A(n14730), .B(n13852), .Z(n14733) );
  XNOR U14586 ( .A(p_input[2137]), .B(n14734), .Z(n13852) );
  AND U14587 ( .A(n286), .B(n14735), .Z(n14734) );
  XOR U14588 ( .A(p_input[2169]), .B(p_input[2137]), .Z(n14735) );
  XNOR U14589 ( .A(n13849), .B(n14730), .Z(n14732) );
  XOR U14590 ( .A(n14736), .B(n14737), .Z(n13849) );
  AND U14591 ( .A(n283), .B(n14738), .Z(n14737) );
  XOR U14592 ( .A(p_input[2105]), .B(p_input[2073]), .Z(n14738) );
  XOR U14593 ( .A(n14739), .B(n14740), .Z(n14730) );
  AND U14594 ( .A(n14741), .B(n14742), .Z(n14740) );
  XOR U14595 ( .A(n14739), .B(n13864), .Z(n14742) );
  XNOR U14596 ( .A(p_input[2136]), .B(n14743), .Z(n13864) );
  AND U14597 ( .A(n286), .B(n14744), .Z(n14743) );
  XOR U14598 ( .A(p_input[2168]), .B(p_input[2136]), .Z(n14744) );
  XNOR U14599 ( .A(n13861), .B(n14739), .Z(n14741) );
  XOR U14600 ( .A(n14745), .B(n14746), .Z(n13861) );
  AND U14601 ( .A(n283), .B(n14747), .Z(n14746) );
  XOR U14602 ( .A(p_input[2104]), .B(p_input[2072]), .Z(n14747) );
  XOR U14603 ( .A(n14748), .B(n14749), .Z(n14739) );
  AND U14604 ( .A(n14750), .B(n14751), .Z(n14749) );
  XOR U14605 ( .A(n14748), .B(n13876), .Z(n14751) );
  XNOR U14606 ( .A(p_input[2135]), .B(n14752), .Z(n13876) );
  AND U14607 ( .A(n286), .B(n14753), .Z(n14752) );
  XOR U14608 ( .A(p_input[2167]), .B(p_input[2135]), .Z(n14753) );
  XNOR U14609 ( .A(n13873), .B(n14748), .Z(n14750) );
  XOR U14610 ( .A(n14754), .B(n14755), .Z(n13873) );
  AND U14611 ( .A(n283), .B(n14756), .Z(n14755) );
  XOR U14612 ( .A(p_input[2103]), .B(p_input[2071]), .Z(n14756) );
  XOR U14613 ( .A(n14757), .B(n14758), .Z(n14748) );
  AND U14614 ( .A(n14759), .B(n14760), .Z(n14758) );
  XOR U14615 ( .A(n14757), .B(n13888), .Z(n14760) );
  XNOR U14616 ( .A(p_input[2134]), .B(n14761), .Z(n13888) );
  AND U14617 ( .A(n286), .B(n14762), .Z(n14761) );
  XOR U14618 ( .A(p_input[2166]), .B(p_input[2134]), .Z(n14762) );
  XNOR U14619 ( .A(n13885), .B(n14757), .Z(n14759) );
  XOR U14620 ( .A(n14763), .B(n14764), .Z(n13885) );
  AND U14621 ( .A(n283), .B(n14765), .Z(n14764) );
  XOR U14622 ( .A(p_input[2102]), .B(p_input[2070]), .Z(n14765) );
  XOR U14623 ( .A(n14766), .B(n14767), .Z(n14757) );
  AND U14624 ( .A(n14768), .B(n14769), .Z(n14767) );
  XOR U14625 ( .A(n14766), .B(n13900), .Z(n14769) );
  XNOR U14626 ( .A(p_input[2133]), .B(n14770), .Z(n13900) );
  AND U14627 ( .A(n286), .B(n14771), .Z(n14770) );
  XOR U14628 ( .A(p_input[2165]), .B(p_input[2133]), .Z(n14771) );
  XNOR U14629 ( .A(n13897), .B(n14766), .Z(n14768) );
  XOR U14630 ( .A(n14772), .B(n14773), .Z(n13897) );
  AND U14631 ( .A(n283), .B(n14774), .Z(n14773) );
  XOR U14632 ( .A(p_input[2101]), .B(p_input[2069]), .Z(n14774) );
  XOR U14633 ( .A(n14775), .B(n14776), .Z(n14766) );
  AND U14634 ( .A(n14777), .B(n14778), .Z(n14776) );
  XOR U14635 ( .A(n14775), .B(n13912), .Z(n14778) );
  XNOR U14636 ( .A(p_input[2132]), .B(n14779), .Z(n13912) );
  AND U14637 ( .A(n286), .B(n14780), .Z(n14779) );
  XOR U14638 ( .A(p_input[2164]), .B(p_input[2132]), .Z(n14780) );
  XNOR U14639 ( .A(n13909), .B(n14775), .Z(n14777) );
  XOR U14640 ( .A(n14781), .B(n14782), .Z(n13909) );
  AND U14641 ( .A(n283), .B(n14783), .Z(n14782) );
  XOR U14642 ( .A(p_input[2100]), .B(p_input[2068]), .Z(n14783) );
  XOR U14643 ( .A(n14784), .B(n14785), .Z(n14775) );
  AND U14644 ( .A(n14786), .B(n14787), .Z(n14785) );
  XOR U14645 ( .A(n14784), .B(n13924), .Z(n14787) );
  XNOR U14646 ( .A(p_input[2131]), .B(n14788), .Z(n13924) );
  AND U14647 ( .A(n286), .B(n14789), .Z(n14788) );
  XOR U14648 ( .A(p_input[2163]), .B(p_input[2131]), .Z(n14789) );
  XNOR U14649 ( .A(n13921), .B(n14784), .Z(n14786) );
  XOR U14650 ( .A(n14790), .B(n14791), .Z(n13921) );
  AND U14651 ( .A(n283), .B(n14792), .Z(n14791) );
  XOR U14652 ( .A(p_input[2099]), .B(p_input[2067]), .Z(n14792) );
  XOR U14653 ( .A(n14793), .B(n14794), .Z(n14784) );
  AND U14654 ( .A(n14795), .B(n14796), .Z(n14794) );
  XOR U14655 ( .A(n14793), .B(n13936), .Z(n14796) );
  XNOR U14656 ( .A(p_input[2130]), .B(n14797), .Z(n13936) );
  AND U14657 ( .A(n286), .B(n14798), .Z(n14797) );
  XOR U14658 ( .A(p_input[2162]), .B(p_input[2130]), .Z(n14798) );
  XNOR U14659 ( .A(n13933), .B(n14793), .Z(n14795) );
  XOR U14660 ( .A(n14799), .B(n14800), .Z(n13933) );
  AND U14661 ( .A(n283), .B(n14801), .Z(n14800) );
  XOR U14662 ( .A(p_input[2098]), .B(p_input[2066]), .Z(n14801) );
  XOR U14663 ( .A(n14802), .B(n14803), .Z(n14793) );
  AND U14664 ( .A(n14804), .B(n14805), .Z(n14803) );
  XOR U14665 ( .A(n14802), .B(n13948), .Z(n14805) );
  XNOR U14666 ( .A(p_input[2129]), .B(n14806), .Z(n13948) );
  AND U14667 ( .A(n286), .B(n14807), .Z(n14806) );
  XOR U14668 ( .A(p_input[2161]), .B(p_input[2129]), .Z(n14807) );
  XNOR U14669 ( .A(n13945), .B(n14802), .Z(n14804) );
  XOR U14670 ( .A(n14808), .B(n14809), .Z(n13945) );
  AND U14671 ( .A(n283), .B(n14810), .Z(n14809) );
  XOR U14672 ( .A(p_input[2097]), .B(p_input[2065]), .Z(n14810) );
  XOR U14673 ( .A(n14811), .B(n14812), .Z(n14802) );
  AND U14674 ( .A(n14813), .B(n14814), .Z(n14812) );
  XOR U14675 ( .A(n14811), .B(n13960), .Z(n14814) );
  XNOR U14676 ( .A(p_input[2128]), .B(n14815), .Z(n13960) );
  AND U14677 ( .A(n286), .B(n14816), .Z(n14815) );
  XOR U14678 ( .A(p_input[2160]), .B(p_input[2128]), .Z(n14816) );
  XNOR U14679 ( .A(n13957), .B(n14811), .Z(n14813) );
  XOR U14680 ( .A(n14817), .B(n14818), .Z(n13957) );
  AND U14681 ( .A(n283), .B(n14819), .Z(n14818) );
  XOR U14682 ( .A(p_input[2096]), .B(p_input[2064]), .Z(n14819) );
  XOR U14683 ( .A(n14820), .B(n14821), .Z(n14811) );
  AND U14684 ( .A(n14822), .B(n14823), .Z(n14821) );
  XOR U14685 ( .A(n14820), .B(n13972), .Z(n14823) );
  XNOR U14686 ( .A(p_input[2127]), .B(n14824), .Z(n13972) );
  AND U14687 ( .A(n286), .B(n14825), .Z(n14824) );
  XOR U14688 ( .A(p_input[2159]), .B(p_input[2127]), .Z(n14825) );
  XNOR U14689 ( .A(n13969), .B(n14820), .Z(n14822) );
  XOR U14690 ( .A(n14826), .B(n14827), .Z(n13969) );
  AND U14691 ( .A(n283), .B(n14828), .Z(n14827) );
  XOR U14692 ( .A(p_input[2095]), .B(p_input[2063]), .Z(n14828) );
  XOR U14693 ( .A(n14829), .B(n14830), .Z(n14820) );
  AND U14694 ( .A(n14831), .B(n14832), .Z(n14830) );
  XOR U14695 ( .A(n14829), .B(n13984), .Z(n14832) );
  XNOR U14696 ( .A(p_input[2126]), .B(n14833), .Z(n13984) );
  AND U14697 ( .A(n286), .B(n14834), .Z(n14833) );
  XOR U14698 ( .A(p_input[2158]), .B(p_input[2126]), .Z(n14834) );
  XNOR U14699 ( .A(n13981), .B(n14829), .Z(n14831) );
  XOR U14700 ( .A(n14835), .B(n14836), .Z(n13981) );
  AND U14701 ( .A(n283), .B(n14837), .Z(n14836) );
  XOR U14702 ( .A(p_input[2094]), .B(p_input[2062]), .Z(n14837) );
  XOR U14703 ( .A(n14838), .B(n14839), .Z(n14829) );
  AND U14704 ( .A(n14840), .B(n14841), .Z(n14839) );
  XOR U14705 ( .A(n14838), .B(n13996), .Z(n14841) );
  XNOR U14706 ( .A(p_input[2125]), .B(n14842), .Z(n13996) );
  AND U14707 ( .A(n286), .B(n14843), .Z(n14842) );
  XOR U14708 ( .A(p_input[2157]), .B(p_input[2125]), .Z(n14843) );
  XNOR U14709 ( .A(n13993), .B(n14838), .Z(n14840) );
  XOR U14710 ( .A(n14844), .B(n14845), .Z(n13993) );
  AND U14711 ( .A(n283), .B(n14846), .Z(n14845) );
  XOR U14712 ( .A(p_input[2093]), .B(p_input[2061]), .Z(n14846) );
  XOR U14713 ( .A(n14847), .B(n14848), .Z(n14838) );
  AND U14714 ( .A(n14849), .B(n14850), .Z(n14848) );
  XOR U14715 ( .A(n14847), .B(n14008), .Z(n14850) );
  XNOR U14716 ( .A(p_input[2124]), .B(n14851), .Z(n14008) );
  AND U14717 ( .A(n286), .B(n14852), .Z(n14851) );
  XOR U14718 ( .A(p_input[2156]), .B(p_input[2124]), .Z(n14852) );
  XNOR U14719 ( .A(n14005), .B(n14847), .Z(n14849) );
  XOR U14720 ( .A(n14853), .B(n14854), .Z(n14005) );
  AND U14721 ( .A(n283), .B(n14855), .Z(n14854) );
  XOR U14722 ( .A(p_input[2092]), .B(p_input[2060]), .Z(n14855) );
  XOR U14723 ( .A(n14856), .B(n14857), .Z(n14847) );
  AND U14724 ( .A(n14858), .B(n14859), .Z(n14857) );
  XOR U14725 ( .A(n14856), .B(n14020), .Z(n14859) );
  XNOR U14726 ( .A(p_input[2123]), .B(n14860), .Z(n14020) );
  AND U14727 ( .A(n286), .B(n14861), .Z(n14860) );
  XOR U14728 ( .A(p_input[2155]), .B(p_input[2123]), .Z(n14861) );
  XNOR U14729 ( .A(n14017), .B(n14856), .Z(n14858) );
  XOR U14730 ( .A(n14862), .B(n14863), .Z(n14017) );
  AND U14731 ( .A(n283), .B(n14864), .Z(n14863) );
  XOR U14732 ( .A(p_input[2091]), .B(p_input[2059]), .Z(n14864) );
  XOR U14733 ( .A(n14865), .B(n14866), .Z(n14856) );
  AND U14734 ( .A(n14867), .B(n14868), .Z(n14866) );
  XOR U14735 ( .A(n14865), .B(n14032), .Z(n14868) );
  XNOR U14736 ( .A(p_input[2122]), .B(n14869), .Z(n14032) );
  AND U14737 ( .A(n286), .B(n14870), .Z(n14869) );
  XOR U14738 ( .A(p_input[2154]), .B(p_input[2122]), .Z(n14870) );
  XNOR U14739 ( .A(n14029), .B(n14865), .Z(n14867) );
  XOR U14740 ( .A(n14871), .B(n14872), .Z(n14029) );
  AND U14741 ( .A(n283), .B(n14873), .Z(n14872) );
  XOR U14742 ( .A(p_input[2090]), .B(p_input[2058]), .Z(n14873) );
  XOR U14743 ( .A(n14874), .B(n14875), .Z(n14865) );
  AND U14744 ( .A(n14876), .B(n14877), .Z(n14875) );
  XOR U14745 ( .A(n14874), .B(n14044), .Z(n14877) );
  XNOR U14746 ( .A(p_input[2121]), .B(n14878), .Z(n14044) );
  AND U14747 ( .A(n286), .B(n14879), .Z(n14878) );
  XOR U14748 ( .A(p_input[2153]), .B(p_input[2121]), .Z(n14879) );
  XNOR U14749 ( .A(n14041), .B(n14874), .Z(n14876) );
  XOR U14750 ( .A(n14880), .B(n14881), .Z(n14041) );
  AND U14751 ( .A(n283), .B(n14882), .Z(n14881) );
  XOR U14752 ( .A(p_input[2089]), .B(p_input[2057]), .Z(n14882) );
  XOR U14753 ( .A(n14883), .B(n14884), .Z(n14874) );
  AND U14754 ( .A(n14885), .B(n14886), .Z(n14884) );
  XOR U14755 ( .A(n14883), .B(n14056), .Z(n14886) );
  XNOR U14756 ( .A(p_input[2120]), .B(n14887), .Z(n14056) );
  AND U14757 ( .A(n286), .B(n14888), .Z(n14887) );
  XOR U14758 ( .A(p_input[2152]), .B(p_input[2120]), .Z(n14888) );
  XNOR U14759 ( .A(n14053), .B(n14883), .Z(n14885) );
  XOR U14760 ( .A(n14889), .B(n14890), .Z(n14053) );
  AND U14761 ( .A(n283), .B(n14891), .Z(n14890) );
  XOR U14762 ( .A(p_input[2088]), .B(p_input[2056]), .Z(n14891) );
  XOR U14763 ( .A(n14892), .B(n14893), .Z(n14883) );
  AND U14764 ( .A(n14894), .B(n14895), .Z(n14893) );
  XOR U14765 ( .A(n14892), .B(n14068), .Z(n14895) );
  XNOR U14766 ( .A(p_input[2119]), .B(n14896), .Z(n14068) );
  AND U14767 ( .A(n286), .B(n14897), .Z(n14896) );
  XOR U14768 ( .A(p_input[2151]), .B(p_input[2119]), .Z(n14897) );
  XNOR U14769 ( .A(n14065), .B(n14892), .Z(n14894) );
  XOR U14770 ( .A(n14898), .B(n14899), .Z(n14065) );
  AND U14771 ( .A(n283), .B(n14900), .Z(n14899) );
  XOR U14772 ( .A(p_input[2087]), .B(p_input[2055]), .Z(n14900) );
  XOR U14773 ( .A(n14901), .B(n14902), .Z(n14892) );
  AND U14774 ( .A(n14903), .B(n14904), .Z(n14902) );
  XOR U14775 ( .A(n14901), .B(n14080), .Z(n14904) );
  XNOR U14776 ( .A(p_input[2118]), .B(n14905), .Z(n14080) );
  AND U14777 ( .A(n286), .B(n14906), .Z(n14905) );
  XOR U14778 ( .A(p_input[2150]), .B(p_input[2118]), .Z(n14906) );
  XNOR U14779 ( .A(n14077), .B(n14901), .Z(n14903) );
  XOR U14780 ( .A(n14907), .B(n14908), .Z(n14077) );
  AND U14781 ( .A(n283), .B(n14909), .Z(n14908) );
  XOR U14782 ( .A(p_input[2086]), .B(p_input[2054]), .Z(n14909) );
  XOR U14783 ( .A(n14910), .B(n14911), .Z(n14901) );
  AND U14784 ( .A(n14912), .B(n14913), .Z(n14911) );
  XOR U14785 ( .A(n14910), .B(n14092), .Z(n14913) );
  XNOR U14786 ( .A(p_input[2117]), .B(n14914), .Z(n14092) );
  AND U14787 ( .A(n286), .B(n14915), .Z(n14914) );
  XOR U14788 ( .A(p_input[2149]), .B(p_input[2117]), .Z(n14915) );
  XNOR U14789 ( .A(n14089), .B(n14910), .Z(n14912) );
  XOR U14790 ( .A(n14916), .B(n14917), .Z(n14089) );
  AND U14791 ( .A(n283), .B(n14918), .Z(n14917) );
  XOR U14792 ( .A(p_input[2085]), .B(p_input[2053]), .Z(n14918) );
  XOR U14793 ( .A(n14919), .B(n14920), .Z(n14910) );
  AND U14794 ( .A(n14921), .B(n14922), .Z(n14920) );
  XOR U14795 ( .A(n14919), .B(n14104), .Z(n14922) );
  XNOR U14796 ( .A(p_input[2116]), .B(n14923), .Z(n14104) );
  AND U14797 ( .A(n286), .B(n14924), .Z(n14923) );
  XOR U14798 ( .A(p_input[2148]), .B(p_input[2116]), .Z(n14924) );
  XNOR U14799 ( .A(n14101), .B(n14919), .Z(n14921) );
  XOR U14800 ( .A(n14925), .B(n14926), .Z(n14101) );
  AND U14801 ( .A(n283), .B(n14927), .Z(n14926) );
  XOR U14802 ( .A(p_input[2084]), .B(p_input[2052]), .Z(n14927) );
  XOR U14803 ( .A(n14928), .B(n14929), .Z(n14919) );
  AND U14804 ( .A(n14930), .B(n14931), .Z(n14929) );
  XOR U14805 ( .A(n14928), .B(n14116), .Z(n14931) );
  XNOR U14806 ( .A(p_input[2115]), .B(n14932), .Z(n14116) );
  AND U14807 ( .A(n286), .B(n14933), .Z(n14932) );
  XOR U14808 ( .A(p_input[2147]), .B(p_input[2115]), .Z(n14933) );
  XNOR U14809 ( .A(n14113), .B(n14928), .Z(n14930) );
  XOR U14810 ( .A(n14934), .B(n14935), .Z(n14113) );
  AND U14811 ( .A(n283), .B(n14936), .Z(n14935) );
  XOR U14812 ( .A(p_input[2083]), .B(p_input[2051]), .Z(n14936) );
  XOR U14813 ( .A(n14937), .B(n14938), .Z(n14928) );
  AND U14814 ( .A(n14939), .B(n14940), .Z(n14938) );
  XOR U14815 ( .A(n14128), .B(n14937), .Z(n14940) );
  XNOR U14816 ( .A(p_input[2114]), .B(n14941), .Z(n14128) );
  AND U14817 ( .A(n286), .B(n14942), .Z(n14941) );
  XOR U14818 ( .A(p_input[2146]), .B(p_input[2114]), .Z(n14942) );
  XNOR U14819 ( .A(n14937), .B(n14125), .Z(n14939) );
  XOR U14820 ( .A(n14943), .B(n14944), .Z(n14125) );
  AND U14821 ( .A(n283), .B(n14945), .Z(n14944) );
  XOR U14822 ( .A(p_input[2082]), .B(p_input[2050]), .Z(n14945) );
  XOR U14823 ( .A(n14946), .B(n14947), .Z(n14937) );
  AND U14824 ( .A(n14948), .B(n14949), .Z(n14947) );
  XNOR U14825 ( .A(n14950), .B(n14141), .Z(n14949) );
  XNOR U14826 ( .A(p_input[2113]), .B(n14951), .Z(n14141) );
  AND U14827 ( .A(n286), .B(n14952), .Z(n14951) );
  XNOR U14828 ( .A(p_input[2145]), .B(n14953), .Z(n14952) );
  IV U14829 ( .A(p_input[2113]), .Z(n14953) );
  XNOR U14830 ( .A(n14138), .B(n14946), .Z(n14948) );
  XNOR U14831 ( .A(p_input[2049]), .B(n14954), .Z(n14138) );
  AND U14832 ( .A(n283), .B(n14955), .Z(n14954) );
  XOR U14833 ( .A(p_input[2081]), .B(p_input[2049]), .Z(n14955) );
  IV U14834 ( .A(n14950), .Z(n14946) );
  AND U14835 ( .A(n14676), .B(n14679), .Z(n14950) );
  XOR U14836 ( .A(p_input[2112]), .B(n14956), .Z(n14679) );
  AND U14837 ( .A(n286), .B(n14957), .Z(n14956) );
  XOR U14838 ( .A(p_input[2144]), .B(p_input[2112]), .Z(n14957) );
  XOR U14839 ( .A(n14958), .B(n14959), .Z(n286) );
  AND U14840 ( .A(n14960), .B(n14961), .Z(n14959) );
  XNOR U14841 ( .A(p_input[2175]), .B(n14958), .Z(n14961) );
  XOR U14842 ( .A(n14958), .B(p_input[2143]), .Z(n14960) );
  XOR U14843 ( .A(n14962), .B(n14963), .Z(n14958) );
  AND U14844 ( .A(n14964), .B(n14965), .Z(n14963) );
  XNOR U14845 ( .A(p_input[2174]), .B(n14962), .Z(n14965) );
  XOR U14846 ( .A(n14962), .B(p_input[2142]), .Z(n14964) );
  XOR U14847 ( .A(n14966), .B(n14967), .Z(n14962) );
  AND U14848 ( .A(n14968), .B(n14969), .Z(n14967) );
  XNOR U14849 ( .A(p_input[2173]), .B(n14966), .Z(n14969) );
  XOR U14850 ( .A(n14966), .B(p_input[2141]), .Z(n14968) );
  XOR U14851 ( .A(n14970), .B(n14971), .Z(n14966) );
  AND U14852 ( .A(n14972), .B(n14973), .Z(n14971) );
  XNOR U14853 ( .A(p_input[2172]), .B(n14970), .Z(n14973) );
  XOR U14854 ( .A(n14970), .B(p_input[2140]), .Z(n14972) );
  XOR U14855 ( .A(n14974), .B(n14975), .Z(n14970) );
  AND U14856 ( .A(n14976), .B(n14977), .Z(n14975) );
  XNOR U14857 ( .A(p_input[2171]), .B(n14974), .Z(n14977) );
  XOR U14858 ( .A(n14974), .B(p_input[2139]), .Z(n14976) );
  XOR U14859 ( .A(n14978), .B(n14979), .Z(n14974) );
  AND U14860 ( .A(n14980), .B(n14981), .Z(n14979) );
  XNOR U14861 ( .A(p_input[2170]), .B(n14978), .Z(n14981) );
  XOR U14862 ( .A(n14978), .B(p_input[2138]), .Z(n14980) );
  XOR U14863 ( .A(n14982), .B(n14983), .Z(n14978) );
  AND U14864 ( .A(n14984), .B(n14985), .Z(n14983) );
  XNOR U14865 ( .A(p_input[2169]), .B(n14982), .Z(n14985) );
  XOR U14866 ( .A(n14982), .B(p_input[2137]), .Z(n14984) );
  XOR U14867 ( .A(n14986), .B(n14987), .Z(n14982) );
  AND U14868 ( .A(n14988), .B(n14989), .Z(n14987) );
  XNOR U14869 ( .A(p_input[2168]), .B(n14986), .Z(n14989) );
  XOR U14870 ( .A(n14986), .B(p_input[2136]), .Z(n14988) );
  XOR U14871 ( .A(n14990), .B(n14991), .Z(n14986) );
  AND U14872 ( .A(n14992), .B(n14993), .Z(n14991) );
  XNOR U14873 ( .A(p_input[2167]), .B(n14990), .Z(n14993) );
  XOR U14874 ( .A(n14990), .B(p_input[2135]), .Z(n14992) );
  XOR U14875 ( .A(n14994), .B(n14995), .Z(n14990) );
  AND U14876 ( .A(n14996), .B(n14997), .Z(n14995) );
  XNOR U14877 ( .A(p_input[2166]), .B(n14994), .Z(n14997) );
  XOR U14878 ( .A(n14994), .B(p_input[2134]), .Z(n14996) );
  XOR U14879 ( .A(n14998), .B(n14999), .Z(n14994) );
  AND U14880 ( .A(n15000), .B(n15001), .Z(n14999) );
  XNOR U14881 ( .A(p_input[2165]), .B(n14998), .Z(n15001) );
  XOR U14882 ( .A(n14998), .B(p_input[2133]), .Z(n15000) );
  XOR U14883 ( .A(n15002), .B(n15003), .Z(n14998) );
  AND U14884 ( .A(n15004), .B(n15005), .Z(n15003) );
  XNOR U14885 ( .A(p_input[2164]), .B(n15002), .Z(n15005) );
  XOR U14886 ( .A(n15002), .B(p_input[2132]), .Z(n15004) );
  XOR U14887 ( .A(n15006), .B(n15007), .Z(n15002) );
  AND U14888 ( .A(n15008), .B(n15009), .Z(n15007) );
  XNOR U14889 ( .A(p_input[2163]), .B(n15006), .Z(n15009) );
  XOR U14890 ( .A(n15006), .B(p_input[2131]), .Z(n15008) );
  XOR U14891 ( .A(n15010), .B(n15011), .Z(n15006) );
  AND U14892 ( .A(n15012), .B(n15013), .Z(n15011) );
  XNOR U14893 ( .A(p_input[2162]), .B(n15010), .Z(n15013) );
  XOR U14894 ( .A(n15010), .B(p_input[2130]), .Z(n15012) );
  XOR U14895 ( .A(n15014), .B(n15015), .Z(n15010) );
  AND U14896 ( .A(n15016), .B(n15017), .Z(n15015) );
  XNOR U14897 ( .A(p_input[2161]), .B(n15014), .Z(n15017) );
  XOR U14898 ( .A(n15014), .B(p_input[2129]), .Z(n15016) );
  XOR U14899 ( .A(n15018), .B(n15019), .Z(n15014) );
  AND U14900 ( .A(n15020), .B(n15021), .Z(n15019) );
  XNOR U14901 ( .A(p_input[2160]), .B(n15018), .Z(n15021) );
  XOR U14902 ( .A(n15018), .B(p_input[2128]), .Z(n15020) );
  XOR U14903 ( .A(n15022), .B(n15023), .Z(n15018) );
  AND U14904 ( .A(n15024), .B(n15025), .Z(n15023) );
  XNOR U14905 ( .A(p_input[2159]), .B(n15022), .Z(n15025) );
  XOR U14906 ( .A(n15022), .B(p_input[2127]), .Z(n15024) );
  XOR U14907 ( .A(n15026), .B(n15027), .Z(n15022) );
  AND U14908 ( .A(n15028), .B(n15029), .Z(n15027) );
  XNOR U14909 ( .A(p_input[2158]), .B(n15026), .Z(n15029) );
  XOR U14910 ( .A(n15026), .B(p_input[2126]), .Z(n15028) );
  XOR U14911 ( .A(n15030), .B(n15031), .Z(n15026) );
  AND U14912 ( .A(n15032), .B(n15033), .Z(n15031) );
  XNOR U14913 ( .A(p_input[2157]), .B(n15030), .Z(n15033) );
  XOR U14914 ( .A(n15030), .B(p_input[2125]), .Z(n15032) );
  XOR U14915 ( .A(n15034), .B(n15035), .Z(n15030) );
  AND U14916 ( .A(n15036), .B(n15037), .Z(n15035) );
  XNOR U14917 ( .A(p_input[2156]), .B(n15034), .Z(n15037) );
  XOR U14918 ( .A(n15034), .B(p_input[2124]), .Z(n15036) );
  XOR U14919 ( .A(n15038), .B(n15039), .Z(n15034) );
  AND U14920 ( .A(n15040), .B(n15041), .Z(n15039) );
  XNOR U14921 ( .A(p_input[2155]), .B(n15038), .Z(n15041) );
  XOR U14922 ( .A(n15038), .B(p_input[2123]), .Z(n15040) );
  XOR U14923 ( .A(n15042), .B(n15043), .Z(n15038) );
  AND U14924 ( .A(n15044), .B(n15045), .Z(n15043) );
  XNOR U14925 ( .A(p_input[2154]), .B(n15042), .Z(n15045) );
  XOR U14926 ( .A(n15042), .B(p_input[2122]), .Z(n15044) );
  XOR U14927 ( .A(n15046), .B(n15047), .Z(n15042) );
  AND U14928 ( .A(n15048), .B(n15049), .Z(n15047) );
  XNOR U14929 ( .A(p_input[2153]), .B(n15046), .Z(n15049) );
  XOR U14930 ( .A(n15046), .B(p_input[2121]), .Z(n15048) );
  XOR U14931 ( .A(n15050), .B(n15051), .Z(n15046) );
  AND U14932 ( .A(n15052), .B(n15053), .Z(n15051) );
  XNOR U14933 ( .A(p_input[2152]), .B(n15050), .Z(n15053) );
  XOR U14934 ( .A(n15050), .B(p_input[2120]), .Z(n15052) );
  XOR U14935 ( .A(n15054), .B(n15055), .Z(n15050) );
  AND U14936 ( .A(n15056), .B(n15057), .Z(n15055) );
  XNOR U14937 ( .A(p_input[2151]), .B(n15054), .Z(n15057) );
  XOR U14938 ( .A(n15054), .B(p_input[2119]), .Z(n15056) );
  XOR U14939 ( .A(n15058), .B(n15059), .Z(n15054) );
  AND U14940 ( .A(n15060), .B(n15061), .Z(n15059) );
  XNOR U14941 ( .A(p_input[2150]), .B(n15058), .Z(n15061) );
  XOR U14942 ( .A(n15058), .B(p_input[2118]), .Z(n15060) );
  XOR U14943 ( .A(n15062), .B(n15063), .Z(n15058) );
  AND U14944 ( .A(n15064), .B(n15065), .Z(n15063) );
  XNOR U14945 ( .A(p_input[2149]), .B(n15062), .Z(n15065) );
  XOR U14946 ( .A(n15062), .B(p_input[2117]), .Z(n15064) );
  XOR U14947 ( .A(n15066), .B(n15067), .Z(n15062) );
  AND U14948 ( .A(n15068), .B(n15069), .Z(n15067) );
  XNOR U14949 ( .A(p_input[2148]), .B(n15066), .Z(n15069) );
  XOR U14950 ( .A(n15066), .B(p_input[2116]), .Z(n15068) );
  XOR U14951 ( .A(n15070), .B(n15071), .Z(n15066) );
  AND U14952 ( .A(n15072), .B(n15073), .Z(n15071) );
  XNOR U14953 ( .A(p_input[2147]), .B(n15070), .Z(n15073) );
  XOR U14954 ( .A(n15070), .B(p_input[2115]), .Z(n15072) );
  XOR U14955 ( .A(n15074), .B(n15075), .Z(n15070) );
  AND U14956 ( .A(n15076), .B(n15077), .Z(n15075) );
  XNOR U14957 ( .A(p_input[2146]), .B(n15074), .Z(n15077) );
  XOR U14958 ( .A(n15074), .B(p_input[2114]), .Z(n15076) );
  XNOR U14959 ( .A(n15078), .B(n15079), .Z(n15074) );
  AND U14960 ( .A(n15080), .B(n15081), .Z(n15079) );
  XOR U14961 ( .A(p_input[2145]), .B(n15078), .Z(n15081) );
  XNOR U14962 ( .A(p_input[2113]), .B(n15078), .Z(n15080) );
  AND U14963 ( .A(p_input[2144]), .B(n15082), .Z(n15078) );
  IV U14964 ( .A(p_input[2112]), .Z(n15082) );
  XNOR U14965 ( .A(p_input[2048]), .B(n15083), .Z(n14676) );
  AND U14966 ( .A(n283), .B(n15084), .Z(n15083) );
  XOR U14967 ( .A(p_input[2080]), .B(p_input[2048]), .Z(n15084) );
  XOR U14968 ( .A(n15085), .B(n15086), .Z(n283) );
  AND U14969 ( .A(n15087), .B(n15088), .Z(n15086) );
  XNOR U14970 ( .A(p_input[2111]), .B(n15085), .Z(n15088) );
  XOR U14971 ( .A(n15085), .B(p_input[2079]), .Z(n15087) );
  XOR U14972 ( .A(n15089), .B(n15090), .Z(n15085) );
  AND U14973 ( .A(n15091), .B(n15092), .Z(n15090) );
  XNOR U14974 ( .A(p_input[2110]), .B(n15089), .Z(n15092) );
  XNOR U14975 ( .A(n15089), .B(n14691), .Z(n15091) );
  IV U14976 ( .A(p_input[2078]), .Z(n14691) );
  XOR U14977 ( .A(n15093), .B(n15094), .Z(n15089) );
  AND U14978 ( .A(n15095), .B(n15096), .Z(n15094) );
  XNOR U14979 ( .A(p_input[2109]), .B(n15093), .Z(n15096) );
  XNOR U14980 ( .A(n15093), .B(n14700), .Z(n15095) );
  IV U14981 ( .A(p_input[2077]), .Z(n14700) );
  XOR U14982 ( .A(n15097), .B(n15098), .Z(n15093) );
  AND U14983 ( .A(n15099), .B(n15100), .Z(n15098) );
  XNOR U14984 ( .A(p_input[2108]), .B(n15097), .Z(n15100) );
  XNOR U14985 ( .A(n15097), .B(n14709), .Z(n15099) );
  IV U14986 ( .A(p_input[2076]), .Z(n14709) );
  XOR U14987 ( .A(n15101), .B(n15102), .Z(n15097) );
  AND U14988 ( .A(n15103), .B(n15104), .Z(n15102) );
  XNOR U14989 ( .A(p_input[2107]), .B(n15101), .Z(n15104) );
  XNOR U14990 ( .A(n15101), .B(n14718), .Z(n15103) );
  IV U14991 ( .A(p_input[2075]), .Z(n14718) );
  XOR U14992 ( .A(n15105), .B(n15106), .Z(n15101) );
  AND U14993 ( .A(n15107), .B(n15108), .Z(n15106) );
  XNOR U14994 ( .A(p_input[2106]), .B(n15105), .Z(n15108) );
  XNOR U14995 ( .A(n15105), .B(n14727), .Z(n15107) );
  IV U14996 ( .A(p_input[2074]), .Z(n14727) );
  XOR U14997 ( .A(n15109), .B(n15110), .Z(n15105) );
  AND U14998 ( .A(n15111), .B(n15112), .Z(n15110) );
  XNOR U14999 ( .A(p_input[2105]), .B(n15109), .Z(n15112) );
  XNOR U15000 ( .A(n15109), .B(n14736), .Z(n15111) );
  IV U15001 ( .A(p_input[2073]), .Z(n14736) );
  XOR U15002 ( .A(n15113), .B(n15114), .Z(n15109) );
  AND U15003 ( .A(n15115), .B(n15116), .Z(n15114) );
  XNOR U15004 ( .A(p_input[2104]), .B(n15113), .Z(n15116) );
  XNOR U15005 ( .A(n15113), .B(n14745), .Z(n15115) );
  IV U15006 ( .A(p_input[2072]), .Z(n14745) );
  XOR U15007 ( .A(n15117), .B(n15118), .Z(n15113) );
  AND U15008 ( .A(n15119), .B(n15120), .Z(n15118) );
  XNOR U15009 ( .A(p_input[2103]), .B(n15117), .Z(n15120) );
  XNOR U15010 ( .A(n15117), .B(n14754), .Z(n15119) );
  IV U15011 ( .A(p_input[2071]), .Z(n14754) );
  XOR U15012 ( .A(n15121), .B(n15122), .Z(n15117) );
  AND U15013 ( .A(n15123), .B(n15124), .Z(n15122) );
  XNOR U15014 ( .A(p_input[2102]), .B(n15121), .Z(n15124) );
  XNOR U15015 ( .A(n15121), .B(n14763), .Z(n15123) );
  IV U15016 ( .A(p_input[2070]), .Z(n14763) );
  XOR U15017 ( .A(n15125), .B(n15126), .Z(n15121) );
  AND U15018 ( .A(n15127), .B(n15128), .Z(n15126) );
  XNOR U15019 ( .A(p_input[2101]), .B(n15125), .Z(n15128) );
  XNOR U15020 ( .A(n15125), .B(n14772), .Z(n15127) );
  IV U15021 ( .A(p_input[2069]), .Z(n14772) );
  XOR U15022 ( .A(n15129), .B(n15130), .Z(n15125) );
  AND U15023 ( .A(n15131), .B(n15132), .Z(n15130) );
  XNOR U15024 ( .A(p_input[2100]), .B(n15129), .Z(n15132) );
  XNOR U15025 ( .A(n15129), .B(n14781), .Z(n15131) );
  IV U15026 ( .A(p_input[2068]), .Z(n14781) );
  XOR U15027 ( .A(n15133), .B(n15134), .Z(n15129) );
  AND U15028 ( .A(n15135), .B(n15136), .Z(n15134) );
  XNOR U15029 ( .A(p_input[2099]), .B(n15133), .Z(n15136) );
  XNOR U15030 ( .A(n15133), .B(n14790), .Z(n15135) );
  IV U15031 ( .A(p_input[2067]), .Z(n14790) );
  XOR U15032 ( .A(n15137), .B(n15138), .Z(n15133) );
  AND U15033 ( .A(n15139), .B(n15140), .Z(n15138) );
  XNOR U15034 ( .A(p_input[2098]), .B(n15137), .Z(n15140) );
  XNOR U15035 ( .A(n15137), .B(n14799), .Z(n15139) );
  IV U15036 ( .A(p_input[2066]), .Z(n14799) );
  XOR U15037 ( .A(n15141), .B(n15142), .Z(n15137) );
  AND U15038 ( .A(n15143), .B(n15144), .Z(n15142) );
  XNOR U15039 ( .A(p_input[2097]), .B(n15141), .Z(n15144) );
  XNOR U15040 ( .A(n15141), .B(n14808), .Z(n15143) );
  IV U15041 ( .A(p_input[2065]), .Z(n14808) );
  XOR U15042 ( .A(n15145), .B(n15146), .Z(n15141) );
  AND U15043 ( .A(n15147), .B(n15148), .Z(n15146) );
  XNOR U15044 ( .A(p_input[2096]), .B(n15145), .Z(n15148) );
  XNOR U15045 ( .A(n15145), .B(n14817), .Z(n15147) );
  IV U15046 ( .A(p_input[2064]), .Z(n14817) );
  XOR U15047 ( .A(n15149), .B(n15150), .Z(n15145) );
  AND U15048 ( .A(n15151), .B(n15152), .Z(n15150) );
  XNOR U15049 ( .A(p_input[2095]), .B(n15149), .Z(n15152) );
  XNOR U15050 ( .A(n15149), .B(n14826), .Z(n15151) );
  IV U15051 ( .A(p_input[2063]), .Z(n14826) );
  XOR U15052 ( .A(n15153), .B(n15154), .Z(n15149) );
  AND U15053 ( .A(n15155), .B(n15156), .Z(n15154) );
  XNOR U15054 ( .A(p_input[2094]), .B(n15153), .Z(n15156) );
  XNOR U15055 ( .A(n15153), .B(n14835), .Z(n15155) );
  IV U15056 ( .A(p_input[2062]), .Z(n14835) );
  XOR U15057 ( .A(n15157), .B(n15158), .Z(n15153) );
  AND U15058 ( .A(n15159), .B(n15160), .Z(n15158) );
  XNOR U15059 ( .A(p_input[2093]), .B(n15157), .Z(n15160) );
  XNOR U15060 ( .A(n15157), .B(n14844), .Z(n15159) );
  IV U15061 ( .A(p_input[2061]), .Z(n14844) );
  XOR U15062 ( .A(n15161), .B(n15162), .Z(n15157) );
  AND U15063 ( .A(n15163), .B(n15164), .Z(n15162) );
  XNOR U15064 ( .A(p_input[2092]), .B(n15161), .Z(n15164) );
  XNOR U15065 ( .A(n15161), .B(n14853), .Z(n15163) );
  IV U15066 ( .A(p_input[2060]), .Z(n14853) );
  XOR U15067 ( .A(n15165), .B(n15166), .Z(n15161) );
  AND U15068 ( .A(n15167), .B(n15168), .Z(n15166) );
  XNOR U15069 ( .A(p_input[2091]), .B(n15165), .Z(n15168) );
  XNOR U15070 ( .A(n15165), .B(n14862), .Z(n15167) );
  IV U15071 ( .A(p_input[2059]), .Z(n14862) );
  XOR U15072 ( .A(n15169), .B(n15170), .Z(n15165) );
  AND U15073 ( .A(n15171), .B(n15172), .Z(n15170) );
  XNOR U15074 ( .A(p_input[2090]), .B(n15169), .Z(n15172) );
  XNOR U15075 ( .A(n15169), .B(n14871), .Z(n15171) );
  IV U15076 ( .A(p_input[2058]), .Z(n14871) );
  XOR U15077 ( .A(n15173), .B(n15174), .Z(n15169) );
  AND U15078 ( .A(n15175), .B(n15176), .Z(n15174) );
  XNOR U15079 ( .A(p_input[2089]), .B(n15173), .Z(n15176) );
  XNOR U15080 ( .A(n15173), .B(n14880), .Z(n15175) );
  IV U15081 ( .A(p_input[2057]), .Z(n14880) );
  XOR U15082 ( .A(n15177), .B(n15178), .Z(n15173) );
  AND U15083 ( .A(n15179), .B(n15180), .Z(n15178) );
  XNOR U15084 ( .A(p_input[2088]), .B(n15177), .Z(n15180) );
  XNOR U15085 ( .A(n15177), .B(n14889), .Z(n15179) );
  IV U15086 ( .A(p_input[2056]), .Z(n14889) );
  XOR U15087 ( .A(n15181), .B(n15182), .Z(n15177) );
  AND U15088 ( .A(n15183), .B(n15184), .Z(n15182) );
  XNOR U15089 ( .A(p_input[2087]), .B(n15181), .Z(n15184) );
  XNOR U15090 ( .A(n15181), .B(n14898), .Z(n15183) );
  IV U15091 ( .A(p_input[2055]), .Z(n14898) );
  XOR U15092 ( .A(n15185), .B(n15186), .Z(n15181) );
  AND U15093 ( .A(n15187), .B(n15188), .Z(n15186) );
  XNOR U15094 ( .A(p_input[2086]), .B(n15185), .Z(n15188) );
  XNOR U15095 ( .A(n15185), .B(n14907), .Z(n15187) );
  IV U15096 ( .A(p_input[2054]), .Z(n14907) );
  XOR U15097 ( .A(n15189), .B(n15190), .Z(n15185) );
  AND U15098 ( .A(n15191), .B(n15192), .Z(n15190) );
  XNOR U15099 ( .A(p_input[2085]), .B(n15189), .Z(n15192) );
  XNOR U15100 ( .A(n15189), .B(n14916), .Z(n15191) );
  IV U15101 ( .A(p_input[2053]), .Z(n14916) );
  XOR U15102 ( .A(n15193), .B(n15194), .Z(n15189) );
  AND U15103 ( .A(n15195), .B(n15196), .Z(n15194) );
  XNOR U15104 ( .A(p_input[2084]), .B(n15193), .Z(n15196) );
  XNOR U15105 ( .A(n15193), .B(n14925), .Z(n15195) );
  IV U15106 ( .A(p_input[2052]), .Z(n14925) );
  XOR U15107 ( .A(n15197), .B(n15198), .Z(n15193) );
  AND U15108 ( .A(n15199), .B(n15200), .Z(n15198) );
  XNOR U15109 ( .A(p_input[2083]), .B(n15197), .Z(n15200) );
  XNOR U15110 ( .A(n15197), .B(n14934), .Z(n15199) );
  IV U15111 ( .A(p_input[2051]), .Z(n14934) );
  XOR U15112 ( .A(n15201), .B(n15202), .Z(n15197) );
  AND U15113 ( .A(n15203), .B(n15204), .Z(n15202) );
  XNOR U15114 ( .A(p_input[2082]), .B(n15201), .Z(n15204) );
  XNOR U15115 ( .A(n15201), .B(n14943), .Z(n15203) );
  IV U15116 ( .A(p_input[2050]), .Z(n14943) );
  XNOR U15117 ( .A(n15205), .B(n15206), .Z(n15201) );
  AND U15118 ( .A(n15207), .B(n15208), .Z(n15206) );
  XOR U15119 ( .A(p_input[2081]), .B(n15205), .Z(n15208) );
  XNOR U15120 ( .A(p_input[2049]), .B(n15205), .Z(n15207) );
  AND U15121 ( .A(p_input[2080]), .B(n15209), .Z(n15205) );
  IV U15122 ( .A(p_input[2048]), .Z(n15209) );
  XOR U15123 ( .A(n15210), .B(n15211), .Z(n11) );
  AND U15124 ( .A(n631), .B(n15212), .Z(n15211) );
  XNOR U15125 ( .A(n15213), .B(n15210), .Z(n15212) );
  XOR U15126 ( .A(n15214), .B(n15215), .Z(n631) );
  AND U15127 ( .A(n15216), .B(n15217), .Z(n15215) );
  XOR U15128 ( .A(n15214), .B(n650), .Z(n15217) );
  XOR U15129 ( .A(n15218), .B(n15219), .Z(n650) );
  AND U15130 ( .A(n622), .B(n15220), .Z(n15219) );
  XOR U15131 ( .A(n15221), .B(n15218), .Z(n15220) );
  XNOR U15132 ( .A(n647), .B(n15214), .Z(n15216) );
  XOR U15133 ( .A(n15222), .B(n15223), .Z(n647) );
  AND U15134 ( .A(n619), .B(n15224), .Z(n15223) );
  XOR U15135 ( .A(n15225), .B(n15222), .Z(n15224) );
  XOR U15136 ( .A(n15226), .B(n15227), .Z(n15214) );
  AND U15137 ( .A(n15228), .B(n15229), .Z(n15227) );
  XOR U15138 ( .A(n15226), .B(n662), .Z(n15229) );
  XOR U15139 ( .A(n15230), .B(n15231), .Z(n662) );
  AND U15140 ( .A(n622), .B(n15232), .Z(n15231) );
  XOR U15141 ( .A(n15233), .B(n15230), .Z(n15232) );
  XNOR U15142 ( .A(n659), .B(n15226), .Z(n15228) );
  XOR U15143 ( .A(n15234), .B(n15235), .Z(n659) );
  AND U15144 ( .A(n619), .B(n15236), .Z(n15235) );
  XOR U15145 ( .A(n15237), .B(n15234), .Z(n15236) );
  XOR U15146 ( .A(n15238), .B(n15239), .Z(n15226) );
  AND U15147 ( .A(n15240), .B(n15241), .Z(n15239) );
  XOR U15148 ( .A(n15238), .B(n674), .Z(n15241) );
  XOR U15149 ( .A(n15242), .B(n15243), .Z(n674) );
  AND U15150 ( .A(n622), .B(n15244), .Z(n15243) );
  XOR U15151 ( .A(n15245), .B(n15242), .Z(n15244) );
  XNOR U15152 ( .A(n671), .B(n15238), .Z(n15240) );
  XOR U15153 ( .A(n15246), .B(n15247), .Z(n671) );
  AND U15154 ( .A(n619), .B(n15248), .Z(n15247) );
  XOR U15155 ( .A(n15249), .B(n15246), .Z(n15248) );
  XOR U15156 ( .A(n15250), .B(n15251), .Z(n15238) );
  AND U15157 ( .A(n15252), .B(n15253), .Z(n15251) );
  XOR U15158 ( .A(n15250), .B(n686), .Z(n15253) );
  XOR U15159 ( .A(n15254), .B(n15255), .Z(n686) );
  AND U15160 ( .A(n622), .B(n15256), .Z(n15255) );
  XOR U15161 ( .A(n15257), .B(n15254), .Z(n15256) );
  XNOR U15162 ( .A(n683), .B(n15250), .Z(n15252) );
  XOR U15163 ( .A(n15258), .B(n15259), .Z(n683) );
  AND U15164 ( .A(n619), .B(n15260), .Z(n15259) );
  XOR U15165 ( .A(n15261), .B(n15258), .Z(n15260) );
  XOR U15166 ( .A(n15262), .B(n15263), .Z(n15250) );
  AND U15167 ( .A(n15264), .B(n15265), .Z(n15263) );
  XOR U15168 ( .A(n15262), .B(n698), .Z(n15265) );
  XOR U15169 ( .A(n15266), .B(n15267), .Z(n698) );
  AND U15170 ( .A(n622), .B(n15268), .Z(n15267) );
  XOR U15171 ( .A(n15269), .B(n15266), .Z(n15268) );
  XNOR U15172 ( .A(n695), .B(n15262), .Z(n15264) );
  XOR U15173 ( .A(n15270), .B(n15271), .Z(n695) );
  AND U15174 ( .A(n619), .B(n15272), .Z(n15271) );
  XOR U15175 ( .A(n15273), .B(n15270), .Z(n15272) );
  XOR U15176 ( .A(n15274), .B(n15275), .Z(n15262) );
  AND U15177 ( .A(n15276), .B(n15277), .Z(n15275) );
  XOR U15178 ( .A(n15274), .B(n710), .Z(n15277) );
  XOR U15179 ( .A(n15278), .B(n15279), .Z(n710) );
  AND U15180 ( .A(n622), .B(n15280), .Z(n15279) );
  XOR U15181 ( .A(n15281), .B(n15278), .Z(n15280) );
  XNOR U15182 ( .A(n707), .B(n15274), .Z(n15276) );
  XOR U15183 ( .A(n15282), .B(n15283), .Z(n707) );
  AND U15184 ( .A(n619), .B(n15284), .Z(n15283) );
  XOR U15185 ( .A(n15285), .B(n15282), .Z(n15284) );
  XOR U15186 ( .A(n15286), .B(n15287), .Z(n15274) );
  AND U15187 ( .A(n15288), .B(n15289), .Z(n15287) );
  XOR U15188 ( .A(n15286), .B(n722), .Z(n15289) );
  XOR U15189 ( .A(n15290), .B(n15291), .Z(n722) );
  AND U15190 ( .A(n622), .B(n15292), .Z(n15291) );
  XOR U15191 ( .A(n15293), .B(n15290), .Z(n15292) );
  XNOR U15192 ( .A(n719), .B(n15286), .Z(n15288) );
  XOR U15193 ( .A(n15294), .B(n15295), .Z(n719) );
  AND U15194 ( .A(n619), .B(n15296), .Z(n15295) );
  XOR U15195 ( .A(n15297), .B(n15294), .Z(n15296) );
  XOR U15196 ( .A(n15298), .B(n15299), .Z(n15286) );
  AND U15197 ( .A(n15300), .B(n15301), .Z(n15299) );
  XOR U15198 ( .A(n15298), .B(n734), .Z(n15301) );
  XOR U15199 ( .A(n15302), .B(n15303), .Z(n734) );
  AND U15200 ( .A(n622), .B(n15304), .Z(n15303) );
  XOR U15201 ( .A(n15305), .B(n15302), .Z(n15304) );
  XNOR U15202 ( .A(n731), .B(n15298), .Z(n15300) );
  XOR U15203 ( .A(n15306), .B(n15307), .Z(n731) );
  AND U15204 ( .A(n619), .B(n15308), .Z(n15307) );
  XOR U15205 ( .A(n15309), .B(n15306), .Z(n15308) );
  XOR U15206 ( .A(n15310), .B(n15311), .Z(n15298) );
  AND U15207 ( .A(n15312), .B(n15313), .Z(n15311) );
  XOR U15208 ( .A(n15310), .B(n746), .Z(n15313) );
  XOR U15209 ( .A(n15314), .B(n15315), .Z(n746) );
  AND U15210 ( .A(n622), .B(n15316), .Z(n15315) );
  XOR U15211 ( .A(n15317), .B(n15314), .Z(n15316) );
  XNOR U15212 ( .A(n743), .B(n15310), .Z(n15312) );
  XOR U15213 ( .A(n15318), .B(n15319), .Z(n743) );
  AND U15214 ( .A(n619), .B(n15320), .Z(n15319) );
  XOR U15215 ( .A(n15321), .B(n15318), .Z(n15320) );
  XOR U15216 ( .A(n15322), .B(n15323), .Z(n15310) );
  AND U15217 ( .A(n15324), .B(n15325), .Z(n15323) );
  XOR U15218 ( .A(n15322), .B(n758), .Z(n15325) );
  XOR U15219 ( .A(n15326), .B(n15327), .Z(n758) );
  AND U15220 ( .A(n622), .B(n15328), .Z(n15327) );
  XOR U15221 ( .A(n15329), .B(n15326), .Z(n15328) );
  XNOR U15222 ( .A(n755), .B(n15322), .Z(n15324) );
  XOR U15223 ( .A(n15330), .B(n15331), .Z(n755) );
  AND U15224 ( .A(n619), .B(n15332), .Z(n15331) );
  XOR U15225 ( .A(n15333), .B(n15330), .Z(n15332) );
  XOR U15226 ( .A(n15334), .B(n15335), .Z(n15322) );
  AND U15227 ( .A(n15336), .B(n15337), .Z(n15335) );
  XOR U15228 ( .A(n15334), .B(n770), .Z(n15337) );
  XOR U15229 ( .A(n15338), .B(n15339), .Z(n770) );
  AND U15230 ( .A(n622), .B(n15340), .Z(n15339) );
  XOR U15231 ( .A(n15341), .B(n15338), .Z(n15340) );
  XNOR U15232 ( .A(n767), .B(n15334), .Z(n15336) );
  XOR U15233 ( .A(n15342), .B(n15343), .Z(n767) );
  AND U15234 ( .A(n619), .B(n15344), .Z(n15343) );
  XOR U15235 ( .A(n15345), .B(n15342), .Z(n15344) );
  XOR U15236 ( .A(n15346), .B(n15347), .Z(n15334) );
  AND U15237 ( .A(n15348), .B(n15349), .Z(n15347) );
  XOR U15238 ( .A(n15346), .B(n782), .Z(n15349) );
  XOR U15239 ( .A(n15350), .B(n15351), .Z(n782) );
  AND U15240 ( .A(n622), .B(n15352), .Z(n15351) );
  XOR U15241 ( .A(n15353), .B(n15350), .Z(n15352) );
  XNOR U15242 ( .A(n779), .B(n15346), .Z(n15348) );
  XOR U15243 ( .A(n15354), .B(n15355), .Z(n779) );
  AND U15244 ( .A(n619), .B(n15356), .Z(n15355) );
  XOR U15245 ( .A(n15357), .B(n15354), .Z(n15356) );
  XOR U15246 ( .A(n15358), .B(n15359), .Z(n15346) );
  AND U15247 ( .A(n15360), .B(n15361), .Z(n15359) );
  XOR U15248 ( .A(n15358), .B(n794), .Z(n15361) );
  XOR U15249 ( .A(n15362), .B(n15363), .Z(n794) );
  AND U15250 ( .A(n622), .B(n15364), .Z(n15363) );
  XOR U15251 ( .A(n15365), .B(n15362), .Z(n15364) );
  XNOR U15252 ( .A(n791), .B(n15358), .Z(n15360) );
  XOR U15253 ( .A(n15366), .B(n15367), .Z(n791) );
  AND U15254 ( .A(n619), .B(n15368), .Z(n15367) );
  XOR U15255 ( .A(n15369), .B(n15366), .Z(n15368) );
  XOR U15256 ( .A(n15370), .B(n15371), .Z(n15358) );
  AND U15257 ( .A(n15372), .B(n15373), .Z(n15371) );
  XOR U15258 ( .A(n15370), .B(n806), .Z(n15373) );
  XOR U15259 ( .A(n15374), .B(n15375), .Z(n806) );
  AND U15260 ( .A(n622), .B(n15376), .Z(n15375) );
  XOR U15261 ( .A(n15377), .B(n15374), .Z(n15376) );
  XNOR U15262 ( .A(n803), .B(n15370), .Z(n15372) );
  XOR U15263 ( .A(n15378), .B(n15379), .Z(n803) );
  AND U15264 ( .A(n619), .B(n15380), .Z(n15379) );
  XOR U15265 ( .A(n15381), .B(n15378), .Z(n15380) );
  XOR U15266 ( .A(n15382), .B(n15383), .Z(n15370) );
  AND U15267 ( .A(n15384), .B(n15385), .Z(n15383) );
  XOR U15268 ( .A(n15382), .B(n818), .Z(n15385) );
  XOR U15269 ( .A(n15386), .B(n15387), .Z(n818) );
  AND U15270 ( .A(n622), .B(n15388), .Z(n15387) );
  XOR U15271 ( .A(n15389), .B(n15386), .Z(n15388) );
  XNOR U15272 ( .A(n815), .B(n15382), .Z(n15384) );
  XOR U15273 ( .A(n15390), .B(n15391), .Z(n815) );
  AND U15274 ( .A(n619), .B(n15392), .Z(n15391) );
  XOR U15275 ( .A(n15393), .B(n15390), .Z(n15392) );
  XOR U15276 ( .A(n15394), .B(n15395), .Z(n15382) );
  AND U15277 ( .A(n15396), .B(n15397), .Z(n15395) );
  XOR U15278 ( .A(n15394), .B(n830), .Z(n15397) );
  XOR U15279 ( .A(n15398), .B(n15399), .Z(n830) );
  AND U15280 ( .A(n622), .B(n15400), .Z(n15399) );
  XOR U15281 ( .A(n15401), .B(n15398), .Z(n15400) );
  XNOR U15282 ( .A(n827), .B(n15394), .Z(n15396) );
  XOR U15283 ( .A(n15402), .B(n15403), .Z(n827) );
  AND U15284 ( .A(n619), .B(n15404), .Z(n15403) );
  XOR U15285 ( .A(n15405), .B(n15402), .Z(n15404) );
  XOR U15286 ( .A(n15406), .B(n15407), .Z(n15394) );
  AND U15287 ( .A(n15408), .B(n15409), .Z(n15407) );
  XOR U15288 ( .A(n15406), .B(n842), .Z(n15409) );
  XOR U15289 ( .A(n15410), .B(n15411), .Z(n842) );
  AND U15290 ( .A(n622), .B(n15412), .Z(n15411) );
  XOR U15291 ( .A(n15413), .B(n15410), .Z(n15412) );
  XNOR U15292 ( .A(n839), .B(n15406), .Z(n15408) );
  XOR U15293 ( .A(n15414), .B(n15415), .Z(n839) );
  AND U15294 ( .A(n619), .B(n15416), .Z(n15415) );
  XOR U15295 ( .A(n15417), .B(n15414), .Z(n15416) );
  XOR U15296 ( .A(n15418), .B(n15419), .Z(n15406) );
  AND U15297 ( .A(n15420), .B(n15421), .Z(n15419) );
  XOR U15298 ( .A(n15418), .B(n854), .Z(n15421) );
  XOR U15299 ( .A(n15422), .B(n15423), .Z(n854) );
  AND U15300 ( .A(n622), .B(n15424), .Z(n15423) );
  XOR U15301 ( .A(n15425), .B(n15422), .Z(n15424) );
  XNOR U15302 ( .A(n851), .B(n15418), .Z(n15420) );
  XOR U15303 ( .A(n15426), .B(n15427), .Z(n851) );
  AND U15304 ( .A(n619), .B(n15428), .Z(n15427) );
  XOR U15305 ( .A(n15429), .B(n15426), .Z(n15428) );
  XOR U15306 ( .A(n15430), .B(n15431), .Z(n15418) );
  AND U15307 ( .A(n15432), .B(n15433), .Z(n15431) );
  XOR U15308 ( .A(n15430), .B(n866), .Z(n15433) );
  XOR U15309 ( .A(n15434), .B(n15435), .Z(n866) );
  AND U15310 ( .A(n622), .B(n15436), .Z(n15435) );
  XOR U15311 ( .A(n15437), .B(n15434), .Z(n15436) );
  XNOR U15312 ( .A(n863), .B(n15430), .Z(n15432) );
  XOR U15313 ( .A(n15438), .B(n15439), .Z(n863) );
  AND U15314 ( .A(n619), .B(n15440), .Z(n15439) );
  XOR U15315 ( .A(n15441), .B(n15438), .Z(n15440) );
  XOR U15316 ( .A(n15442), .B(n15443), .Z(n15430) );
  AND U15317 ( .A(n15444), .B(n15445), .Z(n15443) );
  XOR U15318 ( .A(n15442), .B(n878), .Z(n15445) );
  XOR U15319 ( .A(n15446), .B(n15447), .Z(n878) );
  AND U15320 ( .A(n622), .B(n15448), .Z(n15447) );
  XOR U15321 ( .A(n15449), .B(n15446), .Z(n15448) );
  XNOR U15322 ( .A(n875), .B(n15442), .Z(n15444) );
  XOR U15323 ( .A(n15450), .B(n15451), .Z(n875) );
  AND U15324 ( .A(n619), .B(n15452), .Z(n15451) );
  XOR U15325 ( .A(n15453), .B(n15450), .Z(n15452) );
  XOR U15326 ( .A(n15454), .B(n15455), .Z(n15442) );
  AND U15327 ( .A(n15456), .B(n15457), .Z(n15455) );
  XOR U15328 ( .A(n15454), .B(n890), .Z(n15457) );
  XOR U15329 ( .A(n15458), .B(n15459), .Z(n890) );
  AND U15330 ( .A(n622), .B(n15460), .Z(n15459) );
  XOR U15331 ( .A(n15461), .B(n15458), .Z(n15460) );
  XNOR U15332 ( .A(n887), .B(n15454), .Z(n15456) );
  XOR U15333 ( .A(n15462), .B(n15463), .Z(n887) );
  AND U15334 ( .A(n619), .B(n15464), .Z(n15463) );
  XOR U15335 ( .A(n15465), .B(n15462), .Z(n15464) );
  XOR U15336 ( .A(n15466), .B(n15467), .Z(n15454) );
  AND U15337 ( .A(n15468), .B(n15469), .Z(n15467) );
  XOR U15338 ( .A(n15466), .B(n902), .Z(n15469) );
  XOR U15339 ( .A(n15470), .B(n15471), .Z(n902) );
  AND U15340 ( .A(n622), .B(n15472), .Z(n15471) );
  XOR U15341 ( .A(n15473), .B(n15470), .Z(n15472) );
  XNOR U15342 ( .A(n899), .B(n15466), .Z(n15468) );
  XOR U15343 ( .A(n15474), .B(n15475), .Z(n899) );
  AND U15344 ( .A(n619), .B(n15476), .Z(n15475) );
  XOR U15345 ( .A(n15477), .B(n15474), .Z(n15476) );
  XOR U15346 ( .A(n15478), .B(n15479), .Z(n15466) );
  AND U15347 ( .A(n15480), .B(n15481), .Z(n15479) );
  XOR U15348 ( .A(n15478), .B(n914), .Z(n15481) );
  XOR U15349 ( .A(n15482), .B(n15483), .Z(n914) );
  AND U15350 ( .A(n622), .B(n15484), .Z(n15483) );
  XOR U15351 ( .A(n15485), .B(n15482), .Z(n15484) );
  XNOR U15352 ( .A(n911), .B(n15478), .Z(n15480) );
  XOR U15353 ( .A(n15486), .B(n15487), .Z(n911) );
  AND U15354 ( .A(n619), .B(n15488), .Z(n15487) );
  XOR U15355 ( .A(n15489), .B(n15486), .Z(n15488) );
  XOR U15356 ( .A(n15490), .B(n15491), .Z(n15478) );
  AND U15357 ( .A(n15492), .B(n15493), .Z(n15491) );
  XOR U15358 ( .A(n15490), .B(n926), .Z(n15493) );
  XOR U15359 ( .A(n15494), .B(n15495), .Z(n926) );
  AND U15360 ( .A(n622), .B(n15496), .Z(n15495) );
  XOR U15361 ( .A(n15497), .B(n15494), .Z(n15496) );
  XNOR U15362 ( .A(n923), .B(n15490), .Z(n15492) );
  XOR U15363 ( .A(n15498), .B(n15499), .Z(n923) );
  AND U15364 ( .A(n619), .B(n15500), .Z(n15499) );
  XOR U15365 ( .A(n15501), .B(n15498), .Z(n15500) );
  XOR U15366 ( .A(n15502), .B(n15503), .Z(n15490) );
  AND U15367 ( .A(n15504), .B(n15505), .Z(n15503) );
  XOR U15368 ( .A(n15502), .B(n938), .Z(n15505) );
  XOR U15369 ( .A(n15506), .B(n15507), .Z(n938) );
  AND U15370 ( .A(n622), .B(n15508), .Z(n15507) );
  XOR U15371 ( .A(n15509), .B(n15506), .Z(n15508) );
  XNOR U15372 ( .A(n935), .B(n15502), .Z(n15504) );
  XOR U15373 ( .A(n15510), .B(n15511), .Z(n935) );
  AND U15374 ( .A(n619), .B(n15512), .Z(n15511) );
  XOR U15375 ( .A(n15513), .B(n15510), .Z(n15512) );
  XOR U15376 ( .A(n15514), .B(n15515), .Z(n15502) );
  AND U15377 ( .A(n15516), .B(n15517), .Z(n15515) );
  XOR U15378 ( .A(n15514), .B(n950), .Z(n15517) );
  XOR U15379 ( .A(n15518), .B(n15519), .Z(n950) );
  AND U15380 ( .A(n622), .B(n15520), .Z(n15519) );
  XOR U15381 ( .A(n15521), .B(n15518), .Z(n15520) );
  XNOR U15382 ( .A(n947), .B(n15514), .Z(n15516) );
  XOR U15383 ( .A(n15522), .B(n15523), .Z(n947) );
  AND U15384 ( .A(n619), .B(n15524), .Z(n15523) );
  XOR U15385 ( .A(n15525), .B(n15522), .Z(n15524) );
  XOR U15386 ( .A(n15526), .B(n15527), .Z(n15514) );
  AND U15387 ( .A(n15528), .B(n15529), .Z(n15527) );
  XOR U15388 ( .A(n15526), .B(n962), .Z(n15529) );
  XOR U15389 ( .A(n15530), .B(n15531), .Z(n962) );
  AND U15390 ( .A(n622), .B(n15532), .Z(n15531) );
  XOR U15391 ( .A(n15533), .B(n15530), .Z(n15532) );
  XNOR U15392 ( .A(n959), .B(n15526), .Z(n15528) );
  XOR U15393 ( .A(n15534), .B(n15535), .Z(n959) );
  AND U15394 ( .A(n619), .B(n15536), .Z(n15535) );
  XOR U15395 ( .A(n15537), .B(n15534), .Z(n15536) );
  XOR U15396 ( .A(n15538), .B(n15539), .Z(n15526) );
  AND U15397 ( .A(n15540), .B(n15541), .Z(n15539) );
  XOR U15398 ( .A(n15538), .B(n974), .Z(n15541) );
  XOR U15399 ( .A(n15542), .B(n15543), .Z(n974) );
  AND U15400 ( .A(n622), .B(n15544), .Z(n15543) );
  XOR U15401 ( .A(n15545), .B(n15542), .Z(n15544) );
  XNOR U15402 ( .A(n971), .B(n15538), .Z(n15540) );
  XOR U15403 ( .A(n15546), .B(n15547), .Z(n971) );
  AND U15404 ( .A(n619), .B(n15548), .Z(n15547) );
  XOR U15405 ( .A(n15549), .B(n15546), .Z(n15548) );
  XOR U15406 ( .A(n15550), .B(n15551), .Z(n15538) );
  AND U15407 ( .A(n15552), .B(n15553), .Z(n15551) );
  XOR U15408 ( .A(n15550), .B(n986), .Z(n15553) );
  XOR U15409 ( .A(n15554), .B(n15555), .Z(n986) );
  AND U15410 ( .A(n622), .B(n15556), .Z(n15555) );
  XOR U15411 ( .A(n15557), .B(n15554), .Z(n15556) );
  XNOR U15412 ( .A(n983), .B(n15550), .Z(n15552) );
  XOR U15413 ( .A(n15558), .B(n15559), .Z(n983) );
  AND U15414 ( .A(n619), .B(n15560), .Z(n15559) );
  XOR U15415 ( .A(n15561), .B(n15558), .Z(n15560) );
  XOR U15416 ( .A(n15562), .B(n15563), .Z(n15550) );
  AND U15417 ( .A(n15564), .B(n15565), .Z(n15563) );
  XOR U15418 ( .A(n998), .B(n15562), .Z(n15565) );
  XOR U15419 ( .A(n15566), .B(n15567), .Z(n998) );
  AND U15420 ( .A(n622), .B(n15568), .Z(n15567) );
  XOR U15421 ( .A(n15566), .B(n15569), .Z(n15568) );
  XNOR U15422 ( .A(n15562), .B(n995), .Z(n15564) );
  XOR U15423 ( .A(n15570), .B(n15571), .Z(n995) );
  AND U15424 ( .A(n619), .B(n15572), .Z(n15571) );
  XOR U15425 ( .A(n15570), .B(n15573), .Z(n15572) );
  XOR U15426 ( .A(n15574), .B(n15575), .Z(n15562) );
  AND U15427 ( .A(n15576), .B(n15577), .Z(n15575) );
  XNOR U15428 ( .A(n15578), .B(n1010), .Z(n15577) );
  XOR U15429 ( .A(n15579), .B(n15580), .Z(n1010) );
  AND U15430 ( .A(n622), .B(n15581), .Z(n15580) );
  XOR U15431 ( .A(n15582), .B(n15579), .Z(n15581) );
  XNOR U15432 ( .A(n1007), .B(n15574), .Z(n15576) );
  XOR U15433 ( .A(n15583), .B(n15584), .Z(n1007) );
  AND U15434 ( .A(n619), .B(n15585), .Z(n15584) );
  XOR U15435 ( .A(n15586), .B(n15583), .Z(n15585) );
  IV U15436 ( .A(n15578), .Z(n15574) );
  AND U15437 ( .A(n15210), .B(n15213), .Z(n15578) );
  XNOR U15438 ( .A(n15587), .B(n15588), .Z(n15213) );
  AND U15439 ( .A(n622), .B(n15589), .Z(n15588) );
  XNOR U15440 ( .A(n15590), .B(n15587), .Z(n15589) );
  XOR U15441 ( .A(n15591), .B(n15592), .Z(n622) );
  AND U15442 ( .A(n15593), .B(n15594), .Z(n15592) );
  XOR U15443 ( .A(n15591), .B(n15221), .Z(n15594) );
  XOR U15444 ( .A(n15595), .B(n15596), .Z(n15221) );
  AND U15445 ( .A(n590), .B(n15597), .Z(n15596) );
  XOR U15446 ( .A(n15598), .B(n15595), .Z(n15597) );
  XNOR U15447 ( .A(n15218), .B(n15591), .Z(n15593) );
  XOR U15448 ( .A(n15599), .B(n15600), .Z(n15218) );
  AND U15449 ( .A(n588), .B(n15601), .Z(n15600) );
  XOR U15450 ( .A(n15602), .B(n15599), .Z(n15601) );
  XOR U15451 ( .A(n15603), .B(n15604), .Z(n15591) );
  AND U15452 ( .A(n15605), .B(n15606), .Z(n15604) );
  XOR U15453 ( .A(n15603), .B(n15233), .Z(n15606) );
  XOR U15454 ( .A(n15607), .B(n15608), .Z(n15233) );
  AND U15455 ( .A(n590), .B(n15609), .Z(n15608) );
  XOR U15456 ( .A(n15610), .B(n15607), .Z(n15609) );
  XNOR U15457 ( .A(n15230), .B(n15603), .Z(n15605) );
  XOR U15458 ( .A(n15611), .B(n15612), .Z(n15230) );
  AND U15459 ( .A(n588), .B(n15613), .Z(n15612) );
  XOR U15460 ( .A(n15614), .B(n15611), .Z(n15613) );
  XOR U15461 ( .A(n15615), .B(n15616), .Z(n15603) );
  AND U15462 ( .A(n15617), .B(n15618), .Z(n15616) );
  XOR U15463 ( .A(n15615), .B(n15245), .Z(n15618) );
  XOR U15464 ( .A(n15619), .B(n15620), .Z(n15245) );
  AND U15465 ( .A(n590), .B(n15621), .Z(n15620) );
  XOR U15466 ( .A(n15622), .B(n15619), .Z(n15621) );
  XNOR U15467 ( .A(n15242), .B(n15615), .Z(n15617) );
  XOR U15468 ( .A(n15623), .B(n15624), .Z(n15242) );
  AND U15469 ( .A(n588), .B(n15625), .Z(n15624) );
  XOR U15470 ( .A(n15626), .B(n15623), .Z(n15625) );
  XOR U15471 ( .A(n15627), .B(n15628), .Z(n15615) );
  AND U15472 ( .A(n15629), .B(n15630), .Z(n15628) );
  XOR U15473 ( .A(n15627), .B(n15257), .Z(n15630) );
  XOR U15474 ( .A(n15631), .B(n15632), .Z(n15257) );
  AND U15475 ( .A(n590), .B(n15633), .Z(n15632) );
  XOR U15476 ( .A(n15634), .B(n15631), .Z(n15633) );
  XNOR U15477 ( .A(n15254), .B(n15627), .Z(n15629) );
  XOR U15478 ( .A(n15635), .B(n15636), .Z(n15254) );
  AND U15479 ( .A(n588), .B(n15637), .Z(n15636) );
  XOR U15480 ( .A(n15638), .B(n15635), .Z(n15637) );
  XOR U15481 ( .A(n15639), .B(n15640), .Z(n15627) );
  AND U15482 ( .A(n15641), .B(n15642), .Z(n15640) );
  XOR U15483 ( .A(n15639), .B(n15269), .Z(n15642) );
  XOR U15484 ( .A(n15643), .B(n15644), .Z(n15269) );
  AND U15485 ( .A(n590), .B(n15645), .Z(n15644) );
  XOR U15486 ( .A(n15646), .B(n15643), .Z(n15645) );
  XNOR U15487 ( .A(n15266), .B(n15639), .Z(n15641) );
  XOR U15488 ( .A(n15647), .B(n15648), .Z(n15266) );
  AND U15489 ( .A(n588), .B(n15649), .Z(n15648) );
  XOR U15490 ( .A(n15650), .B(n15647), .Z(n15649) );
  XOR U15491 ( .A(n15651), .B(n15652), .Z(n15639) );
  AND U15492 ( .A(n15653), .B(n15654), .Z(n15652) );
  XOR U15493 ( .A(n15651), .B(n15281), .Z(n15654) );
  XOR U15494 ( .A(n15655), .B(n15656), .Z(n15281) );
  AND U15495 ( .A(n590), .B(n15657), .Z(n15656) );
  XOR U15496 ( .A(n15658), .B(n15655), .Z(n15657) );
  XNOR U15497 ( .A(n15278), .B(n15651), .Z(n15653) );
  XOR U15498 ( .A(n15659), .B(n15660), .Z(n15278) );
  AND U15499 ( .A(n588), .B(n15661), .Z(n15660) );
  XOR U15500 ( .A(n15662), .B(n15659), .Z(n15661) );
  XOR U15501 ( .A(n15663), .B(n15664), .Z(n15651) );
  AND U15502 ( .A(n15665), .B(n15666), .Z(n15664) );
  XOR U15503 ( .A(n15663), .B(n15293), .Z(n15666) );
  XOR U15504 ( .A(n15667), .B(n15668), .Z(n15293) );
  AND U15505 ( .A(n590), .B(n15669), .Z(n15668) );
  XOR U15506 ( .A(n15670), .B(n15667), .Z(n15669) );
  XNOR U15507 ( .A(n15290), .B(n15663), .Z(n15665) );
  XOR U15508 ( .A(n15671), .B(n15672), .Z(n15290) );
  AND U15509 ( .A(n588), .B(n15673), .Z(n15672) );
  XOR U15510 ( .A(n15674), .B(n15671), .Z(n15673) );
  XOR U15511 ( .A(n15675), .B(n15676), .Z(n15663) );
  AND U15512 ( .A(n15677), .B(n15678), .Z(n15676) );
  XOR U15513 ( .A(n15675), .B(n15305), .Z(n15678) );
  XOR U15514 ( .A(n15679), .B(n15680), .Z(n15305) );
  AND U15515 ( .A(n590), .B(n15681), .Z(n15680) );
  XOR U15516 ( .A(n15682), .B(n15679), .Z(n15681) );
  XNOR U15517 ( .A(n15302), .B(n15675), .Z(n15677) );
  XOR U15518 ( .A(n15683), .B(n15684), .Z(n15302) );
  AND U15519 ( .A(n588), .B(n15685), .Z(n15684) );
  XOR U15520 ( .A(n15686), .B(n15683), .Z(n15685) );
  XOR U15521 ( .A(n15687), .B(n15688), .Z(n15675) );
  AND U15522 ( .A(n15689), .B(n15690), .Z(n15688) );
  XOR U15523 ( .A(n15687), .B(n15317), .Z(n15690) );
  XOR U15524 ( .A(n15691), .B(n15692), .Z(n15317) );
  AND U15525 ( .A(n590), .B(n15693), .Z(n15692) );
  XOR U15526 ( .A(n15694), .B(n15691), .Z(n15693) );
  XNOR U15527 ( .A(n15314), .B(n15687), .Z(n15689) );
  XOR U15528 ( .A(n15695), .B(n15696), .Z(n15314) );
  AND U15529 ( .A(n588), .B(n15697), .Z(n15696) );
  XOR U15530 ( .A(n15698), .B(n15695), .Z(n15697) );
  XOR U15531 ( .A(n15699), .B(n15700), .Z(n15687) );
  AND U15532 ( .A(n15701), .B(n15702), .Z(n15700) );
  XOR U15533 ( .A(n15699), .B(n15329), .Z(n15702) );
  XOR U15534 ( .A(n15703), .B(n15704), .Z(n15329) );
  AND U15535 ( .A(n590), .B(n15705), .Z(n15704) );
  XOR U15536 ( .A(n15706), .B(n15703), .Z(n15705) );
  XNOR U15537 ( .A(n15326), .B(n15699), .Z(n15701) );
  XOR U15538 ( .A(n15707), .B(n15708), .Z(n15326) );
  AND U15539 ( .A(n588), .B(n15709), .Z(n15708) );
  XOR U15540 ( .A(n15710), .B(n15707), .Z(n15709) );
  XOR U15541 ( .A(n15711), .B(n15712), .Z(n15699) );
  AND U15542 ( .A(n15713), .B(n15714), .Z(n15712) );
  XOR U15543 ( .A(n15711), .B(n15341), .Z(n15714) );
  XOR U15544 ( .A(n15715), .B(n15716), .Z(n15341) );
  AND U15545 ( .A(n590), .B(n15717), .Z(n15716) );
  XOR U15546 ( .A(n15718), .B(n15715), .Z(n15717) );
  XNOR U15547 ( .A(n15338), .B(n15711), .Z(n15713) );
  XOR U15548 ( .A(n15719), .B(n15720), .Z(n15338) );
  AND U15549 ( .A(n588), .B(n15721), .Z(n15720) );
  XOR U15550 ( .A(n15722), .B(n15719), .Z(n15721) );
  XOR U15551 ( .A(n15723), .B(n15724), .Z(n15711) );
  AND U15552 ( .A(n15725), .B(n15726), .Z(n15724) );
  XOR U15553 ( .A(n15723), .B(n15353), .Z(n15726) );
  XOR U15554 ( .A(n15727), .B(n15728), .Z(n15353) );
  AND U15555 ( .A(n590), .B(n15729), .Z(n15728) );
  XOR U15556 ( .A(n15730), .B(n15727), .Z(n15729) );
  XNOR U15557 ( .A(n15350), .B(n15723), .Z(n15725) );
  XOR U15558 ( .A(n15731), .B(n15732), .Z(n15350) );
  AND U15559 ( .A(n588), .B(n15733), .Z(n15732) );
  XOR U15560 ( .A(n15734), .B(n15731), .Z(n15733) );
  XOR U15561 ( .A(n15735), .B(n15736), .Z(n15723) );
  AND U15562 ( .A(n15737), .B(n15738), .Z(n15736) );
  XOR U15563 ( .A(n15735), .B(n15365), .Z(n15738) );
  XOR U15564 ( .A(n15739), .B(n15740), .Z(n15365) );
  AND U15565 ( .A(n590), .B(n15741), .Z(n15740) );
  XOR U15566 ( .A(n15742), .B(n15739), .Z(n15741) );
  XNOR U15567 ( .A(n15362), .B(n15735), .Z(n15737) );
  XOR U15568 ( .A(n15743), .B(n15744), .Z(n15362) );
  AND U15569 ( .A(n588), .B(n15745), .Z(n15744) );
  XOR U15570 ( .A(n15746), .B(n15743), .Z(n15745) );
  XOR U15571 ( .A(n15747), .B(n15748), .Z(n15735) );
  AND U15572 ( .A(n15749), .B(n15750), .Z(n15748) );
  XOR U15573 ( .A(n15747), .B(n15377), .Z(n15750) );
  XOR U15574 ( .A(n15751), .B(n15752), .Z(n15377) );
  AND U15575 ( .A(n590), .B(n15753), .Z(n15752) );
  XOR U15576 ( .A(n15754), .B(n15751), .Z(n15753) );
  XNOR U15577 ( .A(n15374), .B(n15747), .Z(n15749) );
  XOR U15578 ( .A(n15755), .B(n15756), .Z(n15374) );
  AND U15579 ( .A(n588), .B(n15757), .Z(n15756) );
  XOR U15580 ( .A(n15758), .B(n15755), .Z(n15757) );
  XOR U15581 ( .A(n15759), .B(n15760), .Z(n15747) );
  AND U15582 ( .A(n15761), .B(n15762), .Z(n15760) );
  XOR U15583 ( .A(n15759), .B(n15389), .Z(n15762) );
  XOR U15584 ( .A(n15763), .B(n15764), .Z(n15389) );
  AND U15585 ( .A(n590), .B(n15765), .Z(n15764) );
  XOR U15586 ( .A(n15766), .B(n15763), .Z(n15765) );
  XNOR U15587 ( .A(n15386), .B(n15759), .Z(n15761) );
  XOR U15588 ( .A(n15767), .B(n15768), .Z(n15386) );
  AND U15589 ( .A(n588), .B(n15769), .Z(n15768) );
  XOR U15590 ( .A(n15770), .B(n15767), .Z(n15769) );
  XOR U15591 ( .A(n15771), .B(n15772), .Z(n15759) );
  AND U15592 ( .A(n15773), .B(n15774), .Z(n15772) );
  XOR U15593 ( .A(n15771), .B(n15401), .Z(n15774) );
  XOR U15594 ( .A(n15775), .B(n15776), .Z(n15401) );
  AND U15595 ( .A(n590), .B(n15777), .Z(n15776) );
  XOR U15596 ( .A(n15778), .B(n15775), .Z(n15777) );
  XNOR U15597 ( .A(n15398), .B(n15771), .Z(n15773) );
  XOR U15598 ( .A(n15779), .B(n15780), .Z(n15398) );
  AND U15599 ( .A(n588), .B(n15781), .Z(n15780) );
  XOR U15600 ( .A(n15782), .B(n15779), .Z(n15781) );
  XOR U15601 ( .A(n15783), .B(n15784), .Z(n15771) );
  AND U15602 ( .A(n15785), .B(n15786), .Z(n15784) );
  XOR U15603 ( .A(n15783), .B(n15413), .Z(n15786) );
  XOR U15604 ( .A(n15787), .B(n15788), .Z(n15413) );
  AND U15605 ( .A(n590), .B(n15789), .Z(n15788) );
  XOR U15606 ( .A(n15790), .B(n15787), .Z(n15789) );
  XNOR U15607 ( .A(n15410), .B(n15783), .Z(n15785) );
  XOR U15608 ( .A(n15791), .B(n15792), .Z(n15410) );
  AND U15609 ( .A(n588), .B(n15793), .Z(n15792) );
  XOR U15610 ( .A(n15794), .B(n15791), .Z(n15793) );
  XOR U15611 ( .A(n15795), .B(n15796), .Z(n15783) );
  AND U15612 ( .A(n15797), .B(n15798), .Z(n15796) );
  XOR U15613 ( .A(n15795), .B(n15425), .Z(n15798) );
  XOR U15614 ( .A(n15799), .B(n15800), .Z(n15425) );
  AND U15615 ( .A(n590), .B(n15801), .Z(n15800) );
  XOR U15616 ( .A(n15802), .B(n15799), .Z(n15801) );
  XNOR U15617 ( .A(n15422), .B(n15795), .Z(n15797) );
  XOR U15618 ( .A(n15803), .B(n15804), .Z(n15422) );
  AND U15619 ( .A(n588), .B(n15805), .Z(n15804) );
  XOR U15620 ( .A(n15806), .B(n15803), .Z(n15805) );
  XOR U15621 ( .A(n15807), .B(n15808), .Z(n15795) );
  AND U15622 ( .A(n15809), .B(n15810), .Z(n15808) );
  XOR U15623 ( .A(n15807), .B(n15437), .Z(n15810) );
  XOR U15624 ( .A(n15811), .B(n15812), .Z(n15437) );
  AND U15625 ( .A(n590), .B(n15813), .Z(n15812) );
  XOR U15626 ( .A(n15814), .B(n15811), .Z(n15813) );
  XNOR U15627 ( .A(n15434), .B(n15807), .Z(n15809) );
  XOR U15628 ( .A(n15815), .B(n15816), .Z(n15434) );
  AND U15629 ( .A(n588), .B(n15817), .Z(n15816) );
  XOR U15630 ( .A(n15818), .B(n15815), .Z(n15817) );
  XOR U15631 ( .A(n15819), .B(n15820), .Z(n15807) );
  AND U15632 ( .A(n15821), .B(n15822), .Z(n15820) );
  XOR U15633 ( .A(n15819), .B(n15449), .Z(n15822) );
  XOR U15634 ( .A(n15823), .B(n15824), .Z(n15449) );
  AND U15635 ( .A(n590), .B(n15825), .Z(n15824) );
  XOR U15636 ( .A(n15826), .B(n15823), .Z(n15825) );
  XNOR U15637 ( .A(n15446), .B(n15819), .Z(n15821) );
  XOR U15638 ( .A(n15827), .B(n15828), .Z(n15446) );
  AND U15639 ( .A(n588), .B(n15829), .Z(n15828) );
  XOR U15640 ( .A(n15830), .B(n15827), .Z(n15829) );
  XOR U15641 ( .A(n15831), .B(n15832), .Z(n15819) );
  AND U15642 ( .A(n15833), .B(n15834), .Z(n15832) );
  XOR U15643 ( .A(n15831), .B(n15461), .Z(n15834) );
  XOR U15644 ( .A(n15835), .B(n15836), .Z(n15461) );
  AND U15645 ( .A(n590), .B(n15837), .Z(n15836) );
  XOR U15646 ( .A(n15838), .B(n15835), .Z(n15837) );
  XNOR U15647 ( .A(n15458), .B(n15831), .Z(n15833) );
  XOR U15648 ( .A(n15839), .B(n15840), .Z(n15458) );
  AND U15649 ( .A(n588), .B(n15841), .Z(n15840) );
  XOR U15650 ( .A(n15842), .B(n15839), .Z(n15841) );
  XOR U15651 ( .A(n15843), .B(n15844), .Z(n15831) );
  AND U15652 ( .A(n15845), .B(n15846), .Z(n15844) );
  XOR U15653 ( .A(n15843), .B(n15473), .Z(n15846) );
  XOR U15654 ( .A(n15847), .B(n15848), .Z(n15473) );
  AND U15655 ( .A(n590), .B(n15849), .Z(n15848) );
  XOR U15656 ( .A(n15850), .B(n15847), .Z(n15849) );
  XNOR U15657 ( .A(n15470), .B(n15843), .Z(n15845) );
  XOR U15658 ( .A(n15851), .B(n15852), .Z(n15470) );
  AND U15659 ( .A(n588), .B(n15853), .Z(n15852) );
  XOR U15660 ( .A(n15854), .B(n15851), .Z(n15853) );
  XOR U15661 ( .A(n15855), .B(n15856), .Z(n15843) );
  AND U15662 ( .A(n15857), .B(n15858), .Z(n15856) );
  XOR U15663 ( .A(n15855), .B(n15485), .Z(n15858) );
  XOR U15664 ( .A(n15859), .B(n15860), .Z(n15485) );
  AND U15665 ( .A(n590), .B(n15861), .Z(n15860) );
  XOR U15666 ( .A(n15862), .B(n15859), .Z(n15861) );
  XNOR U15667 ( .A(n15482), .B(n15855), .Z(n15857) );
  XOR U15668 ( .A(n15863), .B(n15864), .Z(n15482) );
  AND U15669 ( .A(n588), .B(n15865), .Z(n15864) );
  XOR U15670 ( .A(n15866), .B(n15863), .Z(n15865) );
  XOR U15671 ( .A(n15867), .B(n15868), .Z(n15855) );
  AND U15672 ( .A(n15869), .B(n15870), .Z(n15868) );
  XOR U15673 ( .A(n15867), .B(n15497), .Z(n15870) );
  XOR U15674 ( .A(n15871), .B(n15872), .Z(n15497) );
  AND U15675 ( .A(n590), .B(n15873), .Z(n15872) );
  XOR U15676 ( .A(n15874), .B(n15871), .Z(n15873) );
  XNOR U15677 ( .A(n15494), .B(n15867), .Z(n15869) );
  XOR U15678 ( .A(n15875), .B(n15876), .Z(n15494) );
  AND U15679 ( .A(n588), .B(n15877), .Z(n15876) );
  XOR U15680 ( .A(n15878), .B(n15875), .Z(n15877) );
  XOR U15681 ( .A(n15879), .B(n15880), .Z(n15867) );
  AND U15682 ( .A(n15881), .B(n15882), .Z(n15880) );
  XOR U15683 ( .A(n15879), .B(n15509), .Z(n15882) );
  XOR U15684 ( .A(n15883), .B(n15884), .Z(n15509) );
  AND U15685 ( .A(n590), .B(n15885), .Z(n15884) );
  XOR U15686 ( .A(n15886), .B(n15883), .Z(n15885) );
  XNOR U15687 ( .A(n15506), .B(n15879), .Z(n15881) );
  XOR U15688 ( .A(n15887), .B(n15888), .Z(n15506) );
  AND U15689 ( .A(n588), .B(n15889), .Z(n15888) );
  XOR U15690 ( .A(n15890), .B(n15887), .Z(n15889) );
  XOR U15691 ( .A(n15891), .B(n15892), .Z(n15879) );
  AND U15692 ( .A(n15893), .B(n15894), .Z(n15892) );
  XOR U15693 ( .A(n15891), .B(n15521), .Z(n15894) );
  XOR U15694 ( .A(n15895), .B(n15896), .Z(n15521) );
  AND U15695 ( .A(n590), .B(n15897), .Z(n15896) );
  XOR U15696 ( .A(n15898), .B(n15895), .Z(n15897) );
  XNOR U15697 ( .A(n15518), .B(n15891), .Z(n15893) );
  XOR U15698 ( .A(n15899), .B(n15900), .Z(n15518) );
  AND U15699 ( .A(n588), .B(n15901), .Z(n15900) );
  XOR U15700 ( .A(n15902), .B(n15899), .Z(n15901) );
  XOR U15701 ( .A(n15903), .B(n15904), .Z(n15891) );
  AND U15702 ( .A(n15905), .B(n15906), .Z(n15904) );
  XOR U15703 ( .A(n15903), .B(n15533), .Z(n15906) );
  XOR U15704 ( .A(n15907), .B(n15908), .Z(n15533) );
  AND U15705 ( .A(n590), .B(n15909), .Z(n15908) );
  XOR U15706 ( .A(n15910), .B(n15907), .Z(n15909) );
  XNOR U15707 ( .A(n15530), .B(n15903), .Z(n15905) );
  XOR U15708 ( .A(n15911), .B(n15912), .Z(n15530) );
  AND U15709 ( .A(n588), .B(n15913), .Z(n15912) );
  XOR U15710 ( .A(n15914), .B(n15911), .Z(n15913) );
  XOR U15711 ( .A(n15915), .B(n15916), .Z(n15903) );
  AND U15712 ( .A(n15917), .B(n15918), .Z(n15916) );
  XOR U15713 ( .A(n15915), .B(n15545), .Z(n15918) );
  XOR U15714 ( .A(n15919), .B(n15920), .Z(n15545) );
  AND U15715 ( .A(n590), .B(n15921), .Z(n15920) );
  XOR U15716 ( .A(n15922), .B(n15919), .Z(n15921) );
  XNOR U15717 ( .A(n15542), .B(n15915), .Z(n15917) );
  XOR U15718 ( .A(n15923), .B(n15924), .Z(n15542) );
  AND U15719 ( .A(n588), .B(n15925), .Z(n15924) );
  XOR U15720 ( .A(n15926), .B(n15923), .Z(n15925) );
  XOR U15721 ( .A(n15927), .B(n15928), .Z(n15915) );
  AND U15722 ( .A(n15929), .B(n15930), .Z(n15928) );
  XOR U15723 ( .A(n15927), .B(n15557), .Z(n15930) );
  XOR U15724 ( .A(n15931), .B(n15932), .Z(n15557) );
  AND U15725 ( .A(n590), .B(n15933), .Z(n15932) );
  XOR U15726 ( .A(n15934), .B(n15931), .Z(n15933) );
  XNOR U15727 ( .A(n15554), .B(n15927), .Z(n15929) );
  XOR U15728 ( .A(n15935), .B(n15936), .Z(n15554) );
  AND U15729 ( .A(n588), .B(n15937), .Z(n15936) );
  XOR U15730 ( .A(n15938), .B(n15935), .Z(n15937) );
  XOR U15731 ( .A(n15939), .B(n15940), .Z(n15927) );
  AND U15732 ( .A(n15941), .B(n15942), .Z(n15940) );
  XOR U15733 ( .A(n15569), .B(n15939), .Z(n15942) );
  XOR U15734 ( .A(n15943), .B(n15944), .Z(n15569) );
  AND U15735 ( .A(n590), .B(n15945), .Z(n15944) );
  XOR U15736 ( .A(n15943), .B(n15946), .Z(n15945) );
  XNOR U15737 ( .A(n15939), .B(n15566), .Z(n15941) );
  XOR U15738 ( .A(n15947), .B(n15948), .Z(n15566) );
  AND U15739 ( .A(n588), .B(n15949), .Z(n15948) );
  XOR U15740 ( .A(n15947), .B(n15950), .Z(n15949) );
  XOR U15741 ( .A(n15951), .B(n15952), .Z(n15939) );
  AND U15742 ( .A(n15953), .B(n15954), .Z(n15952) );
  XNOR U15743 ( .A(n15955), .B(n15582), .Z(n15954) );
  XOR U15744 ( .A(n15956), .B(n15957), .Z(n15582) );
  AND U15745 ( .A(n590), .B(n15958), .Z(n15957) );
  XOR U15746 ( .A(n15959), .B(n15956), .Z(n15958) );
  XNOR U15747 ( .A(n15579), .B(n15951), .Z(n15953) );
  XOR U15748 ( .A(n15960), .B(n15961), .Z(n15579) );
  AND U15749 ( .A(n588), .B(n15962), .Z(n15961) );
  XOR U15750 ( .A(n15963), .B(n15960), .Z(n15962) );
  IV U15751 ( .A(n15955), .Z(n15951) );
  AND U15752 ( .A(n15587), .B(n15590), .Z(n15955) );
  XNOR U15753 ( .A(n15964), .B(n15965), .Z(n15590) );
  AND U15754 ( .A(n590), .B(n15966), .Z(n15965) );
  XNOR U15755 ( .A(n15967), .B(n15964), .Z(n15966) );
  XOR U15756 ( .A(n15968), .B(n15969), .Z(n590) );
  AND U15757 ( .A(n15970), .B(n15971), .Z(n15969) );
  XOR U15758 ( .A(n15968), .B(n15598), .Z(n15971) );
  XOR U15759 ( .A(n15972), .B(n15973), .Z(n15598) );
  AND U15760 ( .A(n518), .B(n15974), .Z(n15973) );
  XOR U15761 ( .A(n15975), .B(n15972), .Z(n15974) );
  XNOR U15762 ( .A(n15595), .B(n15968), .Z(n15970) );
  XOR U15763 ( .A(n15976), .B(n15977), .Z(n15595) );
  AND U15764 ( .A(n516), .B(n15978), .Z(n15977) );
  XOR U15765 ( .A(n15979), .B(n15976), .Z(n15978) );
  XOR U15766 ( .A(n15980), .B(n15981), .Z(n15968) );
  AND U15767 ( .A(n15982), .B(n15983), .Z(n15981) );
  XOR U15768 ( .A(n15980), .B(n15610), .Z(n15983) );
  XOR U15769 ( .A(n15984), .B(n15985), .Z(n15610) );
  AND U15770 ( .A(n518), .B(n15986), .Z(n15985) );
  XOR U15771 ( .A(n15987), .B(n15984), .Z(n15986) );
  XNOR U15772 ( .A(n15607), .B(n15980), .Z(n15982) );
  XOR U15773 ( .A(n15988), .B(n15989), .Z(n15607) );
  AND U15774 ( .A(n516), .B(n15990), .Z(n15989) );
  XOR U15775 ( .A(n15991), .B(n15988), .Z(n15990) );
  XOR U15776 ( .A(n15992), .B(n15993), .Z(n15980) );
  AND U15777 ( .A(n15994), .B(n15995), .Z(n15993) );
  XOR U15778 ( .A(n15992), .B(n15622), .Z(n15995) );
  XOR U15779 ( .A(n15996), .B(n15997), .Z(n15622) );
  AND U15780 ( .A(n518), .B(n15998), .Z(n15997) );
  XOR U15781 ( .A(n15999), .B(n15996), .Z(n15998) );
  XNOR U15782 ( .A(n15619), .B(n15992), .Z(n15994) );
  XOR U15783 ( .A(n16000), .B(n16001), .Z(n15619) );
  AND U15784 ( .A(n516), .B(n16002), .Z(n16001) );
  XOR U15785 ( .A(n16003), .B(n16000), .Z(n16002) );
  XOR U15786 ( .A(n16004), .B(n16005), .Z(n15992) );
  AND U15787 ( .A(n16006), .B(n16007), .Z(n16005) );
  XOR U15788 ( .A(n16004), .B(n15634), .Z(n16007) );
  XOR U15789 ( .A(n16008), .B(n16009), .Z(n15634) );
  AND U15790 ( .A(n518), .B(n16010), .Z(n16009) );
  XOR U15791 ( .A(n16011), .B(n16008), .Z(n16010) );
  XNOR U15792 ( .A(n15631), .B(n16004), .Z(n16006) );
  XOR U15793 ( .A(n16012), .B(n16013), .Z(n15631) );
  AND U15794 ( .A(n516), .B(n16014), .Z(n16013) );
  XOR U15795 ( .A(n16015), .B(n16012), .Z(n16014) );
  XOR U15796 ( .A(n16016), .B(n16017), .Z(n16004) );
  AND U15797 ( .A(n16018), .B(n16019), .Z(n16017) );
  XOR U15798 ( .A(n16016), .B(n15646), .Z(n16019) );
  XOR U15799 ( .A(n16020), .B(n16021), .Z(n15646) );
  AND U15800 ( .A(n518), .B(n16022), .Z(n16021) );
  XOR U15801 ( .A(n16023), .B(n16020), .Z(n16022) );
  XNOR U15802 ( .A(n15643), .B(n16016), .Z(n16018) );
  XOR U15803 ( .A(n16024), .B(n16025), .Z(n15643) );
  AND U15804 ( .A(n516), .B(n16026), .Z(n16025) );
  XOR U15805 ( .A(n16027), .B(n16024), .Z(n16026) );
  XOR U15806 ( .A(n16028), .B(n16029), .Z(n16016) );
  AND U15807 ( .A(n16030), .B(n16031), .Z(n16029) );
  XOR U15808 ( .A(n16028), .B(n15658), .Z(n16031) );
  XOR U15809 ( .A(n16032), .B(n16033), .Z(n15658) );
  AND U15810 ( .A(n518), .B(n16034), .Z(n16033) );
  XOR U15811 ( .A(n16035), .B(n16032), .Z(n16034) );
  XNOR U15812 ( .A(n15655), .B(n16028), .Z(n16030) );
  XOR U15813 ( .A(n16036), .B(n16037), .Z(n15655) );
  AND U15814 ( .A(n516), .B(n16038), .Z(n16037) );
  XOR U15815 ( .A(n16039), .B(n16036), .Z(n16038) );
  XOR U15816 ( .A(n16040), .B(n16041), .Z(n16028) );
  AND U15817 ( .A(n16042), .B(n16043), .Z(n16041) );
  XOR U15818 ( .A(n16040), .B(n15670), .Z(n16043) );
  XOR U15819 ( .A(n16044), .B(n16045), .Z(n15670) );
  AND U15820 ( .A(n518), .B(n16046), .Z(n16045) );
  XOR U15821 ( .A(n16047), .B(n16044), .Z(n16046) );
  XNOR U15822 ( .A(n15667), .B(n16040), .Z(n16042) );
  XOR U15823 ( .A(n16048), .B(n16049), .Z(n15667) );
  AND U15824 ( .A(n516), .B(n16050), .Z(n16049) );
  XOR U15825 ( .A(n16051), .B(n16048), .Z(n16050) );
  XOR U15826 ( .A(n16052), .B(n16053), .Z(n16040) );
  AND U15827 ( .A(n16054), .B(n16055), .Z(n16053) );
  XOR U15828 ( .A(n16052), .B(n15682), .Z(n16055) );
  XOR U15829 ( .A(n16056), .B(n16057), .Z(n15682) );
  AND U15830 ( .A(n518), .B(n16058), .Z(n16057) );
  XOR U15831 ( .A(n16059), .B(n16056), .Z(n16058) );
  XNOR U15832 ( .A(n15679), .B(n16052), .Z(n16054) );
  XOR U15833 ( .A(n16060), .B(n16061), .Z(n15679) );
  AND U15834 ( .A(n516), .B(n16062), .Z(n16061) );
  XOR U15835 ( .A(n16063), .B(n16060), .Z(n16062) );
  XOR U15836 ( .A(n16064), .B(n16065), .Z(n16052) );
  AND U15837 ( .A(n16066), .B(n16067), .Z(n16065) );
  XOR U15838 ( .A(n16064), .B(n15694), .Z(n16067) );
  XOR U15839 ( .A(n16068), .B(n16069), .Z(n15694) );
  AND U15840 ( .A(n518), .B(n16070), .Z(n16069) );
  XOR U15841 ( .A(n16071), .B(n16068), .Z(n16070) );
  XNOR U15842 ( .A(n15691), .B(n16064), .Z(n16066) );
  XOR U15843 ( .A(n16072), .B(n16073), .Z(n15691) );
  AND U15844 ( .A(n516), .B(n16074), .Z(n16073) );
  XOR U15845 ( .A(n16075), .B(n16072), .Z(n16074) );
  XOR U15846 ( .A(n16076), .B(n16077), .Z(n16064) );
  AND U15847 ( .A(n16078), .B(n16079), .Z(n16077) );
  XOR U15848 ( .A(n16076), .B(n15706), .Z(n16079) );
  XOR U15849 ( .A(n16080), .B(n16081), .Z(n15706) );
  AND U15850 ( .A(n518), .B(n16082), .Z(n16081) );
  XOR U15851 ( .A(n16083), .B(n16080), .Z(n16082) );
  XNOR U15852 ( .A(n15703), .B(n16076), .Z(n16078) );
  XOR U15853 ( .A(n16084), .B(n16085), .Z(n15703) );
  AND U15854 ( .A(n516), .B(n16086), .Z(n16085) );
  XOR U15855 ( .A(n16087), .B(n16084), .Z(n16086) );
  XOR U15856 ( .A(n16088), .B(n16089), .Z(n16076) );
  AND U15857 ( .A(n16090), .B(n16091), .Z(n16089) );
  XOR U15858 ( .A(n16088), .B(n15718), .Z(n16091) );
  XOR U15859 ( .A(n16092), .B(n16093), .Z(n15718) );
  AND U15860 ( .A(n518), .B(n16094), .Z(n16093) );
  XOR U15861 ( .A(n16095), .B(n16092), .Z(n16094) );
  XNOR U15862 ( .A(n15715), .B(n16088), .Z(n16090) );
  XOR U15863 ( .A(n16096), .B(n16097), .Z(n15715) );
  AND U15864 ( .A(n516), .B(n16098), .Z(n16097) );
  XOR U15865 ( .A(n16099), .B(n16096), .Z(n16098) );
  XOR U15866 ( .A(n16100), .B(n16101), .Z(n16088) );
  AND U15867 ( .A(n16102), .B(n16103), .Z(n16101) );
  XOR U15868 ( .A(n16100), .B(n15730), .Z(n16103) );
  XOR U15869 ( .A(n16104), .B(n16105), .Z(n15730) );
  AND U15870 ( .A(n518), .B(n16106), .Z(n16105) );
  XOR U15871 ( .A(n16107), .B(n16104), .Z(n16106) );
  XNOR U15872 ( .A(n15727), .B(n16100), .Z(n16102) );
  XOR U15873 ( .A(n16108), .B(n16109), .Z(n15727) );
  AND U15874 ( .A(n516), .B(n16110), .Z(n16109) );
  XOR U15875 ( .A(n16111), .B(n16108), .Z(n16110) );
  XOR U15876 ( .A(n16112), .B(n16113), .Z(n16100) );
  AND U15877 ( .A(n16114), .B(n16115), .Z(n16113) );
  XOR U15878 ( .A(n16112), .B(n15742), .Z(n16115) );
  XOR U15879 ( .A(n16116), .B(n16117), .Z(n15742) );
  AND U15880 ( .A(n518), .B(n16118), .Z(n16117) );
  XOR U15881 ( .A(n16119), .B(n16116), .Z(n16118) );
  XNOR U15882 ( .A(n15739), .B(n16112), .Z(n16114) );
  XOR U15883 ( .A(n16120), .B(n16121), .Z(n15739) );
  AND U15884 ( .A(n516), .B(n16122), .Z(n16121) );
  XOR U15885 ( .A(n16123), .B(n16120), .Z(n16122) );
  XOR U15886 ( .A(n16124), .B(n16125), .Z(n16112) );
  AND U15887 ( .A(n16126), .B(n16127), .Z(n16125) );
  XOR U15888 ( .A(n16124), .B(n15754), .Z(n16127) );
  XOR U15889 ( .A(n16128), .B(n16129), .Z(n15754) );
  AND U15890 ( .A(n518), .B(n16130), .Z(n16129) );
  XOR U15891 ( .A(n16131), .B(n16128), .Z(n16130) );
  XNOR U15892 ( .A(n15751), .B(n16124), .Z(n16126) );
  XOR U15893 ( .A(n16132), .B(n16133), .Z(n15751) );
  AND U15894 ( .A(n516), .B(n16134), .Z(n16133) );
  XOR U15895 ( .A(n16135), .B(n16132), .Z(n16134) );
  XOR U15896 ( .A(n16136), .B(n16137), .Z(n16124) );
  AND U15897 ( .A(n16138), .B(n16139), .Z(n16137) );
  XOR U15898 ( .A(n16136), .B(n15766), .Z(n16139) );
  XOR U15899 ( .A(n16140), .B(n16141), .Z(n15766) );
  AND U15900 ( .A(n518), .B(n16142), .Z(n16141) );
  XOR U15901 ( .A(n16143), .B(n16140), .Z(n16142) );
  XNOR U15902 ( .A(n15763), .B(n16136), .Z(n16138) );
  XOR U15903 ( .A(n16144), .B(n16145), .Z(n15763) );
  AND U15904 ( .A(n516), .B(n16146), .Z(n16145) );
  XOR U15905 ( .A(n16147), .B(n16144), .Z(n16146) );
  XOR U15906 ( .A(n16148), .B(n16149), .Z(n16136) );
  AND U15907 ( .A(n16150), .B(n16151), .Z(n16149) );
  XOR U15908 ( .A(n16148), .B(n15778), .Z(n16151) );
  XOR U15909 ( .A(n16152), .B(n16153), .Z(n15778) );
  AND U15910 ( .A(n518), .B(n16154), .Z(n16153) );
  XOR U15911 ( .A(n16155), .B(n16152), .Z(n16154) );
  XNOR U15912 ( .A(n15775), .B(n16148), .Z(n16150) );
  XOR U15913 ( .A(n16156), .B(n16157), .Z(n15775) );
  AND U15914 ( .A(n516), .B(n16158), .Z(n16157) );
  XOR U15915 ( .A(n16159), .B(n16156), .Z(n16158) );
  XOR U15916 ( .A(n16160), .B(n16161), .Z(n16148) );
  AND U15917 ( .A(n16162), .B(n16163), .Z(n16161) );
  XOR U15918 ( .A(n16160), .B(n15790), .Z(n16163) );
  XOR U15919 ( .A(n16164), .B(n16165), .Z(n15790) );
  AND U15920 ( .A(n518), .B(n16166), .Z(n16165) );
  XOR U15921 ( .A(n16167), .B(n16164), .Z(n16166) );
  XNOR U15922 ( .A(n15787), .B(n16160), .Z(n16162) );
  XOR U15923 ( .A(n16168), .B(n16169), .Z(n15787) );
  AND U15924 ( .A(n516), .B(n16170), .Z(n16169) );
  XOR U15925 ( .A(n16171), .B(n16168), .Z(n16170) );
  XOR U15926 ( .A(n16172), .B(n16173), .Z(n16160) );
  AND U15927 ( .A(n16174), .B(n16175), .Z(n16173) );
  XOR U15928 ( .A(n16172), .B(n15802), .Z(n16175) );
  XOR U15929 ( .A(n16176), .B(n16177), .Z(n15802) );
  AND U15930 ( .A(n518), .B(n16178), .Z(n16177) );
  XOR U15931 ( .A(n16179), .B(n16176), .Z(n16178) );
  XNOR U15932 ( .A(n15799), .B(n16172), .Z(n16174) );
  XOR U15933 ( .A(n16180), .B(n16181), .Z(n15799) );
  AND U15934 ( .A(n516), .B(n16182), .Z(n16181) );
  XOR U15935 ( .A(n16183), .B(n16180), .Z(n16182) );
  XOR U15936 ( .A(n16184), .B(n16185), .Z(n16172) );
  AND U15937 ( .A(n16186), .B(n16187), .Z(n16185) );
  XOR U15938 ( .A(n16184), .B(n15814), .Z(n16187) );
  XOR U15939 ( .A(n16188), .B(n16189), .Z(n15814) );
  AND U15940 ( .A(n518), .B(n16190), .Z(n16189) );
  XOR U15941 ( .A(n16191), .B(n16188), .Z(n16190) );
  XNOR U15942 ( .A(n15811), .B(n16184), .Z(n16186) );
  XOR U15943 ( .A(n16192), .B(n16193), .Z(n15811) );
  AND U15944 ( .A(n516), .B(n16194), .Z(n16193) );
  XOR U15945 ( .A(n16195), .B(n16192), .Z(n16194) );
  XOR U15946 ( .A(n16196), .B(n16197), .Z(n16184) );
  AND U15947 ( .A(n16198), .B(n16199), .Z(n16197) );
  XOR U15948 ( .A(n16196), .B(n15826), .Z(n16199) );
  XOR U15949 ( .A(n16200), .B(n16201), .Z(n15826) );
  AND U15950 ( .A(n518), .B(n16202), .Z(n16201) );
  XOR U15951 ( .A(n16203), .B(n16200), .Z(n16202) );
  XNOR U15952 ( .A(n15823), .B(n16196), .Z(n16198) );
  XOR U15953 ( .A(n16204), .B(n16205), .Z(n15823) );
  AND U15954 ( .A(n516), .B(n16206), .Z(n16205) );
  XOR U15955 ( .A(n16207), .B(n16204), .Z(n16206) );
  XOR U15956 ( .A(n16208), .B(n16209), .Z(n16196) );
  AND U15957 ( .A(n16210), .B(n16211), .Z(n16209) );
  XOR U15958 ( .A(n16208), .B(n15838), .Z(n16211) );
  XOR U15959 ( .A(n16212), .B(n16213), .Z(n15838) );
  AND U15960 ( .A(n518), .B(n16214), .Z(n16213) );
  XOR U15961 ( .A(n16215), .B(n16212), .Z(n16214) );
  XNOR U15962 ( .A(n15835), .B(n16208), .Z(n16210) );
  XOR U15963 ( .A(n16216), .B(n16217), .Z(n15835) );
  AND U15964 ( .A(n516), .B(n16218), .Z(n16217) );
  XOR U15965 ( .A(n16219), .B(n16216), .Z(n16218) );
  XOR U15966 ( .A(n16220), .B(n16221), .Z(n16208) );
  AND U15967 ( .A(n16222), .B(n16223), .Z(n16221) );
  XOR U15968 ( .A(n16220), .B(n15850), .Z(n16223) );
  XOR U15969 ( .A(n16224), .B(n16225), .Z(n15850) );
  AND U15970 ( .A(n518), .B(n16226), .Z(n16225) );
  XOR U15971 ( .A(n16227), .B(n16224), .Z(n16226) );
  XNOR U15972 ( .A(n15847), .B(n16220), .Z(n16222) );
  XOR U15973 ( .A(n16228), .B(n16229), .Z(n15847) );
  AND U15974 ( .A(n516), .B(n16230), .Z(n16229) );
  XOR U15975 ( .A(n16231), .B(n16228), .Z(n16230) );
  XOR U15976 ( .A(n16232), .B(n16233), .Z(n16220) );
  AND U15977 ( .A(n16234), .B(n16235), .Z(n16233) );
  XOR U15978 ( .A(n16232), .B(n15862), .Z(n16235) );
  XOR U15979 ( .A(n16236), .B(n16237), .Z(n15862) );
  AND U15980 ( .A(n518), .B(n16238), .Z(n16237) );
  XOR U15981 ( .A(n16239), .B(n16236), .Z(n16238) );
  XNOR U15982 ( .A(n15859), .B(n16232), .Z(n16234) );
  XOR U15983 ( .A(n16240), .B(n16241), .Z(n15859) );
  AND U15984 ( .A(n516), .B(n16242), .Z(n16241) );
  XOR U15985 ( .A(n16243), .B(n16240), .Z(n16242) );
  XOR U15986 ( .A(n16244), .B(n16245), .Z(n16232) );
  AND U15987 ( .A(n16246), .B(n16247), .Z(n16245) );
  XOR U15988 ( .A(n16244), .B(n15874), .Z(n16247) );
  XOR U15989 ( .A(n16248), .B(n16249), .Z(n15874) );
  AND U15990 ( .A(n518), .B(n16250), .Z(n16249) );
  XOR U15991 ( .A(n16251), .B(n16248), .Z(n16250) );
  XNOR U15992 ( .A(n15871), .B(n16244), .Z(n16246) );
  XOR U15993 ( .A(n16252), .B(n16253), .Z(n15871) );
  AND U15994 ( .A(n516), .B(n16254), .Z(n16253) );
  XOR U15995 ( .A(n16255), .B(n16252), .Z(n16254) );
  XOR U15996 ( .A(n16256), .B(n16257), .Z(n16244) );
  AND U15997 ( .A(n16258), .B(n16259), .Z(n16257) );
  XOR U15998 ( .A(n16256), .B(n15886), .Z(n16259) );
  XOR U15999 ( .A(n16260), .B(n16261), .Z(n15886) );
  AND U16000 ( .A(n518), .B(n16262), .Z(n16261) );
  XOR U16001 ( .A(n16263), .B(n16260), .Z(n16262) );
  XNOR U16002 ( .A(n15883), .B(n16256), .Z(n16258) );
  XOR U16003 ( .A(n16264), .B(n16265), .Z(n15883) );
  AND U16004 ( .A(n516), .B(n16266), .Z(n16265) );
  XOR U16005 ( .A(n16267), .B(n16264), .Z(n16266) );
  XOR U16006 ( .A(n16268), .B(n16269), .Z(n16256) );
  AND U16007 ( .A(n16270), .B(n16271), .Z(n16269) );
  XOR U16008 ( .A(n16268), .B(n15898), .Z(n16271) );
  XOR U16009 ( .A(n16272), .B(n16273), .Z(n15898) );
  AND U16010 ( .A(n518), .B(n16274), .Z(n16273) );
  XOR U16011 ( .A(n16275), .B(n16272), .Z(n16274) );
  XNOR U16012 ( .A(n15895), .B(n16268), .Z(n16270) );
  XOR U16013 ( .A(n16276), .B(n16277), .Z(n15895) );
  AND U16014 ( .A(n516), .B(n16278), .Z(n16277) );
  XOR U16015 ( .A(n16279), .B(n16276), .Z(n16278) );
  XOR U16016 ( .A(n16280), .B(n16281), .Z(n16268) );
  AND U16017 ( .A(n16282), .B(n16283), .Z(n16281) );
  XOR U16018 ( .A(n16280), .B(n15910), .Z(n16283) );
  XOR U16019 ( .A(n16284), .B(n16285), .Z(n15910) );
  AND U16020 ( .A(n518), .B(n16286), .Z(n16285) );
  XOR U16021 ( .A(n16287), .B(n16284), .Z(n16286) );
  XNOR U16022 ( .A(n15907), .B(n16280), .Z(n16282) );
  XOR U16023 ( .A(n16288), .B(n16289), .Z(n15907) );
  AND U16024 ( .A(n516), .B(n16290), .Z(n16289) );
  XOR U16025 ( .A(n16291), .B(n16288), .Z(n16290) );
  XOR U16026 ( .A(n16292), .B(n16293), .Z(n16280) );
  AND U16027 ( .A(n16294), .B(n16295), .Z(n16293) );
  XOR U16028 ( .A(n16292), .B(n15922), .Z(n16295) );
  XOR U16029 ( .A(n16296), .B(n16297), .Z(n15922) );
  AND U16030 ( .A(n518), .B(n16298), .Z(n16297) );
  XOR U16031 ( .A(n16299), .B(n16296), .Z(n16298) );
  XNOR U16032 ( .A(n15919), .B(n16292), .Z(n16294) );
  XOR U16033 ( .A(n16300), .B(n16301), .Z(n15919) );
  AND U16034 ( .A(n516), .B(n16302), .Z(n16301) );
  XOR U16035 ( .A(n16303), .B(n16300), .Z(n16302) );
  XOR U16036 ( .A(n16304), .B(n16305), .Z(n16292) );
  AND U16037 ( .A(n16306), .B(n16307), .Z(n16305) );
  XOR U16038 ( .A(n16304), .B(n15934), .Z(n16307) );
  XOR U16039 ( .A(n16308), .B(n16309), .Z(n15934) );
  AND U16040 ( .A(n518), .B(n16310), .Z(n16309) );
  XOR U16041 ( .A(n16311), .B(n16308), .Z(n16310) );
  XNOR U16042 ( .A(n15931), .B(n16304), .Z(n16306) );
  XOR U16043 ( .A(n16312), .B(n16313), .Z(n15931) );
  AND U16044 ( .A(n516), .B(n16314), .Z(n16313) );
  XOR U16045 ( .A(n16315), .B(n16312), .Z(n16314) );
  XOR U16046 ( .A(n16316), .B(n16317), .Z(n16304) );
  AND U16047 ( .A(n16318), .B(n16319), .Z(n16317) );
  XOR U16048 ( .A(n15946), .B(n16316), .Z(n16319) );
  XOR U16049 ( .A(n16320), .B(n16321), .Z(n15946) );
  AND U16050 ( .A(n518), .B(n16322), .Z(n16321) );
  XOR U16051 ( .A(n16320), .B(n16323), .Z(n16322) );
  XNOR U16052 ( .A(n16316), .B(n15943), .Z(n16318) );
  XOR U16053 ( .A(n16324), .B(n16325), .Z(n15943) );
  AND U16054 ( .A(n516), .B(n16326), .Z(n16325) );
  XOR U16055 ( .A(n16324), .B(n16327), .Z(n16326) );
  XOR U16056 ( .A(n16328), .B(n16329), .Z(n16316) );
  AND U16057 ( .A(n16330), .B(n16331), .Z(n16329) );
  XNOR U16058 ( .A(n16332), .B(n15959), .Z(n16331) );
  XOR U16059 ( .A(n16333), .B(n16334), .Z(n15959) );
  AND U16060 ( .A(n518), .B(n16335), .Z(n16334) );
  XOR U16061 ( .A(n16336), .B(n16333), .Z(n16335) );
  XNOR U16062 ( .A(n15956), .B(n16328), .Z(n16330) );
  XOR U16063 ( .A(n16337), .B(n16338), .Z(n15956) );
  AND U16064 ( .A(n516), .B(n16339), .Z(n16338) );
  XOR U16065 ( .A(n16340), .B(n16337), .Z(n16339) );
  IV U16066 ( .A(n16332), .Z(n16328) );
  AND U16067 ( .A(n15964), .B(n15967), .Z(n16332) );
  XNOR U16068 ( .A(n16341), .B(n16342), .Z(n15967) );
  AND U16069 ( .A(n518), .B(n16343), .Z(n16342) );
  XNOR U16070 ( .A(n16344), .B(n16341), .Z(n16343) );
  XOR U16071 ( .A(n16345), .B(n16346), .Z(n518) );
  AND U16072 ( .A(n16347), .B(n16348), .Z(n16346) );
  XOR U16073 ( .A(n16345), .B(n15975), .Z(n16348) );
  XNOR U16074 ( .A(n16349), .B(n16350), .Z(n15975) );
  AND U16075 ( .A(n16351), .B(n366), .Z(n16350) );
  AND U16076 ( .A(n16349), .B(n16352), .Z(n16351) );
  XNOR U16077 ( .A(n15972), .B(n16345), .Z(n16347) );
  XOR U16078 ( .A(n16353), .B(n16354), .Z(n15972) );
  AND U16079 ( .A(n16355), .B(n364), .Z(n16354) );
  NOR U16080 ( .A(n16353), .B(n16356), .Z(n16355) );
  XOR U16081 ( .A(n16357), .B(n16358), .Z(n16345) );
  AND U16082 ( .A(n16359), .B(n16360), .Z(n16358) );
  XOR U16083 ( .A(n16357), .B(n15987), .Z(n16360) );
  XOR U16084 ( .A(n16361), .B(n16362), .Z(n15987) );
  AND U16085 ( .A(n366), .B(n16363), .Z(n16362) );
  XOR U16086 ( .A(n16364), .B(n16361), .Z(n16363) );
  XNOR U16087 ( .A(n15984), .B(n16357), .Z(n16359) );
  XOR U16088 ( .A(n16365), .B(n16366), .Z(n15984) );
  AND U16089 ( .A(n364), .B(n16367), .Z(n16366) );
  XOR U16090 ( .A(n16368), .B(n16365), .Z(n16367) );
  XOR U16091 ( .A(n16369), .B(n16370), .Z(n16357) );
  AND U16092 ( .A(n16371), .B(n16372), .Z(n16370) );
  XOR U16093 ( .A(n16369), .B(n15999), .Z(n16372) );
  XOR U16094 ( .A(n16373), .B(n16374), .Z(n15999) );
  AND U16095 ( .A(n366), .B(n16375), .Z(n16374) );
  XOR U16096 ( .A(n16376), .B(n16373), .Z(n16375) );
  XNOR U16097 ( .A(n15996), .B(n16369), .Z(n16371) );
  XOR U16098 ( .A(n16377), .B(n16378), .Z(n15996) );
  AND U16099 ( .A(n364), .B(n16379), .Z(n16378) );
  XOR U16100 ( .A(n16380), .B(n16377), .Z(n16379) );
  XOR U16101 ( .A(n16381), .B(n16382), .Z(n16369) );
  AND U16102 ( .A(n16383), .B(n16384), .Z(n16382) );
  XOR U16103 ( .A(n16381), .B(n16011), .Z(n16384) );
  XOR U16104 ( .A(n16385), .B(n16386), .Z(n16011) );
  AND U16105 ( .A(n366), .B(n16387), .Z(n16386) );
  XOR U16106 ( .A(n16388), .B(n16385), .Z(n16387) );
  XNOR U16107 ( .A(n16008), .B(n16381), .Z(n16383) );
  XOR U16108 ( .A(n16389), .B(n16390), .Z(n16008) );
  AND U16109 ( .A(n364), .B(n16391), .Z(n16390) );
  XOR U16110 ( .A(n16392), .B(n16389), .Z(n16391) );
  XOR U16111 ( .A(n16393), .B(n16394), .Z(n16381) );
  AND U16112 ( .A(n16395), .B(n16396), .Z(n16394) );
  XOR U16113 ( .A(n16393), .B(n16023), .Z(n16396) );
  XOR U16114 ( .A(n16397), .B(n16398), .Z(n16023) );
  AND U16115 ( .A(n366), .B(n16399), .Z(n16398) );
  XOR U16116 ( .A(n16400), .B(n16397), .Z(n16399) );
  XNOR U16117 ( .A(n16020), .B(n16393), .Z(n16395) );
  XOR U16118 ( .A(n16401), .B(n16402), .Z(n16020) );
  AND U16119 ( .A(n364), .B(n16403), .Z(n16402) );
  XOR U16120 ( .A(n16404), .B(n16401), .Z(n16403) );
  XOR U16121 ( .A(n16405), .B(n16406), .Z(n16393) );
  AND U16122 ( .A(n16407), .B(n16408), .Z(n16406) );
  XOR U16123 ( .A(n16405), .B(n16035), .Z(n16408) );
  XOR U16124 ( .A(n16409), .B(n16410), .Z(n16035) );
  AND U16125 ( .A(n366), .B(n16411), .Z(n16410) );
  XOR U16126 ( .A(n16412), .B(n16409), .Z(n16411) );
  XNOR U16127 ( .A(n16032), .B(n16405), .Z(n16407) );
  XOR U16128 ( .A(n16413), .B(n16414), .Z(n16032) );
  AND U16129 ( .A(n364), .B(n16415), .Z(n16414) );
  XOR U16130 ( .A(n16416), .B(n16413), .Z(n16415) );
  XOR U16131 ( .A(n16417), .B(n16418), .Z(n16405) );
  AND U16132 ( .A(n16419), .B(n16420), .Z(n16418) );
  XOR U16133 ( .A(n16417), .B(n16047), .Z(n16420) );
  XOR U16134 ( .A(n16421), .B(n16422), .Z(n16047) );
  AND U16135 ( .A(n366), .B(n16423), .Z(n16422) );
  XOR U16136 ( .A(n16424), .B(n16421), .Z(n16423) );
  XNOR U16137 ( .A(n16044), .B(n16417), .Z(n16419) );
  XOR U16138 ( .A(n16425), .B(n16426), .Z(n16044) );
  AND U16139 ( .A(n364), .B(n16427), .Z(n16426) );
  XOR U16140 ( .A(n16428), .B(n16425), .Z(n16427) );
  XOR U16141 ( .A(n16429), .B(n16430), .Z(n16417) );
  AND U16142 ( .A(n16431), .B(n16432), .Z(n16430) );
  XOR U16143 ( .A(n16429), .B(n16059), .Z(n16432) );
  XOR U16144 ( .A(n16433), .B(n16434), .Z(n16059) );
  AND U16145 ( .A(n366), .B(n16435), .Z(n16434) );
  XOR U16146 ( .A(n16436), .B(n16433), .Z(n16435) );
  XNOR U16147 ( .A(n16056), .B(n16429), .Z(n16431) );
  XOR U16148 ( .A(n16437), .B(n16438), .Z(n16056) );
  AND U16149 ( .A(n364), .B(n16439), .Z(n16438) );
  XOR U16150 ( .A(n16440), .B(n16437), .Z(n16439) );
  XOR U16151 ( .A(n16441), .B(n16442), .Z(n16429) );
  AND U16152 ( .A(n16443), .B(n16444), .Z(n16442) );
  XOR U16153 ( .A(n16441), .B(n16071), .Z(n16444) );
  XOR U16154 ( .A(n16445), .B(n16446), .Z(n16071) );
  AND U16155 ( .A(n366), .B(n16447), .Z(n16446) );
  XOR U16156 ( .A(n16448), .B(n16445), .Z(n16447) );
  XNOR U16157 ( .A(n16068), .B(n16441), .Z(n16443) );
  XOR U16158 ( .A(n16449), .B(n16450), .Z(n16068) );
  AND U16159 ( .A(n364), .B(n16451), .Z(n16450) );
  XOR U16160 ( .A(n16452), .B(n16449), .Z(n16451) );
  XOR U16161 ( .A(n16453), .B(n16454), .Z(n16441) );
  AND U16162 ( .A(n16455), .B(n16456), .Z(n16454) );
  XOR U16163 ( .A(n16453), .B(n16083), .Z(n16456) );
  XOR U16164 ( .A(n16457), .B(n16458), .Z(n16083) );
  AND U16165 ( .A(n366), .B(n16459), .Z(n16458) );
  XOR U16166 ( .A(n16460), .B(n16457), .Z(n16459) );
  XNOR U16167 ( .A(n16080), .B(n16453), .Z(n16455) );
  XOR U16168 ( .A(n16461), .B(n16462), .Z(n16080) );
  AND U16169 ( .A(n364), .B(n16463), .Z(n16462) );
  XOR U16170 ( .A(n16464), .B(n16461), .Z(n16463) );
  XOR U16171 ( .A(n16465), .B(n16466), .Z(n16453) );
  AND U16172 ( .A(n16467), .B(n16468), .Z(n16466) );
  XOR U16173 ( .A(n16465), .B(n16095), .Z(n16468) );
  XOR U16174 ( .A(n16469), .B(n16470), .Z(n16095) );
  AND U16175 ( .A(n366), .B(n16471), .Z(n16470) );
  XOR U16176 ( .A(n16472), .B(n16469), .Z(n16471) );
  XNOR U16177 ( .A(n16092), .B(n16465), .Z(n16467) );
  XOR U16178 ( .A(n16473), .B(n16474), .Z(n16092) );
  AND U16179 ( .A(n364), .B(n16475), .Z(n16474) );
  XOR U16180 ( .A(n16476), .B(n16473), .Z(n16475) );
  XOR U16181 ( .A(n16477), .B(n16478), .Z(n16465) );
  AND U16182 ( .A(n16479), .B(n16480), .Z(n16478) );
  XOR U16183 ( .A(n16477), .B(n16107), .Z(n16480) );
  XOR U16184 ( .A(n16481), .B(n16482), .Z(n16107) );
  AND U16185 ( .A(n366), .B(n16483), .Z(n16482) );
  XOR U16186 ( .A(n16484), .B(n16481), .Z(n16483) );
  XNOR U16187 ( .A(n16104), .B(n16477), .Z(n16479) );
  XOR U16188 ( .A(n16485), .B(n16486), .Z(n16104) );
  AND U16189 ( .A(n364), .B(n16487), .Z(n16486) );
  XOR U16190 ( .A(n16488), .B(n16485), .Z(n16487) );
  XOR U16191 ( .A(n16489), .B(n16490), .Z(n16477) );
  AND U16192 ( .A(n16491), .B(n16492), .Z(n16490) );
  XOR U16193 ( .A(n16489), .B(n16119), .Z(n16492) );
  XOR U16194 ( .A(n16493), .B(n16494), .Z(n16119) );
  AND U16195 ( .A(n366), .B(n16495), .Z(n16494) );
  XOR U16196 ( .A(n16496), .B(n16493), .Z(n16495) );
  XNOR U16197 ( .A(n16116), .B(n16489), .Z(n16491) );
  XOR U16198 ( .A(n16497), .B(n16498), .Z(n16116) );
  AND U16199 ( .A(n364), .B(n16499), .Z(n16498) );
  XOR U16200 ( .A(n16500), .B(n16497), .Z(n16499) );
  XOR U16201 ( .A(n16501), .B(n16502), .Z(n16489) );
  AND U16202 ( .A(n16503), .B(n16504), .Z(n16502) );
  XOR U16203 ( .A(n16501), .B(n16131), .Z(n16504) );
  XOR U16204 ( .A(n16505), .B(n16506), .Z(n16131) );
  AND U16205 ( .A(n366), .B(n16507), .Z(n16506) );
  XOR U16206 ( .A(n16508), .B(n16505), .Z(n16507) );
  XNOR U16207 ( .A(n16128), .B(n16501), .Z(n16503) );
  XOR U16208 ( .A(n16509), .B(n16510), .Z(n16128) );
  AND U16209 ( .A(n364), .B(n16511), .Z(n16510) );
  XOR U16210 ( .A(n16512), .B(n16509), .Z(n16511) );
  XOR U16211 ( .A(n16513), .B(n16514), .Z(n16501) );
  AND U16212 ( .A(n16515), .B(n16516), .Z(n16514) );
  XOR U16213 ( .A(n16513), .B(n16143), .Z(n16516) );
  XOR U16214 ( .A(n16517), .B(n16518), .Z(n16143) );
  AND U16215 ( .A(n366), .B(n16519), .Z(n16518) );
  XOR U16216 ( .A(n16520), .B(n16517), .Z(n16519) );
  XNOR U16217 ( .A(n16140), .B(n16513), .Z(n16515) );
  XOR U16218 ( .A(n16521), .B(n16522), .Z(n16140) );
  AND U16219 ( .A(n364), .B(n16523), .Z(n16522) );
  XOR U16220 ( .A(n16524), .B(n16521), .Z(n16523) );
  XOR U16221 ( .A(n16525), .B(n16526), .Z(n16513) );
  AND U16222 ( .A(n16527), .B(n16528), .Z(n16526) );
  XOR U16223 ( .A(n16525), .B(n16155), .Z(n16528) );
  XOR U16224 ( .A(n16529), .B(n16530), .Z(n16155) );
  AND U16225 ( .A(n366), .B(n16531), .Z(n16530) );
  XOR U16226 ( .A(n16532), .B(n16529), .Z(n16531) );
  XNOR U16227 ( .A(n16152), .B(n16525), .Z(n16527) );
  XOR U16228 ( .A(n16533), .B(n16534), .Z(n16152) );
  AND U16229 ( .A(n364), .B(n16535), .Z(n16534) );
  XOR U16230 ( .A(n16536), .B(n16533), .Z(n16535) );
  XOR U16231 ( .A(n16537), .B(n16538), .Z(n16525) );
  AND U16232 ( .A(n16539), .B(n16540), .Z(n16538) );
  XOR U16233 ( .A(n16537), .B(n16167), .Z(n16540) );
  XOR U16234 ( .A(n16541), .B(n16542), .Z(n16167) );
  AND U16235 ( .A(n366), .B(n16543), .Z(n16542) );
  XOR U16236 ( .A(n16544), .B(n16541), .Z(n16543) );
  XNOR U16237 ( .A(n16164), .B(n16537), .Z(n16539) );
  XOR U16238 ( .A(n16545), .B(n16546), .Z(n16164) );
  AND U16239 ( .A(n364), .B(n16547), .Z(n16546) );
  XOR U16240 ( .A(n16548), .B(n16545), .Z(n16547) );
  XOR U16241 ( .A(n16549), .B(n16550), .Z(n16537) );
  AND U16242 ( .A(n16551), .B(n16552), .Z(n16550) );
  XOR U16243 ( .A(n16549), .B(n16179), .Z(n16552) );
  XOR U16244 ( .A(n16553), .B(n16554), .Z(n16179) );
  AND U16245 ( .A(n366), .B(n16555), .Z(n16554) );
  XOR U16246 ( .A(n16556), .B(n16553), .Z(n16555) );
  XNOR U16247 ( .A(n16176), .B(n16549), .Z(n16551) );
  XOR U16248 ( .A(n16557), .B(n16558), .Z(n16176) );
  AND U16249 ( .A(n364), .B(n16559), .Z(n16558) );
  XOR U16250 ( .A(n16560), .B(n16557), .Z(n16559) );
  XOR U16251 ( .A(n16561), .B(n16562), .Z(n16549) );
  AND U16252 ( .A(n16563), .B(n16564), .Z(n16562) );
  XOR U16253 ( .A(n16561), .B(n16191), .Z(n16564) );
  XOR U16254 ( .A(n16565), .B(n16566), .Z(n16191) );
  AND U16255 ( .A(n366), .B(n16567), .Z(n16566) );
  XOR U16256 ( .A(n16568), .B(n16565), .Z(n16567) );
  XNOR U16257 ( .A(n16188), .B(n16561), .Z(n16563) );
  XOR U16258 ( .A(n16569), .B(n16570), .Z(n16188) );
  AND U16259 ( .A(n364), .B(n16571), .Z(n16570) );
  XOR U16260 ( .A(n16572), .B(n16569), .Z(n16571) );
  XOR U16261 ( .A(n16573), .B(n16574), .Z(n16561) );
  AND U16262 ( .A(n16575), .B(n16576), .Z(n16574) );
  XOR U16263 ( .A(n16573), .B(n16203), .Z(n16576) );
  XOR U16264 ( .A(n16577), .B(n16578), .Z(n16203) );
  AND U16265 ( .A(n366), .B(n16579), .Z(n16578) );
  XOR U16266 ( .A(n16580), .B(n16577), .Z(n16579) );
  XNOR U16267 ( .A(n16200), .B(n16573), .Z(n16575) );
  XOR U16268 ( .A(n16581), .B(n16582), .Z(n16200) );
  AND U16269 ( .A(n364), .B(n16583), .Z(n16582) );
  XOR U16270 ( .A(n16584), .B(n16581), .Z(n16583) );
  XOR U16271 ( .A(n16585), .B(n16586), .Z(n16573) );
  AND U16272 ( .A(n16587), .B(n16588), .Z(n16586) );
  XOR U16273 ( .A(n16585), .B(n16215), .Z(n16588) );
  XOR U16274 ( .A(n16589), .B(n16590), .Z(n16215) );
  AND U16275 ( .A(n366), .B(n16591), .Z(n16590) );
  XOR U16276 ( .A(n16592), .B(n16589), .Z(n16591) );
  XNOR U16277 ( .A(n16212), .B(n16585), .Z(n16587) );
  XOR U16278 ( .A(n16593), .B(n16594), .Z(n16212) );
  AND U16279 ( .A(n364), .B(n16595), .Z(n16594) );
  XOR U16280 ( .A(n16596), .B(n16593), .Z(n16595) );
  XOR U16281 ( .A(n16597), .B(n16598), .Z(n16585) );
  AND U16282 ( .A(n16599), .B(n16600), .Z(n16598) );
  XOR U16283 ( .A(n16597), .B(n16227), .Z(n16600) );
  XOR U16284 ( .A(n16601), .B(n16602), .Z(n16227) );
  AND U16285 ( .A(n366), .B(n16603), .Z(n16602) );
  XOR U16286 ( .A(n16604), .B(n16601), .Z(n16603) );
  XNOR U16287 ( .A(n16224), .B(n16597), .Z(n16599) );
  XOR U16288 ( .A(n16605), .B(n16606), .Z(n16224) );
  AND U16289 ( .A(n364), .B(n16607), .Z(n16606) );
  XOR U16290 ( .A(n16608), .B(n16605), .Z(n16607) );
  XOR U16291 ( .A(n16609), .B(n16610), .Z(n16597) );
  AND U16292 ( .A(n16611), .B(n16612), .Z(n16610) );
  XOR U16293 ( .A(n16609), .B(n16239), .Z(n16612) );
  XOR U16294 ( .A(n16613), .B(n16614), .Z(n16239) );
  AND U16295 ( .A(n366), .B(n16615), .Z(n16614) );
  XOR U16296 ( .A(n16616), .B(n16613), .Z(n16615) );
  XNOR U16297 ( .A(n16236), .B(n16609), .Z(n16611) );
  XOR U16298 ( .A(n16617), .B(n16618), .Z(n16236) );
  AND U16299 ( .A(n364), .B(n16619), .Z(n16618) );
  XOR U16300 ( .A(n16620), .B(n16617), .Z(n16619) );
  XOR U16301 ( .A(n16621), .B(n16622), .Z(n16609) );
  AND U16302 ( .A(n16623), .B(n16624), .Z(n16622) );
  XOR U16303 ( .A(n16621), .B(n16251), .Z(n16624) );
  XOR U16304 ( .A(n16625), .B(n16626), .Z(n16251) );
  AND U16305 ( .A(n366), .B(n16627), .Z(n16626) );
  XOR U16306 ( .A(n16628), .B(n16625), .Z(n16627) );
  XNOR U16307 ( .A(n16248), .B(n16621), .Z(n16623) );
  XOR U16308 ( .A(n16629), .B(n16630), .Z(n16248) );
  AND U16309 ( .A(n364), .B(n16631), .Z(n16630) );
  XOR U16310 ( .A(n16632), .B(n16629), .Z(n16631) );
  XOR U16311 ( .A(n16633), .B(n16634), .Z(n16621) );
  AND U16312 ( .A(n16635), .B(n16636), .Z(n16634) );
  XOR U16313 ( .A(n16633), .B(n16263), .Z(n16636) );
  XOR U16314 ( .A(n16637), .B(n16638), .Z(n16263) );
  AND U16315 ( .A(n366), .B(n16639), .Z(n16638) );
  XOR U16316 ( .A(n16640), .B(n16637), .Z(n16639) );
  XNOR U16317 ( .A(n16260), .B(n16633), .Z(n16635) );
  XOR U16318 ( .A(n16641), .B(n16642), .Z(n16260) );
  AND U16319 ( .A(n364), .B(n16643), .Z(n16642) );
  XOR U16320 ( .A(n16644), .B(n16641), .Z(n16643) );
  XOR U16321 ( .A(n16645), .B(n16646), .Z(n16633) );
  AND U16322 ( .A(n16647), .B(n16648), .Z(n16646) );
  XOR U16323 ( .A(n16645), .B(n16275), .Z(n16648) );
  XOR U16324 ( .A(n16649), .B(n16650), .Z(n16275) );
  AND U16325 ( .A(n366), .B(n16651), .Z(n16650) );
  XOR U16326 ( .A(n16652), .B(n16649), .Z(n16651) );
  XNOR U16327 ( .A(n16272), .B(n16645), .Z(n16647) );
  XOR U16328 ( .A(n16653), .B(n16654), .Z(n16272) );
  AND U16329 ( .A(n364), .B(n16655), .Z(n16654) );
  XOR U16330 ( .A(n16656), .B(n16653), .Z(n16655) );
  XOR U16331 ( .A(n16657), .B(n16658), .Z(n16645) );
  AND U16332 ( .A(n16659), .B(n16660), .Z(n16658) );
  XOR U16333 ( .A(n16657), .B(n16287), .Z(n16660) );
  XOR U16334 ( .A(n16661), .B(n16662), .Z(n16287) );
  AND U16335 ( .A(n366), .B(n16663), .Z(n16662) );
  XOR U16336 ( .A(n16664), .B(n16661), .Z(n16663) );
  XNOR U16337 ( .A(n16284), .B(n16657), .Z(n16659) );
  XOR U16338 ( .A(n16665), .B(n16666), .Z(n16284) );
  AND U16339 ( .A(n364), .B(n16667), .Z(n16666) );
  XOR U16340 ( .A(n16668), .B(n16665), .Z(n16667) );
  XOR U16341 ( .A(n16669), .B(n16670), .Z(n16657) );
  AND U16342 ( .A(n16671), .B(n16672), .Z(n16670) );
  XOR U16343 ( .A(n16669), .B(n16299), .Z(n16672) );
  XOR U16344 ( .A(n16673), .B(n16674), .Z(n16299) );
  AND U16345 ( .A(n366), .B(n16675), .Z(n16674) );
  XOR U16346 ( .A(n16676), .B(n16673), .Z(n16675) );
  XNOR U16347 ( .A(n16296), .B(n16669), .Z(n16671) );
  XOR U16348 ( .A(n16677), .B(n16678), .Z(n16296) );
  AND U16349 ( .A(n364), .B(n16679), .Z(n16678) );
  XOR U16350 ( .A(n16680), .B(n16677), .Z(n16679) );
  XOR U16351 ( .A(n16681), .B(n16682), .Z(n16669) );
  AND U16352 ( .A(n16683), .B(n16684), .Z(n16682) );
  XOR U16353 ( .A(n16681), .B(n16311), .Z(n16684) );
  XOR U16354 ( .A(n16685), .B(n16686), .Z(n16311) );
  AND U16355 ( .A(n366), .B(n16687), .Z(n16686) );
  XOR U16356 ( .A(n16688), .B(n16685), .Z(n16687) );
  XNOR U16357 ( .A(n16308), .B(n16681), .Z(n16683) );
  XOR U16358 ( .A(n16689), .B(n16690), .Z(n16308) );
  AND U16359 ( .A(n364), .B(n16691), .Z(n16690) );
  XOR U16360 ( .A(n16692), .B(n16689), .Z(n16691) );
  XOR U16361 ( .A(n16693), .B(n16694), .Z(n16681) );
  AND U16362 ( .A(n16695), .B(n16696), .Z(n16694) );
  XOR U16363 ( .A(n16323), .B(n16693), .Z(n16696) );
  XOR U16364 ( .A(n16697), .B(n16698), .Z(n16323) );
  AND U16365 ( .A(n366), .B(n16699), .Z(n16698) );
  XOR U16366 ( .A(n16697), .B(n16700), .Z(n16699) );
  XNOR U16367 ( .A(n16693), .B(n16320), .Z(n16695) );
  XOR U16368 ( .A(n16701), .B(n16702), .Z(n16320) );
  AND U16369 ( .A(n364), .B(n16703), .Z(n16702) );
  XOR U16370 ( .A(n16701), .B(n16704), .Z(n16703) );
  XOR U16371 ( .A(n16705), .B(n16706), .Z(n16693) );
  AND U16372 ( .A(n16707), .B(n16708), .Z(n16706) );
  XNOR U16373 ( .A(n16709), .B(n16336), .Z(n16708) );
  XOR U16374 ( .A(n16710), .B(n16711), .Z(n16336) );
  AND U16375 ( .A(n366), .B(n16712), .Z(n16711) );
  XOR U16376 ( .A(n16713), .B(n16710), .Z(n16712) );
  XNOR U16377 ( .A(n16333), .B(n16705), .Z(n16707) );
  XOR U16378 ( .A(n16714), .B(n16715), .Z(n16333) );
  AND U16379 ( .A(n364), .B(n16716), .Z(n16715) );
  XOR U16380 ( .A(n16717), .B(n16714), .Z(n16716) );
  IV U16381 ( .A(n16709), .Z(n16705) );
  AND U16382 ( .A(n16341), .B(n16344), .Z(n16709) );
  XNOR U16383 ( .A(n16718), .B(n16719), .Z(n16344) );
  AND U16384 ( .A(n366), .B(n16720), .Z(n16719) );
  XNOR U16385 ( .A(n16721), .B(n16718), .Z(n16720) );
  XOR U16386 ( .A(n16722), .B(n16723), .Z(n366) );
  AND U16387 ( .A(n16724), .B(n16725), .Z(n16723) );
  XOR U16388 ( .A(n16352), .B(n16722), .Z(n16725) );
  IV U16389 ( .A(n16726), .Z(n16352) );
  AND U16390 ( .A(p_input[2047]), .B(p_input[2015]), .Z(n16726) );
  XOR U16391 ( .A(n16722), .B(n16349), .Z(n16724) );
  AND U16392 ( .A(p_input[1951]), .B(p_input[1983]), .Z(n16349) );
  XOR U16393 ( .A(n16727), .B(n16728), .Z(n16722) );
  AND U16394 ( .A(n16729), .B(n16730), .Z(n16728) );
  XOR U16395 ( .A(n16727), .B(n16364), .Z(n16730) );
  XNOR U16396 ( .A(p_input[2014]), .B(n16731), .Z(n16364) );
  AND U16397 ( .A(n430), .B(n16732), .Z(n16731) );
  XOR U16398 ( .A(p_input[2046]), .B(p_input[2014]), .Z(n16732) );
  XNOR U16399 ( .A(n16361), .B(n16727), .Z(n16729) );
  XOR U16400 ( .A(n16733), .B(n16734), .Z(n16361) );
  AND U16401 ( .A(n428), .B(n16735), .Z(n16734) );
  XOR U16402 ( .A(p_input[1982]), .B(p_input[1950]), .Z(n16735) );
  XOR U16403 ( .A(n16736), .B(n16737), .Z(n16727) );
  AND U16404 ( .A(n16738), .B(n16739), .Z(n16737) );
  XOR U16405 ( .A(n16736), .B(n16376), .Z(n16739) );
  XNOR U16406 ( .A(p_input[2013]), .B(n16740), .Z(n16376) );
  AND U16407 ( .A(n430), .B(n16741), .Z(n16740) );
  XOR U16408 ( .A(p_input[2045]), .B(p_input[2013]), .Z(n16741) );
  XNOR U16409 ( .A(n16373), .B(n16736), .Z(n16738) );
  XOR U16410 ( .A(n16742), .B(n16743), .Z(n16373) );
  AND U16411 ( .A(n428), .B(n16744), .Z(n16743) );
  XOR U16412 ( .A(p_input[1981]), .B(p_input[1949]), .Z(n16744) );
  XOR U16413 ( .A(n16745), .B(n16746), .Z(n16736) );
  AND U16414 ( .A(n16747), .B(n16748), .Z(n16746) );
  XOR U16415 ( .A(n16745), .B(n16388), .Z(n16748) );
  XNOR U16416 ( .A(p_input[2012]), .B(n16749), .Z(n16388) );
  AND U16417 ( .A(n430), .B(n16750), .Z(n16749) );
  XOR U16418 ( .A(p_input[2044]), .B(p_input[2012]), .Z(n16750) );
  XNOR U16419 ( .A(n16385), .B(n16745), .Z(n16747) );
  XOR U16420 ( .A(n16751), .B(n16752), .Z(n16385) );
  AND U16421 ( .A(n428), .B(n16753), .Z(n16752) );
  XOR U16422 ( .A(p_input[1980]), .B(p_input[1948]), .Z(n16753) );
  XOR U16423 ( .A(n16754), .B(n16755), .Z(n16745) );
  AND U16424 ( .A(n16756), .B(n16757), .Z(n16755) );
  XOR U16425 ( .A(n16754), .B(n16400), .Z(n16757) );
  XNOR U16426 ( .A(p_input[2011]), .B(n16758), .Z(n16400) );
  AND U16427 ( .A(n430), .B(n16759), .Z(n16758) );
  XOR U16428 ( .A(p_input[2043]), .B(p_input[2011]), .Z(n16759) );
  XNOR U16429 ( .A(n16397), .B(n16754), .Z(n16756) );
  XOR U16430 ( .A(n16760), .B(n16761), .Z(n16397) );
  AND U16431 ( .A(n428), .B(n16762), .Z(n16761) );
  XOR U16432 ( .A(p_input[1979]), .B(p_input[1947]), .Z(n16762) );
  XOR U16433 ( .A(n16763), .B(n16764), .Z(n16754) );
  AND U16434 ( .A(n16765), .B(n16766), .Z(n16764) );
  XOR U16435 ( .A(n16763), .B(n16412), .Z(n16766) );
  XNOR U16436 ( .A(p_input[2010]), .B(n16767), .Z(n16412) );
  AND U16437 ( .A(n430), .B(n16768), .Z(n16767) );
  XOR U16438 ( .A(p_input[2042]), .B(p_input[2010]), .Z(n16768) );
  XNOR U16439 ( .A(n16409), .B(n16763), .Z(n16765) );
  XOR U16440 ( .A(n16769), .B(n16770), .Z(n16409) );
  AND U16441 ( .A(n428), .B(n16771), .Z(n16770) );
  XOR U16442 ( .A(p_input[1978]), .B(p_input[1946]), .Z(n16771) );
  XOR U16443 ( .A(n16772), .B(n16773), .Z(n16763) );
  AND U16444 ( .A(n16774), .B(n16775), .Z(n16773) );
  XOR U16445 ( .A(n16772), .B(n16424), .Z(n16775) );
  XNOR U16446 ( .A(p_input[2009]), .B(n16776), .Z(n16424) );
  AND U16447 ( .A(n430), .B(n16777), .Z(n16776) );
  XOR U16448 ( .A(p_input[2041]), .B(p_input[2009]), .Z(n16777) );
  XNOR U16449 ( .A(n16421), .B(n16772), .Z(n16774) );
  XOR U16450 ( .A(n16778), .B(n16779), .Z(n16421) );
  AND U16451 ( .A(n428), .B(n16780), .Z(n16779) );
  XOR U16452 ( .A(p_input[1977]), .B(p_input[1945]), .Z(n16780) );
  XOR U16453 ( .A(n16781), .B(n16782), .Z(n16772) );
  AND U16454 ( .A(n16783), .B(n16784), .Z(n16782) );
  XOR U16455 ( .A(n16781), .B(n16436), .Z(n16784) );
  XNOR U16456 ( .A(p_input[2008]), .B(n16785), .Z(n16436) );
  AND U16457 ( .A(n430), .B(n16786), .Z(n16785) );
  XOR U16458 ( .A(p_input[2040]), .B(p_input[2008]), .Z(n16786) );
  XNOR U16459 ( .A(n16433), .B(n16781), .Z(n16783) );
  XOR U16460 ( .A(n16787), .B(n16788), .Z(n16433) );
  AND U16461 ( .A(n428), .B(n16789), .Z(n16788) );
  XOR U16462 ( .A(p_input[1976]), .B(p_input[1944]), .Z(n16789) );
  XOR U16463 ( .A(n16790), .B(n16791), .Z(n16781) );
  AND U16464 ( .A(n16792), .B(n16793), .Z(n16791) );
  XOR U16465 ( .A(n16790), .B(n16448), .Z(n16793) );
  XNOR U16466 ( .A(p_input[2007]), .B(n16794), .Z(n16448) );
  AND U16467 ( .A(n430), .B(n16795), .Z(n16794) );
  XOR U16468 ( .A(p_input[2039]), .B(p_input[2007]), .Z(n16795) );
  XNOR U16469 ( .A(n16445), .B(n16790), .Z(n16792) );
  XOR U16470 ( .A(n16796), .B(n16797), .Z(n16445) );
  AND U16471 ( .A(n428), .B(n16798), .Z(n16797) );
  XOR U16472 ( .A(p_input[1975]), .B(p_input[1943]), .Z(n16798) );
  XOR U16473 ( .A(n16799), .B(n16800), .Z(n16790) );
  AND U16474 ( .A(n16801), .B(n16802), .Z(n16800) );
  XOR U16475 ( .A(n16799), .B(n16460), .Z(n16802) );
  XNOR U16476 ( .A(p_input[2006]), .B(n16803), .Z(n16460) );
  AND U16477 ( .A(n430), .B(n16804), .Z(n16803) );
  XOR U16478 ( .A(p_input[2038]), .B(p_input[2006]), .Z(n16804) );
  XNOR U16479 ( .A(n16457), .B(n16799), .Z(n16801) );
  XOR U16480 ( .A(n16805), .B(n16806), .Z(n16457) );
  AND U16481 ( .A(n428), .B(n16807), .Z(n16806) );
  XOR U16482 ( .A(p_input[1974]), .B(p_input[1942]), .Z(n16807) );
  XOR U16483 ( .A(n16808), .B(n16809), .Z(n16799) );
  AND U16484 ( .A(n16810), .B(n16811), .Z(n16809) );
  XOR U16485 ( .A(n16808), .B(n16472), .Z(n16811) );
  XNOR U16486 ( .A(p_input[2005]), .B(n16812), .Z(n16472) );
  AND U16487 ( .A(n430), .B(n16813), .Z(n16812) );
  XOR U16488 ( .A(p_input[2037]), .B(p_input[2005]), .Z(n16813) );
  XNOR U16489 ( .A(n16469), .B(n16808), .Z(n16810) );
  XOR U16490 ( .A(n16814), .B(n16815), .Z(n16469) );
  AND U16491 ( .A(n428), .B(n16816), .Z(n16815) );
  XOR U16492 ( .A(p_input[1973]), .B(p_input[1941]), .Z(n16816) );
  XOR U16493 ( .A(n16817), .B(n16818), .Z(n16808) );
  AND U16494 ( .A(n16819), .B(n16820), .Z(n16818) );
  XOR U16495 ( .A(n16817), .B(n16484), .Z(n16820) );
  XNOR U16496 ( .A(p_input[2004]), .B(n16821), .Z(n16484) );
  AND U16497 ( .A(n430), .B(n16822), .Z(n16821) );
  XOR U16498 ( .A(p_input[2036]), .B(p_input[2004]), .Z(n16822) );
  XNOR U16499 ( .A(n16481), .B(n16817), .Z(n16819) );
  XOR U16500 ( .A(n16823), .B(n16824), .Z(n16481) );
  AND U16501 ( .A(n428), .B(n16825), .Z(n16824) );
  XOR U16502 ( .A(p_input[1972]), .B(p_input[1940]), .Z(n16825) );
  XOR U16503 ( .A(n16826), .B(n16827), .Z(n16817) );
  AND U16504 ( .A(n16828), .B(n16829), .Z(n16827) );
  XOR U16505 ( .A(n16826), .B(n16496), .Z(n16829) );
  XNOR U16506 ( .A(p_input[2003]), .B(n16830), .Z(n16496) );
  AND U16507 ( .A(n430), .B(n16831), .Z(n16830) );
  XOR U16508 ( .A(p_input[2035]), .B(p_input[2003]), .Z(n16831) );
  XNOR U16509 ( .A(n16493), .B(n16826), .Z(n16828) );
  XOR U16510 ( .A(n16832), .B(n16833), .Z(n16493) );
  AND U16511 ( .A(n428), .B(n16834), .Z(n16833) );
  XOR U16512 ( .A(p_input[1971]), .B(p_input[1939]), .Z(n16834) );
  XOR U16513 ( .A(n16835), .B(n16836), .Z(n16826) );
  AND U16514 ( .A(n16837), .B(n16838), .Z(n16836) );
  XOR U16515 ( .A(n16835), .B(n16508), .Z(n16838) );
  XNOR U16516 ( .A(p_input[2002]), .B(n16839), .Z(n16508) );
  AND U16517 ( .A(n430), .B(n16840), .Z(n16839) );
  XOR U16518 ( .A(p_input[2034]), .B(p_input[2002]), .Z(n16840) );
  XNOR U16519 ( .A(n16505), .B(n16835), .Z(n16837) );
  XOR U16520 ( .A(n16841), .B(n16842), .Z(n16505) );
  AND U16521 ( .A(n428), .B(n16843), .Z(n16842) );
  XOR U16522 ( .A(p_input[1970]), .B(p_input[1938]), .Z(n16843) );
  XOR U16523 ( .A(n16844), .B(n16845), .Z(n16835) );
  AND U16524 ( .A(n16846), .B(n16847), .Z(n16845) );
  XOR U16525 ( .A(n16844), .B(n16520), .Z(n16847) );
  XNOR U16526 ( .A(p_input[2001]), .B(n16848), .Z(n16520) );
  AND U16527 ( .A(n430), .B(n16849), .Z(n16848) );
  XOR U16528 ( .A(p_input[2033]), .B(p_input[2001]), .Z(n16849) );
  XNOR U16529 ( .A(n16517), .B(n16844), .Z(n16846) );
  XOR U16530 ( .A(n16850), .B(n16851), .Z(n16517) );
  AND U16531 ( .A(n428), .B(n16852), .Z(n16851) );
  XOR U16532 ( .A(p_input[1969]), .B(p_input[1937]), .Z(n16852) );
  XOR U16533 ( .A(n16853), .B(n16854), .Z(n16844) );
  AND U16534 ( .A(n16855), .B(n16856), .Z(n16854) );
  XOR U16535 ( .A(n16853), .B(n16532), .Z(n16856) );
  XNOR U16536 ( .A(p_input[2000]), .B(n16857), .Z(n16532) );
  AND U16537 ( .A(n430), .B(n16858), .Z(n16857) );
  XOR U16538 ( .A(p_input[2032]), .B(p_input[2000]), .Z(n16858) );
  XNOR U16539 ( .A(n16529), .B(n16853), .Z(n16855) );
  XOR U16540 ( .A(n16859), .B(n16860), .Z(n16529) );
  AND U16541 ( .A(n428), .B(n16861), .Z(n16860) );
  XOR U16542 ( .A(p_input[1968]), .B(p_input[1936]), .Z(n16861) );
  XOR U16543 ( .A(n16862), .B(n16863), .Z(n16853) );
  AND U16544 ( .A(n16864), .B(n16865), .Z(n16863) );
  XOR U16545 ( .A(n16862), .B(n16544), .Z(n16865) );
  XNOR U16546 ( .A(p_input[1999]), .B(n16866), .Z(n16544) );
  AND U16547 ( .A(n430), .B(n16867), .Z(n16866) );
  XOR U16548 ( .A(p_input[2031]), .B(p_input[1999]), .Z(n16867) );
  XNOR U16549 ( .A(n16541), .B(n16862), .Z(n16864) );
  XOR U16550 ( .A(n16868), .B(n16869), .Z(n16541) );
  AND U16551 ( .A(n428), .B(n16870), .Z(n16869) );
  XOR U16552 ( .A(p_input[1967]), .B(p_input[1935]), .Z(n16870) );
  XOR U16553 ( .A(n16871), .B(n16872), .Z(n16862) );
  AND U16554 ( .A(n16873), .B(n16874), .Z(n16872) );
  XOR U16555 ( .A(n16871), .B(n16556), .Z(n16874) );
  XNOR U16556 ( .A(p_input[1998]), .B(n16875), .Z(n16556) );
  AND U16557 ( .A(n430), .B(n16876), .Z(n16875) );
  XOR U16558 ( .A(p_input[2030]), .B(p_input[1998]), .Z(n16876) );
  XNOR U16559 ( .A(n16553), .B(n16871), .Z(n16873) );
  XOR U16560 ( .A(n16877), .B(n16878), .Z(n16553) );
  AND U16561 ( .A(n428), .B(n16879), .Z(n16878) );
  XOR U16562 ( .A(p_input[1966]), .B(p_input[1934]), .Z(n16879) );
  XOR U16563 ( .A(n16880), .B(n16881), .Z(n16871) );
  AND U16564 ( .A(n16882), .B(n16883), .Z(n16881) );
  XOR U16565 ( .A(n16880), .B(n16568), .Z(n16883) );
  XNOR U16566 ( .A(p_input[1997]), .B(n16884), .Z(n16568) );
  AND U16567 ( .A(n430), .B(n16885), .Z(n16884) );
  XOR U16568 ( .A(p_input[2029]), .B(p_input[1997]), .Z(n16885) );
  XNOR U16569 ( .A(n16565), .B(n16880), .Z(n16882) );
  XOR U16570 ( .A(n16886), .B(n16887), .Z(n16565) );
  AND U16571 ( .A(n428), .B(n16888), .Z(n16887) );
  XOR U16572 ( .A(p_input[1965]), .B(p_input[1933]), .Z(n16888) );
  XOR U16573 ( .A(n16889), .B(n16890), .Z(n16880) );
  AND U16574 ( .A(n16891), .B(n16892), .Z(n16890) );
  XOR U16575 ( .A(n16889), .B(n16580), .Z(n16892) );
  XNOR U16576 ( .A(p_input[1996]), .B(n16893), .Z(n16580) );
  AND U16577 ( .A(n430), .B(n16894), .Z(n16893) );
  XOR U16578 ( .A(p_input[2028]), .B(p_input[1996]), .Z(n16894) );
  XNOR U16579 ( .A(n16577), .B(n16889), .Z(n16891) );
  XOR U16580 ( .A(n16895), .B(n16896), .Z(n16577) );
  AND U16581 ( .A(n428), .B(n16897), .Z(n16896) );
  XOR U16582 ( .A(p_input[1964]), .B(p_input[1932]), .Z(n16897) );
  XOR U16583 ( .A(n16898), .B(n16899), .Z(n16889) );
  AND U16584 ( .A(n16900), .B(n16901), .Z(n16899) );
  XOR U16585 ( .A(n16898), .B(n16592), .Z(n16901) );
  XNOR U16586 ( .A(p_input[1995]), .B(n16902), .Z(n16592) );
  AND U16587 ( .A(n430), .B(n16903), .Z(n16902) );
  XOR U16588 ( .A(p_input[2027]), .B(p_input[1995]), .Z(n16903) );
  XNOR U16589 ( .A(n16589), .B(n16898), .Z(n16900) );
  XOR U16590 ( .A(n16904), .B(n16905), .Z(n16589) );
  AND U16591 ( .A(n428), .B(n16906), .Z(n16905) );
  XOR U16592 ( .A(p_input[1963]), .B(p_input[1931]), .Z(n16906) );
  XOR U16593 ( .A(n16907), .B(n16908), .Z(n16898) );
  AND U16594 ( .A(n16909), .B(n16910), .Z(n16908) );
  XOR U16595 ( .A(n16907), .B(n16604), .Z(n16910) );
  XNOR U16596 ( .A(p_input[1994]), .B(n16911), .Z(n16604) );
  AND U16597 ( .A(n430), .B(n16912), .Z(n16911) );
  XOR U16598 ( .A(p_input[2026]), .B(p_input[1994]), .Z(n16912) );
  XNOR U16599 ( .A(n16601), .B(n16907), .Z(n16909) );
  XOR U16600 ( .A(n16913), .B(n16914), .Z(n16601) );
  AND U16601 ( .A(n428), .B(n16915), .Z(n16914) );
  XOR U16602 ( .A(p_input[1962]), .B(p_input[1930]), .Z(n16915) );
  XOR U16603 ( .A(n16916), .B(n16917), .Z(n16907) );
  AND U16604 ( .A(n16918), .B(n16919), .Z(n16917) );
  XOR U16605 ( .A(n16916), .B(n16616), .Z(n16919) );
  XNOR U16606 ( .A(p_input[1993]), .B(n16920), .Z(n16616) );
  AND U16607 ( .A(n430), .B(n16921), .Z(n16920) );
  XOR U16608 ( .A(p_input[2025]), .B(p_input[1993]), .Z(n16921) );
  XNOR U16609 ( .A(n16613), .B(n16916), .Z(n16918) );
  XOR U16610 ( .A(n16922), .B(n16923), .Z(n16613) );
  AND U16611 ( .A(n428), .B(n16924), .Z(n16923) );
  XOR U16612 ( .A(p_input[1961]), .B(p_input[1929]), .Z(n16924) );
  XOR U16613 ( .A(n16925), .B(n16926), .Z(n16916) );
  AND U16614 ( .A(n16927), .B(n16928), .Z(n16926) );
  XOR U16615 ( .A(n16925), .B(n16628), .Z(n16928) );
  XNOR U16616 ( .A(p_input[1992]), .B(n16929), .Z(n16628) );
  AND U16617 ( .A(n430), .B(n16930), .Z(n16929) );
  XOR U16618 ( .A(p_input[2024]), .B(p_input[1992]), .Z(n16930) );
  XNOR U16619 ( .A(n16625), .B(n16925), .Z(n16927) );
  XOR U16620 ( .A(n16931), .B(n16932), .Z(n16625) );
  AND U16621 ( .A(n428), .B(n16933), .Z(n16932) );
  XOR U16622 ( .A(p_input[1960]), .B(p_input[1928]), .Z(n16933) );
  XOR U16623 ( .A(n16934), .B(n16935), .Z(n16925) );
  AND U16624 ( .A(n16936), .B(n16937), .Z(n16935) );
  XOR U16625 ( .A(n16934), .B(n16640), .Z(n16937) );
  XNOR U16626 ( .A(p_input[1991]), .B(n16938), .Z(n16640) );
  AND U16627 ( .A(n430), .B(n16939), .Z(n16938) );
  XOR U16628 ( .A(p_input[2023]), .B(p_input[1991]), .Z(n16939) );
  XNOR U16629 ( .A(n16637), .B(n16934), .Z(n16936) );
  XOR U16630 ( .A(n16940), .B(n16941), .Z(n16637) );
  AND U16631 ( .A(n428), .B(n16942), .Z(n16941) );
  XOR U16632 ( .A(p_input[1959]), .B(p_input[1927]), .Z(n16942) );
  XOR U16633 ( .A(n16943), .B(n16944), .Z(n16934) );
  AND U16634 ( .A(n16945), .B(n16946), .Z(n16944) );
  XOR U16635 ( .A(n16943), .B(n16652), .Z(n16946) );
  XNOR U16636 ( .A(p_input[1990]), .B(n16947), .Z(n16652) );
  AND U16637 ( .A(n430), .B(n16948), .Z(n16947) );
  XOR U16638 ( .A(p_input[2022]), .B(p_input[1990]), .Z(n16948) );
  XNOR U16639 ( .A(n16649), .B(n16943), .Z(n16945) );
  XOR U16640 ( .A(n16949), .B(n16950), .Z(n16649) );
  AND U16641 ( .A(n428), .B(n16951), .Z(n16950) );
  XOR U16642 ( .A(p_input[1958]), .B(p_input[1926]), .Z(n16951) );
  XOR U16643 ( .A(n16952), .B(n16953), .Z(n16943) );
  AND U16644 ( .A(n16954), .B(n16955), .Z(n16953) );
  XOR U16645 ( .A(n16952), .B(n16664), .Z(n16955) );
  XNOR U16646 ( .A(p_input[1989]), .B(n16956), .Z(n16664) );
  AND U16647 ( .A(n430), .B(n16957), .Z(n16956) );
  XOR U16648 ( .A(p_input[2021]), .B(p_input[1989]), .Z(n16957) );
  XNOR U16649 ( .A(n16661), .B(n16952), .Z(n16954) );
  XOR U16650 ( .A(n16958), .B(n16959), .Z(n16661) );
  AND U16651 ( .A(n428), .B(n16960), .Z(n16959) );
  XOR U16652 ( .A(p_input[1957]), .B(p_input[1925]), .Z(n16960) );
  XOR U16653 ( .A(n16961), .B(n16962), .Z(n16952) );
  AND U16654 ( .A(n16963), .B(n16964), .Z(n16962) );
  XOR U16655 ( .A(n16961), .B(n16676), .Z(n16964) );
  XNOR U16656 ( .A(p_input[1988]), .B(n16965), .Z(n16676) );
  AND U16657 ( .A(n430), .B(n16966), .Z(n16965) );
  XOR U16658 ( .A(p_input[2020]), .B(p_input[1988]), .Z(n16966) );
  XNOR U16659 ( .A(n16673), .B(n16961), .Z(n16963) );
  XOR U16660 ( .A(n16967), .B(n16968), .Z(n16673) );
  AND U16661 ( .A(n428), .B(n16969), .Z(n16968) );
  XOR U16662 ( .A(p_input[1956]), .B(p_input[1924]), .Z(n16969) );
  XOR U16663 ( .A(n16970), .B(n16971), .Z(n16961) );
  AND U16664 ( .A(n16972), .B(n16973), .Z(n16971) );
  XOR U16665 ( .A(n16970), .B(n16688), .Z(n16973) );
  XNOR U16666 ( .A(p_input[1987]), .B(n16974), .Z(n16688) );
  AND U16667 ( .A(n430), .B(n16975), .Z(n16974) );
  XOR U16668 ( .A(p_input[2019]), .B(p_input[1987]), .Z(n16975) );
  XNOR U16669 ( .A(n16685), .B(n16970), .Z(n16972) );
  XOR U16670 ( .A(n16976), .B(n16977), .Z(n16685) );
  AND U16671 ( .A(n428), .B(n16978), .Z(n16977) );
  XOR U16672 ( .A(p_input[1955]), .B(p_input[1923]), .Z(n16978) );
  XOR U16673 ( .A(n16979), .B(n16980), .Z(n16970) );
  AND U16674 ( .A(n16981), .B(n16982), .Z(n16980) );
  XOR U16675 ( .A(n16700), .B(n16979), .Z(n16982) );
  XNOR U16676 ( .A(p_input[1986]), .B(n16983), .Z(n16700) );
  AND U16677 ( .A(n430), .B(n16984), .Z(n16983) );
  XOR U16678 ( .A(p_input[2018]), .B(p_input[1986]), .Z(n16984) );
  XNOR U16679 ( .A(n16979), .B(n16697), .Z(n16981) );
  XOR U16680 ( .A(n16985), .B(n16986), .Z(n16697) );
  AND U16681 ( .A(n428), .B(n16987), .Z(n16986) );
  XOR U16682 ( .A(p_input[1954]), .B(p_input[1922]), .Z(n16987) );
  XOR U16683 ( .A(n16988), .B(n16989), .Z(n16979) );
  AND U16684 ( .A(n16990), .B(n16991), .Z(n16989) );
  XNOR U16685 ( .A(n16992), .B(n16713), .Z(n16991) );
  XNOR U16686 ( .A(p_input[1985]), .B(n16993), .Z(n16713) );
  AND U16687 ( .A(n430), .B(n16994), .Z(n16993) );
  XNOR U16688 ( .A(p_input[2017]), .B(n16995), .Z(n16994) );
  IV U16689 ( .A(p_input[1985]), .Z(n16995) );
  XNOR U16690 ( .A(n16710), .B(n16988), .Z(n16990) );
  XNOR U16691 ( .A(p_input[1921]), .B(n16996), .Z(n16710) );
  AND U16692 ( .A(n428), .B(n16997), .Z(n16996) );
  XOR U16693 ( .A(p_input[1953]), .B(p_input[1921]), .Z(n16997) );
  IV U16694 ( .A(n16992), .Z(n16988) );
  AND U16695 ( .A(n16718), .B(n16721), .Z(n16992) );
  XOR U16696 ( .A(p_input[1984]), .B(n16998), .Z(n16721) );
  AND U16697 ( .A(n430), .B(n16999), .Z(n16998) );
  XOR U16698 ( .A(p_input[2016]), .B(p_input[1984]), .Z(n16999) );
  XOR U16699 ( .A(n17000), .B(n17001), .Z(n430) );
  AND U16700 ( .A(n17002), .B(n17003), .Z(n17001) );
  XNOR U16701 ( .A(p_input[2047]), .B(n17000), .Z(n17003) );
  XOR U16702 ( .A(n17000), .B(p_input[2015]), .Z(n17002) );
  XOR U16703 ( .A(n17004), .B(n17005), .Z(n17000) );
  AND U16704 ( .A(n17006), .B(n17007), .Z(n17005) );
  XNOR U16705 ( .A(p_input[2046]), .B(n17004), .Z(n17007) );
  XOR U16706 ( .A(n17004), .B(p_input[2014]), .Z(n17006) );
  XOR U16707 ( .A(n17008), .B(n17009), .Z(n17004) );
  AND U16708 ( .A(n17010), .B(n17011), .Z(n17009) );
  XNOR U16709 ( .A(p_input[2045]), .B(n17008), .Z(n17011) );
  XOR U16710 ( .A(n17008), .B(p_input[2013]), .Z(n17010) );
  XOR U16711 ( .A(n17012), .B(n17013), .Z(n17008) );
  AND U16712 ( .A(n17014), .B(n17015), .Z(n17013) );
  XNOR U16713 ( .A(p_input[2044]), .B(n17012), .Z(n17015) );
  XOR U16714 ( .A(n17012), .B(p_input[2012]), .Z(n17014) );
  XOR U16715 ( .A(n17016), .B(n17017), .Z(n17012) );
  AND U16716 ( .A(n17018), .B(n17019), .Z(n17017) );
  XNOR U16717 ( .A(p_input[2043]), .B(n17016), .Z(n17019) );
  XOR U16718 ( .A(n17016), .B(p_input[2011]), .Z(n17018) );
  XOR U16719 ( .A(n17020), .B(n17021), .Z(n17016) );
  AND U16720 ( .A(n17022), .B(n17023), .Z(n17021) );
  XNOR U16721 ( .A(p_input[2042]), .B(n17020), .Z(n17023) );
  XOR U16722 ( .A(n17020), .B(p_input[2010]), .Z(n17022) );
  XOR U16723 ( .A(n17024), .B(n17025), .Z(n17020) );
  AND U16724 ( .A(n17026), .B(n17027), .Z(n17025) );
  XNOR U16725 ( .A(p_input[2041]), .B(n17024), .Z(n17027) );
  XOR U16726 ( .A(n17024), .B(p_input[2009]), .Z(n17026) );
  XOR U16727 ( .A(n17028), .B(n17029), .Z(n17024) );
  AND U16728 ( .A(n17030), .B(n17031), .Z(n17029) );
  XNOR U16729 ( .A(p_input[2040]), .B(n17028), .Z(n17031) );
  XOR U16730 ( .A(n17028), .B(p_input[2008]), .Z(n17030) );
  XOR U16731 ( .A(n17032), .B(n17033), .Z(n17028) );
  AND U16732 ( .A(n17034), .B(n17035), .Z(n17033) );
  XNOR U16733 ( .A(p_input[2039]), .B(n17032), .Z(n17035) );
  XOR U16734 ( .A(n17032), .B(p_input[2007]), .Z(n17034) );
  XOR U16735 ( .A(n17036), .B(n17037), .Z(n17032) );
  AND U16736 ( .A(n17038), .B(n17039), .Z(n17037) );
  XNOR U16737 ( .A(p_input[2038]), .B(n17036), .Z(n17039) );
  XOR U16738 ( .A(n17036), .B(p_input[2006]), .Z(n17038) );
  XOR U16739 ( .A(n17040), .B(n17041), .Z(n17036) );
  AND U16740 ( .A(n17042), .B(n17043), .Z(n17041) );
  XNOR U16741 ( .A(p_input[2037]), .B(n17040), .Z(n17043) );
  XOR U16742 ( .A(n17040), .B(p_input[2005]), .Z(n17042) );
  XOR U16743 ( .A(n17044), .B(n17045), .Z(n17040) );
  AND U16744 ( .A(n17046), .B(n17047), .Z(n17045) );
  XNOR U16745 ( .A(p_input[2036]), .B(n17044), .Z(n17047) );
  XOR U16746 ( .A(n17044), .B(p_input[2004]), .Z(n17046) );
  XOR U16747 ( .A(n17048), .B(n17049), .Z(n17044) );
  AND U16748 ( .A(n17050), .B(n17051), .Z(n17049) );
  XNOR U16749 ( .A(p_input[2035]), .B(n17048), .Z(n17051) );
  XOR U16750 ( .A(n17048), .B(p_input[2003]), .Z(n17050) );
  XOR U16751 ( .A(n17052), .B(n17053), .Z(n17048) );
  AND U16752 ( .A(n17054), .B(n17055), .Z(n17053) );
  XNOR U16753 ( .A(p_input[2034]), .B(n17052), .Z(n17055) );
  XOR U16754 ( .A(n17052), .B(p_input[2002]), .Z(n17054) );
  XOR U16755 ( .A(n17056), .B(n17057), .Z(n17052) );
  AND U16756 ( .A(n17058), .B(n17059), .Z(n17057) );
  XNOR U16757 ( .A(p_input[2033]), .B(n17056), .Z(n17059) );
  XOR U16758 ( .A(n17056), .B(p_input[2001]), .Z(n17058) );
  XOR U16759 ( .A(n17060), .B(n17061), .Z(n17056) );
  AND U16760 ( .A(n17062), .B(n17063), .Z(n17061) );
  XNOR U16761 ( .A(p_input[2032]), .B(n17060), .Z(n17063) );
  XOR U16762 ( .A(n17060), .B(p_input[2000]), .Z(n17062) );
  XOR U16763 ( .A(n17064), .B(n17065), .Z(n17060) );
  AND U16764 ( .A(n17066), .B(n17067), .Z(n17065) );
  XNOR U16765 ( .A(p_input[2031]), .B(n17064), .Z(n17067) );
  XOR U16766 ( .A(n17064), .B(p_input[1999]), .Z(n17066) );
  XOR U16767 ( .A(n17068), .B(n17069), .Z(n17064) );
  AND U16768 ( .A(n17070), .B(n17071), .Z(n17069) );
  XNOR U16769 ( .A(p_input[2030]), .B(n17068), .Z(n17071) );
  XOR U16770 ( .A(n17068), .B(p_input[1998]), .Z(n17070) );
  XOR U16771 ( .A(n17072), .B(n17073), .Z(n17068) );
  AND U16772 ( .A(n17074), .B(n17075), .Z(n17073) );
  XNOR U16773 ( .A(p_input[2029]), .B(n17072), .Z(n17075) );
  XOR U16774 ( .A(n17072), .B(p_input[1997]), .Z(n17074) );
  XOR U16775 ( .A(n17076), .B(n17077), .Z(n17072) );
  AND U16776 ( .A(n17078), .B(n17079), .Z(n17077) );
  XNOR U16777 ( .A(p_input[2028]), .B(n17076), .Z(n17079) );
  XOR U16778 ( .A(n17076), .B(p_input[1996]), .Z(n17078) );
  XOR U16779 ( .A(n17080), .B(n17081), .Z(n17076) );
  AND U16780 ( .A(n17082), .B(n17083), .Z(n17081) );
  XNOR U16781 ( .A(p_input[2027]), .B(n17080), .Z(n17083) );
  XOR U16782 ( .A(n17080), .B(p_input[1995]), .Z(n17082) );
  XOR U16783 ( .A(n17084), .B(n17085), .Z(n17080) );
  AND U16784 ( .A(n17086), .B(n17087), .Z(n17085) );
  XNOR U16785 ( .A(p_input[2026]), .B(n17084), .Z(n17087) );
  XOR U16786 ( .A(n17084), .B(p_input[1994]), .Z(n17086) );
  XOR U16787 ( .A(n17088), .B(n17089), .Z(n17084) );
  AND U16788 ( .A(n17090), .B(n17091), .Z(n17089) );
  XNOR U16789 ( .A(p_input[2025]), .B(n17088), .Z(n17091) );
  XOR U16790 ( .A(n17088), .B(p_input[1993]), .Z(n17090) );
  XOR U16791 ( .A(n17092), .B(n17093), .Z(n17088) );
  AND U16792 ( .A(n17094), .B(n17095), .Z(n17093) );
  XNOR U16793 ( .A(p_input[2024]), .B(n17092), .Z(n17095) );
  XOR U16794 ( .A(n17092), .B(p_input[1992]), .Z(n17094) );
  XOR U16795 ( .A(n17096), .B(n17097), .Z(n17092) );
  AND U16796 ( .A(n17098), .B(n17099), .Z(n17097) );
  XNOR U16797 ( .A(p_input[2023]), .B(n17096), .Z(n17099) );
  XOR U16798 ( .A(n17096), .B(p_input[1991]), .Z(n17098) );
  XOR U16799 ( .A(n17100), .B(n17101), .Z(n17096) );
  AND U16800 ( .A(n17102), .B(n17103), .Z(n17101) );
  XNOR U16801 ( .A(p_input[2022]), .B(n17100), .Z(n17103) );
  XOR U16802 ( .A(n17100), .B(p_input[1990]), .Z(n17102) );
  XOR U16803 ( .A(n17104), .B(n17105), .Z(n17100) );
  AND U16804 ( .A(n17106), .B(n17107), .Z(n17105) );
  XNOR U16805 ( .A(p_input[2021]), .B(n17104), .Z(n17107) );
  XOR U16806 ( .A(n17104), .B(p_input[1989]), .Z(n17106) );
  XOR U16807 ( .A(n17108), .B(n17109), .Z(n17104) );
  AND U16808 ( .A(n17110), .B(n17111), .Z(n17109) );
  XNOR U16809 ( .A(p_input[2020]), .B(n17108), .Z(n17111) );
  XOR U16810 ( .A(n17108), .B(p_input[1988]), .Z(n17110) );
  XOR U16811 ( .A(n17112), .B(n17113), .Z(n17108) );
  AND U16812 ( .A(n17114), .B(n17115), .Z(n17113) );
  XNOR U16813 ( .A(p_input[2019]), .B(n17112), .Z(n17115) );
  XOR U16814 ( .A(n17112), .B(p_input[1987]), .Z(n17114) );
  XOR U16815 ( .A(n17116), .B(n17117), .Z(n17112) );
  AND U16816 ( .A(n17118), .B(n17119), .Z(n17117) );
  XNOR U16817 ( .A(p_input[2018]), .B(n17116), .Z(n17119) );
  XOR U16818 ( .A(n17116), .B(p_input[1986]), .Z(n17118) );
  XNOR U16819 ( .A(n17120), .B(n17121), .Z(n17116) );
  AND U16820 ( .A(n17122), .B(n17123), .Z(n17121) );
  XOR U16821 ( .A(p_input[2017]), .B(n17120), .Z(n17123) );
  XNOR U16822 ( .A(p_input[1985]), .B(n17120), .Z(n17122) );
  AND U16823 ( .A(p_input[2016]), .B(n17124), .Z(n17120) );
  IV U16824 ( .A(p_input[1984]), .Z(n17124) );
  XNOR U16825 ( .A(p_input[1920]), .B(n17125), .Z(n16718) );
  AND U16826 ( .A(n428), .B(n17126), .Z(n17125) );
  XOR U16827 ( .A(p_input[1952]), .B(p_input[1920]), .Z(n17126) );
  XOR U16828 ( .A(n17127), .B(n17128), .Z(n428) );
  AND U16829 ( .A(n17129), .B(n17130), .Z(n17128) );
  XNOR U16830 ( .A(p_input[1983]), .B(n17127), .Z(n17130) );
  XOR U16831 ( .A(n17127), .B(p_input[1951]), .Z(n17129) );
  XOR U16832 ( .A(n17131), .B(n17132), .Z(n17127) );
  AND U16833 ( .A(n17133), .B(n17134), .Z(n17132) );
  XNOR U16834 ( .A(p_input[1982]), .B(n17131), .Z(n17134) );
  XNOR U16835 ( .A(n17131), .B(n16733), .Z(n17133) );
  IV U16836 ( .A(p_input[1950]), .Z(n16733) );
  XOR U16837 ( .A(n17135), .B(n17136), .Z(n17131) );
  AND U16838 ( .A(n17137), .B(n17138), .Z(n17136) );
  XNOR U16839 ( .A(p_input[1981]), .B(n17135), .Z(n17138) );
  XNOR U16840 ( .A(n17135), .B(n16742), .Z(n17137) );
  IV U16841 ( .A(p_input[1949]), .Z(n16742) );
  XOR U16842 ( .A(n17139), .B(n17140), .Z(n17135) );
  AND U16843 ( .A(n17141), .B(n17142), .Z(n17140) );
  XNOR U16844 ( .A(p_input[1980]), .B(n17139), .Z(n17142) );
  XNOR U16845 ( .A(n17139), .B(n16751), .Z(n17141) );
  IV U16846 ( .A(p_input[1948]), .Z(n16751) );
  XOR U16847 ( .A(n17143), .B(n17144), .Z(n17139) );
  AND U16848 ( .A(n17145), .B(n17146), .Z(n17144) );
  XNOR U16849 ( .A(p_input[1979]), .B(n17143), .Z(n17146) );
  XNOR U16850 ( .A(n17143), .B(n16760), .Z(n17145) );
  IV U16851 ( .A(p_input[1947]), .Z(n16760) );
  XOR U16852 ( .A(n17147), .B(n17148), .Z(n17143) );
  AND U16853 ( .A(n17149), .B(n17150), .Z(n17148) );
  XNOR U16854 ( .A(p_input[1978]), .B(n17147), .Z(n17150) );
  XNOR U16855 ( .A(n17147), .B(n16769), .Z(n17149) );
  IV U16856 ( .A(p_input[1946]), .Z(n16769) );
  XOR U16857 ( .A(n17151), .B(n17152), .Z(n17147) );
  AND U16858 ( .A(n17153), .B(n17154), .Z(n17152) );
  XNOR U16859 ( .A(p_input[1977]), .B(n17151), .Z(n17154) );
  XNOR U16860 ( .A(n17151), .B(n16778), .Z(n17153) );
  IV U16861 ( .A(p_input[1945]), .Z(n16778) );
  XOR U16862 ( .A(n17155), .B(n17156), .Z(n17151) );
  AND U16863 ( .A(n17157), .B(n17158), .Z(n17156) );
  XNOR U16864 ( .A(p_input[1976]), .B(n17155), .Z(n17158) );
  XNOR U16865 ( .A(n17155), .B(n16787), .Z(n17157) );
  IV U16866 ( .A(p_input[1944]), .Z(n16787) );
  XOR U16867 ( .A(n17159), .B(n17160), .Z(n17155) );
  AND U16868 ( .A(n17161), .B(n17162), .Z(n17160) );
  XNOR U16869 ( .A(p_input[1975]), .B(n17159), .Z(n17162) );
  XNOR U16870 ( .A(n17159), .B(n16796), .Z(n17161) );
  IV U16871 ( .A(p_input[1943]), .Z(n16796) );
  XOR U16872 ( .A(n17163), .B(n17164), .Z(n17159) );
  AND U16873 ( .A(n17165), .B(n17166), .Z(n17164) );
  XNOR U16874 ( .A(p_input[1974]), .B(n17163), .Z(n17166) );
  XNOR U16875 ( .A(n17163), .B(n16805), .Z(n17165) );
  IV U16876 ( .A(p_input[1942]), .Z(n16805) );
  XOR U16877 ( .A(n17167), .B(n17168), .Z(n17163) );
  AND U16878 ( .A(n17169), .B(n17170), .Z(n17168) );
  XNOR U16879 ( .A(p_input[1973]), .B(n17167), .Z(n17170) );
  XNOR U16880 ( .A(n17167), .B(n16814), .Z(n17169) );
  IV U16881 ( .A(p_input[1941]), .Z(n16814) );
  XOR U16882 ( .A(n17171), .B(n17172), .Z(n17167) );
  AND U16883 ( .A(n17173), .B(n17174), .Z(n17172) );
  XNOR U16884 ( .A(p_input[1972]), .B(n17171), .Z(n17174) );
  XNOR U16885 ( .A(n17171), .B(n16823), .Z(n17173) );
  IV U16886 ( .A(p_input[1940]), .Z(n16823) );
  XOR U16887 ( .A(n17175), .B(n17176), .Z(n17171) );
  AND U16888 ( .A(n17177), .B(n17178), .Z(n17176) );
  XNOR U16889 ( .A(p_input[1971]), .B(n17175), .Z(n17178) );
  XNOR U16890 ( .A(n17175), .B(n16832), .Z(n17177) );
  IV U16891 ( .A(p_input[1939]), .Z(n16832) );
  XOR U16892 ( .A(n17179), .B(n17180), .Z(n17175) );
  AND U16893 ( .A(n17181), .B(n17182), .Z(n17180) );
  XNOR U16894 ( .A(p_input[1970]), .B(n17179), .Z(n17182) );
  XNOR U16895 ( .A(n17179), .B(n16841), .Z(n17181) );
  IV U16896 ( .A(p_input[1938]), .Z(n16841) );
  XOR U16897 ( .A(n17183), .B(n17184), .Z(n17179) );
  AND U16898 ( .A(n17185), .B(n17186), .Z(n17184) );
  XNOR U16899 ( .A(p_input[1969]), .B(n17183), .Z(n17186) );
  XNOR U16900 ( .A(n17183), .B(n16850), .Z(n17185) );
  IV U16901 ( .A(p_input[1937]), .Z(n16850) );
  XOR U16902 ( .A(n17187), .B(n17188), .Z(n17183) );
  AND U16903 ( .A(n17189), .B(n17190), .Z(n17188) );
  XNOR U16904 ( .A(p_input[1968]), .B(n17187), .Z(n17190) );
  XNOR U16905 ( .A(n17187), .B(n16859), .Z(n17189) );
  IV U16906 ( .A(p_input[1936]), .Z(n16859) );
  XOR U16907 ( .A(n17191), .B(n17192), .Z(n17187) );
  AND U16908 ( .A(n17193), .B(n17194), .Z(n17192) );
  XNOR U16909 ( .A(p_input[1967]), .B(n17191), .Z(n17194) );
  XNOR U16910 ( .A(n17191), .B(n16868), .Z(n17193) );
  IV U16911 ( .A(p_input[1935]), .Z(n16868) );
  XOR U16912 ( .A(n17195), .B(n17196), .Z(n17191) );
  AND U16913 ( .A(n17197), .B(n17198), .Z(n17196) );
  XNOR U16914 ( .A(p_input[1966]), .B(n17195), .Z(n17198) );
  XNOR U16915 ( .A(n17195), .B(n16877), .Z(n17197) );
  IV U16916 ( .A(p_input[1934]), .Z(n16877) );
  XOR U16917 ( .A(n17199), .B(n17200), .Z(n17195) );
  AND U16918 ( .A(n17201), .B(n17202), .Z(n17200) );
  XNOR U16919 ( .A(p_input[1965]), .B(n17199), .Z(n17202) );
  XNOR U16920 ( .A(n17199), .B(n16886), .Z(n17201) );
  IV U16921 ( .A(p_input[1933]), .Z(n16886) );
  XOR U16922 ( .A(n17203), .B(n17204), .Z(n17199) );
  AND U16923 ( .A(n17205), .B(n17206), .Z(n17204) );
  XNOR U16924 ( .A(p_input[1964]), .B(n17203), .Z(n17206) );
  XNOR U16925 ( .A(n17203), .B(n16895), .Z(n17205) );
  IV U16926 ( .A(p_input[1932]), .Z(n16895) );
  XOR U16927 ( .A(n17207), .B(n17208), .Z(n17203) );
  AND U16928 ( .A(n17209), .B(n17210), .Z(n17208) );
  XNOR U16929 ( .A(p_input[1963]), .B(n17207), .Z(n17210) );
  XNOR U16930 ( .A(n17207), .B(n16904), .Z(n17209) );
  IV U16931 ( .A(p_input[1931]), .Z(n16904) );
  XOR U16932 ( .A(n17211), .B(n17212), .Z(n17207) );
  AND U16933 ( .A(n17213), .B(n17214), .Z(n17212) );
  XNOR U16934 ( .A(p_input[1962]), .B(n17211), .Z(n17214) );
  XNOR U16935 ( .A(n17211), .B(n16913), .Z(n17213) );
  IV U16936 ( .A(p_input[1930]), .Z(n16913) );
  XOR U16937 ( .A(n17215), .B(n17216), .Z(n17211) );
  AND U16938 ( .A(n17217), .B(n17218), .Z(n17216) );
  XNOR U16939 ( .A(p_input[1961]), .B(n17215), .Z(n17218) );
  XNOR U16940 ( .A(n17215), .B(n16922), .Z(n17217) );
  IV U16941 ( .A(p_input[1929]), .Z(n16922) );
  XOR U16942 ( .A(n17219), .B(n17220), .Z(n17215) );
  AND U16943 ( .A(n17221), .B(n17222), .Z(n17220) );
  XNOR U16944 ( .A(p_input[1960]), .B(n17219), .Z(n17222) );
  XNOR U16945 ( .A(n17219), .B(n16931), .Z(n17221) );
  IV U16946 ( .A(p_input[1928]), .Z(n16931) );
  XOR U16947 ( .A(n17223), .B(n17224), .Z(n17219) );
  AND U16948 ( .A(n17225), .B(n17226), .Z(n17224) );
  XNOR U16949 ( .A(p_input[1959]), .B(n17223), .Z(n17226) );
  XNOR U16950 ( .A(n17223), .B(n16940), .Z(n17225) );
  IV U16951 ( .A(p_input[1927]), .Z(n16940) );
  XOR U16952 ( .A(n17227), .B(n17228), .Z(n17223) );
  AND U16953 ( .A(n17229), .B(n17230), .Z(n17228) );
  XNOR U16954 ( .A(p_input[1958]), .B(n17227), .Z(n17230) );
  XNOR U16955 ( .A(n17227), .B(n16949), .Z(n17229) );
  IV U16956 ( .A(p_input[1926]), .Z(n16949) );
  XOR U16957 ( .A(n17231), .B(n17232), .Z(n17227) );
  AND U16958 ( .A(n17233), .B(n17234), .Z(n17232) );
  XNOR U16959 ( .A(p_input[1957]), .B(n17231), .Z(n17234) );
  XNOR U16960 ( .A(n17231), .B(n16958), .Z(n17233) );
  IV U16961 ( .A(p_input[1925]), .Z(n16958) );
  XOR U16962 ( .A(n17235), .B(n17236), .Z(n17231) );
  AND U16963 ( .A(n17237), .B(n17238), .Z(n17236) );
  XNOR U16964 ( .A(p_input[1956]), .B(n17235), .Z(n17238) );
  XNOR U16965 ( .A(n17235), .B(n16967), .Z(n17237) );
  IV U16966 ( .A(p_input[1924]), .Z(n16967) );
  XOR U16967 ( .A(n17239), .B(n17240), .Z(n17235) );
  AND U16968 ( .A(n17241), .B(n17242), .Z(n17240) );
  XNOR U16969 ( .A(p_input[1955]), .B(n17239), .Z(n17242) );
  XNOR U16970 ( .A(n17239), .B(n16976), .Z(n17241) );
  IV U16971 ( .A(p_input[1923]), .Z(n16976) );
  XOR U16972 ( .A(n17243), .B(n17244), .Z(n17239) );
  AND U16973 ( .A(n17245), .B(n17246), .Z(n17244) );
  XNOR U16974 ( .A(p_input[1954]), .B(n17243), .Z(n17246) );
  XNOR U16975 ( .A(n17243), .B(n16985), .Z(n17245) );
  IV U16976 ( .A(p_input[1922]), .Z(n16985) );
  XNOR U16977 ( .A(n17247), .B(n17248), .Z(n17243) );
  AND U16978 ( .A(n17249), .B(n17250), .Z(n17248) );
  XOR U16979 ( .A(p_input[1953]), .B(n17247), .Z(n17250) );
  XNOR U16980 ( .A(p_input[1921]), .B(n17247), .Z(n17249) );
  AND U16981 ( .A(p_input[1952]), .B(n17251), .Z(n17247) );
  IV U16982 ( .A(p_input[1920]), .Z(n17251) );
  XOR U16983 ( .A(n17252), .B(n17253), .Z(n16341) );
  AND U16984 ( .A(n364), .B(n17254), .Z(n17253) );
  XNOR U16985 ( .A(n17255), .B(n17252), .Z(n17254) );
  XOR U16986 ( .A(n17256), .B(n17257), .Z(n364) );
  AND U16987 ( .A(n17258), .B(n17259), .Z(n17257) );
  XNOR U16988 ( .A(n16356), .B(n17256), .Z(n17259) );
  AND U16989 ( .A(p_input[1919]), .B(p_input[1887]), .Z(n16356) );
  XNOR U16990 ( .A(n17256), .B(n16353), .Z(n17258) );
  IV U16991 ( .A(n17260), .Z(n16353) );
  AND U16992 ( .A(p_input[1823]), .B(p_input[1855]), .Z(n17260) );
  XOR U16993 ( .A(n17261), .B(n17262), .Z(n17256) );
  AND U16994 ( .A(n17263), .B(n17264), .Z(n17262) );
  XOR U16995 ( .A(n17261), .B(n16368), .Z(n17264) );
  XNOR U16996 ( .A(p_input[1886]), .B(n17265), .Z(n16368) );
  AND U16997 ( .A(n434), .B(n17266), .Z(n17265) );
  XOR U16998 ( .A(p_input[1918]), .B(p_input[1886]), .Z(n17266) );
  XNOR U16999 ( .A(n16365), .B(n17261), .Z(n17263) );
  XOR U17000 ( .A(n17267), .B(n17268), .Z(n16365) );
  AND U17001 ( .A(n431), .B(n17269), .Z(n17268) );
  XOR U17002 ( .A(p_input[1854]), .B(p_input[1822]), .Z(n17269) );
  XOR U17003 ( .A(n17270), .B(n17271), .Z(n17261) );
  AND U17004 ( .A(n17272), .B(n17273), .Z(n17271) );
  XOR U17005 ( .A(n17270), .B(n16380), .Z(n17273) );
  XNOR U17006 ( .A(p_input[1885]), .B(n17274), .Z(n16380) );
  AND U17007 ( .A(n434), .B(n17275), .Z(n17274) );
  XOR U17008 ( .A(p_input[1917]), .B(p_input[1885]), .Z(n17275) );
  XNOR U17009 ( .A(n16377), .B(n17270), .Z(n17272) );
  XOR U17010 ( .A(n17276), .B(n17277), .Z(n16377) );
  AND U17011 ( .A(n431), .B(n17278), .Z(n17277) );
  XOR U17012 ( .A(p_input[1853]), .B(p_input[1821]), .Z(n17278) );
  XOR U17013 ( .A(n17279), .B(n17280), .Z(n17270) );
  AND U17014 ( .A(n17281), .B(n17282), .Z(n17280) );
  XOR U17015 ( .A(n17279), .B(n16392), .Z(n17282) );
  XNOR U17016 ( .A(p_input[1884]), .B(n17283), .Z(n16392) );
  AND U17017 ( .A(n434), .B(n17284), .Z(n17283) );
  XOR U17018 ( .A(p_input[1916]), .B(p_input[1884]), .Z(n17284) );
  XNOR U17019 ( .A(n16389), .B(n17279), .Z(n17281) );
  XOR U17020 ( .A(n17285), .B(n17286), .Z(n16389) );
  AND U17021 ( .A(n431), .B(n17287), .Z(n17286) );
  XOR U17022 ( .A(p_input[1852]), .B(p_input[1820]), .Z(n17287) );
  XOR U17023 ( .A(n17288), .B(n17289), .Z(n17279) );
  AND U17024 ( .A(n17290), .B(n17291), .Z(n17289) );
  XOR U17025 ( .A(n17288), .B(n16404), .Z(n17291) );
  XNOR U17026 ( .A(p_input[1883]), .B(n17292), .Z(n16404) );
  AND U17027 ( .A(n434), .B(n17293), .Z(n17292) );
  XOR U17028 ( .A(p_input[1915]), .B(p_input[1883]), .Z(n17293) );
  XNOR U17029 ( .A(n16401), .B(n17288), .Z(n17290) );
  XOR U17030 ( .A(n17294), .B(n17295), .Z(n16401) );
  AND U17031 ( .A(n431), .B(n17296), .Z(n17295) );
  XOR U17032 ( .A(p_input[1851]), .B(p_input[1819]), .Z(n17296) );
  XOR U17033 ( .A(n17297), .B(n17298), .Z(n17288) );
  AND U17034 ( .A(n17299), .B(n17300), .Z(n17298) );
  XOR U17035 ( .A(n17297), .B(n16416), .Z(n17300) );
  XNOR U17036 ( .A(p_input[1882]), .B(n17301), .Z(n16416) );
  AND U17037 ( .A(n434), .B(n17302), .Z(n17301) );
  XOR U17038 ( .A(p_input[1914]), .B(p_input[1882]), .Z(n17302) );
  XNOR U17039 ( .A(n16413), .B(n17297), .Z(n17299) );
  XOR U17040 ( .A(n17303), .B(n17304), .Z(n16413) );
  AND U17041 ( .A(n431), .B(n17305), .Z(n17304) );
  XOR U17042 ( .A(p_input[1850]), .B(p_input[1818]), .Z(n17305) );
  XOR U17043 ( .A(n17306), .B(n17307), .Z(n17297) );
  AND U17044 ( .A(n17308), .B(n17309), .Z(n17307) );
  XOR U17045 ( .A(n17306), .B(n16428), .Z(n17309) );
  XNOR U17046 ( .A(p_input[1881]), .B(n17310), .Z(n16428) );
  AND U17047 ( .A(n434), .B(n17311), .Z(n17310) );
  XOR U17048 ( .A(p_input[1913]), .B(p_input[1881]), .Z(n17311) );
  XNOR U17049 ( .A(n16425), .B(n17306), .Z(n17308) );
  XOR U17050 ( .A(n17312), .B(n17313), .Z(n16425) );
  AND U17051 ( .A(n431), .B(n17314), .Z(n17313) );
  XOR U17052 ( .A(p_input[1849]), .B(p_input[1817]), .Z(n17314) );
  XOR U17053 ( .A(n17315), .B(n17316), .Z(n17306) );
  AND U17054 ( .A(n17317), .B(n17318), .Z(n17316) );
  XOR U17055 ( .A(n17315), .B(n16440), .Z(n17318) );
  XNOR U17056 ( .A(p_input[1880]), .B(n17319), .Z(n16440) );
  AND U17057 ( .A(n434), .B(n17320), .Z(n17319) );
  XOR U17058 ( .A(p_input[1912]), .B(p_input[1880]), .Z(n17320) );
  XNOR U17059 ( .A(n16437), .B(n17315), .Z(n17317) );
  XOR U17060 ( .A(n17321), .B(n17322), .Z(n16437) );
  AND U17061 ( .A(n431), .B(n17323), .Z(n17322) );
  XOR U17062 ( .A(p_input[1848]), .B(p_input[1816]), .Z(n17323) );
  XOR U17063 ( .A(n17324), .B(n17325), .Z(n17315) );
  AND U17064 ( .A(n17326), .B(n17327), .Z(n17325) );
  XOR U17065 ( .A(n17324), .B(n16452), .Z(n17327) );
  XNOR U17066 ( .A(p_input[1879]), .B(n17328), .Z(n16452) );
  AND U17067 ( .A(n434), .B(n17329), .Z(n17328) );
  XOR U17068 ( .A(p_input[1911]), .B(p_input[1879]), .Z(n17329) );
  XNOR U17069 ( .A(n16449), .B(n17324), .Z(n17326) );
  XOR U17070 ( .A(n17330), .B(n17331), .Z(n16449) );
  AND U17071 ( .A(n431), .B(n17332), .Z(n17331) );
  XOR U17072 ( .A(p_input[1847]), .B(p_input[1815]), .Z(n17332) );
  XOR U17073 ( .A(n17333), .B(n17334), .Z(n17324) );
  AND U17074 ( .A(n17335), .B(n17336), .Z(n17334) );
  XOR U17075 ( .A(n17333), .B(n16464), .Z(n17336) );
  XNOR U17076 ( .A(p_input[1878]), .B(n17337), .Z(n16464) );
  AND U17077 ( .A(n434), .B(n17338), .Z(n17337) );
  XOR U17078 ( .A(p_input[1910]), .B(p_input[1878]), .Z(n17338) );
  XNOR U17079 ( .A(n16461), .B(n17333), .Z(n17335) );
  XOR U17080 ( .A(n17339), .B(n17340), .Z(n16461) );
  AND U17081 ( .A(n431), .B(n17341), .Z(n17340) );
  XOR U17082 ( .A(p_input[1846]), .B(p_input[1814]), .Z(n17341) );
  XOR U17083 ( .A(n17342), .B(n17343), .Z(n17333) );
  AND U17084 ( .A(n17344), .B(n17345), .Z(n17343) );
  XOR U17085 ( .A(n17342), .B(n16476), .Z(n17345) );
  XNOR U17086 ( .A(p_input[1877]), .B(n17346), .Z(n16476) );
  AND U17087 ( .A(n434), .B(n17347), .Z(n17346) );
  XOR U17088 ( .A(p_input[1909]), .B(p_input[1877]), .Z(n17347) );
  XNOR U17089 ( .A(n16473), .B(n17342), .Z(n17344) );
  XOR U17090 ( .A(n17348), .B(n17349), .Z(n16473) );
  AND U17091 ( .A(n431), .B(n17350), .Z(n17349) );
  XOR U17092 ( .A(p_input[1845]), .B(p_input[1813]), .Z(n17350) );
  XOR U17093 ( .A(n17351), .B(n17352), .Z(n17342) );
  AND U17094 ( .A(n17353), .B(n17354), .Z(n17352) );
  XOR U17095 ( .A(n17351), .B(n16488), .Z(n17354) );
  XNOR U17096 ( .A(p_input[1876]), .B(n17355), .Z(n16488) );
  AND U17097 ( .A(n434), .B(n17356), .Z(n17355) );
  XOR U17098 ( .A(p_input[1908]), .B(p_input[1876]), .Z(n17356) );
  XNOR U17099 ( .A(n16485), .B(n17351), .Z(n17353) );
  XOR U17100 ( .A(n17357), .B(n17358), .Z(n16485) );
  AND U17101 ( .A(n431), .B(n17359), .Z(n17358) );
  XOR U17102 ( .A(p_input[1844]), .B(p_input[1812]), .Z(n17359) );
  XOR U17103 ( .A(n17360), .B(n17361), .Z(n17351) );
  AND U17104 ( .A(n17362), .B(n17363), .Z(n17361) );
  XOR U17105 ( .A(n17360), .B(n16500), .Z(n17363) );
  XNOR U17106 ( .A(p_input[1875]), .B(n17364), .Z(n16500) );
  AND U17107 ( .A(n434), .B(n17365), .Z(n17364) );
  XOR U17108 ( .A(p_input[1907]), .B(p_input[1875]), .Z(n17365) );
  XNOR U17109 ( .A(n16497), .B(n17360), .Z(n17362) );
  XOR U17110 ( .A(n17366), .B(n17367), .Z(n16497) );
  AND U17111 ( .A(n431), .B(n17368), .Z(n17367) );
  XOR U17112 ( .A(p_input[1843]), .B(p_input[1811]), .Z(n17368) );
  XOR U17113 ( .A(n17369), .B(n17370), .Z(n17360) );
  AND U17114 ( .A(n17371), .B(n17372), .Z(n17370) );
  XOR U17115 ( .A(n17369), .B(n16512), .Z(n17372) );
  XNOR U17116 ( .A(p_input[1874]), .B(n17373), .Z(n16512) );
  AND U17117 ( .A(n434), .B(n17374), .Z(n17373) );
  XOR U17118 ( .A(p_input[1906]), .B(p_input[1874]), .Z(n17374) );
  XNOR U17119 ( .A(n16509), .B(n17369), .Z(n17371) );
  XOR U17120 ( .A(n17375), .B(n17376), .Z(n16509) );
  AND U17121 ( .A(n431), .B(n17377), .Z(n17376) );
  XOR U17122 ( .A(p_input[1842]), .B(p_input[1810]), .Z(n17377) );
  XOR U17123 ( .A(n17378), .B(n17379), .Z(n17369) );
  AND U17124 ( .A(n17380), .B(n17381), .Z(n17379) );
  XOR U17125 ( .A(n17378), .B(n16524), .Z(n17381) );
  XNOR U17126 ( .A(p_input[1873]), .B(n17382), .Z(n16524) );
  AND U17127 ( .A(n434), .B(n17383), .Z(n17382) );
  XOR U17128 ( .A(p_input[1905]), .B(p_input[1873]), .Z(n17383) );
  XNOR U17129 ( .A(n16521), .B(n17378), .Z(n17380) );
  XOR U17130 ( .A(n17384), .B(n17385), .Z(n16521) );
  AND U17131 ( .A(n431), .B(n17386), .Z(n17385) );
  XOR U17132 ( .A(p_input[1841]), .B(p_input[1809]), .Z(n17386) );
  XOR U17133 ( .A(n17387), .B(n17388), .Z(n17378) );
  AND U17134 ( .A(n17389), .B(n17390), .Z(n17388) );
  XOR U17135 ( .A(n17387), .B(n16536), .Z(n17390) );
  XNOR U17136 ( .A(p_input[1872]), .B(n17391), .Z(n16536) );
  AND U17137 ( .A(n434), .B(n17392), .Z(n17391) );
  XOR U17138 ( .A(p_input[1904]), .B(p_input[1872]), .Z(n17392) );
  XNOR U17139 ( .A(n16533), .B(n17387), .Z(n17389) );
  XOR U17140 ( .A(n17393), .B(n17394), .Z(n16533) );
  AND U17141 ( .A(n431), .B(n17395), .Z(n17394) );
  XOR U17142 ( .A(p_input[1840]), .B(p_input[1808]), .Z(n17395) );
  XOR U17143 ( .A(n17396), .B(n17397), .Z(n17387) );
  AND U17144 ( .A(n17398), .B(n17399), .Z(n17397) );
  XOR U17145 ( .A(n17396), .B(n16548), .Z(n17399) );
  XNOR U17146 ( .A(p_input[1871]), .B(n17400), .Z(n16548) );
  AND U17147 ( .A(n434), .B(n17401), .Z(n17400) );
  XOR U17148 ( .A(p_input[1903]), .B(p_input[1871]), .Z(n17401) );
  XNOR U17149 ( .A(n16545), .B(n17396), .Z(n17398) );
  XOR U17150 ( .A(n17402), .B(n17403), .Z(n16545) );
  AND U17151 ( .A(n431), .B(n17404), .Z(n17403) );
  XOR U17152 ( .A(p_input[1839]), .B(p_input[1807]), .Z(n17404) );
  XOR U17153 ( .A(n17405), .B(n17406), .Z(n17396) );
  AND U17154 ( .A(n17407), .B(n17408), .Z(n17406) );
  XOR U17155 ( .A(n17405), .B(n16560), .Z(n17408) );
  XNOR U17156 ( .A(p_input[1870]), .B(n17409), .Z(n16560) );
  AND U17157 ( .A(n434), .B(n17410), .Z(n17409) );
  XOR U17158 ( .A(p_input[1902]), .B(p_input[1870]), .Z(n17410) );
  XNOR U17159 ( .A(n16557), .B(n17405), .Z(n17407) );
  XOR U17160 ( .A(n17411), .B(n17412), .Z(n16557) );
  AND U17161 ( .A(n431), .B(n17413), .Z(n17412) );
  XOR U17162 ( .A(p_input[1838]), .B(p_input[1806]), .Z(n17413) );
  XOR U17163 ( .A(n17414), .B(n17415), .Z(n17405) );
  AND U17164 ( .A(n17416), .B(n17417), .Z(n17415) );
  XOR U17165 ( .A(n17414), .B(n16572), .Z(n17417) );
  XNOR U17166 ( .A(p_input[1869]), .B(n17418), .Z(n16572) );
  AND U17167 ( .A(n434), .B(n17419), .Z(n17418) );
  XOR U17168 ( .A(p_input[1901]), .B(p_input[1869]), .Z(n17419) );
  XNOR U17169 ( .A(n16569), .B(n17414), .Z(n17416) );
  XOR U17170 ( .A(n17420), .B(n17421), .Z(n16569) );
  AND U17171 ( .A(n431), .B(n17422), .Z(n17421) );
  XOR U17172 ( .A(p_input[1837]), .B(p_input[1805]), .Z(n17422) );
  XOR U17173 ( .A(n17423), .B(n17424), .Z(n17414) );
  AND U17174 ( .A(n17425), .B(n17426), .Z(n17424) );
  XOR U17175 ( .A(n17423), .B(n16584), .Z(n17426) );
  XNOR U17176 ( .A(p_input[1868]), .B(n17427), .Z(n16584) );
  AND U17177 ( .A(n434), .B(n17428), .Z(n17427) );
  XOR U17178 ( .A(p_input[1900]), .B(p_input[1868]), .Z(n17428) );
  XNOR U17179 ( .A(n16581), .B(n17423), .Z(n17425) );
  XOR U17180 ( .A(n17429), .B(n17430), .Z(n16581) );
  AND U17181 ( .A(n431), .B(n17431), .Z(n17430) );
  XOR U17182 ( .A(p_input[1836]), .B(p_input[1804]), .Z(n17431) );
  XOR U17183 ( .A(n17432), .B(n17433), .Z(n17423) );
  AND U17184 ( .A(n17434), .B(n17435), .Z(n17433) );
  XOR U17185 ( .A(n17432), .B(n16596), .Z(n17435) );
  XNOR U17186 ( .A(p_input[1867]), .B(n17436), .Z(n16596) );
  AND U17187 ( .A(n434), .B(n17437), .Z(n17436) );
  XOR U17188 ( .A(p_input[1899]), .B(p_input[1867]), .Z(n17437) );
  XNOR U17189 ( .A(n16593), .B(n17432), .Z(n17434) );
  XOR U17190 ( .A(n17438), .B(n17439), .Z(n16593) );
  AND U17191 ( .A(n431), .B(n17440), .Z(n17439) );
  XOR U17192 ( .A(p_input[1835]), .B(p_input[1803]), .Z(n17440) );
  XOR U17193 ( .A(n17441), .B(n17442), .Z(n17432) );
  AND U17194 ( .A(n17443), .B(n17444), .Z(n17442) );
  XOR U17195 ( .A(n17441), .B(n16608), .Z(n17444) );
  XNOR U17196 ( .A(p_input[1866]), .B(n17445), .Z(n16608) );
  AND U17197 ( .A(n434), .B(n17446), .Z(n17445) );
  XOR U17198 ( .A(p_input[1898]), .B(p_input[1866]), .Z(n17446) );
  XNOR U17199 ( .A(n16605), .B(n17441), .Z(n17443) );
  XOR U17200 ( .A(n17447), .B(n17448), .Z(n16605) );
  AND U17201 ( .A(n431), .B(n17449), .Z(n17448) );
  XOR U17202 ( .A(p_input[1834]), .B(p_input[1802]), .Z(n17449) );
  XOR U17203 ( .A(n17450), .B(n17451), .Z(n17441) );
  AND U17204 ( .A(n17452), .B(n17453), .Z(n17451) );
  XOR U17205 ( .A(n17450), .B(n16620), .Z(n17453) );
  XNOR U17206 ( .A(p_input[1865]), .B(n17454), .Z(n16620) );
  AND U17207 ( .A(n434), .B(n17455), .Z(n17454) );
  XOR U17208 ( .A(p_input[1897]), .B(p_input[1865]), .Z(n17455) );
  XNOR U17209 ( .A(n16617), .B(n17450), .Z(n17452) );
  XOR U17210 ( .A(n17456), .B(n17457), .Z(n16617) );
  AND U17211 ( .A(n431), .B(n17458), .Z(n17457) );
  XOR U17212 ( .A(p_input[1833]), .B(p_input[1801]), .Z(n17458) );
  XOR U17213 ( .A(n17459), .B(n17460), .Z(n17450) );
  AND U17214 ( .A(n17461), .B(n17462), .Z(n17460) );
  XOR U17215 ( .A(n17459), .B(n16632), .Z(n17462) );
  XNOR U17216 ( .A(p_input[1864]), .B(n17463), .Z(n16632) );
  AND U17217 ( .A(n434), .B(n17464), .Z(n17463) );
  XOR U17218 ( .A(p_input[1896]), .B(p_input[1864]), .Z(n17464) );
  XNOR U17219 ( .A(n16629), .B(n17459), .Z(n17461) );
  XOR U17220 ( .A(n17465), .B(n17466), .Z(n16629) );
  AND U17221 ( .A(n431), .B(n17467), .Z(n17466) );
  XOR U17222 ( .A(p_input[1832]), .B(p_input[1800]), .Z(n17467) );
  XOR U17223 ( .A(n17468), .B(n17469), .Z(n17459) );
  AND U17224 ( .A(n17470), .B(n17471), .Z(n17469) );
  XOR U17225 ( .A(n17468), .B(n16644), .Z(n17471) );
  XNOR U17226 ( .A(p_input[1863]), .B(n17472), .Z(n16644) );
  AND U17227 ( .A(n434), .B(n17473), .Z(n17472) );
  XOR U17228 ( .A(p_input[1895]), .B(p_input[1863]), .Z(n17473) );
  XNOR U17229 ( .A(n16641), .B(n17468), .Z(n17470) );
  XOR U17230 ( .A(n17474), .B(n17475), .Z(n16641) );
  AND U17231 ( .A(n431), .B(n17476), .Z(n17475) );
  XOR U17232 ( .A(p_input[1831]), .B(p_input[1799]), .Z(n17476) );
  XOR U17233 ( .A(n17477), .B(n17478), .Z(n17468) );
  AND U17234 ( .A(n17479), .B(n17480), .Z(n17478) );
  XOR U17235 ( .A(n17477), .B(n16656), .Z(n17480) );
  XNOR U17236 ( .A(p_input[1862]), .B(n17481), .Z(n16656) );
  AND U17237 ( .A(n434), .B(n17482), .Z(n17481) );
  XOR U17238 ( .A(p_input[1894]), .B(p_input[1862]), .Z(n17482) );
  XNOR U17239 ( .A(n16653), .B(n17477), .Z(n17479) );
  XOR U17240 ( .A(n17483), .B(n17484), .Z(n16653) );
  AND U17241 ( .A(n431), .B(n17485), .Z(n17484) );
  XOR U17242 ( .A(p_input[1830]), .B(p_input[1798]), .Z(n17485) );
  XOR U17243 ( .A(n17486), .B(n17487), .Z(n17477) );
  AND U17244 ( .A(n17488), .B(n17489), .Z(n17487) );
  XOR U17245 ( .A(n17486), .B(n16668), .Z(n17489) );
  XNOR U17246 ( .A(p_input[1861]), .B(n17490), .Z(n16668) );
  AND U17247 ( .A(n434), .B(n17491), .Z(n17490) );
  XOR U17248 ( .A(p_input[1893]), .B(p_input[1861]), .Z(n17491) );
  XNOR U17249 ( .A(n16665), .B(n17486), .Z(n17488) );
  XOR U17250 ( .A(n17492), .B(n17493), .Z(n16665) );
  AND U17251 ( .A(n431), .B(n17494), .Z(n17493) );
  XOR U17252 ( .A(p_input[1829]), .B(p_input[1797]), .Z(n17494) );
  XOR U17253 ( .A(n17495), .B(n17496), .Z(n17486) );
  AND U17254 ( .A(n17497), .B(n17498), .Z(n17496) );
  XOR U17255 ( .A(n17495), .B(n16680), .Z(n17498) );
  XNOR U17256 ( .A(p_input[1860]), .B(n17499), .Z(n16680) );
  AND U17257 ( .A(n434), .B(n17500), .Z(n17499) );
  XOR U17258 ( .A(p_input[1892]), .B(p_input[1860]), .Z(n17500) );
  XNOR U17259 ( .A(n16677), .B(n17495), .Z(n17497) );
  XOR U17260 ( .A(n17501), .B(n17502), .Z(n16677) );
  AND U17261 ( .A(n431), .B(n17503), .Z(n17502) );
  XOR U17262 ( .A(p_input[1828]), .B(p_input[1796]), .Z(n17503) );
  XOR U17263 ( .A(n17504), .B(n17505), .Z(n17495) );
  AND U17264 ( .A(n17506), .B(n17507), .Z(n17505) );
  XOR U17265 ( .A(n17504), .B(n16692), .Z(n17507) );
  XNOR U17266 ( .A(p_input[1859]), .B(n17508), .Z(n16692) );
  AND U17267 ( .A(n434), .B(n17509), .Z(n17508) );
  XOR U17268 ( .A(p_input[1891]), .B(p_input[1859]), .Z(n17509) );
  XNOR U17269 ( .A(n16689), .B(n17504), .Z(n17506) );
  XOR U17270 ( .A(n17510), .B(n17511), .Z(n16689) );
  AND U17271 ( .A(n431), .B(n17512), .Z(n17511) );
  XOR U17272 ( .A(p_input[1827]), .B(p_input[1795]), .Z(n17512) );
  XOR U17273 ( .A(n17513), .B(n17514), .Z(n17504) );
  AND U17274 ( .A(n17515), .B(n17516), .Z(n17514) );
  XOR U17275 ( .A(n16704), .B(n17513), .Z(n17516) );
  XNOR U17276 ( .A(p_input[1858]), .B(n17517), .Z(n16704) );
  AND U17277 ( .A(n434), .B(n17518), .Z(n17517) );
  XOR U17278 ( .A(p_input[1890]), .B(p_input[1858]), .Z(n17518) );
  XNOR U17279 ( .A(n17513), .B(n16701), .Z(n17515) );
  XOR U17280 ( .A(n17519), .B(n17520), .Z(n16701) );
  AND U17281 ( .A(n431), .B(n17521), .Z(n17520) );
  XOR U17282 ( .A(p_input[1826]), .B(p_input[1794]), .Z(n17521) );
  XOR U17283 ( .A(n17522), .B(n17523), .Z(n17513) );
  AND U17284 ( .A(n17524), .B(n17525), .Z(n17523) );
  XNOR U17285 ( .A(n17526), .B(n16717), .Z(n17525) );
  XNOR U17286 ( .A(p_input[1857]), .B(n17527), .Z(n16717) );
  AND U17287 ( .A(n434), .B(n17528), .Z(n17527) );
  XNOR U17288 ( .A(p_input[1889]), .B(n17529), .Z(n17528) );
  IV U17289 ( .A(p_input[1857]), .Z(n17529) );
  XNOR U17290 ( .A(n16714), .B(n17522), .Z(n17524) );
  XNOR U17291 ( .A(p_input[1793]), .B(n17530), .Z(n16714) );
  AND U17292 ( .A(n431), .B(n17531), .Z(n17530) );
  XOR U17293 ( .A(p_input[1825]), .B(p_input[1793]), .Z(n17531) );
  IV U17294 ( .A(n17526), .Z(n17522) );
  AND U17295 ( .A(n17252), .B(n17255), .Z(n17526) );
  XOR U17296 ( .A(p_input[1856]), .B(n17532), .Z(n17255) );
  AND U17297 ( .A(n434), .B(n17533), .Z(n17532) );
  XOR U17298 ( .A(p_input[1888]), .B(p_input[1856]), .Z(n17533) );
  XOR U17299 ( .A(n17534), .B(n17535), .Z(n434) );
  AND U17300 ( .A(n17536), .B(n17537), .Z(n17535) );
  XNOR U17301 ( .A(p_input[1919]), .B(n17534), .Z(n17537) );
  XOR U17302 ( .A(n17534), .B(p_input[1887]), .Z(n17536) );
  XOR U17303 ( .A(n17538), .B(n17539), .Z(n17534) );
  AND U17304 ( .A(n17540), .B(n17541), .Z(n17539) );
  XNOR U17305 ( .A(p_input[1918]), .B(n17538), .Z(n17541) );
  XOR U17306 ( .A(n17538), .B(p_input[1886]), .Z(n17540) );
  XOR U17307 ( .A(n17542), .B(n17543), .Z(n17538) );
  AND U17308 ( .A(n17544), .B(n17545), .Z(n17543) );
  XNOR U17309 ( .A(p_input[1917]), .B(n17542), .Z(n17545) );
  XOR U17310 ( .A(n17542), .B(p_input[1885]), .Z(n17544) );
  XOR U17311 ( .A(n17546), .B(n17547), .Z(n17542) );
  AND U17312 ( .A(n17548), .B(n17549), .Z(n17547) );
  XNOR U17313 ( .A(p_input[1916]), .B(n17546), .Z(n17549) );
  XOR U17314 ( .A(n17546), .B(p_input[1884]), .Z(n17548) );
  XOR U17315 ( .A(n17550), .B(n17551), .Z(n17546) );
  AND U17316 ( .A(n17552), .B(n17553), .Z(n17551) );
  XNOR U17317 ( .A(p_input[1915]), .B(n17550), .Z(n17553) );
  XOR U17318 ( .A(n17550), .B(p_input[1883]), .Z(n17552) );
  XOR U17319 ( .A(n17554), .B(n17555), .Z(n17550) );
  AND U17320 ( .A(n17556), .B(n17557), .Z(n17555) );
  XNOR U17321 ( .A(p_input[1914]), .B(n17554), .Z(n17557) );
  XOR U17322 ( .A(n17554), .B(p_input[1882]), .Z(n17556) );
  XOR U17323 ( .A(n17558), .B(n17559), .Z(n17554) );
  AND U17324 ( .A(n17560), .B(n17561), .Z(n17559) );
  XNOR U17325 ( .A(p_input[1913]), .B(n17558), .Z(n17561) );
  XOR U17326 ( .A(n17558), .B(p_input[1881]), .Z(n17560) );
  XOR U17327 ( .A(n17562), .B(n17563), .Z(n17558) );
  AND U17328 ( .A(n17564), .B(n17565), .Z(n17563) );
  XNOR U17329 ( .A(p_input[1912]), .B(n17562), .Z(n17565) );
  XOR U17330 ( .A(n17562), .B(p_input[1880]), .Z(n17564) );
  XOR U17331 ( .A(n17566), .B(n17567), .Z(n17562) );
  AND U17332 ( .A(n17568), .B(n17569), .Z(n17567) );
  XNOR U17333 ( .A(p_input[1911]), .B(n17566), .Z(n17569) );
  XOR U17334 ( .A(n17566), .B(p_input[1879]), .Z(n17568) );
  XOR U17335 ( .A(n17570), .B(n17571), .Z(n17566) );
  AND U17336 ( .A(n17572), .B(n17573), .Z(n17571) );
  XNOR U17337 ( .A(p_input[1910]), .B(n17570), .Z(n17573) );
  XOR U17338 ( .A(n17570), .B(p_input[1878]), .Z(n17572) );
  XOR U17339 ( .A(n17574), .B(n17575), .Z(n17570) );
  AND U17340 ( .A(n17576), .B(n17577), .Z(n17575) );
  XNOR U17341 ( .A(p_input[1909]), .B(n17574), .Z(n17577) );
  XOR U17342 ( .A(n17574), .B(p_input[1877]), .Z(n17576) );
  XOR U17343 ( .A(n17578), .B(n17579), .Z(n17574) );
  AND U17344 ( .A(n17580), .B(n17581), .Z(n17579) );
  XNOR U17345 ( .A(p_input[1908]), .B(n17578), .Z(n17581) );
  XOR U17346 ( .A(n17578), .B(p_input[1876]), .Z(n17580) );
  XOR U17347 ( .A(n17582), .B(n17583), .Z(n17578) );
  AND U17348 ( .A(n17584), .B(n17585), .Z(n17583) );
  XNOR U17349 ( .A(p_input[1907]), .B(n17582), .Z(n17585) );
  XOR U17350 ( .A(n17582), .B(p_input[1875]), .Z(n17584) );
  XOR U17351 ( .A(n17586), .B(n17587), .Z(n17582) );
  AND U17352 ( .A(n17588), .B(n17589), .Z(n17587) );
  XNOR U17353 ( .A(p_input[1906]), .B(n17586), .Z(n17589) );
  XOR U17354 ( .A(n17586), .B(p_input[1874]), .Z(n17588) );
  XOR U17355 ( .A(n17590), .B(n17591), .Z(n17586) );
  AND U17356 ( .A(n17592), .B(n17593), .Z(n17591) );
  XNOR U17357 ( .A(p_input[1905]), .B(n17590), .Z(n17593) );
  XOR U17358 ( .A(n17590), .B(p_input[1873]), .Z(n17592) );
  XOR U17359 ( .A(n17594), .B(n17595), .Z(n17590) );
  AND U17360 ( .A(n17596), .B(n17597), .Z(n17595) );
  XNOR U17361 ( .A(p_input[1904]), .B(n17594), .Z(n17597) );
  XOR U17362 ( .A(n17594), .B(p_input[1872]), .Z(n17596) );
  XOR U17363 ( .A(n17598), .B(n17599), .Z(n17594) );
  AND U17364 ( .A(n17600), .B(n17601), .Z(n17599) );
  XNOR U17365 ( .A(p_input[1903]), .B(n17598), .Z(n17601) );
  XOR U17366 ( .A(n17598), .B(p_input[1871]), .Z(n17600) );
  XOR U17367 ( .A(n17602), .B(n17603), .Z(n17598) );
  AND U17368 ( .A(n17604), .B(n17605), .Z(n17603) );
  XNOR U17369 ( .A(p_input[1902]), .B(n17602), .Z(n17605) );
  XOR U17370 ( .A(n17602), .B(p_input[1870]), .Z(n17604) );
  XOR U17371 ( .A(n17606), .B(n17607), .Z(n17602) );
  AND U17372 ( .A(n17608), .B(n17609), .Z(n17607) );
  XNOR U17373 ( .A(p_input[1901]), .B(n17606), .Z(n17609) );
  XOR U17374 ( .A(n17606), .B(p_input[1869]), .Z(n17608) );
  XOR U17375 ( .A(n17610), .B(n17611), .Z(n17606) );
  AND U17376 ( .A(n17612), .B(n17613), .Z(n17611) );
  XNOR U17377 ( .A(p_input[1900]), .B(n17610), .Z(n17613) );
  XOR U17378 ( .A(n17610), .B(p_input[1868]), .Z(n17612) );
  XOR U17379 ( .A(n17614), .B(n17615), .Z(n17610) );
  AND U17380 ( .A(n17616), .B(n17617), .Z(n17615) );
  XNOR U17381 ( .A(p_input[1899]), .B(n17614), .Z(n17617) );
  XOR U17382 ( .A(n17614), .B(p_input[1867]), .Z(n17616) );
  XOR U17383 ( .A(n17618), .B(n17619), .Z(n17614) );
  AND U17384 ( .A(n17620), .B(n17621), .Z(n17619) );
  XNOR U17385 ( .A(p_input[1898]), .B(n17618), .Z(n17621) );
  XOR U17386 ( .A(n17618), .B(p_input[1866]), .Z(n17620) );
  XOR U17387 ( .A(n17622), .B(n17623), .Z(n17618) );
  AND U17388 ( .A(n17624), .B(n17625), .Z(n17623) );
  XNOR U17389 ( .A(p_input[1897]), .B(n17622), .Z(n17625) );
  XOR U17390 ( .A(n17622), .B(p_input[1865]), .Z(n17624) );
  XOR U17391 ( .A(n17626), .B(n17627), .Z(n17622) );
  AND U17392 ( .A(n17628), .B(n17629), .Z(n17627) );
  XNOR U17393 ( .A(p_input[1896]), .B(n17626), .Z(n17629) );
  XOR U17394 ( .A(n17626), .B(p_input[1864]), .Z(n17628) );
  XOR U17395 ( .A(n17630), .B(n17631), .Z(n17626) );
  AND U17396 ( .A(n17632), .B(n17633), .Z(n17631) );
  XNOR U17397 ( .A(p_input[1895]), .B(n17630), .Z(n17633) );
  XOR U17398 ( .A(n17630), .B(p_input[1863]), .Z(n17632) );
  XOR U17399 ( .A(n17634), .B(n17635), .Z(n17630) );
  AND U17400 ( .A(n17636), .B(n17637), .Z(n17635) );
  XNOR U17401 ( .A(p_input[1894]), .B(n17634), .Z(n17637) );
  XOR U17402 ( .A(n17634), .B(p_input[1862]), .Z(n17636) );
  XOR U17403 ( .A(n17638), .B(n17639), .Z(n17634) );
  AND U17404 ( .A(n17640), .B(n17641), .Z(n17639) );
  XNOR U17405 ( .A(p_input[1893]), .B(n17638), .Z(n17641) );
  XOR U17406 ( .A(n17638), .B(p_input[1861]), .Z(n17640) );
  XOR U17407 ( .A(n17642), .B(n17643), .Z(n17638) );
  AND U17408 ( .A(n17644), .B(n17645), .Z(n17643) );
  XNOR U17409 ( .A(p_input[1892]), .B(n17642), .Z(n17645) );
  XOR U17410 ( .A(n17642), .B(p_input[1860]), .Z(n17644) );
  XOR U17411 ( .A(n17646), .B(n17647), .Z(n17642) );
  AND U17412 ( .A(n17648), .B(n17649), .Z(n17647) );
  XNOR U17413 ( .A(p_input[1891]), .B(n17646), .Z(n17649) );
  XOR U17414 ( .A(n17646), .B(p_input[1859]), .Z(n17648) );
  XOR U17415 ( .A(n17650), .B(n17651), .Z(n17646) );
  AND U17416 ( .A(n17652), .B(n17653), .Z(n17651) );
  XNOR U17417 ( .A(p_input[1890]), .B(n17650), .Z(n17653) );
  XOR U17418 ( .A(n17650), .B(p_input[1858]), .Z(n17652) );
  XNOR U17419 ( .A(n17654), .B(n17655), .Z(n17650) );
  AND U17420 ( .A(n17656), .B(n17657), .Z(n17655) );
  XOR U17421 ( .A(p_input[1889]), .B(n17654), .Z(n17657) );
  XNOR U17422 ( .A(p_input[1857]), .B(n17654), .Z(n17656) );
  AND U17423 ( .A(p_input[1888]), .B(n17658), .Z(n17654) );
  IV U17424 ( .A(p_input[1856]), .Z(n17658) );
  XNOR U17425 ( .A(p_input[1792]), .B(n17659), .Z(n17252) );
  AND U17426 ( .A(n431), .B(n17660), .Z(n17659) );
  XOR U17427 ( .A(p_input[1824]), .B(p_input[1792]), .Z(n17660) );
  XOR U17428 ( .A(n17661), .B(n17662), .Z(n431) );
  AND U17429 ( .A(n17663), .B(n17664), .Z(n17662) );
  XNOR U17430 ( .A(p_input[1855]), .B(n17661), .Z(n17664) );
  XOR U17431 ( .A(n17661), .B(p_input[1823]), .Z(n17663) );
  XOR U17432 ( .A(n17665), .B(n17666), .Z(n17661) );
  AND U17433 ( .A(n17667), .B(n17668), .Z(n17666) );
  XNOR U17434 ( .A(p_input[1854]), .B(n17665), .Z(n17668) );
  XNOR U17435 ( .A(n17665), .B(n17267), .Z(n17667) );
  IV U17436 ( .A(p_input[1822]), .Z(n17267) );
  XOR U17437 ( .A(n17669), .B(n17670), .Z(n17665) );
  AND U17438 ( .A(n17671), .B(n17672), .Z(n17670) );
  XNOR U17439 ( .A(p_input[1853]), .B(n17669), .Z(n17672) );
  XNOR U17440 ( .A(n17669), .B(n17276), .Z(n17671) );
  IV U17441 ( .A(p_input[1821]), .Z(n17276) );
  XOR U17442 ( .A(n17673), .B(n17674), .Z(n17669) );
  AND U17443 ( .A(n17675), .B(n17676), .Z(n17674) );
  XNOR U17444 ( .A(p_input[1852]), .B(n17673), .Z(n17676) );
  XNOR U17445 ( .A(n17673), .B(n17285), .Z(n17675) );
  IV U17446 ( .A(p_input[1820]), .Z(n17285) );
  XOR U17447 ( .A(n17677), .B(n17678), .Z(n17673) );
  AND U17448 ( .A(n17679), .B(n17680), .Z(n17678) );
  XNOR U17449 ( .A(p_input[1851]), .B(n17677), .Z(n17680) );
  XNOR U17450 ( .A(n17677), .B(n17294), .Z(n17679) );
  IV U17451 ( .A(p_input[1819]), .Z(n17294) );
  XOR U17452 ( .A(n17681), .B(n17682), .Z(n17677) );
  AND U17453 ( .A(n17683), .B(n17684), .Z(n17682) );
  XNOR U17454 ( .A(p_input[1850]), .B(n17681), .Z(n17684) );
  XNOR U17455 ( .A(n17681), .B(n17303), .Z(n17683) );
  IV U17456 ( .A(p_input[1818]), .Z(n17303) );
  XOR U17457 ( .A(n17685), .B(n17686), .Z(n17681) );
  AND U17458 ( .A(n17687), .B(n17688), .Z(n17686) );
  XNOR U17459 ( .A(p_input[1849]), .B(n17685), .Z(n17688) );
  XNOR U17460 ( .A(n17685), .B(n17312), .Z(n17687) );
  IV U17461 ( .A(p_input[1817]), .Z(n17312) );
  XOR U17462 ( .A(n17689), .B(n17690), .Z(n17685) );
  AND U17463 ( .A(n17691), .B(n17692), .Z(n17690) );
  XNOR U17464 ( .A(p_input[1848]), .B(n17689), .Z(n17692) );
  XNOR U17465 ( .A(n17689), .B(n17321), .Z(n17691) );
  IV U17466 ( .A(p_input[1816]), .Z(n17321) );
  XOR U17467 ( .A(n17693), .B(n17694), .Z(n17689) );
  AND U17468 ( .A(n17695), .B(n17696), .Z(n17694) );
  XNOR U17469 ( .A(p_input[1847]), .B(n17693), .Z(n17696) );
  XNOR U17470 ( .A(n17693), .B(n17330), .Z(n17695) );
  IV U17471 ( .A(p_input[1815]), .Z(n17330) );
  XOR U17472 ( .A(n17697), .B(n17698), .Z(n17693) );
  AND U17473 ( .A(n17699), .B(n17700), .Z(n17698) );
  XNOR U17474 ( .A(p_input[1846]), .B(n17697), .Z(n17700) );
  XNOR U17475 ( .A(n17697), .B(n17339), .Z(n17699) );
  IV U17476 ( .A(p_input[1814]), .Z(n17339) );
  XOR U17477 ( .A(n17701), .B(n17702), .Z(n17697) );
  AND U17478 ( .A(n17703), .B(n17704), .Z(n17702) );
  XNOR U17479 ( .A(p_input[1845]), .B(n17701), .Z(n17704) );
  XNOR U17480 ( .A(n17701), .B(n17348), .Z(n17703) );
  IV U17481 ( .A(p_input[1813]), .Z(n17348) );
  XOR U17482 ( .A(n17705), .B(n17706), .Z(n17701) );
  AND U17483 ( .A(n17707), .B(n17708), .Z(n17706) );
  XNOR U17484 ( .A(p_input[1844]), .B(n17705), .Z(n17708) );
  XNOR U17485 ( .A(n17705), .B(n17357), .Z(n17707) );
  IV U17486 ( .A(p_input[1812]), .Z(n17357) );
  XOR U17487 ( .A(n17709), .B(n17710), .Z(n17705) );
  AND U17488 ( .A(n17711), .B(n17712), .Z(n17710) );
  XNOR U17489 ( .A(p_input[1843]), .B(n17709), .Z(n17712) );
  XNOR U17490 ( .A(n17709), .B(n17366), .Z(n17711) );
  IV U17491 ( .A(p_input[1811]), .Z(n17366) );
  XOR U17492 ( .A(n17713), .B(n17714), .Z(n17709) );
  AND U17493 ( .A(n17715), .B(n17716), .Z(n17714) );
  XNOR U17494 ( .A(p_input[1842]), .B(n17713), .Z(n17716) );
  XNOR U17495 ( .A(n17713), .B(n17375), .Z(n17715) );
  IV U17496 ( .A(p_input[1810]), .Z(n17375) );
  XOR U17497 ( .A(n17717), .B(n17718), .Z(n17713) );
  AND U17498 ( .A(n17719), .B(n17720), .Z(n17718) );
  XNOR U17499 ( .A(p_input[1841]), .B(n17717), .Z(n17720) );
  XNOR U17500 ( .A(n17717), .B(n17384), .Z(n17719) );
  IV U17501 ( .A(p_input[1809]), .Z(n17384) );
  XOR U17502 ( .A(n17721), .B(n17722), .Z(n17717) );
  AND U17503 ( .A(n17723), .B(n17724), .Z(n17722) );
  XNOR U17504 ( .A(p_input[1840]), .B(n17721), .Z(n17724) );
  XNOR U17505 ( .A(n17721), .B(n17393), .Z(n17723) );
  IV U17506 ( .A(p_input[1808]), .Z(n17393) );
  XOR U17507 ( .A(n17725), .B(n17726), .Z(n17721) );
  AND U17508 ( .A(n17727), .B(n17728), .Z(n17726) );
  XNOR U17509 ( .A(p_input[1839]), .B(n17725), .Z(n17728) );
  XNOR U17510 ( .A(n17725), .B(n17402), .Z(n17727) );
  IV U17511 ( .A(p_input[1807]), .Z(n17402) );
  XOR U17512 ( .A(n17729), .B(n17730), .Z(n17725) );
  AND U17513 ( .A(n17731), .B(n17732), .Z(n17730) );
  XNOR U17514 ( .A(p_input[1838]), .B(n17729), .Z(n17732) );
  XNOR U17515 ( .A(n17729), .B(n17411), .Z(n17731) );
  IV U17516 ( .A(p_input[1806]), .Z(n17411) );
  XOR U17517 ( .A(n17733), .B(n17734), .Z(n17729) );
  AND U17518 ( .A(n17735), .B(n17736), .Z(n17734) );
  XNOR U17519 ( .A(p_input[1837]), .B(n17733), .Z(n17736) );
  XNOR U17520 ( .A(n17733), .B(n17420), .Z(n17735) );
  IV U17521 ( .A(p_input[1805]), .Z(n17420) );
  XOR U17522 ( .A(n17737), .B(n17738), .Z(n17733) );
  AND U17523 ( .A(n17739), .B(n17740), .Z(n17738) );
  XNOR U17524 ( .A(p_input[1836]), .B(n17737), .Z(n17740) );
  XNOR U17525 ( .A(n17737), .B(n17429), .Z(n17739) );
  IV U17526 ( .A(p_input[1804]), .Z(n17429) );
  XOR U17527 ( .A(n17741), .B(n17742), .Z(n17737) );
  AND U17528 ( .A(n17743), .B(n17744), .Z(n17742) );
  XNOR U17529 ( .A(p_input[1835]), .B(n17741), .Z(n17744) );
  XNOR U17530 ( .A(n17741), .B(n17438), .Z(n17743) );
  IV U17531 ( .A(p_input[1803]), .Z(n17438) );
  XOR U17532 ( .A(n17745), .B(n17746), .Z(n17741) );
  AND U17533 ( .A(n17747), .B(n17748), .Z(n17746) );
  XNOR U17534 ( .A(p_input[1834]), .B(n17745), .Z(n17748) );
  XNOR U17535 ( .A(n17745), .B(n17447), .Z(n17747) );
  IV U17536 ( .A(p_input[1802]), .Z(n17447) );
  XOR U17537 ( .A(n17749), .B(n17750), .Z(n17745) );
  AND U17538 ( .A(n17751), .B(n17752), .Z(n17750) );
  XNOR U17539 ( .A(p_input[1833]), .B(n17749), .Z(n17752) );
  XNOR U17540 ( .A(n17749), .B(n17456), .Z(n17751) );
  IV U17541 ( .A(p_input[1801]), .Z(n17456) );
  XOR U17542 ( .A(n17753), .B(n17754), .Z(n17749) );
  AND U17543 ( .A(n17755), .B(n17756), .Z(n17754) );
  XNOR U17544 ( .A(p_input[1832]), .B(n17753), .Z(n17756) );
  XNOR U17545 ( .A(n17753), .B(n17465), .Z(n17755) );
  IV U17546 ( .A(p_input[1800]), .Z(n17465) );
  XOR U17547 ( .A(n17757), .B(n17758), .Z(n17753) );
  AND U17548 ( .A(n17759), .B(n17760), .Z(n17758) );
  XNOR U17549 ( .A(p_input[1831]), .B(n17757), .Z(n17760) );
  XNOR U17550 ( .A(n17757), .B(n17474), .Z(n17759) );
  IV U17551 ( .A(p_input[1799]), .Z(n17474) );
  XOR U17552 ( .A(n17761), .B(n17762), .Z(n17757) );
  AND U17553 ( .A(n17763), .B(n17764), .Z(n17762) );
  XNOR U17554 ( .A(p_input[1830]), .B(n17761), .Z(n17764) );
  XNOR U17555 ( .A(n17761), .B(n17483), .Z(n17763) );
  IV U17556 ( .A(p_input[1798]), .Z(n17483) );
  XOR U17557 ( .A(n17765), .B(n17766), .Z(n17761) );
  AND U17558 ( .A(n17767), .B(n17768), .Z(n17766) );
  XNOR U17559 ( .A(p_input[1829]), .B(n17765), .Z(n17768) );
  XNOR U17560 ( .A(n17765), .B(n17492), .Z(n17767) );
  IV U17561 ( .A(p_input[1797]), .Z(n17492) );
  XOR U17562 ( .A(n17769), .B(n17770), .Z(n17765) );
  AND U17563 ( .A(n17771), .B(n17772), .Z(n17770) );
  XNOR U17564 ( .A(p_input[1828]), .B(n17769), .Z(n17772) );
  XNOR U17565 ( .A(n17769), .B(n17501), .Z(n17771) );
  IV U17566 ( .A(p_input[1796]), .Z(n17501) );
  XOR U17567 ( .A(n17773), .B(n17774), .Z(n17769) );
  AND U17568 ( .A(n17775), .B(n17776), .Z(n17774) );
  XNOR U17569 ( .A(p_input[1827]), .B(n17773), .Z(n17776) );
  XNOR U17570 ( .A(n17773), .B(n17510), .Z(n17775) );
  IV U17571 ( .A(p_input[1795]), .Z(n17510) );
  XOR U17572 ( .A(n17777), .B(n17778), .Z(n17773) );
  AND U17573 ( .A(n17779), .B(n17780), .Z(n17778) );
  XNOR U17574 ( .A(p_input[1826]), .B(n17777), .Z(n17780) );
  XNOR U17575 ( .A(n17777), .B(n17519), .Z(n17779) );
  IV U17576 ( .A(p_input[1794]), .Z(n17519) );
  XNOR U17577 ( .A(n17781), .B(n17782), .Z(n17777) );
  AND U17578 ( .A(n17783), .B(n17784), .Z(n17782) );
  XOR U17579 ( .A(p_input[1825]), .B(n17781), .Z(n17784) );
  XNOR U17580 ( .A(p_input[1793]), .B(n17781), .Z(n17783) );
  AND U17581 ( .A(p_input[1824]), .B(n17785), .Z(n17781) );
  IV U17582 ( .A(p_input[1792]), .Z(n17785) );
  XOR U17583 ( .A(n17786), .B(n17787), .Z(n15964) );
  AND U17584 ( .A(n516), .B(n17788), .Z(n17787) );
  XNOR U17585 ( .A(n17789), .B(n17786), .Z(n17788) );
  XOR U17586 ( .A(n17790), .B(n17791), .Z(n516) );
  AND U17587 ( .A(n17792), .B(n17793), .Z(n17791) );
  XOR U17588 ( .A(n17790), .B(n15979), .Z(n17793) );
  XNOR U17589 ( .A(n17794), .B(n17795), .Z(n15979) );
  AND U17590 ( .A(n17796), .B(n370), .Z(n17795) );
  AND U17591 ( .A(n17794), .B(n17797), .Z(n17796) );
  XNOR U17592 ( .A(n15976), .B(n17790), .Z(n17792) );
  XOR U17593 ( .A(n17798), .B(n17799), .Z(n15976) );
  AND U17594 ( .A(n17800), .B(n367), .Z(n17799) );
  NOR U17595 ( .A(n17798), .B(n17801), .Z(n17800) );
  XOR U17596 ( .A(n17802), .B(n17803), .Z(n17790) );
  AND U17597 ( .A(n17804), .B(n17805), .Z(n17803) );
  XOR U17598 ( .A(n17802), .B(n15991), .Z(n17805) );
  XOR U17599 ( .A(n17806), .B(n17807), .Z(n15991) );
  AND U17600 ( .A(n370), .B(n17808), .Z(n17807) );
  XOR U17601 ( .A(n17809), .B(n17806), .Z(n17808) );
  XNOR U17602 ( .A(n15988), .B(n17802), .Z(n17804) );
  XOR U17603 ( .A(n17810), .B(n17811), .Z(n15988) );
  AND U17604 ( .A(n367), .B(n17812), .Z(n17811) );
  XOR U17605 ( .A(n17813), .B(n17810), .Z(n17812) );
  XOR U17606 ( .A(n17814), .B(n17815), .Z(n17802) );
  AND U17607 ( .A(n17816), .B(n17817), .Z(n17815) );
  XOR U17608 ( .A(n17814), .B(n16003), .Z(n17817) );
  XOR U17609 ( .A(n17818), .B(n17819), .Z(n16003) );
  AND U17610 ( .A(n370), .B(n17820), .Z(n17819) );
  XOR U17611 ( .A(n17821), .B(n17818), .Z(n17820) );
  XNOR U17612 ( .A(n16000), .B(n17814), .Z(n17816) );
  XOR U17613 ( .A(n17822), .B(n17823), .Z(n16000) );
  AND U17614 ( .A(n367), .B(n17824), .Z(n17823) );
  XOR U17615 ( .A(n17825), .B(n17822), .Z(n17824) );
  XOR U17616 ( .A(n17826), .B(n17827), .Z(n17814) );
  AND U17617 ( .A(n17828), .B(n17829), .Z(n17827) );
  XOR U17618 ( .A(n17826), .B(n16015), .Z(n17829) );
  XOR U17619 ( .A(n17830), .B(n17831), .Z(n16015) );
  AND U17620 ( .A(n370), .B(n17832), .Z(n17831) );
  XOR U17621 ( .A(n17833), .B(n17830), .Z(n17832) );
  XNOR U17622 ( .A(n16012), .B(n17826), .Z(n17828) );
  XOR U17623 ( .A(n17834), .B(n17835), .Z(n16012) );
  AND U17624 ( .A(n367), .B(n17836), .Z(n17835) );
  XOR U17625 ( .A(n17837), .B(n17834), .Z(n17836) );
  XOR U17626 ( .A(n17838), .B(n17839), .Z(n17826) );
  AND U17627 ( .A(n17840), .B(n17841), .Z(n17839) );
  XOR U17628 ( .A(n17838), .B(n16027), .Z(n17841) );
  XOR U17629 ( .A(n17842), .B(n17843), .Z(n16027) );
  AND U17630 ( .A(n370), .B(n17844), .Z(n17843) );
  XOR U17631 ( .A(n17845), .B(n17842), .Z(n17844) );
  XNOR U17632 ( .A(n16024), .B(n17838), .Z(n17840) );
  XOR U17633 ( .A(n17846), .B(n17847), .Z(n16024) );
  AND U17634 ( .A(n367), .B(n17848), .Z(n17847) );
  XOR U17635 ( .A(n17849), .B(n17846), .Z(n17848) );
  XOR U17636 ( .A(n17850), .B(n17851), .Z(n17838) );
  AND U17637 ( .A(n17852), .B(n17853), .Z(n17851) );
  XOR U17638 ( .A(n17850), .B(n16039), .Z(n17853) );
  XOR U17639 ( .A(n17854), .B(n17855), .Z(n16039) );
  AND U17640 ( .A(n370), .B(n17856), .Z(n17855) );
  XOR U17641 ( .A(n17857), .B(n17854), .Z(n17856) );
  XNOR U17642 ( .A(n16036), .B(n17850), .Z(n17852) );
  XOR U17643 ( .A(n17858), .B(n17859), .Z(n16036) );
  AND U17644 ( .A(n367), .B(n17860), .Z(n17859) );
  XOR U17645 ( .A(n17861), .B(n17858), .Z(n17860) );
  XOR U17646 ( .A(n17862), .B(n17863), .Z(n17850) );
  AND U17647 ( .A(n17864), .B(n17865), .Z(n17863) );
  XOR U17648 ( .A(n17862), .B(n16051), .Z(n17865) );
  XOR U17649 ( .A(n17866), .B(n17867), .Z(n16051) );
  AND U17650 ( .A(n370), .B(n17868), .Z(n17867) );
  XOR U17651 ( .A(n17869), .B(n17866), .Z(n17868) );
  XNOR U17652 ( .A(n16048), .B(n17862), .Z(n17864) );
  XOR U17653 ( .A(n17870), .B(n17871), .Z(n16048) );
  AND U17654 ( .A(n367), .B(n17872), .Z(n17871) );
  XOR U17655 ( .A(n17873), .B(n17870), .Z(n17872) );
  XOR U17656 ( .A(n17874), .B(n17875), .Z(n17862) );
  AND U17657 ( .A(n17876), .B(n17877), .Z(n17875) );
  XOR U17658 ( .A(n17874), .B(n16063), .Z(n17877) );
  XOR U17659 ( .A(n17878), .B(n17879), .Z(n16063) );
  AND U17660 ( .A(n370), .B(n17880), .Z(n17879) );
  XOR U17661 ( .A(n17881), .B(n17878), .Z(n17880) );
  XNOR U17662 ( .A(n16060), .B(n17874), .Z(n17876) );
  XOR U17663 ( .A(n17882), .B(n17883), .Z(n16060) );
  AND U17664 ( .A(n367), .B(n17884), .Z(n17883) );
  XOR U17665 ( .A(n17885), .B(n17882), .Z(n17884) );
  XOR U17666 ( .A(n17886), .B(n17887), .Z(n17874) );
  AND U17667 ( .A(n17888), .B(n17889), .Z(n17887) );
  XOR U17668 ( .A(n17886), .B(n16075), .Z(n17889) );
  XOR U17669 ( .A(n17890), .B(n17891), .Z(n16075) );
  AND U17670 ( .A(n370), .B(n17892), .Z(n17891) );
  XOR U17671 ( .A(n17893), .B(n17890), .Z(n17892) );
  XNOR U17672 ( .A(n16072), .B(n17886), .Z(n17888) );
  XOR U17673 ( .A(n17894), .B(n17895), .Z(n16072) );
  AND U17674 ( .A(n367), .B(n17896), .Z(n17895) );
  XOR U17675 ( .A(n17897), .B(n17894), .Z(n17896) );
  XOR U17676 ( .A(n17898), .B(n17899), .Z(n17886) );
  AND U17677 ( .A(n17900), .B(n17901), .Z(n17899) );
  XOR U17678 ( .A(n17898), .B(n16087), .Z(n17901) );
  XOR U17679 ( .A(n17902), .B(n17903), .Z(n16087) );
  AND U17680 ( .A(n370), .B(n17904), .Z(n17903) );
  XOR U17681 ( .A(n17905), .B(n17902), .Z(n17904) );
  XNOR U17682 ( .A(n16084), .B(n17898), .Z(n17900) );
  XOR U17683 ( .A(n17906), .B(n17907), .Z(n16084) );
  AND U17684 ( .A(n367), .B(n17908), .Z(n17907) );
  XOR U17685 ( .A(n17909), .B(n17906), .Z(n17908) );
  XOR U17686 ( .A(n17910), .B(n17911), .Z(n17898) );
  AND U17687 ( .A(n17912), .B(n17913), .Z(n17911) );
  XOR U17688 ( .A(n17910), .B(n16099), .Z(n17913) );
  XOR U17689 ( .A(n17914), .B(n17915), .Z(n16099) );
  AND U17690 ( .A(n370), .B(n17916), .Z(n17915) );
  XOR U17691 ( .A(n17917), .B(n17914), .Z(n17916) );
  XNOR U17692 ( .A(n16096), .B(n17910), .Z(n17912) );
  XOR U17693 ( .A(n17918), .B(n17919), .Z(n16096) );
  AND U17694 ( .A(n367), .B(n17920), .Z(n17919) );
  XOR U17695 ( .A(n17921), .B(n17918), .Z(n17920) );
  XOR U17696 ( .A(n17922), .B(n17923), .Z(n17910) );
  AND U17697 ( .A(n17924), .B(n17925), .Z(n17923) );
  XOR U17698 ( .A(n17922), .B(n16111), .Z(n17925) );
  XOR U17699 ( .A(n17926), .B(n17927), .Z(n16111) );
  AND U17700 ( .A(n370), .B(n17928), .Z(n17927) );
  XOR U17701 ( .A(n17929), .B(n17926), .Z(n17928) );
  XNOR U17702 ( .A(n16108), .B(n17922), .Z(n17924) );
  XOR U17703 ( .A(n17930), .B(n17931), .Z(n16108) );
  AND U17704 ( .A(n367), .B(n17932), .Z(n17931) );
  XOR U17705 ( .A(n17933), .B(n17930), .Z(n17932) );
  XOR U17706 ( .A(n17934), .B(n17935), .Z(n17922) );
  AND U17707 ( .A(n17936), .B(n17937), .Z(n17935) );
  XOR U17708 ( .A(n17934), .B(n16123), .Z(n17937) );
  XOR U17709 ( .A(n17938), .B(n17939), .Z(n16123) );
  AND U17710 ( .A(n370), .B(n17940), .Z(n17939) );
  XOR U17711 ( .A(n17941), .B(n17938), .Z(n17940) );
  XNOR U17712 ( .A(n16120), .B(n17934), .Z(n17936) );
  XOR U17713 ( .A(n17942), .B(n17943), .Z(n16120) );
  AND U17714 ( .A(n367), .B(n17944), .Z(n17943) );
  XOR U17715 ( .A(n17945), .B(n17942), .Z(n17944) );
  XOR U17716 ( .A(n17946), .B(n17947), .Z(n17934) );
  AND U17717 ( .A(n17948), .B(n17949), .Z(n17947) );
  XOR U17718 ( .A(n17946), .B(n16135), .Z(n17949) );
  XOR U17719 ( .A(n17950), .B(n17951), .Z(n16135) );
  AND U17720 ( .A(n370), .B(n17952), .Z(n17951) );
  XOR U17721 ( .A(n17953), .B(n17950), .Z(n17952) );
  XNOR U17722 ( .A(n16132), .B(n17946), .Z(n17948) );
  XOR U17723 ( .A(n17954), .B(n17955), .Z(n16132) );
  AND U17724 ( .A(n367), .B(n17956), .Z(n17955) );
  XOR U17725 ( .A(n17957), .B(n17954), .Z(n17956) );
  XOR U17726 ( .A(n17958), .B(n17959), .Z(n17946) );
  AND U17727 ( .A(n17960), .B(n17961), .Z(n17959) );
  XOR U17728 ( .A(n17958), .B(n16147), .Z(n17961) );
  XOR U17729 ( .A(n17962), .B(n17963), .Z(n16147) );
  AND U17730 ( .A(n370), .B(n17964), .Z(n17963) );
  XOR U17731 ( .A(n17965), .B(n17962), .Z(n17964) );
  XNOR U17732 ( .A(n16144), .B(n17958), .Z(n17960) );
  XOR U17733 ( .A(n17966), .B(n17967), .Z(n16144) );
  AND U17734 ( .A(n367), .B(n17968), .Z(n17967) );
  XOR U17735 ( .A(n17969), .B(n17966), .Z(n17968) );
  XOR U17736 ( .A(n17970), .B(n17971), .Z(n17958) );
  AND U17737 ( .A(n17972), .B(n17973), .Z(n17971) );
  XOR U17738 ( .A(n17970), .B(n16159), .Z(n17973) );
  XOR U17739 ( .A(n17974), .B(n17975), .Z(n16159) );
  AND U17740 ( .A(n370), .B(n17976), .Z(n17975) );
  XOR U17741 ( .A(n17977), .B(n17974), .Z(n17976) );
  XNOR U17742 ( .A(n16156), .B(n17970), .Z(n17972) );
  XOR U17743 ( .A(n17978), .B(n17979), .Z(n16156) );
  AND U17744 ( .A(n367), .B(n17980), .Z(n17979) );
  XOR U17745 ( .A(n17981), .B(n17978), .Z(n17980) );
  XOR U17746 ( .A(n17982), .B(n17983), .Z(n17970) );
  AND U17747 ( .A(n17984), .B(n17985), .Z(n17983) );
  XOR U17748 ( .A(n17982), .B(n16171), .Z(n17985) );
  XOR U17749 ( .A(n17986), .B(n17987), .Z(n16171) );
  AND U17750 ( .A(n370), .B(n17988), .Z(n17987) );
  XOR U17751 ( .A(n17989), .B(n17986), .Z(n17988) );
  XNOR U17752 ( .A(n16168), .B(n17982), .Z(n17984) );
  XOR U17753 ( .A(n17990), .B(n17991), .Z(n16168) );
  AND U17754 ( .A(n367), .B(n17992), .Z(n17991) );
  XOR U17755 ( .A(n17993), .B(n17990), .Z(n17992) );
  XOR U17756 ( .A(n17994), .B(n17995), .Z(n17982) );
  AND U17757 ( .A(n17996), .B(n17997), .Z(n17995) );
  XOR U17758 ( .A(n17994), .B(n16183), .Z(n17997) );
  XOR U17759 ( .A(n17998), .B(n17999), .Z(n16183) );
  AND U17760 ( .A(n370), .B(n18000), .Z(n17999) );
  XOR U17761 ( .A(n18001), .B(n17998), .Z(n18000) );
  XNOR U17762 ( .A(n16180), .B(n17994), .Z(n17996) );
  XOR U17763 ( .A(n18002), .B(n18003), .Z(n16180) );
  AND U17764 ( .A(n367), .B(n18004), .Z(n18003) );
  XOR U17765 ( .A(n18005), .B(n18002), .Z(n18004) );
  XOR U17766 ( .A(n18006), .B(n18007), .Z(n17994) );
  AND U17767 ( .A(n18008), .B(n18009), .Z(n18007) );
  XOR U17768 ( .A(n18006), .B(n16195), .Z(n18009) );
  XOR U17769 ( .A(n18010), .B(n18011), .Z(n16195) );
  AND U17770 ( .A(n370), .B(n18012), .Z(n18011) );
  XOR U17771 ( .A(n18013), .B(n18010), .Z(n18012) );
  XNOR U17772 ( .A(n16192), .B(n18006), .Z(n18008) );
  XOR U17773 ( .A(n18014), .B(n18015), .Z(n16192) );
  AND U17774 ( .A(n367), .B(n18016), .Z(n18015) );
  XOR U17775 ( .A(n18017), .B(n18014), .Z(n18016) );
  XOR U17776 ( .A(n18018), .B(n18019), .Z(n18006) );
  AND U17777 ( .A(n18020), .B(n18021), .Z(n18019) );
  XOR U17778 ( .A(n18018), .B(n16207), .Z(n18021) );
  XOR U17779 ( .A(n18022), .B(n18023), .Z(n16207) );
  AND U17780 ( .A(n370), .B(n18024), .Z(n18023) );
  XOR U17781 ( .A(n18025), .B(n18022), .Z(n18024) );
  XNOR U17782 ( .A(n16204), .B(n18018), .Z(n18020) );
  XOR U17783 ( .A(n18026), .B(n18027), .Z(n16204) );
  AND U17784 ( .A(n367), .B(n18028), .Z(n18027) );
  XOR U17785 ( .A(n18029), .B(n18026), .Z(n18028) );
  XOR U17786 ( .A(n18030), .B(n18031), .Z(n18018) );
  AND U17787 ( .A(n18032), .B(n18033), .Z(n18031) );
  XOR U17788 ( .A(n18030), .B(n16219), .Z(n18033) );
  XOR U17789 ( .A(n18034), .B(n18035), .Z(n16219) );
  AND U17790 ( .A(n370), .B(n18036), .Z(n18035) );
  XOR U17791 ( .A(n18037), .B(n18034), .Z(n18036) );
  XNOR U17792 ( .A(n16216), .B(n18030), .Z(n18032) );
  XOR U17793 ( .A(n18038), .B(n18039), .Z(n16216) );
  AND U17794 ( .A(n367), .B(n18040), .Z(n18039) );
  XOR U17795 ( .A(n18041), .B(n18038), .Z(n18040) );
  XOR U17796 ( .A(n18042), .B(n18043), .Z(n18030) );
  AND U17797 ( .A(n18044), .B(n18045), .Z(n18043) );
  XOR U17798 ( .A(n18042), .B(n16231), .Z(n18045) );
  XOR U17799 ( .A(n18046), .B(n18047), .Z(n16231) );
  AND U17800 ( .A(n370), .B(n18048), .Z(n18047) );
  XOR U17801 ( .A(n18049), .B(n18046), .Z(n18048) );
  XNOR U17802 ( .A(n16228), .B(n18042), .Z(n18044) );
  XOR U17803 ( .A(n18050), .B(n18051), .Z(n16228) );
  AND U17804 ( .A(n367), .B(n18052), .Z(n18051) );
  XOR U17805 ( .A(n18053), .B(n18050), .Z(n18052) );
  XOR U17806 ( .A(n18054), .B(n18055), .Z(n18042) );
  AND U17807 ( .A(n18056), .B(n18057), .Z(n18055) );
  XOR U17808 ( .A(n18054), .B(n16243), .Z(n18057) );
  XOR U17809 ( .A(n18058), .B(n18059), .Z(n16243) );
  AND U17810 ( .A(n370), .B(n18060), .Z(n18059) );
  XOR U17811 ( .A(n18061), .B(n18058), .Z(n18060) );
  XNOR U17812 ( .A(n16240), .B(n18054), .Z(n18056) );
  XOR U17813 ( .A(n18062), .B(n18063), .Z(n16240) );
  AND U17814 ( .A(n367), .B(n18064), .Z(n18063) );
  XOR U17815 ( .A(n18065), .B(n18062), .Z(n18064) );
  XOR U17816 ( .A(n18066), .B(n18067), .Z(n18054) );
  AND U17817 ( .A(n18068), .B(n18069), .Z(n18067) );
  XOR U17818 ( .A(n18066), .B(n16255), .Z(n18069) );
  XOR U17819 ( .A(n18070), .B(n18071), .Z(n16255) );
  AND U17820 ( .A(n370), .B(n18072), .Z(n18071) );
  XOR U17821 ( .A(n18073), .B(n18070), .Z(n18072) );
  XNOR U17822 ( .A(n16252), .B(n18066), .Z(n18068) );
  XOR U17823 ( .A(n18074), .B(n18075), .Z(n16252) );
  AND U17824 ( .A(n367), .B(n18076), .Z(n18075) );
  XOR U17825 ( .A(n18077), .B(n18074), .Z(n18076) );
  XOR U17826 ( .A(n18078), .B(n18079), .Z(n18066) );
  AND U17827 ( .A(n18080), .B(n18081), .Z(n18079) );
  XOR U17828 ( .A(n18078), .B(n16267), .Z(n18081) );
  XOR U17829 ( .A(n18082), .B(n18083), .Z(n16267) );
  AND U17830 ( .A(n370), .B(n18084), .Z(n18083) );
  XOR U17831 ( .A(n18085), .B(n18082), .Z(n18084) );
  XNOR U17832 ( .A(n16264), .B(n18078), .Z(n18080) );
  XOR U17833 ( .A(n18086), .B(n18087), .Z(n16264) );
  AND U17834 ( .A(n367), .B(n18088), .Z(n18087) );
  XOR U17835 ( .A(n18089), .B(n18086), .Z(n18088) );
  XOR U17836 ( .A(n18090), .B(n18091), .Z(n18078) );
  AND U17837 ( .A(n18092), .B(n18093), .Z(n18091) );
  XOR U17838 ( .A(n18090), .B(n16279), .Z(n18093) );
  XOR U17839 ( .A(n18094), .B(n18095), .Z(n16279) );
  AND U17840 ( .A(n370), .B(n18096), .Z(n18095) );
  XOR U17841 ( .A(n18097), .B(n18094), .Z(n18096) );
  XNOR U17842 ( .A(n16276), .B(n18090), .Z(n18092) );
  XOR U17843 ( .A(n18098), .B(n18099), .Z(n16276) );
  AND U17844 ( .A(n367), .B(n18100), .Z(n18099) );
  XOR U17845 ( .A(n18101), .B(n18098), .Z(n18100) );
  XOR U17846 ( .A(n18102), .B(n18103), .Z(n18090) );
  AND U17847 ( .A(n18104), .B(n18105), .Z(n18103) );
  XOR U17848 ( .A(n18102), .B(n16291), .Z(n18105) );
  XOR U17849 ( .A(n18106), .B(n18107), .Z(n16291) );
  AND U17850 ( .A(n370), .B(n18108), .Z(n18107) );
  XOR U17851 ( .A(n18109), .B(n18106), .Z(n18108) );
  XNOR U17852 ( .A(n16288), .B(n18102), .Z(n18104) );
  XOR U17853 ( .A(n18110), .B(n18111), .Z(n16288) );
  AND U17854 ( .A(n367), .B(n18112), .Z(n18111) );
  XOR U17855 ( .A(n18113), .B(n18110), .Z(n18112) );
  XOR U17856 ( .A(n18114), .B(n18115), .Z(n18102) );
  AND U17857 ( .A(n18116), .B(n18117), .Z(n18115) );
  XOR U17858 ( .A(n18114), .B(n16303), .Z(n18117) );
  XOR U17859 ( .A(n18118), .B(n18119), .Z(n16303) );
  AND U17860 ( .A(n370), .B(n18120), .Z(n18119) );
  XOR U17861 ( .A(n18121), .B(n18118), .Z(n18120) );
  XNOR U17862 ( .A(n16300), .B(n18114), .Z(n18116) );
  XOR U17863 ( .A(n18122), .B(n18123), .Z(n16300) );
  AND U17864 ( .A(n367), .B(n18124), .Z(n18123) );
  XOR U17865 ( .A(n18125), .B(n18122), .Z(n18124) );
  XOR U17866 ( .A(n18126), .B(n18127), .Z(n18114) );
  AND U17867 ( .A(n18128), .B(n18129), .Z(n18127) );
  XOR U17868 ( .A(n18126), .B(n16315), .Z(n18129) );
  XOR U17869 ( .A(n18130), .B(n18131), .Z(n16315) );
  AND U17870 ( .A(n370), .B(n18132), .Z(n18131) );
  XOR U17871 ( .A(n18133), .B(n18130), .Z(n18132) );
  XNOR U17872 ( .A(n16312), .B(n18126), .Z(n18128) );
  XOR U17873 ( .A(n18134), .B(n18135), .Z(n16312) );
  AND U17874 ( .A(n367), .B(n18136), .Z(n18135) );
  XOR U17875 ( .A(n18137), .B(n18134), .Z(n18136) );
  XOR U17876 ( .A(n18138), .B(n18139), .Z(n18126) );
  AND U17877 ( .A(n18140), .B(n18141), .Z(n18139) );
  XOR U17878 ( .A(n16327), .B(n18138), .Z(n18141) );
  XOR U17879 ( .A(n18142), .B(n18143), .Z(n16327) );
  AND U17880 ( .A(n370), .B(n18144), .Z(n18143) );
  XOR U17881 ( .A(n18142), .B(n18145), .Z(n18144) );
  XNOR U17882 ( .A(n18138), .B(n16324), .Z(n18140) );
  XOR U17883 ( .A(n18146), .B(n18147), .Z(n16324) );
  AND U17884 ( .A(n367), .B(n18148), .Z(n18147) );
  XOR U17885 ( .A(n18146), .B(n18149), .Z(n18148) );
  XOR U17886 ( .A(n18150), .B(n18151), .Z(n18138) );
  AND U17887 ( .A(n18152), .B(n18153), .Z(n18151) );
  XNOR U17888 ( .A(n18154), .B(n16340), .Z(n18153) );
  XOR U17889 ( .A(n18155), .B(n18156), .Z(n16340) );
  AND U17890 ( .A(n370), .B(n18157), .Z(n18156) );
  XOR U17891 ( .A(n18158), .B(n18155), .Z(n18157) );
  XNOR U17892 ( .A(n16337), .B(n18150), .Z(n18152) );
  XOR U17893 ( .A(n18159), .B(n18160), .Z(n16337) );
  AND U17894 ( .A(n367), .B(n18161), .Z(n18160) );
  XOR U17895 ( .A(n18162), .B(n18159), .Z(n18161) );
  IV U17896 ( .A(n18154), .Z(n18150) );
  AND U17897 ( .A(n17786), .B(n17789), .Z(n18154) );
  XNOR U17898 ( .A(n18163), .B(n18164), .Z(n17789) );
  AND U17899 ( .A(n370), .B(n18165), .Z(n18164) );
  XNOR U17900 ( .A(n18166), .B(n18163), .Z(n18165) );
  XOR U17901 ( .A(n18167), .B(n18168), .Z(n370) );
  AND U17902 ( .A(n18169), .B(n18170), .Z(n18168) );
  XOR U17903 ( .A(n17797), .B(n18167), .Z(n18170) );
  IV U17904 ( .A(n18171), .Z(n17797) );
  AND U17905 ( .A(p_input[1791]), .B(p_input[1759]), .Z(n18171) );
  XOR U17906 ( .A(n18167), .B(n17794), .Z(n18169) );
  AND U17907 ( .A(p_input[1695]), .B(p_input[1727]), .Z(n17794) );
  XOR U17908 ( .A(n18172), .B(n18173), .Z(n18167) );
  AND U17909 ( .A(n18174), .B(n18175), .Z(n18173) );
  XOR U17910 ( .A(n18172), .B(n17809), .Z(n18175) );
  XNOR U17911 ( .A(p_input[1758]), .B(n18176), .Z(n17809) );
  AND U17912 ( .A(n442), .B(n18177), .Z(n18176) );
  XOR U17913 ( .A(p_input[1790]), .B(p_input[1758]), .Z(n18177) );
  XNOR U17914 ( .A(n17806), .B(n18172), .Z(n18174) );
  XOR U17915 ( .A(n18178), .B(n18179), .Z(n17806) );
  AND U17916 ( .A(n440), .B(n18180), .Z(n18179) );
  XOR U17917 ( .A(p_input[1726]), .B(p_input[1694]), .Z(n18180) );
  XOR U17918 ( .A(n18181), .B(n18182), .Z(n18172) );
  AND U17919 ( .A(n18183), .B(n18184), .Z(n18182) );
  XOR U17920 ( .A(n18181), .B(n17821), .Z(n18184) );
  XNOR U17921 ( .A(p_input[1757]), .B(n18185), .Z(n17821) );
  AND U17922 ( .A(n442), .B(n18186), .Z(n18185) );
  XOR U17923 ( .A(p_input[1789]), .B(p_input[1757]), .Z(n18186) );
  XNOR U17924 ( .A(n17818), .B(n18181), .Z(n18183) );
  XOR U17925 ( .A(n18187), .B(n18188), .Z(n17818) );
  AND U17926 ( .A(n440), .B(n18189), .Z(n18188) );
  XOR U17927 ( .A(p_input[1725]), .B(p_input[1693]), .Z(n18189) );
  XOR U17928 ( .A(n18190), .B(n18191), .Z(n18181) );
  AND U17929 ( .A(n18192), .B(n18193), .Z(n18191) );
  XOR U17930 ( .A(n18190), .B(n17833), .Z(n18193) );
  XNOR U17931 ( .A(p_input[1756]), .B(n18194), .Z(n17833) );
  AND U17932 ( .A(n442), .B(n18195), .Z(n18194) );
  XOR U17933 ( .A(p_input[1788]), .B(p_input[1756]), .Z(n18195) );
  XNOR U17934 ( .A(n17830), .B(n18190), .Z(n18192) );
  XOR U17935 ( .A(n18196), .B(n18197), .Z(n17830) );
  AND U17936 ( .A(n440), .B(n18198), .Z(n18197) );
  XOR U17937 ( .A(p_input[1724]), .B(p_input[1692]), .Z(n18198) );
  XOR U17938 ( .A(n18199), .B(n18200), .Z(n18190) );
  AND U17939 ( .A(n18201), .B(n18202), .Z(n18200) );
  XOR U17940 ( .A(n18199), .B(n17845), .Z(n18202) );
  XNOR U17941 ( .A(p_input[1755]), .B(n18203), .Z(n17845) );
  AND U17942 ( .A(n442), .B(n18204), .Z(n18203) );
  XOR U17943 ( .A(p_input[1787]), .B(p_input[1755]), .Z(n18204) );
  XNOR U17944 ( .A(n17842), .B(n18199), .Z(n18201) );
  XOR U17945 ( .A(n18205), .B(n18206), .Z(n17842) );
  AND U17946 ( .A(n440), .B(n18207), .Z(n18206) );
  XOR U17947 ( .A(p_input[1723]), .B(p_input[1691]), .Z(n18207) );
  XOR U17948 ( .A(n18208), .B(n18209), .Z(n18199) );
  AND U17949 ( .A(n18210), .B(n18211), .Z(n18209) );
  XOR U17950 ( .A(n18208), .B(n17857), .Z(n18211) );
  XNOR U17951 ( .A(p_input[1754]), .B(n18212), .Z(n17857) );
  AND U17952 ( .A(n442), .B(n18213), .Z(n18212) );
  XOR U17953 ( .A(p_input[1786]), .B(p_input[1754]), .Z(n18213) );
  XNOR U17954 ( .A(n17854), .B(n18208), .Z(n18210) );
  XOR U17955 ( .A(n18214), .B(n18215), .Z(n17854) );
  AND U17956 ( .A(n440), .B(n18216), .Z(n18215) );
  XOR U17957 ( .A(p_input[1722]), .B(p_input[1690]), .Z(n18216) );
  XOR U17958 ( .A(n18217), .B(n18218), .Z(n18208) );
  AND U17959 ( .A(n18219), .B(n18220), .Z(n18218) );
  XOR U17960 ( .A(n18217), .B(n17869), .Z(n18220) );
  XNOR U17961 ( .A(p_input[1753]), .B(n18221), .Z(n17869) );
  AND U17962 ( .A(n442), .B(n18222), .Z(n18221) );
  XOR U17963 ( .A(p_input[1785]), .B(p_input[1753]), .Z(n18222) );
  XNOR U17964 ( .A(n17866), .B(n18217), .Z(n18219) );
  XOR U17965 ( .A(n18223), .B(n18224), .Z(n17866) );
  AND U17966 ( .A(n440), .B(n18225), .Z(n18224) );
  XOR U17967 ( .A(p_input[1721]), .B(p_input[1689]), .Z(n18225) );
  XOR U17968 ( .A(n18226), .B(n18227), .Z(n18217) );
  AND U17969 ( .A(n18228), .B(n18229), .Z(n18227) );
  XOR U17970 ( .A(n18226), .B(n17881), .Z(n18229) );
  XNOR U17971 ( .A(p_input[1752]), .B(n18230), .Z(n17881) );
  AND U17972 ( .A(n442), .B(n18231), .Z(n18230) );
  XOR U17973 ( .A(p_input[1784]), .B(p_input[1752]), .Z(n18231) );
  XNOR U17974 ( .A(n17878), .B(n18226), .Z(n18228) );
  XOR U17975 ( .A(n18232), .B(n18233), .Z(n17878) );
  AND U17976 ( .A(n440), .B(n18234), .Z(n18233) );
  XOR U17977 ( .A(p_input[1720]), .B(p_input[1688]), .Z(n18234) );
  XOR U17978 ( .A(n18235), .B(n18236), .Z(n18226) );
  AND U17979 ( .A(n18237), .B(n18238), .Z(n18236) );
  XOR U17980 ( .A(n18235), .B(n17893), .Z(n18238) );
  XNOR U17981 ( .A(p_input[1751]), .B(n18239), .Z(n17893) );
  AND U17982 ( .A(n442), .B(n18240), .Z(n18239) );
  XOR U17983 ( .A(p_input[1783]), .B(p_input[1751]), .Z(n18240) );
  XNOR U17984 ( .A(n17890), .B(n18235), .Z(n18237) );
  XOR U17985 ( .A(n18241), .B(n18242), .Z(n17890) );
  AND U17986 ( .A(n440), .B(n18243), .Z(n18242) );
  XOR U17987 ( .A(p_input[1719]), .B(p_input[1687]), .Z(n18243) );
  XOR U17988 ( .A(n18244), .B(n18245), .Z(n18235) );
  AND U17989 ( .A(n18246), .B(n18247), .Z(n18245) );
  XOR U17990 ( .A(n18244), .B(n17905), .Z(n18247) );
  XNOR U17991 ( .A(p_input[1750]), .B(n18248), .Z(n17905) );
  AND U17992 ( .A(n442), .B(n18249), .Z(n18248) );
  XOR U17993 ( .A(p_input[1782]), .B(p_input[1750]), .Z(n18249) );
  XNOR U17994 ( .A(n17902), .B(n18244), .Z(n18246) );
  XOR U17995 ( .A(n18250), .B(n18251), .Z(n17902) );
  AND U17996 ( .A(n440), .B(n18252), .Z(n18251) );
  XOR U17997 ( .A(p_input[1718]), .B(p_input[1686]), .Z(n18252) );
  XOR U17998 ( .A(n18253), .B(n18254), .Z(n18244) );
  AND U17999 ( .A(n18255), .B(n18256), .Z(n18254) );
  XOR U18000 ( .A(n18253), .B(n17917), .Z(n18256) );
  XNOR U18001 ( .A(p_input[1749]), .B(n18257), .Z(n17917) );
  AND U18002 ( .A(n442), .B(n18258), .Z(n18257) );
  XOR U18003 ( .A(p_input[1781]), .B(p_input[1749]), .Z(n18258) );
  XNOR U18004 ( .A(n17914), .B(n18253), .Z(n18255) );
  XOR U18005 ( .A(n18259), .B(n18260), .Z(n17914) );
  AND U18006 ( .A(n440), .B(n18261), .Z(n18260) );
  XOR U18007 ( .A(p_input[1717]), .B(p_input[1685]), .Z(n18261) );
  XOR U18008 ( .A(n18262), .B(n18263), .Z(n18253) );
  AND U18009 ( .A(n18264), .B(n18265), .Z(n18263) );
  XOR U18010 ( .A(n18262), .B(n17929), .Z(n18265) );
  XNOR U18011 ( .A(p_input[1748]), .B(n18266), .Z(n17929) );
  AND U18012 ( .A(n442), .B(n18267), .Z(n18266) );
  XOR U18013 ( .A(p_input[1780]), .B(p_input[1748]), .Z(n18267) );
  XNOR U18014 ( .A(n17926), .B(n18262), .Z(n18264) );
  XOR U18015 ( .A(n18268), .B(n18269), .Z(n17926) );
  AND U18016 ( .A(n440), .B(n18270), .Z(n18269) );
  XOR U18017 ( .A(p_input[1716]), .B(p_input[1684]), .Z(n18270) );
  XOR U18018 ( .A(n18271), .B(n18272), .Z(n18262) );
  AND U18019 ( .A(n18273), .B(n18274), .Z(n18272) );
  XOR U18020 ( .A(n18271), .B(n17941), .Z(n18274) );
  XNOR U18021 ( .A(p_input[1747]), .B(n18275), .Z(n17941) );
  AND U18022 ( .A(n442), .B(n18276), .Z(n18275) );
  XOR U18023 ( .A(p_input[1779]), .B(p_input[1747]), .Z(n18276) );
  XNOR U18024 ( .A(n17938), .B(n18271), .Z(n18273) );
  XOR U18025 ( .A(n18277), .B(n18278), .Z(n17938) );
  AND U18026 ( .A(n440), .B(n18279), .Z(n18278) );
  XOR U18027 ( .A(p_input[1715]), .B(p_input[1683]), .Z(n18279) );
  XOR U18028 ( .A(n18280), .B(n18281), .Z(n18271) );
  AND U18029 ( .A(n18282), .B(n18283), .Z(n18281) );
  XOR U18030 ( .A(n18280), .B(n17953), .Z(n18283) );
  XNOR U18031 ( .A(p_input[1746]), .B(n18284), .Z(n17953) );
  AND U18032 ( .A(n442), .B(n18285), .Z(n18284) );
  XOR U18033 ( .A(p_input[1778]), .B(p_input[1746]), .Z(n18285) );
  XNOR U18034 ( .A(n17950), .B(n18280), .Z(n18282) );
  XOR U18035 ( .A(n18286), .B(n18287), .Z(n17950) );
  AND U18036 ( .A(n440), .B(n18288), .Z(n18287) );
  XOR U18037 ( .A(p_input[1714]), .B(p_input[1682]), .Z(n18288) );
  XOR U18038 ( .A(n18289), .B(n18290), .Z(n18280) );
  AND U18039 ( .A(n18291), .B(n18292), .Z(n18290) );
  XOR U18040 ( .A(n18289), .B(n17965), .Z(n18292) );
  XNOR U18041 ( .A(p_input[1745]), .B(n18293), .Z(n17965) );
  AND U18042 ( .A(n442), .B(n18294), .Z(n18293) );
  XOR U18043 ( .A(p_input[1777]), .B(p_input[1745]), .Z(n18294) );
  XNOR U18044 ( .A(n17962), .B(n18289), .Z(n18291) );
  XOR U18045 ( .A(n18295), .B(n18296), .Z(n17962) );
  AND U18046 ( .A(n440), .B(n18297), .Z(n18296) );
  XOR U18047 ( .A(p_input[1713]), .B(p_input[1681]), .Z(n18297) );
  XOR U18048 ( .A(n18298), .B(n18299), .Z(n18289) );
  AND U18049 ( .A(n18300), .B(n18301), .Z(n18299) );
  XOR U18050 ( .A(n18298), .B(n17977), .Z(n18301) );
  XNOR U18051 ( .A(p_input[1744]), .B(n18302), .Z(n17977) );
  AND U18052 ( .A(n442), .B(n18303), .Z(n18302) );
  XOR U18053 ( .A(p_input[1776]), .B(p_input[1744]), .Z(n18303) );
  XNOR U18054 ( .A(n17974), .B(n18298), .Z(n18300) );
  XOR U18055 ( .A(n18304), .B(n18305), .Z(n17974) );
  AND U18056 ( .A(n440), .B(n18306), .Z(n18305) );
  XOR U18057 ( .A(p_input[1712]), .B(p_input[1680]), .Z(n18306) );
  XOR U18058 ( .A(n18307), .B(n18308), .Z(n18298) );
  AND U18059 ( .A(n18309), .B(n18310), .Z(n18308) );
  XOR U18060 ( .A(n18307), .B(n17989), .Z(n18310) );
  XNOR U18061 ( .A(p_input[1743]), .B(n18311), .Z(n17989) );
  AND U18062 ( .A(n442), .B(n18312), .Z(n18311) );
  XOR U18063 ( .A(p_input[1775]), .B(p_input[1743]), .Z(n18312) );
  XNOR U18064 ( .A(n17986), .B(n18307), .Z(n18309) );
  XOR U18065 ( .A(n18313), .B(n18314), .Z(n17986) );
  AND U18066 ( .A(n440), .B(n18315), .Z(n18314) );
  XOR U18067 ( .A(p_input[1711]), .B(p_input[1679]), .Z(n18315) );
  XOR U18068 ( .A(n18316), .B(n18317), .Z(n18307) );
  AND U18069 ( .A(n18318), .B(n18319), .Z(n18317) );
  XOR U18070 ( .A(n18316), .B(n18001), .Z(n18319) );
  XNOR U18071 ( .A(p_input[1742]), .B(n18320), .Z(n18001) );
  AND U18072 ( .A(n442), .B(n18321), .Z(n18320) );
  XOR U18073 ( .A(p_input[1774]), .B(p_input[1742]), .Z(n18321) );
  XNOR U18074 ( .A(n17998), .B(n18316), .Z(n18318) );
  XOR U18075 ( .A(n18322), .B(n18323), .Z(n17998) );
  AND U18076 ( .A(n440), .B(n18324), .Z(n18323) );
  XOR U18077 ( .A(p_input[1710]), .B(p_input[1678]), .Z(n18324) );
  XOR U18078 ( .A(n18325), .B(n18326), .Z(n18316) );
  AND U18079 ( .A(n18327), .B(n18328), .Z(n18326) );
  XOR U18080 ( .A(n18325), .B(n18013), .Z(n18328) );
  XNOR U18081 ( .A(p_input[1741]), .B(n18329), .Z(n18013) );
  AND U18082 ( .A(n442), .B(n18330), .Z(n18329) );
  XOR U18083 ( .A(p_input[1773]), .B(p_input[1741]), .Z(n18330) );
  XNOR U18084 ( .A(n18010), .B(n18325), .Z(n18327) );
  XOR U18085 ( .A(n18331), .B(n18332), .Z(n18010) );
  AND U18086 ( .A(n440), .B(n18333), .Z(n18332) );
  XOR U18087 ( .A(p_input[1709]), .B(p_input[1677]), .Z(n18333) );
  XOR U18088 ( .A(n18334), .B(n18335), .Z(n18325) );
  AND U18089 ( .A(n18336), .B(n18337), .Z(n18335) );
  XOR U18090 ( .A(n18334), .B(n18025), .Z(n18337) );
  XNOR U18091 ( .A(p_input[1740]), .B(n18338), .Z(n18025) );
  AND U18092 ( .A(n442), .B(n18339), .Z(n18338) );
  XOR U18093 ( .A(p_input[1772]), .B(p_input[1740]), .Z(n18339) );
  XNOR U18094 ( .A(n18022), .B(n18334), .Z(n18336) );
  XOR U18095 ( .A(n18340), .B(n18341), .Z(n18022) );
  AND U18096 ( .A(n440), .B(n18342), .Z(n18341) );
  XOR U18097 ( .A(p_input[1708]), .B(p_input[1676]), .Z(n18342) );
  XOR U18098 ( .A(n18343), .B(n18344), .Z(n18334) );
  AND U18099 ( .A(n18345), .B(n18346), .Z(n18344) );
  XOR U18100 ( .A(n18343), .B(n18037), .Z(n18346) );
  XNOR U18101 ( .A(p_input[1739]), .B(n18347), .Z(n18037) );
  AND U18102 ( .A(n442), .B(n18348), .Z(n18347) );
  XOR U18103 ( .A(p_input[1771]), .B(p_input[1739]), .Z(n18348) );
  XNOR U18104 ( .A(n18034), .B(n18343), .Z(n18345) );
  XOR U18105 ( .A(n18349), .B(n18350), .Z(n18034) );
  AND U18106 ( .A(n440), .B(n18351), .Z(n18350) );
  XOR U18107 ( .A(p_input[1707]), .B(p_input[1675]), .Z(n18351) );
  XOR U18108 ( .A(n18352), .B(n18353), .Z(n18343) );
  AND U18109 ( .A(n18354), .B(n18355), .Z(n18353) );
  XOR U18110 ( .A(n18352), .B(n18049), .Z(n18355) );
  XNOR U18111 ( .A(p_input[1738]), .B(n18356), .Z(n18049) );
  AND U18112 ( .A(n442), .B(n18357), .Z(n18356) );
  XOR U18113 ( .A(p_input[1770]), .B(p_input[1738]), .Z(n18357) );
  XNOR U18114 ( .A(n18046), .B(n18352), .Z(n18354) );
  XOR U18115 ( .A(n18358), .B(n18359), .Z(n18046) );
  AND U18116 ( .A(n440), .B(n18360), .Z(n18359) );
  XOR U18117 ( .A(p_input[1706]), .B(p_input[1674]), .Z(n18360) );
  XOR U18118 ( .A(n18361), .B(n18362), .Z(n18352) );
  AND U18119 ( .A(n18363), .B(n18364), .Z(n18362) );
  XOR U18120 ( .A(n18361), .B(n18061), .Z(n18364) );
  XNOR U18121 ( .A(p_input[1737]), .B(n18365), .Z(n18061) );
  AND U18122 ( .A(n442), .B(n18366), .Z(n18365) );
  XOR U18123 ( .A(p_input[1769]), .B(p_input[1737]), .Z(n18366) );
  XNOR U18124 ( .A(n18058), .B(n18361), .Z(n18363) );
  XOR U18125 ( .A(n18367), .B(n18368), .Z(n18058) );
  AND U18126 ( .A(n440), .B(n18369), .Z(n18368) );
  XOR U18127 ( .A(p_input[1705]), .B(p_input[1673]), .Z(n18369) );
  XOR U18128 ( .A(n18370), .B(n18371), .Z(n18361) );
  AND U18129 ( .A(n18372), .B(n18373), .Z(n18371) );
  XOR U18130 ( .A(n18370), .B(n18073), .Z(n18373) );
  XNOR U18131 ( .A(p_input[1736]), .B(n18374), .Z(n18073) );
  AND U18132 ( .A(n442), .B(n18375), .Z(n18374) );
  XOR U18133 ( .A(p_input[1768]), .B(p_input[1736]), .Z(n18375) );
  XNOR U18134 ( .A(n18070), .B(n18370), .Z(n18372) );
  XOR U18135 ( .A(n18376), .B(n18377), .Z(n18070) );
  AND U18136 ( .A(n440), .B(n18378), .Z(n18377) );
  XOR U18137 ( .A(p_input[1704]), .B(p_input[1672]), .Z(n18378) );
  XOR U18138 ( .A(n18379), .B(n18380), .Z(n18370) );
  AND U18139 ( .A(n18381), .B(n18382), .Z(n18380) );
  XOR U18140 ( .A(n18379), .B(n18085), .Z(n18382) );
  XNOR U18141 ( .A(p_input[1735]), .B(n18383), .Z(n18085) );
  AND U18142 ( .A(n442), .B(n18384), .Z(n18383) );
  XOR U18143 ( .A(p_input[1767]), .B(p_input[1735]), .Z(n18384) );
  XNOR U18144 ( .A(n18082), .B(n18379), .Z(n18381) );
  XOR U18145 ( .A(n18385), .B(n18386), .Z(n18082) );
  AND U18146 ( .A(n440), .B(n18387), .Z(n18386) );
  XOR U18147 ( .A(p_input[1703]), .B(p_input[1671]), .Z(n18387) );
  XOR U18148 ( .A(n18388), .B(n18389), .Z(n18379) );
  AND U18149 ( .A(n18390), .B(n18391), .Z(n18389) );
  XOR U18150 ( .A(n18388), .B(n18097), .Z(n18391) );
  XNOR U18151 ( .A(p_input[1734]), .B(n18392), .Z(n18097) );
  AND U18152 ( .A(n442), .B(n18393), .Z(n18392) );
  XOR U18153 ( .A(p_input[1766]), .B(p_input[1734]), .Z(n18393) );
  XNOR U18154 ( .A(n18094), .B(n18388), .Z(n18390) );
  XOR U18155 ( .A(n18394), .B(n18395), .Z(n18094) );
  AND U18156 ( .A(n440), .B(n18396), .Z(n18395) );
  XOR U18157 ( .A(p_input[1702]), .B(p_input[1670]), .Z(n18396) );
  XOR U18158 ( .A(n18397), .B(n18398), .Z(n18388) );
  AND U18159 ( .A(n18399), .B(n18400), .Z(n18398) );
  XOR U18160 ( .A(n18397), .B(n18109), .Z(n18400) );
  XNOR U18161 ( .A(p_input[1733]), .B(n18401), .Z(n18109) );
  AND U18162 ( .A(n442), .B(n18402), .Z(n18401) );
  XOR U18163 ( .A(p_input[1765]), .B(p_input[1733]), .Z(n18402) );
  XNOR U18164 ( .A(n18106), .B(n18397), .Z(n18399) );
  XOR U18165 ( .A(n18403), .B(n18404), .Z(n18106) );
  AND U18166 ( .A(n440), .B(n18405), .Z(n18404) );
  XOR U18167 ( .A(p_input[1701]), .B(p_input[1669]), .Z(n18405) );
  XOR U18168 ( .A(n18406), .B(n18407), .Z(n18397) );
  AND U18169 ( .A(n18408), .B(n18409), .Z(n18407) );
  XOR U18170 ( .A(n18406), .B(n18121), .Z(n18409) );
  XNOR U18171 ( .A(p_input[1732]), .B(n18410), .Z(n18121) );
  AND U18172 ( .A(n442), .B(n18411), .Z(n18410) );
  XOR U18173 ( .A(p_input[1764]), .B(p_input[1732]), .Z(n18411) );
  XNOR U18174 ( .A(n18118), .B(n18406), .Z(n18408) );
  XOR U18175 ( .A(n18412), .B(n18413), .Z(n18118) );
  AND U18176 ( .A(n440), .B(n18414), .Z(n18413) );
  XOR U18177 ( .A(p_input[1700]), .B(p_input[1668]), .Z(n18414) );
  XOR U18178 ( .A(n18415), .B(n18416), .Z(n18406) );
  AND U18179 ( .A(n18417), .B(n18418), .Z(n18416) );
  XOR U18180 ( .A(n18415), .B(n18133), .Z(n18418) );
  XNOR U18181 ( .A(p_input[1731]), .B(n18419), .Z(n18133) );
  AND U18182 ( .A(n442), .B(n18420), .Z(n18419) );
  XOR U18183 ( .A(p_input[1763]), .B(p_input[1731]), .Z(n18420) );
  XNOR U18184 ( .A(n18130), .B(n18415), .Z(n18417) );
  XOR U18185 ( .A(n18421), .B(n18422), .Z(n18130) );
  AND U18186 ( .A(n440), .B(n18423), .Z(n18422) );
  XOR U18187 ( .A(p_input[1699]), .B(p_input[1667]), .Z(n18423) );
  XOR U18188 ( .A(n18424), .B(n18425), .Z(n18415) );
  AND U18189 ( .A(n18426), .B(n18427), .Z(n18425) );
  XOR U18190 ( .A(n18145), .B(n18424), .Z(n18427) );
  XNOR U18191 ( .A(p_input[1730]), .B(n18428), .Z(n18145) );
  AND U18192 ( .A(n442), .B(n18429), .Z(n18428) );
  XOR U18193 ( .A(p_input[1762]), .B(p_input[1730]), .Z(n18429) );
  XNOR U18194 ( .A(n18424), .B(n18142), .Z(n18426) );
  XOR U18195 ( .A(n18430), .B(n18431), .Z(n18142) );
  AND U18196 ( .A(n440), .B(n18432), .Z(n18431) );
  XOR U18197 ( .A(p_input[1698]), .B(p_input[1666]), .Z(n18432) );
  XOR U18198 ( .A(n18433), .B(n18434), .Z(n18424) );
  AND U18199 ( .A(n18435), .B(n18436), .Z(n18434) );
  XNOR U18200 ( .A(n18437), .B(n18158), .Z(n18436) );
  XNOR U18201 ( .A(p_input[1729]), .B(n18438), .Z(n18158) );
  AND U18202 ( .A(n442), .B(n18439), .Z(n18438) );
  XNOR U18203 ( .A(p_input[1761]), .B(n18440), .Z(n18439) );
  IV U18204 ( .A(p_input[1729]), .Z(n18440) );
  XNOR U18205 ( .A(n18155), .B(n18433), .Z(n18435) );
  XNOR U18206 ( .A(p_input[1665]), .B(n18441), .Z(n18155) );
  AND U18207 ( .A(n440), .B(n18442), .Z(n18441) );
  XOR U18208 ( .A(p_input[1697]), .B(p_input[1665]), .Z(n18442) );
  IV U18209 ( .A(n18437), .Z(n18433) );
  AND U18210 ( .A(n18163), .B(n18166), .Z(n18437) );
  XOR U18211 ( .A(p_input[1728]), .B(n18443), .Z(n18166) );
  AND U18212 ( .A(n442), .B(n18444), .Z(n18443) );
  XOR U18213 ( .A(p_input[1760]), .B(p_input[1728]), .Z(n18444) );
  XOR U18214 ( .A(n18445), .B(n18446), .Z(n442) );
  AND U18215 ( .A(n18447), .B(n18448), .Z(n18446) );
  XNOR U18216 ( .A(p_input[1791]), .B(n18445), .Z(n18448) );
  XOR U18217 ( .A(n18445), .B(p_input[1759]), .Z(n18447) );
  XOR U18218 ( .A(n18449), .B(n18450), .Z(n18445) );
  AND U18219 ( .A(n18451), .B(n18452), .Z(n18450) );
  XNOR U18220 ( .A(p_input[1790]), .B(n18449), .Z(n18452) );
  XOR U18221 ( .A(n18449), .B(p_input[1758]), .Z(n18451) );
  XOR U18222 ( .A(n18453), .B(n18454), .Z(n18449) );
  AND U18223 ( .A(n18455), .B(n18456), .Z(n18454) );
  XNOR U18224 ( .A(p_input[1789]), .B(n18453), .Z(n18456) );
  XOR U18225 ( .A(n18453), .B(p_input[1757]), .Z(n18455) );
  XOR U18226 ( .A(n18457), .B(n18458), .Z(n18453) );
  AND U18227 ( .A(n18459), .B(n18460), .Z(n18458) );
  XNOR U18228 ( .A(p_input[1788]), .B(n18457), .Z(n18460) );
  XOR U18229 ( .A(n18457), .B(p_input[1756]), .Z(n18459) );
  XOR U18230 ( .A(n18461), .B(n18462), .Z(n18457) );
  AND U18231 ( .A(n18463), .B(n18464), .Z(n18462) );
  XNOR U18232 ( .A(p_input[1787]), .B(n18461), .Z(n18464) );
  XOR U18233 ( .A(n18461), .B(p_input[1755]), .Z(n18463) );
  XOR U18234 ( .A(n18465), .B(n18466), .Z(n18461) );
  AND U18235 ( .A(n18467), .B(n18468), .Z(n18466) );
  XNOR U18236 ( .A(p_input[1786]), .B(n18465), .Z(n18468) );
  XOR U18237 ( .A(n18465), .B(p_input[1754]), .Z(n18467) );
  XOR U18238 ( .A(n18469), .B(n18470), .Z(n18465) );
  AND U18239 ( .A(n18471), .B(n18472), .Z(n18470) );
  XNOR U18240 ( .A(p_input[1785]), .B(n18469), .Z(n18472) );
  XOR U18241 ( .A(n18469), .B(p_input[1753]), .Z(n18471) );
  XOR U18242 ( .A(n18473), .B(n18474), .Z(n18469) );
  AND U18243 ( .A(n18475), .B(n18476), .Z(n18474) );
  XNOR U18244 ( .A(p_input[1784]), .B(n18473), .Z(n18476) );
  XOR U18245 ( .A(n18473), .B(p_input[1752]), .Z(n18475) );
  XOR U18246 ( .A(n18477), .B(n18478), .Z(n18473) );
  AND U18247 ( .A(n18479), .B(n18480), .Z(n18478) );
  XNOR U18248 ( .A(p_input[1783]), .B(n18477), .Z(n18480) );
  XOR U18249 ( .A(n18477), .B(p_input[1751]), .Z(n18479) );
  XOR U18250 ( .A(n18481), .B(n18482), .Z(n18477) );
  AND U18251 ( .A(n18483), .B(n18484), .Z(n18482) );
  XNOR U18252 ( .A(p_input[1782]), .B(n18481), .Z(n18484) );
  XOR U18253 ( .A(n18481), .B(p_input[1750]), .Z(n18483) );
  XOR U18254 ( .A(n18485), .B(n18486), .Z(n18481) );
  AND U18255 ( .A(n18487), .B(n18488), .Z(n18486) );
  XNOR U18256 ( .A(p_input[1781]), .B(n18485), .Z(n18488) );
  XOR U18257 ( .A(n18485), .B(p_input[1749]), .Z(n18487) );
  XOR U18258 ( .A(n18489), .B(n18490), .Z(n18485) );
  AND U18259 ( .A(n18491), .B(n18492), .Z(n18490) );
  XNOR U18260 ( .A(p_input[1780]), .B(n18489), .Z(n18492) );
  XOR U18261 ( .A(n18489), .B(p_input[1748]), .Z(n18491) );
  XOR U18262 ( .A(n18493), .B(n18494), .Z(n18489) );
  AND U18263 ( .A(n18495), .B(n18496), .Z(n18494) );
  XNOR U18264 ( .A(p_input[1779]), .B(n18493), .Z(n18496) );
  XOR U18265 ( .A(n18493), .B(p_input[1747]), .Z(n18495) );
  XOR U18266 ( .A(n18497), .B(n18498), .Z(n18493) );
  AND U18267 ( .A(n18499), .B(n18500), .Z(n18498) );
  XNOR U18268 ( .A(p_input[1778]), .B(n18497), .Z(n18500) );
  XOR U18269 ( .A(n18497), .B(p_input[1746]), .Z(n18499) );
  XOR U18270 ( .A(n18501), .B(n18502), .Z(n18497) );
  AND U18271 ( .A(n18503), .B(n18504), .Z(n18502) );
  XNOR U18272 ( .A(p_input[1777]), .B(n18501), .Z(n18504) );
  XOR U18273 ( .A(n18501), .B(p_input[1745]), .Z(n18503) );
  XOR U18274 ( .A(n18505), .B(n18506), .Z(n18501) );
  AND U18275 ( .A(n18507), .B(n18508), .Z(n18506) );
  XNOR U18276 ( .A(p_input[1776]), .B(n18505), .Z(n18508) );
  XOR U18277 ( .A(n18505), .B(p_input[1744]), .Z(n18507) );
  XOR U18278 ( .A(n18509), .B(n18510), .Z(n18505) );
  AND U18279 ( .A(n18511), .B(n18512), .Z(n18510) );
  XNOR U18280 ( .A(p_input[1775]), .B(n18509), .Z(n18512) );
  XOR U18281 ( .A(n18509), .B(p_input[1743]), .Z(n18511) );
  XOR U18282 ( .A(n18513), .B(n18514), .Z(n18509) );
  AND U18283 ( .A(n18515), .B(n18516), .Z(n18514) );
  XNOR U18284 ( .A(p_input[1774]), .B(n18513), .Z(n18516) );
  XOR U18285 ( .A(n18513), .B(p_input[1742]), .Z(n18515) );
  XOR U18286 ( .A(n18517), .B(n18518), .Z(n18513) );
  AND U18287 ( .A(n18519), .B(n18520), .Z(n18518) );
  XNOR U18288 ( .A(p_input[1773]), .B(n18517), .Z(n18520) );
  XOR U18289 ( .A(n18517), .B(p_input[1741]), .Z(n18519) );
  XOR U18290 ( .A(n18521), .B(n18522), .Z(n18517) );
  AND U18291 ( .A(n18523), .B(n18524), .Z(n18522) );
  XNOR U18292 ( .A(p_input[1772]), .B(n18521), .Z(n18524) );
  XOR U18293 ( .A(n18521), .B(p_input[1740]), .Z(n18523) );
  XOR U18294 ( .A(n18525), .B(n18526), .Z(n18521) );
  AND U18295 ( .A(n18527), .B(n18528), .Z(n18526) );
  XNOR U18296 ( .A(p_input[1771]), .B(n18525), .Z(n18528) );
  XOR U18297 ( .A(n18525), .B(p_input[1739]), .Z(n18527) );
  XOR U18298 ( .A(n18529), .B(n18530), .Z(n18525) );
  AND U18299 ( .A(n18531), .B(n18532), .Z(n18530) );
  XNOR U18300 ( .A(p_input[1770]), .B(n18529), .Z(n18532) );
  XOR U18301 ( .A(n18529), .B(p_input[1738]), .Z(n18531) );
  XOR U18302 ( .A(n18533), .B(n18534), .Z(n18529) );
  AND U18303 ( .A(n18535), .B(n18536), .Z(n18534) );
  XNOR U18304 ( .A(p_input[1769]), .B(n18533), .Z(n18536) );
  XOR U18305 ( .A(n18533), .B(p_input[1737]), .Z(n18535) );
  XOR U18306 ( .A(n18537), .B(n18538), .Z(n18533) );
  AND U18307 ( .A(n18539), .B(n18540), .Z(n18538) );
  XNOR U18308 ( .A(p_input[1768]), .B(n18537), .Z(n18540) );
  XOR U18309 ( .A(n18537), .B(p_input[1736]), .Z(n18539) );
  XOR U18310 ( .A(n18541), .B(n18542), .Z(n18537) );
  AND U18311 ( .A(n18543), .B(n18544), .Z(n18542) );
  XNOR U18312 ( .A(p_input[1767]), .B(n18541), .Z(n18544) );
  XOR U18313 ( .A(n18541), .B(p_input[1735]), .Z(n18543) );
  XOR U18314 ( .A(n18545), .B(n18546), .Z(n18541) );
  AND U18315 ( .A(n18547), .B(n18548), .Z(n18546) );
  XNOR U18316 ( .A(p_input[1766]), .B(n18545), .Z(n18548) );
  XOR U18317 ( .A(n18545), .B(p_input[1734]), .Z(n18547) );
  XOR U18318 ( .A(n18549), .B(n18550), .Z(n18545) );
  AND U18319 ( .A(n18551), .B(n18552), .Z(n18550) );
  XNOR U18320 ( .A(p_input[1765]), .B(n18549), .Z(n18552) );
  XOR U18321 ( .A(n18549), .B(p_input[1733]), .Z(n18551) );
  XOR U18322 ( .A(n18553), .B(n18554), .Z(n18549) );
  AND U18323 ( .A(n18555), .B(n18556), .Z(n18554) );
  XNOR U18324 ( .A(p_input[1764]), .B(n18553), .Z(n18556) );
  XOR U18325 ( .A(n18553), .B(p_input[1732]), .Z(n18555) );
  XOR U18326 ( .A(n18557), .B(n18558), .Z(n18553) );
  AND U18327 ( .A(n18559), .B(n18560), .Z(n18558) );
  XNOR U18328 ( .A(p_input[1763]), .B(n18557), .Z(n18560) );
  XOR U18329 ( .A(n18557), .B(p_input[1731]), .Z(n18559) );
  XOR U18330 ( .A(n18561), .B(n18562), .Z(n18557) );
  AND U18331 ( .A(n18563), .B(n18564), .Z(n18562) );
  XNOR U18332 ( .A(p_input[1762]), .B(n18561), .Z(n18564) );
  XOR U18333 ( .A(n18561), .B(p_input[1730]), .Z(n18563) );
  XNOR U18334 ( .A(n18565), .B(n18566), .Z(n18561) );
  AND U18335 ( .A(n18567), .B(n18568), .Z(n18566) );
  XOR U18336 ( .A(p_input[1761]), .B(n18565), .Z(n18568) );
  XNOR U18337 ( .A(p_input[1729]), .B(n18565), .Z(n18567) );
  AND U18338 ( .A(p_input[1760]), .B(n18569), .Z(n18565) );
  IV U18339 ( .A(p_input[1728]), .Z(n18569) );
  XNOR U18340 ( .A(p_input[1664]), .B(n18570), .Z(n18163) );
  AND U18341 ( .A(n440), .B(n18571), .Z(n18570) );
  XOR U18342 ( .A(p_input[1696]), .B(p_input[1664]), .Z(n18571) );
  XOR U18343 ( .A(n18572), .B(n18573), .Z(n440) );
  AND U18344 ( .A(n18574), .B(n18575), .Z(n18573) );
  XNOR U18345 ( .A(p_input[1727]), .B(n18572), .Z(n18575) );
  XOR U18346 ( .A(n18572), .B(p_input[1695]), .Z(n18574) );
  XOR U18347 ( .A(n18576), .B(n18577), .Z(n18572) );
  AND U18348 ( .A(n18578), .B(n18579), .Z(n18577) );
  XNOR U18349 ( .A(p_input[1726]), .B(n18576), .Z(n18579) );
  XNOR U18350 ( .A(n18576), .B(n18178), .Z(n18578) );
  IV U18351 ( .A(p_input[1694]), .Z(n18178) );
  XOR U18352 ( .A(n18580), .B(n18581), .Z(n18576) );
  AND U18353 ( .A(n18582), .B(n18583), .Z(n18581) );
  XNOR U18354 ( .A(p_input[1725]), .B(n18580), .Z(n18583) );
  XNOR U18355 ( .A(n18580), .B(n18187), .Z(n18582) );
  IV U18356 ( .A(p_input[1693]), .Z(n18187) );
  XOR U18357 ( .A(n18584), .B(n18585), .Z(n18580) );
  AND U18358 ( .A(n18586), .B(n18587), .Z(n18585) );
  XNOR U18359 ( .A(p_input[1724]), .B(n18584), .Z(n18587) );
  XNOR U18360 ( .A(n18584), .B(n18196), .Z(n18586) );
  IV U18361 ( .A(p_input[1692]), .Z(n18196) );
  XOR U18362 ( .A(n18588), .B(n18589), .Z(n18584) );
  AND U18363 ( .A(n18590), .B(n18591), .Z(n18589) );
  XNOR U18364 ( .A(p_input[1723]), .B(n18588), .Z(n18591) );
  XNOR U18365 ( .A(n18588), .B(n18205), .Z(n18590) );
  IV U18366 ( .A(p_input[1691]), .Z(n18205) );
  XOR U18367 ( .A(n18592), .B(n18593), .Z(n18588) );
  AND U18368 ( .A(n18594), .B(n18595), .Z(n18593) );
  XNOR U18369 ( .A(p_input[1722]), .B(n18592), .Z(n18595) );
  XNOR U18370 ( .A(n18592), .B(n18214), .Z(n18594) );
  IV U18371 ( .A(p_input[1690]), .Z(n18214) );
  XOR U18372 ( .A(n18596), .B(n18597), .Z(n18592) );
  AND U18373 ( .A(n18598), .B(n18599), .Z(n18597) );
  XNOR U18374 ( .A(p_input[1721]), .B(n18596), .Z(n18599) );
  XNOR U18375 ( .A(n18596), .B(n18223), .Z(n18598) );
  IV U18376 ( .A(p_input[1689]), .Z(n18223) );
  XOR U18377 ( .A(n18600), .B(n18601), .Z(n18596) );
  AND U18378 ( .A(n18602), .B(n18603), .Z(n18601) );
  XNOR U18379 ( .A(p_input[1720]), .B(n18600), .Z(n18603) );
  XNOR U18380 ( .A(n18600), .B(n18232), .Z(n18602) );
  IV U18381 ( .A(p_input[1688]), .Z(n18232) );
  XOR U18382 ( .A(n18604), .B(n18605), .Z(n18600) );
  AND U18383 ( .A(n18606), .B(n18607), .Z(n18605) );
  XNOR U18384 ( .A(p_input[1719]), .B(n18604), .Z(n18607) );
  XNOR U18385 ( .A(n18604), .B(n18241), .Z(n18606) );
  IV U18386 ( .A(p_input[1687]), .Z(n18241) );
  XOR U18387 ( .A(n18608), .B(n18609), .Z(n18604) );
  AND U18388 ( .A(n18610), .B(n18611), .Z(n18609) );
  XNOR U18389 ( .A(p_input[1718]), .B(n18608), .Z(n18611) );
  XNOR U18390 ( .A(n18608), .B(n18250), .Z(n18610) );
  IV U18391 ( .A(p_input[1686]), .Z(n18250) );
  XOR U18392 ( .A(n18612), .B(n18613), .Z(n18608) );
  AND U18393 ( .A(n18614), .B(n18615), .Z(n18613) );
  XNOR U18394 ( .A(p_input[1717]), .B(n18612), .Z(n18615) );
  XNOR U18395 ( .A(n18612), .B(n18259), .Z(n18614) );
  IV U18396 ( .A(p_input[1685]), .Z(n18259) );
  XOR U18397 ( .A(n18616), .B(n18617), .Z(n18612) );
  AND U18398 ( .A(n18618), .B(n18619), .Z(n18617) );
  XNOR U18399 ( .A(p_input[1716]), .B(n18616), .Z(n18619) );
  XNOR U18400 ( .A(n18616), .B(n18268), .Z(n18618) );
  IV U18401 ( .A(p_input[1684]), .Z(n18268) );
  XOR U18402 ( .A(n18620), .B(n18621), .Z(n18616) );
  AND U18403 ( .A(n18622), .B(n18623), .Z(n18621) );
  XNOR U18404 ( .A(p_input[1715]), .B(n18620), .Z(n18623) );
  XNOR U18405 ( .A(n18620), .B(n18277), .Z(n18622) );
  IV U18406 ( .A(p_input[1683]), .Z(n18277) );
  XOR U18407 ( .A(n18624), .B(n18625), .Z(n18620) );
  AND U18408 ( .A(n18626), .B(n18627), .Z(n18625) );
  XNOR U18409 ( .A(p_input[1714]), .B(n18624), .Z(n18627) );
  XNOR U18410 ( .A(n18624), .B(n18286), .Z(n18626) );
  IV U18411 ( .A(p_input[1682]), .Z(n18286) );
  XOR U18412 ( .A(n18628), .B(n18629), .Z(n18624) );
  AND U18413 ( .A(n18630), .B(n18631), .Z(n18629) );
  XNOR U18414 ( .A(p_input[1713]), .B(n18628), .Z(n18631) );
  XNOR U18415 ( .A(n18628), .B(n18295), .Z(n18630) );
  IV U18416 ( .A(p_input[1681]), .Z(n18295) );
  XOR U18417 ( .A(n18632), .B(n18633), .Z(n18628) );
  AND U18418 ( .A(n18634), .B(n18635), .Z(n18633) );
  XNOR U18419 ( .A(p_input[1712]), .B(n18632), .Z(n18635) );
  XNOR U18420 ( .A(n18632), .B(n18304), .Z(n18634) );
  IV U18421 ( .A(p_input[1680]), .Z(n18304) );
  XOR U18422 ( .A(n18636), .B(n18637), .Z(n18632) );
  AND U18423 ( .A(n18638), .B(n18639), .Z(n18637) );
  XNOR U18424 ( .A(p_input[1711]), .B(n18636), .Z(n18639) );
  XNOR U18425 ( .A(n18636), .B(n18313), .Z(n18638) );
  IV U18426 ( .A(p_input[1679]), .Z(n18313) );
  XOR U18427 ( .A(n18640), .B(n18641), .Z(n18636) );
  AND U18428 ( .A(n18642), .B(n18643), .Z(n18641) );
  XNOR U18429 ( .A(p_input[1710]), .B(n18640), .Z(n18643) );
  XNOR U18430 ( .A(n18640), .B(n18322), .Z(n18642) );
  IV U18431 ( .A(p_input[1678]), .Z(n18322) );
  XOR U18432 ( .A(n18644), .B(n18645), .Z(n18640) );
  AND U18433 ( .A(n18646), .B(n18647), .Z(n18645) );
  XNOR U18434 ( .A(p_input[1709]), .B(n18644), .Z(n18647) );
  XNOR U18435 ( .A(n18644), .B(n18331), .Z(n18646) );
  IV U18436 ( .A(p_input[1677]), .Z(n18331) );
  XOR U18437 ( .A(n18648), .B(n18649), .Z(n18644) );
  AND U18438 ( .A(n18650), .B(n18651), .Z(n18649) );
  XNOR U18439 ( .A(p_input[1708]), .B(n18648), .Z(n18651) );
  XNOR U18440 ( .A(n18648), .B(n18340), .Z(n18650) );
  IV U18441 ( .A(p_input[1676]), .Z(n18340) );
  XOR U18442 ( .A(n18652), .B(n18653), .Z(n18648) );
  AND U18443 ( .A(n18654), .B(n18655), .Z(n18653) );
  XNOR U18444 ( .A(p_input[1707]), .B(n18652), .Z(n18655) );
  XNOR U18445 ( .A(n18652), .B(n18349), .Z(n18654) );
  IV U18446 ( .A(p_input[1675]), .Z(n18349) );
  XOR U18447 ( .A(n18656), .B(n18657), .Z(n18652) );
  AND U18448 ( .A(n18658), .B(n18659), .Z(n18657) );
  XNOR U18449 ( .A(p_input[1706]), .B(n18656), .Z(n18659) );
  XNOR U18450 ( .A(n18656), .B(n18358), .Z(n18658) );
  IV U18451 ( .A(p_input[1674]), .Z(n18358) );
  XOR U18452 ( .A(n18660), .B(n18661), .Z(n18656) );
  AND U18453 ( .A(n18662), .B(n18663), .Z(n18661) );
  XNOR U18454 ( .A(p_input[1705]), .B(n18660), .Z(n18663) );
  XNOR U18455 ( .A(n18660), .B(n18367), .Z(n18662) );
  IV U18456 ( .A(p_input[1673]), .Z(n18367) );
  XOR U18457 ( .A(n18664), .B(n18665), .Z(n18660) );
  AND U18458 ( .A(n18666), .B(n18667), .Z(n18665) );
  XNOR U18459 ( .A(p_input[1704]), .B(n18664), .Z(n18667) );
  XNOR U18460 ( .A(n18664), .B(n18376), .Z(n18666) );
  IV U18461 ( .A(p_input[1672]), .Z(n18376) );
  XOR U18462 ( .A(n18668), .B(n18669), .Z(n18664) );
  AND U18463 ( .A(n18670), .B(n18671), .Z(n18669) );
  XNOR U18464 ( .A(p_input[1703]), .B(n18668), .Z(n18671) );
  XNOR U18465 ( .A(n18668), .B(n18385), .Z(n18670) );
  IV U18466 ( .A(p_input[1671]), .Z(n18385) );
  XOR U18467 ( .A(n18672), .B(n18673), .Z(n18668) );
  AND U18468 ( .A(n18674), .B(n18675), .Z(n18673) );
  XNOR U18469 ( .A(p_input[1702]), .B(n18672), .Z(n18675) );
  XNOR U18470 ( .A(n18672), .B(n18394), .Z(n18674) );
  IV U18471 ( .A(p_input[1670]), .Z(n18394) );
  XOR U18472 ( .A(n18676), .B(n18677), .Z(n18672) );
  AND U18473 ( .A(n18678), .B(n18679), .Z(n18677) );
  XNOR U18474 ( .A(p_input[1701]), .B(n18676), .Z(n18679) );
  XNOR U18475 ( .A(n18676), .B(n18403), .Z(n18678) );
  IV U18476 ( .A(p_input[1669]), .Z(n18403) );
  XOR U18477 ( .A(n18680), .B(n18681), .Z(n18676) );
  AND U18478 ( .A(n18682), .B(n18683), .Z(n18681) );
  XNOR U18479 ( .A(p_input[1700]), .B(n18680), .Z(n18683) );
  XNOR U18480 ( .A(n18680), .B(n18412), .Z(n18682) );
  IV U18481 ( .A(p_input[1668]), .Z(n18412) );
  XOR U18482 ( .A(n18684), .B(n18685), .Z(n18680) );
  AND U18483 ( .A(n18686), .B(n18687), .Z(n18685) );
  XNOR U18484 ( .A(p_input[1699]), .B(n18684), .Z(n18687) );
  XNOR U18485 ( .A(n18684), .B(n18421), .Z(n18686) );
  IV U18486 ( .A(p_input[1667]), .Z(n18421) );
  XOR U18487 ( .A(n18688), .B(n18689), .Z(n18684) );
  AND U18488 ( .A(n18690), .B(n18691), .Z(n18689) );
  XNOR U18489 ( .A(p_input[1698]), .B(n18688), .Z(n18691) );
  XNOR U18490 ( .A(n18688), .B(n18430), .Z(n18690) );
  IV U18491 ( .A(p_input[1666]), .Z(n18430) );
  XNOR U18492 ( .A(n18692), .B(n18693), .Z(n18688) );
  AND U18493 ( .A(n18694), .B(n18695), .Z(n18693) );
  XOR U18494 ( .A(p_input[1697]), .B(n18692), .Z(n18695) );
  XNOR U18495 ( .A(p_input[1665]), .B(n18692), .Z(n18694) );
  AND U18496 ( .A(p_input[1696]), .B(n18696), .Z(n18692) );
  IV U18497 ( .A(p_input[1664]), .Z(n18696) );
  XOR U18498 ( .A(n18697), .B(n18698), .Z(n17786) );
  AND U18499 ( .A(n367), .B(n18699), .Z(n18698) );
  XNOR U18500 ( .A(n18700), .B(n18697), .Z(n18699) );
  XOR U18501 ( .A(n18701), .B(n18702), .Z(n367) );
  AND U18502 ( .A(n18703), .B(n18704), .Z(n18702) );
  XNOR U18503 ( .A(n17801), .B(n18701), .Z(n18704) );
  AND U18504 ( .A(p_input[1663]), .B(p_input[1631]), .Z(n17801) );
  XNOR U18505 ( .A(n18701), .B(n17798), .Z(n18703) );
  IV U18506 ( .A(n18705), .Z(n17798) );
  AND U18507 ( .A(p_input[1567]), .B(p_input[1599]), .Z(n18705) );
  XOR U18508 ( .A(n18706), .B(n18707), .Z(n18701) );
  AND U18509 ( .A(n18708), .B(n18709), .Z(n18707) );
  XOR U18510 ( .A(n18706), .B(n17813), .Z(n18709) );
  XNOR U18511 ( .A(p_input[1630]), .B(n18710), .Z(n17813) );
  AND U18512 ( .A(n446), .B(n18711), .Z(n18710) );
  XOR U18513 ( .A(p_input[1662]), .B(p_input[1630]), .Z(n18711) );
  XNOR U18514 ( .A(n17810), .B(n18706), .Z(n18708) );
  XOR U18515 ( .A(n18712), .B(n18713), .Z(n17810) );
  AND U18516 ( .A(n443), .B(n18714), .Z(n18713) );
  XOR U18517 ( .A(p_input[1598]), .B(p_input[1566]), .Z(n18714) );
  XOR U18518 ( .A(n18715), .B(n18716), .Z(n18706) );
  AND U18519 ( .A(n18717), .B(n18718), .Z(n18716) );
  XOR U18520 ( .A(n18715), .B(n17825), .Z(n18718) );
  XNOR U18521 ( .A(p_input[1629]), .B(n18719), .Z(n17825) );
  AND U18522 ( .A(n446), .B(n18720), .Z(n18719) );
  XOR U18523 ( .A(p_input[1661]), .B(p_input[1629]), .Z(n18720) );
  XNOR U18524 ( .A(n17822), .B(n18715), .Z(n18717) );
  XOR U18525 ( .A(n18721), .B(n18722), .Z(n17822) );
  AND U18526 ( .A(n443), .B(n18723), .Z(n18722) );
  XOR U18527 ( .A(p_input[1597]), .B(p_input[1565]), .Z(n18723) );
  XOR U18528 ( .A(n18724), .B(n18725), .Z(n18715) );
  AND U18529 ( .A(n18726), .B(n18727), .Z(n18725) );
  XOR U18530 ( .A(n18724), .B(n17837), .Z(n18727) );
  XNOR U18531 ( .A(p_input[1628]), .B(n18728), .Z(n17837) );
  AND U18532 ( .A(n446), .B(n18729), .Z(n18728) );
  XOR U18533 ( .A(p_input[1660]), .B(p_input[1628]), .Z(n18729) );
  XNOR U18534 ( .A(n17834), .B(n18724), .Z(n18726) );
  XOR U18535 ( .A(n18730), .B(n18731), .Z(n17834) );
  AND U18536 ( .A(n443), .B(n18732), .Z(n18731) );
  XOR U18537 ( .A(p_input[1596]), .B(p_input[1564]), .Z(n18732) );
  XOR U18538 ( .A(n18733), .B(n18734), .Z(n18724) );
  AND U18539 ( .A(n18735), .B(n18736), .Z(n18734) );
  XOR U18540 ( .A(n18733), .B(n17849), .Z(n18736) );
  XNOR U18541 ( .A(p_input[1627]), .B(n18737), .Z(n17849) );
  AND U18542 ( .A(n446), .B(n18738), .Z(n18737) );
  XOR U18543 ( .A(p_input[1659]), .B(p_input[1627]), .Z(n18738) );
  XNOR U18544 ( .A(n17846), .B(n18733), .Z(n18735) );
  XOR U18545 ( .A(n18739), .B(n18740), .Z(n17846) );
  AND U18546 ( .A(n443), .B(n18741), .Z(n18740) );
  XOR U18547 ( .A(p_input[1595]), .B(p_input[1563]), .Z(n18741) );
  XOR U18548 ( .A(n18742), .B(n18743), .Z(n18733) );
  AND U18549 ( .A(n18744), .B(n18745), .Z(n18743) );
  XOR U18550 ( .A(n18742), .B(n17861), .Z(n18745) );
  XNOR U18551 ( .A(p_input[1626]), .B(n18746), .Z(n17861) );
  AND U18552 ( .A(n446), .B(n18747), .Z(n18746) );
  XOR U18553 ( .A(p_input[1658]), .B(p_input[1626]), .Z(n18747) );
  XNOR U18554 ( .A(n17858), .B(n18742), .Z(n18744) );
  XOR U18555 ( .A(n18748), .B(n18749), .Z(n17858) );
  AND U18556 ( .A(n443), .B(n18750), .Z(n18749) );
  XOR U18557 ( .A(p_input[1594]), .B(p_input[1562]), .Z(n18750) );
  XOR U18558 ( .A(n18751), .B(n18752), .Z(n18742) );
  AND U18559 ( .A(n18753), .B(n18754), .Z(n18752) );
  XOR U18560 ( .A(n18751), .B(n17873), .Z(n18754) );
  XNOR U18561 ( .A(p_input[1625]), .B(n18755), .Z(n17873) );
  AND U18562 ( .A(n446), .B(n18756), .Z(n18755) );
  XOR U18563 ( .A(p_input[1657]), .B(p_input[1625]), .Z(n18756) );
  XNOR U18564 ( .A(n17870), .B(n18751), .Z(n18753) );
  XOR U18565 ( .A(n18757), .B(n18758), .Z(n17870) );
  AND U18566 ( .A(n443), .B(n18759), .Z(n18758) );
  XOR U18567 ( .A(p_input[1593]), .B(p_input[1561]), .Z(n18759) );
  XOR U18568 ( .A(n18760), .B(n18761), .Z(n18751) );
  AND U18569 ( .A(n18762), .B(n18763), .Z(n18761) );
  XOR U18570 ( .A(n18760), .B(n17885), .Z(n18763) );
  XNOR U18571 ( .A(p_input[1624]), .B(n18764), .Z(n17885) );
  AND U18572 ( .A(n446), .B(n18765), .Z(n18764) );
  XOR U18573 ( .A(p_input[1656]), .B(p_input[1624]), .Z(n18765) );
  XNOR U18574 ( .A(n17882), .B(n18760), .Z(n18762) );
  XOR U18575 ( .A(n18766), .B(n18767), .Z(n17882) );
  AND U18576 ( .A(n443), .B(n18768), .Z(n18767) );
  XOR U18577 ( .A(p_input[1592]), .B(p_input[1560]), .Z(n18768) );
  XOR U18578 ( .A(n18769), .B(n18770), .Z(n18760) );
  AND U18579 ( .A(n18771), .B(n18772), .Z(n18770) );
  XOR U18580 ( .A(n18769), .B(n17897), .Z(n18772) );
  XNOR U18581 ( .A(p_input[1623]), .B(n18773), .Z(n17897) );
  AND U18582 ( .A(n446), .B(n18774), .Z(n18773) );
  XOR U18583 ( .A(p_input[1655]), .B(p_input[1623]), .Z(n18774) );
  XNOR U18584 ( .A(n17894), .B(n18769), .Z(n18771) );
  XOR U18585 ( .A(n18775), .B(n18776), .Z(n17894) );
  AND U18586 ( .A(n443), .B(n18777), .Z(n18776) );
  XOR U18587 ( .A(p_input[1591]), .B(p_input[1559]), .Z(n18777) );
  XOR U18588 ( .A(n18778), .B(n18779), .Z(n18769) );
  AND U18589 ( .A(n18780), .B(n18781), .Z(n18779) );
  XOR U18590 ( .A(n18778), .B(n17909), .Z(n18781) );
  XNOR U18591 ( .A(p_input[1622]), .B(n18782), .Z(n17909) );
  AND U18592 ( .A(n446), .B(n18783), .Z(n18782) );
  XOR U18593 ( .A(p_input[1654]), .B(p_input[1622]), .Z(n18783) );
  XNOR U18594 ( .A(n17906), .B(n18778), .Z(n18780) );
  XOR U18595 ( .A(n18784), .B(n18785), .Z(n17906) );
  AND U18596 ( .A(n443), .B(n18786), .Z(n18785) );
  XOR U18597 ( .A(p_input[1590]), .B(p_input[1558]), .Z(n18786) );
  XOR U18598 ( .A(n18787), .B(n18788), .Z(n18778) );
  AND U18599 ( .A(n18789), .B(n18790), .Z(n18788) );
  XOR U18600 ( .A(n18787), .B(n17921), .Z(n18790) );
  XNOR U18601 ( .A(p_input[1621]), .B(n18791), .Z(n17921) );
  AND U18602 ( .A(n446), .B(n18792), .Z(n18791) );
  XOR U18603 ( .A(p_input[1653]), .B(p_input[1621]), .Z(n18792) );
  XNOR U18604 ( .A(n17918), .B(n18787), .Z(n18789) );
  XOR U18605 ( .A(n18793), .B(n18794), .Z(n17918) );
  AND U18606 ( .A(n443), .B(n18795), .Z(n18794) );
  XOR U18607 ( .A(p_input[1589]), .B(p_input[1557]), .Z(n18795) );
  XOR U18608 ( .A(n18796), .B(n18797), .Z(n18787) );
  AND U18609 ( .A(n18798), .B(n18799), .Z(n18797) );
  XOR U18610 ( .A(n18796), .B(n17933), .Z(n18799) );
  XNOR U18611 ( .A(p_input[1620]), .B(n18800), .Z(n17933) );
  AND U18612 ( .A(n446), .B(n18801), .Z(n18800) );
  XOR U18613 ( .A(p_input[1652]), .B(p_input[1620]), .Z(n18801) );
  XNOR U18614 ( .A(n17930), .B(n18796), .Z(n18798) );
  XOR U18615 ( .A(n18802), .B(n18803), .Z(n17930) );
  AND U18616 ( .A(n443), .B(n18804), .Z(n18803) );
  XOR U18617 ( .A(p_input[1588]), .B(p_input[1556]), .Z(n18804) );
  XOR U18618 ( .A(n18805), .B(n18806), .Z(n18796) );
  AND U18619 ( .A(n18807), .B(n18808), .Z(n18806) );
  XOR U18620 ( .A(n18805), .B(n17945), .Z(n18808) );
  XNOR U18621 ( .A(p_input[1619]), .B(n18809), .Z(n17945) );
  AND U18622 ( .A(n446), .B(n18810), .Z(n18809) );
  XOR U18623 ( .A(p_input[1651]), .B(p_input[1619]), .Z(n18810) );
  XNOR U18624 ( .A(n17942), .B(n18805), .Z(n18807) );
  XOR U18625 ( .A(n18811), .B(n18812), .Z(n17942) );
  AND U18626 ( .A(n443), .B(n18813), .Z(n18812) );
  XOR U18627 ( .A(p_input[1587]), .B(p_input[1555]), .Z(n18813) );
  XOR U18628 ( .A(n18814), .B(n18815), .Z(n18805) );
  AND U18629 ( .A(n18816), .B(n18817), .Z(n18815) );
  XOR U18630 ( .A(n18814), .B(n17957), .Z(n18817) );
  XNOR U18631 ( .A(p_input[1618]), .B(n18818), .Z(n17957) );
  AND U18632 ( .A(n446), .B(n18819), .Z(n18818) );
  XOR U18633 ( .A(p_input[1650]), .B(p_input[1618]), .Z(n18819) );
  XNOR U18634 ( .A(n17954), .B(n18814), .Z(n18816) );
  XOR U18635 ( .A(n18820), .B(n18821), .Z(n17954) );
  AND U18636 ( .A(n443), .B(n18822), .Z(n18821) );
  XOR U18637 ( .A(p_input[1586]), .B(p_input[1554]), .Z(n18822) );
  XOR U18638 ( .A(n18823), .B(n18824), .Z(n18814) );
  AND U18639 ( .A(n18825), .B(n18826), .Z(n18824) );
  XOR U18640 ( .A(n18823), .B(n17969), .Z(n18826) );
  XNOR U18641 ( .A(p_input[1617]), .B(n18827), .Z(n17969) );
  AND U18642 ( .A(n446), .B(n18828), .Z(n18827) );
  XOR U18643 ( .A(p_input[1649]), .B(p_input[1617]), .Z(n18828) );
  XNOR U18644 ( .A(n17966), .B(n18823), .Z(n18825) );
  XOR U18645 ( .A(n18829), .B(n18830), .Z(n17966) );
  AND U18646 ( .A(n443), .B(n18831), .Z(n18830) );
  XOR U18647 ( .A(p_input[1585]), .B(p_input[1553]), .Z(n18831) );
  XOR U18648 ( .A(n18832), .B(n18833), .Z(n18823) );
  AND U18649 ( .A(n18834), .B(n18835), .Z(n18833) );
  XOR U18650 ( .A(n18832), .B(n17981), .Z(n18835) );
  XNOR U18651 ( .A(p_input[1616]), .B(n18836), .Z(n17981) );
  AND U18652 ( .A(n446), .B(n18837), .Z(n18836) );
  XOR U18653 ( .A(p_input[1648]), .B(p_input[1616]), .Z(n18837) );
  XNOR U18654 ( .A(n17978), .B(n18832), .Z(n18834) );
  XOR U18655 ( .A(n18838), .B(n18839), .Z(n17978) );
  AND U18656 ( .A(n443), .B(n18840), .Z(n18839) );
  XOR U18657 ( .A(p_input[1584]), .B(p_input[1552]), .Z(n18840) );
  XOR U18658 ( .A(n18841), .B(n18842), .Z(n18832) );
  AND U18659 ( .A(n18843), .B(n18844), .Z(n18842) );
  XOR U18660 ( .A(n18841), .B(n17993), .Z(n18844) );
  XNOR U18661 ( .A(p_input[1615]), .B(n18845), .Z(n17993) );
  AND U18662 ( .A(n446), .B(n18846), .Z(n18845) );
  XOR U18663 ( .A(p_input[1647]), .B(p_input[1615]), .Z(n18846) );
  XNOR U18664 ( .A(n17990), .B(n18841), .Z(n18843) );
  XOR U18665 ( .A(n18847), .B(n18848), .Z(n17990) );
  AND U18666 ( .A(n443), .B(n18849), .Z(n18848) );
  XOR U18667 ( .A(p_input[1583]), .B(p_input[1551]), .Z(n18849) );
  XOR U18668 ( .A(n18850), .B(n18851), .Z(n18841) );
  AND U18669 ( .A(n18852), .B(n18853), .Z(n18851) );
  XOR U18670 ( .A(n18850), .B(n18005), .Z(n18853) );
  XNOR U18671 ( .A(p_input[1614]), .B(n18854), .Z(n18005) );
  AND U18672 ( .A(n446), .B(n18855), .Z(n18854) );
  XOR U18673 ( .A(p_input[1646]), .B(p_input[1614]), .Z(n18855) );
  XNOR U18674 ( .A(n18002), .B(n18850), .Z(n18852) );
  XOR U18675 ( .A(n18856), .B(n18857), .Z(n18002) );
  AND U18676 ( .A(n443), .B(n18858), .Z(n18857) );
  XOR U18677 ( .A(p_input[1582]), .B(p_input[1550]), .Z(n18858) );
  XOR U18678 ( .A(n18859), .B(n18860), .Z(n18850) );
  AND U18679 ( .A(n18861), .B(n18862), .Z(n18860) );
  XOR U18680 ( .A(n18859), .B(n18017), .Z(n18862) );
  XNOR U18681 ( .A(p_input[1613]), .B(n18863), .Z(n18017) );
  AND U18682 ( .A(n446), .B(n18864), .Z(n18863) );
  XOR U18683 ( .A(p_input[1645]), .B(p_input[1613]), .Z(n18864) );
  XNOR U18684 ( .A(n18014), .B(n18859), .Z(n18861) );
  XOR U18685 ( .A(n18865), .B(n18866), .Z(n18014) );
  AND U18686 ( .A(n443), .B(n18867), .Z(n18866) );
  XOR U18687 ( .A(p_input[1581]), .B(p_input[1549]), .Z(n18867) );
  XOR U18688 ( .A(n18868), .B(n18869), .Z(n18859) );
  AND U18689 ( .A(n18870), .B(n18871), .Z(n18869) );
  XOR U18690 ( .A(n18868), .B(n18029), .Z(n18871) );
  XNOR U18691 ( .A(p_input[1612]), .B(n18872), .Z(n18029) );
  AND U18692 ( .A(n446), .B(n18873), .Z(n18872) );
  XOR U18693 ( .A(p_input[1644]), .B(p_input[1612]), .Z(n18873) );
  XNOR U18694 ( .A(n18026), .B(n18868), .Z(n18870) );
  XOR U18695 ( .A(n18874), .B(n18875), .Z(n18026) );
  AND U18696 ( .A(n443), .B(n18876), .Z(n18875) );
  XOR U18697 ( .A(p_input[1580]), .B(p_input[1548]), .Z(n18876) );
  XOR U18698 ( .A(n18877), .B(n18878), .Z(n18868) );
  AND U18699 ( .A(n18879), .B(n18880), .Z(n18878) );
  XOR U18700 ( .A(n18877), .B(n18041), .Z(n18880) );
  XNOR U18701 ( .A(p_input[1611]), .B(n18881), .Z(n18041) );
  AND U18702 ( .A(n446), .B(n18882), .Z(n18881) );
  XOR U18703 ( .A(p_input[1643]), .B(p_input[1611]), .Z(n18882) );
  XNOR U18704 ( .A(n18038), .B(n18877), .Z(n18879) );
  XOR U18705 ( .A(n18883), .B(n18884), .Z(n18038) );
  AND U18706 ( .A(n443), .B(n18885), .Z(n18884) );
  XOR U18707 ( .A(p_input[1579]), .B(p_input[1547]), .Z(n18885) );
  XOR U18708 ( .A(n18886), .B(n18887), .Z(n18877) );
  AND U18709 ( .A(n18888), .B(n18889), .Z(n18887) );
  XOR U18710 ( .A(n18886), .B(n18053), .Z(n18889) );
  XNOR U18711 ( .A(p_input[1610]), .B(n18890), .Z(n18053) );
  AND U18712 ( .A(n446), .B(n18891), .Z(n18890) );
  XOR U18713 ( .A(p_input[1642]), .B(p_input[1610]), .Z(n18891) );
  XNOR U18714 ( .A(n18050), .B(n18886), .Z(n18888) );
  XOR U18715 ( .A(n18892), .B(n18893), .Z(n18050) );
  AND U18716 ( .A(n443), .B(n18894), .Z(n18893) );
  XOR U18717 ( .A(p_input[1578]), .B(p_input[1546]), .Z(n18894) );
  XOR U18718 ( .A(n18895), .B(n18896), .Z(n18886) );
  AND U18719 ( .A(n18897), .B(n18898), .Z(n18896) );
  XOR U18720 ( .A(n18895), .B(n18065), .Z(n18898) );
  XNOR U18721 ( .A(p_input[1609]), .B(n18899), .Z(n18065) );
  AND U18722 ( .A(n446), .B(n18900), .Z(n18899) );
  XOR U18723 ( .A(p_input[1641]), .B(p_input[1609]), .Z(n18900) );
  XNOR U18724 ( .A(n18062), .B(n18895), .Z(n18897) );
  XOR U18725 ( .A(n18901), .B(n18902), .Z(n18062) );
  AND U18726 ( .A(n443), .B(n18903), .Z(n18902) );
  XOR U18727 ( .A(p_input[1577]), .B(p_input[1545]), .Z(n18903) );
  XOR U18728 ( .A(n18904), .B(n18905), .Z(n18895) );
  AND U18729 ( .A(n18906), .B(n18907), .Z(n18905) );
  XOR U18730 ( .A(n18904), .B(n18077), .Z(n18907) );
  XNOR U18731 ( .A(p_input[1608]), .B(n18908), .Z(n18077) );
  AND U18732 ( .A(n446), .B(n18909), .Z(n18908) );
  XOR U18733 ( .A(p_input[1640]), .B(p_input[1608]), .Z(n18909) );
  XNOR U18734 ( .A(n18074), .B(n18904), .Z(n18906) );
  XOR U18735 ( .A(n18910), .B(n18911), .Z(n18074) );
  AND U18736 ( .A(n443), .B(n18912), .Z(n18911) );
  XOR U18737 ( .A(p_input[1576]), .B(p_input[1544]), .Z(n18912) );
  XOR U18738 ( .A(n18913), .B(n18914), .Z(n18904) );
  AND U18739 ( .A(n18915), .B(n18916), .Z(n18914) );
  XOR U18740 ( .A(n18913), .B(n18089), .Z(n18916) );
  XNOR U18741 ( .A(p_input[1607]), .B(n18917), .Z(n18089) );
  AND U18742 ( .A(n446), .B(n18918), .Z(n18917) );
  XOR U18743 ( .A(p_input[1639]), .B(p_input[1607]), .Z(n18918) );
  XNOR U18744 ( .A(n18086), .B(n18913), .Z(n18915) );
  XOR U18745 ( .A(n18919), .B(n18920), .Z(n18086) );
  AND U18746 ( .A(n443), .B(n18921), .Z(n18920) );
  XOR U18747 ( .A(p_input[1575]), .B(p_input[1543]), .Z(n18921) );
  XOR U18748 ( .A(n18922), .B(n18923), .Z(n18913) );
  AND U18749 ( .A(n18924), .B(n18925), .Z(n18923) );
  XOR U18750 ( .A(n18922), .B(n18101), .Z(n18925) );
  XNOR U18751 ( .A(p_input[1606]), .B(n18926), .Z(n18101) );
  AND U18752 ( .A(n446), .B(n18927), .Z(n18926) );
  XOR U18753 ( .A(p_input[1638]), .B(p_input[1606]), .Z(n18927) );
  XNOR U18754 ( .A(n18098), .B(n18922), .Z(n18924) );
  XOR U18755 ( .A(n18928), .B(n18929), .Z(n18098) );
  AND U18756 ( .A(n443), .B(n18930), .Z(n18929) );
  XOR U18757 ( .A(p_input[1574]), .B(p_input[1542]), .Z(n18930) );
  XOR U18758 ( .A(n18931), .B(n18932), .Z(n18922) );
  AND U18759 ( .A(n18933), .B(n18934), .Z(n18932) );
  XOR U18760 ( .A(n18931), .B(n18113), .Z(n18934) );
  XNOR U18761 ( .A(p_input[1605]), .B(n18935), .Z(n18113) );
  AND U18762 ( .A(n446), .B(n18936), .Z(n18935) );
  XOR U18763 ( .A(p_input[1637]), .B(p_input[1605]), .Z(n18936) );
  XNOR U18764 ( .A(n18110), .B(n18931), .Z(n18933) );
  XOR U18765 ( .A(n18937), .B(n18938), .Z(n18110) );
  AND U18766 ( .A(n443), .B(n18939), .Z(n18938) );
  XOR U18767 ( .A(p_input[1573]), .B(p_input[1541]), .Z(n18939) );
  XOR U18768 ( .A(n18940), .B(n18941), .Z(n18931) );
  AND U18769 ( .A(n18942), .B(n18943), .Z(n18941) );
  XOR U18770 ( .A(n18940), .B(n18125), .Z(n18943) );
  XNOR U18771 ( .A(p_input[1604]), .B(n18944), .Z(n18125) );
  AND U18772 ( .A(n446), .B(n18945), .Z(n18944) );
  XOR U18773 ( .A(p_input[1636]), .B(p_input[1604]), .Z(n18945) );
  XNOR U18774 ( .A(n18122), .B(n18940), .Z(n18942) );
  XOR U18775 ( .A(n18946), .B(n18947), .Z(n18122) );
  AND U18776 ( .A(n443), .B(n18948), .Z(n18947) );
  XOR U18777 ( .A(p_input[1572]), .B(p_input[1540]), .Z(n18948) );
  XOR U18778 ( .A(n18949), .B(n18950), .Z(n18940) );
  AND U18779 ( .A(n18951), .B(n18952), .Z(n18950) );
  XOR U18780 ( .A(n18949), .B(n18137), .Z(n18952) );
  XNOR U18781 ( .A(p_input[1603]), .B(n18953), .Z(n18137) );
  AND U18782 ( .A(n446), .B(n18954), .Z(n18953) );
  XOR U18783 ( .A(p_input[1635]), .B(p_input[1603]), .Z(n18954) );
  XNOR U18784 ( .A(n18134), .B(n18949), .Z(n18951) );
  XOR U18785 ( .A(n18955), .B(n18956), .Z(n18134) );
  AND U18786 ( .A(n443), .B(n18957), .Z(n18956) );
  XOR U18787 ( .A(p_input[1571]), .B(p_input[1539]), .Z(n18957) );
  XOR U18788 ( .A(n18958), .B(n18959), .Z(n18949) );
  AND U18789 ( .A(n18960), .B(n18961), .Z(n18959) );
  XOR U18790 ( .A(n18149), .B(n18958), .Z(n18961) );
  XNOR U18791 ( .A(p_input[1602]), .B(n18962), .Z(n18149) );
  AND U18792 ( .A(n446), .B(n18963), .Z(n18962) );
  XOR U18793 ( .A(p_input[1634]), .B(p_input[1602]), .Z(n18963) );
  XNOR U18794 ( .A(n18958), .B(n18146), .Z(n18960) );
  XOR U18795 ( .A(n18964), .B(n18965), .Z(n18146) );
  AND U18796 ( .A(n443), .B(n18966), .Z(n18965) );
  XOR U18797 ( .A(p_input[1570]), .B(p_input[1538]), .Z(n18966) );
  XOR U18798 ( .A(n18967), .B(n18968), .Z(n18958) );
  AND U18799 ( .A(n18969), .B(n18970), .Z(n18968) );
  XNOR U18800 ( .A(n18971), .B(n18162), .Z(n18970) );
  XNOR U18801 ( .A(p_input[1601]), .B(n18972), .Z(n18162) );
  AND U18802 ( .A(n446), .B(n18973), .Z(n18972) );
  XNOR U18803 ( .A(p_input[1633]), .B(n18974), .Z(n18973) );
  IV U18804 ( .A(p_input[1601]), .Z(n18974) );
  XNOR U18805 ( .A(n18159), .B(n18967), .Z(n18969) );
  XNOR U18806 ( .A(p_input[1537]), .B(n18975), .Z(n18159) );
  AND U18807 ( .A(n443), .B(n18976), .Z(n18975) );
  XOR U18808 ( .A(p_input[1569]), .B(p_input[1537]), .Z(n18976) );
  IV U18809 ( .A(n18971), .Z(n18967) );
  AND U18810 ( .A(n18697), .B(n18700), .Z(n18971) );
  XOR U18811 ( .A(p_input[1600]), .B(n18977), .Z(n18700) );
  AND U18812 ( .A(n446), .B(n18978), .Z(n18977) );
  XOR U18813 ( .A(p_input[1632]), .B(p_input[1600]), .Z(n18978) );
  XOR U18814 ( .A(n18979), .B(n18980), .Z(n446) );
  AND U18815 ( .A(n18981), .B(n18982), .Z(n18980) );
  XNOR U18816 ( .A(p_input[1663]), .B(n18979), .Z(n18982) );
  XOR U18817 ( .A(n18979), .B(p_input[1631]), .Z(n18981) );
  XOR U18818 ( .A(n18983), .B(n18984), .Z(n18979) );
  AND U18819 ( .A(n18985), .B(n18986), .Z(n18984) );
  XNOR U18820 ( .A(p_input[1662]), .B(n18983), .Z(n18986) );
  XOR U18821 ( .A(n18983), .B(p_input[1630]), .Z(n18985) );
  XOR U18822 ( .A(n18987), .B(n18988), .Z(n18983) );
  AND U18823 ( .A(n18989), .B(n18990), .Z(n18988) );
  XNOR U18824 ( .A(p_input[1661]), .B(n18987), .Z(n18990) );
  XOR U18825 ( .A(n18987), .B(p_input[1629]), .Z(n18989) );
  XOR U18826 ( .A(n18991), .B(n18992), .Z(n18987) );
  AND U18827 ( .A(n18993), .B(n18994), .Z(n18992) );
  XNOR U18828 ( .A(p_input[1660]), .B(n18991), .Z(n18994) );
  XOR U18829 ( .A(n18991), .B(p_input[1628]), .Z(n18993) );
  XOR U18830 ( .A(n18995), .B(n18996), .Z(n18991) );
  AND U18831 ( .A(n18997), .B(n18998), .Z(n18996) );
  XNOR U18832 ( .A(p_input[1659]), .B(n18995), .Z(n18998) );
  XOR U18833 ( .A(n18995), .B(p_input[1627]), .Z(n18997) );
  XOR U18834 ( .A(n18999), .B(n19000), .Z(n18995) );
  AND U18835 ( .A(n19001), .B(n19002), .Z(n19000) );
  XNOR U18836 ( .A(p_input[1658]), .B(n18999), .Z(n19002) );
  XOR U18837 ( .A(n18999), .B(p_input[1626]), .Z(n19001) );
  XOR U18838 ( .A(n19003), .B(n19004), .Z(n18999) );
  AND U18839 ( .A(n19005), .B(n19006), .Z(n19004) );
  XNOR U18840 ( .A(p_input[1657]), .B(n19003), .Z(n19006) );
  XOR U18841 ( .A(n19003), .B(p_input[1625]), .Z(n19005) );
  XOR U18842 ( .A(n19007), .B(n19008), .Z(n19003) );
  AND U18843 ( .A(n19009), .B(n19010), .Z(n19008) );
  XNOR U18844 ( .A(p_input[1656]), .B(n19007), .Z(n19010) );
  XOR U18845 ( .A(n19007), .B(p_input[1624]), .Z(n19009) );
  XOR U18846 ( .A(n19011), .B(n19012), .Z(n19007) );
  AND U18847 ( .A(n19013), .B(n19014), .Z(n19012) );
  XNOR U18848 ( .A(p_input[1655]), .B(n19011), .Z(n19014) );
  XOR U18849 ( .A(n19011), .B(p_input[1623]), .Z(n19013) );
  XOR U18850 ( .A(n19015), .B(n19016), .Z(n19011) );
  AND U18851 ( .A(n19017), .B(n19018), .Z(n19016) );
  XNOR U18852 ( .A(p_input[1654]), .B(n19015), .Z(n19018) );
  XOR U18853 ( .A(n19015), .B(p_input[1622]), .Z(n19017) );
  XOR U18854 ( .A(n19019), .B(n19020), .Z(n19015) );
  AND U18855 ( .A(n19021), .B(n19022), .Z(n19020) );
  XNOR U18856 ( .A(p_input[1653]), .B(n19019), .Z(n19022) );
  XOR U18857 ( .A(n19019), .B(p_input[1621]), .Z(n19021) );
  XOR U18858 ( .A(n19023), .B(n19024), .Z(n19019) );
  AND U18859 ( .A(n19025), .B(n19026), .Z(n19024) );
  XNOR U18860 ( .A(p_input[1652]), .B(n19023), .Z(n19026) );
  XOR U18861 ( .A(n19023), .B(p_input[1620]), .Z(n19025) );
  XOR U18862 ( .A(n19027), .B(n19028), .Z(n19023) );
  AND U18863 ( .A(n19029), .B(n19030), .Z(n19028) );
  XNOR U18864 ( .A(p_input[1651]), .B(n19027), .Z(n19030) );
  XOR U18865 ( .A(n19027), .B(p_input[1619]), .Z(n19029) );
  XOR U18866 ( .A(n19031), .B(n19032), .Z(n19027) );
  AND U18867 ( .A(n19033), .B(n19034), .Z(n19032) );
  XNOR U18868 ( .A(p_input[1650]), .B(n19031), .Z(n19034) );
  XOR U18869 ( .A(n19031), .B(p_input[1618]), .Z(n19033) );
  XOR U18870 ( .A(n19035), .B(n19036), .Z(n19031) );
  AND U18871 ( .A(n19037), .B(n19038), .Z(n19036) );
  XNOR U18872 ( .A(p_input[1649]), .B(n19035), .Z(n19038) );
  XOR U18873 ( .A(n19035), .B(p_input[1617]), .Z(n19037) );
  XOR U18874 ( .A(n19039), .B(n19040), .Z(n19035) );
  AND U18875 ( .A(n19041), .B(n19042), .Z(n19040) );
  XNOR U18876 ( .A(p_input[1648]), .B(n19039), .Z(n19042) );
  XOR U18877 ( .A(n19039), .B(p_input[1616]), .Z(n19041) );
  XOR U18878 ( .A(n19043), .B(n19044), .Z(n19039) );
  AND U18879 ( .A(n19045), .B(n19046), .Z(n19044) );
  XNOR U18880 ( .A(p_input[1647]), .B(n19043), .Z(n19046) );
  XOR U18881 ( .A(n19043), .B(p_input[1615]), .Z(n19045) );
  XOR U18882 ( .A(n19047), .B(n19048), .Z(n19043) );
  AND U18883 ( .A(n19049), .B(n19050), .Z(n19048) );
  XNOR U18884 ( .A(p_input[1646]), .B(n19047), .Z(n19050) );
  XOR U18885 ( .A(n19047), .B(p_input[1614]), .Z(n19049) );
  XOR U18886 ( .A(n19051), .B(n19052), .Z(n19047) );
  AND U18887 ( .A(n19053), .B(n19054), .Z(n19052) );
  XNOR U18888 ( .A(p_input[1645]), .B(n19051), .Z(n19054) );
  XOR U18889 ( .A(n19051), .B(p_input[1613]), .Z(n19053) );
  XOR U18890 ( .A(n19055), .B(n19056), .Z(n19051) );
  AND U18891 ( .A(n19057), .B(n19058), .Z(n19056) );
  XNOR U18892 ( .A(p_input[1644]), .B(n19055), .Z(n19058) );
  XOR U18893 ( .A(n19055), .B(p_input[1612]), .Z(n19057) );
  XOR U18894 ( .A(n19059), .B(n19060), .Z(n19055) );
  AND U18895 ( .A(n19061), .B(n19062), .Z(n19060) );
  XNOR U18896 ( .A(p_input[1643]), .B(n19059), .Z(n19062) );
  XOR U18897 ( .A(n19059), .B(p_input[1611]), .Z(n19061) );
  XOR U18898 ( .A(n19063), .B(n19064), .Z(n19059) );
  AND U18899 ( .A(n19065), .B(n19066), .Z(n19064) );
  XNOR U18900 ( .A(p_input[1642]), .B(n19063), .Z(n19066) );
  XOR U18901 ( .A(n19063), .B(p_input[1610]), .Z(n19065) );
  XOR U18902 ( .A(n19067), .B(n19068), .Z(n19063) );
  AND U18903 ( .A(n19069), .B(n19070), .Z(n19068) );
  XNOR U18904 ( .A(p_input[1641]), .B(n19067), .Z(n19070) );
  XOR U18905 ( .A(n19067), .B(p_input[1609]), .Z(n19069) );
  XOR U18906 ( .A(n19071), .B(n19072), .Z(n19067) );
  AND U18907 ( .A(n19073), .B(n19074), .Z(n19072) );
  XNOR U18908 ( .A(p_input[1640]), .B(n19071), .Z(n19074) );
  XOR U18909 ( .A(n19071), .B(p_input[1608]), .Z(n19073) );
  XOR U18910 ( .A(n19075), .B(n19076), .Z(n19071) );
  AND U18911 ( .A(n19077), .B(n19078), .Z(n19076) );
  XNOR U18912 ( .A(p_input[1639]), .B(n19075), .Z(n19078) );
  XOR U18913 ( .A(n19075), .B(p_input[1607]), .Z(n19077) );
  XOR U18914 ( .A(n19079), .B(n19080), .Z(n19075) );
  AND U18915 ( .A(n19081), .B(n19082), .Z(n19080) );
  XNOR U18916 ( .A(p_input[1638]), .B(n19079), .Z(n19082) );
  XOR U18917 ( .A(n19079), .B(p_input[1606]), .Z(n19081) );
  XOR U18918 ( .A(n19083), .B(n19084), .Z(n19079) );
  AND U18919 ( .A(n19085), .B(n19086), .Z(n19084) );
  XNOR U18920 ( .A(p_input[1637]), .B(n19083), .Z(n19086) );
  XOR U18921 ( .A(n19083), .B(p_input[1605]), .Z(n19085) );
  XOR U18922 ( .A(n19087), .B(n19088), .Z(n19083) );
  AND U18923 ( .A(n19089), .B(n19090), .Z(n19088) );
  XNOR U18924 ( .A(p_input[1636]), .B(n19087), .Z(n19090) );
  XOR U18925 ( .A(n19087), .B(p_input[1604]), .Z(n19089) );
  XOR U18926 ( .A(n19091), .B(n19092), .Z(n19087) );
  AND U18927 ( .A(n19093), .B(n19094), .Z(n19092) );
  XNOR U18928 ( .A(p_input[1635]), .B(n19091), .Z(n19094) );
  XOR U18929 ( .A(n19091), .B(p_input[1603]), .Z(n19093) );
  XOR U18930 ( .A(n19095), .B(n19096), .Z(n19091) );
  AND U18931 ( .A(n19097), .B(n19098), .Z(n19096) );
  XNOR U18932 ( .A(p_input[1634]), .B(n19095), .Z(n19098) );
  XOR U18933 ( .A(n19095), .B(p_input[1602]), .Z(n19097) );
  XNOR U18934 ( .A(n19099), .B(n19100), .Z(n19095) );
  AND U18935 ( .A(n19101), .B(n19102), .Z(n19100) );
  XOR U18936 ( .A(p_input[1633]), .B(n19099), .Z(n19102) );
  XNOR U18937 ( .A(p_input[1601]), .B(n19099), .Z(n19101) );
  AND U18938 ( .A(p_input[1632]), .B(n19103), .Z(n19099) );
  IV U18939 ( .A(p_input[1600]), .Z(n19103) );
  XNOR U18940 ( .A(p_input[1536]), .B(n19104), .Z(n18697) );
  AND U18941 ( .A(n443), .B(n19105), .Z(n19104) );
  XOR U18942 ( .A(p_input[1568]), .B(p_input[1536]), .Z(n19105) );
  XOR U18943 ( .A(n19106), .B(n19107), .Z(n443) );
  AND U18944 ( .A(n19108), .B(n19109), .Z(n19107) );
  XNOR U18945 ( .A(p_input[1599]), .B(n19106), .Z(n19109) );
  XOR U18946 ( .A(n19106), .B(p_input[1567]), .Z(n19108) );
  XOR U18947 ( .A(n19110), .B(n19111), .Z(n19106) );
  AND U18948 ( .A(n19112), .B(n19113), .Z(n19111) );
  XNOR U18949 ( .A(p_input[1598]), .B(n19110), .Z(n19113) );
  XNOR U18950 ( .A(n19110), .B(n18712), .Z(n19112) );
  IV U18951 ( .A(p_input[1566]), .Z(n18712) );
  XOR U18952 ( .A(n19114), .B(n19115), .Z(n19110) );
  AND U18953 ( .A(n19116), .B(n19117), .Z(n19115) );
  XNOR U18954 ( .A(p_input[1597]), .B(n19114), .Z(n19117) );
  XNOR U18955 ( .A(n19114), .B(n18721), .Z(n19116) );
  IV U18956 ( .A(p_input[1565]), .Z(n18721) );
  XOR U18957 ( .A(n19118), .B(n19119), .Z(n19114) );
  AND U18958 ( .A(n19120), .B(n19121), .Z(n19119) );
  XNOR U18959 ( .A(p_input[1596]), .B(n19118), .Z(n19121) );
  XNOR U18960 ( .A(n19118), .B(n18730), .Z(n19120) );
  IV U18961 ( .A(p_input[1564]), .Z(n18730) );
  XOR U18962 ( .A(n19122), .B(n19123), .Z(n19118) );
  AND U18963 ( .A(n19124), .B(n19125), .Z(n19123) );
  XNOR U18964 ( .A(p_input[1595]), .B(n19122), .Z(n19125) );
  XNOR U18965 ( .A(n19122), .B(n18739), .Z(n19124) );
  IV U18966 ( .A(p_input[1563]), .Z(n18739) );
  XOR U18967 ( .A(n19126), .B(n19127), .Z(n19122) );
  AND U18968 ( .A(n19128), .B(n19129), .Z(n19127) );
  XNOR U18969 ( .A(p_input[1594]), .B(n19126), .Z(n19129) );
  XNOR U18970 ( .A(n19126), .B(n18748), .Z(n19128) );
  IV U18971 ( .A(p_input[1562]), .Z(n18748) );
  XOR U18972 ( .A(n19130), .B(n19131), .Z(n19126) );
  AND U18973 ( .A(n19132), .B(n19133), .Z(n19131) );
  XNOR U18974 ( .A(p_input[1593]), .B(n19130), .Z(n19133) );
  XNOR U18975 ( .A(n19130), .B(n18757), .Z(n19132) );
  IV U18976 ( .A(p_input[1561]), .Z(n18757) );
  XOR U18977 ( .A(n19134), .B(n19135), .Z(n19130) );
  AND U18978 ( .A(n19136), .B(n19137), .Z(n19135) );
  XNOR U18979 ( .A(p_input[1592]), .B(n19134), .Z(n19137) );
  XNOR U18980 ( .A(n19134), .B(n18766), .Z(n19136) );
  IV U18981 ( .A(p_input[1560]), .Z(n18766) );
  XOR U18982 ( .A(n19138), .B(n19139), .Z(n19134) );
  AND U18983 ( .A(n19140), .B(n19141), .Z(n19139) );
  XNOR U18984 ( .A(p_input[1591]), .B(n19138), .Z(n19141) );
  XNOR U18985 ( .A(n19138), .B(n18775), .Z(n19140) );
  IV U18986 ( .A(p_input[1559]), .Z(n18775) );
  XOR U18987 ( .A(n19142), .B(n19143), .Z(n19138) );
  AND U18988 ( .A(n19144), .B(n19145), .Z(n19143) );
  XNOR U18989 ( .A(p_input[1590]), .B(n19142), .Z(n19145) );
  XNOR U18990 ( .A(n19142), .B(n18784), .Z(n19144) );
  IV U18991 ( .A(p_input[1558]), .Z(n18784) );
  XOR U18992 ( .A(n19146), .B(n19147), .Z(n19142) );
  AND U18993 ( .A(n19148), .B(n19149), .Z(n19147) );
  XNOR U18994 ( .A(p_input[1589]), .B(n19146), .Z(n19149) );
  XNOR U18995 ( .A(n19146), .B(n18793), .Z(n19148) );
  IV U18996 ( .A(p_input[1557]), .Z(n18793) );
  XOR U18997 ( .A(n19150), .B(n19151), .Z(n19146) );
  AND U18998 ( .A(n19152), .B(n19153), .Z(n19151) );
  XNOR U18999 ( .A(p_input[1588]), .B(n19150), .Z(n19153) );
  XNOR U19000 ( .A(n19150), .B(n18802), .Z(n19152) );
  IV U19001 ( .A(p_input[1556]), .Z(n18802) );
  XOR U19002 ( .A(n19154), .B(n19155), .Z(n19150) );
  AND U19003 ( .A(n19156), .B(n19157), .Z(n19155) );
  XNOR U19004 ( .A(p_input[1587]), .B(n19154), .Z(n19157) );
  XNOR U19005 ( .A(n19154), .B(n18811), .Z(n19156) );
  IV U19006 ( .A(p_input[1555]), .Z(n18811) );
  XOR U19007 ( .A(n19158), .B(n19159), .Z(n19154) );
  AND U19008 ( .A(n19160), .B(n19161), .Z(n19159) );
  XNOR U19009 ( .A(p_input[1586]), .B(n19158), .Z(n19161) );
  XNOR U19010 ( .A(n19158), .B(n18820), .Z(n19160) );
  IV U19011 ( .A(p_input[1554]), .Z(n18820) );
  XOR U19012 ( .A(n19162), .B(n19163), .Z(n19158) );
  AND U19013 ( .A(n19164), .B(n19165), .Z(n19163) );
  XNOR U19014 ( .A(p_input[1585]), .B(n19162), .Z(n19165) );
  XNOR U19015 ( .A(n19162), .B(n18829), .Z(n19164) );
  IV U19016 ( .A(p_input[1553]), .Z(n18829) );
  XOR U19017 ( .A(n19166), .B(n19167), .Z(n19162) );
  AND U19018 ( .A(n19168), .B(n19169), .Z(n19167) );
  XNOR U19019 ( .A(p_input[1584]), .B(n19166), .Z(n19169) );
  XNOR U19020 ( .A(n19166), .B(n18838), .Z(n19168) );
  IV U19021 ( .A(p_input[1552]), .Z(n18838) );
  XOR U19022 ( .A(n19170), .B(n19171), .Z(n19166) );
  AND U19023 ( .A(n19172), .B(n19173), .Z(n19171) );
  XNOR U19024 ( .A(p_input[1583]), .B(n19170), .Z(n19173) );
  XNOR U19025 ( .A(n19170), .B(n18847), .Z(n19172) );
  IV U19026 ( .A(p_input[1551]), .Z(n18847) );
  XOR U19027 ( .A(n19174), .B(n19175), .Z(n19170) );
  AND U19028 ( .A(n19176), .B(n19177), .Z(n19175) );
  XNOR U19029 ( .A(p_input[1582]), .B(n19174), .Z(n19177) );
  XNOR U19030 ( .A(n19174), .B(n18856), .Z(n19176) );
  IV U19031 ( .A(p_input[1550]), .Z(n18856) );
  XOR U19032 ( .A(n19178), .B(n19179), .Z(n19174) );
  AND U19033 ( .A(n19180), .B(n19181), .Z(n19179) );
  XNOR U19034 ( .A(p_input[1581]), .B(n19178), .Z(n19181) );
  XNOR U19035 ( .A(n19178), .B(n18865), .Z(n19180) );
  IV U19036 ( .A(p_input[1549]), .Z(n18865) );
  XOR U19037 ( .A(n19182), .B(n19183), .Z(n19178) );
  AND U19038 ( .A(n19184), .B(n19185), .Z(n19183) );
  XNOR U19039 ( .A(p_input[1580]), .B(n19182), .Z(n19185) );
  XNOR U19040 ( .A(n19182), .B(n18874), .Z(n19184) );
  IV U19041 ( .A(p_input[1548]), .Z(n18874) );
  XOR U19042 ( .A(n19186), .B(n19187), .Z(n19182) );
  AND U19043 ( .A(n19188), .B(n19189), .Z(n19187) );
  XNOR U19044 ( .A(p_input[1579]), .B(n19186), .Z(n19189) );
  XNOR U19045 ( .A(n19186), .B(n18883), .Z(n19188) );
  IV U19046 ( .A(p_input[1547]), .Z(n18883) );
  XOR U19047 ( .A(n19190), .B(n19191), .Z(n19186) );
  AND U19048 ( .A(n19192), .B(n19193), .Z(n19191) );
  XNOR U19049 ( .A(p_input[1578]), .B(n19190), .Z(n19193) );
  XNOR U19050 ( .A(n19190), .B(n18892), .Z(n19192) );
  IV U19051 ( .A(p_input[1546]), .Z(n18892) );
  XOR U19052 ( .A(n19194), .B(n19195), .Z(n19190) );
  AND U19053 ( .A(n19196), .B(n19197), .Z(n19195) );
  XNOR U19054 ( .A(p_input[1577]), .B(n19194), .Z(n19197) );
  XNOR U19055 ( .A(n19194), .B(n18901), .Z(n19196) );
  IV U19056 ( .A(p_input[1545]), .Z(n18901) );
  XOR U19057 ( .A(n19198), .B(n19199), .Z(n19194) );
  AND U19058 ( .A(n19200), .B(n19201), .Z(n19199) );
  XNOR U19059 ( .A(p_input[1576]), .B(n19198), .Z(n19201) );
  XNOR U19060 ( .A(n19198), .B(n18910), .Z(n19200) );
  IV U19061 ( .A(p_input[1544]), .Z(n18910) );
  XOR U19062 ( .A(n19202), .B(n19203), .Z(n19198) );
  AND U19063 ( .A(n19204), .B(n19205), .Z(n19203) );
  XNOR U19064 ( .A(p_input[1575]), .B(n19202), .Z(n19205) );
  XNOR U19065 ( .A(n19202), .B(n18919), .Z(n19204) );
  IV U19066 ( .A(p_input[1543]), .Z(n18919) );
  XOR U19067 ( .A(n19206), .B(n19207), .Z(n19202) );
  AND U19068 ( .A(n19208), .B(n19209), .Z(n19207) );
  XNOR U19069 ( .A(p_input[1574]), .B(n19206), .Z(n19209) );
  XNOR U19070 ( .A(n19206), .B(n18928), .Z(n19208) );
  IV U19071 ( .A(p_input[1542]), .Z(n18928) );
  XOR U19072 ( .A(n19210), .B(n19211), .Z(n19206) );
  AND U19073 ( .A(n19212), .B(n19213), .Z(n19211) );
  XNOR U19074 ( .A(p_input[1573]), .B(n19210), .Z(n19213) );
  XNOR U19075 ( .A(n19210), .B(n18937), .Z(n19212) );
  IV U19076 ( .A(p_input[1541]), .Z(n18937) );
  XOR U19077 ( .A(n19214), .B(n19215), .Z(n19210) );
  AND U19078 ( .A(n19216), .B(n19217), .Z(n19215) );
  XNOR U19079 ( .A(p_input[1572]), .B(n19214), .Z(n19217) );
  XNOR U19080 ( .A(n19214), .B(n18946), .Z(n19216) );
  IV U19081 ( .A(p_input[1540]), .Z(n18946) );
  XOR U19082 ( .A(n19218), .B(n19219), .Z(n19214) );
  AND U19083 ( .A(n19220), .B(n19221), .Z(n19219) );
  XNOR U19084 ( .A(p_input[1571]), .B(n19218), .Z(n19221) );
  XNOR U19085 ( .A(n19218), .B(n18955), .Z(n19220) );
  IV U19086 ( .A(p_input[1539]), .Z(n18955) );
  XOR U19087 ( .A(n19222), .B(n19223), .Z(n19218) );
  AND U19088 ( .A(n19224), .B(n19225), .Z(n19223) );
  XNOR U19089 ( .A(p_input[1570]), .B(n19222), .Z(n19225) );
  XNOR U19090 ( .A(n19222), .B(n18964), .Z(n19224) );
  IV U19091 ( .A(p_input[1538]), .Z(n18964) );
  XNOR U19092 ( .A(n19226), .B(n19227), .Z(n19222) );
  AND U19093 ( .A(n19228), .B(n19229), .Z(n19227) );
  XOR U19094 ( .A(p_input[1569]), .B(n19226), .Z(n19229) );
  XNOR U19095 ( .A(p_input[1537]), .B(n19226), .Z(n19228) );
  AND U19096 ( .A(p_input[1568]), .B(n19230), .Z(n19226) );
  IV U19097 ( .A(p_input[1536]), .Z(n19230) );
  XOR U19098 ( .A(n19231), .B(n19232), .Z(n15587) );
  AND U19099 ( .A(n588), .B(n19233), .Z(n19232) );
  XNOR U19100 ( .A(n19234), .B(n19231), .Z(n19233) );
  XOR U19101 ( .A(n19235), .B(n19236), .Z(n588) );
  AND U19102 ( .A(n19237), .B(n19238), .Z(n19236) );
  XOR U19103 ( .A(n19235), .B(n15602), .Z(n19238) );
  XOR U19104 ( .A(n19239), .B(n19240), .Z(n15602) );
  AND U19105 ( .A(n522), .B(n19241), .Z(n19240) );
  XOR U19106 ( .A(n19242), .B(n19239), .Z(n19241) );
  XNOR U19107 ( .A(n15599), .B(n19235), .Z(n19237) );
  XOR U19108 ( .A(n19243), .B(n19244), .Z(n15599) );
  AND U19109 ( .A(n519), .B(n19245), .Z(n19244) );
  XOR U19110 ( .A(n19246), .B(n19243), .Z(n19245) );
  XOR U19111 ( .A(n19247), .B(n19248), .Z(n19235) );
  AND U19112 ( .A(n19249), .B(n19250), .Z(n19248) );
  XOR U19113 ( .A(n19247), .B(n15614), .Z(n19250) );
  XOR U19114 ( .A(n19251), .B(n19252), .Z(n15614) );
  AND U19115 ( .A(n522), .B(n19253), .Z(n19252) );
  XOR U19116 ( .A(n19254), .B(n19251), .Z(n19253) );
  XNOR U19117 ( .A(n15611), .B(n19247), .Z(n19249) );
  XOR U19118 ( .A(n19255), .B(n19256), .Z(n15611) );
  AND U19119 ( .A(n519), .B(n19257), .Z(n19256) );
  XOR U19120 ( .A(n19258), .B(n19255), .Z(n19257) );
  XOR U19121 ( .A(n19259), .B(n19260), .Z(n19247) );
  AND U19122 ( .A(n19261), .B(n19262), .Z(n19260) );
  XOR U19123 ( .A(n19259), .B(n15626), .Z(n19262) );
  XOR U19124 ( .A(n19263), .B(n19264), .Z(n15626) );
  AND U19125 ( .A(n522), .B(n19265), .Z(n19264) );
  XOR U19126 ( .A(n19266), .B(n19263), .Z(n19265) );
  XNOR U19127 ( .A(n15623), .B(n19259), .Z(n19261) );
  XOR U19128 ( .A(n19267), .B(n19268), .Z(n15623) );
  AND U19129 ( .A(n519), .B(n19269), .Z(n19268) );
  XOR U19130 ( .A(n19270), .B(n19267), .Z(n19269) );
  XOR U19131 ( .A(n19271), .B(n19272), .Z(n19259) );
  AND U19132 ( .A(n19273), .B(n19274), .Z(n19272) );
  XOR U19133 ( .A(n19271), .B(n15638), .Z(n19274) );
  XOR U19134 ( .A(n19275), .B(n19276), .Z(n15638) );
  AND U19135 ( .A(n522), .B(n19277), .Z(n19276) );
  XOR U19136 ( .A(n19278), .B(n19275), .Z(n19277) );
  XNOR U19137 ( .A(n15635), .B(n19271), .Z(n19273) );
  XOR U19138 ( .A(n19279), .B(n19280), .Z(n15635) );
  AND U19139 ( .A(n519), .B(n19281), .Z(n19280) );
  XOR U19140 ( .A(n19282), .B(n19279), .Z(n19281) );
  XOR U19141 ( .A(n19283), .B(n19284), .Z(n19271) );
  AND U19142 ( .A(n19285), .B(n19286), .Z(n19284) );
  XOR U19143 ( .A(n19283), .B(n15650), .Z(n19286) );
  XOR U19144 ( .A(n19287), .B(n19288), .Z(n15650) );
  AND U19145 ( .A(n522), .B(n19289), .Z(n19288) );
  XOR U19146 ( .A(n19290), .B(n19287), .Z(n19289) );
  XNOR U19147 ( .A(n15647), .B(n19283), .Z(n19285) );
  XOR U19148 ( .A(n19291), .B(n19292), .Z(n15647) );
  AND U19149 ( .A(n519), .B(n19293), .Z(n19292) );
  XOR U19150 ( .A(n19294), .B(n19291), .Z(n19293) );
  XOR U19151 ( .A(n19295), .B(n19296), .Z(n19283) );
  AND U19152 ( .A(n19297), .B(n19298), .Z(n19296) );
  XOR U19153 ( .A(n19295), .B(n15662), .Z(n19298) );
  XOR U19154 ( .A(n19299), .B(n19300), .Z(n15662) );
  AND U19155 ( .A(n522), .B(n19301), .Z(n19300) );
  XOR U19156 ( .A(n19302), .B(n19299), .Z(n19301) );
  XNOR U19157 ( .A(n15659), .B(n19295), .Z(n19297) );
  XOR U19158 ( .A(n19303), .B(n19304), .Z(n15659) );
  AND U19159 ( .A(n519), .B(n19305), .Z(n19304) );
  XOR U19160 ( .A(n19306), .B(n19303), .Z(n19305) );
  XOR U19161 ( .A(n19307), .B(n19308), .Z(n19295) );
  AND U19162 ( .A(n19309), .B(n19310), .Z(n19308) );
  XOR U19163 ( .A(n19307), .B(n15674), .Z(n19310) );
  XOR U19164 ( .A(n19311), .B(n19312), .Z(n15674) );
  AND U19165 ( .A(n522), .B(n19313), .Z(n19312) );
  XOR U19166 ( .A(n19314), .B(n19311), .Z(n19313) );
  XNOR U19167 ( .A(n15671), .B(n19307), .Z(n19309) );
  XOR U19168 ( .A(n19315), .B(n19316), .Z(n15671) );
  AND U19169 ( .A(n519), .B(n19317), .Z(n19316) );
  XOR U19170 ( .A(n19318), .B(n19315), .Z(n19317) );
  XOR U19171 ( .A(n19319), .B(n19320), .Z(n19307) );
  AND U19172 ( .A(n19321), .B(n19322), .Z(n19320) );
  XOR U19173 ( .A(n19319), .B(n15686), .Z(n19322) );
  XOR U19174 ( .A(n19323), .B(n19324), .Z(n15686) );
  AND U19175 ( .A(n522), .B(n19325), .Z(n19324) );
  XOR U19176 ( .A(n19326), .B(n19323), .Z(n19325) );
  XNOR U19177 ( .A(n15683), .B(n19319), .Z(n19321) );
  XOR U19178 ( .A(n19327), .B(n19328), .Z(n15683) );
  AND U19179 ( .A(n519), .B(n19329), .Z(n19328) );
  XOR U19180 ( .A(n19330), .B(n19327), .Z(n19329) );
  XOR U19181 ( .A(n19331), .B(n19332), .Z(n19319) );
  AND U19182 ( .A(n19333), .B(n19334), .Z(n19332) );
  XOR U19183 ( .A(n19331), .B(n15698), .Z(n19334) );
  XOR U19184 ( .A(n19335), .B(n19336), .Z(n15698) );
  AND U19185 ( .A(n522), .B(n19337), .Z(n19336) );
  XOR U19186 ( .A(n19338), .B(n19335), .Z(n19337) );
  XNOR U19187 ( .A(n15695), .B(n19331), .Z(n19333) );
  XOR U19188 ( .A(n19339), .B(n19340), .Z(n15695) );
  AND U19189 ( .A(n519), .B(n19341), .Z(n19340) );
  XOR U19190 ( .A(n19342), .B(n19339), .Z(n19341) );
  XOR U19191 ( .A(n19343), .B(n19344), .Z(n19331) );
  AND U19192 ( .A(n19345), .B(n19346), .Z(n19344) );
  XOR U19193 ( .A(n19343), .B(n15710), .Z(n19346) );
  XOR U19194 ( .A(n19347), .B(n19348), .Z(n15710) );
  AND U19195 ( .A(n522), .B(n19349), .Z(n19348) );
  XOR U19196 ( .A(n19350), .B(n19347), .Z(n19349) );
  XNOR U19197 ( .A(n15707), .B(n19343), .Z(n19345) );
  XOR U19198 ( .A(n19351), .B(n19352), .Z(n15707) );
  AND U19199 ( .A(n519), .B(n19353), .Z(n19352) );
  XOR U19200 ( .A(n19354), .B(n19351), .Z(n19353) );
  XOR U19201 ( .A(n19355), .B(n19356), .Z(n19343) );
  AND U19202 ( .A(n19357), .B(n19358), .Z(n19356) );
  XOR U19203 ( .A(n19355), .B(n15722), .Z(n19358) );
  XOR U19204 ( .A(n19359), .B(n19360), .Z(n15722) );
  AND U19205 ( .A(n522), .B(n19361), .Z(n19360) );
  XOR U19206 ( .A(n19362), .B(n19359), .Z(n19361) );
  XNOR U19207 ( .A(n15719), .B(n19355), .Z(n19357) );
  XOR U19208 ( .A(n19363), .B(n19364), .Z(n15719) );
  AND U19209 ( .A(n519), .B(n19365), .Z(n19364) );
  XOR U19210 ( .A(n19366), .B(n19363), .Z(n19365) );
  XOR U19211 ( .A(n19367), .B(n19368), .Z(n19355) );
  AND U19212 ( .A(n19369), .B(n19370), .Z(n19368) );
  XOR U19213 ( .A(n19367), .B(n15734), .Z(n19370) );
  XOR U19214 ( .A(n19371), .B(n19372), .Z(n15734) );
  AND U19215 ( .A(n522), .B(n19373), .Z(n19372) );
  XOR U19216 ( .A(n19374), .B(n19371), .Z(n19373) );
  XNOR U19217 ( .A(n15731), .B(n19367), .Z(n19369) );
  XOR U19218 ( .A(n19375), .B(n19376), .Z(n15731) );
  AND U19219 ( .A(n519), .B(n19377), .Z(n19376) );
  XOR U19220 ( .A(n19378), .B(n19375), .Z(n19377) );
  XOR U19221 ( .A(n19379), .B(n19380), .Z(n19367) );
  AND U19222 ( .A(n19381), .B(n19382), .Z(n19380) );
  XOR U19223 ( .A(n19379), .B(n15746), .Z(n19382) );
  XOR U19224 ( .A(n19383), .B(n19384), .Z(n15746) );
  AND U19225 ( .A(n522), .B(n19385), .Z(n19384) );
  XOR U19226 ( .A(n19386), .B(n19383), .Z(n19385) );
  XNOR U19227 ( .A(n15743), .B(n19379), .Z(n19381) );
  XOR U19228 ( .A(n19387), .B(n19388), .Z(n15743) );
  AND U19229 ( .A(n519), .B(n19389), .Z(n19388) );
  XOR U19230 ( .A(n19390), .B(n19387), .Z(n19389) );
  XOR U19231 ( .A(n19391), .B(n19392), .Z(n19379) );
  AND U19232 ( .A(n19393), .B(n19394), .Z(n19392) );
  XOR U19233 ( .A(n19391), .B(n15758), .Z(n19394) );
  XOR U19234 ( .A(n19395), .B(n19396), .Z(n15758) );
  AND U19235 ( .A(n522), .B(n19397), .Z(n19396) );
  XOR U19236 ( .A(n19398), .B(n19395), .Z(n19397) );
  XNOR U19237 ( .A(n15755), .B(n19391), .Z(n19393) );
  XOR U19238 ( .A(n19399), .B(n19400), .Z(n15755) );
  AND U19239 ( .A(n519), .B(n19401), .Z(n19400) );
  XOR U19240 ( .A(n19402), .B(n19399), .Z(n19401) );
  XOR U19241 ( .A(n19403), .B(n19404), .Z(n19391) );
  AND U19242 ( .A(n19405), .B(n19406), .Z(n19404) );
  XOR U19243 ( .A(n19403), .B(n15770), .Z(n19406) );
  XOR U19244 ( .A(n19407), .B(n19408), .Z(n15770) );
  AND U19245 ( .A(n522), .B(n19409), .Z(n19408) );
  XOR U19246 ( .A(n19410), .B(n19407), .Z(n19409) );
  XNOR U19247 ( .A(n15767), .B(n19403), .Z(n19405) );
  XOR U19248 ( .A(n19411), .B(n19412), .Z(n15767) );
  AND U19249 ( .A(n519), .B(n19413), .Z(n19412) );
  XOR U19250 ( .A(n19414), .B(n19411), .Z(n19413) );
  XOR U19251 ( .A(n19415), .B(n19416), .Z(n19403) );
  AND U19252 ( .A(n19417), .B(n19418), .Z(n19416) );
  XOR U19253 ( .A(n19415), .B(n15782), .Z(n19418) );
  XOR U19254 ( .A(n19419), .B(n19420), .Z(n15782) );
  AND U19255 ( .A(n522), .B(n19421), .Z(n19420) );
  XOR U19256 ( .A(n19422), .B(n19419), .Z(n19421) );
  XNOR U19257 ( .A(n15779), .B(n19415), .Z(n19417) );
  XOR U19258 ( .A(n19423), .B(n19424), .Z(n15779) );
  AND U19259 ( .A(n519), .B(n19425), .Z(n19424) );
  XOR U19260 ( .A(n19426), .B(n19423), .Z(n19425) );
  XOR U19261 ( .A(n19427), .B(n19428), .Z(n19415) );
  AND U19262 ( .A(n19429), .B(n19430), .Z(n19428) );
  XOR U19263 ( .A(n19427), .B(n15794), .Z(n19430) );
  XOR U19264 ( .A(n19431), .B(n19432), .Z(n15794) );
  AND U19265 ( .A(n522), .B(n19433), .Z(n19432) );
  XOR U19266 ( .A(n19434), .B(n19431), .Z(n19433) );
  XNOR U19267 ( .A(n15791), .B(n19427), .Z(n19429) );
  XOR U19268 ( .A(n19435), .B(n19436), .Z(n15791) );
  AND U19269 ( .A(n519), .B(n19437), .Z(n19436) );
  XOR U19270 ( .A(n19438), .B(n19435), .Z(n19437) );
  XOR U19271 ( .A(n19439), .B(n19440), .Z(n19427) );
  AND U19272 ( .A(n19441), .B(n19442), .Z(n19440) );
  XOR U19273 ( .A(n19439), .B(n15806), .Z(n19442) );
  XOR U19274 ( .A(n19443), .B(n19444), .Z(n15806) );
  AND U19275 ( .A(n522), .B(n19445), .Z(n19444) );
  XOR U19276 ( .A(n19446), .B(n19443), .Z(n19445) );
  XNOR U19277 ( .A(n15803), .B(n19439), .Z(n19441) );
  XOR U19278 ( .A(n19447), .B(n19448), .Z(n15803) );
  AND U19279 ( .A(n519), .B(n19449), .Z(n19448) );
  XOR U19280 ( .A(n19450), .B(n19447), .Z(n19449) );
  XOR U19281 ( .A(n19451), .B(n19452), .Z(n19439) );
  AND U19282 ( .A(n19453), .B(n19454), .Z(n19452) );
  XOR U19283 ( .A(n19451), .B(n15818), .Z(n19454) );
  XOR U19284 ( .A(n19455), .B(n19456), .Z(n15818) );
  AND U19285 ( .A(n522), .B(n19457), .Z(n19456) );
  XOR U19286 ( .A(n19458), .B(n19455), .Z(n19457) );
  XNOR U19287 ( .A(n15815), .B(n19451), .Z(n19453) );
  XOR U19288 ( .A(n19459), .B(n19460), .Z(n15815) );
  AND U19289 ( .A(n519), .B(n19461), .Z(n19460) );
  XOR U19290 ( .A(n19462), .B(n19459), .Z(n19461) );
  XOR U19291 ( .A(n19463), .B(n19464), .Z(n19451) );
  AND U19292 ( .A(n19465), .B(n19466), .Z(n19464) );
  XOR U19293 ( .A(n19463), .B(n15830), .Z(n19466) );
  XOR U19294 ( .A(n19467), .B(n19468), .Z(n15830) );
  AND U19295 ( .A(n522), .B(n19469), .Z(n19468) );
  XOR U19296 ( .A(n19470), .B(n19467), .Z(n19469) );
  XNOR U19297 ( .A(n15827), .B(n19463), .Z(n19465) );
  XOR U19298 ( .A(n19471), .B(n19472), .Z(n15827) );
  AND U19299 ( .A(n519), .B(n19473), .Z(n19472) );
  XOR U19300 ( .A(n19474), .B(n19471), .Z(n19473) );
  XOR U19301 ( .A(n19475), .B(n19476), .Z(n19463) );
  AND U19302 ( .A(n19477), .B(n19478), .Z(n19476) );
  XOR U19303 ( .A(n19475), .B(n15842), .Z(n19478) );
  XOR U19304 ( .A(n19479), .B(n19480), .Z(n15842) );
  AND U19305 ( .A(n522), .B(n19481), .Z(n19480) );
  XOR U19306 ( .A(n19482), .B(n19479), .Z(n19481) );
  XNOR U19307 ( .A(n15839), .B(n19475), .Z(n19477) );
  XOR U19308 ( .A(n19483), .B(n19484), .Z(n15839) );
  AND U19309 ( .A(n519), .B(n19485), .Z(n19484) );
  XOR U19310 ( .A(n19486), .B(n19483), .Z(n19485) );
  XOR U19311 ( .A(n19487), .B(n19488), .Z(n19475) );
  AND U19312 ( .A(n19489), .B(n19490), .Z(n19488) );
  XOR U19313 ( .A(n19487), .B(n15854), .Z(n19490) );
  XOR U19314 ( .A(n19491), .B(n19492), .Z(n15854) );
  AND U19315 ( .A(n522), .B(n19493), .Z(n19492) );
  XOR U19316 ( .A(n19494), .B(n19491), .Z(n19493) );
  XNOR U19317 ( .A(n15851), .B(n19487), .Z(n19489) );
  XOR U19318 ( .A(n19495), .B(n19496), .Z(n15851) );
  AND U19319 ( .A(n519), .B(n19497), .Z(n19496) );
  XOR U19320 ( .A(n19498), .B(n19495), .Z(n19497) );
  XOR U19321 ( .A(n19499), .B(n19500), .Z(n19487) );
  AND U19322 ( .A(n19501), .B(n19502), .Z(n19500) );
  XOR U19323 ( .A(n19499), .B(n15866), .Z(n19502) );
  XOR U19324 ( .A(n19503), .B(n19504), .Z(n15866) );
  AND U19325 ( .A(n522), .B(n19505), .Z(n19504) );
  XOR U19326 ( .A(n19506), .B(n19503), .Z(n19505) );
  XNOR U19327 ( .A(n15863), .B(n19499), .Z(n19501) );
  XOR U19328 ( .A(n19507), .B(n19508), .Z(n15863) );
  AND U19329 ( .A(n519), .B(n19509), .Z(n19508) );
  XOR U19330 ( .A(n19510), .B(n19507), .Z(n19509) );
  XOR U19331 ( .A(n19511), .B(n19512), .Z(n19499) );
  AND U19332 ( .A(n19513), .B(n19514), .Z(n19512) );
  XOR U19333 ( .A(n19511), .B(n15878), .Z(n19514) );
  XOR U19334 ( .A(n19515), .B(n19516), .Z(n15878) );
  AND U19335 ( .A(n522), .B(n19517), .Z(n19516) );
  XOR U19336 ( .A(n19518), .B(n19515), .Z(n19517) );
  XNOR U19337 ( .A(n15875), .B(n19511), .Z(n19513) );
  XOR U19338 ( .A(n19519), .B(n19520), .Z(n15875) );
  AND U19339 ( .A(n519), .B(n19521), .Z(n19520) );
  XOR U19340 ( .A(n19522), .B(n19519), .Z(n19521) );
  XOR U19341 ( .A(n19523), .B(n19524), .Z(n19511) );
  AND U19342 ( .A(n19525), .B(n19526), .Z(n19524) );
  XOR U19343 ( .A(n19523), .B(n15890), .Z(n19526) );
  XOR U19344 ( .A(n19527), .B(n19528), .Z(n15890) );
  AND U19345 ( .A(n522), .B(n19529), .Z(n19528) );
  XOR U19346 ( .A(n19530), .B(n19527), .Z(n19529) );
  XNOR U19347 ( .A(n15887), .B(n19523), .Z(n19525) );
  XOR U19348 ( .A(n19531), .B(n19532), .Z(n15887) );
  AND U19349 ( .A(n519), .B(n19533), .Z(n19532) );
  XOR U19350 ( .A(n19534), .B(n19531), .Z(n19533) );
  XOR U19351 ( .A(n19535), .B(n19536), .Z(n19523) );
  AND U19352 ( .A(n19537), .B(n19538), .Z(n19536) );
  XOR U19353 ( .A(n19535), .B(n15902), .Z(n19538) );
  XOR U19354 ( .A(n19539), .B(n19540), .Z(n15902) );
  AND U19355 ( .A(n522), .B(n19541), .Z(n19540) );
  XOR U19356 ( .A(n19542), .B(n19539), .Z(n19541) );
  XNOR U19357 ( .A(n15899), .B(n19535), .Z(n19537) );
  XOR U19358 ( .A(n19543), .B(n19544), .Z(n15899) );
  AND U19359 ( .A(n519), .B(n19545), .Z(n19544) );
  XOR U19360 ( .A(n19546), .B(n19543), .Z(n19545) );
  XOR U19361 ( .A(n19547), .B(n19548), .Z(n19535) );
  AND U19362 ( .A(n19549), .B(n19550), .Z(n19548) );
  XOR U19363 ( .A(n19547), .B(n15914), .Z(n19550) );
  XOR U19364 ( .A(n19551), .B(n19552), .Z(n15914) );
  AND U19365 ( .A(n522), .B(n19553), .Z(n19552) );
  XOR U19366 ( .A(n19554), .B(n19551), .Z(n19553) );
  XNOR U19367 ( .A(n15911), .B(n19547), .Z(n19549) );
  XOR U19368 ( .A(n19555), .B(n19556), .Z(n15911) );
  AND U19369 ( .A(n519), .B(n19557), .Z(n19556) );
  XOR U19370 ( .A(n19558), .B(n19555), .Z(n19557) );
  XOR U19371 ( .A(n19559), .B(n19560), .Z(n19547) );
  AND U19372 ( .A(n19561), .B(n19562), .Z(n19560) );
  XOR U19373 ( .A(n19559), .B(n15926), .Z(n19562) );
  XOR U19374 ( .A(n19563), .B(n19564), .Z(n15926) );
  AND U19375 ( .A(n522), .B(n19565), .Z(n19564) );
  XOR U19376 ( .A(n19566), .B(n19563), .Z(n19565) );
  XNOR U19377 ( .A(n15923), .B(n19559), .Z(n19561) );
  XOR U19378 ( .A(n19567), .B(n19568), .Z(n15923) );
  AND U19379 ( .A(n519), .B(n19569), .Z(n19568) );
  XOR U19380 ( .A(n19570), .B(n19567), .Z(n19569) );
  XOR U19381 ( .A(n19571), .B(n19572), .Z(n19559) );
  AND U19382 ( .A(n19573), .B(n19574), .Z(n19572) );
  XOR U19383 ( .A(n19571), .B(n15938), .Z(n19574) );
  XOR U19384 ( .A(n19575), .B(n19576), .Z(n15938) );
  AND U19385 ( .A(n522), .B(n19577), .Z(n19576) );
  XOR U19386 ( .A(n19578), .B(n19575), .Z(n19577) );
  XNOR U19387 ( .A(n15935), .B(n19571), .Z(n19573) );
  XOR U19388 ( .A(n19579), .B(n19580), .Z(n15935) );
  AND U19389 ( .A(n519), .B(n19581), .Z(n19580) );
  XOR U19390 ( .A(n19582), .B(n19579), .Z(n19581) );
  XOR U19391 ( .A(n19583), .B(n19584), .Z(n19571) );
  AND U19392 ( .A(n19585), .B(n19586), .Z(n19584) );
  XOR U19393 ( .A(n15950), .B(n19583), .Z(n19586) );
  XOR U19394 ( .A(n19587), .B(n19588), .Z(n15950) );
  AND U19395 ( .A(n522), .B(n19589), .Z(n19588) );
  XOR U19396 ( .A(n19587), .B(n19590), .Z(n19589) );
  XNOR U19397 ( .A(n19583), .B(n15947), .Z(n19585) );
  XOR U19398 ( .A(n19591), .B(n19592), .Z(n15947) );
  AND U19399 ( .A(n519), .B(n19593), .Z(n19592) );
  XOR U19400 ( .A(n19591), .B(n19594), .Z(n19593) );
  XOR U19401 ( .A(n19595), .B(n19596), .Z(n19583) );
  AND U19402 ( .A(n19597), .B(n19598), .Z(n19596) );
  XNOR U19403 ( .A(n19599), .B(n15963), .Z(n19598) );
  XOR U19404 ( .A(n19600), .B(n19601), .Z(n15963) );
  AND U19405 ( .A(n522), .B(n19602), .Z(n19601) );
  XOR U19406 ( .A(n19603), .B(n19600), .Z(n19602) );
  XNOR U19407 ( .A(n15960), .B(n19595), .Z(n19597) );
  XOR U19408 ( .A(n19604), .B(n19605), .Z(n15960) );
  AND U19409 ( .A(n519), .B(n19606), .Z(n19605) );
  XOR U19410 ( .A(n19607), .B(n19604), .Z(n19606) );
  IV U19411 ( .A(n19599), .Z(n19595) );
  AND U19412 ( .A(n19231), .B(n19234), .Z(n19599) );
  XNOR U19413 ( .A(n19608), .B(n19609), .Z(n19234) );
  AND U19414 ( .A(n522), .B(n19610), .Z(n19609) );
  XNOR U19415 ( .A(n19611), .B(n19608), .Z(n19610) );
  XOR U19416 ( .A(n19612), .B(n19613), .Z(n522) );
  AND U19417 ( .A(n19614), .B(n19615), .Z(n19613) );
  XOR U19418 ( .A(n19612), .B(n19242), .Z(n19615) );
  XNOR U19419 ( .A(n19616), .B(n19617), .Z(n19242) );
  AND U19420 ( .A(n19618), .B(n378), .Z(n19617) );
  AND U19421 ( .A(n19616), .B(n19619), .Z(n19618) );
  XNOR U19422 ( .A(n19239), .B(n19612), .Z(n19614) );
  XOR U19423 ( .A(n19620), .B(n19621), .Z(n19239) );
  AND U19424 ( .A(n19622), .B(n376), .Z(n19621) );
  NOR U19425 ( .A(n19620), .B(n19623), .Z(n19622) );
  XOR U19426 ( .A(n19624), .B(n19625), .Z(n19612) );
  AND U19427 ( .A(n19626), .B(n19627), .Z(n19625) );
  XOR U19428 ( .A(n19624), .B(n19254), .Z(n19627) );
  XOR U19429 ( .A(n19628), .B(n19629), .Z(n19254) );
  AND U19430 ( .A(n378), .B(n19630), .Z(n19629) );
  XOR U19431 ( .A(n19631), .B(n19628), .Z(n19630) );
  XNOR U19432 ( .A(n19251), .B(n19624), .Z(n19626) );
  XOR U19433 ( .A(n19632), .B(n19633), .Z(n19251) );
  AND U19434 ( .A(n376), .B(n19634), .Z(n19633) );
  XOR U19435 ( .A(n19635), .B(n19632), .Z(n19634) );
  XOR U19436 ( .A(n19636), .B(n19637), .Z(n19624) );
  AND U19437 ( .A(n19638), .B(n19639), .Z(n19637) );
  XOR U19438 ( .A(n19636), .B(n19266), .Z(n19639) );
  XOR U19439 ( .A(n19640), .B(n19641), .Z(n19266) );
  AND U19440 ( .A(n378), .B(n19642), .Z(n19641) );
  XOR U19441 ( .A(n19643), .B(n19640), .Z(n19642) );
  XNOR U19442 ( .A(n19263), .B(n19636), .Z(n19638) );
  XOR U19443 ( .A(n19644), .B(n19645), .Z(n19263) );
  AND U19444 ( .A(n376), .B(n19646), .Z(n19645) );
  XOR U19445 ( .A(n19647), .B(n19644), .Z(n19646) );
  XOR U19446 ( .A(n19648), .B(n19649), .Z(n19636) );
  AND U19447 ( .A(n19650), .B(n19651), .Z(n19649) );
  XOR U19448 ( .A(n19648), .B(n19278), .Z(n19651) );
  XOR U19449 ( .A(n19652), .B(n19653), .Z(n19278) );
  AND U19450 ( .A(n378), .B(n19654), .Z(n19653) );
  XOR U19451 ( .A(n19655), .B(n19652), .Z(n19654) );
  XNOR U19452 ( .A(n19275), .B(n19648), .Z(n19650) );
  XOR U19453 ( .A(n19656), .B(n19657), .Z(n19275) );
  AND U19454 ( .A(n376), .B(n19658), .Z(n19657) );
  XOR U19455 ( .A(n19659), .B(n19656), .Z(n19658) );
  XOR U19456 ( .A(n19660), .B(n19661), .Z(n19648) );
  AND U19457 ( .A(n19662), .B(n19663), .Z(n19661) );
  XOR U19458 ( .A(n19660), .B(n19290), .Z(n19663) );
  XOR U19459 ( .A(n19664), .B(n19665), .Z(n19290) );
  AND U19460 ( .A(n378), .B(n19666), .Z(n19665) );
  XOR U19461 ( .A(n19667), .B(n19664), .Z(n19666) );
  XNOR U19462 ( .A(n19287), .B(n19660), .Z(n19662) );
  XOR U19463 ( .A(n19668), .B(n19669), .Z(n19287) );
  AND U19464 ( .A(n376), .B(n19670), .Z(n19669) );
  XOR U19465 ( .A(n19671), .B(n19668), .Z(n19670) );
  XOR U19466 ( .A(n19672), .B(n19673), .Z(n19660) );
  AND U19467 ( .A(n19674), .B(n19675), .Z(n19673) );
  XOR U19468 ( .A(n19672), .B(n19302), .Z(n19675) );
  XOR U19469 ( .A(n19676), .B(n19677), .Z(n19302) );
  AND U19470 ( .A(n378), .B(n19678), .Z(n19677) );
  XOR U19471 ( .A(n19679), .B(n19676), .Z(n19678) );
  XNOR U19472 ( .A(n19299), .B(n19672), .Z(n19674) );
  XOR U19473 ( .A(n19680), .B(n19681), .Z(n19299) );
  AND U19474 ( .A(n376), .B(n19682), .Z(n19681) );
  XOR U19475 ( .A(n19683), .B(n19680), .Z(n19682) );
  XOR U19476 ( .A(n19684), .B(n19685), .Z(n19672) );
  AND U19477 ( .A(n19686), .B(n19687), .Z(n19685) );
  XOR U19478 ( .A(n19684), .B(n19314), .Z(n19687) );
  XOR U19479 ( .A(n19688), .B(n19689), .Z(n19314) );
  AND U19480 ( .A(n378), .B(n19690), .Z(n19689) );
  XOR U19481 ( .A(n19691), .B(n19688), .Z(n19690) );
  XNOR U19482 ( .A(n19311), .B(n19684), .Z(n19686) );
  XOR U19483 ( .A(n19692), .B(n19693), .Z(n19311) );
  AND U19484 ( .A(n376), .B(n19694), .Z(n19693) );
  XOR U19485 ( .A(n19695), .B(n19692), .Z(n19694) );
  XOR U19486 ( .A(n19696), .B(n19697), .Z(n19684) );
  AND U19487 ( .A(n19698), .B(n19699), .Z(n19697) );
  XOR U19488 ( .A(n19696), .B(n19326), .Z(n19699) );
  XOR U19489 ( .A(n19700), .B(n19701), .Z(n19326) );
  AND U19490 ( .A(n378), .B(n19702), .Z(n19701) );
  XOR U19491 ( .A(n19703), .B(n19700), .Z(n19702) );
  XNOR U19492 ( .A(n19323), .B(n19696), .Z(n19698) );
  XOR U19493 ( .A(n19704), .B(n19705), .Z(n19323) );
  AND U19494 ( .A(n376), .B(n19706), .Z(n19705) );
  XOR U19495 ( .A(n19707), .B(n19704), .Z(n19706) );
  XOR U19496 ( .A(n19708), .B(n19709), .Z(n19696) );
  AND U19497 ( .A(n19710), .B(n19711), .Z(n19709) );
  XOR U19498 ( .A(n19708), .B(n19338), .Z(n19711) );
  XOR U19499 ( .A(n19712), .B(n19713), .Z(n19338) );
  AND U19500 ( .A(n378), .B(n19714), .Z(n19713) );
  XOR U19501 ( .A(n19715), .B(n19712), .Z(n19714) );
  XNOR U19502 ( .A(n19335), .B(n19708), .Z(n19710) );
  XOR U19503 ( .A(n19716), .B(n19717), .Z(n19335) );
  AND U19504 ( .A(n376), .B(n19718), .Z(n19717) );
  XOR U19505 ( .A(n19719), .B(n19716), .Z(n19718) );
  XOR U19506 ( .A(n19720), .B(n19721), .Z(n19708) );
  AND U19507 ( .A(n19722), .B(n19723), .Z(n19721) );
  XOR U19508 ( .A(n19720), .B(n19350), .Z(n19723) );
  XOR U19509 ( .A(n19724), .B(n19725), .Z(n19350) );
  AND U19510 ( .A(n378), .B(n19726), .Z(n19725) );
  XOR U19511 ( .A(n19727), .B(n19724), .Z(n19726) );
  XNOR U19512 ( .A(n19347), .B(n19720), .Z(n19722) );
  XOR U19513 ( .A(n19728), .B(n19729), .Z(n19347) );
  AND U19514 ( .A(n376), .B(n19730), .Z(n19729) );
  XOR U19515 ( .A(n19731), .B(n19728), .Z(n19730) );
  XOR U19516 ( .A(n19732), .B(n19733), .Z(n19720) );
  AND U19517 ( .A(n19734), .B(n19735), .Z(n19733) );
  XOR U19518 ( .A(n19732), .B(n19362), .Z(n19735) );
  XOR U19519 ( .A(n19736), .B(n19737), .Z(n19362) );
  AND U19520 ( .A(n378), .B(n19738), .Z(n19737) );
  XOR U19521 ( .A(n19739), .B(n19736), .Z(n19738) );
  XNOR U19522 ( .A(n19359), .B(n19732), .Z(n19734) );
  XOR U19523 ( .A(n19740), .B(n19741), .Z(n19359) );
  AND U19524 ( .A(n376), .B(n19742), .Z(n19741) );
  XOR U19525 ( .A(n19743), .B(n19740), .Z(n19742) );
  XOR U19526 ( .A(n19744), .B(n19745), .Z(n19732) );
  AND U19527 ( .A(n19746), .B(n19747), .Z(n19745) );
  XOR U19528 ( .A(n19744), .B(n19374), .Z(n19747) );
  XOR U19529 ( .A(n19748), .B(n19749), .Z(n19374) );
  AND U19530 ( .A(n378), .B(n19750), .Z(n19749) );
  XOR U19531 ( .A(n19751), .B(n19748), .Z(n19750) );
  XNOR U19532 ( .A(n19371), .B(n19744), .Z(n19746) );
  XOR U19533 ( .A(n19752), .B(n19753), .Z(n19371) );
  AND U19534 ( .A(n376), .B(n19754), .Z(n19753) );
  XOR U19535 ( .A(n19755), .B(n19752), .Z(n19754) );
  XOR U19536 ( .A(n19756), .B(n19757), .Z(n19744) );
  AND U19537 ( .A(n19758), .B(n19759), .Z(n19757) );
  XOR U19538 ( .A(n19756), .B(n19386), .Z(n19759) );
  XOR U19539 ( .A(n19760), .B(n19761), .Z(n19386) );
  AND U19540 ( .A(n378), .B(n19762), .Z(n19761) );
  XOR U19541 ( .A(n19763), .B(n19760), .Z(n19762) );
  XNOR U19542 ( .A(n19383), .B(n19756), .Z(n19758) );
  XOR U19543 ( .A(n19764), .B(n19765), .Z(n19383) );
  AND U19544 ( .A(n376), .B(n19766), .Z(n19765) );
  XOR U19545 ( .A(n19767), .B(n19764), .Z(n19766) );
  XOR U19546 ( .A(n19768), .B(n19769), .Z(n19756) );
  AND U19547 ( .A(n19770), .B(n19771), .Z(n19769) );
  XOR U19548 ( .A(n19768), .B(n19398), .Z(n19771) );
  XOR U19549 ( .A(n19772), .B(n19773), .Z(n19398) );
  AND U19550 ( .A(n378), .B(n19774), .Z(n19773) );
  XOR U19551 ( .A(n19775), .B(n19772), .Z(n19774) );
  XNOR U19552 ( .A(n19395), .B(n19768), .Z(n19770) );
  XOR U19553 ( .A(n19776), .B(n19777), .Z(n19395) );
  AND U19554 ( .A(n376), .B(n19778), .Z(n19777) );
  XOR U19555 ( .A(n19779), .B(n19776), .Z(n19778) );
  XOR U19556 ( .A(n19780), .B(n19781), .Z(n19768) );
  AND U19557 ( .A(n19782), .B(n19783), .Z(n19781) );
  XOR U19558 ( .A(n19780), .B(n19410), .Z(n19783) );
  XOR U19559 ( .A(n19784), .B(n19785), .Z(n19410) );
  AND U19560 ( .A(n378), .B(n19786), .Z(n19785) );
  XOR U19561 ( .A(n19787), .B(n19784), .Z(n19786) );
  XNOR U19562 ( .A(n19407), .B(n19780), .Z(n19782) );
  XOR U19563 ( .A(n19788), .B(n19789), .Z(n19407) );
  AND U19564 ( .A(n376), .B(n19790), .Z(n19789) );
  XOR U19565 ( .A(n19791), .B(n19788), .Z(n19790) );
  XOR U19566 ( .A(n19792), .B(n19793), .Z(n19780) );
  AND U19567 ( .A(n19794), .B(n19795), .Z(n19793) );
  XOR U19568 ( .A(n19792), .B(n19422), .Z(n19795) );
  XOR U19569 ( .A(n19796), .B(n19797), .Z(n19422) );
  AND U19570 ( .A(n378), .B(n19798), .Z(n19797) );
  XOR U19571 ( .A(n19799), .B(n19796), .Z(n19798) );
  XNOR U19572 ( .A(n19419), .B(n19792), .Z(n19794) );
  XOR U19573 ( .A(n19800), .B(n19801), .Z(n19419) );
  AND U19574 ( .A(n376), .B(n19802), .Z(n19801) );
  XOR U19575 ( .A(n19803), .B(n19800), .Z(n19802) );
  XOR U19576 ( .A(n19804), .B(n19805), .Z(n19792) );
  AND U19577 ( .A(n19806), .B(n19807), .Z(n19805) );
  XOR U19578 ( .A(n19804), .B(n19434), .Z(n19807) );
  XOR U19579 ( .A(n19808), .B(n19809), .Z(n19434) );
  AND U19580 ( .A(n378), .B(n19810), .Z(n19809) );
  XOR U19581 ( .A(n19811), .B(n19808), .Z(n19810) );
  XNOR U19582 ( .A(n19431), .B(n19804), .Z(n19806) );
  XOR U19583 ( .A(n19812), .B(n19813), .Z(n19431) );
  AND U19584 ( .A(n376), .B(n19814), .Z(n19813) );
  XOR U19585 ( .A(n19815), .B(n19812), .Z(n19814) );
  XOR U19586 ( .A(n19816), .B(n19817), .Z(n19804) );
  AND U19587 ( .A(n19818), .B(n19819), .Z(n19817) );
  XOR U19588 ( .A(n19816), .B(n19446), .Z(n19819) );
  XOR U19589 ( .A(n19820), .B(n19821), .Z(n19446) );
  AND U19590 ( .A(n378), .B(n19822), .Z(n19821) );
  XOR U19591 ( .A(n19823), .B(n19820), .Z(n19822) );
  XNOR U19592 ( .A(n19443), .B(n19816), .Z(n19818) );
  XOR U19593 ( .A(n19824), .B(n19825), .Z(n19443) );
  AND U19594 ( .A(n376), .B(n19826), .Z(n19825) );
  XOR U19595 ( .A(n19827), .B(n19824), .Z(n19826) );
  XOR U19596 ( .A(n19828), .B(n19829), .Z(n19816) );
  AND U19597 ( .A(n19830), .B(n19831), .Z(n19829) );
  XOR U19598 ( .A(n19828), .B(n19458), .Z(n19831) );
  XOR U19599 ( .A(n19832), .B(n19833), .Z(n19458) );
  AND U19600 ( .A(n378), .B(n19834), .Z(n19833) );
  XOR U19601 ( .A(n19835), .B(n19832), .Z(n19834) );
  XNOR U19602 ( .A(n19455), .B(n19828), .Z(n19830) );
  XOR U19603 ( .A(n19836), .B(n19837), .Z(n19455) );
  AND U19604 ( .A(n376), .B(n19838), .Z(n19837) );
  XOR U19605 ( .A(n19839), .B(n19836), .Z(n19838) );
  XOR U19606 ( .A(n19840), .B(n19841), .Z(n19828) );
  AND U19607 ( .A(n19842), .B(n19843), .Z(n19841) );
  XOR U19608 ( .A(n19840), .B(n19470), .Z(n19843) );
  XOR U19609 ( .A(n19844), .B(n19845), .Z(n19470) );
  AND U19610 ( .A(n378), .B(n19846), .Z(n19845) );
  XOR U19611 ( .A(n19847), .B(n19844), .Z(n19846) );
  XNOR U19612 ( .A(n19467), .B(n19840), .Z(n19842) );
  XOR U19613 ( .A(n19848), .B(n19849), .Z(n19467) );
  AND U19614 ( .A(n376), .B(n19850), .Z(n19849) );
  XOR U19615 ( .A(n19851), .B(n19848), .Z(n19850) );
  XOR U19616 ( .A(n19852), .B(n19853), .Z(n19840) );
  AND U19617 ( .A(n19854), .B(n19855), .Z(n19853) );
  XOR U19618 ( .A(n19852), .B(n19482), .Z(n19855) );
  XOR U19619 ( .A(n19856), .B(n19857), .Z(n19482) );
  AND U19620 ( .A(n378), .B(n19858), .Z(n19857) );
  XOR U19621 ( .A(n19859), .B(n19856), .Z(n19858) );
  XNOR U19622 ( .A(n19479), .B(n19852), .Z(n19854) );
  XOR U19623 ( .A(n19860), .B(n19861), .Z(n19479) );
  AND U19624 ( .A(n376), .B(n19862), .Z(n19861) );
  XOR U19625 ( .A(n19863), .B(n19860), .Z(n19862) );
  XOR U19626 ( .A(n19864), .B(n19865), .Z(n19852) );
  AND U19627 ( .A(n19866), .B(n19867), .Z(n19865) );
  XOR U19628 ( .A(n19864), .B(n19494), .Z(n19867) );
  XOR U19629 ( .A(n19868), .B(n19869), .Z(n19494) );
  AND U19630 ( .A(n378), .B(n19870), .Z(n19869) );
  XOR U19631 ( .A(n19871), .B(n19868), .Z(n19870) );
  XNOR U19632 ( .A(n19491), .B(n19864), .Z(n19866) );
  XOR U19633 ( .A(n19872), .B(n19873), .Z(n19491) );
  AND U19634 ( .A(n376), .B(n19874), .Z(n19873) );
  XOR U19635 ( .A(n19875), .B(n19872), .Z(n19874) );
  XOR U19636 ( .A(n19876), .B(n19877), .Z(n19864) );
  AND U19637 ( .A(n19878), .B(n19879), .Z(n19877) );
  XOR U19638 ( .A(n19876), .B(n19506), .Z(n19879) );
  XOR U19639 ( .A(n19880), .B(n19881), .Z(n19506) );
  AND U19640 ( .A(n378), .B(n19882), .Z(n19881) );
  XOR U19641 ( .A(n19883), .B(n19880), .Z(n19882) );
  XNOR U19642 ( .A(n19503), .B(n19876), .Z(n19878) );
  XOR U19643 ( .A(n19884), .B(n19885), .Z(n19503) );
  AND U19644 ( .A(n376), .B(n19886), .Z(n19885) );
  XOR U19645 ( .A(n19887), .B(n19884), .Z(n19886) );
  XOR U19646 ( .A(n19888), .B(n19889), .Z(n19876) );
  AND U19647 ( .A(n19890), .B(n19891), .Z(n19889) );
  XOR U19648 ( .A(n19888), .B(n19518), .Z(n19891) );
  XOR U19649 ( .A(n19892), .B(n19893), .Z(n19518) );
  AND U19650 ( .A(n378), .B(n19894), .Z(n19893) );
  XOR U19651 ( .A(n19895), .B(n19892), .Z(n19894) );
  XNOR U19652 ( .A(n19515), .B(n19888), .Z(n19890) );
  XOR U19653 ( .A(n19896), .B(n19897), .Z(n19515) );
  AND U19654 ( .A(n376), .B(n19898), .Z(n19897) );
  XOR U19655 ( .A(n19899), .B(n19896), .Z(n19898) );
  XOR U19656 ( .A(n19900), .B(n19901), .Z(n19888) );
  AND U19657 ( .A(n19902), .B(n19903), .Z(n19901) );
  XOR U19658 ( .A(n19900), .B(n19530), .Z(n19903) );
  XOR U19659 ( .A(n19904), .B(n19905), .Z(n19530) );
  AND U19660 ( .A(n378), .B(n19906), .Z(n19905) );
  XOR U19661 ( .A(n19907), .B(n19904), .Z(n19906) );
  XNOR U19662 ( .A(n19527), .B(n19900), .Z(n19902) );
  XOR U19663 ( .A(n19908), .B(n19909), .Z(n19527) );
  AND U19664 ( .A(n376), .B(n19910), .Z(n19909) );
  XOR U19665 ( .A(n19911), .B(n19908), .Z(n19910) );
  XOR U19666 ( .A(n19912), .B(n19913), .Z(n19900) );
  AND U19667 ( .A(n19914), .B(n19915), .Z(n19913) );
  XOR U19668 ( .A(n19912), .B(n19542), .Z(n19915) );
  XOR U19669 ( .A(n19916), .B(n19917), .Z(n19542) );
  AND U19670 ( .A(n378), .B(n19918), .Z(n19917) );
  XOR U19671 ( .A(n19919), .B(n19916), .Z(n19918) );
  XNOR U19672 ( .A(n19539), .B(n19912), .Z(n19914) );
  XOR U19673 ( .A(n19920), .B(n19921), .Z(n19539) );
  AND U19674 ( .A(n376), .B(n19922), .Z(n19921) );
  XOR U19675 ( .A(n19923), .B(n19920), .Z(n19922) );
  XOR U19676 ( .A(n19924), .B(n19925), .Z(n19912) );
  AND U19677 ( .A(n19926), .B(n19927), .Z(n19925) );
  XOR U19678 ( .A(n19924), .B(n19554), .Z(n19927) );
  XOR U19679 ( .A(n19928), .B(n19929), .Z(n19554) );
  AND U19680 ( .A(n378), .B(n19930), .Z(n19929) );
  XOR U19681 ( .A(n19931), .B(n19928), .Z(n19930) );
  XNOR U19682 ( .A(n19551), .B(n19924), .Z(n19926) );
  XOR U19683 ( .A(n19932), .B(n19933), .Z(n19551) );
  AND U19684 ( .A(n376), .B(n19934), .Z(n19933) );
  XOR U19685 ( .A(n19935), .B(n19932), .Z(n19934) );
  XOR U19686 ( .A(n19936), .B(n19937), .Z(n19924) );
  AND U19687 ( .A(n19938), .B(n19939), .Z(n19937) );
  XOR U19688 ( .A(n19936), .B(n19566), .Z(n19939) );
  XOR U19689 ( .A(n19940), .B(n19941), .Z(n19566) );
  AND U19690 ( .A(n378), .B(n19942), .Z(n19941) );
  XOR U19691 ( .A(n19943), .B(n19940), .Z(n19942) );
  XNOR U19692 ( .A(n19563), .B(n19936), .Z(n19938) );
  XOR U19693 ( .A(n19944), .B(n19945), .Z(n19563) );
  AND U19694 ( .A(n376), .B(n19946), .Z(n19945) );
  XOR U19695 ( .A(n19947), .B(n19944), .Z(n19946) );
  XOR U19696 ( .A(n19948), .B(n19949), .Z(n19936) );
  AND U19697 ( .A(n19950), .B(n19951), .Z(n19949) );
  XOR U19698 ( .A(n19948), .B(n19578), .Z(n19951) );
  XOR U19699 ( .A(n19952), .B(n19953), .Z(n19578) );
  AND U19700 ( .A(n378), .B(n19954), .Z(n19953) );
  XOR U19701 ( .A(n19955), .B(n19952), .Z(n19954) );
  XNOR U19702 ( .A(n19575), .B(n19948), .Z(n19950) );
  XOR U19703 ( .A(n19956), .B(n19957), .Z(n19575) );
  AND U19704 ( .A(n376), .B(n19958), .Z(n19957) );
  XOR U19705 ( .A(n19959), .B(n19956), .Z(n19958) );
  XOR U19706 ( .A(n19960), .B(n19961), .Z(n19948) );
  AND U19707 ( .A(n19962), .B(n19963), .Z(n19961) );
  XOR U19708 ( .A(n19590), .B(n19960), .Z(n19963) );
  XOR U19709 ( .A(n19964), .B(n19965), .Z(n19590) );
  AND U19710 ( .A(n378), .B(n19966), .Z(n19965) );
  XOR U19711 ( .A(n19964), .B(n19967), .Z(n19966) );
  XNOR U19712 ( .A(n19960), .B(n19587), .Z(n19962) );
  XOR U19713 ( .A(n19968), .B(n19969), .Z(n19587) );
  AND U19714 ( .A(n376), .B(n19970), .Z(n19969) );
  XOR U19715 ( .A(n19968), .B(n19971), .Z(n19970) );
  XOR U19716 ( .A(n19972), .B(n19973), .Z(n19960) );
  AND U19717 ( .A(n19974), .B(n19975), .Z(n19973) );
  XNOR U19718 ( .A(n19976), .B(n19603), .Z(n19975) );
  XOR U19719 ( .A(n19977), .B(n19978), .Z(n19603) );
  AND U19720 ( .A(n378), .B(n19979), .Z(n19978) );
  XOR U19721 ( .A(n19980), .B(n19977), .Z(n19979) );
  XNOR U19722 ( .A(n19600), .B(n19972), .Z(n19974) );
  XOR U19723 ( .A(n19981), .B(n19982), .Z(n19600) );
  AND U19724 ( .A(n376), .B(n19983), .Z(n19982) );
  XOR U19725 ( .A(n19984), .B(n19981), .Z(n19983) );
  IV U19726 ( .A(n19976), .Z(n19972) );
  AND U19727 ( .A(n19608), .B(n19611), .Z(n19976) );
  XNOR U19728 ( .A(n19985), .B(n19986), .Z(n19611) );
  AND U19729 ( .A(n378), .B(n19987), .Z(n19986) );
  XNOR U19730 ( .A(n19988), .B(n19985), .Z(n19987) );
  XOR U19731 ( .A(n19989), .B(n19990), .Z(n378) );
  AND U19732 ( .A(n19991), .B(n19992), .Z(n19990) );
  XOR U19733 ( .A(n19619), .B(n19989), .Z(n19992) );
  IV U19734 ( .A(n19993), .Z(n19619) );
  AND U19735 ( .A(p_input[1535]), .B(p_input[1503]), .Z(n19993) );
  XOR U19736 ( .A(n19989), .B(n19616), .Z(n19991) );
  AND U19737 ( .A(p_input[1439]), .B(p_input[1471]), .Z(n19616) );
  XOR U19738 ( .A(n19994), .B(n19995), .Z(n19989) );
  AND U19739 ( .A(n19996), .B(n19997), .Z(n19995) );
  XOR U19740 ( .A(n19994), .B(n19631), .Z(n19997) );
  XNOR U19741 ( .A(p_input[1502]), .B(n19998), .Z(n19631) );
  AND U19742 ( .A(n458), .B(n19999), .Z(n19998) );
  XOR U19743 ( .A(p_input[1534]), .B(p_input[1502]), .Z(n19999) );
  XNOR U19744 ( .A(n19628), .B(n19994), .Z(n19996) );
  XOR U19745 ( .A(n20000), .B(n20001), .Z(n19628) );
  AND U19746 ( .A(n456), .B(n20002), .Z(n20001) );
  XOR U19747 ( .A(p_input[1470]), .B(p_input[1438]), .Z(n20002) );
  XOR U19748 ( .A(n20003), .B(n20004), .Z(n19994) );
  AND U19749 ( .A(n20005), .B(n20006), .Z(n20004) );
  XOR U19750 ( .A(n20003), .B(n19643), .Z(n20006) );
  XNOR U19751 ( .A(p_input[1501]), .B(n20007), .Z(n19643) );
  AND U19752 ( .A(n458), .B(n20008), .Z(n20007) );
  XOR U19753 ( .A(p_input[1533]), .B(p_input[1501]), .Z(n20008) );
  XNOR U19754 ( .A(n19640), .B(n20003), .Z(n20005) );
  XOR U19755 ( .A(n20009), .B(n20010), .Z(n19640) );
  AND U19756 ( .A(n456), .B(n20011), .Z(n20010) );
  XOR U19757 ( .A(p_input[1469]), .B(p_input[1437]), .Z(n20011) );
  XOR U19758 ( .A(n20012), .B(n20013), .Z(n20003) );
  AND U19759 ( .A(n20014), .B(n20015), .Z(n20013) );
  XOR U19760 ( .A(n20012), .B(n19655), .Z(n20015) );
  XNOR U19761 ( .A(p_input[1500]), .B(n20016), .Z(n19655) );
  AND U19762 ( .A(n458), .B(n20017), .Z(n20016) );
  XOR U19763 ( .A(p_input[1532]), .B(p_input[1500]), .Z(n20017) );
  XNOR U19764 ( .A(n19652), .B(n20012), .Z(n20014) );
  XOR U19765 ( .A(n20018), .B(n20019), .Z(n19652) );
  AND U19766 ( .A(n456), .B(n20020), .Z(n20019) );
  XOR U19767 ( .A(p_input[1468]), .B(p_input[1436]), .Z(n20020) );
  XOR U19768 ( .A(n20021), .B(n20022), .Z(n20012) );
  AND U19769 ( .A(n20023), .B(n20024), .Z(n20022) );
  XOR U19770 ( .A(n20021), .B(n19667), .Z(n20024) );
  XNOR U19771 ( .A(p_input[1499]), .B(n20025), .Z(n19667) );
  AND U19772 ( .A(n458), .B(n20026), .Z(n20025) );
  XOR U19773 ( .A(p_input[1531]), .B(p_input[1499]), .Z(n20026) );
  XNOR U19774 ( .A(n19664), .B(n20021), .Z(n20023) );
  XOR U19775 ( .A(n20027), .B(n20028), .Z(n19664) );
  AND U19776 ( .A(n456), .B(n20029), .Z(n20028) );
  XOR U19777 ( .A(p_input[1467]), .B(p_input[1435]), .Z(n20029) );
  XOR U19778 ( .A(n20030), .B(n20031), .Z(n20021) );
  AND U19779 ( .A(n20032), .B(n20033), .Z(n20031) );
  XOR U19780 ( .A(n20030), .B(n19679), .Z(n20033) );
  XNOR U19781 ( .A(p_input[1498]), .B(n20034), .Z(n19679) );
  AND U19782 ( .A(n458), .B(n20035), .Z(n20034) );
  XOR U19783 ( .A(p_input[1530]), .B(p_input[1498]), .Z(n20035) );
  XNOR U19784 ( .A(n19676), .B(n20030), .Z(n20032) );
  XOR U19785 ( .A(n20036), .B(n20037), .Z(n19676) );
  AND U19786 ( .A(n456), .B(n20038), .Z(n20037) );
  XOR U19787 ( .A(p_input[1466]), .B(p_input[1434]), .Z(n20038) );
  XOR U19788 ( .A(n20039), .B(n20040), .Z(n20030) );
  AND U19789 ( .A(n20041), .B(n20042), .Z(n20040) );
  XOR U19790 ( .A(n20039), .B(n19691), .Z(n20042) );
  XNOR U19791 ( .A(p_input[1497]), .B(n20043), .Z(n19691) );
  AND U19792 ( .A(n458), .B(n20044), .Z(n20043) );
  XOR U19793 ( .A(p_input[1529]), .B(p_input[1497]), .Z(n20044) );
  XNOR U19794 ( .A(n19688), .B(n20039), .Z(n20041) );
  XOR U19795 ( .A(n20045), .B(n20046), .Z(n19688) );
  AND U19796 ( .A(n456), .B(n20047), .Z(n20046) );
  XOR U19797 ( .A(p_input[1465]), .B(p_input[1433]), .Z(n20047) );
  XOR U19798 ( .A(n20048), .B(n20049), .Z(n20039) );
  AND U19799 ( .A(n20050), .B(n20051), .Z(n20049) );
  XOR U19800 ( .A(n20048), .B(n19703), .Z(n20051) );
  XNOR U19801 ( .A(p_input[1496]), .B(n20052), .Z(n19703) );
  AND U19802 ( .A(n458), .B(n20053), .Z(n20052) );
  XOR U19803 ( .A(p_input[1528]), .B(p_input[1496]), .Z(n20053) );
  XNOR U19804 ( .A(n19700), .B(n20048), .Z(n20050) );
  XOR U19805 ( .A(n20054), .B(n20055), .Z(n19700) );
  AND U19806 ( .A(n456), .B(n20056), .Z(n20055) );
  XOR U19807 ( .A(p_input[1464]), .B(p_input[1432]), .Z(n20056) );
  XOR U19808 ( .A(n20057), .B(n20058), .Z(n20048) );
  AND U19809 ( .A(n20059), .B(n20060), .Z(n20058) );
  XOR U19810 ( .A(n20057), .B(n19715), .Z(n20060) );
  XNOR U19811 ( .A(p_input[1495]), .B(n20061), .Z(n19715) );
  AND U19812 ( .A(n458), .B(n20062), .Z(n20061) );
  XOR U19813 ( .A(p_input[1527]), .B(p_input[1495]), .Z(n20062) );
  XNOR U19814 ( .A(n19712), .B(n20057), .Z(n20059) );
  XOR U19815 ( .A(n20063), .B(n20064), .Z(n19712) );
  AND U19816 ( .A(n456), .B(n20065), .Z(n20064) );
  XOR U19817 ( .A(p_input[1463]), .B(p_input[1431]), .Z(n20065) );
  XOR U19818 ( .A(n20066), .B(n20067), .Z(n20057) );
  AND U19819 ( .A(n20068), .B(n20069), .Z(n20067) );
  XOR U19820 ( .A(n20066), .B(n19727), .Z(n20069) );
  XNOR U19821 ( .A(p_input[1494]), .B(n20070), .Z(n19727) );
  AND U19822 ( .A(n458), .B(n20071), .Z(n20070) );
  XOR U19823 ( .A(p_input[1526]), .B(p_input[1494]), .Z(n20071) );
  XNOR U19824 ( .A(n19724), .B(n20066), .Z(n20068) );
  XOR U19825 ( .A(n20072), .B(n20073), .Z(n19724) );
  AND U19826 ( .A(n456), .B(n20074), .Z(n20073) );
  XOR U19827 ( .A(p_input[1462]), .B(p_input[1430]), .Z(n20074) );
  XOR U19828 ( .A(n20075), .B(n20076), .Z(n20066) );
  AND U19829 ( .A(n20077), .B(n20078), .Z(n20076) );
  XOR U19830 ( .A(n20075), .B(n19739), .Z(n20078) );
  XNOR U19831 ( .A(p_input[1493]), .B(n20079), .Z(n19739) );
  AND U19832 ( .A(n458), .B(n20080), .Z(n20079) );
  XOR U19833 ( .A(p_input[1525]), .B(p_input[1493]), .Z(n20080) );
  XNOR U19834 ( .A(n19736), .B(n20075), .Z(n20077) );
  XOR U19835 ( .A(n20081), .B(n20082), .Z(n19736) );
  AND U19836 ( .A(n456), .B(n20083), .Z(n20082) );
  XOR U19837 ( .A(p_input[1461]), .B(p_input[1429]), .Z(n20083) );
  XOR U19838 ( .A(n20084), .B(n20085), .Z(n20075) );
  AND U19839 ( .A(n20086), .B(n20087), .Z(n20085) );
  XOR U19840 ( .A(n20084), .B(n19751), .Z(n20087) );
  XNOR U19841 ( .A(p_input[1492]), .B(n20088), .Z(n19751) );
  AND U19842 ( .A(n458), .B(n20089), .Z(n20088) );
  XOR U19843 ( .A(p_input[1524]), .B(p_input[1492]), .Z(n20089) );
  XNOR U19844 ( .A(n19748), .B(n20084), .Z(n20086) );
  XOR U19845 ( .A(n20090), .B(n20091), .Z(n19748) );
  AND U19846 ( .A(n456), .B(n20092), .Z(n20091) );
  XOR U19847 ( .A(p_input[1460]), .B(p_input[1428]), .Z(n20092) );
  XOR U19848 ( .A(n20093), .B(n20094), .Z(n20084) );
  AND U19849 ( .A(n20095), .B(n20096), .Z(n20094) );
  XOR U19850 ( .A(n20093), .B(n19763), .Z(n20096) );
  XNOR U19851 ( .A(p_input[1491]), .B(n20097), .Z(n19763) );
  AND U19852 ( .A(n458), .B(n20098), .Z(n20097) );
  XOR U19853 ( .A(p_input[1523]), .B(p_input[1491]), .Z(n20098) );
  XNOR U19854 ( .A(n19760), .B(n20093), .Z(n20095) );
  XOR U19855 ( .A(n20099), .B(n20100), .Z(n19760) );
  AND U19856 ( .A(n456), .B(n20101), .Z(n20100) );
  XOR U19857 ( .A(p_input[1459]), .B(p_input[1427]), .Z(n20101) );
  XOR U19858 ( .A(n20102), .B(n20103), .Z(n20093) );
  AND U19859 ( .A(n20104), .B(n20105), .Z(n20103) );
  XOR U19860 ( .A(n20102), .B(n19775), .Z(n20105) );
  XNOR U19861 ( .A(p_input[1490]), .B(n20106), .Z(n19775) );
  AND U19862 ( .A(n458), .B(n20107), .Z(n20106) );
  XOR U19863 ( .A(p_input[1522]), .B(p_input[1490]), .Z(n20107) );
  XNOR U19864 ( .A(n19772), .B(n20102), .Z(n20104) );
  XOR U19865 ( .A(n20108), .B(n20109), .Z(n19772) );
  AND U19866 ( .A(n456), .B(n20110), .Z(n20109) );
  XOR U19867 ( .A(p_input[1458]), .B(p_input[1426]), .Z(n20110) );
  XOR U19868 ( .A(n20111), .B(n20112), .Z(n20102) );
  AND U19869 ( .A(n20113), .B(n20114), .Z(n20112) );
  XOR U19870 ( .A(n20111), .B(n19787), .Z(n20114) );
  XNOR U19871 ( .A(p_input[1489]), .B(n20115), .Z(n19787) );
  AND U19872 ( .A(n458), .B(n20116), .Z(n20115) );
  XOR U19873 ( .A(p_input[1521]), .B(p_input[1489]), .Z(n20116) );
  XNOR U19874 ( .A(n19784), .B(n20111), .Z(n20113) );
  XOR U19875 ( .A(n20117), .B(n20118), .Z(n19784) );
  AND U19876 ( .A(n456), .B(n20119), .Z(n20118) );
  XOR U19877 ( .A(p_input[1457]), .B(p_input[1425]), .Z(n20119) );
  XOR U19878 ( .A(n20120), .B(n20121), .Z(n20111) );
  AND U19879 ( .A(n20122), .B(n20123), .Z(n20121) );
  XOR U19880 ( .A(n20120), .B(n19799), .Z(n20123) );
  XNOR U19881 ( .A(p_input[1488]), .B(n20124), .Z(n19799) );
  AND U19882 ( .A(n458), .B(n20125), .Z(n20124) );
  XOR U19883 ( .A(p_input[1520]), .B(p_input[1488]), .Z(n20125) );
  XNOR U19884 ( .A(n19796), .B(n20120), .Z(n20122) );
  XOR U19885 ( .A(n20126), .B(n20127), .Z(n19796) );
  AND U19886 ( .A(n456), .B(n20128), .Z(n20127) );
  XOR U19887 ( .A(p_input[1456]), .B(p_input[1424]), .Z(n20128) );
  XOR U19888 ( .A(n20129), .B(n20130), .Z(n20120) );
  AND U19889 ( .A(n20131), .B(n20132), .Z(n20130) );
  XOR U19890 ( .A(n20129), .B(n19811), .Z(n20132) );
  XNOR U19891 ( .A(p_input[1487]), .B(n20133), .Z(n19811) );
  AND U19892 ( .A(n458), .B(n20134), .Z(n20133) );
  XOR U19893 ( .A(p_input[1519]), .B(p_input[1487]), .Z(n20134) );
  XNOR U19894 ( .A(n19808), .B(n20129), .Z(n20131) );
  XOR U19895 ( .A(n20135), .B(n20136), .Z(n19808) );
  AND U19896 ( .A(n456), .B(n20137), .Z(n20136) );
  XOR U19897 ( .A(p_input[1455]), .B(p_input[1423]), .Z(n20137) );
  XOR U19898 ( .A(n20138), .B(n20139), .Z(n20129) );
  AND U19899 ( .A(n20140), .B(n20141), .Z(n20139) );
  XOR U19900 ( .A(n20138), .B(n19823), .Z(n20141) );
  XNOR U19901 ( .A(p_input[1486]), .B(n20142), .Z(n19823) );
  AND U19902 ( .A(n458), .B(n20143), .Z(n20142) );
  XOR U19903 ( .A(p_input[1518]), .B(p_input[1486]), .Z(n20143) );
  XNOR U19904 ( .A(n19820), .B(n20138), .Z(n20140) );
  XOR U19905 ( .A(n20144), .B(n20145), .Z(n19820) );
  AND U19906 ( .A(n456), .B(n20146), .Z(n20145) );
  XOR U19907 ( .A(p_input[1454]), .B(p_input[1422]), .Z(n20146) );
  XOR U19908 ( .A(n20147), .B(n20148), .Z(n20138) );
  AND U19909 ( .A(n20149), .B(n20150), .Z(n20148) );
  XOR U19910 ( .A(n20147), .B(n19835), .Z(n20150) );
  XNOR U19911 ( .A(p_input[1485]), .B(n20151), .Z(n19835) );
  AND U19912 ( .A(n458), .B(n20152), .Z(n20151) );
  XOR U19913 ( .A(p_input[1517]), .B(p_input[1485]), .Z(n20152) );
  XNOR U19914 ( .A(n19832), .B(n20147), .Z(n20149) );
  XOR U19915 ( .A(n20153), .B(n20154), .Z(n19832) );
  AND U19916 ( .A(n456), .B(n20155), .Z(n20154) );
  XOR U19917 ( .A(p_input[1453]), .B(p_input[1421]), .Z(n20155) );
  XOR U19918 ( .A(n20156), .B(n20157), .Z(n20147) );
  AND U19919 ( .A(n20158), .B(n20159), .Z(n20157) );
  XOR U19920 ( .A(n20156), .B(n19847), .Z(n20159) );
  XNOR U19921 ( .A(p_input[1484]), .B(n20160), .Z(n19847) );
  AND U19922 ( .A(n458), .B(n20161), .Z(n20160) );
  XOR U19923 ( .A(p_input[1516]), .B(p_input[1484]), .Z(n20161) );
  XNOR U19924 ( .A(n19844), .B(n20156), .Z(n20158) );
  XOR U19925 ( .A(n20162), .B(n20163), .Z(n19844) );
  AND U19926 ( .A(n456), .B(n20164), .Z(n20163) );
  XOR U19927 ( .A(p_input[1452]), .B(p_input[1420]), .Z(n20164) );
  XOR U19928 ( .A(n20165), .B(n20166), .Z(n20156) );
  AND U19929 ( .A(n20167), .B(n20168), .Z(n20166) );
  XOR U19930 ( .A(n20165), .B(n19859), .Z(n20168) );
  XNOR U19931 ( .A(p_input[1483]), .B(n20169), .Z(n19859) );
  AND U19932 ( .A(n458), .B(n20170), .Z(n20169) );
  XOR U19933 ( .A(p_input[1515]), .B(p_input[1483]), .Z(n20170) );
  XNOR U19934 ( .A(n19856), .B(n20165), .Z(n20167) );
  XOR U19935 ( .A(n20171), .B(n20172), .Z(n19856) );
  AND U19936 ( .A(n456), .B(n20173), .Z(n20172) );
  XOR U19937 ( .A(p_input[1451]), .B(p_input[1419]), .Z(n20173) );
  XOR U19938 ( .A(n20174), .B(n20175), .Z(n20165) );
  AND U19939 ( .A(n20176), .B(n20177), .Z(n20175) );
  XOR U19940 ( .A(n20174), .B(n19871), .Z(n20177) );
  XNOR U19941 ( .A(p_input[1482]), .B(n20178), .Z(n19871) );
  AND U19942 ( .A(n458), .B(n20179), .Z(n20178) );
  XOR U19943 ( .A(p_input[1514]), .B(p_input[1482]), .Z(n20179) );
  XNOR U19944 ( .A(n19868), .B(n20174), .Z(n20176) );
  XOR U19945 ( .A(n20180), .B(n20181), .Z(n19868) );
  AND U19946 ( .A(n456), .B(n20182), .Z(n20181) );
  XOR U19947 ( .A(p_input[1450]), .B(p_input[1418]), .Z(n20182) );
  XOR U19948 ( .A(n20183), .B(n20184), .Z(n20174) );
  AND U19949 ( .A(n20185), .B(n20186), .Z(n20184) );
  XOR U19950 ( .A(n20183), .B(n19883), .Z(n20186) );
  XNOR U19951 ( .A(p_input[1481]), .B(n20187), .Z(n19883) );
  AND U19952 ( .A(n458), .B(n20188), .Z(n20187) );
  XOR U19953 ( .A(p_input[1513]), .B(p_input[1481]), .Z(n20188) );
  XNOR U19954 ( .A(n19880), .B(n20183), .Z(n20185) );
  XOR U19955 ( .A(n20189), .B(n20190), .Z(n19880) );
  AND U19956 ( .A(n456), .B(n20191), .Z(n20190) );
  XOR U19957 ( .A(p_input[1449]), .B(p_input[1417]), .Z(n20191) );
  XOR U19958 ( .A(n20192), .B(n20193), .Z(n20183) );
  AND U19959 ( .A(n20194), .B(n20195), .Z(n20193) );
  XOR U19960 ( .A(n20192), .B(n19895), .Z(n20195) );
  XNOR U19961 ( .A(p_input[1480]), .B(n20196), .Z(n19895) );
  AND U19962 ( .A(n458), .B(n20197), .Z(n20196) );
  XOR U19963 ( .A(p_input[1512]), .B(p_input[1480]), .Z(n20197) );
  XNOR U19964 ( .A(n19892), .B(n20192), .Z(n20194) );
  XOR U19965 ( .A(n20198), .B(n20199), .Z(n19892) );
  AND U19966 ( .A(n456), .B(n20200), .Z(n20199) );
  XOR U19967 ( .A(p_input[1448]), .B(p_input[1416]), .Z(n20200) );
  XOR U19968 ( .A(n20201), .B(n20202), .Z(n20192) );
  AND U19969 ( .A(n20203), .B(n20204), .Z(n20202) );
  XOR U19970 ( .A(n20201), .B(n19907), .Z(n20204) );
  XNOR U19971 ( .A(p_input[1479]), .B(n20205), .Z(n19907) );
  AND U19972 ( .A(n458), .B(n20206), .Z(n20205) );
  XOR U19973 ( .A(p_input[1511]), .B(p_input[1479]), .Z(n20206) );
  XNOR U19974 ( .A(n19904), .B(n20201), .Z(n20203) );
  XOR U19975 ( .A(n20207), .B(n20208), .Z(n19904) );
  AND U19976 ( .A(n456), .B(n20209), .Z(n20208) );
  XOR U19977 ( .A(p_input[1447]), .B(p_input[1415]), .Z(n20209) );
  XOR U19978 ( .A(n20210), .B(n20211), .Z(n20201) );
  AND U19979 ( .A(n20212), .B(n20213), .Z(n20211) );
  XOR U19980 ( .A(n20210), .B(n19919), .Z(n20213) );
  XNOR U19981 ( .A(p_input[1478]), .B(n20214), .Z(n19919) );
  AND U19982 ( .A(n458), .B(n20215), .Z(n20214) );
  XOR U19983 ( .A(p_input[1510]), .B(p_input[1478]), .Z(n20215) );
  XNOR U19984 ( .A(n19916), .B(n20210), .Z(n20212) );
  XOR U19985 ( .A(n20216), .B(n20217), .Z(n19916) );
  AND U19986 ( .A(n456), .B(n20218), .Z(n20217) );
  XOR U19987 ( .A(p_input[1446]), .B(p_input[1414]), .Z(n20218) );
  XOR U19988 ( .A(n20219), .B(n20220), .Z(n20210) );
  AND U19989 ( .A(n20221), .B(n20222), .Z(n20220) );
  XOR U19990 ( .A(n20219), .B(n19931), .Z(n20222) );
  XNOR U19991 ( .A(p_input[1477]), .B(n20223), .Z(n19931) );
  AND U19992 ( .A(n458), .B(n20224), .Z(n20223) );
  XOR U19993 ( .A(p_input[1509]), .B(p_input[1477]), .Z(n20224) );
  XNOR U19994 ( .A(n19928), .B(n20219), .Z(n20221) );
  XOR U19995 ( .A(n20225), .B(n20226), .Z(n19928) );
  AND U19996 ( .A(n456), .B(n20227), .Z(n20226) );
  XOR U19997 ( .A(p_input[1445]), .B(p_input[1413]), .Z(n20227) );
  XOR U19998 ( .A(n20228), .B(n20229), .Z(n20219) );
  AND U19999 ( .A(n20230), .B(n20231), .Z(n20229) );
  XOR U20000 ( .A(n20228), .B(n19943), .Z(n20231) );
  XNOR U20001 ( .A(p_input[1476]), .B(n20232), .Z(n19943) );
  AND U20002 ( .A(n458), .B(n20233), .Z(n20232) );
  XOR U20003 ( .A(p_input[1508]), .B(p_input[1476]), .Z(n20233) );
  XNOR U20004 ( .A(n19940), .B(n20228), .Z(n20230) );
  XOR U20005 ( .A(n20234), .B(n20235), .Z(n19940) );
  AND U20006 ( .A(n456), .B(n20236), .Z(n20235) );
  XOR U20007 ( .A(p_input[1444]), .B(p_input[1412]), .Z(n20236) );
  XOR U20008 ( .A(n20237), .B(n20238), .Z(n20228) );
  AND U20009 ( .A(n20239), .B(n20240), .Z(n20238) );
  XOR U20010 ( .A(n20237), .B(n19955), .Z(n20240) );
  XNOR U20011 ( .A(p_input[1475]), .B(n20241), .Z(n19955) );
  AND U20012 ( .A(n458), .B(n20242), .Z(n20241) );
  XOR U20013 ( .A(p_input[1507]), .B(p_input[1475]), .Z(n20242) );
  XNOR U20014 ( .A(n19952), .B(n20237), .Z(n20239) );
  XOR U20015 ( .A(n20243), .B(n20244), .Z(n19952) );
  AND U20016 ( .A(n456), .B(n20245), .Z(n20244) );
  XOR U20017 ( .A(p_input[1443]), .B(p_input[1411]), .Z(n20245) );
  XOR U20018 ( .A(n20246), .B(n20247), .Z(n20237) );
  AND U20019 ( .A(n20248), .B(n20249), .Z(n20247) );
  XOR U20020 ( .A(n19967), .B(n20246), .Z(n20249) );
  XNOR U20021 ( .A(p_input[1474]), .B(n20250), .Z(n19967) );
  AND U20022 ( .A(n458), .B(n20251), .Z(n20250) );
  XOR U20023 ( .A(p_input[1506]), .B(p_input[1474]), .Z(n20251) );
  XNOR U20024 ( .A(n20246), .B(n19964), .Z(n20248) );
  XOR U20025 ( .A(n20252), .B(n20253), .Z(n19964) );
  AND U20026 ( .A(n456), .B(n20254), .Z(n20253) );
  XOR U20027 ( .A(p_input[1442]), .B(p_input[1410]), .Z(n20254) );
  XOR U20028 ( .A(n20255), .B(n20256), .Z(n20246) );
  AND U20029 ( .A(n20257), .B(n20258), .Z(n20256) );
  XNOR U20030 ( .A(n20259), .B(n19980), .Z(n20258) );
  XNOR U20031 ( .A(p_input[1473]), .B(n20260), .Z(n19980) );
  AND U20032 ( .A(n458), .B(n20261), .Z(n20260) );
  XNOR U20033 ( .A(p_input[1505]), .B(n20262), .Z(n20261) );
  IV U20034 ( .A(p_input[1473]), .Z(n20262) );
  XNOR U20035 ( .A(n19977), .B(n20255), .Z(n20257) );
  XNOR U20036 ( .A(p_input[1409]), .B(n20263), .Z(n19977) );
  AND U20037 ( .A(n456), .B(n20264), .Z(n20263) );
  XOR U20038 ( .A(p_input[1441]), .B(p_input[1409]), .Z(n20264) );
  IV U20039 ( .A(n20259), .Z(n20255) );
  AND U20040 ( .A(n19985), .B(n19988), .Z(n20259) );
  XOR U20041 ( .A(p_input[1472]), .B(n20265), .Z(n19988) );
  AND U20042 ( .A(n458), .B(n20266), .Z(n20265) );
  XOR U20043 ( .A(p_input[1504]), .B(p_input[1472]), .Z(n20266) );
  XOR U20044 ( .A(n20267), .B(n20268), .Z(n458) );
  AND U20045 ( .A(n20269), .B(n20270), .Z(n20268) );
  XNOR U20046 ( .A(p_input[1535]), .B(n20267), .Z(n20270) );
  XOR U20047 ( .A(n20267), .B(p_input[1503]), .Z(n20269) );
  XOR U20048 ( .A(n20271), .B(n20272), .Z(n20267) );
  AND U20049 ( .A(n20273), .B(n20274), .Z(n20272) );
  XNOR U20050 ( .A(p_input[1534]), .B(n20271), .Z(n20274) );
  XOR U20051 ( .A(n20271), .B(p_input[1502]), .Z(n20273) );
  XOR U20052 ( .A(n20275), .B(n20276), .Z(n20271) );
  AND U20053 ( .A(n20277), .B(n20278), .Z(n20276) );
  XNOR U20054 ( .A(p_input[1533]), .B(n20275), .Z(n20278) );
  XOR U20055 ( .A(n20275), .B(p_input[1501]), .Z(n20277) );
  XOR U20056 ( .A(n20279), .B(n20280), .Z(n20275) );
  AND U20057 ( .A(n20281), .B(n20282), .Z(n20280) );
  XNOR U20058 ( .A(p_input[1532]), .B(n20279), .Z(n20282) );
  XOR U20059 ( .A(n20279), .B(p_input[1500]), .Z(n20281) );
  XOR U20060 ( .A(n20283), .B(n20284), .Z(n20279) );
  AND U20061 ( .A(n20285), .B(n20286), .Z(n20284) );
  XNOR U20062 ( .A(p_input[1531]), .B(n20283), .Z(n20286) );
  XOR U20063 ( .A(n20283), .B(p_input[1499]), .Z(n20285) );
  XOR U20064 ( .A(n20287), .B(n20288), .Z(n20283) );
  AND U20065 ( .A(n20289), .B(n20290), .Z(n20288) );
  XNOR U20066 ( .A(p_input[1530]), .B(n20287), .Z(n20290) );
  XOR U20067 ( .A(n20287), .B(p_input[1498]), .Z(n20289) );
  XOR U20068 ( .A(n20291), .B(n20292), .Z(n20287) );
  AND U20069 ( .A(n20293), .B(n20294), .Z(n20292) );
  XNOR U20070 ( .A(p_input[1529]), .B(n20291), .Z(n20294) );
  XOR U20071 ( .A(n20291), .B(p_input[1497]), .Z(n20293) );
  XOR U20072 ( .A(n20295), .B(n20296), .Z(n20291) );
  AND U20073 ( .A(n20297), .B(n20298), .Z(n20296) );
  XNOR U20074 ( .A(p_input[1528]), .B(n20295), .Z(n20298) );
  XOR U20075 ( .A(n20295), .B(p_input[1496]), .Z(n20297) );
  XOR U20076 ( .A(n20299), .B(n20300), .Z(n20295) );
  AND U20077 ( .A(n20301), .B(n20302), .Z(n20300) );
  XNOR U20078 ( .A(p_input[1527]), .B(n20299), .Z(n20302) );
  XOR U20079 ( .A(n20299), .B(p_input[1495]), .Z(n20301) );
  XOR U20080 ( .A(n20303), .B(n20304), .Z(n20299) );
  AND U20081 ( .A(n20305), .B(n20306), .Z(n20304) );
  XNOR U20082 ( .A(p_input[1526]), .B(n20303), .Z(n20306) );
  XOR U20083 ( .A(n20303), .B(p_input[1494]), .Z(n20305) );
  XOR U20084 ( .A(n20307), .B(n20308), .Z(n20303) );
  AND U20085 ( .A(n20309), .B(n20310), .Z(n20308) );
  XNOR U20086 ( .A(p_input[1525]), .B(n20307), .Z(n20310) );
  XOR U20087 ( .A(n20307), .B(p_input[1493]), .Z(n20309) );
  XOR U20088 ( .A(n20311), .B(n20312), .Z(n20307) );
  AND U20089 ( .A(n20313), .B(n20314), .Z(n20312) );
  XNOR U20090 ( .A(p_input[1524]), .B(n20311), .Z(n20314) );
  XOR U20091 ( .A(n20311), .B(p_input[1492]), .Z(n20313) );
  XOR U20092 ( .A(n20315), .B(n20316), .Z(n20311) );
  AND U20093 ( .A(n20317), .B(n20318), .Z(n20316) );
  XNOR U20094 ( .A(p_input[1523]), .B(n20315), .Z(n20318) );
  XOR U20095 ( .A(n20315), .B(p_input[1491]), .Z(n20317) );
  XOR U20096 ( .A(n20319), .B(n20320), .Z(n20315) );
  AND U20097 ( .A(n20321), .B(n20322), .Z(n20320) );
  XNOR U20098 ( .A(p_input[1522]), .B(n20319), .Z(n20322) );
  XOR U20099 ( .A(n20319), .B(p_input[1490]), .Z(n20321) );
  XOR U20100 ( .A(n20323), .B(n20324), .Z(n20319) );
  AND U20101 ( .A(n20325), .B(n20326), .Z(n20324) );
  XNOR U20102 ( .A(p_input[1521]), .B(n20323), .Z(n20326) );
  XOR U20103 ( .A(n20323), .B(p_input[1489]), .Z(n20325) );
  XOR U20104 ( .A(n20327), .B(n20328), .Z(n20323) );
  AND U20105 ( .A(n20329), .B(n20330), .Z(n20328) );
  XNOR U20106 ( .A(p_input[1520]), .B(n20327), .Z(n20330) );
  XOR U20107 ( .A(n20327), .B(p_input[1488]), .Z(n20329) );
  XOR U20108 ( .A(n20331), .B(n20332), .Z(n20327) );
  AND U20109 ( .A(n20333), .B(n20334), .Z(n20332) );
  XNOR U20110 ( .A(p_input[1519]), .B(n20331), .Z(n20334) );
  XOR U20111 ( .A(n20331), .B(p_input[1487]), .Z(n20333) );
  XOR U20112 ( .A(n20335), .B(n20336), .Z(n20331) );
  AND U20113 ( .A(n20337), .B(n20338), .Z(n20336) );
  XNOR U20114 ( .A(p_input[1518]), .B(n20335), .Z(n20338) );
  XOR U20115 ( .A(n20335), .B(p_input[1486]), .Z(n20337) );
  XOR U20116 ( .A(n20339), .B(n20340), .Z(n20335) );
  AND U20117 ( .A(n20341), .B(n20342), .Z(n20340) );
  XNOR U20118 ( .A(p_input[1517]), .B(n20339), .Z(n20342) );
  XOR U20119 ( .A(n20339), .B(p_input[1485]), .Z(n20341) );
  XOR U20120 ( .A(n20343), .B(n20344), .Z(n20339) );
  AND U20121 ( .A(n20345), .B(n20346), .Z(n20344) );
  XNOR U20122 ( .A(p_input[1516]), .B(n20343), .Z(n20346) );
  XOR U20123 ( .A(n20343), .B(p_input[1484]), .Z(n20345) );
  XOR U20124 ( .A(n20347), .B(n20348), .Z(n20343) );
  AND U20125 ( .A(n20349), .B(n20350), .Z(n20348) );
  XNOR U20126 ( .A(p_input[1515]), .B(n20347), .Z(n20350) );
  XOR U20127 ( .A(n20347), .B(p_input[1483]), .Z(n20349) );
  XOR U20128 ( .A(n20351), .B(n20352), .Z(n20347) );
  AND U20129 ( .A(n20353), .B(n20354), .Z(n20352) );
  XNOR U20130 ( .A(p_input[1514]), .B(n20351), .Z(n20354) );
  XOR U20131 ( .A(n20351), .B(p_input[1482]), .Z(n20353) );
  XOR U20132 ( .A(n20355), .B(n20356), .Z(n20351) );
  AND U20133 ( .A(n20357), .B(n20358), .Z(n20356) );
  XNOR U20134 ( .A(p_input[1513]), .B(n20355), .Z(n20358) );
  XOR U20135 ( .A(n20355), .B(p_input[1481]), .Z(n20357) );
  XOR U20136 ( .A(n20359), .B(n20360), .Z(n20355) );
  AND U20137 ( .A(n20361), .B(n20362), .Z(n20360) );
  XNOR U20138 ( .A(p_input[1512]), .B(n20359), .Z(n20362) );
  XOR U20139 ( .A(n20359), .B(p_input[1480]), .Z(n20361) );
  XOR U20140 ( .A(n20363), .B(n20364), .Z(n20359) );
  AND U20141 ( .A(n20365), .B(n20366), .Z(n20364) );
  XNOR U20142 ( .A(p_input[1511]), .B(n20363), .Z(n20366) );
  XOR U20143 ( .A(n20363), .B(p_input[1479]), .Z(n20365) );
  XOR U20144 ( .A(n20367), .B(n20368), .Z(n20363) );
  AND U20145 ( .A(n20369), .B(n20370), .Z(n20368) );
  XNOR U20146 ( .A(p_input[1510]), .B(n20367), .Z(n20370) );
  XOR U20147 ( .A(n20367), .B(p_input[1478]), .Z(n20369) );
  XOR U20148 ( .A(n20371), .B(n20372), .Z(n20367) );
  AND U20149 ( .A(n20373), .B(n20374), .Z(n20372) );
  XNOR U20150 ( .A(p_input[1509]), .B(n20371), .Z(n20374) );
  XOR U20151 ( .A(n20371), .B(p_input[1477]), .Z(n20373) );
  XOR U20152 ( .A(n20375), .B(n20376), .Z(n20371) );
  AND U20153 ( .A(n20377), .B(n20378), .Z(n20376) );
  XNOR U20154 ( .A(p_input[1508]), .B(n20375), .Z(n20378) );
  XOR U20155 ( .A(n20375), .B(p_input[1476]), .Z(n20377) );
  XOR U20156 ( .A(n20379), .B(n20380), .Z(n20375) );
  AND U20157 ( .A(n20381), .B(n20382), .Z(n20380) );
  XNOR U20158 ( .A(p_input[1507]), .B(n20379), .Z(n20382) );
  XOR U20159 ( .A(n20379), .B(p_input[1475]), .Z(n20381) );
  XOR U20160 ( .A(n20383), .B(n20384), .Z(n20379) );
  AND U20161 ( .A(n20385), .B(n20386), .Z(n20384) );
  XNOR U20162 ( .A(p_input[1506]), .B(n20383), .Z(n20386) );
  XOR U20163 ( .A(n20383), .B(p_input[1474]), .Z(n20385) );
  XNOR U20164 ( .A(n20387), .B(n20388), .Z(n20383) );
  AND U20165 ( .A(n20389), .B(n20390), .Z(n20388) );
  XOR U20166 ( .A(p_input[1505]), .B(n20387), .Z(n20390) );
  XNOR U20167 ( .A(p_input[1473]), .B(n20387), .Z(n20389) );
  AND U20168 ( .A(p_input[1504]), .B(n20391), .Z(n20387) );
  IV U20169 ( .A(p_input[1472]), .Z(n20391) );
  XNOR U20170 ( .A(p_input[1408]), .B(n20392), .Z(n19985) );
  AND U20171 ( .A(n456), .B(n20393), .Z(n20392) );
  XOR U20172 ( .A(p_input[1440]), .B(p_input[1408]), .Z(n20393) );
  XOR U20173 ( .A(n20394), .B(n20395), .Z(n456) );
  AND U20174 ( .A(n20396), .B(n20397), .Z(n20395) );
  XNOR U20175 ( .A(p_input[1471]), .B(n20394), .Z(n20397) );
  XOR U20176 ( .A(n20394), .B(p_input[1439]), .Z(n20396) );
  XOR U20177 ( .A(n20398), .B(n20399), .Z(n20394) );
  AND U20178 ( .A(n20400), .B(n20401), .Z(n20399) );
  XNOR U20179 ( .A(p_input[1470]), .B(n20398), .Z(n20401) );
  XNOR U20180 ( .A(n20398), .B(n20000), .Z(n20400) );
  IV U20181 ( .A(p_input[1438]), .Z(n20000) );
  XOR U20182 ( .A(n20402), .B(n20403), .Z(n20398) );
  AND U20183 ( .A(n20404), .B(n20405), .Z(n20403) );
  XNOR U20184 ( .A(p_input[1469]), .B(n20402), .Z(n20405) );
  XNOR U20185 ( .A(n20402), .B(n20009), .Z(n20404) );
  IV U20186 ( .A(p_input[1437]), .Z(n20009) );
  XOR U20187 ( .A(n20406), .B(n20407), .Z(n20402) );
  AND U20188 ( .A(n20408), .B(n20409), .Z(n20407) );
  XNOR U20189 ( .A(p_input[1468]), .B(n20406), .Z(n20409) );
  XNOR U20190 ( .A(n20406), .B(n20018), .Z(n20408) );
  IV U20191 ( .A(p_input[1436]), .Z(n20018) );
  XOR U20192 ( .A(n20410), .B(n20411), .Z(n20406) );
  AND U20193 ( .A(n20412), .B(n20413), .Z(n20411) );
  XNOR U20194 ( .A(p_input[1467]), .B(n20410), .Z(n20413) );
  XNOR U20195 ( .A(n20410), .B(n20027), .Z(n20412) );
  IV U20196 ( .A(p_input[1435]), .Z(n20027) );
  XOR U20197 ( .A(n20414), .B(n20415), .Z(n20410) );
  AND U20198 ( .A(n20416), .B(n20417), .Z(n20415) );
  XNOR U20199 ( .A(p_input[1466]), .B(n20414), .Z(n20417) );
  XNOR U20200 ( .A(n20414), .B(n20036), .Z(n20416) );
  IV U20201 ( .A(p_input[1434]), .Z(n20036) );
  XOR U20202 ( .A(n20418), .B(n20419), .Z(n20414) );
  AND U20203 ( .A(n20420), .B(n20421), .Z(n20419) );
  XNOR U20204 ( .A(p_input[1465]), .B(n20418), .Z(n20421) );
  XNOR U20205 ( .A(n20418), .B(n20045), .Z(n20420) );
  IV U20206 ( .A(p_input[1433]), .Z(n20045) );
  XOR U20207 ( .A(n20422), .B(n20423), .Z(n20418) );
  AND U20208 ( .A(n20424), .B(n20425), .Z(n20423) );
  XNOR U20209 ( .A(p_input[1464]), .B(n20422), .Z(n20425) );
  XNOR U20210 ( .A(n20422), .B(n20054), .Z(n20424) );
  IV U20211 ( .A(p_input[1432]), .Z(n20054) );
  XOR U20212 ( .A(n20426), .B(n20427), .Z(n20422) );
  AND U20213 ( .A(n20428), .B(n20429), .Z(n20427) );
  XNOR U20214 ( .A(p_input[1463]), .B(n20426), .Z(n20429) );
  XNOR U20215 ( .A(n20426), .B(n20063), .Z(n20428) );
  IV U20216 ( .A(p_input[1431]), .Z(n20063) );
  XOR U20217 ( .A(n20430), .B(n20431), .Z(n20426) );
  AND U20218 ( .A(n20432), .B(n20433), .Z(n20431) );
  XNOR U20219 ( .A(p_input[1462]), .B(n20430), .Z(n20433) );
  XNOR U20220 ( .A(n20430), .B(n20072), .Z(n20432) );
  IV U20221 ( .A(p_input[1430]), .Z(n20072) );
  XOR U20222 ( .A(n20434), .B(n20435), .Z(n20430) );
  AND U20223 ( .A(n20436), .B(n20437), .Z(n20435) );
  XNOR U20224 ( .A(p_input[1461]), .B(n20434), .Z(n20437) );
  XNOR U20225 ( .A(n20434), .B(n20081), .Z(n20436) );
  IV U20226 ( .A(p_input[1429]), .Z(n20081) );
  XOR U20227 ( .A(n20438), .B(n20439), .Z(n20434) );
  AND U20228 ( .A(n20440), .B(n20441), .Z(n20439) );
  XNOR U20229 ( .A(p_input[1460]), .B(n20438), .Z(n20441) );
  XNOR U20230 ( .A(n20438), .B(n20090), .Z(n20440) );
  IV U20231 ( .A(p_input[1428]), .Z(n20090) );
  XOR U20232 ( .A(n20442), .B(n20443), .Z(n20438) );
  AND U20233 ( .A(n20444), .B(n20445), .Z(n20443) );
  XNOR U20234 ( .A(p_input[1459]), .B(n20442), .Z(n20445) );
  XNOR U20235 ( .A(n20442), .B(n20099), .Z(n20444) );
  IV U20236 ( .A(p_input[1427]), .Z(n20099) );
  XOR U20237 ( .A(n20446), .B(n20447), .Z(n20442) );
  AND U20238 ( .A(n20448), .B(n20449), .Z(n20447) );
  XNOR U20239 ( .A(p_input[1458]), .B(n20446), .Z(n20449) );
  XNOR U20240 ( .A(n20446), .B(n20108), .Z(n20448) );
  IV U20241 ( .A(p_input[1426]), .Z(n20108) );
  XOR U20242 ( .A(n20450), .B(n20451), .Z(n20446) );
  AND U20243 ( .A(n20452), .B(n20453), .Z(n20451) );
  XNOR U20244 ( .A(p_input[1457]), .B(n20450), .Z(n20453) );
  XNOR U20245 ( .A(n20450), .B(n20117), .Z(n20452) );
  IV U20246 ( .A(p_input[1425]), .Z(n20117) );
  XOR U20247 ( .A(n20454), .B(n20455), .Z(n20450) );
  AND U20248 ( .A(n20456), .B(n20457), .Z(n20455) );
  XNOR U20249 ( .A(p_input[1456]), .B(n20454), .Z(n20457) );
  XNOR U20250 ( .A(n20454), .B(n20126), .Z(n20456) );
  IV U20251 ( .A(p_input[1424]), .Z(n20126) );
  XOR U20252 ( .A(n20458), .B(n20459), .Z(n20454) );
  AND U20253 ( .A(n20460), .B(n20461), .Z(n20459) );
  XNOR U20254 ( .A(p_input[1455]), .B(n20458), .Z(n20461) );
  XNOR U20255 ( .A(n20458), .B(n20135), .Z(n20460) );
  IV U20256 ( .A(p_input[1423]), .Z(n20135) );
  XOR U20257 ( .A(n20462), .B(n20463), .Z(n20458) );
  AND U20258 ( .A(n20464), .B(n20465), .Z(n20463) );
  XNOR U20259 ( .A(p_input[1454]), .B(n20462), .Z(n20465) );
  XNOR U20260 ( .A(n20462), .B(n20144), .Z(n20464) );
  IV U20261 ( .A(p_input[1422]), .Z(n20144) );
  XOR U20262 ( .A(n20466), .B(n20467), .Z(n20462) );
  AND U20263 ( .A(n20468), .B(n20469), .Z(n20467) );
  XNOR U20264 ( .A(p_input[1453]), .B(n20466), .Z(n20469) );
  XNOR U20265 ( .A(n20466), .B(n20153), .Z(n20468) );
  IV U20266 ( .A(p_input[1421]), .Z(n20153) );
  XOR U20267 ( .A(n20470), .B(n20471), .Z(n20466) );
  AND U20268 ( .A(n20472), .B(n20473), .Z(n20471) );
  XNOR U20269 ( .A(p_input[1452]), .B(n20470), .Z(n20473) );
  XNOR U20270 ( .A(n20470), .B(n20162), .Z(n20472) );
  IV U20271 ( .A(p_input[1420]), .Z(n20162) );
  XOR U20272 ( .A(n20474), .B(n20475), .Z(n20470) );
  AND U20273 ( .A(n20476), .B(n20477), .Z(n20475) );
  XNOR U20274 ( .A(p_input[1451]), .B(n20474), .Z(n20477) );
  XNOR U20275 ( .A(n20474), .B(n20171), .Z(n20476) );
  IV U20276 ( .A(p_input[1419]), .Z(n20171) );
  XOR U20277 ( .A(n20478), .B(n20479), .Z(n20474) );
  AND U20278 ( .A(n20480), .B(n20481), .Z(n20479) );
  XNOR U20279 ( .A(p_input[1450]), .B(n20478), .Z(n20481) );
  XNOR U20280 ( .A(n20478), .B(n20180), .Z(n20480) );
  IV U20281 ( .A(p_input[1418]), .Z(n20180) );
  XOR U20282 ( .A(n20482), .B(n20483), .Z(n20478) );
  AND U20283 ( .A(n20484), .B(n20485), .Z(n20483) );
  XNOR U20284 ( .A(p_input[1449]), .B(n20482), .Z(n20485) );
  XNOR U20285 ( .A(n20482), .B(n20189), .Z(n20484) );
  IV U20286 ( .A(p_input[1417]), .Z(n20189) );
  XOR U20287 ( .A(n20486), .B(n20487), .Z(n20482) );
  AND U20288 ( .A(n20488), .B(n20489), .Z(n20487) );
  XNOR U20289 ( .A(p_input[1448]), .B(n20486), .Z(n20489) );
  XNOR U20290 ( .A(n20486), .B(n20198), .Z(n20488) );
  IV U20291 ( .A(p_input[1416]), .Z(n20198) );
  XOR U20292 ( .A(n20490), .B(n20491), .Z(n20486) );
  AND U20293 ( .A(n20492), .B(n20493), .Z(n20491) );
  XNOR U20294 ( .A(p_input[1447]), .B(n20490), .Z(n20493) );
  XNOR U20295 ( .A(n20490), .B(n20207), .Z(n20492) );
  IV U20296 ( .A(p_input[1415]), .Z(n20207) );
  XOR U20297 ( .A(n20494), .B(n20495), .Z(n20490) );
  AND U20298 ( .A(n20496), .B(n20497), .Z(n20495) );
  XNOR U20299 ( .A(p_input[1446]), .B(n20494), .Z(n20497) );
  XNOR U20300 ( .A(n20494), .B(n20216), .Z(n20496) );
  IV U20301 ( .A(p_input[1414]), .Z(n20216) );
  XOR U20302 ( .A(n20498), .B(n20499), .Z(n20494) );
  AND U20303 ( .A(n20500), .B(n20501), .Z(n20499) );
  XNOR U20304 ( .A(p_input[1445]), .B(n20498), .Z(n20501) );
  XNOR U20305 ( .A(n20498), .B(n20225), .Z(n20500) );
  IV U20306 ( .A(p_input[1413]), .Z(n20225) );
  XOR U20307 ( .A(n20502), .B(n20503), .Z(n20498) );
  AND U20308 ( .A(n20504), .B(n20505), .Z(n20503) );
  XNOR U20309 ( .A(p_input[1444]), .B(n20502), .Z(n20505) );
  XNOR U20310 ( .A(n20502), .B(n20234), .Z(n20504) );
  IV U20311 ( .A(p_input[1412]), .Z(n20234) );
  XOR U20312 ( .A(n20506), .B(n20507), .Z(n20502) );
  AND U20313 ( .A(n20508), .B(n20509), .Z(n20507) );
  XNOR U20314 ( .A(p_input[1443]), .B(n20506), .Z(n20509) );
  XNOR U20315 ( .A(n20506), .B(n20243), .Z(n20508) );
  IV U20316 ( .A(p_input[1411]), .Z(n20243) );
  XOR U20317 ( .A(n20510), .B(n20511), .Z(n20506) );
  AND U20318 ( .A(n20512), .B(n20513), .Z(n20511) );
  XNOR U20319 ( .A(p_input[1442]), .B(n20510), .Z(n20513) );
  XNOR U20320 ( .A(n20510), .B(n20252), .Z(n20512) );
  IV U20321 ( .A(p_input[1410]), .Z(n20252) );
  XNOR U20322 ( .A(n20514), .B(n20515), .Z(n20510) );
  AND U20323 ( .A(n20516), .B(n20517), .Z(n20515) );
  XOR U20324 ( .A(p_input[1441]), .B(n20514), .Z(n20517) );
  XNOR U20325 ( .A(p_input[1409]), .B(n20514), .Z(n20516) );
  AND U20326 ( .A(p_input[1440]), .B(n20518), .Z(n20514) );
  IV U20327 ( .A(p_input[1408]), .Z(n20518) );
  XOR U20328 ( .A(n20519), .B(n20520), .Z(n19608) );
  AND U20329 ( .A(n376), .B(n20521), .Z(n20520) );
  XNOR U20330 ( .A(n20522), .B(n20519), .Z(n20521) );
  XOR U20331 ( .A(n20523), .B(n20524), .Z(n376) );
  AND U20332 ( .A(n20525), .B(n20526), .Z(n20524) );
  XNOR U20333 ( .A(n19623), .B(n20523), .Z(n20526) );
  AND U20334 ( .A(p_input[1407]), .B(p_input[1375]), .Z(n19623) );
  XNOR U20335 ( .A(n20523), .B(n19620), .Z(n20525) );
  IV U20336 ( .A(n20527), .Z(n19620) );
  AND U20337 ( .A(p_input[1311]), .B(p_input[1343]), .Z(n20527) );
  XOR U20338 ( .A(n20528), .B(n20529), .Z(n20523) );
  AND U20339 ( .A(n20530), .B(n20531), .Z(n20529) );
  XOR U20340 ( .A(n20528), .B(n19635), .Z(n20531) );
  XNOR U20341 ( .A(p_input[1374]), .B(n20532), .Z(n19635) );
  AND U20342 ( .A(n462), .B(n20533), .Z(n20532) );
  XOR U20343 ( .A(p_input[1406]), .B(p_input[1374]), .Z(n20533) );
  XNOR U20344 ( .A(n19632), .B(n20528), .Z(n20530) );
  XOR U20345 ( .A(n20534), .B(n20535), .Z(n19632) );
  AND U20346 ( .A(n459), .B(n20536), .Z(n20535) );
  XOR U20347 ( .A(p_input[1342]), .B(p_input[1310]), .Z(n20536) );
  XOR U20348 ( .A(n20537), .B(n20538), .Z(n20528) );
  AND U20349 ( .A(n20539), .B(n20540), .Z(n20538) );
  XOR U20350 ( .A(n20537), .B(n19647), .Z(n20540) );
  XNOR U20351 ( .A(p_input[1373]), .B(n20541), .Z(n19647) );
  AND U20352 ( .A(n462), .B(n20542), .Z(n20541) );
  XOR U20353 ( .A(p_input[1405]), .B(p_input[1373]), .Z(n20542) );
  XNOR U20354 ( .A(n19644), .B(n20537), .Z(n20539) );
  XOR U20355 ( .A(n20543), .B(n20544), .Z(n19644) );
  AND U20356 ( .A(n459), .B(n20545), .Z(n20544) );
  XOR U20357 ( .A(p_input[1341]), .B(p_input[1309]), .Z(n20545) );
  XOR U20358 ( .A(n20546), .B(n20547), .Z(n20537) );
  AND U20359 ( .A(n20548), .B(n20549), .Z(n20547) );
  XOR U20360 ( .A(n20546), .B(n19659), .Z(n20549) );
  XNOR U20361 ( .A(p_input[1372]), .B(n20550), .Z(n19659) );
  AND U20362 ( .A(n462), .B(n20551), .Z(n20550) );
  XOR U20363 ( .A(p_input[1404]), .B(p_input[1372]), .Z(n20551) );
  XNOR U20364 ( .A(n19656), .B(n20546), .Z(n20548) );
  XOR U20365 ( .A(n20552), .B(n20553), .Z(n19656) );
  AND U20366 ( .A(n459), .B(n20554), .Z(n20553) );
  XOR U20367 ( .A(p_input[1340]), .B(p_input[1308]), .Z(n20554) );
  XOR U20368 ( .A(n20555), .B(n20556), .Z(n20546) );
  AND U20369 ( .A(n20557), .B(n20558), .Z(n20556) );
  XOR U20370 ( .A(n20555), .B(n19671), .Z(n20558) );
  XNOR U20371 ( .A(p_input[1371]), .B(n20559), .Z(n19671) );
  AND U20372 ( .A(n462), .B(n20560), .Z(n20559) );
  XOR U20373 ( .A(p_input[1403]), .B(p_input[1371]), .Z(n20560) );
  XNOR U20374 ( .A(n19668), .B(n20555), .Z(n20557) );
  XOR U20375 ( .A(n20561), .B(n20562), .Z(n19668) );
  AND U20376 ( .A(n459), .B(n20563), .Z(n20562) );
  XOR U20377 ( .A(p_input[1339]), .B(p_input[1307]), .Z(n20563) );
  XOR U20378 ( .A(n20564), .B(n20565), .Z(n20555) );
  AND U20379 ( .A(n20566), .B(n20567), .Z(n20565) );
  XOR U20380 ( .A(n20564), .B(n19683), .Z(n20567) );
  XNOR U20381 ( .A(p_input[1370]), .B(n20568), .Z(n19683) );
  AND U20382 ( .A(n462), .B(n20569), .Z(n20568) );
  XOR U20383 ( .A(p_input[1402]), .B(p_input[1370]), .Z(n20569) );
  XNOR U20384 ( .A(n19680), .B(n20564), .Z(n20566) );
  XOR U20385 ( .A(n20570), .B(n20571), .Z(n19680) );
  AND U20386 ( .A(n459), .B(n20572), .Z(n20571) );
  XOR U20387 ( .A(p_input[1338]), .B(p_input[1306]), .Z(n20572) );
  XOR U20388 ( .A(n20573), .B(n20574), .Z(n20564) );
  AND U20389 ( .A(n20575), .B(n20576), .Z(n20574) );
  XOR U20390 ( .A(n20573), .B(n19695), .Z(n20576) );
  XNOR U20391 ( .A(p_input[1369]), .B(n20577), .Z(n19695) );
  AND U20392 ( .A(n462), .B(n20578), .Z(n20577) );
  XOR U20393 ( .A(p_input[1401]), .B(p_input[1369]), .Z(n20578) );
  XNOR U20394 ( .A(n19692), .B(n20573), .Z(n20575) );
  XOR U20395 ( .A(n20579), .B(n20580), .Z(n19692) );
  AND U20396 ( .A(n459), .B(n20581), .Z(n20580) );
  XOR U20397 ( .A(p_input[1337]), .B(p_input[1305]), .Z(n20581) );
  XOR U20398 ( .A(n20582), .B(n20583), .Z(n20573) );
  AND U20399 ( .A(n20584), .B(n20585), .Z(n20583) );
  XOR U20400 ( .A(n20582), .B(n19707), .Z(n20585) );
  XNOR U20401 ( .A(p_input[1368]), .B(n20586), .Z(n19707) );
  AND U20402 ( .A(n462), .B(n20587), .Z(n20586) );
  XOR U20403 ( .A(p_input[1400]), .B(p_input[1368]), .Z(n20587) );
  XNOR U20404 ( .A(n19704), .B(n20582), .Z(n20584) );
  XOR U20405 ( .A(n20588), .B(n20589), .Z(n19704) );
  AND U20406 ( .A(n459), .B(n20590), .Z(n20589) );
  XOR U20407 ( .A(p_input[1336]), .B(p_input[1304]), .Z(n20590) );
  XOR U20408 ( .A(n20591), .B(n20592), .Z(n20582) );
  AND U20409 ( .A(n20593), .B(n20594), .Z(n20592) );
  XOR U20410 ( .A(n20591), .B(n19719), .Z(n20594) );
  XNOR U20411 ( .A(p_input[1367]), .B(n20595), .Z(n19719) );
  AND U20412 ( .A(n462), .B(n20596), .Z(n20595) );
  XOR U20413 ( .A(p_input[1399]), .B(p_input[1367]), .Z(n20596) );
  XNOR U20414 ( .A(n19716), .B(n20591), .Z(n20593) );
  XOR U20415 ( .A(n20597), .B(n20598), .Z(n19716) );
  AND U20416 ( .A(n459), .B(n20599), .Z(n20598) );
  XOR U20417 ( .A(p_input[1335]), .B(p_input[1303]), .Z(n20599) );
  XOR U20418 ( .A(n20600), .B(n20601), .Z(n20591) );
  AND U20419 ( .A(n20602), .B(n20603), .Z(n20601) );
  XOR U20420 ( .A(n20600), .B(n19731), .Z(n20603) );
  XNOR U20421 ( .A(p_input[1366]), .B(n20604), .Z(n19731) );
  AND U20422 ( .A(n462), .B(n20605), .Z(n20604) );
  XOR U20423 ( .A(p_input[1398]), .B(p_input[1366]), .Z(n20605) );
  XNOR U20424 ( .A(n19728), .B(n20600), .Z(n20602) );
  XOR U20425 ( .A(n20606), .B(n20607), .Z(n19728) );
  AND U20426 ( .A(n459), .B(n20608), .Z(n20607) );
  XOR U20427 ( .A(p_input[1334]), .B(p_input[1302]), .Z(n20608) );
  XOR U20428 ( .A(n20609), .B(n20610), .Z(n20600) );
  AND U20429 ( .A(n20611), .B(n20612), .Z(n20610) );
  XOR U20430 ( .A(n20609), .B(n19743), .Z(n20612) );
  XNOR U20431 ( .A(p_input[1365]), .B(n20613), .Z(n19743) );
  AND U20432 ( .A(n462), .B(n20614), .Z(n20613) );
  XOR U20433 ( .A(p_input[1397]), .B(p_input[1365]), .Z(n20614) );
  XNOR U20434 ( .A(n19740), .B(n20609), .Z(n20611) );
  XOR U20435 ( .A(n20615), .B(n20616), .Z(n19740) );
  AND U20436 ( .A(n459), .B(n20617), .Z(n20616) );
  XOR U20437 ( .A(p_input[1333]), .B(p_input[1301]), .Z(n20617) );
  XOR U20438 ( .A(n20618), .B(n20619), .Z(n20609) );
  AND U20439 ( .A(n20620), .B(n20621), .Z(n20619) );
  XOR U20440 ( .A(n20618), .B(n19755), .Z(n20621) );
  XNOR U20441 ( .A(p_input[1364]), .B(n20622), .Z(n19755) );
  AND U20442 ( .A(n462), .B(n20623), .Z(n20622) );
  XOR U20443 ( .A(p_input[1396]), .B(p_input[1364]), .Z(n20623) );
  XNOR U20444 ( .A(n19752), .B(n20618), .Z(n20620) );
  XOR U20445 ( .A(n20624), .B(n20625), .Z(n19752) );
  AND U20446 ( .A(n459), .B(n20626), .Z(n20625) );
  XOR U20447 ( .A(p_input[1332]), .B(p_input[1300]), .Z(n20626) );
  XOR U20448 ( .A(n20627), .B(n20628), .Z(n20618) );
  AND U20449 ( .A(n20629), .B(n20630), .Z(n20628) );
  XOR U20450 ( .A(n20627), .B(n19767), .Z(n20630) );
  XNOR U20451 ( .A(p_input[1363]), .B(n20631), .Z(n19767) );
  AND U20452 ( .A(n462), .B(n20632), .Z(n20631) );
  XOR U20453 ( .A(p_input[1395]), .B(p_input[1363]), .Z(n20632) );
  XNOR U20454 ( .A(n19764), .B(n20627), .Z(n20629) );
  XOR U20455 ( .A(n20633), .B(n20634), .Z(n19764) );
  AND U20456 ( .A(n459), .B(n20635), .Z(n20634) );
  XOR U20457 ( .A(p_input[1331]), .B(p_input[1299]), .Z(n20635) );
  XOR U20458 ( .A(n20636), .B(n20637), .Z(n20627) );
  AND U20459 ( .A(n20638), .B(n20639), .Z(n20637) );
  XOR U20460 ( .A(n20636), .B(n19779), .Z(n20639) );
  XNOR U20461 ( .A(p_input[1362]), .B(n20640), .Z(n19779) );
  AND U20462 ( .A(n462), .B(n20641), .Z(n20640) );
  XOR U20463 ( .A(p_input[1394]), .B(p_input[1362]), .Z(n20641) );
  XNOR U20464 ( .A(n19776), .B(n20636), .Z(n20638) );
  XOR U20465 ( .A(n20642), .B(n20643), .Z(n19776) );
  AND U20466 ( .A(n459), .B(n20644), .Z(n20643) );
  XOR U20467 ( .A(p_input[1330]), .B(p_input[1298]), .Z(n20644) );
  XOR U20468 ( .A(n20645), .B(n20646), .Z(n20636) );
  AND U20469 ( .A(n20647), .B(n20648), .Z(n20646) );
  XOR U20470 ( .A(n20645), .B(n19791), .Z(n20648) );
  XNOR U20471 ( .A(p_input[1361]), .B(n20649), .Z(n19791) );
  AND U20472 ( .A(n462), .B(n20650), .Z(n20649) );
  XOR U20473 ( .A(p_input[1393]), .B(p_input[1361]), .Z(n20650) );
  XNOR U20474 ( .A(n19788), .B(n20645), .Z(n20647) );
  XOR U20475 ( .A(n20651), .B(n20652), .Z(n19788) );
  AND U20476 ( .A(n459), .B(n20653), .Z(n20652) );
  XOR U20477 ( .A(p_input[1329]), .B(p_input[1297]), .Z(n20653) );
  XOR U20478 ( .A(n20654), .B(n20655), .Z(n20645) );
  AND U20479 ( .A(n20656), .B(n20657), .Z(n20655) );
  XOR U20480 ( .A(n20654), .B(n19803), .Z(n20657) );
  XNOR U20481 ( .A(p_input[1360]), .B(n20658), .Z(n19803) );
  AND U20482 ( .A(n462), .B(n20659), .Z(n20658) );
  XOR U20483 ( .A(p_input[1392]), .B(p_input[1360]), .Z(n20659) );
  XNOR U20484 ( .A(n19800), .B(n20654), .Z(n20656) );
  XOR U20485 ( .A(n20660), .B(n20661), .Z(n19800) );
  AND U20486 ( .A(n459), .B(n20662), .Z(n20661) );
  XOR U20487 ( .A(p_input[1328]), .B(p_input[1296]), .Z(n20662) );
  XOR U20488 ( .A(n20663), .B(n20664), .Z(n20654) );
  AND U20489 ( .A(n20665), .B(n20666), .Z(n20664) );
  XOR U20490 ( .A(n20663), .B(n19815), .Z(n20666) );
  XNOR U20491 ( .A(p_input[1359]), .B(n20667), .Z(n19815) );
  AND U20492 ( .A(n462), .B(n20668), .Z(n20667) );
  XOR U20493 ( .A(p_input[1391]), .B(p_input[1359]), .Z(n20668) );
  XNOR U20494 ( .A(n19812), .B(n20663), .Z(n20665) );
  XOR U20495 ( .A(n20669), .B(n20670), .Z(n19812) );
  AND U20496 ( .A(n459), .B(n20671), .Z(n20670) );
  XOR U20497 ( .A(p_input[1327]), .B(p_input[1295]), .Z(n20671) );
  XOR U20498 ( .A(n20672), .B(n20673), .Z(n20663) );
  AND U20499 ( .A(n20674), .B(n20675), .Z(n20673) );
  XOR U20500 ( .A(n20672), .B(n19827), .Z(n20675) );
  XNOR U20501 ( .A(p_input[1358]), .B(n20676), .Z(n19827) );
  AND U20502 ( .A(n462), .B(n20677), .Z(n20676) );
  XOR U20503 ( .A(p_input[1390]), .B(p_input[1358]), .Z(n20677) );
  XNOR U20504 ( .A(n19824), .B(n20672), .Z(n20674) );
  XOR U20505 ( .A(n20678), .B(n20679), .Z(n19824) );
  AND U20506 ( .A(n459), .B(n20680), .Z(n20679) );
  XOR U20507 ( .A(p_input[1326]), .B(p_input[1294]), .Z(n20680) );
  XOR U20508 ( .A(n20681), .B(n20682), .Z(n20672) );
  AND U20509 ( .A(n20683), .B(n20684), .Z(n20682) );
  XOR U20510 ( .A(n20681), .B(n19839), .Z(n20684) );
  XNOR U20511 ( .A(p_input[1357]), .B(n20685), .Z(n19839) );
  AND U20512 ( .A(n462), .B(n20686), .Z(n20685) );
  XOR U20513 ( .A(p_input[1389]), .B(p_input[1357]), .Z(n20686) );
  XNOR U20514 ( .A(n19836), .B(n20681), .Z(n20683) );
  XOR U20515 ( .A(n20687), .B(n20688), .Z(n19836) );
  AND U20516 ( .A(n459), .B(n20689), .Z(n20688) );
  XOR U20517 ( .A(p_input[1325]), .B(p_input[1293]), .Z(n20689) );
  XOR U20518 ( .A(n20690), .B(n20691), .Z(n20681) );
  AND U20519 ( .A(n20692), .B(n20693), .Z(n20691) );
  XOR U20520 ( .A(n20690), .B(n19851), .Z(n20693) );
  XNOR U20521 ( .A(p_input[1356]), .B(n20694), .Z(n19851) );
  AND U20522 ( .A(n462), .B(n20695), .Z(n20694) );
  XOR U20523 ( .A(p_input[1388]), .B(p_input[1356]), .Z(n20695) );
  XNOR U20524 ( .A(n19848), .B(n20690), .Z(n20692) );
  XOR U20525 ( .A(n20696), .B(n20697), .Z(n19848) );
  AND U20526 ( .A(n459), .B(n20698), .Z(n20697) );
  XOR U20527 ( .A(p_input[1324]), .B(p_input[1292]), .Z(n20698) );
  XOR U20528 ( .A(n20699), .B(n20700), .Z(n20690) );
  AND U20529 ( .A(n20701), .B(n20702), .Z(n20700) );
  XOR U20530 ( .A(n20699), .B(n19863), .Z(n20702) );
  XNOR U20531 ( .A(p_input[1355]), .B(n20703), .Z(n19863) );
  AND U20532 ( .A(n462), .B(n20704), .Z(n20703) );
  XOR U20533 ( .A(p_input[1387]), .B(p_input[1355]), .Z(n20704) );
  XNOR U20534 ( .A(n19860), .B(n20699), .Z(n20701) );
  XOR U20535 ( .A(n20705), .B(n20706), .Z(n19860) );
  AND U20536 ( .A(n459), .B(n20707), .Z(n20706) );
  XOR U20537 ( .A(p_input[1323]), .B(p_input[1291]), .Z(n20707) );
  XOR U20538 ( .A(n20708), .B(n20709), .Z(n20699) );
  AND U20539 ( .A(n20710), .B(n20711), .Z(n20709) );
  XOR U20540 ( .A(n20708), .B(n19875), .Z(n20711) );
  XNOR U20541 ( .A(p_input[1354]), .B(n20712), .Z(n19875) );
  AND U20542 ( .A(n462), .B(n20713), .Z(n20712) );
  XOR U20543 ( .A(p_input[1386]), .B(p_input[1354]), .Z(n20713) );
  XNOR U20544 ( .A(n19872), .B(n20708), .Z(n20710) );
  XOR U20545 ( .A(n20714), .B(n20715), .Z(n19872) );
  AND U20546 ( .A(n459), .B(n20716), .Z(n20715) );
  XOR U20547 ( .A(p_input[1322]), .B(p_input[1290]), .Z(n20716) );
  XOR U20548 ( .A(n20717), .B(n20718), .Z(n20708) );
  AND U20549 ( .A(n20719), .B(n20720), .Z(n20718) );
  XOR U20550 ( .A(n20717), .B(n19887), .Z(n20720) );
  XNOR U20551 ( .A(p_input[1353]), .B(n20721), .Z(n19887) );
  AND U20552 ( .A(n462), .B(n20722), .Z(n20721) );
  XOR U20553 ( .A(p_input[1385]), .B(p_input[1353]), .Z(n20722) );
  XNOR U20554 ( .A(n19884), .B(n20717), .Z(n20719) );
  XOR U20555 ( .A(n20723), .B(n20724), .Z(n19884) );
  AND U20556 ( .A(n459), .B(n20725), .Z(n20724) );
  XOR U20557 ( .A(p_input[1321]), .B(p_input[1289]), .Z(n20725) );
  XOR U20558 ( .A(n20726), .B(n20727), .Z(n20717) );
  AND U20559 ( .A(n20728), .B(n20729), .Z(n20727) );
  XOR U20560 ( .A(n20726), .B(n19899), .Z(n20729) );
  XNOR U20561 ( .A(p_input[1352]), .B(n20730), .Z(n19899) );
  AND U20562 ( .A(n462), .B(n20731), .Z(n20730) );
  XOR U20563 ( .A(p_input[1384]), .B(p_input[1352]), .Z(n20731) );
  XNOR U20564 ( .A(n19896), .B(n20726), .Z(n20728) );
  XOR U20565 ( .A(n20732), .B(n20733), .Z(n19896) );
  AND U20566 ( .A(n459), .B(n20734), .Z(n20733) );
  XOR U20567 ( .A(p_input[1320]), .B(p_input[1288]), .Z(n20734) );
  XOR U20568 ( .A(n20735), .B(n20736), .Z(n20726) );
  AND U20569 ( .A(n20737), .B(n20738), .Z(n20736) );
  XOR U20570 ( .A(n20735), .B(n19911), .Z(n20738) );
  XNOR U20571 ( .A(p_input[1351]), .B(n20739), .Z(n19911) );
  AND U20572 ( .A(n462), .B(n20740), .Z(n20739) );
  XOR U20573 ( .A(p_input[1383]), .B(p_input[1351]), .Z(n20740) );
  XNOR U20574 ( .A(n19908), .B(n20735), .Z(n20737) );
  XOR U20575 ( .A(n20741), .B(n20742), .Z(n19908) );
  AND U20576 ( .A(n459), .B(n20743), .Z(n20742) );
  XOR U20577 ( .A(p_input[1319]), .B(p_input[1287]), .Z(n20743) );
  XOR U20578 ( .A(n20744), .B(n20745), .Z(n20735) );
  AND U20579 ( .A(n20746), .B(n20747), .Z(n20745) );
  XOR U20580 ( .A(n20744), .B(n19923), .Z(n20747) );
  XNOR U20581 ( .A(p_input[1350]), .B(n20748), .Z(n19923) );
  AND U20582 ( .A(n462), .B(n20749), .Z(n20748) );
  XOR U20583 ( .A(p_input[1382]), .B(p_input[1350]), .Z(n20749) );
  XNOR U20584 ( .A(n19920), .B(n20744), .Z(n20746) );
  XOR U20585 ( .A(n20750), .B(n20751), .Z(n19920) );
  AND U20586 ( .A(n459), .B(n20752), .Z(n20751) );
  XOR U20587 ( .A(p_input[1318]), .B(p_input[1286]), .Z(n20752) );
  XOR U20588 ( .A(n20753), .B(n20754), .Z(n20744) );
  AND U20589 ( .A(n20755), .B(n20756), .Z(n20754) );
  XOR U20590 ( .A(n20753), .B(n19935), .Z(n20756) );
  XNOR U20591 ( .A(p_input[1349]), .B(n20757), .Z(n19935) );
  AND U20592 ( .A(n462), .B(n20758), .Z(n20757) );
  XOR U20593 ( .A(p_input[1381]), .B(p_input[1349]), .Z(n20758) );
  XNOR U20594 ( .A(n19932), .B(n20753), .Z(n20755) );
  XOR U20595 ( .A(n20759), .B(n20760), .Z(n19932) );
  AND U20596 ( .A(n459), .B(n20761), .Z(n20760) );
  XOR U20597 ( .A(p_input[1317]), .B(p_input[1285]), .Z(n20761) );
  XOR U20598 ( .A(n20762), .B(n20763), .Z(n20753) );
  AND U20599 ( .A(n20764), .B(n20765), .Z(n20763) );
  XOR U20600 ( .A(n20762), .B(n19947), .Z(n20765) );
  XNOR U20601 ( .A(p_input[1348]), .B(n20766), .Z(n19947) );
  AND U20602 ( .A(n462), .B(n20767), .Z(n20766) );
  XOR U20603 ( .A(p_input[1380]), .B(p_input[1348]), .Z(n20767) );
  XNOR U20604 ( .A(n19944), .B(n20762), .Z(n20764) );
  XOR U20605 ( .A(n20768), .B(n20769), .Z(n19944) );
  AND U20606 ( .A(n459), .B(n20770), .Z(n20769) );
  XOR U20607 ( .A(p_input[1316]), .B(p_input[1284]), .Z(n20770) );
  XOR U20608 ( .A(n20771), .B(n20772), .Z(n20762) );
  AND U20609 ( .A(n20773), .B(n20774), .Z(n20772) );
  XOR U20610 ( .A(n20771), .B(n19959), .Z(n20774) );
  XNOR U20611 ( .A(p_input[1347]), .B(n20775), .Z(n19959) );
  AND U20612 ( .A(n462), .B(n20776), .Z(n20775) );
  XOR U20613 ( .A(p_input[1379]), .B(p_input[1347]), .Z(n20776) );
  XNOR U20614 ( .A(n19956), .B(n20771), .Z(n20773) );
  XOR U20615 ( .A(n20777), .B(n20778), .Z(n19956) );
  AND U20616 ( .A(n459), .B(n20779), .Z(n20778) );
  XOR U20617 ( .A(p_input[1315]), .B(p_input[1283]), .Z(n20779) );
  XOR U20618 ( .A(n20780), .B(n20781), .Z(n20771) );
  AND U20619 ( .A(n20782), .B(n20783), .Z(n20781) );
  XOR U20620 ( .A(n19971), .B(n20780), .Z(n20783) );
  XNOR U20621 ( .A(p_input[1346]), .B(n20784), .Z(n19971) );
  AND U20622 ( .A(n462), .B(n20785), .Z(n20784) );
  XOR U20623 ( .A(p_input[1378]), .B(p_input[1346]), .Z(n20785) );
  XNOR U20624 ( .A(n20780), .B(n19968), .Z(n20782) );
  XOR U20625 ( .A(n20786), .B(n20787), .Z(n19968) );
  AND U20626 ( .A(n459), .B(n20788), .Z(n20787) );
  XOR U20627 ( .A(p_input[1314]), .B(p_input[1282]), .Z(n20788) );
  XOR U20628 ( .A(n20789), .B(n20790), .Z(n20780) );
  AND U20629 ( .A(n20791), .B(n20792), .Z(n20790) );
  XNOR U20630 ( .A(n20793), .B(n19984), .Z(n20792) );
  XNOR U20631 ( .A(p_input[1345]), .B(n20794), .Z(n19984) );
  AND U20632 ( .A(n462), .B(n20795), .Z(n20794) );
  XNOR U20633 ( .A(p_input[1377]), .B(n20796), .Z(n20795) );
  IV U20634 ( .A(p_input[1345]), .Z(n20796) );
  XNOR U20635 ( .A(n19981), .B(n20789), .Z(n20791) );
  XNOR U20636 ( .A(p_input[1281]), .B(n20797), .Z(n19981) );
  AND U20637 ( .A(n459), .B(n20798), .Z(n20797) );
  XOR U20638 ( .A(p_input[1313]), .B(p_input[1281]), .Z(n20798) );
  IV U20639 ( .A(n20793), .Z(n20789) );
  AND U20640 ( .A(n20519), .B(n20522), .Z(n20793) );
  XOR U20641 ( .A(p_input[1344]), .B(n20799), .Z(n20522) );
  AND U20642 ( .A(n462), .B(n20800), .Z(n20799) );
  XOR U20643 ( .A(p_input[1376]), .B(p_input[1344]), .Z(n20800) );
  XOR U20644 ( .A(n20801), .B(n20802), .Z(n462) );
  AND U20645 ( .A(n20803), .B(n20804), .Z(n20802) );
  XNOR U20646 ( .A(p_input[1407]), .B(n20801), .Z(n20804) );
  XOR U20647 ( .A(n20801), .B(p_input[1375]), .Z(n20803) );
  XOR U20648 ( .A(n20805), .B(n20806), .Z(n20801) );
  AND U20649 ( .A(n20807), .B(n20808), .Z(n20806) );
  XNOR U20650 ( .A(p_input[1406]), .B(n20805), .Z(n20808) );
  XOR U20651 ( .A(n20805), .B(p_input[1374]), .Z(n20807) );
  XOR U20652 ( .A(n20809), .B(n20810), .Z(n20805) );
  AND U20653 ( .A(n20811), .B(n20812), .Z(n20810) );
  XNOR U20654 ( .A(p_input[1405]), .B(n20809), .Z(n20812) );
  XOR U20655 ( .A(n20809), .B(p_input[1373]), .Z(n20811) );
  XOR U20656 ( .A(n20813), .B(n20814), .Z(n20809) );
  AND U20657 ( .A(n20815), .B(n20816), .Z(n20814) );
  XNOR U20658 ( .A(p_input[1404]), .B(n20813), .Z(n20816) );
  XOR U20659 ( .A(n20813), .B(p_input[1372]), .Z(n20815) );
  XOR U20660 ( .A(n20817), .B(n20818), .Z(n20813) );
  AND U20661 ( .A(n20819), .B(n20820), .Z(n20818) );
  XNOR U20662 ( .A(p_input[1403]), .B(n20817), .Z(n20820) );
  XOR U20663 ( .A(n20817), .B(p_input[1371]), .Z(n20819) );
  XOR U20664 ( .A(n20821), .B(n20822), .Z(n20817) );
  AND U20665 ( .A(n20823), .B(n20824), .Z(n20822) );
  XNOR U20666 ( .A(p_input[1402]), .B(n20821), .Z(n20824) );
  XOR U20667 ( .A(n20821), .B(p_input[1370]), .Z(n20823) );
  XOR U20668 ( .A(n20825), .B(n20826), .Z(n20821) );
  AND U20669 ( .A(n20827), .B(n20828), .Z(n20826) );
  XNOR U20670 ( .A(p_input[1401]), .B(n20825), .Z(n20828) );
  XOR U20671 ( .A(n20825), .B(p_input[1369]), .Z(n20827) );
  XOR U20672 ( .A(n20829), .B(n20830), .Z(n20825) );
  AND U20673 ( .A(n20831), .B(n20832), .Z(n20830) );
  XNOR U20674 ( .A(p_input[1400]), .B(n20829), .Z(n20832) );
  XOR U20675 ( .A(n20829), .B(p_input[1368]), .Z(n20831) );
  XOR U20676 ( .A(n20833), .B(n20834), .Z(n20829) );
  AND U20677 ( .A(n20835), .B(n20836), .Z(n20834) );
  XNOR U20678 ( .A(p_input[1399]), .B(n20833), .Z(n20836) );
  XOR U20679 ( .A(n20833), .B(p_input[1367]), .Z(n20835) );
  XOR U20680 ( .A(n20837), .B(n20838), .Z(n20833) );
  AND U20681 ( .A(n20839), .B(n20840), .Z(n20838) );
  XNOR U20682 ( .A(p_input[1398]), .B(n20837), .Z(n20840) );
  XOR U20683 ( .A(n20837), .B(p_input[1366]), .Z(n20839) );
  XOR U20684 ( .A(n20841), .B(n20842), .Z(n20837) );
  AND U20685 ( .A(n20843), .B(n20844), .Z(n20842) );
  XNOR U20686 ( .A(p_input[1397]), .B(n20841), .Z(n20844) );
  XOR U20687 ( .A(n20841), .B(p_input[1365]), .Z(n20843) );
  XOR U20688 ( .A(n20845), .B(n20846), .Z(n20841) );
  AND U20689 ( .A(n20847), .B(n20848), .Z(n20846) );
  XNOR U20690 ( .A(p_input[1396]), .B(n20845), .Z(n20848) );
  XOR U20691 ( .A(n20845), .B(p_input[1364]), .Z(n20847) );
  XOR U20692 ( .A(n20849), .B(n20850), .Z(n20845) );
  AND U20693 ( .A(n20851), .B(n20852), .Z(n20850) );
  XNOR U20694 ( .A(p_input[1395]), .B(n20849), .Z(n20852) );
  XOR U20695 ( .A(n20849), .B(p_input[1363]), .Z(n20851) );
  XOR U20696 ( .A(n20853), .B(n20854), .Z(n20849) );
  AND U20697 ( .A(n20855), .B(n20856), .Z(n20854) );
  XNOR U20698 ( .A(p_input[1394]), .B(n20853), .Z(n20856) );
  XOR U20699 ( .A(n20853), .B(p_input[1362]), .Z(n20855) );
  XOR U20700 ( .A(n20857), .B(n20858), .Z(n20853) );
  AND U20701 ( .A(n20859), .B(n20860), .Z(n20858) );
  XNOR U20702 ( .A(p_input[1393]), .B(n20857), .Z(n20860) );
  XOR U20703 ( .A(n20857), .B(p_input[1361]), .Z(n20859) );
  XOR U20704 ( .A(n20861), .B(n20862), .Z(n20857) );
  AND U20705 ( .A(n20863), .B(n20864), .Z(n20862) );
  XNOR U20706 ( .A(p_input[1392]), .B(n20861), .Z(n20864) );
  XOR U20707 ( .A(n20861), .B(p_input[1360]), .Z(n20863) );
  XOR U20708 ( .A(n20865), .B(n20866), .Z(n20861) );
  AND U20709 ( .A(n20867), .B(n20868), .Z(n20866) );
  XNOR U20710 ( .A(p_input[1391]), .B(n20865), .Z(n20868) );
  XOR U20711 ( .A(n20865), .B(p_input[1359]), .Z(n20867) );
  XOR U20712 ( .A(n20869), .B(n20870), .Z(n20865) );
  AND U20713 ( .A(n20871), .B(n20872), .Z(n20870) );
  XNOR U20714 ( .A(p_input[1390]), .B(n20869), .Z(n20872) );
  XOR U20715 ( .A(n20869), .B(p_input[1358]), .Z(n20871) );
  XOR U20716 ( .A(n20873), .B(n20874), .Z(n20869) );
  AND U20717 ( .A(n20875), .B(n20876), .Z(n20874) );
  XNOR U20718 ( .A(p_input[1389]), .B(n20873), .Z(n20876) );
  XOR U20719 ( .A(n20873), .B(p_input[1357]), .Z(n20875) );
  XOR U20720 ( .A(n20877), .B(n20878), .Z(n20873) );
  AND U20721 ( .A(n20879), .B(n20880), .Z(n20878) );
  XNOR U20722 ( .A(p_input[1388]), .B(n20877), .Z(n20880) );
  XOR U20723 ( .A(n20877), .B(p_input[1356]), .Z(n20879) );
  XOR U20724 ( .A(n20881), .B(n20882), .Z(n20877) );
  AND U20725 ( .A(n20883), .B(n20884), .Z(n20882) );
  XNOR U20726 ( .A(p_input[1387]), .B(n20881), .Z(n20884) );
  XOR U20727 ( .A(n20881), .B(p_input[1355]), .Z(n20883) );
  XOR U20728 ( .A(n20885), .B(n20886), .Z(n20881) );
  AND U20729 ( .A(n20887), .B(n20888), .Z(n20886) );
  XNOR U20730 ( .A(p_input[1386]), .B(n20885), .Z(n20888) );
  XOR U20731 ( .A(n20885), .B(p_input[1354]), .Z(n20887) );
  XOR U20732 ( .A(n20889), .B(n20890), .Z(n20885) );
  AND U20733 ( .A(n20891), .B(n20892), .Z(n20890) );
  XNOR U20734 ( .A(p_input[1385]), .B(n20889), .Z(n20892) );
  XOR U20735 ( .A(n20889), .B(p_input[1353]), .Z(n20891) );
  XOR U20736 ( .A(n20893), .B(n20894), .Z(n20889) );
  AND U20737 ( .A(n20895), .B(n20896), .Z(n20894) );
  XNOR U20738 ( .A(p_input[1384]), .B(n20893), .Z(n20896) );
  XOR U20739 ( .A(n20893), .B(p_input[1352]), .Z(n20895) );
  XOR U20740 ( .A(n20897), .B(n20898), .Z(n20893) );
  AND U20741 ( .A(n20899), .B(n20900), .Z(n20898) );
  XNOR U20742 ( .A(p_input[1383]), .B(n20897), .Z(n20900) );
  XOR U20743 ( .A(n20897), .B(p_input[1351]), .Z(n20899) );
  XOR U20744 ( .A(n20901), .B(n20902), .Z(n20897) );
  AND U20745 ( .A(n20903), .B(n20904), .Z(n20902) );
  XNOR U20746 ( .A(p_input[1382]), .B(n20901), .Z(n20904) );
  XOR U20747 ( .A(n20901), .B(p_input[1350]), .Z(n20903) );
  XOR U20748 ( .A(n20905), .B(n20906), .Z(n20901) );
  AND U20749 ( .A(n20907), .B(n20908), .Z(n20906) );
  XNOR U20750 ( .A(p_input[1381]), .B(n20905), .Z(n20908) );
  XOR U20751 ( .A(n20905), .B(p_input[1349]), .Z(n20907) );
  XOR U20752 ( .A(n20909), .B(n20910), .Z(n20905) );
  AND U20753 ( .A(n20911), .B(n20912), .Z(n20910) );
  XNOR U20754 ( .A(p_input[1380]), .B(n20909), .Z(n20912) );
  XOR U20755 ( .A(n20909), .B(p_input[1348]), .Z(n20911) );
  XOR U20756 ( .A(n20913), .B(n20914), .Z(n20909) );
  AND U20757 ( .A(n20915), .B(n20916), .Z(n20914) );
  XNOR U20758 ( .A(p_input[1379]), .B(n20913), .Z(n20916) );
  XOR U20759 ( .A(n20913), .B(p_input[1347]), .Z(n20915) );
  XOR U20760 ( .A(n20917), .B(n20918), .Z(n20913) );
  AND U20761 ( .A(n20919), .B(n20920), .Z(n20918) );
  XNOR U20762 ( .A(p_input[1378]), .B(n20917), .Z(n20920) );
  XOR U20763 ( .A(n20917), .B(p_input[1346]), .Z(n20919) );
  XNOR U20764 ( .A(n20921), .B(n20922), .Z(n20917) );
  AND U20765 ( .A(n20923), .B(n20924), .Z(n20922) );
  XOR U20766 ( .A(p_input[1377]), .B(n20921), .Z(n20924) );
  XNOR U20767 ( .A(p_input[1345]), .B(n20921), .Z(n20923) );
  AND U20768 ( .A(p_input[1376]), .B(n20925), .Z(n20921) );
  IV U20769 ( .A(p_input[1344]), .Z(n20925) );
  XNOR U20770 ( .A(p_input[1280]), .B(n20926), .Z(n20519) );
  AND U20771 ( .A(n459), .B(n20927), .Z(n20926) );
  XOR U20772 ( .A(p_input[1312]), .B(p_input[1280]), .Z(n20927) );
  XOR U20773 ( .A(n20928), .B(n20929), .Z(n459) );
  AND U20774 ( .A(n20930), .B(n20931), .Z(n20929) );
  XNOR U20775 ( .A(p_input[1343]), .B(n20928), .Z(n20931) );
  XOR U20776 ( .A(n20928), .B(p_input[1311]), .Z(n20930) );
  XOR U20777 ( .A(n20932), .B(n20933), .Z(n20928) );
  AND U20778 ( .A(n20934), .B(n20935), .Z(n20933) );
  XNOR U20779 ( .A(p_input[1342]), .B(n20932), .Z(n20935) );
  XNOR U20780 ( .A(n20932), .B(n20534), .Z(n20934) );
  IV U20781 ( .A(p_input[1310]), .Z(n20534) );
  XOR U20782 ( .A(n20936), .B(n20937), .Z(n20932) );
  AND U20783 ( .A(n20938), .B(n20939), .Z(n20937) );
  XNOR U20784 ( .A(p_input[1341]), .B(n20936), .Z(n20939) );
  XNOR U20785 ( .A(n20936), .B(n20543), .Z(n20938) );
  IV U20786 ( .A(p_input[1309]), .Z(n20543) );
  XOR U20787 ( .A(n20940), .B(n20941), .Z(n20936) );
  AND U20788 ( .A(n20942), .B(n20943), .Z(n20941) );
  XNOR U20789 ( .A(p_input[1340]), .B(n20940), .Z(n20943) );
  XNOR U20790 ( .A(n20940), .B(n20552), .Z(n20942) );
  IV U20791 ( .A(p_input[1308]), .Z(n20552) );
  XOR U20792 ( .A(n20944), .B(n20945), .Z(n20940) );
  AND U20793 ( .A(n20946), .B(n20947), .Z(n20945) );
  XNOR U20794 ( .A(p_input[1339]), .B(n20944), .Z(n20947) );
  XNOR U20795 ( .A(n20944), .B(n20561), .Z(n20946) );
  IV U20796 ( .A(p_input[1307]), .Z(n20561) );
  XOR U20797 ( .A(n20948), .B(n20949), .Z(n20944) );
  AND U20798 ( .A(n20950), .B(n20951), .Z(n20949) );
  XNOR U20799 ( .A(p_input[1338]), .B(n20948), .Z(n20951) );
  XNOR U20800 ( .A(n20948), .B(n20570), .Z(n20950) );
  IV U20801 ( .A(p_input[1306]), .Z(n20570) );
  XOR U20802 ( .A(n20952), .B(n20953), .Z(n20948) );
  AND U20803 ( .A(n20954), .B(n20955), .Z(n20953) );
  XNOR U20804 ( .A(p_input[1337]), .B(n20952), .Z(n20955) );
  XNOR U20805 ( .A(n20952), .B(n20579), .Z(n20954) );
  IV U20806 ( .A(p_input[1305]), .Z(n20579) );
  XOR U20807 ( .A(n20956), .B(n20957), .Z(n20952) );
  AND U20808 ( .A(n20958), .B(n20959), .Z(n20957) );
  XNOR U20809 ( .A(p_input[1336]), .B(n20956), .Z(n20959) );
  XNOR U20810 ( .A(n20956), .B(n20588), .Z(n20958) );
  IV U20811 ( .A(p_input[1304]), .Z(n20588) );
  XOR U20812 ( .A(n20960), .B(n20961), .Z(n20956) );
  AND U20813 ( .A(n20962), .B(n20963), .Z(n20961) );
  XNOR U20814 ( .A(p_input[1335]), .B(n20960), .Z(n20963) );
  XNOR U20815 ( .A(n20960), .B(n20597), .Z(n20962) );
  IV U20816 ( .A(p_input[1303]), .Z(n20597) );
  XOR U20817 ( .A(n20964), .B(n20965), .Z(n20960) );
  AND U20818 ( .A(n20966), .B(n20967), .Z(n20965) );
  XNOR U20819 ( .A(p_input[1334]), .B(n20964), .Z(n20967) );
  XNOR U20820 ( .A(n20964), .B(n20606), .Z(n20966) );
  IV U20821 ( .A(p_input[1302]), .Z(n20606) );
  XOR U20822 ( .A(n20968), .B(n20969), .Z(n20964) );
  AND U20823 ( .A(n20970), .B(n20971), .Z(n20969) );
  XNOR U20824 ( .A(p_input[1333]), .B(n20968), .Z(n20971) );
  XNOR U20825 ( .A(n20968), .B(n20615), .Z(n20970) );
  IV U20826 ( .A(p_input[1301]), .Z(n20615) );
  XOR U20827 ( .A(n20972), .B(n20973), .Z(n20968) );
  AND U20828 ( .A(n20974), .B(n20975), .Z(n20973) );
  XNOR U20829 ( .A(p_input[1332]), .B(n20972), .Z(n20975) );
  XNOR U20830 ( .A(n20972), .B(n20624), .Z(n20974) );
  IV U20831 ( .A(p_input[1300]), .Z(n20624) );
  XOR U20832 ( .A(n20976), .B(n20977), .Z(n20972) );
  AND U20833 ( .A(n20978), .B(n20979), .Z(n20977) );
  XNOR U20834 ( .A(p_input[1331]), .B(n20976), .Z(n20979) );
  XNOR U20835 ( .A(n20976), .B(n20633), .Z(n20978) );
  IV U20836 ( .A(p_input[1299]), .Z(n20633) );
  XOR U20837 ( .A(n20980), .B(n20981), .Z(n20976) );
  AND U20838 ( .A(n20982), .B(n20983), .Z(n20981) );
  XNOR U20839 ( .A(p_input[1330]), .B(n20980), .Z(n20983) );
  XNOR U20840 ( .A(n20980), .B(n20642), .Z(n20982) );
  IV U20841 ( .A(p_input[1298]), .Z(n20642) );
  XOR U20842 ( .A(n20984), .B(n20985), .Z(n20980) );
  AND U20843 ( .A(n20986), .B(n20987), .Z(n20985) );
  XNOR U20844 ( .A(p_input[1329]), .B(n20984), .Z(n20987) );
  XNOR U20845 ( .A(n20984), .B(n20651), .Z(n20986) );
  IV U20846 ( .A(p_input[1297]), .Z(n20651) );
  XOR U20847 ( .A(n20988), .B(n20989), .Z(n20984) );
  AND U20848 ( .A(n20990), .B(n20991), .Z(n20989) );
  XNOR U20849 ( .A(p_input[1328]), .B(n20988), .Z(n20991) );
  XNOR U20850 ( .A(n20988), .B(n20660), .Z(n20990) );
  IV U20851 ( .A(p_input[1296]), .Z(n20660) );
  XOR U20852 ( .A(n20992), .B(n20993), .Z(n20988) );
  AND U20853 ( .A(n20994), .B(n20995), .Z(n20993) );
  XNOR U20854 ( .A(p_input[1327]), .B(n20992), .Z(n20995) );
  XNOR U20855 ( .A(n20992), .B(n20669), .Z(n20994) );
  IV U20856 ( .A(p_input[1295]), .Z(n20669) );
  XOR U20857 ( .A(n20996), .B(n20997), .Z(n20992) );
  AND U20858 ( .A(n20998), .B(n20999), .Z(n20997) );
  XNOR U20859 ( .A(p_input[1326]), .B(n20996), .Z(n20999) );
  XNOR U20860 ( .A(n20996), .B(n20678), .Z(n20998) );
  IV U20861 ( .A(p_input[1294]), .Z(n20678) );
  XOR U20862 ( .A(n21000), .B(n21001), .Z(n20996) );
  AND U20863 ( .A(n21002), .B(n21003), .Z(n21001) );
  XNOR U20864 ( .A(p_input[1325]), .B(n21000), .Z(n21003) );
  XNOR U20865 ( .A(n21000), .B(n20687), .Z(n21002) );
  IV U20866 ( .A(p_input[1293]), .Z(n20687) );
  XOR U20867 ( .A(n21004), .B(n21005), .Z(n21000) );
  AND U20868 ( .A(n21006), .B(n21007), .Z(n21005) );
  XNOR U20869 ( .A(p_input[1324]), .B(n21004), .Z(n21007) );
  XNOR U20870 ( .A(n21004), .B(n20696), .Z(n21006) );
  IV U20871 ( .A(p_input[1292]), .Z(n20696) );
  XOR U20872 ( .A(n21008), .B(n21009), .Z(n21004) );
  AND U20873 ( .A(n21010), .B(n21011), .Z(n21009) );
  XNOR U20874 ( .A(p_input[1323]), .B(n21008), .Z(n21011) );
  XNOR U20875 ( .A(n21008), .B(n20705), .Z(n21010) );
  IV U20876 ( .A(p_input[1291]), .Z(n20705) );
  XOR U20877 ( .A(n21012), .B(n21013), .Z(n21008) );
  AND U20878 ( .A(n21014), .B(n21015), .Z(n21013) );
  XNOR U20879 ( .A(p_input[1322]), .B(n21012), .Z(n21015) );
  XNOR U20880 ( .A(n21012), .B(n20714), .Z(n21014) );
  IV U20881 ( .A(p_input[1290]), .Z(n20714) );
  XOR U20882 ( .A(n21016), .B(n21017), .Z(n21012) );
  AND U20883 ( .A(n21018), .B(n21019), .Z(n21017) );
  XNOR U20884 ( .A(p_input[1321]), .B(n21016), .Z(n21019) );
  XNOR U20885 ( .A(n21016), .B(n20723), .Z(n21018) );
  IV U20886 ( .A(p_input[1289]), .Z(n20723) );
  XOR U20887 ( .A(n21020), .B(n21021), .Z(n21016) );
  AND U20888 ( .A(n21022), .B(n21023), .Z(n21021) );
  XNOR U20889 ( .A(p_input[1320]), .B(n21020), .Z(n21023) );
  XNOR U20890 ( .A(n21020), .B(n20732), .Z(n21022) );
  IV U20891 ( .A(p_input[1288]), .Z(n20732) );
  XOR U20892 ( .A(n21024), .B(n21025), .Z(n21020) );
  AND U20893 ( .A(n21026), .B(n21027), .Z(n21025) );
  XNOR U20894 ( .A(p_input[1319]), .B(n21024), .Z(n21027) );
  XNOR U20895 ( .A(n21024), .B(n20741), .Z(n21026) );
  IV U20896 ( .A(p_input[1287]), .Z(n20741) );
  XOR U20897 ( .A(n21028), .B(n21029), .Z(n21024) );
  AND U20898 ( .A(n21030), .B(n21031), .Z(n21029) );
  XNOR U20899 ( .A(p_input[1318]), .B(n21028), .Z(n21031) );
  XNOR U20900 ( .A(n21028), .B(n20750), .Z(n21030) );
  IV U20901 ( .A(p_input[1286]), .Z(n20750) );
  XOR U20902 ( .A(n21032), .B(n21033), .Z(n21028) );
  AND U20903 ( .A(n21034), .B(n21035), .Z(n21033) );
  XNOR U20904 ( .A(p_input[1317]), .B(n21032), .Z(n21035) );
  XNOR U20905 ( .A(n21032), .B(n20759), .Z(n21034) );
  IV U20906 ( .A(p_input[1285]), .Z(n20759) );
  XOR U20907 ( .A(n21036), .B(n21037), .Z(n21032) );
  AND U20908 ( .A(n21038), .B(n21039), .Z(n21037) );
  XNOR U20909 ( .A(p_input[1316]), .B(n21036), .Z(n21039) );
  XNOR U20910 ( .A(n21036), .B(n20768), .Z(n21038) );
  IV U20911 ( .A(p_input[1284]), .Z(n20768) );
  XOR U20912 ( .A(n21040), .B(n21041), .Z(n21036) );
  AND U20913 ( .A(n21042), .B(n21043), .Z(n21041) );
  XNOR U20914 ( .A(p_input[1315]), .B(n21040), .Z(n21043) );
  XNOR U20915 ( .A(n21040), .B(n20777), .Z(n21042) );
  IV U20916 ( .A(p_input[1283]), .Z(n20777) );
  XOR U20917 ( .A(n21044), .B(n21045), .Z(n21040) );
  AND U20918 ( .A(n21046), .B(n21047), .Z(n21045) );
  XNOR U20919 ( .A(p_input[1314]), .B(n21044), .Z(n21047) );
  XNOR U20920 ( .A(n21044), .B(n20786), .Z(n21046) );
  IV U20921 ( .A(p_input[1282]), .Z(n20786) );
  XNOR U20922 ( .A(n21048), .B(n21049), .Z(n21044) );
  AND U20923 ( .A(n21050), .B(n21051), .Z(n21049) );
  XOR U20924 ( .A(p_input[1313]), .B(n21048), .Z(n21051) );
  XNOR U20925 ( .A(p_input[1281]), .B(n21048), .Z(n21050) );
  AND U20926 ( .A(p_input[1312]), .B(n21052), .Z(n21048) );
  IV U20927 ( .A(p_input[1280]), .Z(n21052) );
  XOR U20928 ( .A(n21053), .B(n21054), .Z(n19231) );
  AND U20929 ( .A(n519), .B(n21055), .Z(n21054) );
  XNOR U20930 ( .A(n21056), .B(n21053), .Z(n21055) );
  XOR U20931 ( .A(n21057), .B(n21058), .Z(n519) );
  AND U20932 ( .A(n21059), .B(n21060), .Z(n21058) );
  XOR U20933 ( .A(n21057), .B(n19246), .Z(n21060) );
  XNOR U20934 ( .A(n21061), .B(n21062), .Z(n19246) );
  AND U20935 ( .A(n21063), .B(n382), .Z(n21062) );
  AND U20936 ( .A(n21061), .B(n21064), .Z(n21063) );
  XNOR U20937 ( .A(n19243), .B(n21057), .Z(n21059) );
  XOR U20938 ( .A(n21065), .B(n21066), .Z(n19243) );
  AND U20939 ( .A(n21067), .B(n379), .Z(n21066) );
  NOR U20940 ( .A(n21065), .B(n21068), .Z(n21067) );
  XOR U20941 ( .A(n21069), .B(n21070), .Z(n21057) );
  AND U20942 ( .A(n21071), .B(n21072), .Z(n21070) );
  XOR U20943 ( .A(n21069), .B(n19258), .Z(n21072) );
  XOR U20944 ( .A(n21073), .B(n21074), .Z(n19258) );
  AND U20945 ( .A(n382), .B(n21075), .Z(n21074) );
  XOR U20946 ( .A(n21076), .B(n21073), .Z(n21075) );
  XNOR U20947 ( .A(n19255), .B(n21069), .Z(n21071) );
  XOR U20948 ( .A(n21077), .B(n21078), .Z(n19255) );
  AND U20949 ( .A(n379), .B(n21079), .Z(n21078) );
  XOR U20950 ( .A(n21080), .B(n21077), .Z(n21079) );
  XOR U20951 ( .A(n21081), .B(n21082), .Z(n21069) );
  AND U20952 ( .A(n21083), .B(n21084), .Z(n21082) );
  XOR U20953 ( .A(n21081), .B(n19270), .Z(n21084) );
  XOR U20954 ( .A(n21085), .B(n21086), .Z(n19270) );
  AND U20955 ( .A(n382), .B(n21087), .Z(n21086) );
  XOR U20956 ( .A(n21088), .B(n21085), .Z(n21087) );
  XNOR U20957 ( .A(n19267), .B(n21081), .Z(n21083) );
  XOR U20958 ( .A(n21089), .B(n21090), .Z(n19267) );
  AND U20959 ( .A(n379), .B(n21091), .Z(n21090) );
  XOR U20960 ( .A(n21092), .B(n21089), .Z(n21091) );
  XOR U20961 ( .A(n21093), .B(n21094), .Z(n21081) );
  AND U20962 ( .A(n21095), .B(n21096), .Z(n21094) );
  XOR U20963 ( .A(n21093), .B(n19282), .Z(n21096) );
  XOR U20964 ( .A(n21097), .B(n21098), .Z(n19282) );
  AND U20965 ( .A(n382), .B(n21099), .Z(n21098) );
  XOR U20966 ( .A(n21100), .B(n21097), .Z(n21099) );
  XNOR U20967 ( .A(n19279), .B(n21093), .Z(n21095) );
  XOR U20968 ( .A(n21101), .B(n21102), .Z(n19279) );
  AND U20969 ( .A(n379), .B(n21103), .Z(n21102) );
  XOR U20970 ( .A(n21104), .B(n21101), .Z(n21103) );
  XOR U20971 ( .A(n21105), .B(n21106), .Z(n21093) );
  AND U20972 ( .A(n21107), .B(n21108), .Z(n21106) );
  XOR U20973 ( .A(n21105), .B(n19294), .Z(n21108) );
  XOR U20974 ( .A(n21109), .B(n21110), .Z(n19294) );
  AND U20975 ( .A(n382), .B(n21111), .Z(n21110) );
  XOR U20976 ( .A(n21112), .B(n21109), .Z(n21111) );
  XNOR U20977 ( .A(n19291), .B(n21105), .Z(n21107) );
  XOR U20978 ( .A(n21113), .B(n21114), .Z(n19291) );
  AND U20979 ( .A(n379), .B(n21115), .Z(n21114) );
  XOR U20980 ( .A(n21116), .B(n21113), .Z(n21115) );
  XOR U20981 ( .A(n21117), .B(n21118), .Z(n21105) );
  AND U20982 ( .A(n21119), .B(n21120), .Z(n21118) );
  XOR U20983 ( .A(n21117), .B(n19306), .Z(n21120) );
  XOR U20984 ( .A(n21121), .B(n21122), .Z(n19306) );
  AND U20985 ( .A(n382), .B(n21123), .Z(n21122) );
  XOR U20986 ( .A(n21124), .B(n21121), .Z(n21123) );
  XNOR U20987 ( .A(n19303), .B(n21117), .Z(n21119) );
  XOR U20988 ( .A(n21125), .B(n21126), .Z(n19303) );
  AND U20989 ( .A(n379), .B(n21127), .Z(n21126) );
  XOR U20990 ( .A(n21128), .B(n21125), .Z(n21127) );
  XOR U20991 ( .A(n21129), .B(n21130), .Z(n21117) );
  AND U20992 ( .A(n21131), .B(n21132), .Z(n21130) );
  XOR U20993 ( .A(n21129), .B(n19318), .Z(n21132) );
  XOR U20994 ( .A(n21133), .B(n21134), .Z(n19318) );
  AND U20995 ( .A(n382), .B(n21135), .Z(n21134) );
  XOR U20996 ( .A(n21136), .B(n21133), .Z(n21135) );
  XNOR U20997 ( .A(n19315), .B(n21129), .Z(n21131) );
  XOR U20998 ( .A(n21137), .B(n21138), .Z(n19315) );
  AND U20999 ( .A(n379), .B(n21139), .Z(n21138) );
  XOR U21000 ( .A(n21140), .B(n21137), .Z(n21139) );
  XOR U21001 ( .A(n21141), .B(n21142), .Z(n21129) );
  AND U21002 ( .A(n21143), .B(n21144), .Z(n21142) );
  XOR U21003 ( .A(n21141), .B(n19330), .Z(n21144) );
  XOR U21004 ( .A(n21145), .B(n21146), .Z(n19330) );
  AND U21005 ( .A(n382), .B(n21147), .Z(n21146) );
  XOR U21006 ( .A(n21148), .B(n21145), .Z(n21147) );
  XNOR U21007 ( .A(n19327), .B(n21141), .Z(n21143) );
  XOR U21008 ( .A(n21149), .B(n21150), .Z(n19327) );
  AND U21009 ( .A(n379), .B(n21151), .Z(n21150) );
  XOR U21010 ( .A(n21152), .B(n21149), .Z(n21151) );
  XOR U21011 ( .A(n21153), .B(n21154), .Z(n21141) );
  AND U21012 ( .A(n21155), .B(n21156), .Z(n21154) );
  XOR U21013 ( .A(n21153), .B(n19342), .Z(n21156) );
  XOR U21014 ( .A(n21157), .B(n21158), .Z(n19342) );
  AND U21015 ( .A(n382), .B(n21159), .Z(n21158) );
  XOR U21016 ( .A(n21160), .B(n21157), .Z(n21159) );
  XNOR U21017 ( .A(n19339), .B(n21153), .Z(n21155) );
  XOR U21018 ( .A(n21161), .B(n21162), .Z(n19339) );
  AND U21019 ( .A(n379), .B(n21163), .Z(n21162) );
  XOR U21020 ( .A(n21164), .B(n21161), .Z(n21163) );
  XOR U21021 ( .A(n21165), .B(n21166), .Z(n21153) );
  AND U21022 ( .A(n21167), .B(n21168), .Z(n21166) );
  XOR U21023 ( .A(n21165), .B(n19354), .Z(n21168) );
  XOR U21024 ( .A(n21169), .B(n21170), .Z(n19354) );
  AND U21025 ( .A(n382), .B(n21171), .Z(n21170) );
  XOR U21026 ( .A(n21172), .B(n21169), .Z(n21171) );
  XNOR U21027 ( .A(n19351), .B(n21165), .Z(n21167) );
  XOR U21028 ( .A(n21173), .B(n21174), .Z(n19351) );
  AND U21029 ( .A(n379), .B(n21175), .Z(n21174) );
  XOR U21030 ( .A(n21176), .B(n21173), .Z(n21175) );
  XOR U21031 ( .A(n21177), .B(n21178), .Z(n21165) );
  AND U21032 ( .A(n21179), .B(n21180), .Z(n21178) );
  XOR U21033 ( .A(n21177), .B(n19366), .Z(n21180) );
  XOR U21034 ( .A(n21181), .B(n21182), .Z(n19366) );
  AND U21035 ( .A(n382), .B(n21183), .Z(n21182) );
  XOR U21036 ( .A(n21184), .B(n21181), .Z(n21183) );
  XNOR U21037 ( .A(n19363), .B(n21177), .Z(n21179) );
  XOR U21038 ( .A(n21185), .B(n21186), .Z(n19363) );
  AND U21039 ( .A(n379), .B(n21187), .Z(n21186) );
  XOR U21040 ( .A(n21188), .B(n21185), .Z(n21187) );
  XOR U21041 ( .A(n21189), .B(n21190), .Z(n21177) );
  AND U21042 ( .A(n21191), .B(n21192), .Z(n21190) );
  XOR U21043 ( .A(n21189), .B(n19378), .Z(n21192) );
  XOR U21044 ( .A(n21193), .B(n21194), .Z(n19378) );
  AND U21045 ( .A(n382), .B(n21195), .Z(n21194) );
  XOR U21046 ( .A(n21196), .B(n21193), .Z(n21195) );
  XNOR U21047 ( .A(n19375), .B(n21189), .Z(n21191) );
  XOR U21048 ( .A(n21197), .B(n21198), .Z(n19375) );
  AND U21049 ( .A(n379), .B(n21199), .Z(n21198) );
  XOR U21050 ( .A(n21200), .B(n21197), .Z(n21199) );
  XOR U21051 ( .A(n21201), .B(n21202), .Z(n21189) );
  AND U21052 ( .A(n21203), .B(n21204), .Z(n21202) );
  XOR U21053 ( .A(n21201), .B(n19390), .Z(n21204) );
  XOR U21054 ( .A(n21205), .B(n21206), .Z(n19390) );
  AND U21055 ( .A(n382), .B(n21207), .Z(n21206) );
  XOR U21056 ( .A(n21208), .B(n21205), .Z(n21207) );
  XNOR U21057 ( .A(n19387), .B(n21201), .Z(n21203) );
  XOR U21058 ( .A(n21209), .B(n21210), .Z(n19387) );
  AND U21059 ( .A(n379), .B(n21211), .Z(n21210) );
  XOR U21060 ( .A(n21212), .B(n21209), .Z(n21211) );
  XOR U21061 ( .A(n21213), .B(n21214), .Z(n21201) );
  AND U21062 ( .A(n21215), .B(n21216), .Z(n21214) );
  XOR U21063 ( .A(n21213), .B(n19402), .Z(n21216) );
  XOR U21064 ( .A(n21217), .B(n21218), .Z(n19402) );
  AND U21065 ( .A(n382), .B(n21219), .Z(n21218) );
  XOR U21066 ( .A(n21220), .B(n21217), .Z(n21219) );
  XNOR U21067 ( .A(n19399), .B(n21213), .Z(n21215) );
  XOR U21068 ( .A(n21221), .B(n21222), .Z(n19399) );
  AND U21069 ( .A(n379), .B(n21223), .Z(n21222) );
  XOR U21070 ( .A(n21224), .B(n21221), .Z(n21223) );
  XOR U21071 ( .A(n21225), .B(n21226), .Z(n21213) );
  AND U21072 ( .A(n21227), .B(n21228), .Z(n21226) );
  XOR U21073 ( .A(n21225), .B(n19414), .Z(n21228) );
  XOR U21074 ( .A(n21229), .B(n21230), .Z(n19414) );
  AND U21075 ( .A(n382), .B(n21231), .Z(n21230) );
  XOR U21076 ( .A(n21232), .B(n21229), .Z(n21231) );
  XNOR U21077 ( .A(n19411), .B(n21225), .Z(n21227) );
  XOR U21078 ( .A(n21233), .B(n21234), .Z(n19411) );
  AND U21079 ( .A(n379), .B(n21235), .Z(n21234) );
  XOR U21080 ( .A(n21236), .B(n21233), .Z(n21235) );
  XOR U21081 ( .A(n21237), .B(n21238), .Z(n21225) );
  AND U21082 ( .A(n21239), .B(n21240), .Z(n21238) );
  XOR U21083 ( .A(n21237), .B(n19426), .Z(n21240) );
  XOR U21084 ( .A(n21241), .B(n21242), .Z(n19426) );
  AND U21085 ( .A(n382), .B(n21243), .Z(n21242) );
  XOR U21086 ( .A(n21244), .B(n21241), .Z(n21243) );
  XNOR U21087 ( .A(n19423), .B(n21237), .Z(n21239) );
  XOR U21088 ( .A(n21245), .B(n21246), .Z(n19423) );
  AND U21089 ( .A(n379), .B(n21247), .Z(n21246) );
  XOR U21090 ( .A(n21248), .B(n21245), .Z(n21247) );
  XOR U21091 ( .A(n21249), .B(n21250), .Z(n21237) );
  AND U21092 ( .A(n21251), .B(n21252), .Z(n21250) );
  XOR U21093 ( .A(n21249), .B(n19438), .Z(n21252) );
  XOR U21094 ( .A(n21253), .B(n21254), .Z(n19438) );
  AND U21095 ( .A(n382), .B(n21255), .Z(n21254) );
  XOR U21096 ( .A(n21256), .B(n21253), .Z(n21255) );
  XNOR U21097 ( .A(n19435), .B(n21249), .Z(n21251) );
  XOR U21098 ( .A(n21257), .B(n21258), .Z(n19435) );
  AND U21099 ( .A(n379), .B(n21259), .Z(n21258) );
  XOR U21100 ( .A(n21260), .B(n21257), .Z(n21259) );
  XOR U21101 ( .A(n21261), .B(n21262), .Z(n21249) );
  AND U21102 ( .A(n21263), .B(n21264), .Z(n21262) );
  XOR U21103 ( .A(n21261), .B(n19450), .Z(n21264) );
  XOR U21104 ( .A(n21265), .B(n21266), .Z(n19450) );
  AND U21105 ( .A(n382), .B(n21267), .Z(n21266) );
  XOR U21106 ( .A(n21268), .B(n21265), .Z(n21267) );
  XNOR U21107 ( .A(n19447), .B(n21261), .Z(n21263) );
  XOR U21108 ( .A(n21269), .B(n21270), .Z(n19447) );
  AND U21109 ( .A(n379), .B(n21271), .Z(n21270) );
  XOR U21110 ( .A(n21272), .B(n21269), .Z(n21271) );
  XOR U21111 ( .A(n21273), .B(n21274), .Z(n21261) );
  AND U21112 ( .A(n21275), .B(n21276), .Z(n21274) );
  XOR U21113 ( .A(n21273), .B(n19462), .Z(n21276) );
  XOR U21114 ( .A(n21277), .B(n21278), .Z(n19462) );
  AND U21115 ( .A(n382), .B(n21279), .Z(n21278) );
  XOR U21116 ( .A(n21280), .B(n21277), .Z(n21279) );
  XNOR U21117 ( .A(n19459), .B(n21273), .Z(n21275) );
  XOR U21118 ( .A(n21281), .B(n21282), .Z(n19459) );
  AND U21119 ( .A(n379), .B(n21283), .Z(n21282) );
  XOR U21120 ( .A(n21284), .B(n21281), .Z(n21283) );
  XOR U21121 ( .A(n21285), .B(n21286), .Z(n21273) );
  AND U21122 ( .A(n21287), .B(n21288), .Z(n21286) );
  XOR U21123 ( .A(n21285), .B(n19474), .Z(n21288) );
  XOR U21124 ( .A(n21289), .B(n21290), .Z(n19474) );
  AND U21125 ( .A(n382), .B(n21291), .Z(n21290) );
  XOR U21126 ( .A(n21292), .B(n21289), .Z(n21291) );
  XNOR U21127 ( .A(n19471), .B(n21285), .Z(n21287) );
  XOR U21128 ( .A(n21293), .B(n21294), .Z(n19471) );
  AND U21129 ( .A(n379), .B(n21295), .Z(n21294) );
  XOR U21130 ( .A(n21296), .B(n21293), .Z(n21295) );
  XOR U21131 ( .A(n21297), .B(n21298), .Z(n21285) );
  AND U21132 ( .A(n21299), .B(n21300), .Z(n21298) );
  XOR U21133 ( .A(n21297), .B(n19486), .Z(n21300) );
  XOR U21134 ( .A(n21301), .B(n21302), .Z(n19486) );
  AND U21135 ( .A(n382), .B(n21303), .Z(n21302) );
  XOR U21136 ( .A(n21304), .B(n21301), .Z(n21303) );
  XNOR U21137 ( .A(n19483), .B(n21297), .Z(n21299) );
  XOR U21138 ( .A(n21305), .B(n21306), .Z(n19483) );
  AND U21139 ( .A(n379), .B(n21307), .Z(n21306) );
  XOR U21140 ( .A(n21308), .B(n21305), .Z(n21307) );
  XOR U21141 ( .A(n21309), .B(n21310), .Z(n21297) );
  AND U21142 ( .A(n21311), .B(n21312), .Z(n21310) );
  XOR U21143 ( .A(n21309), .B(n19498), .Z(n21312) );
  XOR U21144 ( .A(n21313), .B(n21314), .Z(n19498) );
  AND U21145 ( .A(n382), .B(n21315), .Z(n21314) );
  XOR U21146 ( .A(n21316), .B(n21313), .Z(n21315) );
  XNOR U21147 ( .A(n19495), .B(n21309), .Z(n21311) );
  XOR U21148 ( .A(n21317), .B(n21318), .Z(n19495) );
  AND U21149 ( .A(n379), .B(n21319), .Z(n21318) );
  XOR U21150 ( .A(n21320), .B(n21317), .Z(n21319) );
  XOR U21151 ( .A(n21321), .B(n21322), .Z(n21309) );
  AND U21152 ( .A(n21323), .B(n21324), .Z(n21322) );
  XOR U21153 ( .A(n21321), .B(n19510), .Z(n21324) );
  XOR U21154 ( .A(n21325), .B(n21326), .Z(n19510) );
  AND U21155 ( .A(n382), .B(n21327), .Z(n21326) );
  XOR U21156 ( .A(n21328), .B(n21325), .Z(n21327) );
  XNOR U21157 ( .A(n19507), .B(n21321), .Z(n21323) );
  XOR U21158 ( .A(n21329), .B(n21330), .Z(n19507) );
  AND U21159 ( .A(n379), .B(n21331), .Z(n21330) );
  XOR U21160 ( .A(n21332), .B(n21329), .Z(n21331) );
  XOR U21161 ( .A(n21333), .B(n21334), .Z(n21321) );
  AND U21162 ( .A(n21335), .B(n21336), .Z(n21334) );
  XOR U21163 ( .A(n21333), .B(n19522), .Z(n21336) );
  XOR U21164 ( .A(n21337), .B(n21338), .Z(n19522) );
  AND U21165 ( .A(n382), .B(n21339), .Z(n21338) );
  XOR U21166 ( .A(n21340), .B(n21337), .Z(n21339) );
  XNOR U21167 ( .A(n19519), .B(n21333), .Z(n21335) );
  XOR U21168 ( .A(n21341), .B(n21342), .Z(n19519) );
  AND U21169 ( .A(n379), .B(n21343), .Z(n21342) );
  XOR U21170 ( .A(n21344), .B(n21341), .Z(n21343) );
  XOR U21171 ( .A(n21345), .B(n21346), .Z(n21333) );
  AND U21172 ( .A(n21347), .B(n21348), .Z(n21346) );
  XOR U21173 ( .A(n21345), .B(n19534), .Z(n21348) );
  XOR U21174 ( .A(n21349), .B(n21350), .Z(n19534) );
  AND U21175 ( .A(n382), .B(n21351), .Z(n21350) );
  XOR U21176 ( .A(n21352), .B(n21349), .Z(n21351) );
  XNOR U21177 ( .A(n19531), .B(n21345), .Z(n21347) );
  XOR U21178 ( .A(n21353), .B(n21354), .Z(n19531) );
  AND U21179 ( .A(n379), .B(n21355), .Z(n21354) );
  XOR U21180 ( .A(n21356), .B(n21353), .Z(n21355) );
  XOR U21181 ( .A(n21357), .B(n21358), .Z(n21345) );
  AND U21182 ( .A(n21359), .B(n21360), .Z(n21358) );
  XOR U21183 ( .A(n21357), .B(n19546), .Z(n21360) );
  XOR U21184 ( .A(n21361), .B(n21362), .Z(n19546) );
  AND U21185 ( .A(n382), .B(n21363), .Z(n21362) );
  XOR U21186 ( .A(n21364), .B(n21361), .Z(n21363) );
  XNOR U21187 ( .A(n19543), .B(n21357), .Z(n21359) );
  XOR U21188 ( .A(n21365), .B(n21366), .Z(n19543) );
  AND U21189 ( .A(n379), .B(n21367), .Z(n21366) );
  XOR U21190 ( .A(n21368), .B(n21365), .Z(n21367) );
  XOR U21191 ( .A(n21369), .B(n21370), .Z(n21357) );
  AND U21192 ( .A(n21371), .B(n21372), .Z(n21370) );
  XOR U21193 ( .A(n21369), .B(n19558), .Z(n21372) );
  XOR U21194 ( .A(n21373), .B(n21374), .Z(n19558) );
  AND U21195 ( .A(n382), .B(n21375), .Z(n21374) );
  XOR U21196 ( .A(n21376), .B(n21373), .Z(n21375) );
  XNOR U21197 ( .A(n19555), .B(n21369), .Z(n21371) );
  XOR U21198 ( .A(n21377), .B(n21378), .Z(n19555) );
  AND U21199 ( .A(n379), .B(n21379), .Z(n21378) );
  XOR U21200 ( .A(n21380), .B(n21377), .Z(n21379) );
  XOR U21201 ( .A(n21381), .B(n21382), .Z(n21369) );
  AND U21202 ( .A(n21383), .B(n21384), .Z(n21382) );
  XOR U21203 ( .A(n21381), .B(n19570), .Z(n21384) );
  XOR U21204 ( .A(n21385), .B(n21386), .Z(n19570) );
  AND U21205 ( .A(n382), .B(n21387), .Z(n21386) );
  XOR U21206 ( .A(n21388), .B(n21385), .Z(n21387) );
  XNOR U21207 ( .A(n19567), .B(n21381), .Z(n21383) );
  XOR U21208 ( .A(n21389), .B(n21390), .Z(n19567) );
  AND U21209 ( .A(n379), .B(n21391), .Z(n21390) );
  XOR U21210 ( .A(n21392), .B(n21389), .Z(n21391) );
  XOR U21211 ( .A(n21393), .B(n21394), .Z(n21381) );
  AND U21212 ( .A(n21395), .B(n21396), .Z(n21394) );
  XOR U21213 ( .A(n21393), .B(n19582), .Z(n21396) );
  XOR U21214 ( .A(n21397), .B(n21398), .Z(n19582) );
  AND U21215 ( .A(n382), .B(n21399), .Z(n21398) );
  XOR U21216 ( .A(n21400), .B(n21397), .Z(n21399) );
  XNOR U21217 ( .A(n19579), .B(n21393), .Z(n21395) );
  XOR U21218 ( .A(n21401), .B(n21402), .Z(n19579) );
  AND U21219 ( .A(n379), .B(n21403), .Z(n21402) );
  XOR U21220 ( .A(n21404), .B(n21401), .Z(n21403) );
  XOR U21221 ( .A(n21405), .B(n21406), .Z(n21393) );
  AND U21222 ( .A(n21407), .B(n21408), .Z(n21406) );
  XOR U21223 ( .A(n19594), .B(n21405), .Z(n21408) );
  XOR U21224 ( .A(n21409), .B(n21410), .Z(n19594) );
  AND U21225 ( .A(n382), .B(n21411), .Z(n21410) );
  XOR U21226 ( .A(n21409), .B(n21412), .Z(n21411) );
  XNOR U21227 ( .A(n21405), .B(n19591), .Z(n21407) );
  XOR U21228 ( .A(n21413), .B(n21414), .Z(n19591) );
  AND U21229 ( .A(n379), .B(n21415), .Z(n21414) );
  XOR U21230 ( .A(n21413), .B(n21416), .Z(n21415) );
  XOR U21231 ( .A(n21417), .B(n21418), .Z(n21405) );
  AND U21232 ( .A(n21419), .B(n21420), .Z(n21418) );
  XNOR U21233 ( .A(n21421), .B(n19607), .Z(n21420) );
  XOR U21234 ( .A(n21422), .B(n21423), .Z(n19607) );
  AND U21235 ( .A(n382), .B(n21424), .Z(n21423) );
  XOR U21236 ( .A(n21425), .B(n21422), .Z(n21424) );
  XNOR U21237 ( .A(n19604), .B(n21417), .Z(n21419) );
  XOR U21238 ( .A(n21426), .B(n21427), .Z(n19604) );
  AND U21239 ( .A(n379), .B(n21428), .Z(n21427) );
  XOR U21240 ( .A(n21429), .B(n21426), .Z(n21428) );
  IV U21241 ( .A(n21421), .Z(n21417) );
  AND U21242 ( .A(n21053), .B(n21056), .Z(n21421) );
  XNOR U21243 ( .A(n21430), .B(n21431), .Z(n21056) );
  AND U21244 ( .A(n382), .B(n21432), .Z(n21431) );
  XNOR U21245 ( .A(n21433), .B(n21430), .Z(n21432) );
  XOR U21246 ( .A(n21434), .B(n21435), .Z(n382) );
  AND U21247 ( .A(n21436), .B(n21437), .Z(n21435) );
  XOR U21248 ( .A(n21064), .B(n21434), .Z(n21437) );
  IV U21249 ( .A(n21438), .Z(n21064) );
  AND U21250 ( .A(p_input[1279]), .B(p_input[1247]), .Z(n21438) );
  XOR U21251 ( .A(n21434), .B(n21061), .Z(n21436) );
  AND U21252 ( .A(p_input[1183]), .B(p_input[1215]), .Z(n21061) );
  XOR U21253 ( .A(n21439), .B(n21440), .Z(n21434) );
  AND U21254 ( .A(n21441), .B(n21442), .Z(n21440) );
  XOR U21255 ( .A(n21439), .B(n21076), .Z(n21442) );
  XNOR U21256 ( .A(p_input[1246]), .B(n21443), .Z(n21076) );
  AND U21257 ( .A(n470), .B(n21444), .Z(n21443) );
  XOR U21258 ( .A(p_input[1278]), .B(p_input[1246]), .Z(n21444) );
  XNOR U21259 ( .A(n21073), .B(n21439), .Z(n21441) );
  XOR U21260 ( .A(n21445), .B(n21446), .Z(n21073) );
  AND U21261 ( .A(n468), .B(n21447), .Z(n21446) );
  XOR U21262 ( .A(p_input[1214]), .B(p_input[1182]), .Z(n21447) );
  XOR U21263 ( .A(n21448), .B(n21449), .Z(n21439) );
  AND U21264 ( .A(n21450), .B(n21451), .Z(n21449) );
  XOR U21265 ( .A(n21448), .B(n21088), .Z(n21451) );
  XNOR U21266 ( .A(p_input[1245]), .B(n21452), .Z(n21088) );
  AND U21267 ( .A(n470), .B(n21453), .Z(n21452) );
  XOR U21268 ( .A(p_input[1277]), .B(p_input[1245]), .Z(n21453) );
  XNOR U21269 ( .A(n21085), .B(n21448), .Z(n21450) );
  XOR U21270 ( .A(n21454), .B(n21455), .Z(n21085) );
  AND U21271 ( .A(n468), .B(n21456), .Z(n21455) );
  XOR U21272 ( .A(p_input[1213]), .B(p_input[1181]), .Z(n21456) );
  XOR U21273 ( .A(n21457), .B(n21458), .Z(n21448) );
  AND U21274 ( .A(n21459), .B(n21460), .Z(n21458) );
  XOR U21275 ( .A(n21457), .B(n21100), .Z(n21460) );
  XNOR U21276 ( .A(p_input[1244]), .B(n21461), .Z(n21100) );
  AND U21277 ( .A(n470), .B(n21462), .Z(n21461) );
  XOR U21278 ( .A(p_input[1276]), .B(p_input[1244]), .Z(n21462) );
  XNOR U21279 ( .A(n21097), .B(n21457), .Z(n21459) );
  XOR U21280 ( .A(n21463), .B(n21464), .Z(n21097) );
  AND U21281 ( .A(n468), .B(n21465), .Z(n21464) );
  XOR U21282 ( .A(p_input[1212]), .B(p_input[1180]), .Z(n21465) );
  XOR U21283 ( .A(n21466), .B(n21467), .Z(n21457) );
  AND U21284 ( .A(n21468), .B(n21469), .Z(n21467) );
  XOR U21285 ( .A(n21466), .B(n21112), .Z(n21469) );
  XNOR U21286 ( .A(p_input[1243]), .B(n21470), .Z(n21112) );
  AND U21287 ( .A(n470), .B(n21471), .Z(n21470) );
  XOR U21288 ( .A(p_input[1275]), .B(p_input[1243]), .Z(n21471) );
  XNOR U21289 ( .A(n21109), .B(n21466), .Z(n21468) );
  XOR U21290 ( .A(n21472), .B(n21473), .Z(n21109) );
  AND U21291 ( .A(n468), .B(n21474), .Z(n21473) );
  XOR U21292 ( .A(p_input[1211]), .B(p_input[1179]), .Z(n21474) );
  XOR U21293 ( .A(n21475), .B(n21476), .Z(n21466) );
  AND U21294 ( .A(n21477), .B(n21478), .Z(n21476) );
  XOR U21295 ( .A(n21475), .B(n21124), .Z(n21478) );
  XNOR U21296 ( .A(p_input[1242]), .B(n21479), .Z(n21124) );
  AND U21297 ( .A(n470), .B(n21480), .Z(n21479) );
  XOR U21298 ( .A(p_input[1274]), .B(p_input[1242]), .Z(n21480) );
  XNOR U21299 ( .A(n21121), .B(n21475), .Z(n21477) );
  XOR U21300 ( .A(n21481), .B(n21482), .Z(n21121) );
  AND U21301 ( .A(n468), .B(n21483), .Z(n21482) );
  XOR U21302 ( .A(p_input[1210]), .B(p_input[1178]), .Z(n21483) );
  XOR U21303 ( .A(n21484), .B(n21485), .Z(n21475) );
  AND U21304 ( .A(n21486), .B(n21487), .Z(n21485) );
  XOR U21305 ( .A(n21484), .B(n21136), .Z(n21487) );
  XNOR U21306 ( .A(p_input[1241]), .B(n21488), .Z(n21136) );
  AND U21307 ( .A(n470), .B(n21489), .Z(n21488) );
  XOR U21308 ( .A(p_input[1273]), .B(p_input[1241]), .Z(n21489) );
  XNOR U21309 ( .A(n21133), .B(n21484), .Z(n21486) );
  XOR U21310 ( .A(n21490), .B(n21491), .Z(n21133) );
  AND U21311 ( .A(n468), .B(n21492), .Z(n21491) );
  XOR U21312 ( .A(p_input[1209]), .B(p_input[1177]), .Z(n21492) );
  XOR U21313 ( .A(n21493), .B(n21494), .Z(n21484) );
  AND U21314 ( .A(n21495), .B(n21496), .Z(n21494) );
  XOR U21315 ( .A(n21493), .B(n21148), .Z(n21496) );
  XNOR U21316 ( .A(p_input[1240]), .B(n21497), .Z(n21148) );
  AND U21317 ( .A(n470), .B(n21498), .Z(n21497) );
  XOR U21318 ( .A(p_input[1272]), .B(p_input[1240]), .Z(n21498) );
  XNOR U21319 ( .A(n21145), .B(n21493), .Z(n21495) );
  XOR U21320 ( .A(n21499), .B(n21500), .Z(n21145) );
  AND U21321 ( .A(n468), .B(n21501), .Z(n21500) );
  XOR U21322 ( .A(p_input[1208]), .B(p_input[1176]), .Z(n21501) );
  XOR U21323 ( .A(n21502), .B(n21503), .Z(n21493) );
  AND U21324 ( .A(n21504), .B(n21505), .Z(n21503) );
  XOR U21325 ( .A(n21502), .B(n21160), .Z(n21505) );
  XNOR U21326 ( .A(p_input[1239]), .B(n21506), .Z(n21160) );
  AND U21327 ( .A(n470), .B(n21507), .Z(n21506) );
  XOR U21328 ( .A(p_input[1271]), .B(p_input[1239]), .Z(n21507) );
  XNOR U21329 ( .A(n21157), .B(n21502), .Z(n21504) );
  XOR U21330 ( .A(n21508), .B(n21509), .Z(n21157) );
  AND U21331 ( .A(n468), .B(n21510), .Z(n21509) );
  XOR U21332 ( .A(p_input[1207]), .B(p_input[1175]), .Z(n21510) );
  XOR U21333 ( .A(n21511), .B(n21512), .Z(n21502) );
  AND U21334 ( .A(n21513), .B(n21514), .Z(n21512) );
  XOR U21335 ( .A(n21511), .B(n21172), .Z(n21514) );
  XNOR U21336 ( .A(p_input[1238]), .B(n21515), .Z(n21172) );
  AND U21337 ( .A(n470), .B(n21516), .Z(n21515) );
  XOR U21338 ( .A(p_input[1270]), .B(p_input[1238]), .Z(n21516) );
  XNOR U21339 ( .A(n21169), .B(n21511), .Z(n21513) );
  XOR U21340 ( .A(n21517), .B(n21518), .Z(n21169) );
  AND U21341 ( .A(n468), .B(n21519), .Z(n21518) );
  XOR U21342 ( .A(p_input[1206]), .B(p_input[1174]), .Z(n21519) );
  XOR U21343 ( .A(n21520), .B(n21521), .Z(n21511) );
  AND U21344 ( .A(n21522), .B(n21523), .Z(n21521) );
  XOR U21345 ( .A(n21520), .B(n21184), .Z(n21523) );
  XNOR U21346 ( .A(p_input[1237]), .B(n21524), .Z(n21184) );
  AND U21347 ( .A(n470), .B(n21525), .Z(n21524) );
  XOR U21348 ( .A(p_input[1269]), .B(p_input[1237]), .Z(n21525) );
  XNOR U21349 ( .A(n21181), .B(n21520), .Z(n21522) );
  XOR U21350 ( .A(n21526), .B(n21527), .Z(n21181) );
  AND U21351 ( .A(n468), .B(n21528), .Z(n21527) );
  XOR U21352 ( .A(p_input[1205]), .B(p_input[1173]), .Z(n21528) );
  XOR U21353 ( .A(n21529), .B(n21530), .Z(n21520) );
  AND U21354 ( .A(n21531), .B(n21532), .Z(n21530) );
  XOR U21355 ( .A(n21529), .B(n21196), .Z(n21532) );
  XNOR U21356 ( .A(p_input[1236]), .B(n21533), .Z(n21196) );
  AND U21357 ( .A(n470), .B(n21534), .Z(n21533) );
  XOR U21358 ( .A(p_input[1268]), .B(p_input[1236]), .Z(n21534) );
  XNOR U21359 ( .A(n21193), .B(n21529), .Z(n21531) );
  XOR U21360 ( .A(n21535), .B(n21536), .Z(n21193) );
  AND U21361 ( .A(n468), .B(n21537), .Z(n21536) );
  XOR U21362 ( .A(p_input[1204]), .B(p_input[1172]), .Z(n21537) );
  XOR U21363 ( .A(n21538), .B(n21539), .Z(n21529) );
  AND U21364 ( .A(n21540), .B(n21541), .Z(n21539) );
  XOR U21365 ( .A(n21538), .B(n21208), .Z(n21541) );
  XNOR U21366 ( .A(p_input[1235]), .B(n21542), .Z(n21208) );
  AND U21367 ( .A(n470), .B(n21543), .Z(n21542) );
  XOR U21368 ( .A(p_input[1267]), .B(p_input[1235]), .Z(n21543) );
  XNOR U21369 ( .A(n21205), .B(n21538), .Z(n21540) );
  XOR U21370 ( .A(n21544), .B(n21545), .Z(n21205) );
  AND U21371 ( .A(n468), .B(n21546), .Z(n21545) );
  XOR U21372 ( .A(p_input[1203]), .B(p_input[1171]), .Z(n21546) );
  XOR U21373 ( .A(n21547), .B(n21548), .Z(n21538) );
  AND U21374 ( .A(n21549), .B(n21550), .Z(n21548) );
  XOR U21375 ( .A(n21547), .B(n21220), .Z(n21550) );
  XNOR U21376 ( .A(p_input[1234]), .B(n21551), .Z(n21220) );
  AND U21377 ( .A(n470), .B(n21552), .Z(n21551) );
  XOR U21378 ( .A(p_input[1266]), .B(p_input[1234]), .Z(n21552) );
  XNOR U21379 ( .A(n21217), .B(n21547), .Z(n21549) );
  XOR U21380 ( .A(n21553), .B(n21554), .Z(n21217) );
  AND U21381 ( .A(n468), .B(n21555), .Z(n21554) );
  XOR U21382 ( .A(p_input[1202]), .B(p_input[1170]), .Z(n21555) );
  XOR U21383 ( .A(n21556), .B(n21557), .Z(n21547) );
  AND U21384 ( .A(n21558), .B(n21559), .Z(n21557) );
  XOR U21385 ( .A(n21556), .B(n21232), .Z(n21559) );
  XNOR U21386 ( .A(p_input[1233]), .B(n21560), .Z(n21232) );
  AND U21387 ( .A(n470), .B(n21561), .Z(n21560) );
  XOR U21388 ( .A(p_input[1265]), .B(p_input[1233]), .Z(n21561) );
  XNOR U21389 ( .A(n21229), .B(n21556), .Z(n21558) );
  XOR U21390 ( .A(n21562), .B(n21563), .Z(n21229) );
  AND U21391 ( .A(n468), .B(n21564), .Z(n21563) );
  XOR U21392 ( .A(p_input[1201]), .B(p_input[1169]), .Z(n21564) );
  XOR U21393 ( .A(n21565), .B(n21566), .Z(n21556) );
  AND U21394 ( .A(n21567), .B(n21568), .Z(n21566) );
  XOR U21395 ( .A(n21565), .B(n21244), .Z(n21568) );
  XNOR U21396 ( .A(p_input[1232]), .B(n21569), .Z(n21244) );
  AND U21397 ( .A(n470), .B(n21570), .Z(n21569) );
  XOR U21398 ( .A(p_input[1264]), .B(p_input[1232]), .Z(n21570) );
  XNOR U21399 ( .A(n21241), .B(n21565), .Z(n21567) );
  XOR U21400 ( .A(n21571), .B(n21572), .Z(n21241) );
  AND U21401 ( .A(n468), .B(n21573), .Z(n21572) );
  XOR U21402 ( .A(p_input[1200]), .B(p_input[1168]), .Z(n21573) );
  XOR U21403 ( .A(n21574), .B(n21575), .Z(n21565) );
  AND U21404 ( .A(n21576), .B(n21577), .Z(n21575) );
  XOR U21405 ( .A(n21574), .B(n21256), .Z(n21577) );
  XNOR U21406 ( .A(p_input[1231]), .B(n21578), .Z(n21256) );
  AND U21407 ( .A(n470), .B(n21579), .Z(n21578) );
  XOR U21408 ( .A(p_input[1263]), .B(p_input[1231]), .Z(n21579) );
  XNOR U21409 ( .A(n21253), .B(n21574), .Z(n21576) );
  XOR U21410 ( .A(n21580), .B(n21581), .Z(n21253) );
  AND U21411 ( .A(n468), .B(n21582), .Z(n21581) );
  XOR U21412 ( .A(p_input[1199]), .B(p_input[1167]), .Z(n21582) );
  XOR U21413 ( .A(n21583), .B(n21584), .Z(n21574) );
  AND U21414 ( .A(n21585), .B(n21586), .Z(n21584) );
  XOR U21415 ( .A(n21583), .B(n21268), .Z(n21586) );
  XNOR U21416 ( .A(p_input[1230]), .B(n21587), .Z(n21268) );
  AND U21417 ( .A(n470), .B(n21588), .Z(n21587) );
  XOR U21418 ( .A(p_input[1262]), .B(p_input[1230]), .Z(n21588) );
  XNOR U21419 ( .A(n21265), .B(n21583), .Z(n21585) );
  XOR U21420 ( .A(n21589), .B(n21590), .Z(n21265) );
  AND U21421 ( .A(n468), .B(n21591), .Z(n21590) );
  XOR U21422 ( .A(p_input[1198]), .B(p_input[1166]), .Z(n21591) );
  XOR U21423 ( .A(n21592), .B(n21593), .Z(n21583) );
  AND U21424 ( .A(n21594), .B(n21595), .Z(n21593) );
  XOR U21425 ( .A(n21592), .B(n21280), .Z(n21595) );
  XNOR U21426 ( .A(p_input[1229]), .B(n21596), .Z(n21280) );
  AND U21427 ( .A(n470), .B(n21597), .Z(n21596) );
  XOR U21428 ( .A(p_input[1261]), .B(p_input[1229]), .Z(n21597) );
  XNOR U21429 ( .A(n21277), .B(n21592), .Z(n21594) );
  XOR U21430 ( .A(n21598), .B(n21599), .Z(n21277) );
  AND U21431 ( .A(n468), .B(n21600), .Z(n21599) );
  XOR U21432 ( .A(p_input[1197]), .B(p_input[1165]), .Z(n21600) );
  XOR U21433 ( .A(n21601), .B(n21602), .Z(n21592) );
  AND U21434 ( .A(n21603), .B(n21604), .Z(n21602) );
  XOR U21435 ( .A(n21601), .B(n21292), .Z(n21604) );
  XNOR U21436 ( .A(p_input[1228]), .B(n21605), .Z(n21292) );
  AND U21437 ( .A(n470), .B(n21606), .Z(n21605) );
  XOR U21438 ( .A(p_input[1260]), .B(p_input[1228]), .Z(n21606) );
  XNOR U21439 ( .A(n21289), .B(n21601), .Z(n21603) );
  XOR U21440 ( .A(n21607), .B(n21608), .Z(n21289) );
  AND U21441 ( .A(n468), .B(n21609), .Z(n21608) );
  XOR U21442 ( .A(p_input[1196]), .B(p_input[1164]), .Z(n21609) );
  XOR U21443 ( .A(n21610), .B(n21611), .Z(n21601) );
  AND U21444 ( .A(n21612), .B(n21613), .Z(n21611) );
  XOR U21445 ( .A(n21610), .B(n21304), .Z(n21613) );
  XNOR U21446 ( .A(p_input[1227]), .B(n21614), .Z(n21304) );
  AND U21447 ( .A(n470), .B(n21615), .Z(n21614) );
  XOR U21448 ( .A(p_input[1259]), .B(p_input[1227]), .Z(n21615) );
  XNOR U21449 ( .A(n21301), .B(n21610), .Z(n21612) );
  XOR U21450 ( .A(n21616), .B(n21617), .Z(n21301) );
  AND U21451 ( .A(n468), .B(n21618), .Z(n21617) );
  XOR U21452 ( .A(p_input[1195]), .B(p_input[1163]), .Z(n21618) );
  XOR U21453 ( .A(n21619), .B(n21620), .Z(n21610) );
  AND U21454 ( .A(n21621), .B(n21622), .Z(n21620) );
  XOR U21455 ( .A(n21619), .B(n21316), .Z(n21622) );
  XNOR U21456 ( .A(p_input[1226]), .B(n21623), .Z(n21316) );
  AND U21457 ( .A(n470), .B(n21624), .Z(n21623) );
  XOR U21458 ( .A(p_input[1258]), .B(p_input[1226]), .Z(n21624) );
  XNOR U21459 ( .A(n21313), .B(n21619), .Z(n21621) );
  XOR U21460 ( .A(n21625), .B(n21626), .Z(n21313) );
  AND U21461 ( .A(n468), .B(n21627), .Z(n21626) );
  XOR U21462 ( .A(p_input[1194]), .B(p_input[1162]), .Z(n21627) );
  XOR U21463 ( .A(n21628), .B(n21629), .Z(n21619) );
  AND U21464 ( .A(n21630), .B(n21631), .Z(n21629) );
  XOR U21465 ( .A(n21628), .B(n21328), .Z(n21631) );
  XNOR U21466 ( .A(p_input[1225]), .B(n21632), .Z(n21328) );
  AND U21467 ( .A(n470), .B(n21633), .Z(n21632) );
  XOR U21468 ( .A(p_input[1257]), .B(p_input[1225]), .Z(n21633) );
  XNOR U21469 ( .A(n21325), .B(n21628), .Z(n21630) );
  XOR U21470 ( .A(n21634), .B(n21635), .Z(n21325) );
  AND U21471 ( .A(n468), .B(n21636), .Z(n21635) );
  XOR U21472 ( .A(p_input[1193]), .B(p_input[1161]), .Z(n21636) );
  XOR U21473 ( .A(n21637), .B(n21638), .Z(n21628) );
  AND U21474 ( .A(n21639), .B(n21640), .Z(n21638) );
  XOR U21475 ( .A(n21637), .B(n21340), .Z(n21640) );
  XNOR U21476 ( .A(p_input[1224]), .B(n21641), .Z(n21340) );
  AND U21477 ( .A(n470), .B(n21642), .Z(n21641) );
  XOR U21478 ( .A(p_input[1256]), .B(p_input[1224]), .Z(n21642) );
  XNOR U21479 ( .A(n21337), .B(n21637), .Z(n21639) );
  XOR U21480 ( .A(n21643), .B(n21644), .Z(n21337) );
  AND U21481 ( .A(n468), .B(n21645), .Z(n21644) );
  XOR U21482 ( .A(p_input[1192]), .B(p_input[1160]), .Z(n21645) );
  XOR U21483 ( .A(n21646), .B(n21647), .Z(n21637) );
  AND U21484 ( .A(n21648), .B(n21649), .Z(n21647) );
  XOR U21485 ( .A(n21646), .B(n21352), .Z(n21649) );
  XNOR U21486 ( .A(p_input[1223]), .B(n21650), .Z(n21352) );
  AND U21487 ( .A(n470), .B(n21651), .Z(n21650) );
  XOR U21488 ( .A(p_input[1255]), .B(p_input[1223]), .Z(n21651) );
  XNOR U21489 ( .A(n21349), .B(n21646), .Z(n21648) );
  XOR U21490 ( .A(n21652), .B(n21653), .Z(n21349) );
  AND U21491 ( .A(n468), .B(n21654), .Z(n21653) );
  XOR U21492 ( .A(p_input[1191]), .B(p_input[1159]), .Z(n21654) );
  XOR U21493 ( .A(n21655), .B(n21656), .Z(n21646) );
  AND U21494 ( .A(n21657), .B(n21658), .Z(n21656) );
  XOR U21495 ( .A(n21655), .B(n21364), .Z(n21658) );
  XNOR U21496 ( .A(p_input[1222]), .B(n21659), .Z(n21364) );
  AND U21497 ( .A(n470), .B(n21660), .Z(n21659) );
  XOR U21498 ( .A(p_input[1254]), .B(p_input[1222]), .Z(n21660) );
  XNOR U21499 ( .A(n21361), .B(n21655), .Z(n21657) );
  XOR U21500 ( .A(n21661), .B(n21662), .Z(n21361) );
  AND U21501 ( .A(n468), .B(n21663), .Z(n21662) );
  XOR U21502 ( .A(p_input[1190]), .B(p_input[1158]), .Z(n21663) );
  XOR U21503 ( .A(n21664), .B(n21665), .Z(n21655) );
  AND U21504 ( .A(n21666), .B(n21667), .Z(n21665) );
  XOR U21505 ( .A(n21664), .B(n21376), .Z(n21667) );
  XNOR U21506 ( .A(p_input[1221]), .B(n21668), .Z(n21376) );
  AND U21507 ( .A(n470), .B(n21669), .Z(n21668) );
  XOR U21508 ( .A(p_input[1253]), .B(p_input[1221]), .Z(n21669) );
  XNOR U21509 ( .A(n21373), .B(n21664), .Z(n21666) );
  XOR U21510 ( .A(n21670), .B(n21671), .Z(n21373) );
  AND U21511 ( .A(n468), .B(n21672), .Z(n21671) );
  XOR U21512 ( .A(p_input[1189]), .B(p_input[1157]), .Z(n21672) );
  XOR U21513 ( .A(n21673), .B(n21674), .Z(n21664) );
  AND U21514 ( .A(n21675), .B(n21676), .Z(n21674) );
  XOR U21515 ( .A(n21673), .B(n21388), .Z(n21676) );
  XNOR U21516 ( .A(p_input[1220]), .B(n21677), .Z(n21388) );
  AND U21517 ( .A(n470), .B(n21678), .Z(n21677) );
  XOR U21518 ( .A(p_input[1252]), .B(p_input[1220]), .Z(n21678) );
  XNOR U21519 ( .A(n21385), .B(n21673), .Z(n21675) );
  XOR U21520 ( .A(n21679), .B(n21680), .Z(n21385) );
  AND U21521 ( .A(n468), .B(n21681), .Z(n21680) );
  XOR U21522 ( .A(p_input[1188]), .B(p_input[1156]), .Z(n21681) );
  XOR U21523 ( .A(n21682), .B(n21683), .Z(n21673) );
  AND U21524 ( .A(n21684), .B(n21685), .Z(n21683) );
  XOR U21525 ( .A(n21682), .B(n21400), .Z(n21685) );
  XNOR U21526 ( .A(p_input[1219]), .B(n21686), .Z(n21400) );
  AND U21527 ( .A(n470), .B(n21687), .Z(n21686) );
  XOR U21528 ( .A(p_input[1251]), .B(p_input[1219]), .Z(n21687) );
  XNOR U21529 ( .A(n21397), .B(n21682), .Z(n21684) );
  XOR U21530 ( .A(n21688), .B(n21689), .Z(n21397) );
  AND U21531 ( .A(n468), .B(n21690), .Z(n21689) );
  XOR U21532 ( .A(p_input[1187]), .B(p_input[1155]), .Z(n21690) );
  XOR U21533 ( .A(n21691), .B(n21692), .Z(n21682) );
  AND U21534 ( .A(n21693), .B(n21694), .Z(n21692) );
  XOR U21535 ( .A(n21412), .B(n21691), .Z(n21694) );
  XNOR U21536 ( .A(p_input[1218]), .B(n21695), .Z(n21412) );
  AND U21537 ( .A(n470), .B(n21696), .Z(n21695) );
  XOR U21538 ( .A(p_input[1250]), .B(p_input[1218]), .Z(n21696) );
  XNOR U21539 ( .A(n21691), .B(n21409), .Z(n21693) );
  XOR U21540 ( .A(n21697), .B(n21698), .Z(n21409) );
  AND U21541 ( .A(n468), .B(n21699), .Z(n21698) );
  XOR U21542 ( .A(p_input[1186]), .B(p_input[1154]), .Z(n21699) );
  XOR U21543 ( .A(n21700), .B(n21701), .Z(n21691) );
  AND U21544 ( .A(n21702), .B(n21703), .Z(n21701) );
  XNOR U21545 ( .A(n21704), .B(n21425), .Z(n21703) );
  XNOR U21546 ( .A(p_input[1217]), .B(n21705), .Z(n21425) );
  AND U21547 ( .A(n470), .B(n21706), .Z(n21705) );
  XNOR U21548 ( .A(p_input[1249]), .B(n21707), .Z(n21706) );
  IV U21549 ( .A(p_input[1217]), .Z(n21707) );
  XNOR U21550 ( .A(n21422), .B(n21700), .Z(n21702) );
  XNOR U21551 ( .A(p_input[1153]), .B(n21708), .Z(n21422) );
  AND U21552 ( .A(n468), .B(n21709), .Z(n21708) );
  XOR U21553 ( .A(p_input[1185]), .B(p_input[1153]), .Z(n21709) );
  IV U21554 ( .A(n21704), .Z(n21700) );
  AND U21555 ( .A(n21430), .B(n21433), .Z(n21704) );
  XOR U21556 ( .A(p_input[1216]), .B(n21710), .Z(n21433) );
  AND U21557 ( .A(n470), .B(n21711), .Z(n21710) );
  XOR U21558 ( .A(p_input[1248]), .B(p_input[1216]), .Z(n21711) );
  XOR U21559 ( .A(n21712), .B(n21713), .Z(n470) );
  AND U21560 ( .A(n21714), .B(n21715), .Z(n21713) );
  XNOR U21561 ( .A(p_input[1279]), .B(n21712), .Z(n21715) );
  XOR U21562 ( .A(n21712), .B(p_input[1247]), .Z(n21714) );
  XOR U21563 ( .A(n21716), .B(n21717), .Z(n21712) );
  AND U21564 ( .A(n21718), .B(n21719), .Z(n21717) );
  XNOR U21565 ( .A(p_input[1278]), .B(n21716), .Z(n21719) );
  XOR U21566 ( .A(n21716), .B(p_input[1246]), .Z(n21718) );
  XOR U21567 ( .A(n21720), .B(n21721), .Z(n21716) );
  AND U21568 ( .A(n21722), .B(n21723), .Z(n21721) );
  XNOR U21569 ( .A(p_input[1277]), .B(n21720), .Z(n21723) );
  XOR U21570 ( .A(n21720), .B(p_input[1245]), .Z(n21722) );
  XOR U21571 ( .A(n21724), .B(n21725), .Z(n21720) );
  AND U21572 ( .A(n21726), .B(n21727), .Z(n21725) );
  XNOR U21573 ( .A(p_input[1276]), .B(n21724), .Z(n21727) );
  XOR U21574 ( .A(n21724), .B(p_input[1244]), .Z(n21726) );
  XOR U21575 ( .A(n21728), .B(n21729), .Z(n21724) );
  AND U21576 ( .A(n21730), .B(n21731), .Z(n21729) );
  XNOR U21577 ( .A(p_input[1275]), .B(n21728), .Z(n21731) );
  XOR U21578 ( .A(n21728), .B(p_input[1243]), .Z(n21730) );
  XOR U21579 ( .A(n21732), .B(n21733), .Z(n21728) );
  AND U21580 ( .A(n21734), .B(n21735), .Z(n21733) );
  XNOR U21581 ( .A(p_input[1274]), .B(n21732), .Z(n21735) );
  XOR U21582 ( .A(n21732), .B(p_input[1242]), .Z(n21734) );
  XOR U21583 ( .A(n21736), .B(n21737), .Z(n21732) );
  AND U21584 ( .A(n21738), .B(n21739), .Z(n21737) );
  XNOR U21585 ( .A(p_input[1273]), .B(n21736), .Z(n21739) );
  XOR U21586 ( .A(n21736), .B(p_input[1241]), .Z(n21738) );
  XOR U21587 ( .A(n21740), .B(n21741), .Z(n21736) );
  AND U21588 ( .A(n21742), .B(n21743), .Z(n21741) );
  XNOR U21589 ( .A(p_input[1272]), .B(n21740), .Z(n21743) );
  XOR U21590 ( .A(n21740), .B(p_input[1240]), .Z(n21742) );
  XOR U21591 ( .A(n21744), .B(n21745), .Z(n21740) );
  AND U21592 ( .A(n21746), .B(n21747), .Z(n21745) );
  XNOR U21593 ( .A(p_input[1271]), .B(n21744), .Z(n21747) );
  XOR U21594 ( .A(n21744), .B(p_input[1239]), .Z(n21746) );
  XOR U21595 ( .A(n21748), .B(n21749), .Z(n21744) );
  AND U21596 ( .A(n21750), .B(n21751), .Z(n21749) );
  XNOR U21597 ( .A(p_input[1270]), .B(n21748), .Z(n21751) );
  XOR U21598 ( .A(n21748), .B(p_input[1238]), .Z(n21750) );
  XOR U21599 ( .A(n21752), .B(n21753), .Z(n21748) );
  AND U21600 ( .A(n21754), .B(n21755), .Z(n21753) );
  XNOR U21601 ( .A(p_input[1269]), .B(n21752), .Z(n21755) );
  XOR U21602 ( .A(n21752), .B(p_input[1237]), .Z(n21754) );
  XOR U21603 ( .A(n21756), .B(n21757), .Z(n21752) );
  AND U21604 ( .A(n21758), .B(n21759), .Z(n21757) );
  XNOR U21605 ( .A(p_input[1268]), .B(n21756), .Z(n21759) );
  XOR U21606 ( .A(n21756), .B(p_input[1236]), .Z(n21758) );
  XOR U21607 ( .A(n21760), .B(n21761), .Z(n21756) );
  AND U21608 ( .A(n21762), .B(n21763), .Z(n21761) );
  XNOR U21609 ( .A(p_input[1267]), .B(n21760), .Z(n21763) );
  XOR U21610 ( .A(n21760), .B(p_input[1235]), .Z(n21762) );
  XOR U21611 ( .A(n21764), .B(n21765), .Z(n21760) );
  AND U21612 ( .A(n21766), .B(n21767), .Z(n21765) );
  XNOR U21613 ( .A(p_input[1266]), .B(n21764), .Z(n21767) );
  XOR U21614 ( .A(n21764), .B(p_input[1234]), .Z(n21766) );
  XOR U21615 ( .A(n21768), .B(n21769), .Z(n21764) );
  AND U21616 ( .A(n21770), .B(n21771), .Z(n21769) );
  XNOR U21617 ( .A(p_input[1265]), .B(n21768), .Z(n21771) );
  XOR U21618 ( .A(n21768), .B(p_input[1233]), .Z(n21770) );
  XOR U21619 ( .A(n21772), .B(n21773), .Z(n21768) );
  AND U21620 ( .A(n21774), .B(n21775), .Z(n21773) );
  XNOR U21621 ( .A(p_input[1264]), .B(n21772), .Z(n21775) );
  XOR U21622 ( .A(n21772), .B(p_input[1232]), .Z(n21774) );
  XOR U21623 ( .A(n21776), .B(n21777), .Z(n21772) );
  AND U21624 ( .A(n21778), .B(n21779), .Z(n21777) );
  XNOR U21625 ( .A(p_input[1263]), .B(n21776), .Z(n21779) );
  XOR U21626 ( .A(n21776), .B(p_input[1231]), .Z(n21778) );
  XOR U21627 ( .A(n21780), .B(n21781), .Z(n21776) );
  AND U21628 ( .A(n21782), .B(n21783), .Z(n21781) );
  XNOR U21629 ( .A(p_input[1262]), .B(n21780), .Z(n21783) );
  XOR U21630 ( .A(n21780), .B(p_input[1230]), .Z(n21782) );
  XOR U21631 ( .A(n21784), .B(n21785), .Z(n21780) );
  AND U21632 ( .A(n21786), .B(n21787), .Z(n21785) );
  XNOR U21633 ( .A(p_input[1261]), .B(n21784), .Z(n21787) );
  XOR U21634 ( .A(n21784), .B(p_input[1229]), .Z(n21786) );
  XOR U21635 ( .A(n21788), .B(n21789), .Z(n21784) );
  AND U21636 ( .A(n21790), .B(n21791), .Z(n21789) );
  XNOR U21637 ( .A(p_input[1260]), .B(n21788), .Z(n21791) );
  XOR U21638 ( .A(n21788), .B(p_input[1228]), .Z(n21790) );
  XOR U21639 ( .A(n21792), .B(n21793), .Z(n21788) );
  AND U21640 ( .A(n21794), .B(n21795), .Z(n21793) );
  XNOR U21641 ( .A(p_input[1259]), .B(n21792), .Z(n21795) );
  XOR U21642 ( .A(n21792), .B(p_input[1227]), .Z(n21794) );
  XOR U21643 ( .A(n21796), .B(n21797), .Z(n21792) );
  AND U21644 ( .A(n21798), .B(n21799), .Z(n21797) );
  XNOR U21645 ( .A(p_input[1258]), .B(n21796), .Z(n21799) );
  XOR U21646 ( .A(n21796), .B(p_input[1226]), .Z(n21798) );
  XOR U21647 ( .A(n21800), .B(n21801), .Z(n21796) );
  AND U21648 ( .A(n21802), .B(n21803), .Z(n21801) );
  XNOR U21649 ( .A(p_input[1257]), .B(n21800), .Z(n21803) );
  XOR U21650 ( .A(n21800), .B(p_input[1225]), .Z(n21802) );
  XOR U21651 ( .A(n21804), .B(n21805), .Z(n21800) );
  AND U21652 ( .A(n21806), .B(n21807), .Z(n21805) );
  XNOR U21653 ( .A(p_input[1256]), .B(n21804), .Z(n21807) );
  XOR U21654 ( .A(n21804), .B(p_input[1224]), .Z(n21806) );
  XOR U21655 ( .A(n21808), .B(n21809), .Z(n21804) );
  AND U21656 ( .A(n21810), .B(n21811), .Z(n21809) );
  XNOR U21657 ( .A(p_input[1255]), .B(n21808), .Z(n21811) );
  XOR U21658 ( .A(n21808), .B(p_input[1223]), .Z(n21810) );
  XOR U21659 ( .A(n21812), .B(n21813), .Z(n21808) );
  AND U21660 ( .A(n21814), .B(n21815), .Z(n21813) );
  XNOR U21661 ( .A(p_input[1254]), .B(n21812), .Z(n21815) );
  XOR U21662 ( .A(n21812), .B(p_input[1222]), .Z(n21814) );
  XOR U21663 ( .A(n21816), .B(n21817), .Z(n21812) );
  AND U21664 ( .A(n21818), .B(n21819), .Z(n21817) );
  XNOR U21665 ( .A(p_input[1253]), .B(n21816), .Z(n21819) );
  XOR U21666 ( .A(n21816), .B(p_input[1221]), .Z(n21818) );
  XOR U21667 ( .A(n21820), .B(n21821), .Z(n21816) );
  AND U21668 ( .A(n21822), .B(n21823), .Z(n21821) );
  XNOR U21669 ( .A(p_input[1252]), .B(n21820), .Z(n21823) );
  XOR U21670 ( .A(n21820), .B(p_input[1220]), .Z(n21822) );
  XOR U21671 ( .A(n21824), .B(n21825), .Z(n21820) );
  AND U21672 ( .A(n21826), .B(n21827), .Z(n21825) );
  XNOR U21673 ( .A(p_input[1251]), .B(n21824), .Z(n21827) );
  XOR U21674 ( .A(n21824), .B(p_input[1219]), .Z(n21826) );
  XOR U21675 ( .A(n21828), .B(n21829), .Z(n21824) );
  AND U21676 ( .A(n21830), .B(n21831), .Z(n21829) );
  XNOR U21677 ( .A(p_input[1250]), .B(n21828), .Z(n21831) );
  XOR U21678 ( .A(n21828), .B(p_input[1218]), .Z(n21830) );
  XNOR U21679 ( .A(n21832), .B(n21833), .Z(n21828) );
  AND U21680 ( .A(n21834), .B(n21835), .Z(n21833) );
  XOR U21681 ( .A(p_input[1249]), .B(n21832), .Z(n21835) );
  XNOR U21682 ( .A(p_input[1217]), .B(n21832), .Z(n21834) );
  AND U21683 ( .A(p_input[1248]), .B(n21836), .Z(n21832) );
  IV U21684 ( .A(p_input[1216]), .Z(n21836) );
  XNOR U21685 ( .A(p_input[1152]), .B(n21837), .Z(n21430) );
  AND U21686 ( .A(n468), .B(n21838), .Z(n21837) );
  XOR U21687 ( .A(p_input[1184]), .B(p_input[1152]), .Z(n21838) );
  XOR U21688 ( .A(n21839), .B(n21840), .Z(n468) );
  AND U21689 ( .A(n21841), .B(n21842), .Z(n21840) );
  XNOR U21690 ( .A(p_input[1215]), .B(n21839), .Z(n21842) );
  XOR U21691 ( .A(n21839), .B(p_input[1183]), .Z(n21841) );
  XOR U21692 ( .A(n21843), .B(n21844), .Z(n21839) );
  AND U21693 ( .A(n21845), .B(n21846), .Z(n21844) );
  XNOR U21694 ( .A(p_input[1214]), .B(n21843), .Z(n21846) );
  XNOR U21695 ( .A(n21843), .B(n21445), .Z(n21845) );
  IV U21696 ( .A(p_input[1182]), .Z(n21445) );
  XOR U21697 ( .A(n21847), .B(n21848), .Z(n21843) );
  AND U21698 ( .A(n21849), .B(n21850), .Z(n21848) );
  XNOR U21699 ( .A(p_input[1213]), .B(n21847), .Z(n21850) );
  XNOR U21700 ( .A(n21847), .B(n21454), .Z(n21849) );
  IV U21701 ( .A(p_input[1181]), .Z(n21454) );
  XOR U21702 ( .A(n21851), .B(n21852), .Z(n21847) );
  AND U21703 ( .A(n21853), .B(n21854), .Z(n21852) );
  XNOR U21704 ( .A(p_input[1212]), .B(n21851), .Z(n21854) );
  XNOR U21705 ( .A(n21851), .B(n21463), .Z(n21853) );
  IV U21706 ( .A(p_input[1180]), .Z(n21463) );
  XOR U21707 ( .A(n21855), .B(n21856), .Z(n21851) );
  AND U21708 ( .A(n21857), .B(n21858), .Z(n21856) );
  XNOR U21709 ( .A(p_input[1211]), .B(n21855), .Z(n21858) );
  XNOR U21710 ( .A(n21855), .B(n21472), .Z(n21857) );
  IV U21711 ( .A(p_input[1179]), .Z(n21472) );
  XOR U21712 ( .A(n21859), .B(n21860), .Z(n21855) );
  AND U21713 ( .A(n21861), .B(n21862), .Z(n21860) );
  XNOR U21714 ( .A(p_input[1210]), .B(n21859), .Z(n21862) );
  XNOR U21715 ( .A(n21859), .B(n21481), .Z(n21861) );
  IV U21716 ( .A(p_input[1178]), .Z(n21481) );
  XOR U21717 ( .A(n21863), .B(n21864), .Z(n21859) );
  AND U21718 ( .A(n21865), .B(n21866), .Z(n21864) );
  XNOR U21719 ( .A(p_input[1209]), .B(n21863), .Z(n21866) );
  XNOR U21720 ( .A(n21863), .B(n21490), .Z(n21865) );
  IV U21721 ( .A(p_input[1177]), .Z(n21490) );
  XOR U21722 ( .A(n21867), .B(n21868), .Z(n21863) );
  AND U21723 ( .A(n21869), .B(n21870), .Z(n21868) );
  XNOR U21724 ( .A(p_input[1208]), .B(n21867), .Z(n21870) );
  XNOR U21725 ( .A(n21867), .B(n21499), .Z(n21869) );
  IV U21726 ( .A(p_input[1176]), .Z(n21499) );
  XOR U21727 ( .A(n21871), .B(n21872), .Z(n21867) );
  AND U21728 ( .A(n21873), .B(n21874), .Z(n21872) );
  XNOR U21729 ( .A(p_input[1207]), .B(n21871), .Z(n21874) );
  XNOR U21730 ( .A(n21871), .B(n21508), .Z(n21873) );
  IV U21731 ( .A(p_input[1175]), .Z(n21508) );
  XOR U21732 ( .A(n21875), .B(n21876), .Z(n21871) );
  AND U21733 ( .A(n21877), .B(n21878), .Z(n21876) );
  XNOR U21734 ( .A(p_input[1206]), .B(n21875), .Z(n21878) );
  XNOR U21735 ( .A(n21875), .B(n21517), .Z(n21877) );
  IV U21736 ( .A(p_input[1174]), .Z(n21517) );
  XOR U21737 ( .A(n21879), .B(n21880), .Z(n21875) );
  AND U21738 ( .A(n21881), .B(n21882), .Z(n21880) );
  XNOR U21739 ( .A(p_input[1205]), .B(n21879), .Z(n21882) );
  XNOR U21740 ( .A(n21879), .B(n21526), .Z(n21881) );
  IV U21741 ( .A(p_input[1173]), .Z(n21526) );
  XOR U21742 ( .A(n21883), .B(n21884), .Z(n21879) );
  AND U21743 ( .A(n21885), .B(n21886), .Z(n21884) );
  XNOR U21744 ( .A(p_input[1204]), .B(n21883), .Z(n21886) );
  XNOR U21745 ( .A(n21883), .B(n21535), .Z(n21885) );
  IV U21746 ( .A(p_input[1172]), .Z(n21535) );
  XOR U21747 ( .A(n21887), .B(n21888), .Z(n21883) );
  AND U21748 ( .A(n21889), .B(n21890), .Z(n21888) );
  XNOR U21749 ( .A(p_input[1203]), .B(n21887), .Z(n21890) );
  XNOR U21750 ( .A(n21887), .B(n21544), .Z(n21889) );
  IV U21751 ( .A(p_input[1171]), .Z(n21544) );
  XOR U21752 ( .A(n21891), .B(n21892), .Z(n21887) );
  AND U21753 ( .A(n21893), .B(n21894), .Z(n21892) );
  XNOR U21754 ( .A(p_input[1202]), .B(n21891), .Z(n21894) );
  XNOR U21755 ( .A(n21891), .B(n21553), .Z(n21893) );
  IV U21756 ( .A(p_input[1170]), .Z(n21553) );
  XOR U21757 ( .A(n21895), .B(n21896), .Z(n21891) );
  AND U21758 ( .A(n21897), .B(n21898), .Z(n21896) );
  XNOR U21759 ( .A(p_input[1201]), .B(n21895), .Z(n21898) );
  XNOR U21760 ( .A(n21895), .B(n21562), .Z(n21897) );
  IV U21761 ( .A(p_input[1169]), .Z(n21562) );
  XOR U21762 ( .A(n21899), .B(n21900), .Z(n21895) );
  AND U21763 ( .A(n21901), .B(n21902), .Z(n21900) );
  XNOR U21764 ( .A(p_input[1200]), .B(n21899), .Z(n21902) );
  XNOR U21765 ( .A(n21899), .B(n21571), .Z(n21901) );
  IV U21766 ( .A(p_input[1168]), .Z(n21571) );
  XOR U21767 ( .A(n21903), .B(n21904), .Z(n21899) );
  AND U21768 ( .A(n21905), .B(n21906), .Z(n21904) );
  XNOR U21769 ( .A(p_input[1199]), .B(n21903), .Z(n21906) );
  XNOR U21770 ( .A(n21903), .B(n21580), .Z(n21905) );
  IV U21771 ( .A(p_input[1167]), .Z(n21580) );
  XOR U21772 ( .A(n21907), .B(n21908), .Z(n21903) );
  AND U21773 ( .A(n21909), .B(n21910), .Z(n21908) );
  XNOR U21774 ( .A(p_input[1198]), .B(n21907), .Z(n21910) );
  XNOR U21775 ( .A(n21907), .B(n21589), .Z(n21909) );
  IV U21776 ( .A(p_input[1166]), .Z(n21589) );
  XOR U21777 ( .A(n21911), .B(n21912), .Z(n21907) );
  AND U21778 ( .A(n21913), .B(n21914), .Z(n21912) );
  XNOR U21779 ( .A(p_input[1197]), .B(n21911), .Z(n21914) );
  XNOR U21780 ( .A(n21911), .B(n21598), .Z(n21913) );
  IV U21781 ( .A(p_input[1165]), .Z(n21598) );
  XOR U21782 ( .A(n21915), .B(n21916), .Z(n21911) );
  AND U21783 ( .A(n21917), .B(n21918), .Z(n21916) );
  XNOR U21784 ( .A(p_input[1196]), .B(n21915), .Z(n21918) );
  XNOR U21785 ( .A(n21915), .B(n21607), .Z(n21917) );
  IV U21786 ( .A(p_input[1164]), .Z(n21607) );
  XOR U21787 ( .A(n21919), .B(n21920), .Z(n21915) );
  AND U21788 ( .A(n21921), .B(n21922), .Z(n21920) );
  XNOR U21789 ( .A(p_input[1195]), .B(n21919), .Z(n21922) );
  XNOR U21790 ( .A(n21919), .B(n21616), .Z(n21921) );
  IV U21791 ( .A(p_input[1163]), .Z(n21616) );
  XOR U21792 ( .A(n21923), .B(n21924), .Z(n21919) );
  AND U21793 ( .A(n21925), .B(n21926), .Z(n21924) );
  XNOR U21794 ( .A(p_input[1194]), .B(n21923), .Z(n21926) );
  XNOR U21795 ( .A(n21923), .B(n21625), .Z(n21925) );
  IV U21796 ( .A(p_input[1162]), .Z(n21625) );
  XOR U21797 ( .A(n21927), .B(n21928), .Z(n21923) );
  AND U21798 ( .A(n21929), .B(n21930), .Z(n21928) );
  XNOR U21799 ( .A(p_input[1193]), .B(n21927), .Z(n21930) );
  XNOR U21800 ( .A(n21927), .B(n21634), .Z(n21929) );
  IV U21801 ( .A(p_input[1161]), .Z(n21634) );
  XOR U21802 ( .A(n21931), .B(n21932), .Z(n21927) );
  AND U21803 ( .A(n21933), .B(n21934), .Z(n21932) );
  XNOR U21804 ( .A(p_input[1192]), .B(n21931), .Z(n21934) );
  XNOR U21805 ( .A(n21931), .B(n21643), .Z(n21933) );
  IV U21806 ( .A(p_input[1160]), .Z(n21643) );
  XOR U21807 ( .A(n21935), .B(n21936), .Z(n21931) );
  AND U21808 ( .A(n21937), .B(n21938), .Z(n21936) );
  XNOR U21809 ( .A(p_input[1191]), .B(n21935), .Z(n21938) );
  XNOR U21810 ( .A(n21935), .B(n21652), .Z(n21937) );
  IV U21811 ( .A(p_input[1159]), .Z(n21652) );
  XOR U21812 ( .A(n21939), .B(n21940), .Z(n21935) );
  AND U21813 ( .A(n21941), .B(n21942), .Z(n21940) );
  XNOR U21814 ( .A(p_input[1190]), .B(n21939), .Z(n21942) );
  XNOR U21815 ( .A(n21939), .B(n21661), .Z(n21941) );
  IV U21816 ( .A(p_input[1158]), .Z(n21661) );
  XOR U21817 ( .A(n21943), .B(n21944), .Z(n21939) );
  AND U21818 ( .A(n21945), .B(n21946), .Z(n21944) );
  XNOR U21819 ( .A(p_input[1189]), .B(n21943), .Z(n21946) );
  XNOR U21820 ( .A(n21943), .B(n21670), .Z(n21945) );
  IV U21821 ( .A(p_input[1157]), .Z(n21670) );
  XOR U21822 ( .A(n21947), .B(n21948), .Z(n21943) );
  AND U21823 ( .A(n21949), .B(n21950), .Z(n21948) );
  XNOR U21824 ( .A(p_input[1188]), .B(n21947), .Z(n21950) );
  XNOR U21825 ( .A(n21947), .B(n21679), .Z(n21949) );
  IV U21826 ( .A(p_input[1156]), .Z(n21679) );
  XOR U21827 ( .A(n21951), .B(n21952), .Z(n21947) );
  AND U21828 ( .A(n21953), .B(n21954), .Z(n21952) );
  XNOR U21829 ( .A(p_input[1187]), .B(n21951), .Z(n21954) );
  XNOR U21830 ( .A(n21951), .B(n21688), .Z(n21953) );
  IV U21831 ( .A(p_input[1155]), .Z(n21688) );
  XOR U21832 ( .A(n21955), .B(n21956), .Z(n21951) );
  AND U21833 ( .A(n21957), .B(n21958), .Z(n21956) );
  XNOR U21834 ( .A(p_input[1186]), .B(n21955), .Z(n21958) );
  XNOR U21835 ( .A(n21955), .B(n21697), .Z(n21957) );
  IV U21836 ( .A(p_input[1154]), .Z(n21697) );
  XNOR U21837 ( .A(n21959), .B(n21960), .Z(n21955) );
  AND U21838 ( .A(n21961), .B(n21962), .Z(n21960) );
  XOR U21839 ( .A(p_input[1185]), .B(n21959), .Z(n21962) );
  XNOR U21840 ( .A(p_input[1153]), .B(n21959), .Z(n21961) );
  AND U21841 ( .A(p_input[1184]), .B(n21963), .Z(n21959) );
  IV U21842 ( .A(p_input[1152]), .Z(n21963) );
  XOR U21843 ( .A(n21964), .B(n21965), .Z(n21053) );
  AND U21844 ( .A(n379), .B(n21966), .Z(n21965) );
  XNOR U21845 ( .A(n21967), .B(n21964), .Z(n21966) );
  XOR U21846 ( .A(n21968), .B(n21969), .Z(n379) );
  AND U21847 ( .A(n21970), .B(n21971), .Z(n21969) );
  XNOR U21848 ( .A(n21068), .B(n21968), .Z(n21971) );
  AND U21849 ( .A(p_input[1151]), .B(p_input[1119]), .Z(n21068) );
  XNOR U21850 ( .A(n21968), .B(n21065), .Z(n21970) );
  IV U21851 ( .A(n21972), .Z(n21065) );
  AND U21852 ( .A(p_input[1055]), .B(p_input[1087]), .Z(n21972) );
  XOR U21853 ( .A(n21973), .B(n21974), .Z(n21968) );
  AND U21854 ( .A(n21975), .B(n21976), .Z(n21974) );
  XOR U21855 ( .A(n21973), .B(n21080), .Z(n21976) );
  XNOR U21856 ( .A(p_input[1118]), .B(n21977), .Z(n21080) );
  AND U21857 ( .A(n474), .B(n21978), .Z(n21977) );
  XOR U21858 ( .A(p_input[1150]), .B(p_input[1118]), .Z(n21978) );
  XNOR U21859 ( .A(n21077), .B(n21973), .Z(n21975) );
  XOR U21860 ( .A(n21979), .B(n21980), .Z(n21077) );
  AND U21861 ( .A(n471), .B(n21981), .Z(n21980) );
  XOR U21862 ( .A(p_input[1086]), .B(p_input[1054]), .Z(n21981) );
  XOR U21863 ( .A(n21982), .B(n21983), .Z(n21973) );
  AND U21864 ( .A(n21984), .B(n21985), .Z(n21983) );
  XOR U21865 ( .A(n21982), .B(n21092), .Z(n21985) );
  XNOR U21866 ( .A(p_input[1117]), .B(n21986), .Z(n21092) );
  AND U21867 ( .A(n474), .B(n21987), .Z(n21986) );
  XOR U21868 ( .A(p_input[1149]), .B(p_input[1117]), .Z(n21987) );
  XNOR U21869 ( .A(n21089), .B(n21982), .Z(n21984) );
  XOR U21870 ( .A(n21988), .B(n21989), .Z(n21089) );
  AND U21871 ( .A(n471), .B(n21990), .Z(n21989) );
  XOR U21872 ( .A(p_input[1085]), .B(p_input[1053]), .Z(n21990) );
  XOR U21873 ( .A(n21991), .B(n21992), .Z(n21982) );
  AND U21874 ( .A(n21993), .B(n21994), .Z(n21992) );
  XOR U21875 ( .A(n21991), .B(n21104), .Z(n21994) );
  XNOR U21876 ( .A(p_input[1116]), .B(n21995), .Z(n21104) );
  AND U21877 ( .A(n474), .B(n21996), .Z(n21995) );
  XOR U21878 ( .A(p_input[1148]), .B(p_input[1116]), .Z(n21996) );
  XNOR U21879 ( .A(n21101), .B(n21991), .Z(n21993) );
  XOR U21880 ( .A(n21997), .B(n21998), .Z(n21101) );
  AND U21881 ( .A(n471), .B(n21999), .Z(n21998) );
  XOR U21882 ( .A(p_input[1084]), .B(p_input[1052]), .Z(n21999) );
  XOR U21883 ( .A(n22000), .B(n22001), .Z(n21991) );
  AND U21884 ( .A(n22002), .B(n22003), .Z(n22001) );
  XOR U21885 ( .A(n22000), .B(n21116), .Z(n22003) );
  XNOR U21886 ( .A(p_input[1115]), .B(n22004), .Z(n21116) );
  AND U21887 ( .A(n474), .B(n22005), .Z(n22004) );
  XOR U21888 ( .A(p_input[1147]), .B(p_input[1115]), .Z(n22005) );
  XNOR U21889 ( .A(n21113), .B(n22000), .Z(n22002) );
  XOR U21890 ( .A(n22006), .B(n22007), .Z(n21113) );
  AND U21891 ( .A(n471), .B(n22008), .Z(n22007) );
  XOR U21892 ( .A(p_input[1083]), .B(p_input[1051]), .Z(n22008) );
  XOR U21893 ( .A(n22009), .B(n22010), .Z(n22000) );
  AND U21894 ( .A(n22011), .B(n22012), .Z(n22010) );
  XOR U21895 ( .A(n22009), .B(n21128), .Z(n22012) );
  XNOR U21896 ( .A(p_input[1114]), .B(n22013), .Z(n21128) );
  AND U21897 ( .A(n474), .B(n22014), .Z(n22013) );
  XOR U21898 ( .A(p_input[1146]), .B(p_input[1114]), .Z(n22014) );
  XNOR U21899 ( .A(n21125), .B(n22009), .Z(n22011) );
  XOR U21900 ( .A(n22015), .B(n22016), .Z(n21125) );
  AND U21901 ( .A(n471), .B(n22017), .Z(n22016) );
  XOR U21902 ( .A(p_input[1082]), .B(p_input[1050]), .Z(n22017) );
  XOR U21903 ( .A(n22018), .B(n22019), .Z(n22009) );
  AND U21904 ( .A(n22020), .B(n22021), .Z(n22019) );
  XOR U21905 ( .A(n22018), .B(n21140), .Z(n22021) );
  XNOR U21906 ( .A(p_input[1113]), .B(n22022), .Z(n21140) );
  AND U21907 ( .A(n474), .B(n22023), .Z(n22022) );
  XOR U21908 ( .A(p_input[1145]), .B(p_input[1113]), .Z(n22023) );
  XNOR U21909 ( .A(n21137), .B(n22018), .Z(n22020) );
  XOR U21910 ( .A(n22024), .B(n22025), .Z(n21137) );
  AND U21911 ( .A(n471), .B(n22026), .Z(n22025) );
  XOR U21912 ( .A(p_input[1081]), .B(p_input[1049]), .Z(n22026) );
  XOR U21913 ( .A(n22027), .B(n22028), .Z(n22018) );
  AND U21914 ( .A(n22029), .B(n22030), .Z(n22028) );
  XOR U21915 ( .A(n22027), .B(n21152), .Z(n22030) );
  XNOR U21916 ( .A(p_input[1112]), .B(n22031), .Z(n21152) );
  AND U21917 ( .A(n474), .B(n22032), .Z(n22031) );
  XOR U21918 ( .A(p_input[1144]), .B(p_input[1112]), .Z(n22032) );
  XNOR U21919 ( .A(n21149), .B(n22027), .Z(n22029) );
  XOR U21920 ( .A(n22033), .B(n22034), .Z(n21149) );
  AND U21921 ( .A(n471), .B(n22035), .Z(n22034) );
  XOR U21922 ( .A(p_input[1080]), .B(p_input[1048]), .Z(n22035) );
  XOR U21923 ( .A(n22036), .B(n22037), .Z(n22027) );
  AND U21924 ( .A(n22038), .B(n22039), .Z(n22037) );
  XOR U21925 ( .A(n22036), .B(n21164), .Z(n22039) );
  XNOR U21926 ( .A(p_input[1111]), .B(n22040), .Z(n21164) );
  AND U21927 ( .A(n474), .B(n22041), .Z(n22040) );
  XOR U21928 ( .A(p_input[1143]), .B(p_input[1111]), .Z(n22041) );
  XNOR U21929 ( .A(n21161), .B(n22036), .Z(n22038) );
  XOR U21930 ( .A(n22042), .B(n22043), .Z(n21161) );
  AND U21931 ( .A(n471), .B(n22044), .Z(n22043) );
  XOR U21932 ( .A(p_input[1079]), .B(p_input[1047]), .Z(n22044) );
  XOR U21933 ( .A(n22045), .B(n22046), .Z(n22036) );
  AND U21934 ( .A(n22047), .B(n22048), .Z(n22046) );
  XOR U21935 ( .A(n22045), .B(n21176), .Z(n22048) );
  XNOR U21936 ( .A(p_input[1110]), .B(n22049), .Z(n21176) );
  AND U21937 ( .A(n474), .B(n22050), .Z(n22049) );
  XOR U21938 ( .A(p_input[1142]), .B(p_input[1110]), .Z(n22050) );
  XNOR U21939 ( .A(n21173), .B(n22045), .Z(n22047) );
  XOR U21940 ( .A(n22051), .B(n22052), .Z(n21173) );
  AND U21941 ( .A(n471), .B(n22053), .Z(n22052) );
  XOR U21942 ( .A(p_input[1078]), .B(p_input[1046]), .Z(n22053) );
  XOR U21943 ( .A(n22054), .B(n22055), .Z(n22045) );
  AND U21944 ( .A(n22056), .B(n22057), .Z(n22055) );
  XOR U21945 ( .A(n22054), .B(n21188), .Z(n22057) );
  XNOR U21946 ( .A(p_input[1109]), .B(n22058), .Z(n21188) );
  AND U21947 ( .A(n474), .B(n22059), .Z(n22058) );
  XOR U21948 ( .A(p_input[1141]), .B(p_input[1109]), .Z(n22059) );
  XNOR U21949 ( .A(n21185), .B(n22054), .Z(n22056) );
  XOR U21950 ( .A(n22060), .B(n22061), .Z(n21185) );
  AND U21951 ( .A(n471), .B(n22062), .Z(n22061) );
  XOR U21952 ( .A(p_input[1077]), .B(p_input[1045]), .Z(n22062) );
  XOR U21953 ( .A(n22063), .B(n22064), .Z(n22054) );
  AND U21954 ( .A(n22065), .B(n22066), .Z(n22064) );
  XOR U21955 ( .A(n22063), .B(n21200), .Z(n22066) );
  XNOR U21956 ( .A(p_input[1108]), .B(n22067), .Z(n21200) );
  AND U21957 ( .A(n474), .B(n22068), .Z(n22067) );
  XOR U21958 ( .A(p_input[1140]), .B(p_input[1108]), .Z(n22068) );
  XNOR U21959 ( .A(n21197), .B(n22063), .Z(n22065) );
  XOR U21960 ( .A(n22069), .B(n22070), .Z(n21197) );
  AND U21961 ( .A(n471), .B(n22071), .Z(n22070) );
  XOR U21962 ( .A(p_input[1076]), .B(p_input[1044]), .Z(n22071) );
  XOR U21963 ( .A(n22072), .B(n22073), .Z(n22063) );
  AND U21964 ( .A(n22074), .B(n22075), .Z(n22073) );
  XOR U21965 ( .A(n22072), .B(n21212), .Z(n22075) );
  XNOR U21966 ( .A(p_input[1107]), .B(n22076), .Z(n21212) );
  AND U21967 ( .A(n474), .B(n22077), .Z(n22076) );
  XOR U21968 ( .A(p_input[1139]), .B(p_input[1107]), .Z(n22077) );
  XNOR U21969 ( .A(n21209), .B(n22072), .Z(n22074) );
  XOR U21970 ( .A(n22078), .B(n22079), .Z(n21209) );
  AND U21971 ( .A(n471), .B(n22080), .Z(n22079) );
  XOR U21972 ( .A(p_input[1075]), .B(p_input[1043]), .Z(n22080) );
  XOR U21973 ( .A(n22081), .B(n22082), .Z(n22072) );
  AND U21974 ( .A(n22083), .B(n22084), .Z(n22082) );
  XOR U21975 ( .A(n22081), .B(n21224), .Z(n22084) );
  XNOR U21976 ( .A(p_input[1106]), .B(n22085), .Z(n21224) );
  AND U21977 ( .A(n474), .B(n22086), .Z(n22085) );
  XOR U21978 ( .A(p_input[1138]), .B(p_input[1106]), .Z(n22086) );
  XNOR U21979 ( .A(n21221), .B(n22081), .Z(n22083) );
  XOR U21980 ( .A(n22087), .B(n22088), .Z(n21221) );
  AND U21981 ( .A(n471), .B(n22089), .Z(n22088) );
  XOR U21982 ( .A(p_input[1074]), .B(p_input[1042]), .Z(n22089) );
  XOR U21983 ( .A(n22090), .B(n22091), .Z(n22081) );
  AND U21984 ( .A(n22092), .B(n22093), .Z(n22091) );
  XOR U21985 ( .A(n22090), .B(n21236), .Z(n22093) );
  XNOR U21986 ( .A(p_input[1105]), .B(n22094), .Z(n21236) );
  AND U21987 ( .A(n474), .B(n22095), .Z(n22094) );
  XOR U21988 ( .A(p_input[1137]), .B(p_input[1105]), .Z(n22095) );
  XNOR U21989 ( .A(n21233), .B(n22090), .Z(n22092) );
  XOR U21990 ( .A(n22096), .B(n22097), .Z(n21233) );
  AND U21991 ( .A(n471), .B(n22098), .Z(n22097) );
  XOR U21992 ( .A(p_input[1073]), .B(p_input[1041]), .Z(n22098) );
  XOR U21993 ( .A(n22099), .B(n22100), .Z(n22090) );
  AND U21994 ( .A(n22101), .B(n22102), .Z(n22100) );
  XOR U21995 ( .A(n22099), .B(n21248), .Z(n22102) );
  XNOR U21996 ( .A(p_input[1104]), .B(n22103), .Z(n21248) );
  AND U21997 ( .A(n474), .B(n22104), .Z(n22103) );
  XOR U21998 ( .A(p_input[1136]), .B(p_input[1104]), .Z(n22104) );
  XNOR U21999 ( .A(n21245), .B(n22099), .Z(n22101) );
  XOR U22000 ( .A(n22105), .B(n22106), .Z(n21245) );
  AND U22001 ( .A(n471), .B(n22107), .Z(n22106) );
  XOR U22002 ( .A(p_input[1072]), .B(p_input[1040]), .Z(n22107) );
  XOR U22003 ( .A(n22108), .B(n22109), .Z(n22099) );
  AND U22004 ( .A(n22110), .B(n22111), .Z(n22109) );
  XOR U22005 ( .A(n22108), .B(n21260), .Z(n22111) );
  XNOR U22006 ( .A(p_input[1103]), .B(n22112), .Z(n21260) );
  AND U22007 ( .A(n474), .B(n22113), .Z(n22112) );
  XOR U22008 ( .A(p_input[1135]), .B(p_input[1103]), .Z(n22113) );
  XNOR U22009 ( .A(n21257), .B(n22108), .Z(n22110) );
  XOR U22010 ( .A(n22114), .B(n22115), .Z(n21257) );
  AND U22011 ( .A(n471), .B(n22116), .Z(n22115) );
  XOR U22012 ( .A(p_input[1071]), .B(p_input[1039]), .Z(n22116) );
  XOR U22013 ( .A(n22117), .B(n22118), .Z(n22108) );
  AND U22014 ( .A(n22119), .B(n22120), .Z(n22118) );
  XOR U22015 ( .A(n22117), .B(n21272), .Z(n22120) );
  XNOR U22016 ( .A(p_input[1102]), .B(n22121), .Z(n21272) );
  AND U22017 ( .A(n474), .B(n22122), .Z(n22121) );
  XOR U22018 ( .A(p_input[1134]), .B(p_input[1102]), .Z(n22122) );
  XNOR U22019 ( .A(n21269), .B(n22117), .Z(n22119) );
  XOR U22020 ( .A(n22123), .B(n22124), .Z(n21269) );
  AND U22021 ( .A(n471), .B(n22125), .Z(n22124) );
  XOR U22022 ( .A(p_input[1070]), .B(p_input[1038]), .Z(n22125) );
  XOR U22023 ( .A(n22126), .B(n22127), .Z(n22117) );
  AND U22024 ( .A(n22128), .B(n22129), .Z(n22127) );
  XOR U22025 ( .A(n22126), .B(n21284), .Z(n22129) );
  XNOR U22026 ( .A(p_input[1101]), .B(n22130), .Z(n21284) );
  AND U22027 ( .A(n474), .B(n22131), .Z(n22130) );
  XOR U22028 ( .A(p_input[1133]), .B(p_input[1101]), .Z(n22131) );
  XNOR U22029 ( .A(n21281), .B(n22126), .Z(n22128) );
  XOR U22030 ( .A(n22132), .B(n22133), .Z(n21281) );
  AND U22031 ( .A(n471), .B(n22134), .Z(n22133) );
  XOR U22032 ( .A(p_input[1069]), .B(p_input[1037]), .Z(n22134) );
  XOR U22033 ( .A(n22135), .B(n22136), .Z(n22126) );
  AND U22034 ( .A(n22137), .B(n22138), .Z(n22136) );
  XOR U22035 ( .A(n22135), .B(n21296), .Z(n22138) );
  XNOR U22036 ( .A(p_input[1100]), .B(n22139), .Z(n21296) );
  AND U22037 ( .A(n474), .B(n22140), .Z(n22139) );
  XOR U22038 ( .A(p_input[1132]), .B(p_input[1100]), .Z(n22140) );
  XNOR U22039 ( .A(n21293), .B(n22135), .Z(n22137) );
  XOR U22040 ( .A(n22141), .B(n22142), .Z(n21293) );
  AND U22041 ( .A(n471), .B(n22143), .Z(n22142) );
  XOR U22042 ( .A(p_input[1068]), .B(p_input[1036]), .Z(n22143) );
  XOR U22043 ( .A(n22144), .B(n22145), .Z(n22135) );
  AND U22044 ( .A(n22146), .B(n22147), .Z(n22145) );
  XOR U22045 ( .A(n22144), .B(n21308), .Z(n22147) );
  XNOR U22046 ( .A(p_input[1099]), .B(n22148), .Z(n21308) );
  AND U22047 ( .A(n474), .B(n22149), .Z(n22148) );
  XOR U22048 ( .A(p_input[1131]), .B(p_input[1099]), .Z(n22149) );
  XNOR U22049 ( .A(n21305), .B(n22144), .Z(n22146) );
  XOR U22050 ( .A(n22150), .B(n22151), .Z(n21305) );
  AND U22051 ( .A(n471), .B(n22152), .Z(n22151) );
  XOR U22052 ( .A(p_input[1067]), .B(p_input[1035]), .Z(n22152) );
  XOR U22053 ( .A(n22153), .B(n22154), .Z(n22144) );
  AND U22054 ( .A(n22155), .B(n22156), .Z(n22154) );
  XOR U22055 ( .A(n22153), .B(n21320), .Z(n22156) );
  XNOR U22056 ( .A(p_input[1098]), .B(n22157), .Z(n21320) );
  AND U22057 ( .A(n474), .B(n22158), .Z(n22157) );
  XOR U22058 ( .A(p_input[1130]), .B(p_input[1098]), .Z(n22158) );
  XNOR U22059 ( .A(n21317), .B(n22153), .Z(n22155) );
  XOR U22060 ( .A(n22159), .B(n22160), .Z(n21317) );
  AND U22061 ( .A(n471), .B(n22161), .Z(n22160) );
  XOR U22062 ( .A(p_input[1066]), .B(p_input[1034]), .Z(n22161) );
  XOR U22063 ( .A(n22162), .B(n22163), .Z(n22153) );
  AND U22064 ( .A(n22164), .B(n22165), .Z(n22163) );
  XOR U22065 ( .A(n22162), .B(n21332), .Z(n22165) );
  XNOR U22066 ( .A(p_input[1097]), .B(n22166), .Z(n21332) );
  AND U22067 ( .A(n474), .B(n22167), .Z(n22166) );
  XOR U22068 ( .A(p_input[1129]), .B(p_input[1097]), .Z(n22167) );
  XNOR U22069 ( .A(n21329), .B(n22162), .Z(n22164) );
  XOR U22070 ( .A(n22168), .B(n22169), .Z(n21329) );
  AND U22071 ( .A(n471), .B(n22170), .Z(n22169) );
  XOR U22072 ( .A(p_input[1065]), .B(p_input[1033]), .Z(n22170) );
  XOR U22073 ( .A(n22171), .B(n22172), .Z(n22162) );
  AND U22074 ( .A(n22173), .B(n22174), .Z(n22172) );
  XOR U22075 ( .A(n22171), .B(n21344), .Z(n22174) );
  XNOR U22076 ( .A(p_input[1096]), .B(n22175), .Z(n21344) );
  AND U22077 ( .A(n474), .B(n22176), .Z(n22175) );
  XOR U22078 ( .A(p_input[1128]), .B(p_input[1096]), .Z(n22176) );
  XNOR U22079 ( .A(n21341), .B(n22171), .Z(n22173) );
  XOR U22080 ( .A(n22177), .B(n22178), .Z(n21341) );
  AND U22081 ( .A(n471), .B(n22179), .Z(n22178) );
  XOR U22082 ( .A(p_input[1064]), .B(p_input[1032]), .Z(n22179) );
  XOR U22083 ( .A(n22180), .B(n22181), .Z(n22171) );
  AND U22084 ( .A(n22182), .B(n22183), .Z(n22181) );
  XOR U22085 ( .A(n22180), .B(n21356), .Z(n22183) );
  XNOR U22086 ( .A(p_input[1095]), .B(n22184), .Z(n21356) );
  AND U22087 ( .A(n474), .B(n22185), .Z(n22184) );
  XOR U22088 ( .A(p_input[1127]), .B(p_input[1095]), .Z(n22185) );
  XNOR U22089 ( .A(n21353), .B(n22180), .Z(n22182) );
  XOR U22090 ( .A(n22186), .B(n22187), .Z(n21353) );
  AND U22091 ( .A(n471), .B(n22188), .Z(n22187) );
  XOR U22092 ( .A(p_input[1063]), .B(p_input[1031]), .Z(n22188) );
  XOR U22093 ( .A(n22189), .B(n22190), .Z(n22180) );
  AND U22094 ( .A(n22191), .B(n22192), .Z(n22190) );
  XOR U22095 ( .A(n22189), .B(n21368), .Z(n22192) );
  XNOR U22096 ( .A(p_input[1094]), .B(n22193), .Z(n21368) );
  AND U22097 ( .A(n474), .B(n22194), .Z(n22193) );
  XOR U22098 ( .A(p_input[1126]), .B(p_input[1094]), .Z(n22194) );
  XNOR U22099 ( .A(n21365), .B(n22189), .Z(n22191) );
  XOR U22100 ( .A(n22195), .B(n22196), .Z(n21365) );
  AND U22101 ( .A(n471), .B(n22197), .Z(n22196) );
  XOR U22102 ( .A(p_input[1062]), .B(p_input[1030]), .Z(n22197) );
  XOR U22103 ( .A(n22198), .B(n22199), .Z(n22189) );
  AND U22104 ( .A(n22200), .B(n22201), .Z(n22199) );
  XOR U22105 ( .A(n22198), .B(n21380), .Z(n22201) );
  XNOR U22106 ( .A(p_input[1093]), .B(n22202), .Z(n21380) );
  AND U22107 ( .A(n474), .B(n22203), .Z(n22202) );
  XOR U22108 ( .A(p_input[1125]), .B(p_input[1093]), .Z(n22203) );
  XNOR U22109 ( .A(n21377), .B(n22198), .Z(n22200) );
  XOR U22110 ( .A(n22204), .B(n22205), .Z(n21377) );
  AND U22111 ( .A(n471), .B(n22206), .Z(n22205) );
  XOR U22112 ( .A(p_input[1061]), .B(p_input[1029]), .Z(n22206) );
  XOR U22113 ( .A(n22207), .B(n22208), .Z(n22198) );
  AND U22114 ( .A(n22209), .B(n22210), .Z(n22208) );
  XOR U22115 ( .A(n22207), .B(n21392), .Z(n22210) );
  XNOR U22116 ( .A(p_input[1092]), .B(n22211), .Z(n21392) );
  AND U22117 ( .A(n474), .B(n22212), .Z(n22211) );
  XOR U22118 ( .A(p_input[1124]), .B(p_input[1092]), .Z(n22212) );
  XNOR U22119 ( .A(n21389), .B(n22207), .Z(n22209) );
  XOR U22120 ( .A(n22213), .B(n22214), .Z(n21389) );
  AND U22121 ( .A(n471), .B(n22215), .Z(n22214) );
  XOR U22122 ( .A(p_input[1060]), .B(p_input[1028]), .Z(n22215) );
  XOR U22123 ( .A(n22216), .B(n22217), .Z(n22207) );
  AND U22124 ( .A(n22218), .B(n22219), .Z(n22217) );
  XOR U22125 ( .A(n22216), .B(n21404), .Z(n22219) );
  XNOR U22126 ( .A(p_input[1091]), .B(n22220), .Z(n21404) );
  AND U22127 ( .A(n474), .B(n22221), .Z(n22220) );
  XOR U22128 ( .A(p_input[1123]), .B(p_input[1091]), .Z(n22221) );
  XNOR U22129 ( .A(n21401), .B(n22216), .Z(n22218) );
  XOR U22130 ( .A(n22222), .B(n22223), .Z(n21401) );
  AND U22131 ( .A(n471), .B(n22224), .Z(n22223) );
  XOR U22132 ( .A(p_input[1059]), .B(p_input[1027]), .Z(n22224) );
  XOR U22133 ( .A(n22225), .B(n22226), .Z(n22216) );
  AND U22134 ( .A(n22227), .B(n22228), .Z(n22226) );
  XOR U22135 ( .A(n21416), .B(n22225), .Z(n22228) );
  XNOR U22136 ( .A(p_input[1090]), .B(n22229), .Z(n21416) );
  AND U22137 ( .A(n474), .B(n22230), .Z(n22229) );
  XOR U22138 ( .A(p_input[1122]), .B(p_input[1090]), .Z(n22230) );
  XNOR U22139 ( .A(n22225), .B(n21413), .Z(n22227) );
  XOR U22140 ( .A(n22231), .B(n22232), .Z(n21413) );
  AND U22141 ( .A(n471), .B(n22233), .Z(n22232) );
  XOR U22142 ( .A(p_input[1058]), .B(p_input[1026]), .Z(n22233) );
  XOR U22143 ( .A(n22234), .B(n22235), .Z(n22225) );
  AND U22144 ( .A(n22236), .B(n22237), .Z(n22235) );
  XNOR U22145 ( .A(n22238), .B(n21429), .Z(n22237) );
  XNOR U22146 ( .A(p_input[1089]), .B(n22239), .Z(n21429) );
  AND U22147 ( .A(n474), .B(n22240), .Z(n22239) );
  XNOR U22148 ( .A(p_input[1121]), .B(n22241), .Z(n22240) );
  IV U22149 ( .A(p_input[1089]), .Z(n22241) );
  XNOR U22150 ( .A(n21426), .B(n22234), .Z(n22236) );
  XNOR U22151 ( .A(p_input[1025]), .B(n22242), .Z(n21426) );
  AND U22152 ( .A(n471), .B(n22243), .Z(n22242) );
  XOR U22153 ( .A(p_input[1057]), .B(p_input[1025]), .Z(n22243) );
  IV U22154 ( .A(n22238), .Z(n22234) );
  AND U22155 ( .A(n21964), .B(n21967), .Z(n22238) );
  XOR U22156 ( .A(p_input[1088]), .B(n22244), .Z(n21967) );
  AND U22157 ( .A(n474), .B(n22245), .Z(n22244) );
  XOR U22158 ( .A(p_input[1120]), .B(p_input[1088]), .Z(n22245) );
  XOR U22159 ( .A(n22246), .B(n22247), .Z(n474) );
  AND U22160 ( .A(n22248), .B(n22249), .Z(n22247) );
  XNOR U22161 ( .A(p_input[1151]), .B(n22246), .Z(n22249) );
  XOR U22162 ( .A(n22246), .B(p_input[1119]), .Z(n22248) );
  XOR U22163 ( .A(n22250), .B(n22251), .Z(n22246) );
  AND U22164 ( .A(n22252), .B(n22253), .Z(n22251) );
  XNOR U22165 ( .A(p_input[1150]), .B(n22250), .Z(n22253) );
  XOR U22166 ( .A(n22250), .B(p_input[1118]), .Z(n22252) );
  XOR U22167 ( .A(n22254), .B(n22255), .Z(n22250) );
  AND U22168 ( .A(n22256), .B(n22257), .Z(n22255) );
  XNOR U22169 ( .A(p_input[1149]), .B(n22254), .Z(n22257) );
  XOR U22170 ( .A(n22254), .B(p_input[1117]), .Z(n22256) );
  XOR U22171 ( .A(n22258), .B(n22259), .Z(n22254) );
  AND U22172 ( .A(n22260), .B(n22261), .Z(n22259) );
  XNOR U22173 ( .A(p_input[1148]), .B(n22258), .Z(n22261) );
  XOR U22174 ( .A(n22258), .B(p_input[1116]), .Z(n22260) );
  XOR U22175 ( .A(n22262), .B(n22263), .Z(n22258) );
  AND U22176 ( .A(n22264), .B(n22265), .Z(n22263) );
  XNOR U22177 ( .A(p_input[1147]), .B(n22262), .Z(n22265) );
  XOR U22178 ( .A(n22262), .B(p_input[1115]), .Z(n22264) );
  XOR U22179 ( .A(n22266), .B(n22267), .Z(n22262) );
  AND U22180 ( .A(n22268), .B(n22269), .Z(n22267) );
  XNOR U22181 ( .A(p_input[1146]), .B(n22266), .Z(n22269) );
  XOR U22182 ( .A(n22266), .B(p_input[1114]), .Z(n22268) );
  XOR U22183 ( .A(n22270), .B(n22271), .Z(n22266) );
  AND U22184 ( .A(n22272), .B(n22273), .Z(n22271) );
  XNOR U22185 ( .A(p_input[1145]), .B(n22270), .Z(n22273) );
  XOR U22186 ( .A(n22270), .B(p_input[1113]), .Z(n22272) );
  XOR U22187 ( .A(n22274), .B(n22275), .Z(n22270) );
  AND U22188 ( .A(n22276), .B(n22277), .Z(n22275) );
  XNOR U22189 ( .A(p_input[1144]), .B(n22274), .Z(n22277) );
  XOR U22190 ( .A(n22274), .B(p_input[1112]), .Z(n22276) );
  XOR U22191 ( .A(n22278), .B(n22279), .Z(n22274) );
  AND U22192 ( .A(n22280), .B(n22281), .Z(n22279) );
  XNOR U22193 ( .A(p_input[1143]), .B(n22278), .Z(n22281) );
  XOR U22194 ( .A(n22278), .B(p_input[1111]), .Z(n22280) );
  XOR U22195 ( .A(n22282), .B(n22283), .Z(n22278) );
  AND U22196 ( .A(n22284), .B(n22285), .Z(n22283) );
  XNOR U22197 ( .A(p_input[1142]), .B(n22282), .Z(n22285) );
  XOR U22198 ( .A(n22282), .B(p_input[1110]), .Z(n22284) );
  XOR U22199 ( .A(n22286), .B(n22287), .Z(n22282) );
  AND U22200 ( .A(n22288), .B(n22289), .Z(n22287) );
  XNOR U22201 ( .A(p_input[1141]), .B(n22286), .Z(n22289) );
  XOR U22202 ( .A(n22286), .B(p_input[1109]), .Z(n22288) );
  XOR U22203 ( .A(n22290), .B(n22291), .Z(n22286) );
  AND U22204 ( .A(n22292), .B(n22293), .Z(n22291) );
  XNOR U22205 ( .A(p_input[1140]), .B(n22290), .Z(n22293) );
  XOR U22206 ( .A(n22290), .B(p_input[1108]), .Z(n22292) );
  XOR U22207 ( .A(n22294), .B(n22295), .Z(n22290) );
  AND U22208 ( .A(n22296), .B(n22297), .Z(n22295) );
  XNOR U22209 ( .A(p_input[1139]), .B(n22294), .Z(n22297) );
  XOR U22210 ( .A(n22294), .B(p_input[1107]), .Z(n22296) );
  XOR U22211 ( .A(n22298), .B(n22299), .Z(n22294) );
  AND U22212 ( .A(n22300), .B(n22301), .Z(n22299) );
  XNOR U22213 ( .A(p_input[1138]), .B(n22298), .Z(n22301) );
  XOR U22214 ( .A(n22298), .B(p_input[1106]), .Z(n22300) );
  XOR U22215 ( .A(n22302), .B(n22303), .Z(n22298) );
  AND U22216 ( .A(n22304), .B(n22305), .Z(n22303) );
  XNOR U22217 ( .A(p_input[1137]), .B(n22302), .Z(n22305) );
  XOR U22218 ( .A(n22302), .B(p_input[1105]), .Z(n22304) );
  XOR U22219 ( .A(n22306), .B(n22307), .Z(n22302) );
  AND U22220 ( .A(n22308), .B(n22309), .Z(n22307) );
  XNOR U22221 ( .A(p_input[1136]), .B(n22306), .Z(n22309) );
  XOR U22222 ( .A(n22306), .B(p_input[1104]), .Z(n22308) );
  XOR U22223 ( .A(n22310), .B(n22311), .Z(n22306) );
  AND U22224 ( .A(n22312), .B(n22313), .Z(n22311) );
  XNOR U22225 ( .A(p_input[1135]), .B(n22310), .Z(n22313) );
  XOR U22226 ( .A(n22310), .B(p_input[1103]), .Z(n22312) );
  XOR U22227 ( .A(n22314), .B(n22315), .Z(n22310) );
  AND U22228 ( .A(n22316), .B(n22317), .Z(n22315) );
  XNOR U22229 ( .A(p_input[1134]), .B(n22314), .Z(n22317) );
  XOR U22230 ( .A(n22314), .B(p_input[1102]), .Z(n22316) );
  XOR U22231 ( .A(n22318), .B(n22319), .Z(n22314) );
  AND U22232 ( .A(n22320), .B(n22321), .Z(n22319) );
  XNOR U22233 ( .A(p_input[1133]), .B(n22318), .Z(n22321) );
  XOR U22234 ( .A(n22318), .B(p_input[1101]), .Z(n22320) );
  XOR U22235 ( .A(n22322), .B(n22323), .Z(n22318) );
  AND U22236 ( .A(n22324), .B(n22325), .Z(n22323) );
  XNOR U22237 ( .A(p_input[1132]), .B(n22322), .Z(n22325) );
  XOR U22238 ( .A(n22322), .B(p_input[1100]), .Z(n22324) );
  XOR U22239 ( .A(n22326), .B(n22327), .Z(n22322) );
  AND U22240 ( .A(n22328), .B(n22329), .Z(n22327) );
  XNOR U22241 ( .A(p_input[1131]), .B(n22326), .Z(n22329) );
  XOR U22242 ( .A(n22326), .B(p_input[1099]), .Z(n22328) );
  XOR U22243 ( .A(n22330), .B(n22331), .Z(n22326) );
  AND U22244 ( .A(n22332), .B(n22333), .Z(n22331) );
  XNOR U22245 ( .A(p_input[1130]), .B(n22330), .Z(n22333) );
  XOR U22246 ( .A(n22330), .B(p_input[1098]), .Z(n22332) );
  XOR U22247 ( .A(n22334), .B(n22335), .Z(n22330) );
  AND U22248 ( .A(n22336), .B(n22337), .Z(n22335) );
  XNOR U22249 ( .A(p_input[1129]), .B(n22334), .Z(n22337) );
  XOR U22250 ( .A(n22334), .B(p_input[1097]), .Z(n22336) );
  XOR U22251 ( .A(n22338), .B(n22339), .Z(n22334) );
  AND U22252 ( .A(n22340), .B(n22341), .Z(n22339) );
  XNOR U22253 ( .A(p_input[1128]), .B(n22338), .Z(n22341) );
  XOR U22254 ( .A(n22338), .B(p_input[1096]), .Z(n22340) );
  XOR U22255 ( .A(n22342), .B(n22343), .Z(n22338) );
  AND U22256 ( .A(n22344), .B(n22345), .Z(n22343) );
  XNOR U22257 ( .A(p_input[1127]), .B(n22342), .Z(n22345) );
  XOR U22258 ( .A(n22342), .B(p_input[1095]), .Z(n22344) );
  XOR U22259 ( .A(n22346), .B(n22347), .Z(n22342) );
  AND U22260 ( .A(n22348), .B(n22349), .Z(n22347) );
  XNOR U22261 ( .A(p_input[1126]), .B(n22346), .Z(n22349) );
  XOR U22262 ( .A(n22346), .B(p_input[1094]), .Z(n22348) );
  XOR U22263 ( .A(n22350), .B(n22351), .Z(n22346) );
  AND U22264 ( .A(n22352), .B(n22353), .Z(n22351) );
  XNOR U22265 ( .A(p_input[1125]), .B(n22350), .Z(n22353) );
  XOR U22266 ( .A(n22350), .B(p_input[1093]), .Z(n22352) );
  XOR U22267 ( .A(n22354), .B(n22355), .Z(n22350) );
  AND U22268 ( .A(n22356), .B(n22357), .Z(n22355) );
  XNOR U22269 ( .A(p_input[1124]), .B(n22354), .Z(n22357) );
  XOR U22270 ( .A(n22354), .B(p_input[1092]), .Z(n22356) );
  XOR U22271 ( .A(n22358), .B(n22359), .Z(n22354) );
  AND U22272 ( .A(n22360), .B(n22361), .Z(n22359) );
  XNOR U22273 ( .A(p_input[1123]), .B(n22358), .Z(n22361) );
  XOR U22274 ( .A(n22358), .B(p_input[1091]), .Z(n22360) );
  XOR U22275 ( .A(n22362), .B(n22363), .Z(n22358) );
  AND U22276 ( .A(n22364), .B(n22365), .Z(n22363) );
  XNOR U22277 ( .A(p_input[1122]), .B(n22362), .Z(n22365) );
  XOR U22278 ( .A(n22362), .B(p_input[1090]), .Z(n22364) );
  XNOR U22279 ( .A(n22366), .B(n22367), .Z(n22362) );
  AND U22280 ( .A(n22368), .B(n22369), .Z(n22367) );
  XOR U22281 ( .A(p_input[1121]), .B(n22366), .Z(n22369) );
  XNOR U22282 ( .A(p_input[1089]), .B(n22366), .Z(n22368) );
  AND U22283 ( .A(p_input[1120]), .B(n22370), .Z(n22366) );
  IV U22284 ( .A(p_input[1088]), .Z(n22370) );
  XNOR U22285 ( .A(p_input[1024]), .B(n22371), .Z(n21964) );
  AND U22286 ( .A(n471), .B(n22372), .Z(n22371) );
  XOR U22287 ( .A(p_input[1056]), .B(p_input[1024]), .Z(n22372) );
  XOR U22288 ( .A(n22373), .B(n22374), .Z(n471) );
  AND U22289 ( .A(n22375), .B(n22376), .Z(n22374) );
  XNOR U22290 ( .A(p_input[1087]), .B(n22373), .Z(n22376) );
  XOR U22291 ( .A(n22373), .B(p_input[1055]), .Z(n22375) );
  XOR U22292 ( .A(n22377), .B(n22378), .Z(n22373) );
  AND U22293 ( .A(n22379), .B(n22380), .Z(n22378) );
  XNOR U22294 ( .A(p_input[1086]), .B(n22377), .Z(n22380) );
  XNOR U22295 ( .A(n22377), .B(n21979), .Z(n22379) );
  IV U22296 ( .A(p_input[1054]), .Z(n21979) );
  XOR U22297 ( .A(n22381), .B(n22382), .Z(n22377) );
  AND U22298 ( .A(n22383), .B(n22384), .Z(n22382) );
  XNOR U22299 ( .A(p_input[1085]), .B(n22381), .Z(n22384) );
  XNOR U22300 ( .A(n22381), .B(n21988), .Z(n22383) );
  IV U22301 ( .A(p_input[1053]), .Z(n21988) );
  XOR U22302 ( .A(n22385), .B(n22386), .Z(n22381) );
  AND U22303 ( .A(n22387), .B(n22388), .Z(n22386) );
  XNOR U22304 ( .A(p_input[1084]), .B(n22385), .Z(n22388) );
  XNOR U22305 ( .A(n22385), .B(n21997), .Z(n22387) );
  IV U22306 ( .A(p_input[1052]), .Z(n21997) );
  XOR U22307 ( .A(n22389), .B(n22390), .Z(n22385) );
  AND U22308 ( .A(n22391), .B(n22392), .Z(n22390) );
  XNOR U22309 ( .A(p_input[1083]), .B(n22389), .Z(n22392) );
  XNOR U22310 ( .A(n22389), .B(n22006), .Z(n22391) );
  IV U22311 ( .A(p_input[1051]), .Z(n22006) );
  XOR U22312 ( .A(n22393), .B(n22394), .Z(n22389) );
  AND U22313 ( .A(n22395), .B(n22396), .Z(n22394) );
  XNOR U22314 ( .A(p_input[1082]), .B(n22393), .Z(n22396) );
  XNOR U22315 ( .A(n22393), .B(n22015), .Z(n22395) );
  IV U22316 ( .A(p_input[1050]), .Z(n22015) );
  XOR U22317 ( .A(n22397), .B(n22398), .Z(n22393) );
  AND U22318 ( .A(n22399), .B(n22400), .Z(n22398) );
  XNOR U22319 ( .A(p_input[1081]), .B(n22397), .Z(n22400) );
  XNOR U22320 ( .A(n22397), .B(n22024), .Z(n22399) );
  IV U22321 ( .A(p_input[1049]), .Z(n22024) );
  XOR U22322 ( .A(n22401), .B(n22402), .Z(n22397) );
  AND U22323 ( .A(n22403), .B(n22404), .Z(n22402) );
  XNOR U22324 ( .A(p_input[1080]), .B(n22401), .Z(n22404) );
  XNOR U22325 ( .A(n22401), .B(n22033), .Z(n22403) );
  IV U22326 ( .A(p_input[1048]), .Z(n22033) );
  XOR U22327 ( .A(n22405), .B(n22406), .Z(n22401) );
  AND U22328 ( .A(n22407), .B(n22408), .Z(n22406) );
  XNOR U22329 ( .A(p_input[1079]), .B(n22405), .Z(n22408) );
  XNOR U22330 ( .A(n22405), .B(n22042), .Z(n22407) );
  IV U22331 ( .A(p_input[1047]), .Z(n22042) );
  XOR U22332 ( .A(n22409), .B(n22410), .Z(n22405) );
  AND U22333 ( .A(n22411), .B(n22412), .Z(n22410) );
  XNOR U22334 ( .A(p_input[1078]), .B(n22409), .Z(n22412) );
  XNOR U22335 ( .A(n22409), .B(n22051), .Z(n22411) );
  IV U22336 ( .A(p_input[1046]), .Z(n22051) );
  XOR U22337 ( .A(n22413), .B(n22414), .Z(n22409) );
  AND U22338 ( .A(n22415), .B(n22416), .Z(n22414) );
  XNOR U22339 ( .A(p_input[1077]), .B(n22413), .Z(n22416) );
  XNOR U22340 ( .A(n22413), .B(n22060), .Z(n22415) );
  IV U22341 ( .A(p_input[1045]), .Z(n22060) );
  XOR U22342 ( .A(n22417), .B(n22418), .Z(n22413) );
  AND U22343 ( .A(n22419), .B(n22420), .Z(n22418) );
  XNOR U22344 ( .A(p_input[1076]), .B(n22417), .Z(n22420) );
  XNOR U22345 ( .A(n22417), .B(n22069), .Z(n22419) );
  IV U22346 ( .A(p_input[1044]), .Z(n22069) );
  XOR U22347 ( .A(n22421), .B(n22422), .Z(n22417) );
  AND U22348 ( .A(n22423), .B(n22424), .Z(n22422) );
  XNOR U22349 ( .A(p_input[1075]), .B(n22421), .Z(n22424) );
  XNOR U22350 ( .A(n22421), .B(n22078), .Z(n22423) );
  IV U22351 ( .A(p_input[1043]), .Z(n22078) );
  XOR U22352 ( .A(n22425), .B(n22426), .Z(n22421) );
  AND U22353 ( .A(n22427), .B(n22428), .Z(n22426) );
  XNOR U22354 ( .A(p_input[1074]), .B(n22425), .Z(n22428) );
  XNOR U22355 ( .A(n22425), .B(n22087), .Z(n22427) );
  IV U22356 ( .A(p_input[1042]), .Z(n22087) );
  XOR U22357 ( .A(n22429), .B(n22430), .Z(n22425) );
  AND U22358 ( .A(n22431), .B(n22432), .Z(n22430) );
  XNOR U22359 ( .A(p_input[1073]), .B(n22429), .Z(n22432) );
  XNOR U22360 ( .A(n22429), .B(n22096), .Z(n22431) );
  IV U22361 ( .A(p_input[1041]), .Z(n22096) );
  XOR U22362 ( .A(n22433), .B(n22434), .Z(n22429) );
  AND U22363 ( .A(n22435), .B(n22436), .Z(n22434) );
  XNOR U22364 ( .A(p_input[1072]), .B(n22433), .Z(n22436) );
  XNOR U22365 ( .A(n22433), .B(n22105), .Z(n22435) );
  IV U22366 ( .A(p_input[1040]), .Z(n22105) );
  XOR U22367 ( .A(n22437), .B(n22438), .Z(n22433) );
  AND U22368 ( .A(n22439), .B(n22440), .Z(n22438) );
  XNOR U22369 ( .A(p_input[1071]), .B(n22437), .Z(n22440) );
  XNOR U22370 ( .A(n22437), .B(n22114), .Z(n22439) );
  IV U22371 ( .A(p_input[1039]), .Z(n22114) );
  XOR U22372 ( .A(n22441), .B(n22442), .Z(n22437) );
  AND U22373 ( .A(n22443), .B(n22444), .Z(n22442) );
  XNOR U22374 ( .A(p_input[1070]), .B(n22441), .Z(n22444) );
  XNOR U22375 ( .A(n22441), .B(n22123), .Z(n22443) );
  IV U22376 ( .A(p_input[1038]), .Z(n22123) );
  XOR U22377 ( .A(n22445), .B(n22446), .Z(n22441) );
  AND U22378 ( .A(n22447), .B(n22448), .Z(n22446) );
  XNOR U22379 ( .A(p_input[1069]), .B(n22445), .Z(n22448) );
  XNOR U22380 ( .A(n22445), .B(n22132), .Z(n22447) );
  IV U22381 ( .A(p_input[1037]), .Z(n22132) );
  XOR U22382 ( .A(n22449), .B(n22450), .Z(n22445) );
  AND U22383 ( .A(n22451), .B(n22452), .Z(n22450) );
  XNOR U22384 ( .A(p_input[1068]), .B(n22449), .Z(n22452) );
  XNOR U22385 ( .A(n22449), .B(n22141), .Z(n22451) );
  IV U22386 ( .A(p_input[1036]), .Z(n22141) );
  XOR U22387 ( .A(n22453), .B(n22454), .Z(n22449) );
  AND U22388 ( .A(n22455), .B(n22456), .Z(n22454) );
  XNOR U22389 ( .A(p_input[1067]), .B(n22453), .Z(n22456) );
  XNOR U22390 ( .A(n22453), .B(n22150), .Z(n22455) );
  IV U22391 ( .A(p_input[1035]), .Z(n22150) );
  XOR U22392 ( .A(n22457), .B(n22458), .Z(n22453) );
  AND U22393 ( .A(n22459), .B(n22460), .Z(n22458) );
  XNOR U22394 ( .A(p_input[1066]), .B(n22457), .Z(n22460) );
  XNOR U22395 ( .A(n22457), .B(n22159), .Z(n22459) );
  IV U22396 ( .A(p_input[1034]), .Z(n22159) );
  XOR U22397 ( .A(n22461), .B(n22462), .Z(n22457) );
  AND U22398 ( .A(n22463), .B(n22464), .Z(n22462) );
  XNOR U22399 ( .A(p_input[1065]), .B(n22461), .Z(n22464) );
  XNOR U22400 ( .A(n22461), .B(n22168), .Z(n22463) );
  IV U22401 ( .A(p_input[1033]), .Z(n22168) );
  XOR U22402 ( .A(n22465), .B(n22466), .Z(n22461) );
  AND U22403 ( .A(n22467), .B(n22468), .Z(n22466) );
  XNOR U22404 ( .A(p_input[1064]), .B(n22465), .Z(n22468) );
  XNOR U22405 ( .A(n22465), .B(n22177), .Z(n22467) );
  IV U22406 ( .A(p_input[1032]), .Z(n22177) );
  XOR U22407 ( .A(n22469), .B(n22470), .Z(n22465) );
  AND U22408 ( .A(n22471), .B(n22472), .Z(n22470) );
  XNOR U22409 ( .A(p_input[1063]), .B(n22469), .Z(n22472) );
  XNOR U22410 ( .A(n22469), .B(n22186), .Z(n22471) );
  IV U22411 ( .A(p_input[1031]), .Z(n22186) );
  XOR U22412 ( .A(n22473), .B(n22474), .Z(n22469) );
  AND U22413 ( .A(n22475), .B(n22476), .Z(n22474) );
  XNOR U22414 ( .A(p_input[1062]), .B(n22473), .Z(n22476) );
  XNOR U22415 ( .A(n22473), .B(n22195), .Z(n22475) );
  IV U22416 ( .A(p_input[1030]), .Z(n22195) );
  XOR U22417 ( .A(n22477), .B(n22478), .Z(n22473) );
  AND U22418 ( .A(n22479), .B(n22480), .Z(n22478) );
  XNOR U22419 ( .A(p_input[1061]), .B(n22477), .Z(n22480) );
  XNOR U22420 ( .A(n22477), .B(n22204), .Z(n22479) );
  IV U22421 ( .A(p_input[1029]), .Z(n22204) );
  XOR U22422 ( .A(n22481), .B(n22482), .Z(n22477) );
  AND U22423 ( .A(n22483), .B(n22484), .Z(n22482) );
  XNOR U22424 ( .A(p_input[1060]), .B(n22481), .Z(n22484) );
  XNOR U22425 ( .A(n22481), .B(n22213), .Z(n22483) );
  IV U22426 ( .A(p_input[1028]), .Z(n22213) );
  XOR U22427 ( .A(n22485), .B(n22486), .Z(n22481) );
  AND U22428 ( .A(n22487), .B(n22488), .Z(n22486) );
  XNOR U22429 ( .A(p_input[1059]), .B(n22485), .Z(n22488) );
  XNOR U22430 ( .A(n22485), .B(n22222), .Z(n22487) );
  IV U22431 ( .A(p_input[1027]), .Z(n22222) );
  XOR U22432 ( .A(n22489), .B(n22490), .Z(n22485) );
  AND U22433 ( .A(n22491), .B(n22492), .Z(n22490) );
  XNOR U22434 ( .A(p_input[1058]), .B(n22489), .Z(n22492) );
  XNOR U22435 ( .A(n22489), .B(n22231), .Z(n22491) );
  IV U22436 ( .A(p_input[1026]), .Z(n22231) );
  XNOR U22437 ( .A(n22493), .B(n22494), .Z(n22489) );
  AND U22438 ( .A(n22495), .B(n22496), .Z(n22494) );
  XOR U22439 ( .A(p_input[1057]), .B(n22493), .Z(n22496) );
  XNOR U22440 ( .A(p_input[1025]), .B(n22493), .Z(n22495) );
  AND U22441 ( .A(p_input[1056]), .B(n22497), .Z(n22493) );
  IV U22442 ( .A(p_input[1024]), .Z(n22497) );
  XOR U22443 ( .A(n22498), .B(n22499), .Z(n15210) );
  AND U22444 ( .A(n619), .B(n22500), .Z(n22499) );
  XNOR U22445 ( .A(n22501), .B(n22498), .Z(n22500) );
  XOR U22446 ( .A(n22502), .B(n22503), .Z(n619) );
  AND U22447 ( .A(n22504), .B(n22505), .Z(n22503) );
  XOR U22448 ( .A(n22502), .B(n15225), .Z(n22505) );
  XOR U22449 ( .A(n22506), .B(n22507), .Z(n15225) );
  AND U22450 ( .A(n594), .B(n22508), .Z(n22507) );
  XOR U22451 ( .A(n22509), .B(n22506), .Z(n22508) );
  XNOR U22452 ( .A(n15222), .B(n22502), .Z(n22504) );
  XOR U22453 ( .A(n22510), .B(n22511), .Z(n15222) );
  AND U22454 ( .A(n591), .B(n22512), .Z(n22511) );
  XOR U22455 ( .A(n22513), .B(n22510), .Z(n22512) );
  XOR U22456 ( .A(n22514), .B(n22515), .Z(n22502) );
  AND U22457 ( .A(n22516), .B(n22517), .Z(n22515) );
  XOR U22458 ( .A(n22514), .B(n15237), .Z(n22517) );
  XOR U22459 ( .A(n22518), .B(n22519), .Z(n15237) );
  AND U22460 ( .A(n594), .B(n22520), .Z(n22519) );
  XOR U22461 ( .A(n22521), .B(n22518), .Z(n22520) );
  XNOR U22462 ( .A(n15234), .B(n22514), .Z(n22516) );
  XOR U22463 ( .A(n22522), .B(n22523), .Z(n15234) );
  AND U22464 ( .A(n591), .B(n22524), .Z(n22523) );
  XOR U22465 ( .A(n22525), .B(n22522), .Z(n22524) );
  XOR U22466 ( .A(n22526), .B(n22527), .Z(n22514) );
  AND U22467 ( .A(n22528), .B(n22529), .Z(n22527) );
  XOR U22468 ( .A(n22526), .B(n15249), .Z(n22529) );
  XOR U22469 ( .A(n22530), .B(n22531), .Z(n15249) );
  AND U22470 ( .A(n594), .B(n22532), .Z(n22531) );
  XOR U22471 ( .A(n22533), .B(n22530), .Z(n22532) );
  XNOR U22472 ( .A(n15246), .B(n22526), .Z(n22528) );
  XOR U22473 ( .A(n22534), .B(n22535), .Z(n15246) );
  AND U22474 ( .A(n591), .B(n22536), .Z(n22535) );
  XOR U22475 ( .A(n22537), .B(n22534), .Z(n22536) );
  XOR U22476 ( .A(n22538), .B(n22539), .Z(n22526) );
  AND U22477 ( .A(n22540), .B(n22541), .Z(n22539) );
  XOR U22478 ( .A(n22538), .B(n15261), .Z(n22541) );
  XOR U22479 ( .A(n22542), .B(n22543), .Z(n15261) );
  AND U22480 ( .A(n594), .B(n22544), .Z(n22543) );
  XOR U22481 ( .A(n22545), .B(n22542), .Z(n22544) );
  XNOR U22482 ( .A(n15258), .B(n22538), .Z(n22540) );
  XOR U22483 ( .A(n22546), .B(n22547), .Z(n15258) );
  AND U22484 ( .A(n591), .B(n22548), .Z(n22547) );
  XOR U22485 ( .A(n22549), .B(n22546), .Z(n22548) );
  XOR U22486 ( .A(n22550), .B(n22551), .Z(n22538) );
  AND U22487 ( .A(n22552), .B(n22553), .Z(n22551) );
  XOR U22488 ( .A(n22550), .B(n15273), .Z(n22553) );
  XOR U22489 ( .A(n22554), .B(n22555), .Z(n15273) );
  AND U22490 ( .A(n594), .B(n22556), .Z(n22555) );
  XOR U22491 ( .A(n22557), .B(n22554), .Z(n22556) );
  XNOR U22492 ( .A(n15270), .B(n22550), .Z(n22552) );
  XOR U22493 ( .A(n22558), .B(n22559), .Z(n15270) );
  AND U22494 ( .A(n591), .B(n22560), .Z(n22559) );
  XOR U22495 ( .A(n22561), .B(n22558), .Z(n22560) );
  XOR U22496 ( .A(n22562), .B(n22563), .Z(n22550) );
  AND U22497 ( .A(n22564), .B(n22565), .Z(n22563) );
  XOR U22498 ( .A(n22562), .B(n15285), .Z(n22565) );
  XOR U22499 ( .A(n22566), .B(n22567), .Z(n15285) );
  AND U22500 ( .A(n594), .B(n22568), .Z(n22567) );
  XOR U22501 ( .A(n22569), .B(n22566), .Z(n22568) );
  XNOR U22502 ( .A(n15282), .B(n22562), .Z(n22564) );
  XOR U22503 ( .A(n22570), .B(n22571), .Z(n15282) );
  AND U22504 ( .A(n591), .B(n22572), .Z(n22571) );
  XOR U22505 ( .A(n22573), .B(n22570), .Z(n22572) );
  XOR U22506 ( .A(n22574), .B(n22575), .Z(n22562) );
  AND U22507 ( .A(n22576), .B(n22577), .Z(n22575) );
  XOR U22508 ( .A(n22574), .B(n15297), .Z(n22577) );
  XOR U22509 ( .A(n22578), .B(n22579), .Z(n15297) );
  AND U22510 ( .A(n594), .B(n22580), .Z(n22579) );
  XOR U22511 ( .A(n22581), .B(n22578), .Z(n22580) );
  XNOR U22512 ( .A(n15294), .B(n22574), .Z(n22576) );
  XOR U22513 ( .A(n22582), .B(n22583), .Z(n15294) );
  AND U22514 ( .A(n591), .B(n22584), .Z(n22583) );
  XOR U22515 ( .A(n22585), .B(n22582), .Z(n22584) );
  XOR U22516 ( .A(n22586), .B(n22587), .Z(n22574) );
  AND U22517 ( .A(n22588), .B(n22589), .Z(n22587) );
  XOR U22518 ( .A(n22586), .B(n15309), .Z(n22589) );
  XOR U22519 ( .A(n22590), .B(n22591), .Z(n15309) );
  AND U22520 ( .A(n594), .B(n22592), .Z(n22591) );
  XOR U22521 ( .A(n22593), .B(n22590), .Z(n22592) );
  XNOR U22522 ( .A(n15306), .B(n22586), .Z(n22588) );
  XOR U22523 ( .A(n22594), .B(n22595), .Z(n15306) );
  AND U22524 ( .A(n591), .B(n22596), .Z(n22595) );
  XOR U22525 ( .A(n22597), .B(n22594), .Z(n22596) );
  XOR U22526 ( .A(n22598), .B(n22599), .Z(n22586) );
  AND U22527 ( .A(n22600), .B(n22601), .Z(n22599) );
  XOR U22528 ( .A(n22598), .B(n15321), .Z(n22601) );
  XOR U22529 ( .A(n22602), .B(n22603), .Z(n15321) );
  AND U22530 ( .A(n594), .B(n22604), .Z(n22603) );
  XOR U22531 ( .A(n22605), .B(n22602), .Z(n22604) );
  XNOR U22532 ( .A(n15318), .B(n22598), .Z(n22600) );
  XOR U22533 ( .A(n22606), .B(n22607), .Z(n15318) );
  AND U22534 ( .A(n591), .B(n22608), .Z(n22607) );
  XOR U22535 ( .A(n22609), .B(n22606), .Z(n22608) );
  XOR U22536 ( .A(n22610), .B(n22611), .Z(n22598) );
  AND U22537 ( .A(n22612), .B(n22613), .Z(n22611) );
  XOR U22538 ( .A(n22610), .B(n15333), .Z(n22613) );
  XOR U22539 ( .A(n22614), .B(n22615), .Z(n15333) );
  AND U22540 ( .A(n594), .B(n22616), .Z(n22615) );
  XOR U22541 ( .A(n22617), .B(n22614), .Z(n22616) );
  XNOR U22542 ( .A(n15330), .B(n22610), .Z(n22612) );
  XOR U22543 ( .A(n22618), .B(n22619), .Z(n15330) );
  AND U22544 ( .A(n591), .B(n22620), .Z(n22619) );
  XOR U22545 ( .A(n22621), .B(n22618), .Z(n22620) );
  XOR U22546 ( .A(n22622), .B(n22623), .Z(n22610) );
  AND U22547 ( .A(n22624), .B(n22625), .Z(n22623) );
  XOR U22548 ( .A(n22622), .B(n15345), .Z(n22625) );
  XOR U22549 ( .A(n22626), .B(n22627), .Z(n15345) );
  AND U22550 ( .A(n594), .B(n22628), .Z(n22627) );
  XOR U22551 ( .A(n22629), .B(n22626), .Z(n22628) );
  XNOR U22552 ( .A(n15342), .B(n22622), .Z(n22624) );
  XOR U22553 ( .A(n22630), .B(n22631), .Z(n15342) );
  AND U22554 ( .A(n591), .B(n22632), .Z(n22631) );
  XOR U22555 ( .A(n22633), .B(n22630), .Z(n22632) );
  XOR U22556 ( .A(n22634), .B(n22635), .Z(n22622) );
  AND U22557 ( .A(n22636), .B(n22637), .Z(n22635) );
  XOR U22558 ( .A(n22634), .B(n15357), .Z(n22637) );
  XOR U22559 ( .A(n22638), .B(n22639), .Z(n15357) );
  AND U22560 ( .A(n594), .B(n22640), .Z(n22639) );
  XOR U22561 ( .A(n22641), .B(n22638), .Z(n22640) );
  XNOR U22562 ( .A(n15354), .B(n22634), .Z(n22636) );
  XOR U22563 ( .A(n22642), .B(n22643), .Z(n15354) );
  AND U22564 ( .A(n591), .B(n22644), .Z(n22643) );
  XOR U22565 ( .A(n22645), .B(n22642), .Z(n22644) );
  XOR U22566 ( .A(n22646), .B(n22647), .Z(n22634) );
  AND U22567 ( .A(n22648), .B(n22649), .Z(n22647) );
  XOR U22568 ( .A(n22646), .B(n15369), .Z(n22649) );
  XOR U22569 ( .A(n22650), .B(n22651), .Z(n15369) );
  AND U22570 ( .A(n594), .B(n22652), .Z(n22651) );
  XOR U22571 ( .A(n22653), .B(n22650), .Z(n22652) );
  XNOR U22572 ( .A(n15366), .B(n22646), .Z(n22648) );
  XOR U22573 ( .A(n22654), .B(n22655), .Z(n15366) );
  AND U22574 ( .A(n591), .B(n22656), .Z(n22655) );
  XOR U22575 ( .A(n22657), .B(n22654), .Z(n22656) );
  XOR U22576 ( .A(n22658), .B(n22659), .Z(n22646) );
  AND U22577 ( .A(n22660), .B(n22661), .Z(n22659) );
  XOR U22578 ( .A(n22658), .B(n15381), .Z(n22661) );
  XOR U22579 ( .A(n22662), .B(n22663), .Z(n15381) );
  AND U22580 ( .A(n594), .B(n22664), .Z(n22663) );
  XOR U22581 ( .A(n22665), .B(n22662), .Z(n22664) );
  XNOR U22582 ( .A(n15378), .B(n22658), .Z(n22660) );
  XOR U22583 ( .A(n22666), .B(n22667), .Z(n15378) );
  AND U22584 ( .A(n591), .B(n22668), .Z(n22667) );
  XOR U22585 ( .A(n22669), .B(n22666), .Z(n22668) );
  XOR U22586 ( .A(n22670), .B(n22671), .Z(n22658) );
  AND U22587 ( .A(n22672), .B(n22673), .Z(n22671) );
  XOR U22588 ( .A(n22670), .B(n15393), .Z(n22673) );
  XOR U22589 ( .A(n22674), .B(n22675), .Z(n15393) );
  AND U22590 ( .A(n594), .B(n22676), .Z(n22675) );
  XOR U22591 ( .A(n22677), .B(n22674), .Z(n22676) );
  XNOR U22592 ( .A(n15390), .B(n22670), .Z(n22672) );
  XOR U22593 ( .A(n22678), .B(n22679), .Z(n15390) );
  AND U22594 ( .A(n591), .B(n22680), .Z(n22679) );
  XOR U22595 ( .A(n22681), .B(n22678), .Z(n22680) );
  XOR U22596 ( .A(n22682), .B(n22683), .Z(n22670) );
  AND U22597 ( .A(n22684), .B(n22685), .Z(n22683) );
  XOR U22598 ( .A(n22682), .B(n15405), .Z(n22685) );
  XOR U22599 ( .A(n22686), .B(n22687), .Z(n15405) );
  AND U22600 ( .A(n594), .B(n22688), .Z(n22687) );
  XOR U22601 ( .A(n22689), .B(n22686), .Z(n22688) );
  XNOR U22602 ( .A(n15402), .B(n22682), .Z(n22684) );
  XOR U22603 ( .A(n22690), .B(n22691), .Z(n15402) );
  AND U22604 ( .A(n591), .B(n22692), .Z(n22691) );
  XOR U22605 ( .A(n22693), .B(n22690), .Z(n22692) );
  XOR U22606 ( .A(n22694), .B(n22695), .Z(n22682) );
  AND U22607 ( .A(n22696), .B(n22697), .Z(n22695) );
  XOR U22608 ( .A(n22694), .B(n15417), .Z(n22697) );
  XOR U22609 ( .A(n22698), .B(n22699), .Z(n15417) );
  AND U22610 ( .A(n594), .B(n22700), .Z(n22699) );
  XOR U22611 ( .A(n22701), .B(n22698), .Z(n22700) );
  XNOR U22612 ( .A(n15414), .B(n22694), .Z(n22696) );
  XOR U22613 ( .A(n22702), .B(n22703), .Z(n15414) );
  AND U22614 ( .A(n591), .B(n22704), .Z(n22703) );
  XOR U22615 ( .A(n22705), .B(n22702), .Z(n22704) );
  XOR U22616 ( .A(n22706), .B(n22707), .Z(n22694) );
  AND U22617 ( .A(n22708), .B(n22709), .Z(n22707) );
  XOR U22618 ( .A(n22706), .B(n15429), .Z(n22709) );
  XOR U22619 ( .A(n22710), .B(n22711), .Z(n15429) );
  AND U22620 ( .A(n594), .B(n22712), .Z(n22711) );
  XOR U22621 ( .A(n22713), .B(n22710), .Z(n22712) );
  XNOR U22622 ( .A(n15426), .B(n22706), .Z(n22708) );
  XOR U22623 ( .A(n22714), .B(n22715), .Z(n15426) );
  AND U22624 ( .A(n591), .B(n22716), .Z(n22715) );
  XOR U22625 ( .A(n22717), .B(n22714), .Z(n22716) );
  XOR U22626 ( .A(n22718), .B(n22719), .Z(n22706) );
  AND U22627 ( .A(n22720), .B(n22721), .Z(n22719) );
  XOR U22628 ( .A(n22718), .B(n15441), .Z(n22721) );
  XOR U22629 ( .A(n22722), .B(n22723), .Z(n15441) );
  AND U22630 ( .A(n594), .B(n22724), .Z(n22723) );
  XOR U22631 ( .A(n22725), .B(n22722), .Z(n22724) );
  XNOR U22632 ( .A(n15438), .B(n22718), .Z(n22720) );
  XOR U22633 ( .A(n22726), .B(n22727), .Z(n15438) );
  AND U22634 ( .A(n591), .B(n22728), .Z(n22727) );
  XOR U22635 ( .A(n22729), .B(n22726), .Z(n22728) );
  XOR U22636 ( .A(n22730), .B(n22731), .Z(n22718) );
  AND U22637 ( .A(n22732), .B(n22733), .Z(n22731) );
  XOR U22638 ( .A(n22730), .B(n15453), .Z(n22733) );
  XOR U22639 ( .A(n22734), .B(n22735), .Z(n15453) );
  AND U22640 ( .A(n594), .B(n22736), .Z(n22735) );
  XOR U22641 ( .A(n22737), .B(n22734), .Z(n22736) );
  XNOR U22642 ( .A(n15450), .B(n22730), .Z(n22732) );
  XOR U22643 ( .A(n22738), .B(n22739), .Z(n15450) );
  AND U22644 ( .A(n591), .B(n22740), .Z(n22739) );
  XOR U22645 ( .A(n22741), .B(n22738), .Z(n22740) );
  XOR U22646 ( .A(n22742), .B(n22743), .Z(n22730) );
  AND U22647 ( .A(n22744), .B(n22745), .Z(n22743) );
  XOR U22648 ( .A(n22742), .B(n15465), .Z(n22745) );
  XOR U22649 ( .A(n22746), .B(n22747), .Z(n15465) );
  AND U22650 ( .A(n594), .B(n22748), .Z(n22747) );
  XOR U22651 ( .A(n22749), .B(n22746), .Z(n22748) );
  XNOR U22652 ( .A(n15462), .B(n22742), .Z(n22744) );
  XOR U22653 ( .A(n22750), .B(n22751), .Z(n15462) );
  AND U22654 ( .A(n591), .B(n22752), .Z(n22751) );
  XOR U22655 ( .A(n22753), .B(n22750), .Z(n22752) );
  XOR U22656 ( .A(n22754), .B(n22755), .Z(n22742) );
  AND U22657 ( .A(n22756), .B(n22757), .Z(n22755) );
  XOR U22658 ( .A(n22754), .B(n15477), .Z(n22757) );
  XOR U22659 ( .A(n22758), .B(n22759), .Z(n15477) );
  AND U22660 ( .A(n594), .B(n22760), .Z(n22759) );
  XOR U22661 ( .A(n22761), .B(n22758), .Z(n22760) );
  XNOR U22662 ( .A(n15474), .B(n22754), .Z(n22756) );
  XOR U22663 ( .A(n22762), .B(n22763), .Z(n15474) );
  AND U22664 ( .A(n591), .B(n22764), .Z(n22763) );
  XOR U22665 ( .A(n22765), .B(n22762), .Z(n22764) );
  XOR U22666 ( .A(n22766), .B(n22767), .Z(n22754) );
  AND U22667 ( .A(n22768), .B(n22769), .Z(n22767) );
  XOR U22668 ( .A(n22766), .B(n15489), .Z(n22769) );
  XOR U22669 ( .A(n22770), .B(n22771), .Z(n15489) );
  AND U22670 ( .A(n594), .B(n22772), .Z(n22771) );
  XOR U22671 ( .A(n22773), .B(n22770), .Z(n22772) );
  XNOR U22672 ( .A(n15486), .B(n22766), .Z(n22768) );
  XOR U22673 ( .A(n22774), .B(n22775), .Z(n15486) );
  AND U22674 ( .A(n591), .B(n22776), .Z(n22775) );
  XOR U22675 ( .A(n22777), .B(n22774), .Z(n22776) );
  XOR U22676 ( .A(n22778), .B(n22779), .Z(n22766) );
  AND U22677 ( .A(n22780), .B(n22781), .Z(n22779) );
  XOR U22678 ( .A(n22778), .B(n15501), .Z(n22781) );
  XOR U22679 ( .A(n22782), .B(n22783), .Z(n15501) );
  AND U22680 ( .A(n594), .B(n22784), .Z(n22783) );
  XOR U22681 ( .A(n22785), .B(n22782), .Z(n22784) );
  XNOR U22682 ( .A(n15498), .B(n22778), .Z(n22780) );
  XOR U22683 ( .A(n22786), .B(n22787), .Z(n15498) );
  AND U22684 ( .A(n591), .B(n22788), .Z(n22787) );
  XOR U22685 ( .A(n22789), .B(n22786), .Z(n22788) );
  XOR U22686 ( .A(n22790), .B(n22791), .Z(n22778) );
  AND U22687 ( .A(n22792), .B(n22793), .Z(n22791) );
  XOR U22688 ( .A(n22790), .B(n15513), .Z(n22793) );
  XOR U22689 ( .A(n22794), .B(n22795), .Z(n15513) );
  AND U22690 ( .A(n594), .B(n22796), .Z(n22795) );
  XOR U22691 ( .A(n22797), .B(n22794), .Z(n22796) );
  XNOR U22692 ( .A(n15510), .B(n22790), .Z(n22792) );
  XOR U22693 ( .A(n22798), .B(n22799), .Z(n15510) );
  AND U22694 ( .A(n591), .B(n22800), .Z(n22799) );
  XOR U22695 ( .A(n22801), .B(n22798), .Z(n22800) );
  XOR U22696 ( .A(n22802), .B(n22803), .Z(n22790) );
  AND U22697 ( .A(n22804), .B(n22805), .Z(n22803) );
  XOR U22698 ( .A(n22802), .B(n15525), .Z(n22805) );
  XOR U22699 ( .A(n22806), .B(n22807), .Z(n15525) );
  AND U22700 ( .A(n594), .B(n22808), .Z(n22807) );
  XOR U22701 ( .A(n22809), .B(n22806), .Z(n22808) );
  XNOR U22702 ( .A(n15522), .B(n22802), .Z(n22804) );
  XOR U22703 ( .A(n22810), .B(n22811), .Z(n15522) );
  AND U22704 ( .A(n591), .B(n22812), .Z(n22811) );
  XOR U22705 ( .A(n22813), .B(n22810), .Z(n22812) );
  XOR U22706 ( .A(n22814), .B(n22815), .Z(n22802) );
  AND U22707 ( .A(n22816), .B(n22817), .Z(n22815) );
  XOR U22708 ( .A(n22814), .B(n15537), .Z(n22817) );
  XOR U22709 ( .A(n22818), .B(n22819), .Z(n15537) );
  AND U22710 ( .A(n594), .B(n22820), .Z(n22819) );
  XOR U22711 ( .A(n22821), .B(n22818), .Z(n22820) );
  XNOR U22712 ( .A(n15534), .B(n22814), .Z(n22816) );
  XOR U22713 ( .A(n22822), .B(n22823), .Z(n15534) );
  AND U22714 ( .A(n591), .B(n22824), .Z(n22823) );
  XOR U22715 ( .A(n22825), .B(n22822), .Z(n22824) );
  XOR U22716 ( .A(n22826), .B(n22827), .Z(n22814) );
  AND U22717 ( .A(n22828), .B(n22829), .Z(n22827) );
  XOR U22718 ( .A(n22826), .B(n15549), .Z(n22829) );
  XOR U22719 ( .A(n22830), .B(n22831), .Z(n15549) );
  AND U22720 ( .A(n594), .B(n22832), .Z(n22831) );
  XOR U22721 ( .A(n22833), .B(n22830), .Z(n22832) );
  XNOR U22722 ( .A(n15546), .B(n22826), .Z(n22828) );
  XOR U22723 ( .A(n22834), .B(n22835), .Z(n15546) );
  AND U22724 ( .A(n591), .B(n22836), .Z(n22835) );
  XOR U22725 ( .A(n22837), .B(n22834), .Z(n22836) );
  XOR U22726 ( .A(n22838), .B(n22839), .Z(n22826) );
  AND U22727 ( .A(n22840), .B(n22841), .Z(n22839) );
  XOR U22728 ( .A(n22838), .B(n15561), .Z(n22841) );
  XOR U22729 ( .A(n22842), .B(n22843), .Z(n15561) );
  AND U22730 ( .A(n594), .B(n22844), .Z(n22843) );
  XOR U22731 ( .A(n22845), .B(n22842), .Z(n22844) );
  XNOR U22732 ( .A(n15558), .B(n22838), .Z(n22840) );
  XOR U22733 ( .A(n22846), .B(n22847), .Z(n15558) );
  AND U22734 ( .A(n591), .B(n22848), .Z(n22847) );
  XOR U22735 ( .A(n22849), .B(n22846), .Z(n22848) );
  XOR U22736 ( .A(n22850), .B(n22851), .Z(n22838) );
  AND U22737 ( .A(n22852), .B(n22853), .Z(n22851) );
  XOR U22738 ( .A(n15573), .B(n22850), .Z(n22853) );
  XOR U22739 ( .A(n22854), .B(n22855), .Z(n15573) );
  AND U22740 ( .A(n594), .B(n22856), .Z(n22855) );
  XOR U22741 ( .A(n22854), .B(n22857), .Z(n22856) );
  XNOR U22742 ( .A(n22850), .B(n15570), .Z(n22852) );
  XOR U22743 ( .A(n22858), .B(n22859), .Z(n15570) );
  AND U22744 ( .A(n591), .B(n22860), .Z(n22859) );
  XOR U22745 ( .A(n22858), .B(n22861), .Z(n22860) );
  XOR U22746 ( .A(n22862), .B(n22863), .Z(n22850) );
  AND U22747 ( .A(n22864), .B(n22865), .Z(n22863) );
  XNOR U22748 ( .A(n22866), .B(n15586), .Z(n22865) );
  XOR U22749 ( .A(n22867), .B(n22868), .Z(n15586) );
  AND U22750 ( .A(n594), .B(n22869), .Z(n22868) );
  XOR U22751 ( .A(n22870), .B(n22867), .Z(n22869) );
  XNOR U22752 ( .A(n15583), .B(n22862), .Z(n22864) );
  XOR U22753 ( .A(n22871), .B(n22872), .Z(n15583) );
  AND U22754 ( .A(n591), .B(n22873), .Z(n22872) );
  XOR U22755 ( .A(n22874), .B(n22871), .Z(n22873) );
  IV U22756 ( .A(n22866), .Z(n22862) );
  AND U22757 ( .A(n22498), .B(n22501), .Z(n22866) );
  XNOR U22758 ( .A(n22875), .B(n22876), .Z(n22501) );
  AND U22759 ( .A(n594), .B(n22877), .Z(n22876) );
  XNOR U22760 ( .A(n22878), .B(n22875), .Z(n22877) );
  XOR U22761 ( .A(n22879), .B(n22880), .Z(n594) );
  AND U22762 ( .A(n22881), .B(n22882), .Z(n22880) );
  XOR U22763 ( .A(n22879), .B(n22509), .Z(n22882) );
  XOR U22764 ( .A(n22883), .B(n22884), .Z(n22509) );
  AND U22765 ( .A(n530), .B(n22885), .Z(n22884) );
  XOR U22766 ( .A(n22886), .B(n22883), .Z(n22885) );
  XNOR U22767 ( .A(n22506), .B(n22879), .Z(n22881) );
  XOR U22768 ( .A(n22887), .B(n22888), .Z(n22506) );
  AND U22769 ( .A(n528), .B(n22889), .Z(n22888) );
  XOR U22770 ( .A(n22890), .B(n22887), .Z(n22889) );
  XOR U22771 ( .A(n22891), .B(n22892), .Z(n22879) );
  AND U22772 ( .A(n22893), .B(n22894), .Z(n22892) );
  XOR U22773 ( .A(n22891), .B(n22521), .Z(n22894) );
  XOR U22774 ( .A(n22895), .B(n22896), .Z(n22521) );
  AND U22775 ( .A(n530), .B(n22897), .Z(n22896) );
  XOR U22776 ( .A(n22898), .B(n22895), .Z(n22897) );
  XNOR U22777 ( .A(n22518), .B(n22891), .Z(n22893) );
  XOR U22778 ( .A(n22899), .B(n22900), .Z(n22518) );
  AND U22779 ( .A(n528), .B(n22901), .Z(n22900) );
  XOR U22780 ( .A(n22902), .B(n22899), .Z(n22901) );
  XOR U22781 ( .A(n22903), .B(n22904), .Z(n22891) );
  AND U22782 ( .A(n22905), .B(n22906), .Z(n22904) );
  XOR U22783 ( .A(n22903), .B(n22533), .Z(n22906) );
  XOR U22784 ( .A(n22907), .B(n22908), .Z(n22533) );
  AND U22785 ( .A(n530), .B(n22909), .Z(n22908) );
  XOR U22786 ( .A(n22910), .B(n22907), .Z(n22909) );
  XNOR U22787 ( .A(n22530), .B(n22903), .Z(n22905) );
  XOR U22788 ( .A(n22911), .B(n22912), .Z(n22530) );
  AND U22789 ( .A(n528), .B(n22913), .Z(n22912) );
  XOR U22790 ( .A(n22914), .B(n22911), .Z(n22913) );
  XOR U22791 ( .A(n22915), .B(n22916), .Z(n22903) );
  AND U22792 ( .A(n22917), .B(n22918), .Z(n22916) );
  XOR U22793 ( .A(n22915), .B(n22545), .Z(n22918) );
  XOR U22794 ( .A(n22919), .B(n22920), .Z(n22545) );
  AND U22795 ( .A(n530), .B(n22921), .Z(n22920) );
  XOR U22796 ( .A(n22922), .B(n22919), .Z(n22921) );
  XNOR U22797 ( .A(n22542), .B(n22915), .Z(n22917) );
  XOR U22798 ( .A(n22923), .B(n22924), .Z(n22542) );
  AND U22799 ( .A(n528), .B(n22925), .Z(n22924) );
  XOR U22800 ( .A(n22926), .B(n22923), .Z(n22925) );
  XOR U22801 ( .A(n22927), .B(n22928), .Z(n22915) );
  AND U22802 ( .A(n22929), .B(n22930), .Z(n22928) );
  XOR U22803 ( .A(n22927), .B(n22557), .Z(n22930) );
  XOR U22804 ( .A(n22931), .B(n22932), .Z(n22557) );
  AND U22805 ( .A(n530), .B(n22933), .Z(n22932) );
  XOR U22806 ( .A(n22934), .B(n22931), .Z(n22933) );
  XNOR U22807 ( .A(n22554), .B(n22927), .Z(n22929) );
  XOR U22808 ( .A(n22935), .B(n22936), .Z(n22554) );
  AND U22809 ( .A(n528), .B(n22937), .Z(n22936) );
  XOR U22810 ( .A(n22938), .B(n22935), .Z(n22937) );
  XOR U22811 ( .A(n22939), .B(n22940), .Z(n22927) );
  AND U22812 ( .A(n22941), .B(n22942), .Z(n22940) );
  XOR U22813 ( .A(n22939), .B(n22569), .Z(n22942) );
  XOR U22814 ( .A(n22943), .B(n22944), .Z(n22569) );
  AND U22815 ( .A(n530), .B(n22945), .Z(n22944) );
  XOR U22816 ( .A(n22946), .B(n22943), .Z(n22945) );
  XNOR U22817 ( .A(n22566), .B(n22939), .Z(n22941) );
  XOR U22818 ( .A(n22947), .B(n22948), .Z(n22566) );
  AND U22819 ( .A(n528), .B(n22949), .Z(n22948) );
  XOR U22820 ( .A(n22950), .B(n22947), .Z(n22949) );
  XOR U22821 ( .A(n22951), .B(n22952), .Z(n22939) );
  AND U22822 ( .A(n22953), .B(n22954), .Z(n22952) );
  XOR U22823 ( .A(n22951), .B(n22581), .Z(n22954) );
  XOR U22824 ( .A(n22955), .B(n22956), .Z(n22581) );
  AND U22825 ( .A(n530), .B(n22957), .Z(n22956) );
  XOR U22826 ( .A(n22958), .B(n22955), .Z(n22957) );
  XNOR U22827 ( .A(n22578), .B(n22951), .Z(n22953) );
  XOR U22828 ( .A(n22959), .B(n22960), .Z(n22578) );
  AND U22829 ( .A(n528), .B(n22961), .Z(n22960) );
  XOR U22830 ( .A(n22962), .B(n22959), .Z(n22961) );
  XOR U22831 ( .A(n22963), .B(n22964), .Z(n22951) );
  AND U22832 ( .A(n22965), .B(n22966), .Z(n22964) );
  XOR U22833 ( .A(n22963), .B(n22593), .Z(n22966) );
  XOR U22834 ( .A(n22967), .B(n22968), .Z(n22593) );
  AND U22835 ( .A(n530), .B(n22969), .Z(n22968) );
  XOR U22836 ( .A(n22970), .B(n22967), .Z(n22969) );
  XNOR U22837 ( .A(n22590), .B(n22963), .Z(n22965) );
  XOR U22838 ( .A(n22971), .B(n22972), .Z(n22590) );
  AND U22839 ( .A(n528), .B(n22973), .Z(n22972) );
  XOR U22840 ( .A(n22974), .B(n22971), .Z(n22973) );
  XOR U22841 ( .A(n22975), .B(n22976), .Z(n22963) );
  AND U22842 ( .A(n22977), .B(n22978), .Z(n22976) );
  XOR U22843 ( .A(n22975), .B(n22605), .Z(n22978) );
  XOR U22844 ( .A(n22979), .B(n22980), .Z(n22605) );
  AND U22845 ( .A(n530), .B(n22981), .Z(n22980) );
  XOR U22846 ( .A(n22982), .B(n22979), .Z(n22981) );
  XNOR U22847 ( .A(n22602), .B(n22975), .Z(n22977) );
  XOR U22848 ( .A(n22983), .B(n22984), .Z(n22602) );
  AND U22849 ( .A(n528), .B(n22985), .Z(n22984) );
  XOR U22850 ( .A(n22986), .B(n22983), .Z(n22985) );
  XOR U22851 ( .A(n22987), .B(n22988), .Z(n22975) );
  AND U22852 ( .A(n22989), .B(n22990), .Z(n22988) );
  XOR U22853 ( .A(n22987), .B(n22617), .Z(n22990) );
  XOR U22854 ( .A(n22991), .B(n22992), .Z(n22617) );
  AND U22855 ( .A(n530), .B(n22993), .Z(n22992) );
  XOR U22856 ( .A(n22994), .B(n22991), .Z(n22993) );
  XNOR U22857 ( .A(n22614), .B(n22987), .Z(n22989) );
  XOR U22858 ( .A(n22995), .B(n22996), .Z(n22614) );
  AND U22859 ( .A(n528), .B(n22997), .Z(n22996) );
  XOR U22860 ( .A(n22998), .B(n22995), .Z(n22997) );
  XOR U22861 ( .A(n22999), .B(n23000), .Z(n22987) );
  AND U22862 ( .A(n23001), .B(n23002), .Z(n23000) );
  XOR U22863 ( .A(n22999), .B(n22629), .Z(n23002) );
  XOR U22864 ( .A(n23003), .B(n23004), .Z(n22629) );
  AND U22865 ( .A(n530), .B(n23005), .Z(n23004) );
  XOR U22866 ( .A(n23006), .B(n23003), .Z(n23005) );
  XNOR U22867 ( .A(n22626), .B(n22999), .Z(n23001) );
  XOR U22868 ( .A(n23007), .B(n23008), .Z(n22626) );
  AND U22869 ( .A(n528), .B(n23009), .Z(n23008) );
  XOR U22870 ( .A(n23010), .B(n23007), .Z(n23009) );
  XOR U22871 ( .A(n23011), .B(n23012), .Z(n22999) );
  AND U22872 ( .A(n23013), .B(n23014), .Z(n23012) );
  XOR U22873 ( .A(n23011), .B(n22641), .Z(n23014) );
  XOR U22874 ( .A(n23015), .B(n23016), .Z(n22641) );
  AND U22875 ( .A(n530), .B(n23017), .Z(n23016) );
  XOR U22876 ( .A(n23018), .B(n23015), .Z(n23017) );
  XNOR U22877 ( .A(n22638), .B(n23011), .Z(n23013) );
  XOR U22878 ( .A(n23019), .B(n23020), .Z(n22638) );
  AND U22879 ( .A(n528), .B(n23021), .Z(n23020) );
  XOR U22880 ( .A(n23022), .B(n23019), .Z(n23021) );
  XOR U22881 ( .A(n23023), .B(n23024), .Z(n23011) );
  AND U22882 ( .A(n23025), .B(n23026), .Z(n23024) );
  XOR U22883 ( .A(n23023), .B(n22653), .Z(n23026) );
  XOR U22884 ( .A(n23027), .B(n23028), .Z(n22653) );
  AND U22885 ( .A(n530), .B(n23029), .Z(n23028) );
  XOR U22886 ( .A(n23030), .B(n23027), .Z(n23029) );
  XNOR U22887 ( .A(n22650), .B(n23023), .Z(n23025) );
  XOR U22888 ( .A(n23031), .B(n23032), .Z(n22650) );
  AND U22889 ( .A(n528), .B(n23033), .Z(n23032) );
  XOR U22890 ( .A(n23034), .B(n23031), .Z(n23033) );
  XOR U22891 ( .A(n23035), .B(n23036), .Z(n23023) );
  AND U22892 ( .A(n23037), .B(n23038), .Z(n23036) );
  XOR U22893 ( .A(n23035), .B(n22665), .Z(n23038) );
  XOR U22894 ( .A(n23039), .B(n23040), .Z(n22665) );
  AND U22895 ( .A(n530), .B(n23041), .Z(n23040) );
  XOR U22896 ( .A(n23042), .B(n23039), .Z(n23041) );
  XNOR U22897 ( .A(n22662), .B(n23035), .Z(n23037) );
  XOR U22898 ( .A(n23043), .B(n23044), .Z(n22662) );
  AND U22899 ( .A(n528), .B(n23045), .Z(n23044) );
  XOR U22900 ( .A(n23046), .B(n23043), .Z(n23045) );
  XOR U22901 ( .A(n23047), .B(n23048), .Z(n23035) );
  AND U22902 ( .A(n23049), .B(n23050), .Z(n23048) );
  XOR U22903 ( .A(n23047), .B(n22677), .Z(n23050) );
  XOR U22904 ( .A(n23051), .B(n23052), .Z(n22677) );
  AND U22905 ( .A(n530), .B(n23053), .Z(n23052) );
  XOR U22906 ( .A(n23054), .B(n23051), .Z(n23053) );
  XNOR U22907 ( .A(n22674), .B(n23047), .Z(n23049) );
  XOR U22908 ( .A(n23055), .B(n23056), .Z(n22674) );
  AND U22909 ( .A(n528), .B(n23057), .Z(n23056) );
  XOR U22910 ( .A(n23058), .B(n23055), .Z(n23057) );
  XOR U22911 ( .A(n23059), .B(n23060), .Z(n23047) );
  AND U22912 ( .A(n23061), .B(n23062), .Z(n23060) );
  XOR U22913 ( .A(n23059), .B(n22689), .Z(n23062) );
  XOR U22914 ( .A(n23063), .B(n23064), .Z(n22689) );
  AND U22915 ( .A(n530), .B(n23065), .Z(n23064) );
  XOR U22916 ( .A(n23066), .B(n23063), .Z(n23065) );
  XNOR U22917 ( .A(n22686), .B(n23059), .Z(n23061) );
  XOR U22918 ( .A(n23067), .B(n23068), .Z(n22686) );
  AND U22919 ( .A(n528), .B(n23069), .Z(n23068) );
  XOR U22920 ( .A(n23070), .B(n23067), .Z(n23069) );
  XOR U22921 ( .A(n23071), .B(n23072), .Z(n23059) );
  AND U22922 ( .A(n23073), .B(n23074), .Z(n23072) );
  XOR U22923 ( .A(n23071), .B(n22701), .Z(n23074) );
  XOR U22924 ( .A(n23075), .B(n23076), .Z(n22701) );
  AND U22925 ( .A(n530), .B(n23077), .Z(n23076) );
  XOR U22926 ( .A(n23078), .B(n23075), .Z(n23077) );
  XNOR U22927 ( .A(n22698), .B(n23071), .Z(n23073) );
  XOR U22928 ( .A(n23079), .B(n23080), .Z(n22698) );
  AND U22929 ( .A(n528), .B(n23081), .Z(n23080) );
  XOR U22930 ( .A(n23082), .B(n23079), .Z(n23081) );
  XOR U22931 ( .A(n23083), .B(n23084), .Z(n23071) );
  AND U22932 ( .A(n23085), .B(n23086), .Z(n23084) );
  XOR U22933 ( .A(n23083), .B(n22713), .Z(n23086) );
  XOR U22934 ( .A(n23087), .B(n23088), .Z(n22713) );
  AND U22935 ( .A(n530), .B(n23089), .Z(n23088) );
  XOR U22936 ( .A(n23090), .B(n23087), .Z(n23089) );
  XNOR U22937 ( .A(n22710), .B(n23083), .Z(n23085) );
  XOR U22938 ( .A(n23091), .B(n23092), .Z(n22710) );
  AND U22939 ( .A(n528), .B(n23093), .Z(n23092) );
  XOR U22940 ( .A(n23094), .B(n23091), .Z(n23093) );
  XOR U22941 ( .A(n23095), .B(n23096), .Z(n23083) );
  AND U22942 ( .A(n23097), .B(n23098), .Z(n23096) );
  XOR U22943 ( .A(n23095), .B(n22725), .Z(n23098) );
  XOR U22944 ( .A(n23099), .B(n23100), .Z(n22725) );
  AND U22945 ( .A(n530), .B(n23101), .Z(n23100) );
  XOR U22946 ( .A(n23102), .B(n23099), .Z(n23101) );
  XNOR U22947 ( .A(n22722), .B(n23095), .Z(n23097) );
  XOR U22948 ( .A(n23103), .B(n23104), .Z(n22722) );
  AND U22949 ( .A(n528), .B(n23105), .Z(n23104) );
  XOR U22950 ( .A(n23106), .B(n23103), .Z(n23105) );
  XOR U22951 ( .A(n23107), .B(n23108), .Z(n23095) );
  AND U22952 ( .A(n23109), .B(n23110), .Z(n23108) );
  XOR U22953 ( .A(n23107), .B(n22737), .Z(n23110) );
  XOR U22954 ( .A(n23111), .B(n23112), .Z(n22737) );
  AND U22955 ( .A(n530), .B(n23113), .Z(n23112) );
  XOR U22956 ( .A(n23114), .B(n23111), .Z(n23113) );
  XNOR U22957 ( .A(n22734), .B(n23107), .Z(n23109) );
  XOR U22958 ( .A(n23115), .B(n23116), .Z(n22734) );
  AND U22959 ( .A(n528), .B(n23117), .Z(n23116) );
  XOR U22960 ( .A(n23118), .B(n23115), .Z(n23117) );
  XOR U22961 ( .A(n23119), .B(n23120), .Z(n23107) );
  AND U22962 ( .A(n23121), .B(n23122), .Z(n23120) );
  XOR U22963 ( .A(n23119), .B(n22749), .Z(n23122) );
  XOR U22964 ( .A(n23123), .B(n23124), .Z(n22749) );
  AND U22965 ( .A(n530), .B(n23125), .Z(n23124) );
  XOR U22966 ( .A(n23126), .B(n23123), .Z(n23125) );
  XNOR U22967 ( .A(n22746), .B(n23119), .Z(n23121) );
  XOR U22968 ( .A(n23127), .B(n23128), .Z(n22746) );
  AND U22969 ( .A(n528), .B(n23129), .Z(n23128) );
  XOR U22970 ( .A(n23130), .B(n23127), .Z(n23129) );
  XOR U22971 ( .A(n23131), .B(n23132), .Z(n23119) );
  AND U22972 ( .A(n23133), .B(n23134), .Z(n23132) );
  XOR U22973 ( .A(n23131), .B(n22761), .Z(n23134) );
  XOR U22974 ( .A(n23135), .B(n23136), .Z(n22761) );
  AND U22975 ( .A(n530), .B(n23137), .Z(n23136) );
  XOR U22976 ( .A(n23138), .B(n23135), .Z(n23137) );
  XNOR U22977 ( .A(n22758), .B(n23131), .Z(n23133) );
  XOR U22978 ( .A(n23139), .B(n23140), .Z(n22758) );
  AND U22979 ( .A(n528), .B(n23141), .Z(n23140) );
  XOR U22980 ( .A(n23142), .B(n23139), .Z(n23141) );
  XOR U22981 ( .A(n23143), .B(n23144), .Z(n23131) );
  AND U22982 ( .A(n23145), .B(n23146), .Z(n23144) );
  XOR U22983 ( .A(n23143), .B(n22773), .Z(n23146) );
  XOR U22984 ( .A(n23147), .B(n23148), .Z(n22773) );
  AND U22985 ( .A(n530), .B(n23149), .Z(n23148) );
  XOR U22986 ( .A(n23150), .B(n23147), .Z(n23149) );
  XNOR U22987 ( .A(n22770), .B(n23143), .Z(n23145) );
  XOR U22988 ( .A(n23151), .B(n23152), .Z(n22770) );
  AND U22989 ( .A(n528), .B(n23153), .Z(n23152) );
  XOR U22990 ( .A(n23154), .B(n23151), .Z(n23153) );
  XOR U22991 ( .A(n23155), .B(n23156), .Z(n23143) );
  AND U22992 ( .A(n23157), .B(n23158), .Z(n23156) );
  XOR U22993 ( .A(n23155), .B(n22785), .Z(n23158) );
  XOR U22994 ( .A(n23159), .B(n23160), .Z(n22785) );
  AND U22995 ( .A(n530), .B(n23161), .Z(n23160) );
  XOR U22996 ( .A(n23162), .B(n23159), .Z(n23161) );
  XNOR U22997 ( .A(n22782), .B(n23155), .Z(n23157) );
  XOR U22998 ( .A(n23163), .B(n23164), .Z(n22782) );
  AND U22999 ( .A(n528), .B(n23165), .Z(n23164) );
  XOR U23000 ( .A(n23166), .B(n23163), .Z(n23165) );
  XOR U23001 ( .A(n23167), .B(n23168), .Z(n23155) );
  AND U23002 ( .A(n23169), .B(n23170), .Z(n23168) );
  XOR U23003 ( .A(n23167), .B(n22797), .Z(n23170) );
  XOR U23004 ( .A(n23171), .B(n23172), .Z(n22797) );
  AND U23005 ( .A(n530), .B(n23173), .Z(n23172) );
  XOR U23006 ( .A(n23174), .B(n23171), .Z(n23173) );
  XNOR U23007 ( .A(n22794), .B(n23167), .Z(n23169) );
  XOR U23008 ( .A(n23175), .B(n23176), .Z(n22794) );
  AND U23009 ( .A(n528), .B(n23177), .Z(n23176) );
  XOR U23010 ( .A(n23178), .B(n23175), .Z(n23177) );
  XOR U23011 ( .A(n23179), .B(n23180), .Z(n23167) );
  AND U23012 ( .A(n23181), .B(n23182), .Z(n23180) );
  XOR U23013 ( .A(n23179), .B(n22809), .Z(n23182) );
  XOR U23014 ( .A(n23183), .B(n23184), .Z(n22809) );
  AND U23015 ( .A(n530), .B(n23185), .Z(n23184) );
  XOR U23016 ( .A(n23186), .B(n23183), .Z(n23185) );
  XNOR U23017 ( .A(n22806), .B(n23179), .Z(n23181) );
  XOR U23018 ( .A(n23187), .B(n23188), .Z(n22806) );
  AND U23019 ( .A(n528), .B(n23189), .Z(n23188) );
  XOR U23020 ( .A(n23190), .B(n23187), .Z(n23189) );
  XOR U23021 ( .A(n23191), .B(n23192), .Z(n23179) );
  AND U23022 ( .A(n23193), .B(n23194), .Z(n23192) );
  XOR U23023 ( .A(n23191), .B(n22821), .Z(n23194) );
  XOR U23024 ( .A(n23195), .B(n23196), .Z(n22821) );
  AND U23025 ( .A(n530), .B(n23197), .Z(n23196) );
  XOR U23026 ( .A(n23198), .B(n23195), .Z(n23197) );
  XNOR U23027 ( .A(n22818), .B(n23191), .Z(n23193) );
  XOR U23028 ( .A(n23199), .B(n23200), .Z(n22818) );
  AND U23029 ( .A(n528), .B(n23201), .Z(n23200) );
  XOR U23030 ( .A(n23202), .B(n23199), .Z(n23201) );
  XOR U23031 ( .A(n23203), .B(n23204), .Z(n23191) );
  AND U23032 ( .A(n23205), .B(n23206), .Z(n23204) );
  XOR U23033 ( .A(n23203), .B(n22833), .Z(n23206) );
  XOR U23034 ( .A(n23207), .B(n23208), .Z(n22833) );
  AND U23035 ( .A(n530), .B(n23209), .Z(n23208) );
  XOR U23036 ( .A(n23210), .B(n23207), .Z(n23209) );
  XNOR U23037 ( .A(n22830), .B(n23203), .Z(n23205) );
  XOR U23038 ( .A(n23211), .B(n23212), .Z(n22830) );
  AND U23039 ( .A(n528), .B(n23213), .Z(n23212) );
  XOR U23040 ( .A(n23214), .B(n23211), .Z(n23213) );
  XOR U23041 ( .A(n23215), .B(n23216), .Z(n23203) );
  AND U23042 ( .A(n23217), .B(n23218), .Z(n23216) );
  XOR U23043 ( .A(n23215), .B(n22845), .Z(n23218) );
  XOR U23044 ( .A(n23219), .B(n23220), .Z(n22845) );
  AND U23045 ( .A(n530), .B(n23221), .Z(n23220) );
  XOR U23046 ( .A(n23222), .B(n23219), .Z(n23221) );
  XNOR U23047 ( .A(n22842), .B(n23215), .Z(n23217) );
  XOR U23048 ( .A(n23223), .B(n23224), .Z(n22842) );
  AND U23049 ( .A(n528), .B(n23225), .Z(n23224) );
  XOR U23050 ( .A(n23226), .B(n23223), .Z(n23225) );
  XOR U23051 ( .A(n23227), .B(n23228), .Z(n23215) );
  AND U23052 ( .A(n23229), .B(n23230), .Z(n23228) );
  XOR U23053 ( .A(n22857), .B(n23227), .Z(n23230) );
  XOR U23054 ( .A(n23231), .B(n23232), .Z(n22857) );
  AND U23055 ( .A(n530), .B(n23233), .Z(n23232) );
  XOR U23056 ( .A(n23231), .B(n23234), .Z(n23233) );
  XNOR U23057 ( .A(n23227), .B(n22854), .Z(n23229) );
  XOR U23058 ( .A(n23235), .B(n23236), .Z(n22854) );
  AND U23059 ( .A(n528), .B(n23237), .Z(n23236) );
  XOR U23060 ( .A(n23235), .B(n23238), .Z(n23237) );
  XOR U23061 ( .A(n23239), .B(n23240), .Z(n23227) );
  AND U23062 ( .A(n23241), .B(n23242), .Z(n23240) );
  XNOR U23063 ( .A(n23243), .B(n22870), .Z(n23242) );
  XOR U23064 ( .A(n23244), .B(n23245), .Z(n22870) );
  AND U23065 ( .A(n530), .B(n23246), .Z(n23245) );
  XOR U23066 ( .A(n23247), .B(n23244), .Z(n23246) );
  XNOR U23067 ( .A(n22867), .B(n23239), .Z(n23241) );
  XOR U23068 ( .A(n23248), .B(n23249), .Z(n22867) );
  AND U23069 ( .A(n528), .B(n23250), .Z(n23249) );
  XOR U23070 ( .A(n23251), .B(n23248), .Z(n23250) );
  IV U23071 ( .A(n23243), .Z(n23239) );
  AND U23072 ( .A(n22875), .B(n22878), .Z(n23243) );
  XNOR U23073 ( .A(n23252), .B(n23253), .Z(n22878) );
  AND U23074 ( .A(n530), .B(n23254), .Z(n23253) );
  XNOR U23075 ( .A(n23255), .B(n23252), .Z(n23254) );
  XOR U23076 ( .A(n23256), .B(n23257), .Z(n530) );
  AND U23077 ( .A(n23258), .B(n23259), .Z(n23257) );
  XOR U23078 ( .A(n23256), .B(n22886), .Z(n23259) );
  XNOR U23079 ( .A(n23260), .B(n23261), .Z(n22886) );
  AND U23080 ( .A(n23262), .B(n394), .Z(n23261) );
  AND U23081 ( .A(n23260), .B(n23263), .Z(n23262) );
  XNOR U23082 ( .A(n22883), .B(n23256), .Z(n23258) );
  XOR U23083 ( .A(n23264), .B(n23265), .Z(n22883) );
  AND U23084 ( .A(n23266), .B(n392), .Z(n23265) );
  NOR U23085 ( .A(n23264), .B(n23267), .Z(n23266) );
  XOR U23086 ( .A(n23268), .B(n23269), .Z(n23256) );
  AND U23087 ( .A(n23270), .B(n23271), .Z(n23269) );
  XOR U23088 ( .A(n23268), .B(n22898), .Z(n23271) );
  XOR U23089 ( .A(n23272), .B(n23273), .Z(n22898) );
  AND U23090 ( .A(n394), .B(n23274), .Z(n23273) );
  XOR U23091 ( .A(n23275), .B(n23272), .Z(n23274) );
  XNOR U23092 ( .A(n22895), .B(n23268), .Z(n23270) );
  XOR U23093 ( .A(n23276), .B(n23277), .Z(n22895) );
  AND U23094 ( .A(n392), .B(n23278), .Z(n23277) );
  XOR U23095 ( .A(n23279), .B(n23276), .Z(n23278) );
  XOR U23096 ( .A(n23280), .B(n23281), .Z(n23268) );
  AND U23097 ( .A(n23282), .B(n23283), .Z(n23281) );
  XOR U23098 ( .A(n23280), .B(n22910), .Z(n23283) );
  XOR U23099 ( .A(n23284), .B(n23285), .Z(n22910) );
  AND U23100 ( .A(n394), .B(n23286), .Z(n23285) );
  XOR U23101 ( .A(n23287), .B(n23284), .Z(n23286) );
  XNOR U23102 ( .A(n22907), .B(n23280), .Z(n23282) );
  XOR U23103 ( .A(n23288), .B(n23289), .Z(n22907) );
  AND U23104 ( .A(n392), .B(n23290), .Z(n23289) );
  XOR U23105 ( .A(n23291), .B(n23288), .Z(n23290) );
  XOR U23106 ( .A(n23292), .B(n23293), .Z(n23280) );
  AND U23107 ( .A(n23294), .B(n23295), .Z(n23293) );
  XOR U23108 ( .A(n23292), .B(n22922), .Z(n23295) );
  XOR U23109 ( .A(n23296), .B(n23297), .Z(n22922) );
  AND U23110 ( .A(n394), .B(n23298), .Z(n23297) );
  XOR U23111 ( .A(n23299), .B(n23296), .Z(n23298) );
  XNOR U23112 ( .A(n22919), .B(n23292), .Z(n23294) );
  XOR U23113 ( .A(n23300), .B(n23301), .Z(n22919) );
  AND U23114 ( .A(n392), .B(n23302), .Z(n23301) );
  XOR U23115 ( .A(n23303), .B(n23300), .Z(n23302) );
  XOR U23116 ( .A(n23304), .B(n23305), .Z(n23292) );
  AND U23117 ( .A(n23306), .B(n23307), .Z(n23305) );
  XOR U23118 ( .A(n23304), .B(n22934), .Z(n23307) );
  XOR U23119 ( .A(n23308), .B(n23309), .Z(n22934) );
  AND U23120 ( .A(n394), .B(n23310), .Z(n23309) );
  XOR U23121 ( .A(n23311), .B(n23308), .Z(n23310) );
  XNOR U23122 ( .A(n22931), .B(n23304), .Z(n23306) );
  XOR U23123 ( .A(n23312), .B(n23313), .Z(n22931) );
  AND U23124 ( .A(n392), .B(n23314), .Z(n23313) );
  XOR U23125 ( .A(n23315), .B(n23312), .Z(n23314) );
  XOR U23126 ( .A(n23316), .B(n23317), .Z(n23304) );
  AND U23127 ( .A(n23318), .B(n23319), .Z(n23317) );
  XOR U23128 ( .A(n23316), .B(n22946), .Z(n23319) );
  XOR U23129 ( .A(n23320), .B(n23321), .Z(n22946) );
  AND U23130 ( .A(n394), .B(n23322), .Z(n23321) );
  XOR U23131 ( .A(n23323), .B(n23320), .Z(n23322) );
  XNOR U23132 ( .A(n22943), .B(n23316), .Z(n23318) );
  XOR U23133 ( .A(n23324), .B(n23325), .Z(n22943) );
  AND U23134 ( .A(n392), .B(n23326), .Z(n23325) );
  XOR U23135 ( .A(n23327), .B(n23324), .Z(n23326) );
  XOR U23136 ( .A(n23328), .B(n23329), .Z(n23316) );
  AND U23137 ( .A(n23330), .B(n23331), .Z(n23329) );
  XOR U23138 ( .A(n23328), .B(n22958), .Z(n23331) );
  XOR U23139 ( .A(n23332), .B(n23333), .Z(n22958) );
  AND U23140 ( .A(n394), .B(n23334), .Z(n23333) );
  XOR U23141 ( .A(n23335), .B(n23332), .Z(n23334) );
  XNOR U23142 ( .A(n22955), .B(n23328), .Z(n23330) );
  XOR U23143 ( .A(n23336), .B(n23337), .Z(n22955) );
  AND U23144 ( .A(n392), .B(n23338), .Z(n23337) );
  XOR U23145 ( .A(n23339), .B(n23336), .Z(n23338) );
  XOR U23146 ( .A(n23340), .B(n23341), .Z(n23328) );
  AND U23147 ( .A(n23342), .B(n23343), .Z(n23341) );
  XOR U23148 ( .A(n23340), .B(n22970), .Z(n23343) );
  XOR U23149 ( .A(n23344), .B(n23345), .Z(n22970) );
  AND U23150 ( .A(n394), .B(n23346), .Z(n23345) );
  XOR U23151 ( .A(n23347), .B(n23344), .Z(n23346) );
  XNOR U23152 ( .A(n22967), .B(n23340), .Z(n23342) );
  XOR U23153 ( .A(n23348), .B(n23349), .Z(n22967) );
  AND U23154 ( .A(n392), .B(n23350), .Z(n23349) );
  XOR U23155 ( .A(n23351), .B(n23348), .Z(n23350) );
  XOR U23156 ( .A(n23352), .B(n23353), .Z(n23340) );
  AND U23157 ( .A(n23354), .B(n23355), .Z(n23353) );
  XOR U23158 ( .A(n23352), .B(n22982), .Z(n23355) );
  XOR U23159 ( .A(n23356), .B(n23357), .Z(n22982) );
  AND U23160 ( .A(n394), .B(n23358), .Z(n23357) );
  XOR U23161 ( .A(n23359), .B(n23356), .Z(n23358) );
  XNOR U23162 ( .A(n22979), .B(n23352), .Z(n23354) );
  XOR U23163 ( .A(n23360), .B(n23361), .Z(n22979) );
  AND U23164 ( .A(n392), .B(n23362), .Z(n23361) );
  XOR U23165 ( .A(n23363), .B(n23360), .Z(n23362) );
  XOR U23166 ( .A(n23364), .B(n23365), .Z(n23352) );
  AND U23167 ( .A(n23366), .B(n23367), .Z(n23365) );
  XOR U23168 ( .A(n23364), .B(n22994), .Z(n23367) );
  XOR U23169 ( .A(n23368), .B(n23369), .Z(n22994) );
  AND U23170 ( .A(n394), .B(n23370), .Z(n23369) );
  XOR U23171 ( .A(n23371), .B(n23368), .Z(n23370) );
  XNOR U23172 ( .A(n22991), .B(n23364), .Z(n23366) );
  XOR U23173 ( .A(n23372), .B(n23373), .Z(n22991) );
  AND U23174 ( .A(n392), .B(n23374), .Z(n23373) );
  XOR U23175 ( .A(n23375), .B(n23372), .Z(n23374) );
  XOR U23176 ( .A(n23376), .B(n23377), .Z(n23364) );
  AND U23177 ( .A(n23378), .B(n23379), .Z(n23377) );
  XOR U23178 ( .A(n23376), .B(n23006), .Z(n23379) );
  XOR U23179 ( .A(n23380), .B(n23381), .Z(n23006) );
  AND U23180 ( .A(n394), .B(n23382), .Z(n23381) );
  XOR U23181 ( .A(n23383), .B(n23380), .Z(n23382) );
  XNOR U23182 ( .A(n23003), .B(n23376), .Z(n23378) );
  XOR U23183 ( .A(n23384), .B(n23385), .Z(n23003) );
  AND U23184 ( .A(n392), .B(n23386), .Z(n23385) );
  XOR U23185 ( .A(n23387), .B(n23384), .Z(n23386) );
  XOR U23186 ( .A(n23388), .B(n23389), .Z(n23376) );
  AND U23187 ( .A(n23390), .B(n23391), .Z(n23389) );
  XOR U23188 ( .A(n23388), .B(n23018), .Z(n23391) );
  XOR U23189 ( .A(n23392), .B(n23393), .Z(n23018) );
  AND U23190 ( .A(n394), .B(n23394), .Z(n23393) );
  XOR U23191 ( .A(n23395), .B(n23392), .Z(n23394) );
  XNOR U23192 ( .A(n23015), .B(n23388), .Z(n23390) );
  XOR U23193 ( .A(n23396), .B(n23397), .Z(n23015) );
  AND U23194 ( .A(n392), .B(n23398), .Z(n23397) );
  XOR U23195 ( .A(n23399), .B(n23396), .Z(n23398) );
  XOR U23196 ( .A(n23400), .B(n23401), .Z(n23388) );
  AND U23197 ( .A(n23402), .B(n23403), .Z(n23401) );
  XOR U23198 ( .A(n23400), .B(n23030), .Z(n23403) );
  XOR U23199 ( .A(n23404), .B(n23405), .Z(n23030) );
  AND U23200 ( .A(n394), .B(n23406), .Z(n23405) );
  XOR U23201 ( .A(n23407), .B(n23404), .Z(n23406) );
  XNOR U23202 ( .A(n23027), .B(n23400), .Z(n23402) );
  XOR U23203 ( .A(n23408), .B(n23409), .Z(n23027) );
  AND U23204 ( .A(n392), .B(n23410), .Z(n23409) );
  XOR U23205 ( .A(n23411), .B(n23408), .Z(n23410) );
  XOR U23206 ( .A(n23412), .B(n23413), .Z(n23400) );
  AND U23207 ( .A(n23414), .B(n23415), .Z(n23413) );
  XOR U23208 ( .A(n23412), .B(n23042), .Z(n23415) );
  XOR U23209 ( .A(n23416), .B(n23417), .Z(n23042) );
  AND U23210 ( .A(n394), .B(n23418), .Z(n23417) );
  XOR U23211 ( .A(n23419), .B(n23416), .Z(n23418) );
  XNOR U23212 ( .A(n23039), .B(n23412), .Z(n23414) );
  XOR U23213 ( .A(n23420), .B(n23421), .Z(n23039) );
  AND U23214 ( .A(n392), .B(n23422), .Z(n23421) );
  XOR U23215 ( .A(n23423), .B(n23420), .Z(n23422) );
  XOR U23216 ( .A(n23424), .B(n23425), .Z(n23412) );
  AND U23217 ( .A(n23426), .B(n23427), .Z(n23425) );
  XOR U23218 ( .A(n23424), .B(n23054), .Z(n23427) );
  XOR U23219 ( .A(n23428), .B(n23429), .Z(n23054) );
  AND U23220 ( .A(n394), .B(n23430), .Z(n23429) );
  XOR U23221 ( .A(n23431), .B(n23428), .Z(n23430) );
  XNOR U23222 ( .A(n23051), .B(n23424), .Z(n23426) );
  XOR U23223 ( .A(n23432), .B(n23433), .Z(n23051) );
  AND U23224 ( .A(n392), .B(n23434), .Z(n23433) );
  XOR U23225 ( .A(n23435), .B(n23432), .Z(n23434) );
  XOR U23226 ( .A(n23436), .B(n23437), .Z(n23424) );
  AND U23227 ( .A(n23438), .B(n23439), .Z(n23437) );
  XOR U23228 ( .A(n23436), .B(n23066), .Z(n23439) );
  XOR U23229 ( .A(n23440), .B(n23441), .Z(n23066) );
  AND U23230 ( .A(n394), .B(n23442), .Z(n23441) );
  XOR U23231 ( .A(n23443), .B(n23440), .Z(n23442) );
  XNOR U23232 ( .A(n23063), .B(n23436), .Z(n23438) );
  XOR U23233 ( .A(n23444), .B(n23445), .Z(n23063) );
  AND U23234 ( .A(n392), .B(n23446), .Z(n23445) );
  XOR U23235 ( .A(n23447), .B(n23444), .Z(n23446) );
  XOR U23236 ( .A(n23448), .B(n23449), .Z(n23436) );
  AND U23237 ( .A(n23450), .B(n23451), .Z(n23449) );
  XOR U23238 ( .A(n23448), .B(n23078), .Z(n23451) );
  XOR U23239 ( .A(n23452), .B(n23453), .Z(n23078) );
  AND U23240 ( .A(n394), .B(n23454), .Z(n23453) );
  XOR U23241 ( .A(n23455), .B(n23452), .Z(n23454) );
  XNOR U23242 ( .A(n23075), .B(n23448), .Z(n23450) );
  XOR U23243 ( .A(n23456), .B(n23457), .Z(n23075) );
  AND U23244 ( .A(n392), .B(n23458), .Z(n23457) );
  XOR U23245 ( .A(n23459), .B(n23456), .Z(n23458) );
  XOR U23246 ( .A(n23460), .B(n23461), .Z(n23448) );
  AND U23247 ( .A(n23462), .B(n23463), .Z(n23461) );
  XOR U23248 ( .A(n23460), .B(n23090), .Z(n23463) );
  XOR U23249 ( .A(n23464), .B(n23465), .Z(n23090) );
  AND U23250 ( .A(n394), .B(n23466), .Z(n23465) );
  XOR U23251 ( .A(n23467), .B(n23464), .Z(n23466) );
  XNOR U23252 ( .A(n23087), .B(n23460), .Z(n23462) );
  XOR U23253 ( .A(n23468), .B(n23469), .Z(n23087) );
  AND U23254 ( .A(n392), .B(n23470), .Z(n23469) );
  XOR U23255 ( .A(n23471), .B(n23468), .Z(n23470) );
  XOR U23256 ( .A(n23472), .B(n23473), .Z(n23460) );
  AND U23257 ( .A(n23474), .B(n23475), .Z(n23473) );
  XOR U23258 ( .A(n23472), .B(n23102), .Z(n23475) );
  XOR U23259 ( .A(n23476), .B(n23477), .Z(n23102) );
  AND U23260 ( .A(n394), .B(n23478), .Z(n23477) );
  XOR U23261 ( .A(n23479), .B(n23476), .Z(n23478) );
  XNOR U23262 ( .A(n23099), .B(n23472), .Z(n23474) );
  XOR U23263 ( .A(n23480), .B(n23481), .Z(n23099) );
  AND U23264 ( .A(n392), .B(n23482), .Z(n23481) );
  XOR U23265 ( .A(n23483), .B(n23480), .Z(n23482) );
  XOR U23266 ( .A(n23484), .B(n23485), .Z(n23472) );
  AND U23267 ( .A(n23486), .B(n23487), .Z(n23485) );
  XOR U23268 ( .A(n23484), .B(n23114), .Z(n23487) );
  XOR U23269 ( .A(n23488), .B(n23489), .Z(n23114) );
  AND U23270 ( .A(n394), .B(n23490), .Z(n23489) );
  XOR U23271 ( .A(n23491), .B(n23488), .Z(n23490) );
  XNOR U23272 ( .A(n23111), .B(n23484), .Z(n23486) );
  XOR U23273 ( .A(n23492), .B(n23493), .Z(n23111) );
  AND U23274 ( .A(n392), .B(n23494), .Z(n23493) );
  XOR U23275 ( .A(n23495), .B(n23492), .Z(n23494) );
  XOR U23276 ( .A(n23496), .B(n23497), .Z(n23484) );
  AND U23277 ( .A(n23498), .B(n23499), .Z(n23497) );
  XOR U23278 ( .A(n23496), .B(n23126), .Z(n23499) );
  XOR U23279 ( .A(n23500), .B(n23501), .Z(n23126) );
  AND U23280 ( .A(n394), .B(n23502), .Z(n23501) );
  XOR U23281 ( .A(n23503), .B(n23500), .Z(n23502) );
  XNOR U23282 ( .A(n23123), .B(n23496), .Z(n23498) );
  XOR U23283 ( .A(n23504), .B(n23505), .Z(n23123) );
  AND U23284 ( .A(n392), .B(n23506), .Z(n23505) );
  XOR U23285 ( .A(n23507), .B(n23504), .Z(n23506) );
  XOR U23286 ( .A(n23508), .B(n23509), .Z(n23496) );
  AND U23287 ( .A(n23510), .B(n23511), .Z(n23509) );
  XOR U23288 ( .A(n23508), .B(n23138), .Z(n23511) );
  XOR U23289 ( .A(n23512), .B(n23513), .Z(n23138) );
  AND U23290 ( .A(n394), .B(n23514), .Z(n23513) );
  XOR U23291 ( .A(n23515), .B(n23512), .Z(n23514) );
  XNOR U23292 ( .A(n23135), .B(n23508), .Z(n23510) );
  XOR U23293 ( .A(n23516), .B(n23517), .Z(n23135) );
  AND U23294 ( .A(n392), .B(n23518), .Z(n23517) );
  XOR U23295 ( .A(n23519), .B(n23516), .Z(n23518) );
  XOR U23296 ( .A(n23520), .B(n23521), .Z(n23508) );
  AND U23297 ( .A(n23522), .B(n23523), .Z(n23521) );
  XOR U23298 ( .A(n23520), .B(n23150), .Z(n23523) );
  XOR U23299 ( .A(n23524), .B(n23525), .Z(n23150) );
  AND U23300 ( .A(n394), .B(n23526), .Z(n23525) );
  XOR U23301 ( .A(n23527), .B(n23524), .Z(n23526) );
  XNOR U23302 ( .A(n23147), .B(n23520), .Z(n23522) );
  XOR U23303 ( .A(n23528), .B(n23529), .Z(n23147) );
  AND U23304 ( .A(n392), .B(n23530), .Z(n23529) );
  XOR U23305 ( .A(n23531), .B(n23528), .Z(n23530) );
  XOR U23306 ( .A(n23532), .B(n23533), .Z(n23520) );
  AND U23307 ( .A(n23534), .B(n23535), .Z(n23533) );
  XOR U23308 ( .A(n23532), .B(n23162), .Z(n23535) );
  XOR U23309 ( .A(n23536), .B(n23537), .Z(n23162) );
  AND U23310 ( .A(n394), .B(n23538), .Z(n23537) );
  XOR U23311 ( .A(n23539), .B(n23536), .Z(n23538) );
  XNOR U23312 ( .A(n23159), .B(n23532), .Z(n23534) );
  XOR U23313 ( .A(n23540), .B(n23541), .Z(n23159) );
  AND U23314 ( .A(n392), .B(n23542), .Z(n23541) );
  XOR U23315 ( .A(n23543), .B(n23540), .Z(n23542) );
  XOR U23316 ( .A(n23544), .B(n23545), .Z(n23532) );
  AND U23317 ( .A(n23546), .B(n23547), .Z(n23545) );
  XOR U23318 ( .A(n23544), .B(n23174), .Z(n23547) );
  XOR U23319 ( .A(n23548), .B(n23549), .Z(n23174) );
  AND U23320 ( .A(n394), .B(n23550), .Z(n23549) );
  XOR U23321 ( .A(n23551), .B(n23548), .Z(n23550) );
  XNOR U23322 ( .A(n23171), .B(n23544), .Z(n23546) );
  XOR U23323 ( .A(n23552), .B(n23553), .Z(n23171) );
  AND U23324 ( .A(n392), .B(n23554), .Z(n23553) );
  XOR U23325 ( .A(n23555), .B(n23552), .Z(n23554) );
  XOR U23326 ( .A(n23556), .B(n23557), .Z(n23544) );
  AND U23327 ( .A(n23558), .B(n23559), .Z(n23557) );
  XOR U23328 ( .A(n23556), .B(n23186), .Z(n23559) );
  XOR U23329 ( .A(n23560), .B(n23561), .Z(n23186) );
  AND U23330 ( .A(n394), .B(n23562), .Z(n23561) );
  XOR U23331 ( .A(n23563), .B(n23560), .Z(n23562) );
  XNOR U23332 ( .A(n23183), .B(n23556), .Z(n23558) );
  XOR U23333 ( .A(n23564), .B(n23565), .Z(n23183) );
  AND U23334 ( .A(n392), .B(n23566), .Z(n23565) );
  XOR U23335 ( .A(n23567), .B(n23564), .Z(n23566) );
  XOR U23336 ( .A(n23568), .B(n23569), .Z(n23556) );
  AND U23337 ( .A(n23570), .B(n23571), .Z(n23569) );
  XOR U23338 ( .A(n23568), .B(n23198), .Z(n23571) );
  XOR U23339 ( .A(n23572), .B(n23573), .Z(n23198) );
  AND U23340 ( .A(n394), .B(n23574), .Z(n23573) );
  XOR U23341 ( .A(n23575), .B(n23572), .Z(n23574) );
  XNOR U23342 ( .A(n23195), .B(n23568), .Z(n23570) );
  XOR U23343 ( .A(n23576), .B(n23577), .Z(n23195) );
  AND U23344 ( .A(n392), .B(n23578), .Z(n23577) );
  XOR U23345 ( .A(n23579), .B(n23576), .Z(n23578) );
  XOR U23346 ( .A(n23580), .B(n23581), .Z(n23568) );
  AND U23347 ( .A(n23582), .B(n23583), .Z(n23581) );
  XOR U23348 ( .A(n23580), .B(n23210), .Z(n23583) );
  XOR U23349 ( .A(n23584), .B(n23585), .Z(n23210) );
  AND U23350 ( .A(n394), .B(n23586), .Z(n23585) );
  XOR U23351 ( .A(n23587), .B(n23584), .Z(n23586) );
  XNOR U23352 ( .A(n23207), .B(n23580), .Z(n23582) );
  XOR U23353 ( .A(n23588), .B(n23589), .Z(n23207) );
  AND U23354 ( .A(n392), .B(n23590), .Z(n23589) );
  XOR U23355 ( .A(n23591), .B(n23588), .Z(n23590) );
  XOR U23356 ( .A(n23592), .B(n23593), .Z(n23580) );
  AND U23357 ( .A(n23594), .B(n23595), .Z(n23593) );
  XOR U23358 ( .A(n23592), .B(n23222), .Z(n23595) );
  XOR U23359 ( .A(n23596), .B(n23597), .Z(n23222) );
  AND U23360 ( .A(n394), .B(n23598), .Z(n23597) );
  XOR U23361 ( .A(n23599), .B(n23596), .Z(n23598) );
  XNOR U23362 ( .A(n23219), .B(n23592), .Z(n23594) );
  XOR U23363 ( .A(n23600), .B(n23601), .Z(n23219) );
  AND U23364 ( .A(n392), .B(n23602), .Z(n23601) );
  XOR U23365 ( .A(n23603), .B(n23600), .Z(n23602) );
  XOR U23366 ( .A(n23604), .B(n23605), .Z(n23592) );
  AND U23367 ( .A(n23606), .B(n23607), .Z(n23605) );
  XOR U23368 ( .A(n23234), .B(n23604), .Z(n23607) );
  XOR U23369 ( .A(n23608), .B(n23609), .Z(n23234) );
  AND U23370 ( .A(n394), .B(n23610), .Z(n23609) );
  XOR U23371 ( .A(n23608), .B(n23611), .Z(n23610) );
  XNOR U23372 ( .A(n23604), .B(n23231), .Z(n23606) );
  XOR U23373 ( .A(n23612), .B(n23613), .Z(n23231) );
  AND U23374 ( .A(n392), .B(n23614), .Z(n23613) );
  XOR U23375 ( .A(n23612), .B(n23615), .Z(n23614) );
  XOR U23376 ( .A(n23616), .B(n23617), .Z(n23604) );
  AND U23377 ( .A(n23618), .B(n23619), .Z(n23617) );
  XNOR U23378 ( .A(n23620), .B(n23247), .Z(n23619) );
  XOR U23379 ( .A(n23621), .B(n23622), .Z(n23247) );
  AND U23380 ( .A(n394), .B(n23623), .Z(n23622) );
  XOR U23381 ( .A(n23624), .B(n23621), .Z(n23623) );
  XNOR U23382 ( .A(n23244), .B(n23616), .Z(n23618) );
  XOR U23383 ( .A(n23625), .B(n23626), .Z(n23244) );
  AND U23384 ( .A(n392), .B(n23627), .Z(n23626) );
  XOR U23385 ( .A(n23628), .B(n23625), .Z(n23627) );
  IV U23386 ( .A(n23620), .Z(n23616) );
  AND U23387 ( .A(n23252), .B(n23255), .Z(n23620) );
  XNOR U23388 ( .A(n23629), .B(n23630), .Z(n23255) );
  AND U23389 ( .A(n394), .B(n23631), .Z(n23630) );
  XNOR U23390 ( .A(n23632), .B(n23629), .Z(n23631) );
  XOR U23391 ( .A(n23633), .B(n23634), .Z(n394) );
  AND U23392 ( .A(n23635), .B(n23636), .Z(n23634) );
  XOR U23393 ( .A(n23263), .B(n23633), .Z(n23636) );
  IV U23394 ( .A(n23637), .Z(n23263) );
  AND U23395 ( .A(p_input[991]), .B(p_input[1023]), .Z(n23637) );
  XOR U23396 ( .A(n23633), .B(n23260), .Z(n23635) );
  AND U23397 ( .A(p_input[927]), .B(p_input[959]), .Z(n23260) );
  XOR U23398 ( .A(n23638), .B(n23639), .Z(n23633) );
  AND U23399 ( .A(n23640), .B(n23641), .Z(n23639) );
  XOR U23400 ( .A(n23638), .B(n23275), .Z(n23641) );
  XNOR U23401 ( .A(p_input[990]), .B(n23642), .Z(n23275) );
  AND U23402 ( .A(n550), .B(n23643), .Z(n23642) );
  XOR U23403 ( .A(p_input[990]), .B(p_input[1022]), .Z(n23643) );
  XNOR U23404 ( .A(n23272), .B(n23638), .Z(n23640) );
  XOR U23405 ( .A(n23644), .B(n23645), .Z(n23272) );
  AND U23406 ( .A(n548), .B(n23646), .Z(n23645) );
  XOR U23407 ( .A(p_input[958]), .B(p_input[926]), .Z(n23646) );
  XOR U23408 ( .A(n23647), .B(n23648), .Z(n23638) );
  AND U23409 ( .A(n23649), .B(n23650), .Z(n23648) );
  XOR U23410 ( .A(n23647), .B(n23287), .Z(n23650) );
  XNOR U23411 ( .A(p_input[989]), .B(n23651), .Z(n23287) );
  AND U23412 ( .A(n550), .B(n23652), .Z(n23651) );
  XOR U23413 ( .A(p_input[989]), .B(p_input[1021]), .Z(n23652) );
  XNOR U23414 ( .A(n23284), .B(n23647), .Z(n23649) );
  XOR U23415 ( .A(n23653), .B(n23654), .Z(n23284) );
  AND U23416 ( .A(n548), .B(n23655), .Z(n23654) );
  XOR U23417 ( .A(p_input[957]), .B(p_input[925]), .Z(n23655) );
  XOR U23418 ( .A(n23656), .B(n23657), .Z(n23647) );
  AND U23419 ( .A(n23658), .B(n23659), .Z(n23657) );
  XOR U23420 ( .A(n23656), .B(n23299), .Z(n23659) );
  XNOR U23421 ( .A(p_input[988]), .B(n23660), .Z(n23299) );
  AND U23422 ( .A(n550), .B(n23661), .Z(n23660) );
  XOR U23423 ( .A(p_input[988]), .B(p_input[1020]), .Z(n23661) );
  XNOR U23424 ( .A(n23296), .B(n23656), .Z(n23658) );
  XOR U23425 ( .A(n23662), .B(n23663), .Z(n23296) );
  AND U23426 ( .A(n548), .B(n23664), .Z(n23663) );
  XOR U23427 ( .A(p_input[956]), .B(p_input[924]), .Z(n23664) );
  XOR U23428 ( .A(n23665), .B(n23666), .Z(n23656) );
  AND U23429 ( .A(n23667), .B(n23668), .Z(n23666) );
  XOR U23430 ( .A(n23665), .B(n23311), .Z(n23668) );
  XNOR U23431 ( .A(p_input[987]), .B(n23669), .Z(n23311) );
  AND U23432 ( .A(n550), .B(n23670), .Z(n23669) );
  XOR U23433 ( .A(p_input[987]), .B(p_input[1019]), .Z(n23670) );
  XNOR U23434 ( .A(n23308), .B(n23665), .Z(n23667) );
  XOR U23435 ( .A(n23671), .B(n23672), .Z(n23308) );
  AND U23436 ( .A(n548), .B(n23673), .Z(n23672) );
  XOR U23437 ( .A(p_input[955]), .B(p_input[923]), .Z(n23673) );
  XOR U23438 ( .A(n23674), .B(n23675), .Z(n23665) );
  AND U23439 ( .A(n23676), .B(n23677), .Z(n23675) );
  XOR U23440 ( .A(n23674), .B(n23323), .Z(n23677) );
  XNOR U23441 ( .A(p_input[986]), .B(n23678), .Z(n23323) );
  AND U23442 ( .A(n550), .B(n23679), .Z(n23678) );
  XOR U23443 ( .A(p_input[986]), .B(p_input[1018]), .Z(n23679) );
  XNOR U23444 ( .A(n23320), .B(n23674), .Z(n23676) );
  XOR U23445 ( .A(n23680), .B(n23681), .Z(n23320) );
  AND U23446 ( .A(n548), .B(n23682), .Z(n23681) );
  XOR U23447 ( .A(p_input[954]), .B(p_input[922]), .Z(n23682) );
  XOR U23448 ( .A(n23683), .B(n23684), .Z(n23674) );
  AND U23449 ( .A(n23685), .B(n23686), .Z(n23684) );
  XOR U23450 ( .A(n23683), .B(n23335), .Z(n23686) );
  XNOR U23451 ( .A(p_input[985]), .B(n23687), .Z(n23335) );
  AND U23452 ( .A(n550), .B(n23688), .Z(n23687) );
  XOR U23453 ( .A(p_input[985]), .B(p_input[1017]), .Z(n23688) );
  XNOR U23454 ( .A(n23332), .B(n23683), .Z(n23685) );
  XOR U23455 ( .A(n23689), .B(n23690), .Z(n23332) );
  AND U23456 ( .A(n548), .B(n23691), .Z(n23690) );
  XOR U23457 ( .A(p_input[953]), .B(p_input[921]), .Z(n23691) );
  XOR U23458 ( .A(n23692), .B(n23693), .Z(n23683) );
  AND U23459 ( .A(n23694), .B(n23695), .Z(n23693) );
  XOR U23460 ( .A(n23692), .B(n23347), .Z(n23695) );
  XNOR U23461 ( .A(p_input[984]), .B(n23696), .Z(n23347) );
  AND U23462 ( .A(n550), .B(n23697), .Z(n23696) );
  XOR U23463 ( .A(p_input[984]), .B(p_input[1016]), .Z(n23697) );
  XNOR U23464 ( .A(n23344), .B(n23692), .Z(n23694) );
  XOR U23465 ( .A(n23698), .B(n23699), .Z(n23344) );
  AND U23466 ( .A(n548), .B(n23700), .Z(n23699) );
  XOR U23467 ( .A(p_input[952]), .B(p_input[920]), .Z(n23700) );
  XOR U23468 ( .A(n23701), .B(n23702), .Z(n23692) );
  AND U23469 ( .A(n23703), .B(n23704), .Z(n23702) );
  XOR U23470 ( .A(n23701), .B(n23359), .Z(n23704) );
  XNOR U23471 ( .A(p_input[983]), .B(n23705), .Z(n23359) );
  AND U23472 ( .A(n550), .B(n23706), .Z(n23705) );
  XOR U23473 ( .A(p_input[983]), .B(p_input[1015]), .Z(n23706) );
  XNOR U23474 ( .A(n23356), .B(n23701), .Z(n23703) );
  XOR U23475 ( .A(n23707), .B(n23708), .Z(n23356) );
  AND U23476 ( .A(n548), .B(n23709), .Z(n23708) );
  XOR U23477 ( .A(p_input[951]), .B(p_input[919]), .Z(n23709) );
  XOR U23478 ( .A(n23710), .B(n23711), .Z(n23701) );
  AND U23479 ( .A(n23712), .B(n23713), .Z(n23711) );
  XOR U23480 ( .A(n23710), .B(n23371), .Z(n23713) );
  XNOR U23481 ( .A(p_input[982]), .B(n23714), .Z(n23371) );
  AND U23482 ( .A(n550), .B(n23715), .Z(n23714) );
  XOR U23483 ( .A(p_input[982]), .B(p_input[1014]), .Z(n23715) );
  XNOR U23484 ( .A(n23368), .B(n23710), .Z(n23712) );
  XOR U23485 ( .A(n23716), .B(n23717), .Z(n23368) );
  AND U23486 ( .A(n548), .B(n23718), .Z(n23717) );
  XOR U23487 ( .A(p_input[950]), .B(p_input[918]), .Z(n23718) );
  XOR U23488 ( .A(n23719), .B(n23720), .Z(n23710) );
  AND U23489 ( .A(n23721), .B(n23722), .Z(n23720) );
  XOR U23490 ( .A(n23719), .B(n23383), .Z(n23722) );
  XNOR U23491 ( .A(p_input[981]), .B(n23723), .Z(n23383) );
  AND U23492 ( .A(n550), .B(n23724), .Z(n23723) );
  XOR U23493 ( .A(p_input[981]), .B(p_input[1013]), .Z(n23724) );
  XNOR U23494 ( .A(n23380), .B(n23719), .Z(n23721) );
  XOR U23495 ( .A(n23725), .B(n23726), .Z(n23380) );
  AND U23496 ( .A(n548), .B(n23727), .Z(n23726) );
  XOR U23497 ( .A(p_input[949]), .B(p_input[917]), .Z(n23727) );
  XOR U23498 ( .A(n23728), .B(n23729), .Z(n23719) );
  AND U23499 ( .A(n23730), .B(n23731), .Z(n23729) );
  XOR U23500 ( .A(n23728), .B(n23395), .Z(n23731) );
  XNOR U23501 ( .A(p_input[980]), .B(n23732), .Z(n23395) );
  AND U23502 ( .A(n550), .B(n23733), .Z(n23732) );
  XOR U23503 ( .A(p_input[980]), .B(p_input[1012]), .Z(n23733) );
  XNOR U23504 ( .A(n23392), .B(n23728), .Z(n23730) );
  XOR U23505 ( .A(n23734), .B(n23735), .Z(n23392) );
  AND U23506 ( .A(n548), .B(n23736), .Z(n23735) );
  XOR U23507 ( .A(p_input[948]), .B(p_input[916]), .Z(n23736) );
  XOR U23508 ( .A(n23737), .B(n23738), .Z(n23728) );
  AND U23509 ( .A(n23739), .B(n23740), .Z(n23738) );
  XOR U23510 ( .A(n23737), .B(n23407), .Z(n23740) );
  XNOR U23511 ( .A(p_input[979]), .B(n23741), .Z(n23407) );
  AND U23512 ( .A(n550), .B(n23742), .Z(n23741) );
  XOR U23513 ( .A(p_input[979]), .B(p_input[1011]), .Z(n23742) );
  XNOR U23514 ( .A(n23404), .B(n23737), .Z(n23739) );
  XOR U23515 ( .A(n23743), .B(n23744), .Z(n23404) );
  AND U23516 ( .A(n548), .B(n23745), .Z(n23744) );
  XOR U23517 ( .A(p_input[947]), .B(p_input[915]), .Z(n23745) );
  XOR U23518 ( .A(n23746), .B(n23747), .Z(n23737) );
  AND U23519 ( .A(n23748), .B(n23749), .Z(n23747) );
  XOR U23520 ( .A(n23746), .B(n23419), .Z(n23749) );
  XNOR U23521 ( .A(p_input[978]), .B(n23750), .Z(n23419) );
  AND U23522 ( .A(n550), .B(n23751), .Z(n23750) );
  XOR U23523 ( .A(p_input[978]), .B(p_input[1010]), .Z(n23751) );
  XNOR U23524 ( .A(n23416), .B(n23746), .Z(n23748) );
  XOR U23525 ( .A(n23752), .B(n23753), .Z(n23416) );
  AND U23526 ( .A(n548), .B(n23754), .Z(n23753) );
  XOR U23527 ( .A(p_input[946]), .B(p_input[914]), .Z(n23754) );
  XOR U23528 ( .A(n23755), .B(n23756), .Z(n23746) );
  AND U23529 ( .A(n23757), .B(n23758), .Z(n23756) );
  XOR U23530 ( .A(n23755), .B(n23431), .Z(n23758) );
  XNOR U23531 ( .A(p_input[977]), .B(n23759), .Z(n23431) );
  AND U23532 ( .A(n550), .B(n23760), .Z(n23759) );
  XOR U23533 ( .A(p_input[977]), .B(p_input[1009]), .Z(n23760) );
  XNOR U23534 ( .A(n23428), .B(n23755), .Z(n23757) );
  XOR U23535 ( .A(n23761), .B(n23762), .Z(n23428) );
  AND U23536 ( .A(n548), .B(n23763), .Z(n23762) );
  XOR U23537 ( .A(p_input[945]), .B(p_input[913]), .Z(n23763) );
  XOR U23538 ( .A(n23764), .B(n23765), .Z(n23755) );
  AND U23539 ( .A(n23766), .B(n23767), .Z(n23765) );
  XOR U23540 ( .A(n23764), .B(n23443), .Z(n23767) );
  XNOR U23541 ( .A(p_input[976]), .B(n23768), .Z(n23443) );
  AND U23542 ( .A(n550), .B(n23769), .Z(n23768) );
  XOR U23543 ( .A(p_input[976]), .B(p_input[1008]), .Z(n23769) );
  XNOR U23544 ( .A(n23440), .B(n23764), .Z(n23766) );
  XOR U23545 ( .A(n23770), .B(n23771), .Z(n23440) );
  AND U23546 ( .A(n548), .B(n23772), .Z(n23771) );
  XOR U23547 ( .A(p_input[944]), .B(p_input[912]), .Z(n23772) );
  XOR U23548 ( .A(n23773), .B(n23774), .Z(n23764) );
  AND U23549 ( .A(n23775), .B(n23776), .Z(n23774) );
  XOR U23550 ( .A(n23773), .B(n23455), .Z(n23776) );
  XNOR U23551 ( .A(p_input[975]), .B(n23777), .Z(n23455) );
  AND U23552 ( .A(n550), .B(n23778), .Z(n23777) );
  XOR U23553 ( .A(p_input[975]), .B(p_input[1007]), .Z(n23778) );
  XNOR U23554 ( .A(n23452), .B(n23773), .Z(n23775) );
  XOR U23555 ( .A(n23779), .B(n23780), .Z(n23452) );
  AND U23556 ( .A(n548), .B(n23781), .Z(n23780) );
  XOR U23557 ( .A(p_input[943]), .B(p_input[911]), .Z(n23781) );
  XOR U23558 ( .A(n23782), .B(n23783), .Z(n23773) );
  AND U23559 ( .A(n23784), .B(n23785), .Z(n23783) );
  XOR U23560 ( .A(n23782), .B(n23467), .Z(n23785) );
  XNOR U23561 ( .A(p_input[974]), .B(n23786), .Z(n23467) );
  AND U23562 ( .A(n550), .B(n23787), .Z(n23786) );
  XOR U23563 ( .A(p_input[974]), .B(p_input[1006]), .Z(n23787) );
  XNOR U23564 ( .A(n23464), .B(n23782), .Z(n23784) );
  XOR U23565 ( .A(n23788), .B(n23789), .Z(n23464) );
  AND U23566 ( .A(n548), .B(n23790), .Z(n23789) );
  XOR U23567 ( .A(p_input[942]), .B(p_input[910]), .Z(n23790) );
  XOR U23568 ( .A(n23791), .B(n23792), .Z(n23782) );
  AND U23569 ( .A(n23793), .B(n23794), .Z(n23792) );
  XOR U23570 ( .A(n23791), .B(n23479), .Z(n23794) );
  XNOR U23571 ( .A(p_input[973]), .B(n23795), .Z(n23479) );
  AND U23572 ( .A(n550), .B(n23796), .Z(n23795) );
  XOR U23573 ( .A(p_input[973]), .B(p_input[1005]), .Z(n23796) );
  XNOR U23574 ( .A(n23476), .B(n23791), .Z(n23793) );
  XOR U23575 ( .A(n23797), .B(n23798), .Z(n23476) );
  AND U23576 ( .A(n548), .B(n23799), .Z(n23798) );
  XOR U23577 ( .A(p_input[941]), .B(p_input[909]), .Z(n23799) );
  XOR U23578 ( .A(n23800), .B(n23801), .Z(n23791) );
  AND U23579 ( .A(n23802), .B(n23803), .Z(n23801) );
  XOR U23580 ( .A(n23800), .B(n23491), .Z(n23803) );
  XNOR U23581 ( .A(p_input[972]), .B(n23804), .Z(n23491) );
  AND U23582 ( .A(n550), .B(n23805), .Z(n23804) );
  XOR U23583 ( .A(p_input[972]), .B(p_input[1004]), .Z(n23805) );
  XNOR U23584 ( .A(n23488), .B(n23800), .Z(n23802) );
  XOR U23585 ( .A(n23806), .B(n23807), .Z(n23488) );
  AND U23586 ( .A(n548), .B(n23808), .Z(n23807) );
  XOR U23587 ( .A(p_input[940]), .B(p_input[908]), .Z(n23808) );
  XOR U23588 ( .A(n23809), .B(n23810), .Z(n23800) );
  AND U23589 ( .A(n23811), .B(n23812), .Z(n23810) );
  XOR U23590 ( .A(n23809), .B(n23503), .Z(n23812) );
  XNOR U23591 ( .A(p_input[971]), .B(n23813), .Z(n23503) );
  AND U23592 ( .A(n550), .B(n23814), .Z(n23813) );
  XOR U23593 ( .A(p_input[971]), .B(p_input[1003]), .Z(n23814) );
  XNOR U23594 ( .A(n23500), .B(n23809), .Z(n23811) );
  XOR U23595 ( .A(n23815), .B(n23816), .Z(n23500) );
  AND U23596 ( .A(n548), .B(n23817), .Z(n23816) );
  XOR U23597 ( .A(p_input[939]), .B(p_input[907]), .Z(n23817) );
  XOR U23598 ( .A(n23818), .B(n23819), .Z(n23809) );
  AND U23599 ( .A(n23820), .B(n23821), .Z(n23819) );
  XOR U23600 ( .A(n23818), .B(n23515), .Z(n23821) );
  XNOR U23601 ( .A(p_input[970]), .B(n23822), .Z(n23515) );
  AND U23602 ( .A(n550), .B(n23823), .Z(n23822) );
  XOR U23603 ( .A(p_input[970]), .B(p_input[1002]), .Z(n23823) );
  XNOR U23604 ( .A(n23512), .B(n23818), .Z(n23820) );
  XOR U23605 ( .A(n23824), .B(n23825), .Z(n23512) );
  AND U23606 ( .A(n548), .B(n23826), .Z(n23825) );
  XOR U23607 ( .A(p_input[938]), .B(p_input[906]), .Z(n23826) );
  XOR U23608 ( .A(n23827), .B(n23828), .Z(n23818) );
  AND U23609 ( .A(n23829), .B(n23830), .Z(n23828) );
  XOR U23610 ( .A(n23827), .B(n23527), .Z(n23830) );
  XNOR U23611 ( .A(p_input[969]), .B(n23831), .Z(n23527) );
  AND U23612 ( .A(n550), .B(n23832), .Z(n23831) );
  XOR U23613 ( .A(p_input[969]), .B(p_input[1001]), .Z(n23832) );
  XNOR U23614 ( .A(n23524), .B(n23827), .Z(n23829) );
  XOR U23615 ( .A(n23833), .B(n23834), .Z(n23524) );
  AND U23616 ( .A(n548), .B(n23835), .Z(n23834) );
  XOR U23617 ( .A(p_input[937]), .B(p_input[905]), .Z(n23835) );
  XOR U23618 ( .A(n23836), .B(n23837), .Z(n23827) );
  AND U23619 ( .A(n23838), .B(n23839), .Z(n23837) );
  XOR U23620 ( .A(n23836), .B(n23539), .Z(n23839) );
  XNOR U23621 ( .A(p_input[968]), .B(n23840), .Z(n23539) );
  AND U23622 ( .A(n550), .B(n23841), .Z(n23840) );
  XOR U23623 ( .A(p_input[968]), .B(p_input[1000]), .Z(n23841) );
  XNOR U23624 ( .A(n23536), .B(n23836), .Z(n23838) );
  XOR U23625 ( .A(n23842), .B(n23843), .Z(n23536) );
  AND U23626 ( .A(n548), .B(n23844), .Z(n23843) );
  XOR U23627 ( .A(p_input[936]), .B(p_input[904]), .Z(n23844) );
  XOR U23628 ( .A(n23845), .B(n23846), .Z(n23836) );
  AND U23629 ( .A(n23847), .B(n23848), .Z(n23846) );
  XOR U23630 ( .A(n23845), .B(n23551), .Z(n23848) );
  XNOR U23631 ( .A(p_input[967]), .B(n23849), .Z(n23551) );
  AND U23632 ( .A(n550), .B(n23850), .Z(n23849) );
  XOR U23633 ( .A(p_input[999]), .B(p_input[967]), .Z(n23850) );
  XNOR U23634 ( .A(n23548), .B(n23845), .Z(n23847) );
  XOR U23635 ( .A(n23851), .B(n23852), .Z(n23548) );
  AND U23636 ( .A(n548), .B(n23853), .Z(n23852) );
  XOR U23637 ( .A(p_input[935]), .B(p_input[903]), .Z(n23853) );
  XOR U23638 ( .A(n23854), .B(n23855), .Z(n23845) );
  AND U23639 ( .A(n23856), .B(n23857), .Z(n23855) );
  XOR U23640 ( .A(n23854), .B(n23563), .Z(n23857) );
  XNOR U23641 ( .A(p_input[966]), .B(n23858), .Z(n23563) );
  AND U23642 ( .A(n550), .B(n23859), .Z(n23858) );
  XOR U23643 ( .A(p_input[998]), .B(p_input[966]), .Z(n23859) );
  XNOR U23644 ( .A(n23560), .B(n23854), .Z(n23856) );
  XOR U23645 ( .A(n23860), .B(n23861), .Z(n23560) );
  AND U23646 ( .A(n548), .B(n23862), .Z(n23861) );
  XOR U23647 ( .A(p_input[934]), .B(p_input[902]), .Z(n23862) );
  XOR U23648 ( .A(n23863), .B(n23864), .Z(n23854) );
  AND U23649 ( .A(n23865), .B(n23866), .Z(n23864) );
  XOR U23650 ( .A(n23863), .B(n23575), .Z(n23866) );
  XNOR U23651 ( .A(p_input[965]), .B(n23867), .Z(n23575) );
  AND U23652 ( .A(n550), .B(n23868), .Z(n23867) );
  XOR U23653 ( .A(p_input[997]), .B(p_input[965]), .Z(n23868) );
  XNOR U23654 ( .A(n23572), .B(n23863), .Z(n23865) );
  XOR U23655 ( .A(n23869), .B(n23870), .Z(n23572) );
  AND U23656 ( .A(n548), .B(n23871), .Z(n23870) );
  XOR U23657 ( .A(p_input[933]), .B(p_input[901]), .Z(n23871) );
  XOR U23658 ( .A(n23872), .B(n23873), .Z(n23863) );
  AND U23659 ( .A(n23874), .B(n23875), .Z(n23873) );
  XOR U23660 ( .A(n23872), .B(n23587), .Z(n23875) );
  XNOR U23661 ( .A(p_input[964]), .B(n23876), .Z(n23587) );
  AND U23662 ( .A(n550), .B(n23877), .Z(n23876) );
  XOR U23663 ( .A(p_input[996]), .B(p_input[964]), .Z(n23877) );
  XNOR U23664 ( .A(n23584), .B(n23872), .Z(n23874) );
  XOR U23665 ( .A(n23878), .B(n23879), .Z(n23584) );
  AND U23666 ( .A(n548), .B(n23880), .Z(n23879) );
  XOR U23667 ( .A(p_input[932]), .B(p_input[900]), .Z(n23880) );
  XOR U23668 ( .A(n23881), .B(n23882), .Z(n23872) );
  AND U23669 ( .A(n23883), .B(n23884), .Z(n23882) );
  XOR U23670 ( .A(n23881), .B(n23599), .Z(n23884) );
  XNOR U23671 ( .A(p_input[963]), .B(n23885), .Z(n23599) );
  AND U23672 ( .A(n550), .B(n23886), .Z(n23885) );
  XOR U23673 ( .A(p_input[995]), .B(p_input[963]), .Z(n23886) );
  XNOR U23674 ( .A(n23596), .B(n23881), .Z(n23883) );
  XOR U23675 ( .A(n23887), .B(n23888), .Z(n23596) );
  AND U23676 ( .A(n548), .B(n23889), .Z(n23888) );
  XOR U23677 ( .A(p_input[931]), .B(p_input[899]), .Z(n23889) );
  XOR U23678 ( .A(n23890), .B(n23891), .Z(n23881) );
  AND U23679 ( .A(n23892), .B(n23893), .Z(n23891) );
  XOR U23680 ( .A(n23611), .B(n23890), .Z(n23893) );
  XNOR U23681 ( .A(p_input[962]), .B(n23894), .Z(n23611) );
  AND U23682 ( .A(n550), .B(n23895), .Z(n23894) );
  XOR U23683 ( .A(p_input[994]), .B(p_input[962]), .Z(n23895) );
  XNOR U23684 ( .A(n23890), .B(n23608), .Z(n23892) );
  XOR U23685 ( .A(n23896), .B(n23897), .Z(n23608) );
  AND U23686 ( .A(n548), .B(n23898), .Z(n23897) );
  XOR U23687 ( .A(p_input[930]), .B(p_input[898]), .Z(n23898) );
  XOR U23688 ( .A(n23899), .B(n23900), .Z(n23890) );
  AND U23689 ( .A(n23901), .B(n23902), .Z(n23900) );
  XNOR U23690 ( .A(n23903), .B(n23624), .Z(n23902) );
  XNOR U23691 ( .A(p_input[961]), .B(n23904), .Z(n23624) );
  AND U23692 ( .A(n550), .B(n23905), .Z(n23904) );
  XNOR U23693 ( .A(p_input[993]), .B(n23906), .Z(n23905) );
  IV U23694 ( .A(p_input[961]), .Z(n23906) );
  XNOR U23695 ( .A(n23621), .B(n23899), .Z(n23901) );
  XNOR U23696 ( .A(p_input[897]), .B(n23907), .Z(n23621) );
  AND U23697 ( .A(n548), .B(n23908), .Z(n23907) );
  XOR U23698 ( .A(p_input[929]), .B(p_input[897]), .Z(n23908) );
  IV U23699 ( .A(n23903), .Z(n23899) );
  AND U23700 ( .A(n23629), .B(n23632), .Z(n23903) );
  XOR U23701 ( .A(p_input[960]), .B(n23909), .Z(n23632) );
  AND U23702 ( .A(n550), .B(n23910), .Z(n23909) );
  XOR U23703 ( .A(p_input[992]), .B(p_input[960]), .Z(n23910) );
  XOR U23704 ( .A(n23911), .B(n23912), .Z(n550) );
  AND U23705 ( .A(n23913), .B(n23914), .Z(n23912) );
  XNOR U23706 ( .A(p_input[1023]), .B(n23911), .Z(n23914) );
  XOR U23707 ( .A(n23911), .B(p_input[991]), .Z(n23913) );
  XOR U23708 ( .A(n23915), .B(n23916), .Z(n23911) );
  AND U23709 ( .A(n23917), .B(n23918), .Z(n23916) );
  XNOR U23710 ( .A(p_input[1022]), .B(n23915), .Z(n23918) );
  XOR U23711 ( .A(n23915), .B(p_input[990]), .Z(n23917) );
  XOR U23712 ( .A(n23919), .B(n23920), .Z(n23915) );
  AND U23713 ( .A(n23921), .B(n23922), .Z(n23920) );
  XNOR U23714 ( .A(p_input[1021]), .B(n23919), .Z(n23922) );
  XOR U23715 ( .A(n23919), .B(p_input[989]), .Z(n23921) );
  XOR U23716 ( .A(n23923), .B(n23924), .Z(n23919) );
  AND U23717 ( .A(n23925), .B(n23926), .Z(n23924) );
  XNOR U23718 ( .A(p_input[1020]), .B(n23923), .Z(n23926) );
  XOR U23719 ( .A(n23923), .B(p_input[988]), .Z(n23925) );
  XOR U23720 ( .A(n23927), .B(n23928), .Z(n23923) );
  AND U23721 ( .A(n23929), .B(n23930), .Z(n23928) );
  XNOR U23722 ( .A(p_input[1019]), .B(n23927), .Z(n23930) );
  XOR U23723 ( .A(n23927), .B(p_input[987]), .Z(n23929) );
  XOR U23724 ( .A(n23931), .B(n23932), .Z(n23927) );
  AND U23725 ( .A(n23933), .B(n23934), .Z(n23932) );
  XNOR U23726 ( .A(p_input[1018]), .B(n23931), .Z(n23934) );
  XOR U23727 ( .A(n23931), .B(p_input[986]), .Z(n23933) );
  XOR U23728 ( .A(n23935), .B(n23936), .Z(n23931) );
  AND U23729 ( .A(n23937), .B(n23938), .Z(n23936) );
  XNOR U23730 ( .A(p_input[1017]), .B(n23935), .Z(n23938) );
  XOR U23731 ( .A(n23935), .B(p_input[985]), .Z(n23937) );
  XOR U23732 ( .A(n23939), .B(n23940), .Z(n23935) );
  AND U23733 ( .A(n23941), .B(n23942), .Z(n23940) );
  XNOR U23734 ( .A(p_input[1016]), .B(n23939), .Z(n23942) );
  XOR U23735 ( .A(n23939), .B(p_input[984]), .Z(n23941) );
  XOR U23736 ( .A(n23943), .B(n23944), .Z(n23939) );
  AND U23737 ( .A(n23945), .B(n23946), .Z(n23944) );
  XNOR U23738 ( .A(p_input[1015]), .B(n23943), .Z(n23946) );
  XOR U23739 ( .A(n23943), .B(p_input[983]), .Z(n23945) );
  XOR U23740 ( .A(n23947), .B(n23948), .Z(n23943) );
  AND U23741 ( .A(n23949), .B(n23950), .Z(n23948) );
  XNOR U23742 ( .A(p_input[1014]), .B(n23947), .Z(n23950) );
  XOR U23743 ( .A(n23947), .B(p_input[982]), .Z(n23949) );
  XOR U23744 ( .A(n23951), .B(n23952), .Z(n23947) );
  AND U23745 ( .A(n23953), .B(n23954), .Z(n23952) );
  XNOR U23746 ( .A(p_input[1013]), .B(n23951), .Z(n23954) );
  XOR U23747 ( .A(n23951), .B(p_input[981]), .Z(n23953) );
  XOR U23748 ( .A(n23955), .B(n23956), .Z(n23951) );
  AND U23749 ( .A(n23957), .B(n23958), .Z(n23956) );
  XNOR U23750 ( .A(p_input[1012]), .B(n23955), .Z(n23958) );
  XOR U23751 ( .A(n23955), .B(p_input[980]), .Z(n23957) );
  XOR U23752 ( .A(n23959), .B(n23960), .Z(n23955) );
  AND U23753 ( .A(n23961), .B(n23962), .Z(n23960) );
  XNOR U23754 ( .A(p_input[1011]), .B(n23959), .Z(n23962) );
  XOR U23755 ( .A(n23959), .B(p_input[979]), .Z(n23961) );
  XOR U23756 ( .A(n23963), .B(n23964), .Z(n23959) );
  AND U23757 ( .A(n23965), .B(n23966), .Z(n23964) );
  XNOR U23758 ( .A(p_input[1010]), .B(n23963), .Z(n23966) );
  XOR U23759 ( .A(n23963), .B(p_input[978]), .Z(n23965) );
  XOR U23760 ( .A(n23967), .B(n23968), .Z(n23963) );
  AND U23761 ( .A(n23969), .B(n23970), .Z(n23968) );
  XNOR U23762 ( .A(p_input[1009]), .B(n23967), .Z(n23970) );
  XOR U23763 ( .A(n23967), .B(p_input[977]), .Z(n23969) );
  XOR U23764 ( .A(n23971), .B(n23972), .Z(n23967) );
  AND U23765 ( .A(n23973), .B(n23974), .Z(n23972) );
  XNOR U23766 ( .A(p_input[1008]), .B(n23971), .Z(n23974) );
  XOR U23767 ( .A(n23971), .B(p_input[976]), .Z(n23973) );
  XOR U23768 ( .A(n23975), .B(n23976), .Z(n23971) );
  AND U23769 ( .A(n23977), .B(n23978), .Z(n23976) );
  XNOR U23770 ( .A(p_input[1007]), .B(n23975), .Z(n23978) );
  XOR U23771 ( .A(n23975), .B(p_input[975]), .Z(n23977) );
  XOR U23772 ( .A(n23979), .B(n23980), .Z(n23975) );
  AND U23773 ( .A(n23981), .B(n23982), .Z(n23980) );
  XNOR U23774 ( .A(p_input[1006]), .B(n23979), .Z(n23982) );
  XOR U23775 ( .A(n23979), .B(p_input[974]), .Z(n23981) );
  XOR U23776 ( .A(n23983), .B(n23984), .Z(n23979) );
  AND U23777 ( .A(n23985), .B(n23986), .Z(n23984) );
  XNOR U23778 ( .A(p_input[1005]), .B(n23983), .Z(n23986) );
  XOR U23779 ( .A(n23983), .B(p_input[973]), .Z(n23985) );
  XOR U23780 ( .A(n23987), .B(n23988), .Z(n23983) );
  AND U23781 ( .A(n23989), .B(n23990), .Z(n23988) );
  XNOR U23782 ( .A(p_input[1004]), .B(n23987), .Z(n23990) );
  XOR U23783 ( .A(n23987), .B(p_input[972]), .Z(n23989) );
  XOR U23784 ( .A(n23991), .B(n23992), .Z(n23987) );
  AND U23785 ( .A(n23993), .B(n23994), .Z(n23992) );
  XNOR U23786 ( .A(p_input[1003]), .B(n23991), .Z(n23994) );
  XOR U23787 ( .A(n23991), .B(p_input[971]), .Z(n23993) );
  XOR U23788 ( .A(n23995), .B(n23996), .Z(n23991) );
  AND U23789 ( .A(n23997), .B(n23998), .Z(n23996) );
  XNOR U23790 ( .A(p_input[1002]), .B(n23995), .Z(n23998) );
  XOR U23791 ( .A(n23995), .B(p_input[970]), .Z(n23997) );
  XOR U23792 ( .A(n23999), .B(n24000), .Z(n23995) );
  AND U23793 ( .A(n24001), .B(n24002), .Z(n24000) );
  XNOR U23794 ( .A(p_input[1001]), .B(n23999), .Z(n24002) );
  XOR U23795 ( .A(n23999), .B(p_input[969]), .Z(n24001) );
  XOR U23796 ( .A(n24003), .B(n24004), .Z(n23999) );
  AND U23797 ( .A(n24005), .B(n24006), .Z(n24004) );
  XNOR U23798 ( .A(p_input[1000]), .B(n24003), .Z(n24006) );
  XOR U23799 ( .A(n24003), .B(p_input[968]), .Z(n24005) );
  XOR U23800 ( .A(n24007), .B(n24008), .Z(n24003) );
  AND U23801 ( .A(n24009), .B(n24010), .Z(n24008) );
  XNOR U23802 ( .A(p_input[999]), .B(n24007), .Z(n24010) );
  XOR U23803 ( .A(n24007), .B(p_input[967]), .Z(n24009) );
  XOR U23804 ( .A(n24011), .B(n24012), .Z(n24007) );
  AND U23805 ( .A(n24013), .B(n24014), .Z(n24012) );
  XNOR U23806 ( .A(p_input[998]), .B(n24011), .Z(n24014) );
  XOR U23807 ( .A(n24011), .B(p_input[966]), .Z(n24013) );
  XOR U23808 ( .A(n24015), .B(n24016), .Z(n24011) );
  AND U23809 ( .A(n24017), .B(n24018), .Z(n24016) );
  XNOR U23810 ( .A(p_input[997]), .B(n24015), .Z(n24018) );
  XOR U23811 ( .A(n24015), .B(p_input[965]), .Z(n24017) );
  XOR U23812 ( .A(n24019), .B(n24020), .Z(n24015) );
  AND U23813 ( .A(n24021), .B(n24022), .Z(n24020) );
  XNOR U23814 ( .A(p_input[996]), .B(n24019), .Z(n24022) );
  XOR U23815 ( .A(n24019), .B(p_input[964]), .Z(n24021) );
  XOR U23816 ( .A(n24023), .B(n24024), .Z(n24019) );
  AND U23817 ( .A(n24025), .B(n24026), .Z(n24024) );
  XNOR U23818 ( .A(p_input[995]), .B(n24023), .Z(n24026) );
  XOR U23819 ( .A(n24023), .B(p_input[963]), .Z(n24025) );
  XOR U23820 ( .A(n24027), .B(n24028), .Z(n24023) );
  AND U23821 ( .A(n24029), .B(n24030), .Z(n24028) );
  XNOR U23822 ( .A(p_input[994]), .B(n24027), .Z(n24030) );
  XOR U23823 ( .A(n24027), .B(p_input[962]), .Z(n24029) );
  XNOR U23824 ( .A(n24031), .B(n24032), .Z(n24027) );
  AND U23825 ( .A(n24033), .B(n24034), .Z(n24032) );
  XOR U23826 ( .A(p_input[993]), .B(n24031), .Z(n24034) );
  XNOR U23827 ( .A(p_input[961]), .B(n24031), .Z(n24033) );
  AND U23828 ( .A(p_input[992]), .B(n24035), .Z(n24031) );
  IV U23829 ( .A(p_input[960]), .Z(n24035) );
  XNOR U23830 ( .A(p_input[896]), .B(n24036), .Z(n23629) );
  AND U23831 ( .A(n548), .B(n24037), .Z(n24036) );
  XOR U23832 ( .A(p_input[928]), .B(p_input[896]), .Z(n24037) );
  XOR U23833 ( .A(n24038), .B(n24039), .Z(n548) );
  AND U23834 ( .A(n24040), .B(n24041), .Z(n24039) );
  XNOR U23835 ( .A(p_input[959]), .B(n24038), .Z(n24041) );
  XOR U23836 ( .A(n24038), .B(p_input[927]), .Z(n24040) );
  XOR U23837 ( .A(n24042), .B(n24043), .Z(n24038) );
  AND U23838 ( .A(n24044), .B(n24045), .Z(n24043) );
  XNOR U23839 ( .A(p_input[958]), .B(n24042), .Z(n24045) );
  XNOR U23840 ( .A(n24042), .B(n23644), .Z(n24044) );
  IV U23841 ( .A(p_input[926]), .Z(n23644) );
  XOR U23842 ( .A(n24046), .B(n24047), .Z(n24042) );
  AND U23843 ( .A(n24048), .B(n24049), .Z(n24047) );
  XNOR U23844 ( .A(p_input[957]), .B(n24046), .Z(n24049) );
  XNOR U23845 ( .A(n24046), .B(n23653), .Z(n24048) );
  IV U23846 ( .A(p_input[925]), .Z(n23653) );
  XOR U23847 ( .A(n24050), .B(n24051), .Z(n24046) );
  AND U23848 ( .A(n24052), .B(n24053), .Z(n24051) );
  XNOR U23849 ( .A(p_input[956]), .B(n24050), .Z(n24053) );
  XNOR U23850 ( .A(n24050), .B(n23662), .Z(n24052) );
  IV U23851 ( .A(p_input[924]), .Z(n23662) );
  XOR U23852 ( .A(n24054), .B(n24055), .Z(n24050) );
  AND U23853 ( .A(n24056), .B(n24057), .Z(n24055) );
  XNOR U23854 ( .A(p_input[955]), .B(n24054), .Z(n24057) );
  XNOR U23855 ( .A(n24054), .B(n23671), .Z(n24056) );
  IV U23856 ( .A(p_input[923]), .Z(n23671) );
  XOR U23857 ( .A(n24058), .B(n24059), .Z(n24054) );
  AND U23858 ( .A(n24060), .B(n24061), .Z(n24059) );
  XNOR U23859 ( .A(p_input[954]), .B(n24058), .Z(n24061) );
  XNOR U23860 ( .A(n24058), .B(n23680), .Z(n24060) );
  IV U23861 ( .A(p_input[922]), .Z(n23680) );
  XOR U23862 ( .A(n24062), .B(n24063), .Z(n24058) );
  AND U23863 ( .A(n24064), .B(n24065), .Z(n24063) );
  XNOR U23864 ( .A(p_input[953]), .B(n24062), .Z(n24065) );
  XNOR U23865 ( .A(n24062), .B(n23689), .Z(n24064) );
  IV U23866 ( .A(p_input[921]), .Z(n23689) );
  XOR U23867 ( .A(n24066), .B(n24067), .Z(n24062) );
  AND U23868 ( .A(n24068), .B(n24069), .Z(n24067) );
  XNOR U23869 ( .A(p_input[952]), .B(n24066), .Z(n24069) );
  XNOR U23870 ( .A(n24066), .B(n23698), .Z(n24068) );
  IV U23871 ( .A(p_input[920]), .Z(n23698) );
  XOR U23872 ( .A(n24070), .B(n24071), .Z(n24066) );
  AND U23873 ( .A(n24072), .B(n24073), .Z(n24071) );
  XNOR U23874 ( .A(p_input[951]), .B(n24070), .Z(n24073) );
  XNOR U23875 ( .A(n24070), .B(n23707), .Z(n24072) );
  IV U23876 ( .A(p_input[919]), .Z(n23707) );
  XOR U23877 ( .A(n24074), .B(n24075), .Z(n24070) );
  AND U23878 ( .A(n24076), .B(n24077), .Z(n24075) );
  XNOR U23879 ( .A(p_input[950]), .B(n24074), .Z(n24077) );
  XNOR U23880 ( .A(n24074), .B(n23716), .Z(n24076) );
  IV U23881 ( .A(p_input[918]), .Z(n23716) );
  XOR U23882 ( .A(n24078), .B(n24079), .Z(n24074) );
  AND U23883 ( .A(n24080), .B(n24081), .Z(n24079) );
  XNOR U23884 ( .A(p_input[949]), .B(n24078), .Z(n24081) );
  XNOR U23885 ( .A(n24078), .B(n23725), .Z(n24080) );
  IV U23886 ( .A(p_input[917]), .Z(n23725) );
  XOR U23887 ( .A(n24082), .B(n24083), .Z(n24078) );
  AND U23888 ( .A(n24084), .B(n24085), .Z(n24083) );
  XNOR U23889 ( .A(p_input[948]), .B(n24082), .Z(n24085) );
  XNOR U23890 ( .A(n24082), .B(n23734), .Z(n24084) );
  IV U23891 ( .A(p_input[916]), .Z(n23734) );
  XOR U23892 ( .A(n24086), .B(n24087), .Z(n24082) );
  AND U23893 ( .A(n24088), .B(n24089), .Z(n24087) );
  XNOR U23894 ( .A(p_input[947]), .B(n24086), .Z(n24089) );
  XNOR U23895 ( .A(n24086), .B(n23743), .Z(n24088) );
  IV U23896 ( .A(p_input[915]), .Z(n23743) );
  XOR U23897 ( .A(n24090), .B(n24091), .Z(n24086) );
  AND U23898 ( .A(n24092), .B(n24093), .Z(n24091) );
  XNOR U23899 ( .A(p_input[946]), .B(n24090), .Z(n24093) );
  XNOR U23900 ( .A(n24090), .B(n23752), .Z(n24092) );
  IV U23901 ( .A(p_input[914]), .Z(n23752) );
  XOR U23902 ( .A(n24094), .B(n24095), .Z(n24090) );
  AND U23903 ( .A(n24096), .B(n24097), .Z(n24095) );
  XNOR U23904 ( .A(p_input[945]), .B(n24094), .Z(n24097) );
  XNOR U23905 ( .A(n24094), .B(n23761), .Z(n24096) );
  IV U23906 ( .A(p_input[913]), .Z(n23761) );
  XOR U23907 ( .A(n24098), .B(n24099), .Z(n24094) );
  AND U23908 ( .A(n24100), .B(n24101), .Z(n24099) );
  XNOR U23909 ( .A(p_input[944]), .B(n24098), .Z(n24101) );
  XNOR U23910 ( .A(n24098), .B(n23770), .Z(n24100) );
  IV U23911 ( .A(p_input[912]), .Z(n23770) );
  XOR U23912 ( .A(n24102), .B(n24103), .Z(n24098) );
  AND U23913 ( .A(n24104), .B(n24105), .Z(n24103) );
  XNOR U23914 ( .A(p_input[943]), .B(n24102), .Z(n24105) );
  XNOR U23915 ( .A(n24102), .B(n23779), .Z(n24104) );
  IV U23916 ( .A(p_input[911]), .Z(n23779) );
  XOR U23917 ( .A(n24106), .B(n24107), .Z(n24102) );
  AND U23918 ( .A(n24108), .B(n24109), .Z(n24107) );
  XNOR U23919 ( .A(p_input[942]), .B(n24106), .Z(n24109) );
  XNOR U23920 ( .A(n24106), .B(n23788), .Z(n24108) );
  IV U23921 ( .A(p_input[910]), .Z(n23788) );
  XOR U23922 ( .A(n24110), .B(n24111), .Z(n24106) );
  AND U23923 ( .A(n24112), .B(n24113), .Z(n24111) );
  XNOR U23924 ( .A(p_input[941]), .B(n24110), .Z(n24113) );
  XNOR U23925 ( .A(n24110), .B(n23797), .Z(n24112) );
  IV U23926 ( .A(p_input[909]), .Z(n23797) );
  XOR U23927 ( .A(n24114), .B(n24115), .Z(n24110) );
  AND U23928 ( .A(n24116), .B(n24117), .Z(n24115) );
  XNOR U23929 ( .A(p_input[940]), .B(n24114), .Z(n24117) );
  XNOR U23930 ( .A(n24114), .B(n23806), .Z(n24116) );
  IV U23931 ( .A(p_input[908]), .Z(n23806) );
  XOR U23932 ( .A(n24118), .B(n24119), .Z(n24114) );
  AND U23933 ( .A(n24120), .B(n24121), .Z(n24119) );
  XNOR U23934 ( .A(p_input[939]), .B(n24118), .Z(n24121) );
  XNOR U23935 ( .A(n24118), .B(n23815), .Z(n24120) );
  IV U23936 ( .A(p_input[907]), .Z(n23815) );
  XOR U23937 ( .A(n24122), .B(n24123), .Z(n24118) );
  AND U23938 ( .A(n24124), .B(n24125), .Z(n24123) );
  XNOR U23939 ( .A(p_input[938]), .B(n24122), .Z(n24125) );
  XNOR U23940 ( .A(n24122), .B(n23824), .Z(n24124) );
  IV U23941 ( .A(p_input[906]), .Z(n23824) );
  XOR U23942 ( .A(n24126), .B(n24127), .Z(n24122) );
  AND U23943 ( .A(n24128), .B(n24129), .Z(n24127) );
  XNOR U23944 ( .A(p_input[937]), .B(n24126), .Z(n24129) );
  XNOR U23945 ( .A(n24126), .B(n23833), .Z(n24128) );
  IV U23946 ( .A(p_input[905]), .Z(n23833) );
  XOR U23947 ( .A(n24130), .B(n24131), .Z(n24126) );
  AND U23948 ( .A(n24132), .B(n24133), .Z(n24131) );
  XNOR U23949 ( .A(p_input[936]), .B(n24130), .Z(n24133) );
  XNOR U23950 ( .A(n24130), .B(n23842), .Z(n24132) );
  IV U23951 ( .A(p_input[904]), .Z(n23842) );
  XOR U23952 ( .A(n24134), .B(n24135), .Z(n24130) );
  AND U23953 ( .A(n24136), .B(n24137), .Z(n24135) );
  XNOR U23954 ( .A(p_input[935]), .B(n24134), .Z(n24137) );
  XNOR U23955 ( .A(n24134), .B(n23851), .Z(n24136) );
  IV U23956 ( .A(p_input[903]), .Z(n23851) );
  XOR U23957 ( .A(n24138), .B(n24139), .Z(n24134) );
  AND U23958 ( .A(n24140), .B(n24141), .Z(n24139) );
  XNOR U23959 ( .A(p_input[934]), .B(n24138), .Z(n24141) );
  XNOR U23960 ( .A(n24138), .B(n23860), .Z(n24140) );
  IV U23961 ( .A(p_input[902]), .Z(n23860) );
  XOR U23962 ( .A(n24142), .B(n24143), .Z(n24138) );
  AND U23963 ( .A(n24144), .B(n24145), .Z(n24143) );
  XNOR U23964 ( .A(p_input[933]), .B(n24142), .Z(n24145) );
  XNOR U23965 ( .A(n24142), .B(n23869), .Z(n24144) );
  IV U23966 ( .A(p_input[901]), .Z(n23869) );
  XOR U23967 ( .A(n24146), .B(n24147), .Z(n24142) );
  AND U23968 ( .A(n24148), .B(n24149), .Z(n24147) );
  XNOR U23969 ( .A(p_input[932]), .B(n24146), .Z(n24149) );
  XNOR U23970 ( .A(n24146), .B(n23878), .Z(n24148) );
  IV U23971 ( .A(p_input[900]), .Z(n23878) );
  XOR U23972 ( .A(n24150), .B(n24151), .Z(n24146) );
  AND U23973 ( .A(n24152), .B(n24153), .Z(n24151) );
  XNOR U23974 ( .A(p_input[931]), .B(n24150), .Z(n24153) );
  XNOR U23975 ( .A(n24150), .B(n23887), .Z(n24152) );
  IV U23976 ( .A(p_input[899]), .Z(n23887) );
  XOR U23977 ( .A(n24154), .B(n24155), .Z(n24150) );
  AND U23978 ( .A(n24156), .B(n24157), .Z(n24155) );
  XNOR U23979 ( .A(p_input[930]), .B(n24154), .Z(n24157) );
  XNOR U23980 ( .A(n24154), .B(n23896), .Z(n24156) );
  IV U23981 ( .A(p_input[898]), .Z(n23896) );
  XNOR U23982 ( .A(n24158), .B(n24159), .Z(n24154) );
  AND U23983 ( .A(n24160), .B(n24161), .Z(n24159) );
  XOR U23984 ( .A(p_input[929]), .B(n24158), .Z(n24161) );
  XNOR U23985 ( .A(p_input[897]), .B(n24158), .Z(n24160) );
  AND U23986 ( .A(p_input[928]), .B(n24162), .Z(n24158) );
  IV U23987 ( .A(p_input[896]), .Z(n24162) );
  XOR U23988 ( .A(n24163), .B(n24164), .Z(n23252) );
  AND U23989 ( .A(n392), .B(n24165), .Z(n24164) );
  XNOR U23990 ( .A(n24166), .B(n24163), .Z(n24165) );
  XOR U23991 ( .A(n24167), .B(n24168), .Z(n392) );
  AND U23992 ( .A(n24169), .B(n24170), .Z(n24168) );
  XNOR U23993 ( .A(n23267), .B(n24167), .Z(n24170) );
  AND U23994 ( .A(p_input[895]), .B(p_input[863]), .Z(n23267) );
  XNOR U23995 ( .A(n24167), .B(n23264), .Z(n24169) );
  IV U23996 ( .A(n24171), .Z(n23264) );
  AND U23997 ( .A(p_input[799]), .B(p_input[831]), .Z(n24171) );
  XOR U23998 ( .A(n24172), .B(n24173), .Z(n24167) );
  AND U23999 ( .A(n24174), .B(n24175), .Z(n24173) );
  XOR U24000 ( .A(n24172), .B(n23279), .Z(n24175) );
  XNOR U24001 ( .A(p_input[862]), .B(n24176), .Z(n23279) );
  AND U24002 ( .A(n554), .B(n24177), .Z(n24176) );
  XOR U24003 ( .A(p_input[894]), .B(p_input[862]), .Z(n24177) );
  XNOR U24004 ( .A(n23276), .B(n24172), .Z(n24174) );
  XOR U24005 ( .A(n24178), .B(n24179), .Z(n23276) );
  AND U24006 ( .A(n551), .B(n24180), .Z(n24179) );
  XOR U24007 ( .A(p_input[830]), .B(p_input[798]), .Z(n24180) );
  XOR U24008 ( .A(n24181), .B(n24182), .Z(n24172) );
  AND U24009 ( .A(n24183), .B(n24184), .Z(n24182) );
  XOR U24010 ( .A(n24181), .B(n23291), .Z(n24184) );
  XNOR U24011 ( .A(p_input[861]), .B(n24185), .Z(n23291) );
  AND U24012 ( .A(n554), .B(n24186), .Z(n24185) );
  XOR U24013 ( .A(p_input[893]), .B(p_input[861]), .Z(n24186) );
  XNOR U24014 ( .A(n23288), .B(n24181), .Z(n24183) );
  XOR U24015 ( .A(n24187), .B(n24188), .Z(n23288) );
  AND U24016 ( .A(n551), .B(n24189), .Z(n24188) );
  XOR U24017 ( .A(p_input[829]), .B(p_input[797]), .Z(n24189) );
  XOR U24018 ( .A(n24190), .B(n24191), .Z(n24181) );
  AND U24019 ( .A(n24192), .B(n24193), .Z(n24191) );
  XOR U24020 ( .A(n24190), .B(n23303), .Z(n24193) );
  XNOR U24021 ( .A(p_input[860]), .B(n24194), .Z(n23303) );
  AND U24022 ( .A(n554), .B(n24195), .Z(n24194) );
  XOR U24023 ( .A(p_input[892]), .B(p_input[860]), .Z(n24195) );
  XNOR U24024 ( .A(n23300), .B(n24190), .Z(n24192) );
  XOR U24025 ( .A(n24196), .B(n24197), .Z(n23300) );
  AND U24026 ( .A(n551), .B(n24198), .Z(n24197) );
  XOR U24027 ( .A(p_input[828]), .B(p_input[796]), .Z(n24198) );
  XOR U24028 ( .A(n24199), .B(n24200), .Z(n24190) );
  AND U24029 ( .A(n24201), .B(n24202), .Z(n24200) );
  XOR U24030 ( .A(n24199), .B(n23315), .Z(n24202) );
  XNOR U24031 ( .A(p_input[859]), .B(n24203), .Z(n23315) );
  AND U24032 ( .A(n554), .B(n24204), .Z(n24203) );
  XOR U24033 ( .A(p_input[891]), .B(p_input[859]), .Z(n24204) );
  XNOR U24034 ( .A(n23312), .B(n24199), .Z(n24201) );
  XOR U24035 ( .A(n24205), .B(n24206), .Z(n23312) );
  AND U24036 ( .A(n551), .B(n24207), .Z(n24206) );
  XOR U24037 ( .A(p_input[827]), .B(p_input[795]), .Z(n24207) );
  XOR U24038 ( .A(n24208), .B(n24209), .Z(n24199) );
  AND U24039 ( .A(n24210), .B(n24211), .Z(n24209) );
  XOR U24040 ( .A(n24208), .B(n23327), .Z(n24211) );
  XNOR U24041 ( .A(p_input[858]), .B(n24212), .Z(n23327) );
  AND U24042 ( .A(n554), .B(n24213), .Z(n24212) );
  XOR U24043 ( .A(p_input[890]), .B(p_input[858]), .Z(n24213) );
  XNOR U24044 ( .A(n23324), .B(n24208), .Z(n24210) );
  XOR U24045 ( .A(n24214), .B(n24215), .Z(n23324) );
  AND U24046 ( .A(n551), .B(n24216), .Z(n24215) );
  XOR U24047 ( .A(p_input[826]), .B(p_input[794]), .Z(n24216) );
  XOR U24048 ( .A(n24217), .B(n24218), .Z(n24208) );
  AND U24049 ( .A(n24219), .B(n24220), .Z(n24218) );
  XOR U24050 ( .A(n24217), .B(n23339), .Z(n24220) );
  XNOR U24051 ( .A(p_input[857]), .B(n24221), .Z(n23339) );
  AND U24052 ( .A(n554), .B(n24222), .Z(n24221) );
  XOR U24053 ( .A(p_input[889]), .B(p_input[857]), .Z(n24222) );
  XNOR U24054 ( .A(n23336), .B(n24217), .Z(n24219) );
  XOR U24055 ( .A(n24223), .B(n24224), .Z(n23336) );
  AND U24056 ( .A(n551), .B(n24225), .Z(n24224) );
  XOR U24057 ( .A(p_input[825]), .B(p_input[793]), .Z(n24225) );
  XOR U24058 ( .A(n24226), .B(n24227), .Z(n24217) );
  AND U24059 ( .A(n24228), .B(n24229), .Z(n24227) );
  XOR U24060 ( .A(n24226), .B(n23351), .Z(n24229) );
  XNOR U24061 ( .A(p_input[856]), .B(n24230), .Z(n23351) );
  AND U24062 ( .A(n554), .B(n24231), .Z(n24230) );
  XOR U24063 ( .A(p_input[888]), .B(p_input[856]), .Z(n24231) );
  XNOR U24064 ( .A(n23348), .B(n24226), .Z(n24228) );
  XOR U24065 ( .A(n24232), .B(n24233), .Z(n23348) );
  AND U24066 ( .A(n551), .B(n24234), .Z(n24233) );
  XOR U24067 ( .A(p_input[824]), .B(p_input[792]), .Z(n24234) );
  XOR U24068 ( .A(n24235), .B(n24236), .Z(n24226) );
  AND U24069 ( .A(n24237), .B(n24238), .Z(n24236) );
  XOR U24070 ( .A(n24235), .B(n23363), .Z(n24238) );
  XNOR U24071 ( .A(p_input[855]), .B(n24239), .Z(n23363) );
  AND U24072 ( .A(n554), .B(n24240), .Z(n24239) );
  XOR U24073 ( .A(p_input[887]), .B(p_input[855]), .Z(n24240) );
  XNOR U24074 ( .A(n23360), .B(n24235), .Z(n24237) );
  XOR U24075 ( .A(n24241), .B(n24242), .Z(n23360) );
  AND U24076 ( .A(n551), .B(n24243), .Z(n24242) );
  XOR U24077 ( .A(p_input[823]), .B(p_input[791]), .Z(n24243) );
  XOR U24078 ( .A(n24244), .B(n24245), .Z(n24235) );
  AND U24079 ( .A(n24246), .B(n24247), .Z(n24245) );
  XOR U24080 ( .A(n24244), .B(n23375), .Z(n24247) );
  XNOR U24081 ( .A(p_input[854]), .B(n24248), .Z(n23375) );
  AND U24082 ( .A(n554), .B(n24249), .Z(n24248) );
  XOR U24083 ( .A(p_input[886]), .B(p_input[854]), .Z(n24249) );
  XNOR U24084 ( .A(n23372), .B(n24244), .Z(n24246) );
  XOR U24085 ( .A(n24250), .B(n24251), .Z(n23372) );
  AND U24086 ( .A(n551), .B(n24252), .Z(n24251) );
  XOR U24087 ( .A(p_input[822]), .B(p_input[790]), .Z(n24252) );
  XOR U24088 ( .A(n24253), .B(n24254), .Z(n24244) );
  AND U24089 ( .A(n24255), .B(n24256), .Z(n24254) );
  XOR U24090 ( .A(n24253), .B(n23387), .Z(n24256) );
  XNOR U24091 ( .A(p_input[853]), .B(n24257), .Z(n23387) );
  AND U24092 ( .A(n554), .B(n24258), .Z(n24257) );
  XOR U24093 ( .A(p_input[885]), .B(p_input[853]), .Z(n24258) );
  XNOR U24094 ( .A(n23384), .B(n24253), .Z(n24255) );
  XOR U24095 ( .A(n24259), .B(n24260), .Z(n23384) );
  AND U24096 ( .A(n551), .B(n24261), .Z(n24260) );
  XOR U24097 ( .A(p_input[821]), .B(p_input[789]), .Z(n24261) );
  XOR U24098 ( .A(n24262), .B(n24263), .Z(n24253) );
  AND U24099 ( .A(n24264), .B(n24265), .Z(n24263) );
  XOR U24100 ( .A(n24262), .B(n23399), .Z(n24265) );
  XNOR U24101 ( .A(p_input[852]), .B(n24266), .Z(n23399) );
  AND U24102 ( .A(n554), .B(n24267), .Z(n24266) );
  XOR U24103 ( .A(p_input[884]), .B(p_input[852]), .Z(n24267) );
  XNOR U24104 ( .A(n23396), .B(n24262), .Z(n24264) );
  XOR U24105 ( .A(n24268), .B(n24269), .Z(n23396) );
  AND U24106 ( .A(n551), .B(n24270), .Z(n24269) );
  XOR U24107 ( .A(p_input[820]), .B(p_input[788]), .Z(n24270) );
  XOR U24108 ( .A(n24271), .B(n24272), .Z(n24262) );
  AND U24109 ( .A(n24273), .B(n24274), .Z(n24272) );
  XOR U24110 ( .A(n24271), .B(n23411), .Z(n24274) );
  XNOR U24111 ( .A(p_input[851]), .B(n24275), .Z(n23411) );
  AND U24112 ( .A(n554), .B(n24276), .Z(n24275) );
  XOR U24113 ( .A(p_input[883]), .B(p_input[851]), .Z(n24276) );
  XNOR U24114 ( .A(n23408), .B(n24271), .Z(n24273) );
  XOR U24115 ( .A(n24277), .B(n24278), .Z(n23408) );
  AND U24116 ( .A(n551), .B(n24279), .Z(n24278) );
  XOR U24117 ( .A(p_input[819]), .B(p_input[787]), .Z(n24279) );
  XOR U24118 ( .A(n24280), .B(n24281), .Z(n24271) );
  AND U24119 ( .A(n24282), .B(n24283), .Z(n24281) );
  XOR U24120 ( .A(n24280), .B(n23423), .Z(n24283) );
  XNOR U24121 ( .A(p_input[850]), .B(n24284), .Z(n23423) );
  AND U24122 ( .A(n554), .B(n24285), .Z(n24284) );
  XOR U24123 ( .A(p_input[882]), .B(p_input[850]), .Z(n24285) );
  XNOR U24124 ( .A(n23420), .B(n24280), .Z(n24282) );
  XOR U24125 ( .A(n24286), .B(n24287), .Z(n23420) );
  AND U24126 ( .A(n551), .B(n24288), .Z(n24287) );
  XOR U24127 ( .A(p_input[818]), .B(p_input[786]), .Z(n24288) );
  XOR U24128 ( .A(n24289), .B(n24290), .Z(n24280) );
  AND U24129 ( .A(n24291), .B(n24292), .Z(n24290) );
  XOR U24130 ( .A(n24289), .B(n23435), .Z(n24292) );
  XNOR U24131 ( .A(p_input[849]), .B(n24293), .Z(n23435) );
  AND U24132 ( .A(n554), .B(n24294), .Z(n24293) );
  XOR U24133 ( .A(p_input[881]), .B(p_input[849]), .Z(n24294) );
  XNOR U24134 ( .A(n23432), .B(n24289), .Z(n24291) );
  XOR U24135 ( .A(n24295), .B(n24296), .Z(n23432) );
  AND U24136 ( .A(n551), .B(n24297), .Z(n24296) );
  XOR U24137 ( .A(p_input[817]), .B(p_input[785]), .Z(n24297) );
  XOR U24138 ( .A(n24298), .B(n24299), .Z(n24289) );
  AND U24139 ( .A(n24300), .B(n24301), .Z(n24299) );
  XOR U24140 ( .A(n24298), .B(n23447), .Z(n24301) );
  XNOR U24141 ( .A(p_input[848]), .B(n24302), .Z(n23447) );
  AND U24142 ( .A(n554), .B(n24303), .Z(n24302) );
  XOR U24143 ( .A(p_input[880]), .B(p_input[848]), .Z(n24303) );
  XNOR U24144 ( .A(n23444), .B(n24298), .Z(n24300) );
  XOR U24145 ( .A(n24304), .B(n24305), .Z(n23444) );
  AND U24146 ( .A(n551), .B(n24306), .Z(n24305) );
  XOR U24147 ( .A(p_input[816]), .B(p_input[784]), .Z(n24306) );
  XOR U24148 ( .A(n24307), .B(n24308), .Z(n24298) );
  AND U24149 ( .A(n24309), .B(n24310), .Z(n24308) );
  XOR U24150 ( .A(n24307), .B(n23459), .Z(n24310) );
  XNOR U24151 ( .A(p_input[847]), .B(n24311), .Z(n23459) );
  AND U24152 ( .A(n554), .B(n24312), .Z(n24311) );
  XOR U24153 ( .A(p_input[879]), .B(p_input[847]), .Z(n24312) );
  XNOR U24154 ( .A(n23456), .B(n24307), .Z(n24309) );
  XOR U24155 ( .A(n24313), .B(n24314), .Z(n23456) );
  AND U24156 ( .A(n551), .B(n24315), .Z(n24314) );
  XOR U24157 ( .A(p_input[815]), .B(p_input[783]), .Z(n24315) );
  XOR U24158 ( .A(n24316), .B(n24317), .Z(n24307) );
  AND U24159 ( .A(n24318), .B(n24319), .Z(n24317) );
  XOR U24160 ( .A(n24316), .B(n23471), .Z(n24319) );
  XNOR U24161 ( .A(p_input[846]), .B(n24320), .Z(n23471) );
  AND U24162 ( .A(n554), .B(n24321), .Z(n24320) );
  XOR U24163 ( .A(p_input[878]), .B(p_input[846]), .Z(n24321) );
  XNOR U24164 ( .A(n23468), .B(n24316), .Z(n24318) );
  XOR U24165 ( .A(n24322), .B(n24323), .Z(n23468) );
  AND U24166 ( .A(n551), .B(n24324), .Z(n24323) );
  XOR U24167 ( .A(p_input[814]), .B(p_input[782]), .Z(n24324) );
  XOR U24168 ( .A(n24325), .B(n24326), .Z(n24316) );
  AND U24169 ( .A(n24327), .B(n24328), .Z(n24326) );
  XOR U24170 ( .A(n24325), .B(n23483), .Z(n24328) );
  XNOR U24171 ( .A(p_input[845]), .B(n24329), .Z(n23483) );
  AND U24172 ( .A(n554), .B(n24330), .Z(n24329) );
  XOR U24173 ( .A(p_input[877]), .B(p_input[845]), .Z(n24330) );
  XNOR U24174 ( .A(n23480), .B(n24325), .Z(n24327) );
  XOR U24175 ( .A(n24331), .B(n24332), .Z(n23480) );
  AND U24176 ( .A(n551), .B(n24333), .Z(n24332) );
  XOR U24177 ( .A(p_input[813]), .B(p_input[781]), .Z(n24333) );
  XOR U24178 ( .A(n24334), .B(n24335), .Z(n24325) );
  AND U24179 ( .A(n24336), .B(n24337), .Z(n24335) );
  XOR U24180 ( .A(n24334), .B(n23495), .Z(n24337) );
  XNOR U24181 ( .A(p_input[844]), .B(n24338), .Z(n23495) );
  AND U24182 ( .A(n554), .B(n24339), .Z(n24338) );
  XOR U24183 ( .A(p_input[876]), .B(p_input[844]), .Z(n24339) );
  XNOR U24184 ( .A(n23492), .B(n24334), .Z(n24336) );
  XOR U24185 ( .A(n24340), .B(n24341), .Z(n23492) );
  AND U24186 ( .A(n551), .B(n24342), .Z(n24341) );
  XOR U24187 ( .A(p_input[812]), .B(p_input[780]), .Z(n24342) );
  XOR U24188 ( .A(n24343), .B(n24344), .Z(n24334) );
  AND U24189 ( .A(n24345), .B(n24346), .Z(n24344) );
  XOR U24190 ( .A(n24343), .B(n23507), .Z(n24346) );
  XNOR U24191 ( .A(p_input[843]), .B(n24347), .Z(n23507) );
  AND U24192 ( .A(n554), .B(n24348), .Z(n24347) );
  XOR U24193 ( .A(p_input[875]), .B(p_input[843]), .Z(n24348) );
  XNOR U24194 ( .A(n23504), .B(n24343), .Z(n24345) );
  XOR U24195 ( .A(n24349), .B(n24350), .Z(n23504) );
  AND U24196 ( .A(n551), .B(n24351), .Z(n24350) );
  XOR U24197 ( .A(p_input[811]), .B(p_input[779]), .Z(n24351) );
  XOR U24198 ( .A(n24352), .B(n24353), .Z(n24343) );
  AND U24199 ( .A(n24354), .B(n24355), .Z(n24353) );
  XOR U24200 ( .A(n24352), .B(n23519), .Z(n24355) );
  XNOR U24201 ( .A(p_input[842]), .B(n24356), .Z(n23519) );
  AND U24202 ( .A(n554), .B(n24357), .Z(n24356) );
  XOR U24203 ( .A(p_input[874]), .B(p_input[842]), .Z(n24357) );
  XNOR U24204 ( .A(n23516), .B(n24352), .Z(n24354) );
  XOR U24205 ( .A(n24358), .B(n24359), .Z(n23516) );
  AND U24206 ( .A(n551), .B(n24360), .Z(n24359) );
  XOR U24207 ( .A(p_input[810]), .B(p_input[778]), .Z(n24360) );
  XOR U24208 ( .A(n24361), .B(n24362), .Z(n24352) );
  AND U24209 ( .A(n24363), .B(n24364), .Z(n24362) );
  XOR U24210 ( .A(n24361), .B(n23531), .Z(n24364) );
  XNOR U24211 ( .A(p_input[841]), .B(n24365), .Z(n23531) );
  AND U24212 ( .A(n554), .B(n24366), .Z(n24365) );
  XOR U24213 ( .A(p_input[873]), .B(p_input[841]), .Z(n24366) );
  XNOR U24214 ( .A(n23528), .B(n24361), .Z(n24363) );
  XOR U24215 ( .A(n24367), .B(n24368), .Z(n23528) );
  AND U24216 ( .A(n551), .B(n24369), .Z(n24368) );
  XOR U24217 ( .A(p_input[809]), .B(p_input[777]), .Z(n24369) );
  XOR U24218 ( .A(n24370), .B(n24371), .Z(n24361) );
  AND U24219 ( .A(n24372), .B(n24373), .Z(n24371) );
  XOR U24220 ( .A(n24370), .B(n23543), .Z(n24373) );
  XNOR U24221 ( .A(p_input[840]), .B(n24374), .Z(n23543) );
  AND U24222 ( .A(n554), .B(n24375), .Z(n24374) );
  XOR U24223 ( .A(p_input[872]), .B(p_input[840]), .Z(n24375) );
  XNOR U24224 ( .A(n23540), .B(n24370), .Z(n24372) );
  XOR U24225 ( .A(n24376), .B(n24377), .Z(n23540) );
  AND U24226 ( .A(n551), .B(n24378), .Z(n24377) );
  XOR U24227 ( .A(p_input[808]), .B(p_input[776]), .Z(n24378) );
  XOR U24228 ( .A(n24379), .B(n24380), .Z(n24370) );
  AND U24229 ( .A(n24381), .B(n24382), .Z(n24380) );
  XOR U24230 ( .A(n24379), .B(n23555), .Z(n24382) );
  XNOR U24231 ( .A(p_input[839]), .B(n24383), .Z(n23555) );
  AND U24232 ( .A(n554), .B(n24384), .Z(n24383) );
  XOR U24233 ( .A(p_input[871]), .B(p_input[839]), .Z(n24384) );
  XNOR U24234 ( .A(n23552), .B(n24379), .Z(n24381) );
  XOR U24235 ( .A(n24385), .B(n24386), .Z(n23552) );
  AND U24236 ( .A(n551), .B(n24387), .Z(n24386) );
  XOR U24237 ( .A(p_input[807]), .B(p_input[775]), .Z(n24387) );
  XOR U24238 ( .A(n24388), .B(n24389), .Z(n24379) );
  AND U24239 ( .A(n24390), .B(n24391), .Z(n24389) );
  XOR U24240 ( .A(n24388), .B(n23567), .Z(n24391) );
  XNOR U24241 ( .A(p_input[838]), .B(n24392), .Z(n23567) );
  AND U24242 ( .A(n554), .B(n24393), .Z(n24392) );
  XOR U24243 ( .A(p_input[870]), .B(p_input[838]), .Z(n24393) );
  XNOR U24244 ( .A(n23564), .B(n24388), .Z(n24390) );
  XOR U24245 ( .A(n24394), .B(n24395), .Z(n23564) );
  AND U24246 ( .A(n551), .B(n24396), .Z(n24395) );
  XOR U24247 ( .A(p_input[806]), .B(p_input[774]), .Z(n24396) );
  XOR U24248 ( .A(n24397), .B(n24398), .Z(n24388) );
  AND U24249 ( .A(n24399), .B(n24400), .Z(n24398) );
  XOR U24250 ( .A(n24397), .B(n23579), .Z(n24400) );
  XNOR U24251 ( .A(p_input[837]), .B(n24401), .Z(n23579) );
  AND U24252 ( .A(n554), .B(n24402), .Z(n24401) );
  XOR U24253 ( .A(p_input[869]), .B(p_input[837]), .Z(n24402) );
  XNOR U24254 ( .A(n23576), .B(n24397), .Z(n24399) );
  XOR U24255 ( .A(n24403), .B(n24404), .Z(n23576) );
  AND U24256 ( .A(n551), .B(n24405), .Z(n24404) );
  XOR U24257 ( .A(p_input[805]), .B(p_input[773]), .Z(n24405) );
  XOR U24258 ( .A(n24406), .B(n24407), .Z(n24397) );
  AND U24259 ( .A(n24408), .B(n24409), .Z(n24407) );
  XOR U24260 ( .A(n24406), .B(n23591), .Z(n24409) );
  XNOR U24261 ( .A(p_input[836]), .B(n24410), .Z(n23591) );
  AND U24262 ( .A(n554), .B(n24411), .Z(n24410) );
  XOR U24263 ( .A(p_input[868]), .B(p_input[836]), .Z(n24411) );
  XNOR U24264 ( .A(n23588), .B(n24406), .Z(n24408) );
  XOR U24265 ( .A(n24412), .B(n24413), .Z(n23588) );
  AND U24266 ( .A(n551), .B(n24414), .Z(n24413) );
  XOR U24267 ( .A(p_input[804]), .B(p_input[772]), .Z(n24414) );
  XOR U24268 ( .A(n24415), .B(n24416), .Z(n24406) );
  AND U24269 ( .A(n24417), .B(n24418), .Z(n24416) );
  XOR U24270 ( .A(n24415), .B(n23603), .Z(n24418) );
  XNOR U24271 ( .A(p_input[835]), .B(n24419), .Z(n23603) );
  AND U24272 ( .A(n554), .B(n24420), .Z(n24419) );
  XOR U24273 ( .A(p_input[867]), .B(p_input[835]), .Z(n24420) );
  XNOR U24274 ( .A(n23600), .B(n24415), .Z(n24417) );
  XOR U24275 ( .A(n24421), .B(n24422), .Z(n23600) );
  AND U24276 ( .A(n551), .B(n24423), .Z(n24422) );
  XOR U24277 ( .A(p_input[803]), .B(p_input[771]), .Z(n24423) );
  XOR U24278 ( .A(n24424), .B(n24425), .Z(n24415) );
  AND U24279 ( .A(n24426), .B(n24427), .Z(n24425) );
  XOR U24280 ( .A(n23615), .B(n24424), .Z(n24427) );
  XNOR U24281 ( .A(p_input[834]), .B(n24428), .Z(n23615) );
  AND U24282 ( .A(n554), .B(n24429), .Z(n24428) );
  XOR U24283 ( .A(p_input[866]), .B(p_input[834]), .Z(n24429) );
  XNOR U24284 ( .A(n24424), .B(n23612), .Z(n24426) );
  XOR U24285 ( .A(n24430), .B(n24431), .Z(n23612) );
  AND U24286 ( .A(n551), .B(n24432), .Z(n24431) );
  XOR U24287 ( .A(p_input[802]), .B(p_input[770]), .Z(n24432) );
  XOR U24288 ( .A(n24433), .B(n24434), .Z(n24424) );
  AND U24289 ( .A(n24435), .B(n24436), .Z(n24434) );
  XNOR U24290 ( .A(n24437), .B(n23628), .Z(n24436) );
  XNOR U24291 ( .A(p_input[833]), .B(n24438), .Z(n23628) );
  AND U24292 ( .A(n554), .B(n24439), .Z(n24438) );
  XNOR U24293 ( .A(p_input[865]), .B(n24440), .Z(n24439) );
  IV U24294 ( .A(p_input[833]), .Z(n24440) );
  XNOR U24295 ( .A(n23625), .B(n24433), .Z(n24435) );
  XNOR U24296 ( .A(p_input[769]), .B(n24441), .Z(n23625) );
  AND U24297 ( .A(n551), .B(n24442), .Z(n24441) );
  XOR U24298 ( .A(p_input[801]), .B(p_input[769]), .Z(n24442) );
  IV U24299 ( .A(n24437), .Z(n24433) );
  AND U24300 ( .A(n24163), .B(n24166), .Z(n24437) );
  XOR U24301 ( .A(p_input[832]), .B(n24443), .Z(n24166) );
  AND U24302 ( .A(n554), .B(n24444), .Z(n24443) );
  XOR U24303 ( .A(p_input[864]), .B(p_input[832]), .Z(n24444) );
  XOR U24304 ( .A(n24445), .B(n24446), .Z(n554) );
  AND U24305 ( .A(n24447), .B(n24448), .Z(n24446) );
  XNOR U24306 ( .A(p_input[895]), .B(n24445), .Z(n24448) );
  XOR U24307 ( .A(n24445), .B(p_input[863]), .Z(n24447) );
  XOR U24308 ( .A(n24449), .B(n24450), .Z(n24445) );
  AND U24309 ( .A(n24451), .B(n24452), .Z(n24450) );
  XNOR U24310 ( .A(p_input[894]), .B(n24449), .Z(n24452) );
  XOR U24311 ( .A(n24449), .B(p_input[862]), .Z(n24451) );
  XOR U24312 ( .A(n24453), .B(n24454), .Z(n24449) );
  AND U24313 ( .A(n24455), .B(n24456), .Z(n24454) );
  XNOR U24314 ( .A(p_input[893]), .B(n24453), .Z(n24456) );
  XOR U24315 ( .A(n24453), .B(p_input[861]), .Z(n24455) );
  XOR U24316 ( .A(n24457), .B(n24458), .Z(n24453) );
  AND U24317 ( .A(n24459), .B(n24460), .Z(n24458) );
  XNOR U24318 ( .A(p_input[892]), .B(n24457), .Z(n24460) );
  XOR U24319 ( .A(n24457), .B(p_input[860]), .Z(n24459) );
  XOR U24320 ( .A(n24461), .B(n24462), .Z(n24457) );
  AND U24321 ( .A(n24463), .B(n24464), .Z(n24462) );
  XNOR U24322 ( .A(p_input[891]), .B(n24461), .Z(n24464) );
  XOR U24323 ( .A(n24461), .B(p_input[859]), .Z(n24463) );
  XOR U24324 ( .A(n24465), .B(n24466), .Z(n24461) );
  AND U24325 ( .A(n24467), .B(n24468), .Z(n24466) );
  XNOR U24326 ( .A(p_input[890]), .B(n24465), .Z(n24468) );
  XOR U24327 ( .A(n24465), .B(p_input[858]), .Z(n24467) );
  XOR U24328 ( .A(n24469), .B(n24470), .Z(n24465) );
  AND U24329 ( .A(n24471), .B(n24472), .Z(n24470) );
  XNOR U24330 ( .A(p_input[889]), .B(n24469), .Z(n24472) );
  XOR U24331 ( .A(n24469), .B(p_input[857]), .Z(n24471) );
  XOR U24332 ( .A(n24473), .B(n24474), .Z(n24469) );
  AND U24333 ( .A(n24475), .B(n24476), .Z(n24474) );
  XNOR U24334 ( .A(p_input[888]), .B(n24473), .Z(n24476) );
  XOR U24335 ( .A(n24473), .B(p_input[856]), .Z(n24475) );
  XOR U24336 ( .A(n24477), .B(n24478), .Z(n24473) );
  AND U24337 ( .A(n24479), .B(n24480), .Z(n24478) );
  XNOR U24338 ( .A(p_input[887]), .B(n24477), .Z(n24480) );
  XOR U24339 ( .A(n24477), .B(p_input[855]), .Z(n24479) );
  XOR U24340 ( .A(n24481), .B(n24482), .Z(n24477) );
  AND U24341 ( .A(n24483), .B(n24484), .Z(n24482) );
  XNOR U24342 ( .A(p_input[886]), .B(n24481), .Z(n24484) );
  XOR U24343 ( .A(n24481), .B(p_input[854]), .Z(n24483) );
  XOR U24344 ( .A(n24485), .B(n24486), .Z(n24481) );
  AND U24345 ( .A(n24487), .B(n24488), .Z(n24486) );
  XNOR U24346 ( .A(p_input[885]), .B(n24485), .Z(n24488) );
  XOR U24347 ( .A(n24485), .B(p_input[853]), .Z(n24487) );
  XOR U24348 ( .A(n24489), .B(n24490), .Z(n24485) );
  AND U24349 ( .A(n24491), .B(n24492), .Z(n24490) );
  XNOR U24350 ( .A(p_input[884]), .B(n24489), .Z(n24492) );
  XOR U24351 ( .A(n24489), .B(p_input[852]), .Z(n24491) );
  XOR U24352 ( .A(n24493), .B(n24494), .Z(n24489) );
  AND U24353 ( .A(n24495), .B(n24496), .Z(n24494) );
  XNOR U24354 ( .A(p_input[883]), .B(n24493), .Z(n24496) );
  XOR U24355 ( .A(n24493), .B(p_input[851]), .Z(n24495) );
  XOR U24356 ( .A(n24497), .B(n24498), .Z(n24493) );
  AND U24357 ( .A(n24499), .B(n24500), .Z(n24498) );
  XNOR U24358 ( .A(p_input[882]), .B(n24497), .Z(n24500) );
  XOR U24359 ( .A(n24497), .B(p_input[850]), .Z(n24499) );
  XOR U24360 ( .A(n24501), .B(n24502), .Z(n24497) );
  AND U24361 ( .A(n24503), .B(n24504), .Z(n24502) );
  XNOR U24362 ( .A(p_input[881]), .B(n24501), .Z(n24504) );
  XOR U24363 ( .A(n24501), .B(p_input[849]), .Z(n24503) );
  XOR U24364 ( .A(n24505), .B(n24506), .Z(n24501) );
  AND U24365 ( .A(n24507), .B(n24508), .Z(n24506) );
  XNOR U24366 ( .A(p_input[880]), .B(n24505), .Z(n24508) );
  XOR U24367 ( .A(n24505), .B(p_input[848]), .Z(n24507) );
  XOR U24368 ( .A(n24509), .B(n24510), .Z(n24505) );
  AND U24369 ( .A(n24511), .B(n24512), .Z(n24510) );
  XNOR U24370 ( .A(p_input[879]), .B(n24509), .Z(n24512) );
  XOR U24371 ( .A(n24509), .B(p_input[847]), .Z(n24511) );
  XOR U24372 ( .A(n24513), .B(n24514), .Z(n24509) );
  AND U24373 ( .A(n24515), .B(n24516), .Z(n24514) );
  XNOR U24374 ( .A(p_input[878]), .B(n24513), .Z(n24516) );
  XOR U24375 ( .A(n24513), .B(p_input[846]), .Z(n24515) );
  XOR U24376 ( .A(n24517), .B(n24518), .Z(n24513) );
  AND U24377 ( .A(n24519), .B(n24520), .Z(n24518) );
  XNOR U24378 ( .A(p_input[877]), .B(n24517), .Z(n24520) );
  XOR U24379 ( .A(n24517), .B(p_input[845]), .Z(n24519) );
  XOR U24380 ( .A(n24521), .B(n24522), .Z(n24517) );
  AND U24381 ( .A(n24523), .B(n24524), .Z(n24522) );
  XNOR U24382 ( .A(p_input[876]), .B(n24521), .Z(n24524) );
  XOR U24383 ( .A(n24521), .B(p_input[844]), .Z(n24523) );
  XOR U24384 ( .A(n24525), .B(n24526), .Z(n24521) );
  AND U24385 ( .A(n24527), .B(n24528), .Z(n24526) );
  XNOR U24386 ( .A(p_input[875]), .B(n24525), .Z(n24528) );
  XOR U24387 ( .A(n24525), .B(p_input[843]), .Z(n24527) );
  XOR U24388 ( .A(n24529), .B(n24530), .Z(n24525) );
  AND U24389 ( .A(n24531), .B(n24532), .Z(n24530) );
  XNOR U24390 ( .A(p_input[874]), .B(n24529), .Z(n24532) );
  XOR U24391 ( .A(n24529), .B(p_input[842]), .Z(n24531) );
  XOR U24392 ( .A(n24533), .B(n24534), .Z(n24529) );
  AND U24393 ( .A(n24535), .B(n24536), .Z(n24534) );
  XNOR U24394 ( .A(p_input[873]), .B(n24533), .Z(n24536) );
  XOR U24395 ( .A(n24533), .B(p_input[841]), .Z(n24535) );
  XOR U24396 ( .A(n24537), .B(n24538), .Z(n24533) );
  AND U24397 ( .A(n24539), .B(n24540), .Z(n24538) );
  XNOR U24398 ( .A(p_input[872]), .B(n24537), .Z(n24540) );
  XOR U24399 ( .A(n24537), .B(p_input[840]), .Z(n24539) );
  XOR U24400 ( .A(n24541), .B(n24542), .Z(n24537) );
  AND U24401 ( .A(n24543), .B(n24544), .Z(n24542) );
  XNOR U24402 ( .A(p_input[871]), .B(n24541), .Z(n24544) );
  XOR U24403 ( .A(n24541), .B(p_input[839]), .Z(n24543) );
  XOR U24404 ( .A(n24545), .B(n24546), .Z(n24541) );
  AND U24405 ( .A(n24547), .B(n24548), .Z(n24546) );
  XNOR U24406 ( .A(p_input[870]), .B(n24545), .Z(n24548) );
  XOR U24407 ( .A(n24545), .B(p_input[838]), .Z(n24547) );
  XOR U24408 ( .A(n24549), .B(n24550), .Z(n24545) );
  AND U24409 ( .A(n24551), .B(n24552), .Z(n24550) );
  XNOR U24410 ( .A(p_input[869]), .B(n24549), .Z(n24552) );
  XOR U24411 ( .A(n24549), .B(p_input[837]), .Z(n24551) );
  XOR U24412 ( .A(n24553), .B(n24554), .Z(n24549) );
  AND U24413 ( .A(n24555), .B(n24556), .Z(n24554) );
  XNOR U24414 ( .A(p_input[868]), .B(n24553), .Z(n24556) );
  XOR U24415 ( .A(n24553), .B(p_input[836]), .Z(n24555) );
  XOR U24416 ( .A(n24557), .B(n24558), .Z(n24553) );
  AND U24417 ( .A(n24559), .B(n24560), .Z(n24558) );
  XNOR U24418 ( .A(p_input[867]), .B(n24557), .Z(n24560) );
  XOR U24419 ( .A(n24557), .B(p_input[835]), .Z(n24559) );
  XOR U24420 ( .A(n24561), .B(n24562), .Z(n24557) );
  AND U24421 ( .A(n24563), .B(n24564), .Z(n24562) );
  XNOR U24422 ( .A(p_input[866]), .B(n24561), .Z(n24564) );
  XOR U24423 ( .A(n24561), .B(p_input[834]), .Z(n24563) );
  XNOR U24424 ( .A(n24565), .B(n24566), .Z(n24561) );
  AND U24425 ( .A(n24567), .B(n24568), .Z(n24566) );
  XOR U24426 ( .A(p_input[865]), .B(n24565), .Z(n24568) );
  XNOR U24427 ( .A(p_input[833]), .B(n24565), .Z(n24567) );
  AND U24428 ( .A(p_input[864]), .B(n24569), .Z(n24565) );
  IV U24429 ( .A(p_input[832]), .Z(n24569) );
  XNOR U24430 ( .A(p_input[768]), .B(n24570), .Z(n24163) );
  AND U24431 ( .A(n551), .B(n24571), .Z(n24570) );
  XOR U24432 ( .A(p_input[800]), .B(p_input[768]), .Z(n24571) );
  XOR U24433 ( .A(n24572), .B(n24573), .Z(n551) );
  AND U24434 ( .A(n24574), .B(n24575), .Z(n24573) );
  XNOR U24435 ( .A(p_input[831]), .B(n24572), .Z(n24575) );
  XOR U24436 ( .A(n24572), .B(p_input[799]), .Z(n24574) );
  XOR U24437 ( .A(n24576), .B(n24577), .Z(n24572) );
  AND U24438 ( .A(n24578), .B(n24579), .Z(n24577) );
  XNOR U24439 ( .A(p_input[830]), .B(n24576), .Z(n24579) );
  XNOR U24440 ( .A(n24576), .B(n24178), .Z(n24578) );
  IV U24441 ( .A(p_input[798]), .Z(n24178) );
  XOR U24442 ( .A(n24580), .B(n24581), .Z(n24576) );
  AND U24443 ( .A(n24582), .B(n24583), .Z(n24581) );
  XNOR U24444 ( .A(p_input[829]), .B(n24580), .Z(n24583) );
  XNOR U24445 ( .A(n24580), .B(n24187), .Z(n24582) );
  IV U24446 ( .A(p_input[797]), .Z(n24187) );
  XOR U24447 ( .A(n24584), .B(n24585), .Z(n24580) );
  AND U24448 ( .A(n24586), .B(n24587), .Z(n24585) );
  XNOR U24449 ( .A(p_input[828]), .B(n24584), .Z(n24587) );
  XNOR U24450 ( .A(n24584), .B(n24196), .Z(n24586) );
  IV U24451 ( .A(p_input[796]), .Z(n24196) );
  XOR U24452 ( .A(n24588), .B(n24589), .Z(n24584) );
  AND U24453 ( .A(n24590), .B(n24591), .Z(n24589) );
  XNOR U24454 ( .A(p_input[827]), .B(n24588), .Z(n24591) );
  XNOR U24455 ( .A(n24588), .B(n24205), .Z(n24590) );
  IV U24456 ( .A(p_input[795]), .Z(n24205) );
  XOR U24457 ( .A(n24592), .B(n24593), .Z(n24588) );
  AND U24458 ( .A(n24594), .B(n24595), .Z(n24593) );
  XNOR U24459 ( .A(p_input[826]), .B(n24592), .Z(n24595) );
  XNOR U24460 ( .A(n24592), .B(n24214), .Z(n24594) );
  IV U24461 ( .A(p_input[794]), .Z(n24214) );
  XOR U24462 ( .A(n24596), .B(n24597), .Z(n24592) );
  AND U24463 ( .A(n24598), .B(n24599), .Z(n24597) );
  XNOR U24464 ( .A(p_input[825]), .B(n24596), .Z(n24599) );
  XNOR U24465 ( .A(n24596), .B(n24223), .Z(n24598) );
  IV U24466 ( .A(p_input[793]), .Z(n24223) );
  XOR U24467 ( .A(n24600), .B(n24601), .Z(n24596) );
  AND U24468 ( .A(n24602), .B(n24603), .Z(n24601) );
  XNOR U24469 ( .A(p_input[824]), .B(n24600), .Z(n24603) );
  XNOR U24470 ( .A(n24600), .B(n24232), .Z(n24602) );
  IV U24471 ( .A(p_input[792]), .Z(n24232) );
  XOR U24472 ( .A(n24604), .B(n24605), .Z(n24600) );
  AND U24473 ( .A(n24606), .B(n24607), .Z(n24605) );
  XNOR U24474 ( .A(p_input[823]), .B(n24604), .Z(n24607) );
  XNOR U24475 ( .A(n24604), .B(n24241), .Z(n24606) );
  IV U24476 ( .A(p_input[791]), .Z(n24241) );
  XOR U24477 ( .A(n24608), .B(n24609), .Z(n24604) );
  AND U24478 ( .A(n24610), .B(n24611), .Z(n24609) );
  XNOR U24479 ( .A(p_input[822]), .B(n24608), .Z(n24611) );
  XNOR U24480 ( .A(n24608), .B(n24250), .Z(n24610) );
  IV U24481 ( .A(p_input[790]), .Z(n24250) );
  XOR U24482 ( .A(n24612), .B(n24613), .Z(n24608) );
  AND U24483 ( .A(n24614), .B(n24615), .Z(n24613) );
  XNOR U24484 ( .A(p_input[821]), .B(n24612), .Z(n24615) );
  XNOR U24485 ( .A(n24612), .B(n24259), .Z(n24614) );
  IV U24486 ( .A(p_input[789]), .Z(n24259) );
  XOR U24487 ( .A(n24616), .B(n24617), .Z(n24612) );
  AND U24488 ( .A(n24618), .B(n24619), .Z(n24617) );
  XNOR U24489 ( .A(p_input[820]), .B(n24616), .Z(n24619) );
  XNOR U24490 ( .A(n24616), .B(n24268), .Z(n24618) );
  IV U24491 ( .A(p_input[788]), .Z(n24268) );
  XOR U24492 ( .A(n24620), .B(n24621), .Z(n24616) );
  AND U24493 ( .A(n24622), .B(n24623), .Z(n24621) );
  XNOR U24494 ( .A(p_input[819]), .B(n24620), .Z(n24623) );
  XNOR U24495 ( .A(n24620), .B(n24277), .Z(n24622) );
  IV U24496 ( .A(p_input[787]), .Z(n24277) );
  XOR U24497 ( .A(n24624), .B(n24625), .Z(n24620) );
  AND U24498 ( .A(n24626), .B(n24627), .Z(n24625) );
  XNOR U24499 ( .A(p_input[818]), .B(n24624), .Z(n24627) );
  XNOR U24500 ( .A(n24624), .B(n24286), .Z(n24626) );
  IV U24501 ( .A(p_input[786]), .Z(n24286) );
  XOR U24502 ( .A(n24628), .B(n24629), .Z(n24624) );
  AND U24503 ( .A(n24630), .B(n24631), .Z(n24629) );
  XNOR U24504 ( .A(p_input[817]), .B(n24628), .Z(n24631) );
  XNOR U24505 ( .A(n24628), .B(n24295), .Z(n24630) );
  IV U24506 ( .A(p_input[785]), .Z(n24295) );
  XOR U24507 ( .A(n24632), .B(n24633), .Z(n24628) );
  AND U24508 ( .A(n24634), .B(n24635), .Z(n24633) );
  XNOR U24509 ( .A(p_input[816]), .B(n24632), .Z(n24635) );
  XNOR U24510 ( .A(n24632), .B(n24304), .Z(n24634) );
  IV U24511 ( .A(p_input[784]), .Z(n24304) );
  XOR U24512 ( .A(n24636), .B(n24637), .Z(n24632) );
  AND U24513 ( .A(n24638), .B(n24639), .Z(n24637) );
  XNOR U24514 ( .A(p_input[815]), .B(n24636), .Z(n24639) );
  XNOR U24515 ( .A(n24636), .B(n24313), .Z(n24638) );
  IV U24516 ( .A(p_input[783]), .Z(n24313) );
  XOR U24517 ( .A(n24640), .B(n24641), .Z(n24636) );
  AND U24518 ( .A(n24642), .B(n24643), .Z(n24641) );
  XNOR U24519 ( .A(p_input[814]), .B(n24640), .Z(n24643) );
  XNOR U24520 ( .A(n24640), .B(n24322), .Z(n24642) );
  IV U24521 ( .A(p_input[782]), .Z(n24322) );
  XOR U24522 ( .A(n24644), .B(n24645), .Z(n24640) );
  AND U24523 ( .A(n24646), .B(n24647), .Z(n24645) );
  XNOR U24524 ( .A(p_input[813]), .B(n24644), .Z(n24647) );
  XNOR U24525 ( .A(n24644), .B(n24331), .Z(n24646) );
  IV U24526 ( .A(p_input[781]), .Z(n24331) );
  XOR U24527 ( .A(n24648), .B(n24649), .Z(n24644) );
  AND U24528 ( .A(n24650), .B(n24651), .Z(n24649) );
  XNOR U24529 ( .A(p_input[812]), .B(n24648), .Z(n24651) );
  XNOR U24530 ( .A(n24648), .B(n24340), .Z(n24650) );
  IV U24531 ( .A(p_input[780]), .Z(n24340) );
  XOR U24532 ( .A(n24652), .B(n24653), .Z(n24648) );
  AND U24533 ( .A(n24654), .B(n24655), .Z(n24653) );
  XNOR U24534 ( .A(p_input[811]), .B(n24652), .Z(n24655) );
  XNOR U24535 ( .A(n24652), .B(n24349), .Z(n24654) );
  IV U24536 ( .A(p_input[779]), .Z(n24349) );
  XOR U24537 ( .A(n24656), .B(n24657), .Z(n24652) );
  AND U24538 ( .A(n24658), .B(n24659), .Z(n24657) );
  XNOR U24539 ( .A(p_input[810]), .B(n24656), .Z(n24659) );
  XNOR U24540 ( .A(n24656), .B(n24358), .Z(n24658) );
  IV U24541 ( .A(p_input[778]), .Z(n24358) );
  XOR U24542 ( .A(n24660), .B(n24661), .Z(n24656) );
  AND U24543 ( .A(n24662), .B(n24663), .Z(n24661) );
  XNOR U24544 ( .A(p_input[809]), .B(n24660), .Z(n24663) );
  XNOR U24545 ( .A(n24660), .B(n24367), .Z(n24662) );
  IV U24546 ( .A(p_input[777]), .Z(n24367) );
  XOR U24547 ( .A(n24664), .B(n24665), .Z(n24660) );
  AND U24548 ( .A(n24666), .B(n24667), .Z(n24665) );
  XNOR U24549 ( .A(p_input[808]), .B(n24664), .Z(n24667) );
  XNOR U24550 ( .A(n24664), .B(n24376), .Z(n24666) );
  IV U24551 ( .A(p_input[776]), .Z(n24376) );
  XOR U24552 ( .A(n24668), .B(n24669), .Z(n24664) );
  AND U24553 ( .A(n24670), .B(n24671), .Z(n24669) );
  XNOR U24554 ( .A(p_input[807]), .B(n24668), .Z(n24671) );
  XNOR U24555 ( .A(n24668), .B(n24385), .Z(n24670) );
  IV U24556 ( .A(p_input[775]), .Z(n24385) );
  XOR U24557 ( .A(n24672), .B(n24673), .Z(n24668) );
  AND U24558 ( .A(n24674), .B(n24675), .Z(n24673) );
  XNOR U24559 ( .A(p_input[806]), .B(n24672), .Z(n24675) );
  XNOR U24560 ( .A(n24672), .B(n24394), .Z(n24674) );
  IV U24561 ( .A(p_input[774]), .Z(n24394) );
  XOR U24562 ( .A(n24676), .B(n24677), .Z(n24672) );
  AND U24563 ( .A(n24678), .B(n24679), .Z(n24677) );
  XNOR U24564 ( .A(p_input[805]), .B(n24676), .Z(n24679) );
  XNOR U24565 ( .A(n24676), .B(n24403), .Z(n24678) );
  IV U24566 ( .A(p_input[773]), .Z(n24403) );
  XOR U24567 ( .A(n24680), .B(n24681), .Z(n24676) );
  AND U24568 ( .A(n24682), .B(n24683), .Z(n24681) );
  XNOR U24569 ( .A(p_input[804]), .B(n24680), .Z(n24683) );
  XNOR U24570 ( .A(n24680), .B(n24412), .Z(n24682) );
  IV U24571 ( .A(p_input[772]), .Z(n24412) );
  XOR U24572 ( .A(n24684), .B(n24685), .Z(n24680) );
  AND U24573 ( .A(n24686), .B(n24687), .Z(n24685) );
  XNOR U24574 ( .A(p_input[803]), .B(n24684), .Z(n24687) );
  XNOR U24575 ( .A(n24684), .B(n24421), .Z(n24686) );
  IV U24576 ( .A(p_input[771]), .Z(n24421) );
  XOR U24577 ( .A(n24688), .B(n24689), .Z(n24684) );
  AND U24578 ( .A(n24690), .B(n24691), .Z(n24689) );
  XNOR U24579 ( .A(p_input[802]), .B(n24688), .Z(n24691) );
  XNOR U24580 ( .A(n24688), .B(n24430), .Z(n24690) );
  IV U24581 ( .A(p_input[770]), .Z(n24430) );
  XNOR U24582 ( .A(n24692), .B(n24693), .Z(n24688) );
  AND U24583 ( .A(n24694), .B(n24695), .Z(n24693) );
  XOR U24584 ( .A(p_input[801]), .B(n24692), .Z(n24695) );
  XNOR U24585 ( .A(p_input[769]), .B(n24692), .Z(n24694) );
  AND U24586 ( .A(p_input[800]), .B(n24696), .Z(n24692) );
  IV U24587 ( .A(p_input[768]), .Z(n24696) );
  XOR U24588 ( .A(n24697), .B(n24698), .Z(n22875) );
  AND U24589 ( .A(n528), .B(n24699), .Z(n24698) );
  XNOR U24590 ( .A(n24700), .B(n24697), .Z(n24699) );
  XOR U24591 ( .A(n24701), .B(n24702), .Z(n528) );
  AND U24592 ( .A(n24703), .B(n24704), .Z(n24702) );
  XOR U24593 ( .A(n24701), .B(n22890), .Z(n24704) );
  XNOR U24594 ( .A(n24705), .B(n24706), .Z(n22890) );
  AND U24595 ( .A(n24707), .B(n398), .Z(n24706) );
  AND U24596 ( .A(n24705), .B(n24708), .Z(n24707) );
  XNOR U24597 ( .A(n22887), .B(n24701), .Z(n24703) );
  XOR U24598 ( .A(n24709), .B(n24710), .Z(n22887) );
  AND U24599 ( .A(n24711), .B(n395), .Z(n24710) );
  NOR U24600 ( .A(n24709), .B(n24712), .Z(n24711) );
  XOR U24601 ( .A(n24713), .B(n24714), .Z(n24701) );
  AND U24602 ( .A(n24715), .B(n24716), .Z(n24714) );
  XOR U24603 ( .A(n24713), .B(n22902), .Z(n24716) );
  XOR U24604 ( .A(n24717), .B(n24718), .Z(n22902) );
  AND U24605 ( .A(n398), .B(n24719), .Z(n24718) );
  XOR U24606 ( .A(n24720), .B(n24717), .Z(n24719) );
  XNOR U24607 ( .A(n22899), .B(n24713), .Z(n24715) );
  XOR U24608 ( .A(n24721), .B(n24722), .Z(n22899) );
  AND U24609 ( .A(n395), .B(n24723), .Z(n24722) );
  XOR U24610 ( .A(n24724), .B(n24721), .Z(n24723) );
  XOR U24611 ( .A(n24725), .B(n24726), .Z(n24713) );
  AND U24612 ( .A(n24727), .B(n24728), .Z(n24726) );
  XOR U24613 ( .A(n24725), .B(n22914), .Z(n24728) );
  XOR U24614 ( .A(n24729), .B(n24730), .Z(n22914) );
  AND U24615 ( .A(n398), .B(n24731), .Z(n24730) );
  XOR U24616 ( .A(n24732), .B(n24729), .Z(n24731) );
  XNOR U24617 ( .A(n22911), .B(n24725), .Z(n24727) );
  XOR U24618 ( .A(n24733), .B(n24734), .Z(n22911) );
  AND U24619 ( .A(n395), .B(n24735), .Z(n24734) );
  XOR U24620 ( .A(n24736), .B(n24733), .Z(n24735) );
  XOR U24621 ( .A(n24737), .B(n24738), .Z(n24725) );
  AND U24622 ( .A(n24739), .B(n24740), .Z(n24738) );
  XOR U24623 ( .A(n24737), .B(n22926), .Z(n24740) );
  XOR U24624 ( .A(n24741), .B(n24742), .Z(n22926) );
  AND U24625 ( .A(n398), .B(n24743), .Z(n24742) );
  XOR U24626 ( .A(n24744), .B(n24741), .Z(n24743) );
  XNOR U24627 ( .A(n22923), .B(n24737), .Z(n24739) );
  XOR U24628 ( .A(n24745), .B(n24746), .Z(n22923) );
  AND U24629 ( .A(n395), .B(n24747), .Z(n24746) );
  XOR U24630 ( .A(n24748), .B(n24745), .Z(n24747) );
  XOR U24631 ( .A(n24749), .B(n24750), .Z(n24737) );
  AND U24632 ( .A(n24751), .B(n24752), .Z(n24750) );
  XOR U24633 ( .A(n24749), .B(n22938), .Z(n24752) );
  XOR U24634 ( .A(n24753), .B(n24754), .Z(n22938) );
  AND U24635 ( .A(n398), .B(n24755), .Z(n24754) );
  XOR U24636 ( .A(n24756), .B(n24753), .Z(n24755) );
  XNOR U24637 ( .A(n22935), .B(n24749), .Z(n24751) );
  XOR U24638 ( .A(n24757), .B(n24758), .Z(n22935) );
  AND U24639 ( .A(n395), .B(n24759), .Z(n24758) );
  XOR U24640 ( .A(n24760), .B(n24757), .Z(n24759) );
  XOR U24641 ( .A(n24761), .B(n24762), .Z(n24749) );
  AND U24642 ( .A(n24763), .B(n24764), .Z(n24762) );
  XOR U24643 ( .A(n24761), .B(n22950), .Z(n24764) );
  XOR U24644 ( .A(n24765), .B(n24766), .Z(n22950) );
  AND U24645 ( .A(n398), .B(n24767), .Z(n24766) );
  XOR U24646 ( .A(n24768), .B(n24765), .Z(n24767) );
  XNOR U24647 ( .A(n22947), .B(n24761), .Z(n24763) );
  XOR U24648 ( .A(n24769), .B(n24770), .Z(n22947) );
  AND U24649 ( .A(n395), .B(n24771), .Z(n24770) );
  XOR U24650 ( .A(n24772), .B(n24769), .Z(n24771) );
  XOR U24651 ( .A(n24773), .B(n24774), .Z(n24761) );
  AND U24652 ( .A(n24775), .B(n24776), .Z(n24774) );
  XOR U24653 ( .A(n24773), .B(n22962), .Z(n24776) );
  XOR U24654 ( .A(n24777), .B(n24778), .Z(n22962) );
  AND U24655 ( .A(n398), .B(n24779), .Z(n24778) );
  XOR U24656 ( .A(n24780), .B(n24777), .Z(n24779) );
  XNOR U24657 ( .A(n22959), .B(n24773), .Z(n24775) );
  XOR U24658 ( .A(n24781), .B(n24782), .Z(n22959) );
  AND U24659 ( .A(n395), .B(n24783), .Z(n24782) );
  XOR U24660 ( .A(n24784), .B(n24781), .Z(n24783) );
  XOR U24661 ( .A(n24785), .B(n24786), .Z(n24773) );
  AND U24662 ( .A(n24787), .B(n24788), .Z(n24786) );
  XOR U24663 ( .A(n24785), .B(n22974), .Z(n24788) );
  XOR U24664 ( .A(n24789), .B(n24790), .Z(n22974) );
  AND U24665 ( .A(n398), .B(n24791), .Z(n24790) );
  XOR U24666 ( .A(n24792), .B(n24789), .Z(n24791) );
  XNOR U24667 ( .A(n22971), .B(n24785), .Z(n24787) );
  XOR U24668 ( .A(n24793), .B(n24794), .Z(n22971) );
  AND U24669 ( .A(n395), .B(n24795), .Z(n24794) );
  XOR U24670 ( .A(n24796), .B(n24793), .Z(n24795) );
  XOR U24671 ( .A(n24797), .B(n24798), .Z(n24785) );
  AND U24672 ( .A(n24799), .B(n24800), .Z(n24798) );
  XOR U24673 ( .A(n24797), .B(n22986), .Z(n24800) );
  XOR U24674 ( .A(n24801), .B(n24802), .Z(n22986) );
  AND U24675 ( .A(n398), .B(n24803), .Z(n24802) );
  XOR U24676 ( .A(n24804), .B(n24801), .Z(n24803) );
  XNOR U24677 ( .A(n22983), .B(n24797), .Z(n24799) );
  XOR U24678 ( .A(n24805), .B(n24806), .Z(n22983) );
  AND U24679 ( .A(n395), .B(n24807), .Z(n24806) );
  XOR U24680 ( .A(n24808), .B(n24805), .Z(n24807) );
  XOR U24681 ( .A(n24809), .B(n24810), .Z(n24797) );
  AND U24682 ( .A(n24811), .B(n24812), .Z(n24810) );
  XOR U24683 ( .A(n24809), .B(n22998), .Z(n24812) );
  XOR U24684 ( .A(n24813), .B(n24814), .Z(n22998) );
  AND U24685 ( .A(n398), .B(n24815), .Z(n24814) );
  XOR U24686 ( .A(n24816), .B(n24813), .Z(n24815) );
  XNOR U24687 ( .A(n22995), .B(n24809), .Z(n24811) );
  XOR U24688 ( .A(n24817), .B(n24818), .Z(n22995) );
  AND U24689 ( .A(n395), .B(n24819), .Z(n24818) );
  XOR U24690 ( .A(n24820), .B(n24817), .Z(n24819) );
  XOR U24691 ( .A(n24821), .B(n24822), .Z(n24809) );
  AND U24692 ( .A(n24823), .B(n24824), .Z(n24822) );
  XOR U24693 ( .A(n24821), .B(n23010), .Z(n24824) );
  XOR U24694 ( .A(n24825), .B(n24826), .Z(n23010) );
  AND U24695 ( .A(n398), .B(n24827), .Z(n24826) );
  XOR U24696 ( .A(n24828), .B(n24825), .Z(n24827) );
  XNOR U24697 ( .A(n23007), .B(n24821), .Z(n24823) );
  XOR U24698 ( .A(n24829), .B(n24830), .Z(n23007) );
  AND U24699 ( .A(n395), .B(n24831), .Z(n24830) );
  XOR U24700 ( .A(n24832), .B(n24829), .Z(n24831) );
  XOR U24701 ( .A(n24833), .B(n24834), .Z(n24821) );
  AND U24702 ( .A(n24835), .B(n24836), .Z(n24834) );
  XOR U24703 ( .A(n24833), .B(n23022), .Z(n24836) );
  XOR U24704 ( .A(n24837), .B(n24838), .Z(n23022) );
  AND U24705 ( .A(n398), .B(n24839), .Z(n24838) );
  XOR U24706 ( .A(n24840), .B(n24837), .Z(n24839) );
  XNOR U24707 ( .A(n23019), .B(n24833), .Z(n24835) );
  XOR U24708 ( .A(n24841), .B(n24842), .Z(n23019) );
  AND U24709 ( .A(n395), .B(n24843), .Z(n24842) );
  XOR U24710 ( .A(n24844), .B(n24841), .Z(n24843) );
  XOR U24711 ( .A(n24845), .B(n24846), .Z(n24833) );
  AND U24712 ( .A(n24847), .B(n24848), .Z(n24846) );
  XOR U24713 ( .A(n24845), .B(n23034), .Z(n24848) );
  XOR U24714 ( .A(n24849), .B(n24850), .Z(n23034) );
  AND U24715 ( .A(n398), .B(n24851), .Z(n24850) );
  XOR U24716 ( .A(n24852), .B(n24849), .Z(n24851) );
  XNOR U24717 ( .A(n23031), .B(n24845), .Z(n24847) );
  XOR U24718 ( .A(n24853), .B(n24854), .Z(n23031) );
  AND U24719 ( .A(n395), .B(n24855), .Z(n24854) );
  XOR U24720 ( .A(n24856), .B(n24853), .Z(n24855) );
  XOR U24721 ( .A(n24857), .B(n24858), .Z(n24845) );
  AND U24722 ( .A(n24859), .B(n24860), .Z(n24858) );
  XOR U24723 ( .A(n24857), .B(n23046), .Z(n24860) );
  XOR U24724 ( .A(n24861), .B(n24862), .Z(n23046) );
  AND U24725 ( .A(n398), .B(n24863), .Z(n24862) );
  XOR U24726 ( .A(n24864), .B(n24861), .Z(n24863) );
  XNOR U24727 ( .A(n23043), .B(n24857), .Z(n24859) );
  XOR U24728 ( .A(n24865), .B(n24866), .Z(n23043) );
  AND U24729 ( .A(n395), .B(n24867), .Z(n24866) );
  XOR U24730 ( .A(n24868), .B(n24865), .Z(n24867) );
  XOR U24731 ( .A(n24869), .B(n24870), .Z(n24857) );
  AND U24732 ( .A(n24871), .B(n24872), .Z(n24870) );
  XOR U24733 ( .A(n24869), .B(n23058), .Z(n24872) );
  XOR U24734 ( .A(n24873), .B(n24874), .Z(n23058) );
  AND U24735 ( .A(n398), .B(n24875), .Z(n24874) );
  XOR U24736 ( .A(n24876), .B(n24873), .Z(n24875) );
  XNOR U24737 ( .A(n23055), .B(n24869), .Z(n24871) );
  XOR U24738 ( .A(n24877), .B(n24878), .Z(n23055) );
  AND U24739 ( .A(n395), .B(n24879), .Z(n24878) );
  XOR U24740 ( .A(n24880), .B(n24877), .Z(n24879) );
  XOR U24741 ( .A(n24881), .B(n24882), .Z(n24869) );
  AND U24742 ( .A(n24883), .B(n24884), .Z(n24882) );
  XOR U24743 ( .A(n24881), .B(n23070), .Z(n24884) );
  XOR U24744 ( .A(n24885), .B(n24886), .Z(n23070) );
  AND U24745 ( .A(n398), .B(n24887), .Z(n24886) );
  XOR U24746 ( .A(n24888), .B(n24885), .Z(n24887) );
  XNOR U24747 ( .A(n23067), .B(n24881), .Z(n24883) );
  XOR U24748 ( .A(n24889), .B(n24890), .Z(n23067) );
  AND U24749 ( .A(n395), .B(n24891), .Z(n24890) );
  XOR U24750 ( .A(n24892), .B(n24889), .Z(n24891) );
  XOR U24751 ( .A(n24893), .B(n24894), .Z(n24881) );
  AND U24752 ( .A(n24895), .B(n24896), .Z(n24894) );
  XOR U24753 ( .A(n24893), .B(n23082), .Z(n24896) );
  XOR U24754 ( .A(n24897), .B(n24898), .Z(n23082) );
  AND U24755 ( .A(n398), .B(n24899), .Z(n24898) );
  XOR U24756 ( .A(n24900), .B(n24897), .Z(n24899) );
  XNOR U24757 ( .A(n23079), .B(n24893), .Z(n24895) );
  XOR U24758 ( .A(n24901), .B(n24902), .Z(n23079) );
  AND U24759 ( .A(n395), .B(n24903), .Z(n24902) );
  XOR U24760 ( .A(n24904), .B(n24901), .Z(n24903) );
  XOR U24761 ( .A(n24905), .B(n24906), .Z(n24893) );
  AND U24762 ( .A(n24907), .B(n24908), .Z(n24906) );
  XOR U24763 ( .A(n24905), .B(n23094), .Z(n24908) );
  XOR U24764 ( .A(n24909), .B(n24910), .Z(n23094) );
  AND U24765 ( .A(n398), .B(n24911), .Z(n24910) );
  XOR U24766 ( .A(n24912), .B(n24909), .Z(n24911) );
  XNOR U24767 ( .A(n23091), .B(n24905), .Z(n24907) );
  XOR U24768 ( .A(n24913), .B(n24914), .Z(n23091) );
  AND U24769 ( .A(n395), .B(n24915), .Z(n24914) );
  XOR U24770 ( .A(n24916), .B(n24913), .Z(n24915) );
  XOR U24771 ( .A(n24917), .B(n24918), .Z(n24905) );
  AND U24772 ( .A(n24919), .B(n24920), .Z(n24918) );
  XOR U24773 ( .A(n24917), .B(n23106), .Z(n24920) );
  XOR U24774 ( .A(n24921), .B(n24922), .Z(n23106) );
  AND U24775 ( .A(n398), .B(n24923), .Z(n24922) );
  XOR U24776 ( .A(n24924), .B(n24921), .Z(n24923) );
  XNOR U24777 ( .A(n23103), .B(n24917), .Z(n24919) );
  XOR U24778 ( .A(n24925), .B(n24926), .Z(n23103) );
  AND U24779 ( .A(n395), .B(n24927), .Z(n24926) );
  XOR U24780 ( .A(n24928), .B(n24925), .Z(n24927) );
  XOR U24781 ( .A(n24929), .B(n24930), .Z(n24917) );
  AND U24782 ( .A(n24931), .B(n24932), .Z(n24930) );
  XOR U24783 ( .A(n24929), .B(n23118), .Z(n24932) );
  XOR U24784 ( .A(n24933), .B(n24934), .Z(n23118) );
  AND U24785 ( .A(n398), .B(n24935), .Z(n24934) );
  XOR U24786 ( .A(n24936), .B(n24933), .Z(n24935) );
  XNOR U24787 ( .A(n23115), .B(n24929), .Z(n24931) );
  XOR U24788 ( .A(n24937), .B(n24938), .Z(n23115) );
  AND U24789 ( .A(n395), .B(n24939), .Z(n24938) );
  XOR U24790 ( .A(n24940), .B(n24937), .Z(n24939) );
  XOR U24791 ( .A(n24941), .B(n24942), .Z(n24929) );
  AND U24792 ( .A(n24943), .B(n24944), .Z(n24942) );
  XOR U24793 ( .A(n24941), .B(n23130), .Z(n24944) );
  XOR U24794 ( .A(n24945), .B(n24946), .Z(n23130) );
  AND U24795 ( .A(n398), .B(n24947), .Z(n24946) );
  XOR U24796 ( .A(n24948), .B(n24945), .Z(n24947) );
  XNOR U24797 ( .A(n23127), .B(n24941), .Z(n24943) );
  XOR U24798 ( .A(n24949), .B(n24950), .Z(n23127) );
  AND U24799 ( .A(n395), .B(n24951), .Z(n24950) );
  XOR U24800 ( .A(n24952), .B(n24949), .Z(n24951) );
  XOR U24801 ( .A(n24953), .B(n24954), .Z(n24941) );
  AND U24802 ( .A(n24955), .B(n24956), .Z(n24954) );
  XOR U24803 ( .A(n24953), .B(n23142), .Z(n24956) );
  XOR U24804 ( .A(n24957), .B(n24958), .Z(n23142) );
  AND U24805 ( .A(n398), .B(n24959), .Z(n24958) );
  XOR U24806 ( .A(n24960), .B(n24957), .Z(n24959) );
  XNOR U24807 ( .A(n23139), .B(n24953), .Z(n24955) );
  XOR U24808 ( .A(n24961), .B(n24962), .Z(n23139) );
  AND U24809 ( .A(n395), .B(n24963), .Z(n24962) );
  XOR U24810 ( .A(n24964), .B(n24961), .Z(n24963) );
  XOR U24811 ( .A(n24965), .B(n24966), .Z(n24953) );
  AND U24812 ( .A(n24967), .B(n24968), .Z(n24966) );
  XOR U24813 ( .A(n24965), .B(n23154), .Z(n24968) );
  XOR U24814 ( .A(n24969), .B(n24970), .Z(n23154) );
  AND U24815 ( .A(n398), .B(n24971), .Z(n24970) );
  XOR U24816 ( .A(n24972), .B(n24969), .Z(n24971) );
  XNOR U24817 ( .A(n23151), .B(n24965), .Z(n24967) );
  XOR U24818 ( .A(n24973), .B(n24974), .Z(n23151) );
  AND U24819 ( .A(n395), .B(n24975), .Z(n24974) );
  XOR U24820 ( .A(n24976), .B(n24973), .Z(n24975) );
  XOR U24821 ( .A(n24977), .B(n24978), .Z(n24965) );
  AND U24822 ( .A(n24979), .B(n24980), .Z(n24978) );
  XOR U24823 ( .A(n24977), .B(n23166), .Z(n24980) );
  XOR U24824 ( .A(n24981), .B(n24982), .Z(n23166) );
  AND U24825 ( .A(n398), .B(n24983), .Z(n24982) );
  XOR U24826 ( .A(n24984), .B(n24981), .Z(n24983) );
  XNOR U24827 ( .A(n23163), .B(n24977), .Z(n24979) );
  XOR U24828 ( .A(n24985), .B(n24986), .Z(n23163) );
  AND U24829 ( .A(n395), .B(n24987), .Z(n24986) );
  XOR U24830 ( .A(n24988), .B(n24985), .Z(n24987) );
  XOR U24831 ( .A(n24989), .B(n24990), .Z(n24977) );
  AND U24832 ( .A(n24991), .B(n24992), .Z(n24990) );
  XOR U24833 ( .A(n24989), .B(n23178), .Z(n24992) );
  XOR U24834 ( .A(n24993), .B(n24994), .Z(n23178) );
  AND U24835 ( .A(n398), .B(n24995), .Z(n24994) );
  XOR U24836 ( .A(n24996), .B(n24993), .Z(n24995) );
  XNOR U24837 ( .A(n23175), .B(n24989), .Z(n24991) );
  XOR U24838 ( .A(n24997), .B(n24998), .Z(n23175) );
  AND U24839 ( .A(n395), .B(n24999), .Z(n24998) );
  XOR U24840 ( .A(n25000), .B(n24997), .Z(n24999) );
  XOR U24841 ( .A(n25001), .B(n25002), .Z(n24989) );
  AND U24842 ( .A(n25003), .B(n25004), .Z(n25002) );
  XOR U24843 ( .A(n25001), .B(n23190), .Z(n25004) );
  XOR U24844 ( .A(n25005), .B(n25006), .Z(n23190) );
  AND U24845 ( .A(n398), .B(n25007), .Z(n25006) );
  XOR U24846 ( .A(n25008), .B(n25005), .Z(n25007) );
  XNOR U24847 ( .A(n23187), .B(n25001), .Z(n25003) );
  XOR U24848 ( .A(n25009), .B(n25010), .Z(n23187) );
  AND U24849 ( .A(n395), .B(n25011), .Z(n25010) );
  XOR U24850 ( .A(n25012), .B(n25009), .Z(n25011) );
  XOR U24851 ( .A(n25013), .B(n25014), .Z(n25001) );
  AND U24852 ( .A(n25015), .B(n25016), .Z(n25014) );
  XOR U24853 ( .A(n25013), .B(n23202), .Z(n25016) );
  XOR U24854 ( .A(n25017), .B(n25018), .Z(n23202) );
  AND U24855 ( .A(n398), .B(n25019), .Z(n25018) );
  XOR U24856 ( .A(n25020), .B(n25017), .Z(n25019) );
  XNOR U24857 ( .A(n23199), .B(n25013), .Z(n25015) );
  XOR U24858 ( .A(n25021), .B(n25022), .Z(n23199) );
  AND U24859 ( .A(n395), .B(n25023), .Z(n25022) );
  XOR U24860 ( .A(n25024), .B(n25021), .Z(n25023) );
  XOR U24861 ( .A(n25025), .B(n25026), .Z(n25013) );
  AND U24862 ( .A(n25027), .B(n25028), .Z(n25026) );
  XOR U24863 ( .A(n25025), .B(n23214), .Z(n25028) );
  XOR U24864 ( .A(n25029), .B(n25030), .Z(n23214) );
  AND U24865 ( .A(n398), .B(n25031), .Z(n25030) );
  XOR U24866 ( .A(n25032), .B(n25029), .Z(n25031) );
  XNOR U24867 ( .A(n23211), .B(n25025), .Z(n25027) );
  XOR U24868 ( .A(n25033), .B(n25034), .Z(n23211) );
  AND U24869 ( .A(n395), .B(n25035), .Z(n25034) );
  XOR U24870 ( .A(n25036), .B(n25033), .Z(n25035) );
  XOR U24871 ( .A(n25037), .B(n25038), .Z(n25025) );
  AND U24872 ( .A(n25039), .B(n25040), .Z(n25038) );
  XOR U24873 ( .A(n25037), .B(n23226), .Z(n25040) );
  XOR U24874 ( .A(n25041), .B(n25042), .Z(n23226) );
  AND U24875 ( .A(n398), .B(n25043), .Z(n25042) );
  XOR U24876 ( .A(n25044), .B(n25041), .Z(n25043) );
  XNOR U24877 ( .A(n23223), .B(n25037), .Z(n25039) );
  XOR U24878 ( .A(n25045), .B(n25046), .Z(n23223) );
  AND U24879 ( .A(n395), .B(n25047), .Z(n25046) );
  XOR U24880 ( .A(n25048), .B(n25045), .Z(n25047) );
  XOR U24881 ( .A(n25049), .B(n25050), .Z(n25037) );
  AND U24882 ( .A(n25051), .B(n25052), .Z(n25050) );
  XOR U24883 ( .A(n23238), .B(n25049), .Z(n25052) );
  XOR U24884 ( .A(n25053), .B(n25054), .Z(n23238) );
  AND U24885 ( .A(n398), .B(n25055), .Z(n25054) );
  XOR U24886 ( .A(n25053), .B(n25056), .Z(n25055) );
  XNOR U24887 ( .A(n25049), .B(n23235), .Z(n25051) );
  XOR U24888 ( .A(n25057), .B(n25058), .Z(n23235) );
  AND U24889 ( .A(n395), .B(n25059), .Z(n25058) );
  XOR U24890 ( .A(n25057), .B(n25060), .Z(n25059) );
  XOR U24891 ( .A(n25061), .B(n25062), .Z(n25049) );
  AND U24892 ( .A(n25063), .B(n25064), .Z(n25062) );
  XNOR U24893 ( .A(n25065), .B(n23251), .Z(n25064) );
  XOR U24894 ( .A(n25066), .B(n25067), .Z(n23251) );
  AND U24895 ( .A(n398), .B(n25068), .Z(n25067) );
  XOR U24896 ( .A(n25069), .B(n25066), .Z(n25068) );
  XNOR U24897 ( .A(n23248), .B(n25061), .Z(n25063) );
  XOR U24898 ( .A(n25070), .B(n25071), .Z(n23248) );
  AND U24899 ( .A(n395), .B(n25072), .Z(n25071) );
  XOR U24900 ( .A(n25073), .B(n25070), .Z(n25072) );
  IV U24901 ( .A(n25065), .Z(n25061) );
  AND U24902 ( .A(n24697), .B(n24700), .Z(n25065) );
  XNOR U24903 ( .A(n25074), .B(n25075), .Z(n24700) );
  AND U24904 ( .A(n398), .B(n25076), .Z(n25075) );
  XNOR U24905 ( .A(n25077), .B(n25074), .Z(n25076) );
  XOR U24906 ( .A(n25078), .B(n25079), .Z(n398) );
  AND U24907 ( .A(n25080), .B(n25081), .Z(n25079) );
  XOR U24908 ( .A(n24708), .B(n25078), .Z(n25081) );
  IV U24909 ( .A(n25082), .Z(n24708) );
  AND U24910 ( .A(p_input[767]), .B(p_input[735]), .Z(n25082) );
  XOR U24911 ( .A(n25078), .B(n24705), .Z(n25080) );
  AND U24912 ( .A(p_input[671]), .B(p_input[703]), .Z(n24705) );
  XOR U24913 ( .A(n25083), .B(n25084), .Z(n25078) );
  AND U24914 ( .A(n25085), .B(n25086), .Z(n25084) );
  XOR U24915 ( .A(n25083), .B(n24720), .Z(n25086) );
  XNOR U24916 ( .A(p_input[734]), .B(n25087), .Z(n24720) );
  AND U24917 ( .A(n562), .B(n25088), .Z(n25087) );
  XOR U24918 ( .A(p_input[766]), .B(p_input[734]), .Z(n25088) );
  XNOR U24919 ( .A(n24717), .B(n25083), .Z(n25085) );
  XOR U24920 ( .A(n25089), .B(n25090), .Z(n24717) );
  AND U24921 ( .A(n560), .B(n25091), .Z(n25090) );
  XOR U24922 ( .A(p_input[702]), .B(p_input[670]), .Z(n25091) );
  XOR U24923 ( .A(n25092), .B(n25093), .Z(n25083) );
  AND U24924 ( .A(n25094), .B(n25095), .Z(n25093) );
  XOR U24925 ( .A(n25092), .B(n24732), .Z(n25095) );
  XNOR U24926 ( .A(p_input[733]), .B(n25096), .Z(n24732) );
  AND U24927 ( .A(n562), .B(n25097), .Z(n25096) );
  XOR U24928 ( .A(p_input[765]), .B(p_input[733]), .Z(n25097) );
  XNOR U24929 ( .A(n24729), .B(n25092), .Z(n25094) );
  XOR U24930 ( .A(n25098), .B(n25099), .Z(n24729) );
  AND U24931 ( .A(n560), .B(n25100), .Z(n25099) );
  XOR U24932 ( .A(p_input[701]), .B(p_input[669]), .Z(n25100) );
  XOR U24933 ( .A(n25101), .B(n25102), .Z(n25092) );
  AND U24934 ( .A(n25103), .B(n25104), .Z(n25102) );
  XOR U24935 ( .A(n25101), .B(n24744), .Z(n25104) );
  XNOR U24936 ( .A(p_input[732]), .B(n25105), .Z(n24744) );
  AND U24937 ( .A(n562), .B(n25106), .Z(n25105) );
  XOR U24938 ( .A(p_input[764]), .B(p_input[732]), .Z(n25106) );
  XNOR U24939 ( .A(n24741), .B(n25101), .Z(n25103) );
  XOR U24940 ( .A(n25107), .B(n25108), .Z(n24741) );
  AND U24941 ( .A(n560), .B(n25109), .Z(n25108) );
  XOR U24942 ( .A(p_input[700]), .B(p_input[668]), .Z(n25109) );
  XOR U24943 ( .A(n25110), .B(n25111), .Z(n25101) );
  AND U24944 ( .A(n25112), .B(n25113), .Z(n25111) );
  XOR U24945 ( .A(n25110), .B(n24756), .Z(n25113) );
  XNOR U24946 ( .A(p_input[731]), .B(n25114), .Z(n24756) );
  AND U24947 ( .A(n562), .B(n25115), .Z(n25114) );
  XOR U24948 ( .A(p_input[763]), .B(p_input[731]), .Z(n25115) );
  XNOR U24949 ( .A(n24753), .B(n25110), .Z(n25112) );
  XOR U24950 ( .A(n25116), .B(n25117), .Z(n24753) );
  AND U24951 ( .A(n560), .B(n25118), .Z(n25117) );
  XOR U24952 ( .A(p_input[699]), .B(p_input[667]), .Z(n25118) );
  XOR U24953 ( .A(n25119), .B(n25120), .Z(n25110) );
  AND U24954 ( .A(n25121), .B(n25122), .Z(n25120) );
  XOR U24955 ( .A(n25119), .B(n24768), .Z(n25122) );
  XNOR U24956 ( .A(p_input[730]), .B(n25123), .Z(n24768) );
  AND U24957 ( .A(n562), .B(n25124), .Z(n25123) );
  XOR U24958 ( .A(p_input[762]), .B(p_input[730]), .Z(n25124) );
  XNOR U24959 ( .A(n24765), .B(n25119), .Z(n25121) );
  XOR U24960 ( .A(n25125), .B(n25126), .Z(n24765) );
  AND U24961 ( .A(n560), .B(n25127), .Z(n25126) );
  XOR U24962 ( .A(p_input[698]), .B(p_input[666]), .Z(n25127) );
  XOR U24963 ( .A(n25128), .B(n25129), .Z(n25119) );
  AND U24964 ( .A(n25130), .B(n25131), .Z(n25129) );
  XOR U24965 ( .A(n25128), .B(n24780), .Z(n25131) );
  XNOR U24966 ( .A(p_input[729]), .B(n25132), .Z(n24780) );
  AND U24967 ( .A(n562), .B(n25133), .Z(n25132) );
  XOR U24968 ( .A(p_input[761]), .B(p_input[729]), .Z(n25133) );
  XNOR U24969 ( .A(n24777), .B(n25128), .Z(n25130) );
  XOR U24970 ( .A(n25134), .B(n25135), .Z(n24777) );
  AND U24971 ( .A(n560), .B(n25136), .Z(n25135) );
  XOR U24972 ( .A(p_input[697]), .B(p_input[665]), .Z(n25136) );
  XOR U24973 ( .A(n25137), .B(n25138), .Z(n25128) );
  AND U24974 ( .A(n25139), .B(n25140), .Z(n25138) );
  XOR U24975 ( .A(n25137), .B(n24792), .Z(n25140) );
  XNOR U24976 ( .A(p_input[728]), .B(n25141), .Z(n24792) );
  AND U24977 ( .A(n562), .B(n25142), .Z(n25141) );
  XOR U24978 ( .A(p_input[760]), .B(p_input[728]), .Z(n25142) );
  XNOR U24979 ( .A(n24789), .B(n25137), .Z(n25139) );
  XOR U24980 ( .A(n25143), .B(n25144), .Z(n24789) );
  AND U24981 ( .A(n560), .B(n25145), .Z(n25144) );
  XOR U24982 ( .A(p_input[696]), .B(p_input[664]), .Z(n25145) );
  XOR U24983 ( .A(n25146), .B(n25147), .Z(n25137) );
  AND U24984 ( .A(n25148), .B(n25149), .Z(n25147) );
  XOR U24985 ( .A(n25146), .B(n24804), .Z(n25149) );
  XNOR U24986 ( .A(p_input[727]), .B(n25150), .Z(n24804) );
  AND U24987 ( .A(n562), .B(n25151), .Z(n25150) );
  XOR U24988 ( .A(p_input[759]), .B(p_input[727]), .Z(n25151) );
  XNOR U24989 ( .A(n24801), .B(n25146), .Z(n25148) );
  XOR U24990 ( .A(n25152), .B(n25153), .Z(n24801) );
  AND U24991 ( .A(n560), .B(n25154), .Z(n25153) );
  XOR U24992 ( .A(p_input[695]), .B(p_input[663]), .Z(n25154) );
  XOR U24993 ( .A(n25155), .B(n25156), .Z(n25146) );
  AND U24994 ( .A(n25157), .B(n25158), .Z(n25156) );
  XOR U24995 ( .A(n25155), .B(n24816), .Z(n25158) );
  XNOR U24996 ( .A(p_input[726]), .B(n25159), .Z(n24816) );
  AND U24997 ( .A(n562), .B(n25160), .Z(n25159) );
  XOR U24998 ( .A(p_input[758]), .B(p_input[726]), .Z(n25160) );
  XNOR U24999 ( .A(n24813), .B(n25155), .Z(n25157) );
  XOR U25000 ( .A(n25161), .B(n25162), .Z(n24813) );
  AND U25001 ( .A(n560), .B(n25163), .Z(n25162) );
  XOR U25002 ( .A(p_input[694]), .B(p_input[662]), .Z(n25163) );
  XOR U25003 ( .A(n25164), .B(n25165), .Z(n25155) );
  AND U25004 ( .A(n25166), .B(n25167), .Z(n25165) );
  XOR U25005 ( .A(n25164), .B(n24828), .Z(n25167) );
  XNOR U25006 ( .A(p_input[725]), .B(n25168), .Z(n24828) );
  AND U25007 ( .A(n562), .B(n25169), .Z(n25168) );
  XOR U25008 ( .A(p_input[757]), .B(p_input[725]), .Z(n25169) );
  XNOR U25009 ( .A(n24825), .B(n25164), .Z(n25166) );
  XOR U25010 ( .A(n25170), .B(n25171), .Z(n24825) );
  AND U25011 ( .A(n560), .B(n25172), .Z(n25171) );
  XOR U25012 ( .A(p_input[693]), .B(p_input[661]), .Z(n25172) );
  XOR U25013 ( .A(n25173), .B(n25174), .Z(n25164) );
  AND U25014 ( .A(n25175), .B(n25176), .Z(n25174) );
  XOR U25015 ( .A(n25173), .B(n24840), .Z(n25176) );
  XNOR U25016 ( .A(p_input[724]), .B(n25177), .Z(n24840) );
  AND U25017 ( .A(n562), .B(n25178), .Z(n25177) );
  XOR U25018 ( .A(p_input[756]), .B(p_input[724]), .Z(n25178) );
  XNOR U25019 ( .A(n24837), .B(n25173), .Z(n25175) );
  XOR U25020 ( .A(n25179), .B(n25180), .Z(n24837) );
  AND U25021 ( .A(n560), .B(n25181), .Z(n25180) );
  XOR U25022 ( .A(p_input[692]), .B(p_input[660]), .Z(n25181) );
  XOR U25023 ( .A(n25182), .B(n25183), .Z(n25173) );
  AND U25024 ( .A(n25184), .B(n25185), .Z(n25183) );
  XOR U25025 ( .A(n25182), .B(n24852), .Z(n25185) );
  XNOR U25026 ( .A(p_input[723]), .B(n25186), .Z(n24852) );
  AND U25027 ( .A(n562), .B(n25187), .Z(n25186) );
  XOR U25028 ( .A(p_input[755]), .B(p_input[723]), .Z(n25187) );
  XNOR U25029 ( .A(n24849), .B(n25182), .Z(n25184) );
  XOR U25030 ( .A(n25188), .B(n25189), .Z(n24849) );
  AND U25031 ( .A(n560), .B(n25190), .Z(n25189) );
  XOR U25032 ( .A(p_input[691]), .B(p_input[659]), .Z(n25190) );
  XOR U25033 ( .A(n25191), .B(n25192), .Z(n25182) );
  AND U25034 ( .A(n25193), .B(n25194), .Z(n25192) );
  XOR U25035 ( .A(n25191), .B(n24864), .Z(n25194) );
  XNOR U25036 ( .A(p_input[722]), .B(n25195), .Z(n24864) );
  AND U25037 ( .A(n562), .B(n25196), .Z(n25195) );
  XOR U25038 ( .A(p_input[754]), .B(p_input[722]), .Z(n25196) );
  XNOR U25039 ( .A(n24861), .B(n25191), .Z(n25193) );
  XOR U25040 ( .A(n25197), .B(n25198), .Z(n24861) );
  AND U25041 ( .A(n560), .B(n25199), .Z(n25198) );
  XOR U25042 ( .A(p_input[690]), .B(p_input[658]), .Z(n25199) );
  XOR U25043 ( .A(n25200), .B(n25201), .Z(n25191) );
  AND U25044 ( .A(n25202), .B(n25203), .Z(n25201) );
  XOR U25045 ( .A(n25200), .B(n24876), .Z(n25203) );
  XNOR U25046 ( .A(p_input[721]), .B(n25204), .Z(n24876) );
  AND U25047 ( .A(n562), .B(n25205), .Z(n25204) );
  XOR U25048 ( .A(p_input[753]), .B(p_input[721]), .Z(n25205) );
  XNOR U25049 ( .A(n24873), .B(n25200), .Z(n25202) );
  XOR U25050 ( .A(n25206), .B(n25207), .Z(n24873) );
  AND U25051 ( .A(n560), .B(n25208), .Z(n25207) );
  XOR U25052 ( .A(p_input[689]), .B(p_input[657]), .Z(n25208) );
  XOR U25053 ( .A(n25209), .B(n25210), .Z(n25200) );
  AND U25054 ( .A(n25211), .B(n25212), .Z(n25210) );
  XOR U25055 ( .A(n25209), .B(n24888), .Z(n25212) );
  XNOR U25056 ( .A(p_input[720]), .B(n25213), .Z(n24888) );
  AND U25057 ( .A(n562), .B(n25214), .Z(n25213) );
  XOR U25058 ( .A(p_input[752]), .B(p_input[720]), .Z(n25214) );
  XNOR U25059 ( .A(n24885), .B(n25209), .Z(n25211) );
  XOR U25060 ( .A(n25215), .B(n25216), .Z(n24885) );
  AND U25061 ( .A(n560), .B(n25217), .Z(n25216) );
  XOR U25062 ( .A(p_input[688]), .B(p_input[656]), .Z(n25217) );
  XOR U25063 ( .A(n25218), .B(n25219), .Z(n25209) );
  AND U25064 ( .A(n25220), .B(n25221), .Z(n25219) );
  XOR U25065 ( .A(n25218), .B(n24900), .Z(n25221) );
  XNOR U25066 ( .A(p_input[719]), .B(n25222), .Z(n24900) );
  AND U25067 ( .A(n562), .B(n25223), .Z(n25222) );
  XOR U25068 ( .A(p_input[751]), .B(p_input[719]), .Z(n25223) );
  XNOR U25069 ( .A(n24897), .B(n25218), .Z(n25220) );
  XOR U25070 ( .A(n25224), .B(n25225), .Z(n24897) );
  AND U25071 ( .A(n560), .B(n25226), .Z(n25225) );
  XOR U25072 ( .A(p_input[687]), .B(p_input[655]), .Z(n25226) );
  XOR U25073 ( .A(n25227), .B(n25228), .Z(n25218) );
  AND U25074 ( .A(n25229), .B(n25230), .Z(n25228) );
  XOR U25075 ( .A(n25227), .B(n24912), .Z(n25230) );
  XNOR U25076 ( .A(p_input[718]), .B(n25231), .Z(n24912) );
  AND U25077 ( .A(n562), .B(n25232), .Z(n25231) );
  XOR U25078 ( .A(p_input[750]), .B(p_input[718]), .Z(n25232) );
  XNOR U25079 ( .A(n24909), .B(n25227), .Z(n25229) );
  XOR U25080 ( .A(n25233), .B(n25234), .Z(n24909) );
  AND U25081 ( .A(n560), .B(n25235), .Z(n25234) );
  XOR U25082 ( .A(p_input[686]), .B(p_input[654]), .Z(n25235) );
  XOR U25083 ( .A(n25236), .B(n25237), .Z(n25227) );
  AND U25084 ( .A(n25238), .B(n25239), .Z(n25237) );
  XOR U25085 ( .A(n25236), .B(n24924), .Z(n25239) );
  XNOR U25086 ( .A(p_input[717]), .B(n25240), .Z(n24924) );
  AND U25087 ( .A(n562), .B(n25241), .Z(n25240) );
  XOR U25088 ( .A(p_input[749]), .B(p_input[717]), .Z(n25241) );
  XNOR U25089 ( .A(n24921), .B(n25236), .Z(n25238) );
  XOR U25090 ( .A(n25242), .B(n25243), .Z(n24921) );
  AND U25091 ( .A(n560), .B(n25244), .Z(n25243) );
  XOR U25092 ( .A(p_input[685]), .B(p_input[653]), .Z(n25244) );
  XOR U25093 ( .A(n25245), .B(n25246), .Z(n25236) );
  AND U25094 ( .A(n25247), .B(n25248), .Z(n25246) );
  XOR U25095 ( .A(n25245), .B(n24936), .Z(n25248) );
  XNOR U25096 ( .A(p_input[716]), .B(n25249), .Z(n24936) );
  AND U25097 ( .A(n562), .B(n25250), .Z(n25249) );
  XOR U25098 ( .A(p_input[748]), .B(p_input[716]), .Z(n25250) );
  XNOR U25099 ( .A(n24933), .B(n25245), .Z(n25247) );
  XOR U25100 ( .A(n25251), .B(n25252), .Z(n24933) );
  AND U25101 ( .A(n560), .B(n25253), .Z(n25252) );
  XOR U25102 ( .A(p_input[684]), .B(p_input[652]), .Z(n25253) );
  XOR U25103 ( .A(n25254), .B(n25255), .Z(n25245) );
  AND U25104 ( .A(n25256), .B(n25257), .Z(n25255) );
  XOR U25105 ( .A(n25254), .B(n24948), .Z(n25257) );
  XNOR U25106 ( .A(p_input[715]), .B(n25258), .Z(n24948) );
  AND U25107 ( .A(n562), .B(n25259), .Z(n25258) );
  XOR U25108 ( .A(p_input[747]), .B(p_input[715]), .Z(n25259) );
  XNOR U25109 ( .A(n24945), .B(n25254), .Z(n25256) );
  XOR U25110 ( .A(n25260), .B(n25261), .Z(n24945) );
  AND U25111 ( .A(n560), .B(n25262), .Z(n25261) );
  XOR U25112 ( .A(p_input[683]), .B(p_input[651]), .Z(n25262) );
  XOR U25113 ( .A(n25263), .B(n25264), .Z(n25254) );
  AND U25114 ( .A(n25265), .B(n25266), .Z(n25264) );
  XOR U25115 ( .A(n25263), .B(n24960), .Z(n25266) );
  XNOR U25116 ( .A(p_input[714]), .B(n25267), .Z(n24960) );
  AND U25117 ( .A(n562), .B(n25268), .Z(n25267) );
  XOR U25118 ( .A(p_input[746]), .B(p_input[714]), .Z(n25268) );
  XNOR U25119 ( .A(n24957), .B(n25263), .Z(n25265) );
  XOR U25120 ( .A(n25269), .B(n25270), .Z(n24957) );
  AND U25121 ( .A(n560), .B(n25271), .Z(n25270) );
  XOR U25122 ( .A(p_input[682]), .B(p_input[650]), .Z(n25271) );
  XOR U25123 ( .A(n25272), .B(n25273), .Z(n25263) );
  AND U25124 ( .A(n25274), .B(n25275), .Z(n25273) );
  XOR U25125 ( .A(n25272), .B(n24972), .Z(n25275) );
  XNOR U25126 ( .A(p_input[713]), .B(n25276), .Z(n24972) );
  AND U25127 ( .A(n562), .B(n25277), .Z(n25276) );
  XOR U25128 ( .A(p_input[745]), .B(p_input[713]), .Z(n25277) );
  XNOR U25129 ( .A(n24969), .B(n25272), .Z(n25274) );
  XOR U25130 ( .A(n25278), .B(n25279), .Z(n24969) );
  AND U25131 ( .A(n560), .B(n25280), .Z(n25279) );
  XOR U25132 ( .A(p_input[681]), .B(p_input[649]), .Z(n25280) );
  XOR U25133 ( .A(n25281), .B(n25282), .Z(n25272) );
  AND U25134 ( .A(n25283), .B(n25284), .Z(n25282) );
  XOR U25135 ( .A(n25281), .B(n24984), .Z(n25284) );
  XNOR U25136 ( .A(p_input[712]), .B(n25285), .Z(n24984) );
  AND U25137 ( .A(n562), .B(n25286), .Z(n25285) );
  XOR U25138 ( .A(p_input[744]), .B(p_input[712]), .Z(n25286) );
  XNOR U25139 ( .A(n24981), .B(n25281), .Z(n25283) );
  XOR U25140 ( .A(n25287), .B(n25288), .Z(n24981) );
  AND U25141 ( .A(n560), .B(n25289), .Z(n25288) );
  XOR U25142 ( .A(p_input[680]), .B(p_input[648]), .Z(n25289) );
  XOR U25143 ( .A(n25290), .B(n25291), .Z(n25281) );
  AND U25144 ( .A(n25292), .B(n25293), .Z(n25291) );
  XOR U25145 ( .A(n25290), .B(n24996), .Z(n25293) );
  XNOR U25146 ( .A(p_input[711]), .B(n25294), .Z(n24996) );
  AND U25147 ( .A(n562), .B(n25295), .Z(n25294) );
  XOR U25148 ( .A(p_input[743]), .B(p_input[711]), .Z(n25295) );
  XNOR U25149 ( .A(n24993), .B(n25290), .Z(n25292) );
  XOR U25150 ( .A(n25296), .B(n25297), .Z(n24993) );
  AND U25151 ( .A(n560), .B(n25298), .Z(n25297) );
  XOR U25152 ( .A(p_input[679]), .B(p_input[647]), .Z(n25298) );
  XOR U25153 ( .A(n25299), .B(n25300), .Z(n25290) );
  AND U25154 ( .A(n25301), .B(n25302), .Z(n25300) );
  XOR U25155 ( .A(n25299), .B(n25008), .Z(n25302) );
  XNOR U25156 ( .A(p_input[710]), .B(n25303), .Z(n25008) );
  AND U25157 ( .A(n562), .B(n25304), .Z(n25303) );
  XOR U25158 ( .A(p_input[742]), .B(p_input[710]), .Z(n25304) );
  XNOR U25159 ( .A(n25005), .B(n25299), .Z(n25301) );
  XOR U25160 ( .A(n25305), .B(n25306), .Z(n25005) );
  AND U25161 ( .A(n560), .B(n25307), .Z(n25306) );
  XOR U25162 ( .A(p_input[678]), .B(p_input[646]), .Z(n25307) );
  XOR U25163 ( .A(n25308), .B(n25309), .Z(n25299) );
  AND U25164 ( .A(n25310), .B(n25311), .Z(n25309) );
  XOR U25165 ( .A(n25308), .B(n25020), .Z(n25311) );
  XNOR U25166 ( .A(p_input[709]), .B(n25312), .Z(n25020) );
  AND U25167 ( .A(n562), .B(n25313), .Z(n25312) );
  XOR U25168 ( .A(p_input[741]), .B(p_input[709]), .Z(n25313) );
  XNOR U25169 ( .A(n25017), .B(n25308), .Z(n25310) );
  XOR U25170 ( .A(n25314), .B(n25315), .Z(n25017) );
  AND U25171 ( .A(n560), .B(n25316), .Z(n25315) );
  XOR U25172 ( .A(p_input[677]), .B(p_input[645]), .Z(n25316) );
  XOR U25173 ( .A(n25317), .B(n25318), .Z(n25308) );
  AND U25174 ( .A(n25319), .B(n25320), .Z(n25318) );
  XOR U25175 ( .A(n25317), .B(n25032), .Z(n25320) );
  XNOR U25176 ( .A(p_input[708]), .B(n25321), .Z(n25032) );
  AND U25177 ( .A(n562), .B(n25322), .Z(n25321) );
  XOR U25178 ( .A(p_input[740]), .B(p_input[708]), .Z(n25322) );
  XNOR U25179 ( .A(n25029), .B(n25317), .Z(n25319) );
  XOR U25180 ( .A(n25323), .B(n25324), .Z(n25029) );
  AND U25181 ( .A(n560), .B(n25325), .Z(n25324) );
  XOR U25182 ( .A(p_input[676]), .B(p_input[644]), .Z(n25325) );
  XOR U25183 ( .A(n25326), .B(n25327), .Z(n25317) );
  AND U25184 ( .A(n25328), .B(n25329), .Z(n25327) );
  XOR U25185 ( .A(n25326), .B(n25044), .Z(n25329) );
  XNOR U25186 ( .A(p_input[707]), .B(n25330), .Z(n25044) );
  AND U25187 ( .A(n562), .B(n25331), .Z(n25330) );
  XOR U25188 ( .A(p_input[739]), .B(p_input[707]), .Z(n25331) );
  XNOR U25189 ( .A(n25041), .B(n25326), .Z(n25328) );
  XOR U25190 ( .A(n25332), .B(n25333), .Z(n25041) );
  AND U25191 ( .A(n560), .B(n25334), .Z(n25333) );
  XOR U25192 ( .A(p_input[675]), .B(p_input[643]), .Z(n25334) );
  XOR U25193 ( .A(n25335), .B(n25336), .Z(n25326) );
  AND U25194 ( .A(n25337), .B(n25338), .Z(n25336) );
  XOR U25195 ( .A(n25056), .B(n25335), .Z(n25338) );
  XNOR U25196 ( .A(p_input[706]), .B(n25339), .Z(n25056) );
  AND U25197 ( .A(n562), .B(n25340), .Z(n25339) );
  XOR U25198 ( .A(p_input[738]), .B(p_input[706]), .Z(n25340) );
  XNOR U25199 ( .A(n25335), .B(n25053), .Z(n25337) );
  XOR U25200 ( .A(n25341), .B(n25342), .Z(n25053) );
  AND U25201 ( .A(n560), .B(n25343), .Z(n25342) );
  XOR U25202 ( .A(p_input[674]), .B(p_input[642]), .Z(n25343) );
  XOR U25203 ( .A(n25344), .B(n25345), .Z(n25335) );
  AND U25204 ( .A(n25346), .B(n25347), .Z(n25345) );
  XNOR U25205 ( .A(n25348), .B(n25069), .Z(n25347) );
  XNOR U25206 ( .A(p_input[705]), .B(n25349), .Z(n25069) );
  AND U25207 ( .A(n562), .B(n25350), .Z(n25349) );
  XNOR U25208 ( .A(p_input[737]), .B(n25351), .Z(n25350) );
  IV U25209 ( .A(p_input[705]), .Z(n25351) );
  XNOR U25210 ( .A(n25066), .B(n25344), .Z(n25346) );
  XNOR U25211 ( .A(p_input[641]), .B(n25352), .Z(n25066) );
  AND U25212 ( .A(n560), .B(n25353), .Z(n25352) );
  XOR U25213 ( .A(p_input[673]), .B(p_input[641]), .Z(n25353) );
  IV U25214 ( .A(n25348), .Z(n25344) );
  AND U25215 ( .A(n25074), .B(n25077), .Z(n25348) );
  XOR U25216 ( .A(p_input[704]), .B(n25354), .Z(n25077) );
  AND U25217 ( .A(n562), .B(n25355), .Z(n25354) );
  XOR U25218 ( .A(p_input[736]), .B(p_input[704]), .Z(n25355) );
  XOR U25219 ( .A(n25356), .B(n25357), .Z(n562) );
  AND U25220 ( .A(n25358), .B(n25359), .Z(n25357) );
  XNOR U25221 ( .A(p_input[767]), .B(n25356), .Z(n25359) );
  XOR U25222 ( .A(n25356), .B(p_input[735]), .Z(n25358) );
  XOR U25223 ( .A(n25360), .B(n25361), .Z(n25356) );
  AND U25224 ( .A(n25362), .B(n25363), .Z(n25361) );
  XNOR U25225 ( .A(p_input[766]), .B(n25360), .Z(n25363) );
  XOR U25226 ( .A(n25360), .B(p_input[734]), .Z(n25362) );
  XOR U25227 ( .A(n25364), .B(n25365), .Z(n25360) );
  AND U25228 ( .A(n25366), .B(n25367), .Z(n25365) );
  XNOR U25229 ( .A(p_input[765]), .B(n25364), .Z(n25367) );
  XOR U25230 ( .A(n25364), .B(p_input[733]), .Z(n25366) );
  XOR U25231 ( .A(n25368), .B(n25369), .Z(n25364) );
  AND U25232 ( .A(n25370), .B(n25371), .Z(n25369) );
  XNOR U25233 ( .A(p_input[764]), .B(n25368), .Z(n25371) );
  XOR U25234 ( .A(n25368), .B(p_input[732]), .Z(n25370) );
  XOR U25235 ( .A(n25372), .B(n25373), .Z(n25368) );
  AND U25236 ( .A(n25374), .B(n25375), .Z(n25373) );
  XNOR U25237 ( .A(p_input[763]), .B(n25372), .Z(n25375) );
  XOR U25238 ( .A(n25372), .B(p_input[731]), .Z(n25374) );
  XOR U25239 ( .A(n25376), .B(n25377), .Z(n25372) );
  AND U25240 ( .A(n25378), .B(n25379), .Z(n25377) );
  XNOR U25241 ( .A(p_input[762]), .B(n25376), .Z(n25379) );
  XOR U25242 ( .A(n25376), .B(p_input[730]), .Z(n25378) );
  XOR U25243 ( .A(n25380), .B(n25381), .Z(n25376) );
  AND U25244 ( .A(n25382), .B(n25383), .Z(n25381) );
  XNOR U25245 ( .A(p_input[761]), .B(n25380), .Z(n25383) );
  XOR U25246 ( .A(n25380), .B(p_input[729]), .Z(n25382) );
  XOR U25247 ( .A(n25384), .B(n25385), .Z(n25380) );
  AND U25248 ( .A(n25386), .B(n25387), .Z(n25385) );
  XNOR U25249 ( .A(p_input[760]), .B(n25384), .Z(n25387) );
  XOR U25250 ( .A(n25384), .B(p_input[728]), .Z(n25386) );
  XOR U25251 ( .A(n25388), .B(n25389), .Z(n25384) );
  AND U25252 ( .A(n25390), .B(n25391), .Z(n25389) );
  XNOR U25253 ( .A(p_input[759]), .B(n25388), .Z(n25391) );
  XOR U25254 ( .A(n25388), .B(p_input[727]), .Z(n25390) );
  XOR U25255 ( .A(n25392), .B(n25393), .Z(n25388) );
  AND U25256 ( .A(n25394), .B(n25395), .Z(n25393) );
  XNOR U25257 ( .A(p_input[758]), .B(n25392), .Z(n25395) );
  XOR U25258 ( .A(n25392), .B(p_input[726]), .Z(n25394) );
  XOR U25259 ( .A(n25396), .B(n25397), .Z(n25392) );
  AND U25260 ( .A(n25398), .B(n25399), .Z(n25397) );
  XNOR U25261 ( .A(p_input[757]), .B(n25396), .Z(n25399) );
  XOR U25262 ( .A(n25396), .B(p_input[725]), .Z(n25398) );
  XOR U25263 ( .A(n25400), .B(n25401), .Z(n25396) );
  AND U25264 ( .A(n25402), .B(n25403), .Z(n25401) );
  XNOR U25265 ( .A(p_input[756]), .B(n25400), .Z(n25403) );
  XOR U25266 ( .A(n25400), .B(p_input[724]), .Z(n25402) );
  XOR U25267 ( .A(n25404), .B(n25405), .Z(n25400) );
  AND U25268 ( .A(n25406), .B(n25407), .Z(n25405) );
  XNOR U25269 ( .A(p_input[755]), .B(n25404), .Z(n25407) );
  XOR U25270 ( .A(n25404), .B(p_input[723]), .Z(n25406) );
  XOR U25271 ( .A(n25408), .B(n25409), .Z(n25404) );
  AND U25272 ( .A(n25410), .B(n25411), .Z(n25409) );
  XNOR U25273 ( .A(p_input[754]), .B(n25408), .Z(n25411) );
  XOR U25274 ( .A(n25408), .B(p_input[722]), .Z(n25410) );
  XOR U25275 ( .A(n25412), .B(n25413), .Z(n25408) );
  AND U25276 ( .A(n25414), .B(n25415), .Z(n25413) );
  XNOR U25277 ( .A(p_input[753]), .B(n25412), .Z(n25415) );
  XOR U25278 ( .A(n25412), .B(p_input[721]), .Z(n25414) );
  XOR U25279 ( .A(n25416), .B(n25417), .Z(n25412) );
  AND U25280 ( .A(n25418), .B(n25419), .Z(n25417) );
  XNOR U25281 ( .A(p_input[752]), .B(n25416), .Z(n25419) );
  XOR U25282 ( .A(n25416), .B(p_input[720]), .Z(n25418) );
  XOR U25283 ( .A(n25420), .B(n25421), .Z(n25416) );
  AND U25284 ( .A(n25422), .B(n25423), .Z(n25421) );
  XNOR U25285 ( .A(p_input[751]), .B(n25420), .Z(n25423) );
  XOR U25286 ( .A(n25420), .B(p_input[719]), .Z(n25422) );
  XOR U25287 ( .A(n25424), .B(n25425), .Z(n25420) );
  AND U25288 ( .A(n25426), .B(n25427), .Z(n25425) );
  XNOR U25289 ( .A(p_input[750]), .B(n25424), .Z(n25427) );
  XOR U25290 ( .A(n25424), .B(p_input[718]), .Z(n25426) );
  XOR U25291 ( .A(n25428), .B(n25429), .Z(n25424) );
  AND U25292 ( .A(n25430), .B(n25431), .Z(n25429) );
  XNOR U25293 ( .A(p_input[749]), .B(n25428), .Z(n25431) );
  XOR U25294 ( .A(n25428), .B(p_input[717]), .Z(n25430) );
  XOR U25295 ( .A(n25432), .B(n25433), .Z(n25428) );
  AND U25296 ( .A(n25434), .B(n25435), .Z(n25433) );
  XNOR U25297 ( .A(p_input[748]), .B(n25432), .Z(n25435) );
  XOR U25298 ( .A(n25432), .B(p_input[716]), .Z(n25434) );
  XOR U25299 ( .A(n25436), .B(n25437), .Z(n25432) );
  AND U25300 ( .A(n25438), .B(n25439), .Z(n25437) );
  XNOR U25301 ( .A(p_input[747]), .B(n25436), .Z(n25439) );
  XOR U25302 ( .A(n25436), .B(p_input[715]), .Z(n25438) );
  XOR U25303 ( .A(n25440), .B(n25441), .Z(n25436) );
  AND U25304 ( .A(n25442), .B(n25443), .Z(n25441) );
  XNOR U25305 ( .A(p_input[746]), .B(n25440), .Z(n25443) );
  XOR U25306 ( .A(n25440), .B(p_input[714]), .Z(n25442) );
  XOR U25307 ( .A(n25444), .B(n25445), .Z(n25440) );
  AND U25308 ( .A(n25446), .B(n25447), .Z(n25445) );
  XNOR U25309 ( .A(p_input[745]), .B(n25444), .Z(n25447) );
  XOR U25310 ( .A(n25444), .B(p_input[713]), .Z(n25446) );
  XOR U25311 ( .A(n25448), .B(n25449), .Z(n25444) );
  AND U25312 ( .A(n25450), .B(n25451), .Z(n25449) );
  XNOR U25313 ( .A(p_input[744]), .B(n25448), .Z(n25451) );
  XOR U25314 ( .A(n25448), .B(p_input[712]), .Z(n25450) );
  XOR U25315 ( .A(n25452), .B(n25453), .Z(n25448) );
  AND U25316 ( .A(n25454), .B(n25455), .Z(n25453) );
  XNOR U25317 ( .A(p_input[743]), .B(n25452), .Z(n25455) );
  XOR U25318 ( .A(n25452), .B(p_input[711]), .Z(n25454) );
  XOR U25319 ( .A(n25456), .B(n25457), .Z(n25452) );
  AND U25320 ( .A(n25458), .B(n25459), .Z(n25457) );
  XNOR U25321 ( .A(p_input[742]), .B(n25456), .Z(n25459) );
  XOR U25322 ( .A(n25456), .B(p_input[710]), .Z(n25458) );
  XOR U25323 ( .A(n25460), .B(n25461), .Z(n25456) );
  AND U25324 ( .A(n25462), .B(n25463), .Z(n25461) );
  XNOR U25325 ( .A(p_input[741]), .B(n25460), .Z(n25463) );
  XOR U25326 ( .A(n25460), .B(p_input[709]), .Z(n25462) );
  XOR U25327 ( .A(n25464), .B(n25465), .Z(n25460) );
  AND U25328 ( .A(n25466), .B(n25467), .Z(n25465) );
  XNOR U25329 ( .A(p_input[740]), .B(n25464), .Z(n25467) );
  XOR U25330 ( .A(n25464), .B(p_input[708]), .Z(n25466) );
  XOR U25331 ( .A(n25468), .B(n25469), .Z(n25464) );
  AND U25332 ( .A(n25470), .B(n25471), .Z(n25469) );
  XNOR U25333 ( .A(p_input[739]), .B(n25468), .Z(n25471) );
  XOR U25334 ( .A(n25468), .B(p_input[707]), .Z(n25470) );
  XOR U25335 ( .A(n25472), .B(n25473), .Z(n25468) );
  AND U25336 ( .A(n25474), .B(n25475), .Z(n25473) );
  XNOR U25337 ( .A(p_input[738]), .B(n25472), .Z(n25475) );
  XOR U25338 ( .A(n25472), .B(p_input[706]), .Z(n25474) );
  XNOR U25339 ( .A(n25476), .B(n25477), .Z(n25472) );
  AND U25340 ( .A(n25478), .B(n25479), .Z(n25477) );
  XOR U25341 ( .A(p_input[737]), .B(n25476), .Z(n25479) );
  XNOR U25342 ( .A(p_input[705]), .B(n25476), .Z(n25478) );
  AND U25343 ( .A(p_input[736]), .B(n25480), .Z(n25476) );
  IV U25344 ( .A(p_input[704]), .Z(n25480) );
  XNOR U25345 ( .A(p_input[640]), .B(n25481), .Z(n25074) );
  AND U25346 ( .A(n560), .B(n25482), .Z(n25481) );
  XOR U25347 ( .A(p_input[672]), .B(p_input[640]), .Z(n25482) );
  XOR U25348 ( .A(n25483), .B(n25484), .Z(n560) );
  AND U25349 ( .A(n25485), .B(n25486), .Z(n25484) );
  XNOR U25350 ( .A(p_input[703]), .B(n25483), .Z(n25486) );
  XOR U25351 ( .A(n25483), .B(p_input[671]), .Z(n25485) );
  XOR U25352 ( .A(n25487), .B(n25488), .Z(n25483) );
  AND U25353 ( .A(n25489), .B(n25490), .Z(n25488) );
  XNOR U25354 ( .A(p_input[702]), .B(n25487), .Z(n25490) );
  XNOR U25355 ( .A(n25487), .B(n25089), .Z(n25489) );
  IV U25356 ( .A(p_input[670]), .Z(n25089) );
  XOR U25357 ( .A(n25491), .B(n25492), .Z(n25487) );
  AND U25358 ( .A(n25493), .B(n25494), .Z(n25492) );
  XNOR U25359 ( .A(p_input[701]), .B(n25491), .Z(n25494) );
  XNOR U25360 ( .A(n25491), .B(n25098), .Z(n25493) );
  IV U25361 ( .A(p_input[669]), .Z(n25098) );
  XOR U25362 ( .A(n25495), .B(n25496), .Z(n25491) );
  AND U25363 ( .A(n25497), .B(n25498), .Z(n25496) );
  XNOR U25364 ( .A(p_input[700]), .B(n25495), .Z(n25498) );
  XNOR U25365 ( .A(n25495), .B(n25107), .Z(n25497) );
  IV U25366 ( .A(p_input[668]), .Z(n25107) );
  XOR U25367 ( .A(n25499), .B(n25500), .Z(n25495) );
  AND U25368 ( .A(n25501), .B(n25502), .Z(n25500) );
  XNOR U25369 ( .A(p_input[699]), .B(n25499), .Z(n25502) );
  XNOR U25370 ( .A(n25499), .B(n25116), .Z(n25501) );
  IV U25371 ( .A(p_input[667]), .Z(n25116) );
  XOR U25372 ( .A(n25503), .B(n25504), .Z(n25499) );
  AND U25373 ( .A(n25505), .B(n25506), .Z(n25504) );
  XNOR U25374 ( .A(p_input[698]), .B(n25503), .Z(n25506) );
  XNOR U25375 ( .A(n25503), .B(n25125), .Z(n25505) );
  IV U25376 ( .A(p_input[666]), .Z(n25125) );
  XOR U25377 ( .A(n25507), .B(n25508), .Z(n25503) );
  AND U25378 ( .A(n25509), .B(n25510), .Z(n25508) );
  XNOR U25379 ( .A(p_input[697]), .B(n25507), .Z(n25510) );
  XNOR U25380 ( .A(n25507), .B(n25134), .Z(n25509) );
  IV U25381 ( .A(p_input[665]), .Z(n25134) );
  XOR U25382 ( .A(n25511), .B(n25512), .Z(n25507) );
  AND U25383 ( .A(n25513), .B(n25514), .Z(n25512) );
  XNOR U25384 ( .A(p_input[696]), .B(n25511), .Z(n25514) );
  XNOR U25385 ( .A(n25511), .B(n25143), .Z(n25513) );
  IV U25386 ( .A(p_input[664]), .Z(n25143) );
  XOR U25387 ( .A(n25515), .B(n25516), .Z(n25511) );
  AND U25388 ( .A(n25517), .B(n25518), .Z(n25516) );
  XNOR U25389 ( .A(p_input[695]), .B(n25515), .Z(n25518) );
  XNOR U25390 ( .A(n25515), .B(n25152), .Z(n25517) );
  IV U25391 ( .A(p_input[663]), .Z(n25152) );
  XOR U25392 ( .A(n25519), .B(n25520), .Z(n25515) );
  AND U25393 ( .A(n25521), .B(n25522), .Z(n25520) );
  XNOR U25394 ( .A(p_input[694]), .B(n25519), .Z(n25522) );
  XNOR U25395 ( .A(n25519), .B(n25161), .Z(n25521) );
  IV U25396 ( .A(p_input[662]), .Z(n25161) );
  XOR U25397 ( .A(n25523), .B(n25524), .Z(n25519) );
  AND U25398 ( .A(n25525), .B(n25526), .Z(n25524) );
  XNOR U25399 ( .A(p_input[693]), .B(n25523), .Z(n25526) );
  XNOR U25400 ( .A(n25523), .B(n25170), .Z(n25525) );
  IV U25401 ( .A(p_input[661]), .Z(n25170) );
  XOR U25402 ( .A(n25527), .B(n25528), .Z(n25523) );
  AND U25403 ( .A(n25529), .B(n25530), .Z(n25528) );
  XNOR U25404 ( .A(p_input[692]), .B(n25527), .Z(n25530) );
  XNOR U25405 ( .A(n25527), .B(n25179), .Z(n25529) );
  IV U25406 ( .A(p_input[660]), .Z(n25179) );
  XOR U25407 ( .A(n25531), .B(n25532), .Z(n25527) );
  AND U25408 ( .A(n25533), .B(n25534), .Z(n25532) );
  XNOR U25409 ( .A(p_input[691]), .B(n25531), .Z(n25534) );
  XNOR U25410 ( .A(n25531), .B(n25188), .Z(n25533) );
  IV U25411 ( .A(p_input[659]), .Z(n25188) );
  XOR U25412 ( .A(n25535), .B(n25536), .Z(n25531) );
  AND U25413 ( .A(n25537), .B(n25538), .Z(n25536) );
  XNOR U25414 ( .A(p_input[690]), .B(n25535), .Z(n25538) );
  XNOR U25415 ( .A(n25535), .B(n25197), .Z(n25537) );
  IV U25416 ( .A(p_input[658]), .Z(n25197) );
  XOR U25417 ( .A(n25539), .B(n25540), .Z(n25535) );
  AND U25418 ( .A(n25541), .B(n25542), .Z(n25540) );
  XNOR U25419 ( .A(p_input[689]), .B(n25539), .Z(n25542) );
  XNOR U25420 ( .A(n25539), .B(n25206), .Z(n25541) );
  IV U25421 ( .A(p_input[657]), .Z(n25206) );
  XOR U25422 ( .A(n25543), .B(n25544), .Z(n25539) );
  AND U25423 ( .A(n25545), .B(n25546), .Z(n25544) );
  XNOR U25424 ( .A(p_input[688]), .B(n25543), .Z(n25546) );
  XNOR U25425 ( .A(n25543), .B(n25215), .Z(n25545) );
  IV U25426 ( .A(p_input[656]), .Z(n25215) );
  XOR U25427 ( .A(n25547), .B(n25548), .Z(n25543) );
  AND U25428 ( .A(n25549), .B(n25550), .Z(n25548) );
  XNOR U25429 ( .A(p_input[687]), .B(n25547), .Z(n25550) );
  XNOR U25430 ( .A(n25547), .B(n25224), .Z(n25549) );
  IV U25431 ( .A(p_input[655]), .Z(n25224) );
  XOR U25432 ( .A(n25551), .B(n25552), .Z(n25547) );
  AND U25433 ( .A(n25553), .B(n25554), .Z(n25552) );
  XNOR U25434 ( .A(p_input[686]), .B(n25551), .Z(n25554) );
  XNOR U25435 ( .A(n25551), .B(n25233), .Z(n25553) );
  IV U25436 ( .A(p_input[654]), .Z(n25233) );
  XOR U25437 ( .A(n25555), .B(n25556), .Z(n25551) );
  AND U25438 ( .A(n25557), .B(n25558), .Z(n25556) );
  XNOR U25439 ( .A(p_input[685]), .B(n25555), .Z(n25558) );
  XNOR U25440 ( .A(n25555), .B(n25242), .Z(n25557) );
  IV U25441 ( .A(p_input[653]), .Z(n25242) );
  XOR U25442 ( .A(n25559), .B(n25560), .Z(n25555) );
  AND U25443 ( .A(n25561), .B(n25562), .Z(n25560) );
  XNOR U25444 ( .A(p_input[684]), .B(n25559), .Z(n25562) );
  XNOR U25445 ( .A(n25559), .B(n25251), .Z(n25561) );
  IV U25446 ( .A(p_input[652]), .Z(n25251) );
  XOR U25447 ( .A(n25563), .B(n25564), .Z(n25559) );
  AND U25448 ( .A(n25565), .B(n25566), .Z(n25564) );
  XNOR U25449 ( .A(p_input[683]), .B(n25563), .Z(n25566) );
  XNOR U25450 ( .A(n25563), .B(n25260), .Z(n25565) );
  IV U25451 ( .A(p_input[651]), .Z(n25260) );
  XOR U25452 ( .A(n25567), .B(n25568), .Z(n25563) );
  AND U25453 ( .A(n25569), .B(n25570), .Z(n25568) );
  XNOR U25454 ( .A(p_input[682]), .B(n25567), .Z(n25570) );
  XNOR U25455 ( .A(n25567), .B(n25269), .Z(n25569) );
  IV U25456 ( .A(p_input[650]), .Z(n25269) );
  XOR U25457 ( .A(n25571), .B(n25572), .Z(n25567) );
  AND U25458 ( .A(n25573), .B(n25574), .Z(n25572) );
  XNOR U25459 ( .A(p_input[681]), .B(n25571), .Z(n25574) );
  XNOR U25460 ( .A(n25571), .B(n25278), .Z(n25573) );
  IV U25461 ( .A(p_input[649]), .Z(n25278) );
  XOR U25462 ( .A(n25575), .B(n25576), .Z(n25571) );
  AND U25463 ( .A(n25577), .B(n25578), .Z(n25576) );
  XNOR U25464 ( .A(p_input[680]), .B(n25575), .Z(n25578) );
  XNOR U25465 ( .A(n25575), .B(n25287), .Z(n25577) );
  IV U25466 ( .A(p_input[648]), .Z(n25287) );
  XOR U25467 ( .A(n25579), .B(n25580), .Z(n25575) );
  AND U25468 ( .A(n25581), .B(n25582), .Z(n25580) );
  XNOR U25469 ( .A(p_input[679]), .B(n25579), .Z(n25582) );
  XNOR U25470 ( .A(n25579), .B(n25296), .Z(n25581) );
  IV U25471 ( .A(p_input[647]), .Z(n25296) );
  XOR U25472 ( .A(n25583), .B(n25584), .Z(n25579) );
  AND U25473 ( .A(n25585), .B(n25586), .Z(n25584) );
  XNOR U25474 ( .A(p_input[678]), .B(n25583), .Z(n25586) );
  XNOR U25475 ( .A(n25583), .B(n25305), .Z(n25585) );
  IV U25476 ( .A(p_input[646]), .Z(n25305) );
  XOR U25477 ( .A(n25587), .B(n25588), .Z(n25583) );
  AND U25478 ( .A(n25589), .B(n25590), .Z(n25588) );
  XNOR U25479 ( .A(p_input[677]), .B(n25587), .Z(n25590) );
  XNOR U25480 ( .A(n25587), .B(n25314), .Z(n25589) );
  IV U25481 ( .A(p_input[645]), .Z(n25314) );
  XOR U25482 ( .A(n25591), .B(n25592), .Z(n25587) );
  AND U25483 ( .A(n25593), .B(n25594), .Z(n25592) );
  XNOR U25484 ( .A(p_input[676]), .B(n25591), .Z(n25594) );
  XNOR U25485 ( .A(n25591), .B(n25323), .Z(n25593) );
  IV U25486 ( .A(p_input[644]), .Z(n25323) );
  XOR U25487 ( .A(n25595), .B(n25596), .Z(n25591) );
  AND U25488 ( .A(n25597), .B(n25598), .Z(n25596) );
  XNOR U25489 ( .A(p_input[675]), .B(n25595), .Z(n25598) );
  XNOR U25490 ( .A(n25595), .B(n25332), .Z(n25597) );
  IV U25491 ( .A(p_input[643]), .Z(n25332) );
  XOR U25492 ( .A(n25599), .B(n25600), .Z(n25595) );
  AND U25493 ( .A(n25601), .B(n25602), .Z(n25600) );
  XNOR U25494 ( .A(p_input[674]), .B(n25599), .Z(n25602) );
  XNOR U25495 ( .A(n25599), .B(n25341), .Z(n25601) );
  IV U25496 ( .A(p_input[642]), .Z(n25341) );
  XNOR U25497 ( .A(n25603), .B(n25604), .Z(n25599) );
  AND U25498 ( .A(n25605), .B(n25606), .Z(n25604) );
  XOR U25499 ( .A(p_input[673]), .B(n25603), .Z(n25606) );
  XNOR U25500 ( .A(p_input[641]), .B(n25603), .Z(n25605) );
  AND U25501 ( .A(p_input[672]), .B(n25607), .Z(n25603) );
  IV U25502 ( .A(p_input[640]), .Z(n25607) );
  XOR U25503 ( .A(n25608), .B(n25609), .Z(n24697) );
  AND U25504 ( .A(n395), .B(n25610), .Z(n25609) );
  XNOR U25505 ( .A(n25611), .B(n25608), .Z(n25610) );
  XOR U25506 ( .A(n25612), .B(n25613), .Z(n395) );
  AND U25507 ( .A(n25614), .B(n25615), .Z(n25613) );
  XNOR U25508 ( .A(n24712), .B(n25612), .Z(n25615) );
  AND U25509 ( .A(p_input[639]), .B(p_input[607]), .Z(n24712) );
  XNOR U25510 ( .A(n25612), .B(n24709), .Z(n25614) );
  IV U25511 ( .A(n25616), .Z(n24709) );
  AND U25512 ( .A(p_input[543]), .B(p_input[575]), .Z(n25616) );
  XOR U25513 ( .A(n25617), .B(n25618), .Z(n25612) );
  AND U25514 ( .A(n25619), .B(n25620), .Z(n25618) );
  XOR U25515 ( .A(n25617), .B(n24724), .Z(n25620) );
  XNOR U25516 ( .A(p_input[606]), .B(n25621), .Z(n24724) );
  AND U25517 ( .A(n566), .B(n25622), .Z(n25621) );
  XOR U25518 ( .A(p_input[638]), .B(p_input[606]), .Z(n25622) );
  XNOR U25519 ( .A(n24721), .B(n25617), .Z(n25619) );
  XOR U25520 ( .A(n25623), .B(n25624), .Z(n24721) );
  AND U25521 ( .A(n563), .B(n25625), .Z(n25624) );
  XOR U25522 ( .A(p_input[574]), .B(p_input[542]), .Z(n25625) );
  XOR U25523 ( .A(n25626), .B(n25627), .Z(n25617) );
  AND U25524 ( .A(n25628), .B(n25629), .Z(n25627) );
  XOR U25525 ( .A(n25626), .B(n24736), .Z(n25629) );
  XNOR U25526 ( .A(p_input[605]), .B(n25630), .Z(n24736) );
  AND U25527 ( .A(n566), .B(n25631), .Z(n25630) );
  XOR U25528 ( .A(p_input[637]), .B(p_input[605]), .Z(n25631) );
  XNOR U25529 ( .A(n24733), .B(n25626), .Z(n25628) );
  XOR U25530 ( .A(n25632), .B(n25633), .Z(n24733) );
  AND U25531 ( .A(n563), .B(n25634), .Z(n25633) );
  XOR U25532 ( .A(p_input[573]), .B(p_input[541]), .Z(n25634) );
  XOR U25533 ( .A(n25635), .B(n25636), .Z(n25626) );
  AND U25534 ( .A(n25637), .B(n25638), .Z(n25636) );
  XOR U25535 ( .A(n25635), .B(n24748), .Z(n25638) );
  XNOR U25536 ( .A(p_input[604]), .B(n25639), .Z(n24748) );
  AND U25537 ( .A(n566), .B(n25640), .Z(n25639) );
  XOR U25538 ( .A(p_input[636]), .B(p_input[604]), .Z(n25640) );
  XNOR U25539 ( .A(n24745), .B(n25635), .Z(n25637) );
  XOR U25540 ( .A(n25641), .B(n25642), .Z(n24745) );
  AND U25541 ( .A(n563), .B(n25643), .Z(n25642) );
  XOR U25542 ( .A(p_input[572]), .B(p_input[540]), .Z(n25643) );
  XOR U25543 ( .A(n25644), .B(n25645), .Z(n25635) );
  AND U25544 ( .A(n25646), .B(n25647), .Z(n25645) );
  XOR U25545 ( .A(n25644), .B(n24760), .Z(n25647) );
  XNOR U25546 ( .A(p_input[603]), .B(n25648), .Z(n24760) );
  AND U25547 ( .A(n566), .B(n25649), .Z(n25648) );
  XOR U25548 ( .A(p_input[635]), .B(p_input[603]), .Z(n25649) );
  XNOR U25549 ( .A(n24757), .B(n25644), .Z(n25646) );
  XOR U25550 ( .A(n25650), .B(n25651), .Z(n24757) );
  AND U25551 ( .A(n563), .B(n25652), .Z(n25651) );
  XOR U25552 ( .A(p_input[571]), .B(p_input[539]), .Z(n25652) );
  XOR U25553 ( .A(n25653), .B(n25654), .Z(n25644) );
  AND U25554 ( .A(n25655), .B(n25656), .Z(n25654) );
  XOR U25555 ( .A(n25653), .B(n24772), .Z(n25656) );
  XNOR U25556 ( .A(p_input[602]), .B(n25657), .Z(n24772) );
  AND U25557 ( .A(n566), .B(n25658), .Z(n25657) );
  XOR U25558 ( .A(p_input[634]), .B(p_input[602]), .Z(n25658) );
  XNOR U25559 ( .A(n24769), .B(n25653), .Z(n25655) );
  XOR U25560 ( .A(n25659), .B(n25660), .Z(n24769) );
  AND U25561 ( .A(n563), .B(n25661), .Z(n25660) );
  XOR U25562 ( .A(p_input[570]), .B(p_input[538]), .Z(n25661) );
  XOR U25563 ( .A(n25662), .B(n25663), .Z(n25653) );
  AND U25564 ( .A(n25664), .B(n25665), .Z(n25663) );
  XOR U25565 ( .A(n25662), .B(n24784), .Z(n25665) );
  XNOR U25566 ( .A(p_input[601]), .B(n25666), .Z(n24784) );
  AND U25567 ( .A(n566), .B(n25667), .Z(n25666) );
  XOR U25568 ( .A(p_input[633]), .B(p_input[601]), .Z(n25667) );
  XNOR U25569 ( .A(n24781), .B(n25662), .Z(n25664) );
  XOR U25570 ( .A(n25668), .B(n25669), .Z(n24781) );
  AND U25571 ( .A(n563), .B(n25670), .Z(n25669) );
  XOR U25572 ( .A(p_input[569]), .B(p_input[537]), .Z(n25670) );
  XOR U25573 ( .A(n25671), .B(n25672), .Z(n25662) );
  AND U25574 ( .A(n25673), .B(n25674), .Z(n25672) );
  XOR U25575 ( .A(n25671), .B(n24796), .Z(n25674) );
  XNOR U25576 ( .A(p_input[600]), .B(n25675), .Z(n24796) );
  AND U25577 ( .A(n566), .B(n25676), .Z(n25675) );
  XOR U25578 ( .A(p_input[632]), .B(p_input[600]), .Z(n25676) );
  XNOR U25579 ( .A(n24793), .B(n25671), .Z(n25673) );
  XOR U25580 ( .A(n25677), .B(n25678), .Z(n24793) );
  AND U25581 ( .A(n563), .B(n25679), .Z(n25678) );
  XOR U25582 ( .A(p_input[568]), .B(p_input[536]), .Z(n25679) );
  XOR U25583 ( .A(n25680), .B(n25681), .Z(n25671) );
  AND U25584 ( .A(n25682), .B(n25683), .Z(n25681) );
  XOR U25585 ( .A(n25680), .B(n24808), .Z(n25683) );
  XNOR U25586 ( .A(p_input[599]), .B(n25684), .Z(n24808) );
  AND U25587 ( .A(n566), .B(n25685), .Z(n25684) );
  XOR U25588 ( .A(p_input[631]), .B(p_input[599]), .Z(n25685) );
  XNOR U25589 ( .A(n24805), .B(n25680), .Z(n25682) );
  XOR U25590 ( .A(n25686), .B(n25687), .Z(n24805) );
  AND U25591 ( .A(n563), .B(n25688), .Z(n25687) );
  XOR U25592 ( .A(p_input[567]), .B(p_input[535]), .Z(n25688) );
  XOR U25593 ( .A(n25689), .B(n25690), .Z(n25680) );
  AND U25594 ( .A(n25691), .B(n25692), .Z(n25690) );
  XOR U25595 ( .A(n25689), .B(n24820), .Z(n25692) );
  XNOR U25596 ( .A(p_input[598]), .B(n25693), .Z(n24820) );
  AND U25597 ( .A(n566), .B(n25694), .Z(n25693) );
  XOR U25598 ( .A(p_input[630]), .B(p_input[598]), .Z(n25694) );
  XNOR U25599 ( .A(n24817), .B(n25689), .Z(n25691) );
  XOR U25600 ( .A(n25695), .B(n25696), .Z(n24817) );
  AND U25601 ( .A(n563), .B(n25697), .Z(n25696) );
  XOR U25602 ( .A(p_input[566]), .B(p_input[534]), .Z(n25697) );
  XOR U25603 ( .A(n25698), .B(n25699), .Z(n25689) );
  AND U25604 ( .A(n25700), .B(n25701), .Z(n25699) );
  XOR U25605 ( .A(n25698), .B(n24832), .Z(n25701) );
  XNOR U25606 ( .A(p_input[597]), .B(n25702), .Z(n24832) );
  AND U25607 ( .A(n566), .B(n25703), .Z(n25702) );
  XOR U25608 ( .A(p_input[629]), .B(p_input[597]), .Z(n25703) );
  XNOR U25609 ( .A(n24829), .B(n25698), .Z(n25700) );
  XOR U25610 ( .A(n25704), .B(n25705), .Z(n24829) );
  AND U25611 ( .A(n563), .B(n25706), .Z(n25705) );
  XOR U25612 ( .A(p_input[565]), .B(p_input[533]), .Z(n25706) );
  XOR U25613 ( .A(n25707), .B(n25708), .Z(n25698) );
  AND U25614 ( .A(n25709), .B(n25710), .Z(n25708) );
  XOR U25615 ( .A(n25707), .B(n24844), .Z(n25710) );
  XNOR U25616 ( .A(p_input[596]), .B(n25711), .Z(n24844) );
  AND U25617 ( .A(n566), .B(n25712), .Z(n25711) );
  XOR U25618 ( .A(p_input[628]), .B(p_input[596]), .Z(n25712) );
  XNOR U25619 ( .A(n24841), .B(n25707), .Z(n25709) );
  XOR U25620 ( .A(n25713), .B(n25714), .Z(n24841) );
  AND U25621 ( .A(n563), .B(n25715), .Z(n25714) );
  XOR U25622 ( .A(p_input[564]), .B(p_input[532]), .Z(n25715) );
  XOR U25623 ( .A(n25716), .B(n25717), .Z(n25707) );
  AND U25624 ( .A(n25718), .B(n25719), .Z(n25717) );
  XOR U25625 ( .A(n25716), .B(n24856), .Z(n25719) );
  XNOR U25626 ( .A(p_input[595]), .B(n25720), .Z(n24856) );
  AND U25627 ( .A(n566), .B(n25721), .Z(n25720) );
  XOR U25628 ( .A(p_input[627]), .B(p_input[595]), .Z(n25721) );
  XNOR U25629 ( .A(n24853), .B(n25716), .Z(n25718) );
  XOR U25630 ( .A(n25722), .B(n25723), .Z(n24853) );
  AND U25631 ( .A(n563), .B(n25724), .Z(n25723) );
  XOR U25632 ( .A(p_input[563]), .B(p_input[531]), .Z(n25724) );
  XOR U25633 ( .A(n25725), .B(n25726), .Z(n25716) );
  AND U25634 ( .A(n25727), .B(n25728), .Z(n25726) );
  XOR U25635 ( .A(n25725), .B(n24868), .Z(n25728) );
  XNOR U25636 ( .A(p_input[594]), .B(n25729), .Z(n24868) );
  AND U25637 ( .A(n566), .B(n25730), .Z(n25729) );
  XOR U25638 ( .A(p_input[626]), .B(p_input[594]), .Z(n25730) );
  XNOR U25639 ( .A(n24865), .B(n25725), .Z(n25727) );
  XOR U25640 ( .A(n25731), .B(n25732), .Z(n24865) );
  AND U25641 ( .A(n563), .B(n25733), .Z(n25732) );
  XOR U25642 ( .A(p_input[562]), .B(p_input[530]), .Z(n25733) );
  XOR U25643 ( .A(n25734), .B(n25735), .Z(n25725) );
  AND U25644 ( .A(n25736), .B(n25737), .Z(n25735) );
  XOR U25645 ( .A(n25734), .B(n24880), .Z(n25737) );
  XNOR U25646 ( .A(p_input[593]), .B(n25738), .Z(n24880) );
  AND U25647 ( .A(n566), .B(n25739), .Z(n25738) );
  XOR U25648 ( .A(p_input[625]), .B(p_input[593]), .Z(n25739) );
  XNOR U25649 ( .A(n24877), .B(n25734), .Z(n25736) );
  XOR U25650 ( .A(n25740), .B(n25741), .Z(n24877) );
  AND U25651 ( .A(n563), .B(n25742), .Z(n25741) );
  XOR U25652 ( .A(p_input[561]), .B(p_input[529]), .Z(n25742) );
  XOR U25653 ( .A(n25743), .B(n25744), .Z(n25734) );
  AND U25654 ( .A(n25745), .B(n25746), .Z(n25744) );
  XOR U25655 ( .A(n25743), .B(n24892), .Z(n25746) );
  XNOR U25656 ( .A(p_input[592]), .B(n25747), .Z(n24892) );
  AND U25657 ( .A(n566), .B(n25748), .Z(n25747) );
  XOR U25658 ( .A(p_input[624]), .B(p_input[592]), .Z(n25748) );
  XNOR U25659 ( .A(n24889), .B(n25743), .Z(n25745) );
  XOR U25660 ( .A(n25749), .B(n25750), .Z(n24889) );
  AND U25661 ( .A(n563), .B(n25751), .Z(n25750) );
  XOR U25662 ( .A(p_input[560]), .B(p_input[528]), .Z(n25751) );
  XOR U25663 ( .A(n25752), .B(n25753), .Z(n25743) );
  AND U25664 ( .A(n25754), .B(n25755), .Z(n25753) );
  XOR U25665 ( .A(n25752), .B(n24904), .Z(n25755) );
  XNOR U25666 ( .A(p_input[591]), .B(n25756), .Z(n24904) );
  AND U25667 ( .A(n566), .B(n25757), .Z(n25756) );
  XOR U25668 ( .A(p_input[623]), .B(p_input[591]), .Z(n25757) );
  XNOR U25669 ( .A(n24901), .B(n25752), .Z(n25754) );
  XOR U25670 ( .A(n25758), .B(n25759), .Z(n24901) );
  AND U25671 ( .A(n563), .B(n25760), .Z(n25759) );
  XOR U25672 ( .A(p_input[559]), .B(p_input[527]), .Z(n25760) );
  XOR U25673 ( .A(n25761), .B(n25762), .Z(n25752) );
  AND U25674 ( .A(n25763), .B(n25764), .Z(n25762) );
  XOR U25675 ( .A(n25761), .B(n24916), .Z(n25764) );
  XNOR U25676 ( .A(p_input[590]), .B(n25765), .Z(n24916) );
  AND U25677 ( .A(n566), .B(n25766), .Z(n25765) );
  XOR U25678 ( .A(p_input[622]), .B(p_input[590]), .Z(n25766) );
  XNOR U25679 ( .A(n24913), .B(n25761), .Z(n25763) );
  XOR U25680 ( .A(n25767), .B(n25768), .Z(n24913) );
  AND U25681 ( .A(n563), .B(n25769), .Z(n25768) );
  XOR U25682 ( .A(p_input[558]), .B(p_input[526]), .Z(n25769) );
  XOR U25683 ( .A(n25770), .B(n25771), .Z(n25761) );
  AND U25684 ( .A(n25772), .B(n25773), .Z(n25771) );
  XOR U25685 ( .A(n25770), .B(n24928), .Z(n25773) );
  XNOR U25686 ( .A(p_input[589]), .B(n25774), .Z(n24928) );
  AND U25687 ( .A(n566), .B(n25775), .Z(n25774) );
  XOR U25688 ( .A(p_input[621]), .B(p_input[589]), .Z(n25775) );
  XNOR U25689 ( .A(n24925), .B(n25770), .Z(n25772) );
  XOR U25690 ( .A(n25776), .B(n25777), .Z(n24925) );
  AND U25691 ( .A(n563), .B(n25778), .Z(n25777) );
  XOR U25692 ( .A(p_input[557]), .B(p_input[525]), .Z(n25778) );
  XOR U25693 ( .A(n25779), .B(n25780), .Z(n25770) );
  AND U25694 ( .A(n25781), .B(n25782), .Z(n25780) );
  XOR U25695 ( .A(n25779), .B(n24940), .Z(n25782) );
  XNOR U25696 ( .A(p_input[588]), .B(n25783), .Z(n24940) );
  AND U25697 ( .A(n566), .B(n25784), .Z(n25783) );
  XOR U25698 ( .A(p_input[620]), .B(p_input[588]), .Z(n25784) );
  XNOR U25699 ( .A(n24937), .B(n25779), .Z(n25781) );
  XOR U25700 ( .A(n25785), .B(n25786), .Z(n24937) );
  AND U25701 ( .A(n563), .B(n25787), .Z(n25786) );
  XOR U25702 ( .A(p_input[556]), .B(p_input[524]), .Z(n25787) );
  XOR U25703 ( .A(n25788), .B(n25789), .Z(n25779) );
  AND U25704 ( .A(n25790), .B(n25791), .Z(n25789) );
  XOR U25705 ( .A(n25788), .B(n24952), .Z(n25791) );
  XNOR U25706 ( .A(p_input[587]), .B(n25792), .Z(n24952) );
  AND U25707 ( .A(n566), .B(n25793), .Z(n25792) );
  XOR U25708 ( .A(p_input[619]), .B(p_input[587]), .Z(n25793) );
  XNOR U25709 ( .A(n24949), .B(n25788), .Z(n25790) );
  XOR U25710 ( .A(n25794), .B(n25795), .Z(n24949) );
  AND U25711 ( .A(n563), .B(n25796), .Z(n25795) );
  XOR U25712 ( .A(p_input[555]), .B(p_input[523]), .Z(n25796) );
  XOR U25713 ( .A(n25797), .B(n25798), .Z(n25788) );
  AND U25714 ( .A(n25799), .B(n25800), .Z(n25798) );
  XOR U25715 ( .A(n25797), .B(n24964), .Z(n25800) );
  XNOR U25716 ( .A(p_input[586]), .B(n25801), .Z(n24964) );
  AND U25717 ( .A(n566), .B(n25802), .Z(n25801) );
  XOR U25718 ( .A(p_input[618]), .B(p_input[586]), .Z(n25802) );
  XNOR U25719 ( .A(n24961), .B(n25797), .Z(n25799) );
  XOR U25720 ( .A(n25803), .B(n25804), .Z(n24961) );
  AND U25721 ( .A(n563), .B(n25805), .Z(n25804) );
  XOR U25722 ( .A(p_input[554]), .B(p_input[522]), .Z(n25805) );
  XOR U25723 ( .A(n25806), .B(n25807), .Z(n25797) );
  AND U25724 ( .A(n25808), .B(n25809), .Z(n25807) );
  XOR U25725 ( .A(n25806), .B(n24976), .Z(n25809) );
  XNOR U25726 ( .A(p_input[585]), .B(n25810), .Z(n24976) );
  AND U25727 ( .A(n566), .B(n25811), .Z(n25810) );
  XOR U25728 ( .A(p_input[617]), .B(p_input[585]), .Z(n25811) );
  XNOR U25729 ( .A(n24973), .B(n25806), .Z(n25808) );
  XOR U25730 ( .A(n25812), .B(n25813), .Z(n24973) );
  AND U25731 ( .A(n563), .B(n25814), .Z(n25813) );
  XOR U25732 ( .A(p_input[553]), .B(p_input[521]), .Z(n25814) );
  XOR U25733 ( .A(n25815), .B(n25816), .Z(n25806) );
  AND U25734 ( .A(n25817), .B(n25818), .Z(n25816) );
  XOR U25735 ( .A(n25815), .B(n24988), .Z(n25818) );
  XNOR U25736 ( .A(p_input[584]), .B(n25819), .Z(n24988) );
  AND U25737 ( .A(n566), .B(n25820), .Z(n25819) );
  XOR U25738 ( .A(p_input[616]), .B(p_input[584]), .Z(n25820) );
  XNOR U25739 ( .A(n24985), .B(n25815), .Z(n25817) );
  XOR U25740 ( .A(n25821), .B(n25822), .Z(n24985) );
  AND U25741 ( .A(n563), .B(n25823), .Z(n25822) );
  XOR U25742 ( .A(p_input[552]), .B(p_input[520]), .Z(n25823) );
  XOR U25743 ( .A(n25824), .B(n25825), .Z(n25815) );
  AND U25744 ( .A(n25826), .B(n25827), .Z(n25825) );
  XOR U25745 ( .A(n25824), .B(n25000), .Z(n25827) );
  XNOR U25746 ( .A(p_input[583]), .B(n25828), .Z(n25000) );
  AND U25747 ( .A(n566), .B(n25829), .Z(n25828) );
  XOR U25748 ( .A(p_input[615]), .B(p_input[583]), .Z(n25829) );
  XNOR U25749 ( .A(n24997), .B(n25824), .Z(n25826) );
  XOR U25750 ( .A(n25830), .B(n25831), .Z(n24997) );
  AND U25751 ( .A(n563), .B(n25832), .Z(n25831) );
  XOR U25752 ( .A(p_input[551]), .B(p_input[519]), .Z(n25832) );
  XOR U25753 ( .A(n25833), .B(n25834), .Z(n25824) );
  AND U25754 ( .A(n25835), .B(n25836), .Z(n25834) );
  XOR U25755 ( .A(n25833), .B(n25012), .Z(n25836) );
  XNOR U25756 ( .A(p_input[582]), .B(n25837), .Z(n25012) );
  AND U25757 ( .A(n566), .B(n25838), .Z(n25837) );
  XOR U25758 ( .A(p_input[614]), .B(p_input[582]), .Z(n25838) );
  XNOR U25759 ( .A(n25009), .B(n25833), .Z(n25835) );
  XOR U25760 ( .A(n25839), .B(n25840), .Z(n25009) );
  AND U25761 ( .A(n563), .B(n25841), .Z(n25840) );
  XOR U25762 ( .A(p_input[550]), .B(p_input[518]), .Z(n25841) );
  XOR U25763 ( .A(n25842), .B(n25843), .Z(n25833) );
  AND U25764 ( .A(n25844), .B(n25845), .Z(n25843) );
  XOR U25765 ( .A(n25842), .B(n25024), .Z(n25845) );
  XNOR U25766 ( .A(p_input[581]), .B(n25846), .Z(n25024) );
  AND U25767 ( .A(n566), .B(n25847), .Z(n25846) );
  XOR U25768 ( .A(p_input[613]), .B(p_input[581]), .Z(n25847) );
  XNOR U25769 ( .A(n25021), .B(n25842), .Z(n25844) );
  XOR U25770 ( .A(n25848), .B(n25849), .Z(n25021) );
  AND U25771 ( .A(n563), .B(n25850), .Z(n25849) );
  XOR U25772 ( .A(p_input[549]), .B(p_input[517]), .Z(n25850) );
  XOR U25773 ( .A(n25851), .B(n25852), .Z(n25842) );
  AND U25774 ( .A(n25853), .B(n25854), .Z(n25852) );
  XOR U25775 ( .A(n25851), .B(n25036), .Z(n25854) );
  XNOR U25776 ( .A(p_input[580]), .B(n25855), .Z(n25036) );
  AND U25777 ( .A(n566), .B(n25856), .Z(n25855) );
  XOR U25778 ( .A(p_input[612]), .B(p_input[580]), .Z(n25856) );
  XNOR U25779 ( .A(n25033), .B(n25851), .Z(n25853) );
  XOR U25780 ( .A(n25857), .B(n25858), .Z(n25033) );
  AND U25781 ( .A(n563), .B(n25859), .Z(n25858) );
  XOR U25782 ( .A(p_input[548]), .B(p_input[516]), .Z(n25859) );
  XOR U25783 ( .A(n25860), .B(n25861), .Z(n25851) );
  AND U25784 ( .A(n25862), .B(n25863), .Z(n25861) );
  XOR U25785 ( .A(n25860), .B(n25048), .Z(n25863) );
  XNOR U25786 ( .A(p_input[579]), .B(n25864), .Z(n25048) );
  AND U25787 ( .A(n566), .B(n25865), .Z(n25864) );
  XOR U25788 ( .A(p_input[611]), .B(p_input[579]), .Z(n25865) );
  XNOR U25789 ( .A(n25045), .B(n25860), .Z(n25862) );
  XOR U25790 ( .A(n25866), .B(n25867), .Z(n25045) );
  AND U25791 ( .A(n563), .B(n25868), .Z(n25867) );
  XOR U25792 ( .A(p_input[547]), .B(p_input[515]), .Z(n25868) );
  XOR U25793 ( .A(n25869), .B(n25870), .Z(n25860) );
  AND U25794 ( .A(n25871), .B(n25872), .Z(n25870) );
  XOR U25795 ( .A(n25060), .B(n25869), .Z(n25872) );
  XNOR U25796 ( .A(p_input[578]), .B(n25873), .Z(n25060) );
  AND U25797 ( .A(n566), .B(n25874), .Z(n25873) );
  XOR U25798 ( .A(p_input[610]), .B(p_input[578]), .Z(n25874) );
  XNOR U25799 ( .A(n25869), .B(n25057), .Z(n25871) );
  XOR U25800 ( .A(n25875), .B(n25876), .Z(n25057) );
  AND U25801 ( .A(n563), .B(n25877), .Z(n25876) );
  XOR U25802 ( .A(p_input[546]), .B(p_input[514]), .Z(n25877) );
  XOR U25803 ( .A(n25878), .B(n25879), .Z(n25869) );
  AND U25804 ( .A(n25880), .B(n25881), .Z(n25879) );
  XNOR U25805 ( .A(n25882), .B(n25073), .Z(n25881) );
  XNOR U25806 ( .A(p_input[577]), .B(n25883), .Z(n25073) );
  AND U25807 ( .A(n566), .B(n25884), .Z(n25883) );
  XNOR U25808 ( .A(p_input[609]), .B(n25885), .Z(n25884) );
  IV U25809 ( .A(p_input[577]), .Z(n25885) );
  XNOR U25810 ( .A(n25070), .B(n25878), .Z(n25880) );
  XNOR U25811 ( .A(p_input[513]), .B(n25886), .Z(n25070) );
  AND U25812 ( .A(n563), .B(n25887), .Z(n25886) );
  XOR U25813 ( .A(p_input[545]), .B(p_input[513]), .Z(n25887) );
  IV U25814 ( .A(n25882), .Z(n25878) );
  AND U25815 ( .A(n25608), .B(n25611), .Z(n25882) );
  XOR U25816 ( .A(p_input[576]), .B(n25888), .Z(n25611) );
  AND U25817 ( .A(n566), .B(n25889), .Z(n25888) );
  XOR U25818 ( .A(p_input[608]), .B(p_input[576]), .Z(n25889) );
  XOR U25819 ( .A(n25890), .B(n25891), .Z(n566) );
  AND U25820 ( .A(n25892), .B(n25893), .Z(n25891) );
  XNOR U25821 ( .A(p_input[639]), .B(n25890), .Z(n25893) );
  XOR U25822 ( .A(n25890), .B(p_input[607]), .Z(n25892) );
  XOR U25823 ( .A(n25894), .B(n25895), .Z(n25890) );
  AND U25824 ( .A(n25896), .B(n25897), .Z(n25895) );
  XNOR U25825 ( .A(p_input[638]), .B(n25894), .Z(n25897) );
  XOR U25826 ( .A(n25894), .B(p_input[606]), .Z(n25896) );
  XOR U25827 ( .A(n25898), .B(n25899), .Z(n25894) );
  AND U25828 ( .A(n25900), .B(n25901), .Z(n25899) );
  XNOR U25829 ( .A(p_input[637]), .B(n25898), .Z(n25901) );
  XOR U25830 ( .A(n25898), .B(p_input[605]), .Z(n25900) );
  XOR U25831 ( .A(n25902), .B(n25903), .Z(n25898) );
  AND U25832 ( .A(n25904), .B(n25905), .Z(n25903) );
  XNOR U25833 ( .A(p_input[636]), .B(n25902), .Z(n25905) );
  XOR U25834 ( .A(n25902), .B(p_input[604]), .Z(n25904) );
  XOR U25835 ( .A(n25906), .B(n25907), .Z(n25902) );
  AND U25836 ( .A(n25908), .B(n25909), .Z(n25907) );
  XNOR U25837 ( .A(p_input[635]), .B(n25906), .Z(n25909) );
  XOR U25838 ( .A(n25906), .B(p_input[603]), .Z(n25908) );
  XOR U25839 ( .A(n25910), .B(n25911), .Z(n25906) );
  AND U25840 ( .A(n25912), .B(n25913), .Z(n25911) );
  XNOR U25841 ( .A(p_input[634]), .B(n25910), .Z(n25913) );
  XOR U25842 ( .A(n25910), .B(p_input[602]), .Z(n25912) );
  XOR U25843 ( .A(n25914), .B(n25915), .Z(n25910) );
  AND U25844 ( .A(n25916), .B(n25917), .Z(n25915) );
  XNOR U25845 ( .A(p_input[633]), .B(n25914), .Z(n25917) );
  XOR U25846 ( .A(n25914), .B(p_input[601]), .Z(n25916) );
  XOR U25847 ( .A(n25918), .B(n25919), .Z(n25914) );
  AND U25848 ( .A(n25920), .B(n25921), .Z(n25919) );
  XNOR U25849 ( .A(p_input[632]), .B(n25918), .Z(n25921) );
  XOR U25850 ( .A(n25918), .B(p_input[600]), .Z(n25920) );
  XOR U25851 ( .A(n25922), .B(n25923), .Z(n25918) );
  AND U25852 ( .A(n25924), .B(n25925), .Z(n25923) );
  XNOR U25853 ( .A(p_input[631]), .B(n25922), .Z(n25925) );
  XOR U25854 ( .A(n25922), .B(p_input[599]), .Z(n25924) );
  XOR U25855 ( .A(n25926), .B(n25927), .Z(n25922) );
  AND U25856 ( .A(n25928), .B(n25929), .Z(n25927) );
  XNOR U25857 ( .A(p_input[630]), .B(n25926), .Z(n25929) );
  XOR U25858 ( .A(n25926), .B(p_input[598]), .Z(n25928) );
  XOR U25859 ( .A(n25930), .B(n25931), .Z(n25926) );
  AND U25860 ( .A(n25932), .B(n25933), .Z(n25931) );
  XNOR U25861 ( .A(p_input[629]), .B(n25930), .Z(n25933) );
  XOR U25862 ( .A(n25930), .B(p_input[597]), .Z(n25932) );
  XOR U25863 ( .A(n25934), .B(n25935), .Z(n25930) );
  AND U25864 ( .A(n25936), .B(n25937), .Z(n25935) );
  XNOR U25865 ( .A(p_input[628]), .B(n25934), .Z(n25937) );
  XOR U25866 ( .A(n25934), .B(p_input[596]), .Z(n25936) );
  XOR U25867 ( .A(n25938), .B(n25939), .Z(n25934) );
  AND U25868 ( .A(n25940), .B(n25941), .Z(n25939) );
  XNOR U25869 ( .A(p_input[627]), .B(n25938), .Z(n25941) );
  XOR U25870 ( .A(n25938), .B(p_input[595]), .Z(n25940) );
  XOR U25871 ( .A(n25942), .B(n25943), .Z(n25938) );
  AND U25872 ( .A(n25944), .B(n25945), .Z(n25943) );
  XNOR U25873 ( .A(p_input[626]), .B(n25942), .Z(n25945) );
  XOR U25874 ( .A(n25942), .B(p_input[594]), .Z(n25944) );
  XOR U25875 ( .A(n25946), .B(n25947), .Z(n25942) );
  AND U25876 ( .A(n25948), .B(n25949), .Z(n25947) );
  XNOR U25877 ( .A(p_input[625]), .B(n25946), .Z(n25949) );
  XOR U25878 ( .A(n25946), .B(p_input[593]), .Z(n25948) );
  XOR U25879 ( .A(n25950), .B(n25951), .Z(n25946) );
  AND U25880 ( .A(n25952), .B(n25953), .Z(n25951) );
  XNOR U25881 ( .A(p_input[624]), .B(n25950), .Z(n25953) );
  XOR U25882 ( .A(n25950), .B(p_input[592]), .Z(n25952) );
  XOR U25883 ( .A(n25954), .B(n25955), .Z(n25950) );
  AND U25884 ( .A(n25956), .B(n25957), .Z(n25955) );
  XNOR U25885 ( .A(p_input[623]), .B(n25954), .Z(n25957) );
  XOR U25886 ( .A(n25954), .B(p_input[591]), .Z(n25956) );
  XOR U25887 ( .A(n25958), .B(n25959), .Z(n25954) );
  AND U25888 ( .A(n25960), .B(n25961), .Z(n25959) );
  XNOR U25889 ( .A(p_input[622]), .B(n25958), .Z(n25961) );
  XOR U25890 ( .A(n25958), .B(p_input[590]), .Z(n25960) );
  XOR U25891 ( .A(n25962), .B(n25963), .Z(n25958) );
  AND U25892 ( .A(n25964), .B(n25965), .Z(n25963) );
  XNOR U25893 ( .A(p_input[621]), .B(n25962), .Z(n25965) );
  XOR U25894 ( .A(n25962), .B(p_input[589]), .Z(n25964) );
  XOR U25895 ( .A(n25966), .B(n25967), .Z(n25962) );
  AND U25896 ( .A(n25968), .B(n25969), .Z(n25967) );
  XNOR U25897 ( .A(p_input[620]), .B(n25966), .Z(n25969) );
  XOR U25898 ( .A(n25966), .B(p_input[588]), .Z(n25968) );
  XOR U25899 ( .A(n25970), .B(n25971), .Z(n25966) );
  AND U25900 ( .A(n25972), .B(n25973), .Z(n25971) );
  XNOR U25901 ( .A(p_input[619]), .B(n25970), .Z(n25973) );
  XOR U25902 ( .A(n25970), .B(p_input[587]), .Z(n25972) );
  XOR U25903 ( .A(n25974), .B(n25975), .Z(n25970) );
  AND U25904 ( .A(n25976), .B(n25977), .Z(n25975) );
  XNOR U25905 ( .A(p_input[618]), .B(n25974), .Z(n25977) );
  XOR U25906 ( .A(n25974), .B(p_input[586]), .Z(n25976) );
  XOR U25907 ( .A(n25978), .B(n25979), .Z(n25974) );
  AND U25908 ( .A(n25980), .B(n25981), .Z(n25979) );
  XNOR U25909 ( .A(p_input[617]), .B(n25978), .Z(n25981) );
  XOR U25910 ( .A(n25978), .B(p_input[585]), .Z(n25980) );
  XOR U25911 ( .A(n25982), .B(n25983), .Z(n25978) );
  AND U25912 ( .A(n25984), .B(n25985), .Z(n25983) );
  XNOR U25913 ( .A(p_input[616]), .B(n25982), .Z(n25985) );
  XOR U25914 ( .A(n25982), .B(p_input[584]), .Z(n25984) );
  XOR U25915 ( .A(n25986), .B(n25987), .Z(n25982) );
  AND U25916 ( .A(n25988), .B(n25989), .Z(n25987) );
  XNOR U25917 ( .A(p_input[615]), .B(n25986), .Z(n25989) );
  XOR U25918 ( .A(n25986), .B(p_input[583]), .Z(n25988) );
  XOR U25919 ( .A(n25990), .B(n25991), .Z(n25986) );
  AND U25920 ( .A(n25992), .B(n25993), .Z(n25991) );
  XNOR U25921 ( .A(p_input[614]), .B(n25990), .Z(n25993) );
  XOR U25922 ( .A(n25990), .B(p_input[582]), .Z(n25992) );
  XOR U25923 ( .A(n25994), .B(n25995), .Z(n25990) );
  AND U25924 ( .A(n25996), .B(n25997), .Z(n25995) );
  XNOR U25925 ( .A(p_input[613]), .B(n25994), .Z(n25997) );
  XOR U25926 ( .A(n25994), .B(p_input[581]), .Z(n25996) );
  XOR U25927 ( .A(n25998), .B(n25999), .Z(n25994) );
  AND U25928 ( .A(n26000), .B(n26001), .Z(n25999) );
  XNOR U25929 ( .A(p_input[612]), .B(n25998), .Z(n26001) );
  XOR U25930 ( .A(n25998), .B(p_input[580]), .Z(n26000) );
  XOR U25931 ( .A(n26002), .B(n26003), .Z(n25998) );
  AND U25932 ( .A(n26004), .B(n26005), .Z(n26003) );
  XNOR U25933 ( .A(p_input[611]), .B(n26002), .Z(n26005) );
  XOR U25934 ( .A(n26002), .B(p_input[579]), .Z(n26004) );
  XOR U25935 ( .A(n26006), .B(n26007), .Z(n26002) );
  AND U25936 ( .A(n26008), .B(n26009), .Z(n26007) );
  XNOR U25937 ( .A(p_input[610]), .B(n26006), .Z(n26009) );
  XOR U25938 ( .A(n26006), .B(p_input[578]), .Z(n26008) );
  XNOR U25939 ( .A(n26010), .B(n26011), .Z(n26006) );
  AND U25940 ( .A(n26012), .B(n26013), .Z(n26011) );
  XOR U25941 ( .A(p_input[609]), .B(n26010), .Z(n26013) );
  XNOR U25942 ( .A(p_input[577]), .B(n26010), .Z(n26012) );
  AND U25943 ( .A(p_input[608]), .B(n26014), .Z(n26010) );
  IV U25944 ( .A(p_input[576]), .Z(n26014) );
  XNOR U25945 ( .A(p_input[512]), .B(n26015), .Z(n25608) );
  AND U25946 ( .A(n563), .B(n26016), .Z(n26015) );
  XOR U25947 ( .A(p_input[544]), .B(p_input[512]), .Z(n26016) );
  XOR U25948 ( .A(n26017), .B(n26018), .Z(n563) );
  AND U25949 ( .A(n26019), .B(n26020), .Z(n26018) );
  XNOR U25950 ( .A(p_input[575]), .B(n26017), .Z(n26020) );
  XOR U25951 ( .A(n26017), .B(p_input[543]), .Z(n26019) );
  XOR U25952 ( .A(n26021), .B(n26022), .Z(n26017) );
  AND U25953 ( .A(n26023), .B(n26024), .Z(n26022) );
  XNOR U25954 ( .A(p_input[574]), .B(n26021), .Z(n26024) );
  XNOR U25955 ( .A(n26021), .B(n25623), .Z(n26023) );
  IV U25956 ( .A(p_input[542]), .Z(n25623) );
  XOR U25957 ( .A(n26025), .B(n26026), .Z(n26021) );
  AND U25958 ( .A(n26027), .B(n26028), .Z(n26026) );
  XNOR U25959 ( .A(p_input[573]), .B(n26025), .Z(n26028) );
  XNOR U25960 ( .A(n26025), .B(n25632), .Z(n26027) );
  IV U25961 ( .A(p_input[541]), .Z(n25632) );
  XOR U25962 ( .A(n26029), .B(n26030), .Z(n26025) );
  AND U25963 ( .A(n26031), .B(n26032), .Z(n26030) );
  XNOR U25964 ( .A(p_input[572]), .B(n26029), .Z(n26032) );
  XNOR U25965 ( .A(n26029), .B(n25641), .Z(n26031) );
  IV U25966 ( .A(p_input[540]), .Z(n25641) );
  XOR U25967 ( .A(n26033), .B(n26034), .Z(n26029) );
  AND U25968 ( .A(n26035), .B(n26036), .Z(n26034) );
  XNOR U25969 ( .A(p_input[571]), .B(n26033), .Z(n26036) );
  XNOR U25970 ( .A(n26033), .B(n25650), .Z(n26035) );
  IV U25971 ( .A(p_input[539]), .Z(n25650) );
  XOR U25972 ( .A(n26037), .B(n26038), .Z(n26033) );
  AND U25973 ( .A(n26039), .B(n26040), .Z(n26038) );
  XNOR U25974 ( .A(p_input[570]), .B(n26037), .Z(n26040) );
  XNOR U25975 ( .A(n26037), .B(n25659), .Z(n26039) );
  IV U25976 ( .A(p_input[538]), .Z(n25659) );
  XOR U25977 ( .A(n26041), .B(n26042), .Z(n26037) );
  AND U25978 ( .A(n26043), .B(n26044), .Z(n26042) );
  XNOR U25979 ( .A(p_input[569]), .B(n26041), .Z(n26044) );
  XNOR U25980 ( .A(n26041), .B(n25668), .Z(n26043) );
  IV U25981 ( .A(p_input[537]), .Z(n25668) );
  XOR U25982 ( .A(n26045), .B(n26046), .Z(n26041) );
  AND U25983 ( .A(n26047), .B(n26048), .Z(n26046) );
  XNOR U25984 ( .A(p_input[568]), .B(n26045), .Z(n26048) );
  XNOR U25985 ( .A(n26045), .B(n25677), .Z(n26047) );
  IV U25986 ( .A(p_input[536]), .Z(n25677) );
  XOR U25987 ( .A(n26049), .B(n26050), .Z(n26045) );
  AND U25988 ( .A(n26051), .B(n26052), .Z(n26050) );
  XNOR U25989 ( .A(p_input[567]), .B(n26049), .Z(n26052) );
  XNOR U25990 ( .A(n26049), .B(n25686), .Z(n26051) );
  IV U25991 ( .A(p_input[535]), .Z(n25686) );
  XOR U25992 ( .A(n26053), .B(n26054), .Z(n26049) );
  AND U25993 ( .A(n26055), .B(n26056), .Z(n26054) );
  XNOR U25994 ( .A(p_input[566]), .B(n26053), .Z(n26056) );
  XNOR U25995 ( .A(n26053), .B(n25695), .Z(n26055) );
  IV U25996 ( .A(p_input[534]), .Z(n25695) );
  XOR U25997 ( .A(n26057), .B(n26058), .Z(n26053) );
  AND U25998 ( .A(n26059), .B(n26060), .Z(n26058) );
  XNOR U25999 ( .A(p_input[565]), .B(n26057), .Z(n26060) );
  XNOR U26000 ( .A(n26057), .B(n25704), .Z(n26059) );
  IV U26001 ( .A(p_input[533]), .Z(n25704) );
  XOR U26002 ( .A(n26061), .B(n26062), .Z(n26057) );
  AND U26003 ( .A(n26063), .B(n26064), .Z(n26062) );
  XNOR U26004 ( .A(p_input[564]), .B(n26061), .Z(n26064) );
  XNOR U26005 ( .A(n26061), .B(n25713), .Z(n26063) );
  IV U26006 ( .A(p_input[532]), .Z(n25713) );
  XOR U26007 ( .A(n26065), .B(n26066), .Z(n26061) );
  AND U26008 ( .A(n26067), .B(n26068), .Z(n26066) );
  XNOR U26009 ( .A(p_input[563]), .B(n26065), .Z(n26068) );
  XNOR U26010 ( .A(n26065), .B(n25722), .Z(n26067) );
  IV U26011 ( .A(p_input[531]), .Z(n25722) );
  XOR U26012 ( .A(n26069), .B(n26070), .Z(n26065) );
  AND U26013 ( .A(n26071), .B(n26072), .Z(n26070) );
  XNOR U26014 ( .A(p_input[562]), .B(n26069), .Z(n26072) );
  XNOR U26015 ( .A(n26069), .B(n25731), .Z(n26071) );
  IV U26016 ( .A(p_input[530]), .Z(n25731) );
  XOR U26017 ( .A(n26073), .B(n26074), .Z(n26069) );
  AND U26018 ( .A(n26075), .B(n26076), .Z(n26074) );
  XNOR U26019 ( .A(p_input[561]), .B(n26073), .Z(n26076) );
  XNOR U26020 ( .A(n26073), .B(n25740), .Z(n26075) );
  IV U26021 ( .A(p_input[529]), .Z(n25740) );
  XOR U26022 ( .A(n26077), .B(n26078), .Z(n26073) );
  AND U26023 ( .A(n26079), .B(n26080), .Z(n26078) );
  XNOR U26024 ( .A(p_input[560]), .B(n26077), .Z(n26080) );
  XNOR U26025 ( .A(n26077), .B(n25749), .Z(n26079) );
  IV U26026 ( .A(p_input[528]), .Z(n25749) );
  XOR U26027 ( .A(n26081), .B(n26082), .Z(n26077) );
  AND U26028 ( .A(n26083), .B(n26084), .Z(n26082) );
  XNOR U26029 ( .A(p_input[559]), .B(n26081), .Z(n26084) );
  XNOR U26030 ( .A(n26081), .B(n25758), .Z(n26083) );
  IV U26031 ( .A(p_input[527]), .Z(n25758) );
  XOR U26032 ( .A(n26085), .B(n26086), .Z(n26081) );
  AND U26033 ( .A(n26087), .B(n26088), .Z(n26086) );
  XNOR U26034 ( .A(p_input[558]), .B(n26085), .Z(n26088) );
  XNOR U26035 ( .A(n26085), .B(n25767), .Z(n26087) );
  IV U26036 ( .A(p_input[526]), .Z(n25767) );
  XOR U26037 ( .A(n26089), .B(n26090), .Z(n26085) );
  AND U26038 ( .A(n26091), .B(n26092), .Z(n26090) );
  XNOR U26039 ( .A(p_input[557]), .B(n26089), .Z(n26092) );
  XNOR U26040 ( .A(n26089), .B(n25776), .Z(n26091) );
  IV U26041 ( .A(p_input[525]), .Z(n25776) );
  XOR U26042 ( .A(n26093), .B(n26094), .Z(n26089) );
  AND U26043 ( .A(n26095), .B(n26096), .Z(n26094) );
  XNOR U26044 ( .A(p_input[556]), .B(n26093), .Z(n26096) );
  XNOR U26045 ( .A(n26093), .B(n25785), .Z(n26095) );
  IV U26046 ( .A(p_input[524]), .Z(n25785) );
  XOR U26047 ( .A(n26097), .B(n26098), .Z(n26093) );
  AND U26048 ( .A(n26099), .B(n26100), .Z(n26098) );
  XNOR U26049 ( .A(p_input[555]), .B(n26097), .Z(n26100) );
  XNOR U26050 ( .A(n26097), .B(n25794), .Z(n26099) );
  IV U26051 ( .A(p_input[523]), .Z(n25794) );
  XOR U26052 ( .A(n26101), .B(n26102), .Z(n26097) );
  AND U26053 ( .A(n26103), .B(n26104), .Z(n26102) );
  XNOR U26054 ( .A(p_input[554]), .B(n26101), .Z(n26104) );
  XNOR U26055 ( .A(n26101), .B(n25803), .Z(n26103) );
  IV U26056 ( .A(p_input[522]), .Z(n25803) );
  XOR U26057 ( .A(n26105), .B(n26106), .Z(n26101) );
  AND U26058 ( .A(n26107), .B(n26108), .Z(n26106) );
  XNOR U26059 ( .A(p_input[553]), .B(n26105), .Z(n26108) );
  XNOR U26060 ( .A(n26105), .B(n25812), .Z(n26107) );
  IV U26061 ( .A(p_input[521]), .Z(n25812) );
  XOR U26062 ( .A(n26109), .B(n26110), .Z(n26105) );
  AND U26063 ( .A(n26111), .B(n26112), .Z(n26110) );
  XNOR U26064 ( .A(p_input[552]), .B(n26109), .Z(n26112) );
  XNOR U26065 ( .A(n26109), .B(n25821), .Z(n26111) );
  IV U26066 ( .A(p_input[520]), .Z(n25821) );
  XOR U26067 ( .A(n26113), .B(n26114), .Z(n26109) );
  AND U26068 ( .A(n26115), .B(n26116), .Z(n26114) );
  XNOR U26069 ( .A(p_input[551]), .B(n26113), .Z(n26116) );
  XNOR U26070 ( .A(n26113), .B(n25830), .Z(n26115) );
  IV U26071 ( .A(p_input[519]), .Z(n25830) );
  XOR U26072 ( .A(n26117), .B(n26118), .Z(n26113) );
  AND U26073 ( .A(n26119), .B(n26120), .Z(n26118) );
  XNOR U26074 ( .A(p_input[550]), .B(n26117), .Z(n26120) );
  XNOR U26075 ( .A(n26117), .B(n25839), .Z(n26119) );
  IV U26076 ( .A(p_input[518]), .Z(n25839) );
  XOR U26077 ( .A(n26121), .B(n26122), .Z(n26117) );
  AND U26078 ( .A(n26123), .B(n26124), .Z(n26122) );
  XNOR U26079 ( .A(p_input[549]), .B(n26121), .Z(n26124) );
  XNOR U26080 ( .A(n26121), .B(n25848), .Z(n26123) );
  IV U26081 ( .A(p_input[517]), .Z(n25848) );
  XOR U26082 ( .A(n26125), .B(n26126), .Z(n26121) );
  AND U26083 ( .A(n26127), .B(n26128), .Z(n26126) );
  XNOR U26084 ( .A(p_input[548]), .B(n26125), .Z(n26128) );
  XNOR U26085 ( .A(n26125), .B(n25857), .Z(n26127) );
  IV U26086 ( .A(p_input[516]), .Z(n25857) );
  XOR U26087 ( .A(n26129), .B(n26130), .Z(n26125) );
  AND U26088 ( .A(n26131), .B(n26132), .Z(n26130) );
  XNOR U26089 ( .A(p_input[547]), .B(n26129), .Z(n26132) );
  XNOR U26090 ( .A(n26129), .B(n25866), .Z(n26131) );
  IV U26091 ( .A(p_input[515]), .Z(n25866) );
  XOR U26092 ( .A(n26133), .B(n26134), .Z(n26129) );
  AND U26093 ( .A(n26135), .B(n26136), .Z(n26134) );
  XNOR U26094 ( .A(p_input[546]), .B(n26133), .Z(n26136) );
  XNOR U26095 ( .A(n26133), .B(n25875), .Z(n26135) );
  IV U26096 ( .A(p_input[514]), .Z(n25875) );
  XNOR U26097 ( .A(n26137), .B(n26138), .Z(n26133) );
  AND U26098 ( .A(n26139), .B(n26140), .Z(n26138) );
  XOR U26099 ( .A(p_input[545]), .B(n26137), .Z(n26140) );
  XNOR U26100 ( .A(p_input[513]), .B(n26137), .Z(n26139) );
  AND U26101 ( .A(p_input[544]), .B(n26141), .Z(n26137) );
  IV U26102 ( .A(p_input[512]), .Z(n26141) );
  XOR U26103 ( .A(n26142), .B(n26143), .Z(n22498) );
  AND U26104 ( .A(n591), .B(n26144), .Z(n26143) );
  XNOR U26105 ( .A(n26145), .B(n26142), .Z(n26144) );
  XOR U26106 ( .A(n26146), .B(n26147), .Z(n591) );
  AND U26107 ( .A(n26148), .B(n26149), .Z(n26147) );
  XOR U26108 ( .A(n26146), .B(n22513), .Z(n26149) );
  XOR U26109 ( .A(n26150), .B(n26151), .Z(n22513) );
  AND U26110 ( .A(n534), .B(n26152), .Z(n26151) );
  XOR U26111 ( .A(n26153), .B(n26150), .Z(n26152) );
  XNOR U26112 ( .A(n22510), .B(n26146), .Z(n26148) );
  XOR U26113 ( .A(n26154), .B(n26155), .Z(n22510) );
  AND U26114 ( .A(n531), .B(n26156), .Z(n26155) );
  XOR U26115 ( .A(n26157), .B(n26154), .Z(n26156) );
  XOR U26116 ( .A(n26158), .B(n26159), .Z(n26146) );
  AND U26117 ( .A(n26160), .B(n26161), .Z(n26159) );
  XOR U26118 ( .A(n26158), .B(n22525), .Z(n26161) );
  XOR U26119 ( .A(n26162), .B(n26163), .Z(n22525) );
  AND U26120 ( .A(n534), .B(n26164), .Z(n26163) );
  XOR U26121 ( .A(n26165), .B(n26162), .Z(n26164) );
  XNOR U26122 ( .A(n22522), .B(n26158), .Z(n26160) );
  XOR U26123 ( .A(n26166), .B(n26167), .Z(n22522) );
  AND U26124 ( .A(n531), .B(n26168), .Z(n26167) );
  XOR U26125 ( .A(n26169), .B(n26166), .Z(n26168) );
  XOR U26126 ( .A(n26170), .B(n26171), .Z(n26158) );
  AND U26127 ( .A(n26172), .B(n26173), .Z(n26171) );
  XOR U26128 ( .A(n26170), .B(n22537), .Z(n26173) );
  XOR U26129 ( .A(n26174), .B(n26175), .Z(n22537) );
  AND U26130 ( .A(n534), .B(n26176), .Z(n26175) );
  XOR U26131 ( .A(n26177), .B(n26174), .Z(n26176) );
  XNOR U26132 ( .A(n22534), .B(n26170), .Z(n26172) );
  XOR U26133 ( .A(n26178), .B(n26179), .Z(n22534) );
  AND U26134 ( .A(n531), .B(n26180), .Z(n26179) );
  XOR U26135 ( .A(n26181), .B(n26178), .Z(n26180) );
  XOR U26136 ( .A(n26182), .B(n26183), .Z(n26170) );
  AND U26137 ( .A(n26184), .B(n26185), .Z(n26183) );
  XOR U26138 ( .A(n26182), .B(n22549), .Z(n26185) );
  XOR U26139 ( .A(n26186), .B(n26187), .Z(n22549) );
  AND U26140 ( .A(n534), .B(n26188), .Z(n26187) );
  XOR U26141 ( .A(n26189), .B(n26186), .Z(n26188) );
  XNOR U26142 ( .A(n22546), .B(n26182), .Z(n26184) );
  XOR U26143 ( .A(n26190), .B(n26191), .Z(n22546) );
  AND U26144 ( .A(n531), .B(n26192), .Z(n26191) );
  XOR U26145 ( .A(n26193), .B(n26190), .Z(n26192) );
  XOR U26146 ( .A(n26194), .B(n26195), .Z(n26182) );
  AND U26147 ( .A(n26196), .B(n26197), .Z(n26195) );
  XOR U26148 ( .A(n26194), .B(n22561), .Z(n26197) );
  XOR U26149 ( .A(n26198), .B(n26199), .Z(n22561) );
  AND U26150 ( .A(n534), .B(n26200), .Z(n26199) );
  XOR U26151 ( .A(n26201), .B(n26198), .Z(n26200) );
  XNOR U26152 ( .A(n22558), .B(n26194), .Z(n26196) );
  XOR U26153 ( .A(n26202), .B(n26203), .Z(n22558) );
  AND U26154 ( .A(n531), .B(n26204), .Z(n26203) );
  XOR U26155 ( .A(n26205), .B(n26202), .Z(n26204) );
  XOR U26156 ( .A(n26206), .B(n26207), .Z(n26194) );
  AND U26157 ( .A(n26208), .B(n26209), .Z(n26207) );
  XOR U26158 ( .A(n26206), .B(n22573), .Z(n26209) );
  XOR U26159 ( .A(n26210), .B(n26211), .Z(n22573) );
  AND U26160 ( .A(n534), .B(n26212), .Z(n26211) );
  XOR U26161 ( .A(n26213), .B(n26210), .Z(n26212) );
  XNOR U26162 ( .A(n22570), .B(n26206), .Z(n26208) );
  XOR U26163 ( .A(n26214), .B(n26215), .Z(n22570) );
  AND U26164 ( .A(n531), .B(n26216), .Z(n26215) );
  XOR U26165 ( .A(n26217), .B(n26214), .Z(n26216) );
  XOR U26166 ( .A(n26218), .B(n26219), .Z(n26206) );
  AND U26167 ( .A(n26220), .B(n26221), .Z(n26219) );
  XOR U26168 ( .A(n26218), .B(n22585), .Z(n26221) );
  XOR U26169 ( .A(n26222), .B(n26223), .Z(n22585) );
  AND U26170 ( .A(n534), .B(n26224), .Z(n26223) );
  XOR U26171 ( .A(n26225), .B(n26222), .Z(n26224) );
  XNOR U26172 ( .A(n22582), .B(n26218), .Z(n26220) );
  XOR U26173 ( .A(n26226), .B(n26227), .Z(n22582) );
  AND U26174 ( .A(n531), .B(n26228), .Z(n26227) );
  XOR U26175 ( .A(n26229), .B(n26226), .Z(n26228) );
  XOR U26176 ( .A(n26230), .B(n26231), .Z(n26218) );
  AND U26177 ( .A(n26232), .B(n26233), .Z(n26231) );
  XOR U26178 ( .A(n26230), .B(n22597), .Z(n26233) );
  XOR U26179 ( .A(n26234), .B(n26235), .Z(n22597) );
  AND U26180 ( .A(n534), .B(n26236), .Z(n26235) );
  XOR U26181 ( .A(n26237), .B(n26234), .Z(n26236) );
  XNOR U26182 ( .A(n22594), .B(n26230), .Z(n26232) );
  XOR U26183 ( .A(n26238), .B(n26239), .Z(n22594) );
  AND U26184 ( .A(n531), .B(n26240), .Z(n26239) );
  XOR U26185 ( .A(n26241), .B(n26238), .Z(n26240) );
  XOR U26186 ( .A(n26242), .B(n26243), .Z(n26230) );
  AND U26187 ( .A(n26244), .B(n26245), .Z(n26243) );
  XOR U26188 ( .A(n26242), .B(n22609), .Z(n26245) );
  XOR U26189 ( .A(n26246), .B(n26247), .Z(n22609) );
  AND U26190 ( .A(n534), .B(n26248), .Z(n26247) );
  XOR U26191 ( .A(n26249), .B(n26246), .Z(n26248) );
  XNOR U26192 ( .A(n22606), .B(n26242), .Z(n26244) );
  XOR U26193 ( .A(n26250), .B(n26251), .Z(n22606) );
  AND U26194 ( .A(n531), .B(n26252), .Z(n26251) );
  XOR U26195 ( .A(n26253), .B(n26250), .Z(n26252) );
  XOR U26196 ( .A(n26254), .B(n26255), .Z(n26242) );
  AND U26197 ( .A(n26256), .B(n26257), .Z(n26255) );
  XOR U26198 ( .A(n26254), .B(n22621), .Z(n26257) );
  XOR U26199 ( .A(n26258), .B(n26259), .Z(n22621) );
  AND U26200 ( .A(n534), .B(n26260), .Z(n26259) );
  XOR U26201 ( .A(n26261), .B(n26258), .Z(n26260) );
  XNOR U26202 ( .A(n22618), .B(n26254), .Z(n26256) );
  XOR U26203 ( .A(n26262), .B(n26263), .Z(n22618) );
  AND U26204 ( .A(n531), .B(n26264), .Z(n26263) );
  XOR U26205 ( .A(n26265), .B(n26262), .Z(n26264) );
  XOR U26206 ( .A(n26266), .B(n26267), .Z(n26254) );
  AND U26207 ( .A(n26268), .B(n26269), .Z(n26267) );
  XOR U26208 ( .A(n26266), .B(n22633), .Z(n26269) );
  XOR U26209 ( .A(n26270), .B(n26271), .Z(n22633) );
  AND U26210 ( .A(n534), .B(n26272), .Z(n26271) );
  XOR U26211 ( .A(n26273), .B(n26270), .Z(n26272) );
  XNOR U26212 ( .A(n22630), .B(n26266), .Z(n26268) );
  XOR U26213 ( .A(n26274), .B(n26275), .Z(n22630) );
  AND U26214 ( .A(n531), .B(n26276), .Z(n26275) );
  XOR U26215 ( .A(n26277), .B(n26274), .Z(n26276) );
  XOR U26216 ( .A(n26278), .B(n26279), .Z(n26266) );
  AND U26217 ( .A(n26280), .B(n26281), .Z(n26279) );
  XOR U26218 ( .A(n26278), .B(n22645), .Z(n26281) );
  XOR U26219 ( .A(n26282), .B(n26283), .Z(n22645) );
  AND U26220 ( .A(n534), .B(n26284), .Z(n26283) );
  XOR U26221 ( .A(n26285), .B(n26282), .Z(n26284) );
  XNOR U26222 ( .A(n22642), .B(n26278), .Z(n26280) );
  XOR U26223 ( .A(n26286), .B(n26287), .Z(n22642) );
  AND U26224 ( .A(n531), .B(n26288), .Z(n26287) );
  XOR U26225 ( .A(n26289), .B(n26286), .Z(n26288) );
  XOR U26226 ( .A(n26290), .B(n26291), .Z(n26278) );
  AND U26227 ( .A(n26292), .B(n26293), .Z(n26291) );
  XOR U26228 ( .A(n26290), .B(n22657), .Z(n26293) );
  XOR U26229 ( .A(n26294), .B(n26295), .Z(n22657) );
  AND U26230 ( .A(n534), .B(n26296), .Z(n26295) );
  XOR U26231 ( .A(n26297), .B(n26294), .Z(n26296) );
  XNOR U26232 ( .A(n22654), .B(n26290), .Z(n26292) );
  XOR U26233 ( .A(n26298), .B(n26299), .Z(n22654) );
  AND U26234 ( .A(n531), .B(n26300), .Z(n26299) );
  XOR U26235 ( .A(n26301), .B(n26298), .Z(n26300) );
  XOR U26236 ( .A(n26302), .B(n26303), .Z(n26290) );
  AND U26237 ( .A(n26304), .B(n26305), .Z(n26303) );
  XOR U26238 ( .A(n26302), .B(n22669), .Z(n26305) );
  XOR U26239 ( .A(n26306), .B(n26307), .Z(n22669) );
  AND U26240 ( .A(n534), .B(n26308), .Z(n26307) );
  XOR U26241 ( .A(n26309), .B(n26306), .Z(n26308) );
  XNOR U26242 ( .A(n22666), .B(n26302), .Z(n26304) );
  XOR U26243 ( .A(n26310), .B(n26311), .Z(n22666) );
  AND U26244 ( .A(n531), .B(n26312), .Z(n26311) );
  XOR U26245 ( .A(n26313), .B(n26310), .Z(n26312) );
  XOR U26246 ( .A(n26314), .B(n26315), .Z(n26302) );
  AND U26247 ( .A(n26316), .B(n26317), .Z(n26315) );
  XOR U26248 ( .A(n26314), .B(n22681), .Z(n26317) );
  XOR U26249 ( .A(n26318), .B(n26319), .Z(n22681) );
  AND U26250 ( .A(n534), .B(n26320), .Z(n26319) );
  XOR U26251 ( .A(n26321), .B(n26318), .Z(n26320) );
  XNOR U26252 ( .A(n22678), .B(n26314), .Z(n26316) );
  XOR U26253 ( .A(n26322), .B(n26323), .Z(n22678) );
  AND U26254 ( .A(n531), .B(n26324), .Z(n26323) );
  XOR U26255 ( .A(n26325), .B(n26322), .Z(n26324) );
  XOR U26256 ( .A(n26326), .B(n26327), .Z(n26314) );
  AND U26257 ( .A(n26328), .B(n26329), .Z(n26327) );
  XOR U26258 ( .A(n26326), .B(n22693), .Z(n26329) );
  XOR U26259 ( .A(n26330), .B(n26331), .Z(n22693) );
  AND U26260 ( .A(n534), .B(n26332), .Z(n26331) );
  XOR U26261 ( .A(n26333), .B(n26330), .Z(n26332) );
  XNOR U26262 ( .A(n22690), .B(n26326), .Z(n26328) );
  XOR U26263 ( .A(n26334), .B(n26335), .Z(n22690) );
  AND U26264 ( .A(n531), .B(n26336), .Z(n26335) );
  XOR U26265 ( .A(n26337), .B(n26334), .Z(n26336) );
  XOR U26266 ( .A(n26338), .B(n26339), .Z(n26326) );
  AND U26267 ( .A(n26340), .B(n26341), .Z(n26339) );
  XOR U26268 ( .A(n26338), .B(n22705), .Z(n26341) );
  XOR U26269 ( .A(n26342), .B(n26343), .Z(n22705) );
  AND U26270 ( .A(n534), .B(n26344), .Z(n26343) );
  XOR U26271 ( .A(n26345), .B(n26342), .Z(n26344) );
  XNOR U26272 ( .A(n22702), .B(n26338), .Z(n26340) );
  XOR U26273 ( .A(n26346), .B(n26347), .Z(n22702) );
  AND U26274 ( .A(n531), .B(n26348), .Z(n26347) );
  XOR U26275 ( .A(n26349), .B(n26346), .Z(n26348) );
  XOR U26276 ( .A(n26350), .B(n26351), .Z(n26338) );
  AND U26277 ( .A(n26352), .B(n26353), .Z(n26351) );
  XOR U26278 ( .A(n26350), .B(n22717), .Z(n26353) );
  XOR U26279 ( .A(n26354), .B(n26355), .Z(n22717) );
  AND U26280 ( .A(n534), .B(n26356), .Z(n26355) );
  XOR U26281 ( .A(n26357), .B(n26354), .Z(n26356) );
  XNOR U26282 ( .A(n22714), .B(n26350), .Z(n26352) );
  XOR U26283 ( .A(n26358), .B(n26359), .Z(n22714) );
  AND U26284 ( .A(n531), .B(n26360), .Z(n26359) );
  XOR U26285 ( .A(n26361), .B(n26358), .Z(n26360) );
  XOR U26286 ( .A(n26362), .B(n26363), .Z(n26350) );
  AND U26287 ( .A(n26364), .B(n26365), .Z(n26363) );
  XOR U26288 ( .A(n26362), .B(n22729), .Z(n26365) );
  XOR U26289 ( .A(n26366), .B(n26367), .Z(n22729) );
  AND U26290 ( .A(n534), .B(n26368), .Z(n26367) );
  XOR U26291 ( .A(n26369), .B(n26366), .Z(n26368) );
  XNOR U26292 ( .A(n22726), .B(n26362), .Z(n26364) );
  XOR U26293 ( .A(n26370), .B(n26371), .Z(n22726) );
  AND U26294 ( .A(n531), .B(n26372), .Z(n26371) );
  XOR U26295 ( .A(n26373), .B(n26370), .Z(n26372) );
  XOR U26296 ( .A(n26374), .B(n26375), .Z(n26362) );
  AND U26297 ( .A(n26376), .B(n26377), .Z(n26375) );
  XOR U26298 ( .A(n26374), .B(n22741), .Z(n26377) );
  XOR U26299 ( .A(n26378), .B(n26379), .Z(n22741) );
  AND U26300 ( .A(n534), .B(n26380), .Z(n26379) );
  XOR U26301 ( .A(n26381), .B(n26378), .Z(n26380) );
  XNOR U26302 ( .A(n22738), .B(n26374), .Z(n26376) );
  XOR U26303 ( .A(n26382), .B(n26383), .Z(n22738) );
  AND U26304 ( .A(n531), .B(n26384), .Z(n26383) );
  XOR U26305 ( .A(n26385), .B(n26382), .Z(n26384) );
  XOR U26306 ( .A(n26386), .B(n26387), .Z(n26374) );
  AND U26307 ( .A(n26388), .B(n26389), .Z(n26387) );
  XOR U26308 ( .A(n26386), .B(n22753), .Z(n26389) );
  XOR U26309 ( .A(n26390), .B(n26391), .Z(n22753) );
  AND U26310 ( .A(n534), .B(n26392), .Z(n26391) );
  XOR U26311 ( .A(n26393), .B(n26390), .Z(n26392) );
  XNOR U26312 ( .A(n22750), .B(n26386), .Z(n26388) );
  XOR U26313 ( .A(n26394), .B(n26395), .Z(n22750) );
  AND U26314 ( .A(n531), .B(n26396), .Z(n26395) );
  XOR U26315 ( .A(n26397), .B(n26394), .Z(n26396) );
  XOR U26316 ( .A(n26398), .B(n26399), .Z(n26386) );
  AND U26317 ( .A(n26400), .B(n26401), .Z(n26399) );
  XOR U26318 ( .A(n26398), .B(n22765), .Z(n26401) );
  XOR U26319 ( .A(n26402), .B(n26403), .Z(n22765) );
  AND U26320 ( .A(n534), .B(n26404), .Z(n26403) );
  XOR U26321 ( .A(n26405), .B(n26402), .Z(n26404) );
  XNOR U26322 ( .A(n22762), .B(n26398), .Z(n26400) );
  XOR U26323 ( .A(n26406), .B(n26407), .Z(n22762) );
  AND U26324 ( .A(n531), .B(n26408), .Z(n26407) );
  XOR U26325 ( .A(n26409), .B(n26406), .Z(n26408) );
  XOR U26326 ( .A(n26410), .B(n26411), .Z(n26398) );
  AND U26327 ( .A(n26412), .B(n26413), .Z(n26411) );
  XOR U26328 ( .A(n26410), .B(n22777), .Z(n26413) );
  XOR U26329 ( .A(n26414), .B(n26415), .Z(n22777) );
  AND U26330 ( .A(n534), .B(n26416), .Z(n26415) );
  XOR U26331 ( .A(n26417), .B(n26414), .Z(n26416) );
  XNOR U26332 ( .A(n22774), .B(n26410), .Z(n26412) );
  XOR U26333 ( .A(n26418), .B(n26419), .Z(n22774) );
  AND U26334 ( .A(n531), .B(n26420), .Z(n26419) );
  XOR U26335 ( .A(n26421), .B(n26418), .Z(n26420) );
  XOR U26336 ( .A(n26422), .B(n26423), .Z(n26410) );
  AND U26337 ( .A(n26424), .B(n26425), .Z(n26423) );
  XOR U26338 ( .A(n26422), .B(n22789), .Z(n26425) );
  XOR U26339 ( .A(n26426), .B(n26427), .Z(n22789) );
  AND U26340 ( .A(n534), .B(n26428), .Z(n26427) );
  XOR U26341 ( .A(n26429), .B(n26426), .Z(n26428) );
  XNOR U26342 ( .A(n22786), .B(n26422), .Z(n26424) );
  XOR U26343 ( .A(n26430), .B(n26431), .Z(n22786) );
  AND U26344 ( .A(n531), .B(n26432), .Z(n26431) );
  XOR U26345 ( .A(n26433), .B(n26430), .Z(n26432) );
  XOR U26346 ( .A(n26434), .B(n26435), .Z(n26422) );
  AND U26347 ( .A(n26436), .B(n26437), .Z(n26435) );
  XOR U26348 ( .A(n26434), .B(n22801), .Z(n26437) );
  XOR U26349 ( .A(n26438), .B(n26439), .Z(n22801) );
  AND U26350 ( .A(n534), .B(n26440), .Z(n26439) );
  XOR U26351 ( .A(n26441), .B(n26438), .Z(n26440) );
  XNOR U26352 ( .A(n22798), .B(n26434), .Z(n26436) );
  XOR U26353 ( .A(n26442), .B(n26443), .Z(n22798) );
  AND U26354 ( .A(n531), .B(n26444), .Z(n26443) );
  XOR U26355 ( .A(n26445), .B(n26442), .Z(n26444) );
  XOR U26356 ( .A(n26446), .B(n26447), .Z(n26434) );
  AND U26357 ( .A(n26448), .B(n26449), .Z(n26447) );
  XOR U26358 ( .A(n26446), .B(n22813), .Z(n26449) );
  XOR U26359 ( .A(n26450), .B(n26451), .Z(n22813) );
  AND U26360 ( .A(n534), .B(n26452), .Z(n26451) );
  XOR U26361 ( .A(n26453), .B(n26450), .Z(n26452) );
  XNOR U26362 ( .A(n22810), .B(n26446), .Z(n26448) );
  XOR U26363 ( .A(n26454), .B(n26455), .Z(n22810) );
  AND U26364 ( .A(n531), .B(n26456), .Z(n26455) );
  XOR U26365 ( .A(n26457), .B(n26454), .Z(n26456) );
  XOR U26366 ( .A(n26458), .B(n26459), .Z(n26446) );
  AND U26367 ( .A(n26460), .B(n26461), .Z(n26459) );
  XOR U26368 ( .A(n26458), .B(n22825), .Z(n26461) );
  XOR U26369 ( .A(n26462), .B(n26463), .Z(n22825) );
  AND U26370 ( .A(n534), .B(n26464), .Z(n26463) );
  XOR U26371 ( .A(n26465), .B(n26462), .Z(n26464) );
  XNOR U26372 ( .A(n22822), .B(n26458), .Z(n26460) );
  XOR U26373 ( .A(n26466), .B(n26467), .Z(n22822) );
  AND U26374 ( .A(n531), .B(n26468), .Z(n26467) );
  XOR U26375 ( .A(n26469), .B(n26466), .Z(n26468) );
  XOR U26376 ( .A(n26470), .B(n26471), .Z(n26458) );
  AND U26377 ( .A(n26472), .B(n26473), .Z(n26471) );
  XOR U26378 ( .A(n26470), .B(n22837), .Z(n26473) );
  XOR U26379 ( .A(n26474), .B(n26475), .Z(n22837) );
  AND U26380 ( .A(n534), .B(n26476), .Z(n26475) );
  XOR U26381 ( .A(n26477), .B(n26474), .Z(n26476) );
  XNOR U26382 ( .A(n22834), .B(n26470), .Z(n26472) );
  XOR U26383 ( .A(n26478), .B(n26479), .Z(n22834) );
  AND U26384 ( .A(n531), .B(n26480), .Z(n26479) );
  XOR U26385 ( .A(n26481), .B(n26478), .Z(n26480) );
  XOR U26386 ( .A(n26482), .B(n26483), .Z(n26470) );
  AND U26387 ( .A(n26484), .B(n26485), .Z(n26483) );
  XOR U26388 ( .A(n26482), .B(n22849), .Z(n26485) );
  XOR U26389 ( .A(n26486), .B(n26487), .Z(n22849) );
  AND U26390 ( .A(n534), .B(n26488), .Z(n26487) );
  XOR U26391 ( .A(n26489), .B(n26486), .Z(n26488) );
  XNOR U26392 ( .A(n22846), .B(n26482), .Z(n26484) );
  XOR U26393 ( .A(n26490), .B(n26491), .Z(n22846) );
  AND U26394 ( .A(n531), .B(n26492), .Z(n26491) );
  XOR U26395 ( .A(n26493), .B(n26490), .Z(n26492) );
  XOR U26396 ( .A(n26494), .B(n26495), .Z(n26482) );
  AND U26397 ( .A(n26496), .B(n26497), .Z(n26495) );
  XOR U26398 ( .A(n22861), .B(n26494), .Z(n26497) );
  XOR U26399 ( .A(n26498), .B(n26499), .Z(n22861) );
  AND U26400 ( .A(n534), .B(n26500), .Z(n26499) );
  XOR U26401 ( .A(n26498), .B(n26501), .Z(n26500) );
  XNOR U26402 ( .A(n26494), .B(n22858), .Z(n26496) );
  XOR U26403 ( .A(n26502), .B(n26503), .Z(n22858) );
  AND U26404 ( .A(n531), .B(n26504), .Z(n26503) );
  XOR U26405 ( .A(n26502), .B(n26505), .Z(n26504) );
  XOR U26406 ( .A(n26506), .B(n26507), .Z(n26494) );
  AND U26407 ( .A(n26508), .B(n26509), .Z(n26507) );
  XNOR U26408 ( .A(n26510), .B(n22874), .Z(n26509) );
  XOR U26409 ( .A(n26511), .B(n26512), .Z(n22874) );
  AND U26410 ( .A(n534), .B(n26513), .Z(n26512) );
  XOR U26411 ( .A(n26514), .B(n26511), .Z(n26513) );
  XNOR U26412 ( .A(n22871), .B(n26506), .Z(n26508) );
  XOR U26413 ( .A(n26515), .B(n26516), .Z(n22871) );
  AND U26414 ( .A(n531), .B(n26517), .Z(n26516) );
  XOR U26415 ( .A(n26518), .B(n26515), .Z(n26517) );
  IV U26416 ( .A(n26510), .Z(n26506) );
  AND U26417 ( .A(n26142), .B(n26145), .Z(n26510) );
  XNOR U26418 ( .A(n26519), .B(n26520), .Z(n26145) );
  AND U26419 ( .A(n534), .B(n26521), .Z(n26520) );
  XNOR U26420 ( .A(n26522), .B(n26519), .Z(n26521) );
  XOR U26421 ( .A(n26523), .B(n26524), .Z(n534) );
  AND U26422 ( .A(n26525), .B(n26526), .Z(n26524) );
  XOR U26423 ( .A(n26523), .B(n26153), .Z(n26526) );
  XNOR U26424 ( .A(n26527), .B(n26528), .Z(n26153) );
  AND U26425 ( .A(n26529), .B(n406), .Z(n26528) );
  AND U26426 ( .A(n26527), .B(n26530), .Z(n26529) );
  XNOR U26427 ( .A(n26150), .B(n26523), .Z(n26525) );
  XOR U26428 ( .A(n26531), .B(n26532), .Z(n26150) );
  AND U26429 ( .A(n26533), .B(n404), .Z(n26532) );
  NOR U26430 ( .A(n26531), .B(n26534), .Z(n26533) );
  XOR U26431 ( .A(n26535), .B(n26536), .Z(n26523) );
  AND U26432 ( .A(n26537), .B(n26538), .Z(n26536) );
  XOR U26433 ( .A(n26535), .B(n26165), .Z(n26538) );
  XOR U26434 ( .A(n26539), .B(n26540), .Z(n26165) );
  AND U26435 ( .A(n406), .B(n26541), .Z(n26540) );
  XOR U26436 ( .A(n26542), .B(n26539), .Z(n26541) );
  XNOR U26437 ( .A(n26162), .B(n26535), .Z(n26537) );
  XOR U26438 ( .A(n26543), .B(n26544), .Z(n26162) );
  AND U26439 ( .A(n404), .B(n26545), .Z(n26544) );
  XOR U26440 ( .A(n26546), .B(n26543), .Z(n26545) );
  XOR U26441 ( .A(n26547), .B(n26548), .Z(n26535) );
  AND U26442 ( .A(n26549), .B(n26550), .Z(n26548) );
  XOR U26443 ( .A(n26547), .B(n26177), .Z(n26550) );
  XOR U26444 ( .A(n26551), .B(n26552), .Z(n26177) );
  AND U26445 ( .A(n406), .B(n26553), .Z(n26552) );
  XOR U26446 ( .A(n26554), .B(n26551), .Z(n26553) );
  XNOR U26447 ( .A(n26174), .B(n26547), .Z(n26549) );
  XOR U26448 ( .A(n26555), .B(n26556), .Z(n26174) );
  AND U26449 ( .A(n404), .B(n26557), .Z(n26556) );
  XOR U26450 ( .A(n26558), .B(n26555), .Z(n26557) );
  XOR U26451 ( .A(n26559), .B(n26560), .Z(n26547) );
  AND U26452 ( .A(n26561), .B(n26562), .Z(n26560) );
  XOR U26453 ( .A(n26559), .B(n26189), .Z(n26562) );
  XOR U26454 ( .A(n26563), .B(n26564), .Z(n26189) );
  AND U26455 ( .A(n406), .B(n26565), .Z(n26564) );
  XOR U26456 ( .A(n26566), .B(n26563), .Z(n26565) );
  XNOR U26457 ( .A(n26186), .B(n26559), .Z(n26561) );
  XOR U26458 ( .A(n26567), .B(n26568), .Z(n26186) );
  AND U26459 ( .A(n404), .B(n26569), .Z(n26568) );
  XOR U26460 ( .A(n26570), .B(n26567), .Z(n26569) );
  XOR U26461 ( .A(n26571), .B(n26572), .Z(n26559) );
  AND U26462 ( .A(n26573), .B(n26574), .Z(n26572) );
  XOR U26463 ( .A(n26571), .B(n26201), .Z(n26574) );
  XOR U26464 ( .A(n26575), .B(n26576), .Z(n26201) );
  AND U26465 ( .A(n406), .B(n26577), .Z(n26576) );
  XOR U26466 ( .A(n26578), .B(n26575), .Z(n26577) );
  XNOR U26467 ( .A(n26198), .B(n26571), .Z(n26573) );
  XOR U26468 ( .A(n26579), .B(n26580), .Z(n26198) );
  AND U26469 ( .A(n404), .B(n26581), .Z(n26580) );
  XOR U26470 ( .A(n26582), .B(n26579), .Z(n26581) );
  XOR U26471 ( .A(n26583), .B(n26584), .Z(n26571) );
  AND U26472 ( .A(n26585), .B(n26586), .Z(n26584) );
  XOR U26473 ( .A(n26583), .B(n26213), .Z(n26586) );
  XOR U26474 ( .A(n26587), .B(n26588), .Z(n26213) );
  AND U26475 ( .A(n406), .B(n26589), .Z(n26588) );
  XOR U26476 ( .A(n26590), .B(n26587), .Z(n26589) );
  XNOR U26477 ( .A(n26210), .B(n26583), .Z(n26585) );
  XOR U26478 ( .A(n26591), .B(n26592), .Z(n26210) );
  AND U26479 ( .A(n404), .B(n26593), .Z(n26592) );
  XOR U26480 ( .A(n26594), .B(n26591), .Z(n26593) );
  XOR U26481 ( .A(n26595), .B(n26596), .Z(n26583) );
  AND U26482 ( .A(n26597), .B(n26598), .Z(n26596) );
  XOR U26483 ( .A(n26595), .B(n26225), .Z(n26598) );
  XOR U26484 ( .A(n26599), .B(n26600), .Z(n26225) );
  AND U26485 ( .A(n406), .B(n26601), .Z(n26600) );
  XOR U26486 ( .A(n26602), .B(n26599), .Z(n26601) );
  XNOR U26487 ( .A(n26222), .B(n26595), .Z(n26597) );
  XOR U26488 ( .A(n26603), .B(n26604), .Z(n26222) );
  AND U26489 ( .A(n404), .B(n26605), .Z(n26604) );
  XOR U26490 ( .A(n26606), .B(n26603), .Z(n26605) );
  XOR U26491 ( .A(n26607), .B(n26608), .Z(n26595) );
  AND U26492 ( .A(n26609), .B(n26610), .Z(n26608) );
  XOR U26493 ( .A(n26607), .B(n26237), .Z(n26610) );
  XOR U26494 ( .A(n26611), .B(n26612), .Z(n26237) );
  AND U26495 ( .A(n406), .B(n26613), .Z(n26612) );
  XOR U26496 ( .A(n26614), .B(n26611), .Z(n26613) );
  XNOR U26497 ( .A(n26234), .B(n26607), .Z(n26609) );
  XOR U26498 ( .A(n26615), .B(n26616), .Z(n26234) );
  AND U26499 ( .A(n404), .B(n26617), .Z(n26616) );
  XOR U26500 ( .A(n26618), .B(n26615), .Z(n26617) );
  XOR U26501 ( .A(n26619), .B(n26620), .Z(n26607) );
  AND U26502 ( .A(n26621), .B(n26622), .Z(n26620) );
  XOR U26503 ( .A(n26619), .B(n26249), .Z(n26622) );
  XOR U26504 ( .A(n26623), .B(n26624), .Z(n26249) );
  AND U26505 ( .A(n406), .B(n26625), .Z(n26624) );
  XOR U26506 ( .A(n26626), .B(n26623), .Z(n26625) );
  XNOR U26507 ( .A(n26246), .B(n26619), .Z(n26621) );
  XOR U26508 ( .A(n26627), .B(n26628), .Z(n26246) );
  AND U26509 ( .A(n404), .B(n26629), .Z(n26628) );
  XOR U26510 ( .A(n26630), .B(n26627), .Z(n26629) );
  XOR U26511 ( .A(n26631), .B(n26632), .Z(n26619) );
  AND U26512 ( .A(n26633), .B(n26634), .Z(n26632) );
  XOR U26513 ( .A(n26631), .B(n26261), .Z(n26634) );
  XOR U26514 ( .A(n26635), .B(n26636), .Z(n26261) );
  AND U26515 ( .A(n406), .B(n26637), .Z(n26636) );
  XOR U26516 ( .A(n26638), .B(n26635), .Z(n26637) );
  XNOR U26517 ( .A(n26258), .B(n26631), .Z(n26633) );
  XOR U26518 ( .A(n26639), .B(n26640), .Z(n26258) );
  AND U26519 ( .A(n404), .B(n26641), .Z(n26640) );
  XOR U26520 ( .A(n26642), .B(n26639), .Z(n26641) );
  XOR U26521 ( .A(n26643), .B(n26644), .Z(n26631) );
  AND U26522 ( .A(n26645), .B(n26646), .Z(n26644) );
  XOR U26523 ( .A(n26643), .B(n26273), .Z(n26646) );
  XOR U26524 ( .A(n26647), .B(n26648), .Z(n26273) );
  AND U26525 ( .A(n406), .B(n26649), .Z(n26648) );
  XOR U26526 ( .A(n26650), .B(n26647), .Z(n26649) );
  XNOR U26527 ( .A(n26270), .B(n26643), .Z(n26645) );
  XOR U26528 ( .A(n26651), .B(n26652), .Z(n26270) );
  AND U26529 ( .A(n404), .B(n26653), .Z(n26652) );
  XOR U26530 ( .A(n26654), .B(n26651), .Z(n26653) );
  XOR U26531 ( .A(n26655), .B(n26656), .Z(n26643) );
  AND U26532 ( .A(n26657), .B(n26658), .Z(n26656) );
  XOR U26533 ( .A(n26655), .B(n26285), .Z(n26658) );
  XOR U26534 ( .A(n26659), .B(n26660), .Z(n26285) );
  AND U26535 ( .A(n406), .B(n26661), .Z(n26660) );
  XOR U26536 ( .A(n26662), .B(n26659), .Z(n26661) );
  XNOR U26537 ( .A(n26282), .B(n26655), .Z(n26657) );
  XOR U26538 ( .A(n26663), .B(n26664), .Z(n26282) );
  AND U26539 ( .A(n404), .B(n26665), .Z(n26664) );
  XOR U26540 ( .A(n26666), .B(n26663), .Z(n26665) );
  XOR U26541 ( .A(n26667), .B(n26668), .Z(n26655) );
  AND U26542 ( .A(n26669), .B(n26670), .Z(n26668) );
  XOR U26543 ( .A(n26667), .B(n26297), .Z(n26670) );
  XOR U26544 ( .A(n26671), .B(n26672), .Z(n26297) );
  AND U26545 ( .A(n406), .B(n26673), .Z(n26672) );
  XOR U26546 ( .A(n26674), .B(n26671), .Z(n26673) );
  XNOR U26547 ( .A(n26294), .B(n26667), .Z(n26669) );
  XOR U26548 ( .A(n26675), .B(n26676), .Z(n26294) );
  AND U26549 ( .A(n404), .B(n26677), .Z(n26676) );
  XOR U26550 ( .A(n26678), .B(n26675), .Z(n26677) );
  XOR U26551 ( .A(n26679), .B(n26680), .Z(n26667) );
  AND U26552 ( .A(n26681), .B(n26682), .Z(n26680) );
  XOR U26553 ( .A(n26679), .B(n26309), .Z(n26682) );
  XOR U26554 ( .A(n26683), .B(n26684), .Z(n26309) );
  AND U26555 ( .A(n406), .B(n26685), .Z(n26684) );
  XOR U26556 ( .A(n26686), .B(n26683), .Z(n26685) );
  XNOR U26557 ( .A(n26306), .B(n26679), .Z(n26681) );
  XOR U26558 ( .A(n26687), .B(n26688), .Z(n26306) );
  AND U26559 ( .A(n404), .B(n26689), .Z(n26688) );
  XOR U26560 ( .A(n26690), .B(n26687), .Z(n26689) );
  XOR U26561 ( .A(n26691), .B(n26692), .Z(n26679) );
  AND U26562 ( .A(n26693), .B(n26694), .Z(n26692) );
  XOR U26563 ( .A(n26691), .B(n26321), .Z(n26694) );
  XOR U26564 ( .A(n26695), .B(n26696), .Z(n26321) );
  AND U26565 ( .A(n406), .B(n26697), .Z(n26696) );
  XOR U26566 ( .A(n26698), .B(n26695), .Z(n26697) );
  XNOR U26567 ( .A(n26318), .B(n26691), .Z(n26693) );
  XOR U26568 ( .A(n26699), .B(n26700), .Z(n26318) );
  AND U26569 ( .A(n404), .B(n26701), .Z(n26700) );
  XOR U26570 ( .A(n26702), .B(n26699), .Z(n26701) );
  XOR U26571 ( .A(n26703), .B(n26704), .Z(n26691) );
  AND U26572 ( .A(n26705), .B(n26706), .Z(n26704) );
  XOR U26573 ( .A(n26703), .B(n26333), .Z(n26706) );
  XOR U26574 ( .A(n26707), .B(n26708), .Z(n26333) );
  AND U26575 ( .A(n406), .B(n26709), .Z(n26708) );
  XOR U26576 ( .A(n26710), .B(n26707), .Z(n26709) );
  XNOR U26577 ( .A(n26330), .B(n26703), .Z(n26705) );
  XOR U26578 ( .A(n26711), .B(n26712), .Z(n26330) );
  AND U26579 ( .A(n404), .B(n26713), .Z(n26712) );
  XOR U26580 ( .A(n26714), .B(n26711), .Z(n26713) );
  XOR U26581 ( .A(n26715), .B(n26716), .Z(n26703) );
  AND U26582 ( .A(n26717), .B(n26718), .Z(n26716) );
  XOR U26583 ( .A(n26715), .B(n26345), .Z(n26718) );
  XOR U26584 ( .A(n26719), .B(n26720), .Z(n26345) );
  AND U26585 ( .A(n406), .B(n26721), .Z(n26720) );
  XOR U26586 ( .A(n26722), .B(n26719), .Z(n26721) );
  XNOR U26587 ( .A(n26342), .B(n26715), .Z(n26717) );
  XOR U26588 ( .A(n26723), .B(n26724), .Z(n26342) );
  AND U26589 ( .A(n404), .B(n26725), .Z(n26724) );
  XOR U26590 ( .A(n26726), .B(n26723), .Z(n26725) );
  XOR U26591 ( .A(n26727), .B(n26728), .Z(n26715) );
  AND U26592 ( .A(n26729), .B(n26730), .Z(n26728) );
  XOR U26593 ( .A(n26727), .B(n26357), .Z(n26730) );
  XOR U26594 ( .A(n26731), .B(n26732), .Z(n26357) );
  AND U26595 ( .A(n406), .B(n26733), .Z(n26732) );
  XOR U26596 ( .A(n26734), .B(n26731), .Z(n26733) );
  XNOR U26597 ( .A(n26354), .B(n26727), .Z(n26729) );
  XOR U26598 ( .A(n26735), .B(n26736), .Z(n26354) );
  AND U26599 ( .A(n404), .B(n26737), .Z(n26736) );
  XOR U26600 ( .A(n26738), .B(n26735), .Z(n26737) );
  XOR U26601 ( .A(n26739), .B(n26740), .Z(n26727) );
  AND U26602 ( .A(n26741), .B(n26742), .Z(n26740) );
  XOR U26603 ( .A(n26739), .B(n26369), .Z(n26742) );
  XOR U26604 ( .A(n26743), .B(n26744), .Z(n26369) );
  AND U26605 ( .A(n406), .B(n26745), .Z(n26744) );
  XOR U26606 ( .A(n26746), .B(n26743), .Z(n26745) );
  XNOR U26607 ( .A(n26366), .B(n26739), .Z(n26741) );
  XOR U26608 ( .A(n26747), .B(n26748), .Z(n26366) );
  AND U26609 ( .A(n404), .B(n26749), .Z(n26748) );
  XOR U26610 ( .A(n26750), .B(n26747), .Z(n26749) );
  XOR U26611 ( .A(n26751), .B(n26752), .Z(n26739) );
  AND U26612 ( .A(n26753), .B(n26754), .Z(n26752) );
  XOR U26613 ( .A(n26751), .B(n26381), .Z(n26754) );
  XOR U26614 ( .A(n26755), .B(n26756), .Z(n26381) );
  AND U26615 ( .A(n406), .B(n26757), .Z(n26756) );
  XOR U26616 ( .A(n26758), .B(n26755), .Z(n26757) );
  XNOR U26617 ( .A(n26378), .B(n26751), .Z(n26753) );
  XOR U26618 ( .A(n26759), .B(n26760), .Z(n26378) );
  AND U26619 ( .A(n404), .B(n26761), .Z(n26760) );
  XOR U26620 ( .A(n26762), .B(n26759), .Z(n26761) );
  XOR U26621 ( .A(n26763), .B(n26764), .Z(n26751) );
  AND U26622 ( .A(n26765), .B(n26766), .Z(n26764) );
  XOR U26623 ( .A(n26763), .B(n26393), .Z(n26766) );
  XOR U26624 ( .A(n26767), .B(n26768), .Z(n26393) );
  AND U26625 ( .A(n406), .B(n26769), .Z(n26768) );
  XOR U26626 ( .A(n26770), .B(n26767), .Z(n26769) );
  XNOR U26627 ( .A(n26390), .B(n26763), .Z(n26765) );
  XOR U26628 ( .A(n26771), .B(n26772), .Z(n26390) );
  AND U26629 ( .A(n404), .B(n26773), .Z(n26772) );
  XOR U26630 ( .A(n26774), .B(n26771), .Z(n26773) );
  XOR U26631 ( .A(n26775), .B(n26776), .Z(n26763) );
  AND U26632 ( .A(n26777), .B(n26778), .Z(n26776) );
  XOR U26633 ( .A(n26775), .B(n26405), .Z(n26778) );
  XOR U26634 ( .A(n26779), .B(n26780), .Z(n26405) );
  AND U26635 ( .A(n406), .B(n26781), .Z(n26780) );
  XOR U26636 ( .A(n26782), .B(n26779), .Z(n26781) );
  XNOR U26637 ( .A(n26402), .B(n26775), .Z(n26777) );
  XOR U26638 ( .A(n26783), .B(n26784), .Z(n26402) );
  AND U26639 ( .A(n404), .B(n26785), .Z(n26784) );
  XOR U26640 ( .A(n26786), .B(n26783), .Z(n26785) );
  XOR U26641 ( .A(n26787), .B(n26788), .Z(n26775) );
  AND U26642 ( .A(n26789), .B(n26790), .Z(n26788) );
  XOR U26643 ( .A(n26787), .B(n26417), .Z(n26790) );
  XOR U26644 ( .A(n26791), .B(n26792), .Z(n26417) );
  AND U26645 ( .A(n406), .B(n26793), .Z(n26792) );
  XOR U26646 ( .A(n26794), .B(n26791), .Z(n26793) );
  XNOR U26647 ( .A(n26414), .B(n26787), .Z(n26789) );
  XOR U26648 ( .A(n26795), .B(n26796), .Z(n26414) );
  AND U26649 ( .A(n404), .B(n26797), .Z(n26796) );
  XOR U26650 ( .A(n26798), .B(n26795), .Z(n26797) );
  XOR U26651 ( .A(n26799), .B(n26800), .Z(n26787) );
  AND U26652 ( .A(n26801), .B(n26802), .Z(n26800) );
  XOR U26653 ( .A(n26799), .B(n26429), .Z(n26802) );
  XOR U26654 ( .A(n26803), .B(n26804), .Z(n26429) );
  AND U26655 ( .A(n406), .B(n26805), .Z(n26804) );
  XOR U26656 ( .A(n26806), .B(n26803), .Z(n26805) );
  XNOR U26657 ( .A(n26426), .B(n26799), .Z(n26801) );
  XOR U26658 ( .A(n26807), .B(n26808), .Z(n26426) );
  AND U26659 ( .A(n404), .B(n26809), .Z(n26808) );
  XOR U26660 ( .A(n26810), .B(n26807), .Z(n26809) );
  XOR U26661 ( .A(n26811), .B(n26812), .Z(n26799) );
  AND U26662 ( .A(n26813), .B(n26814), .Z(n26812) );
  XOR U26663 ( .A(n26811), .B(n26441), .Z(n26814) );
  XOR U26664 ( .A(n26815), .B(n26816), .Z(n26441) );
  AND U26665 ( .A(n406), .B(n26817), .Z(n26816) );
  XOR U26666 ( .A(n26818), .B(n26815), .Z(n26817) );
  XNOR U26667 ( .A(n26438), .B(n26811), .Z(n26813) );
  XOR U26668 ( .A(n26819), .B(n26820), .Z(n26438) );
  AND U26669 ( .A(n404), .B(n26821), .Z(n26820) );
  XOR U26670 ( .A(n26822), .B(n26819), .Z(n26821) );
  XOR U26671 ( .A(n26823), .B(n26824), .Z(n26811) );
  AND U26672 ( .A(n26825), .B(n26826), .Z(n26824) );
  XOR U26673 ( .A(n26823), .B(n26453), .Z(n26826) );
  XOR U26674 ( .A(n26827), .B(n26828), .Z(n26453) );
  AND U26675 ( .A(n406), .B(n26829), .Z(n26828) );
  XOR U26676 ( .A(n26830), .B(n26827), .Z(n26829) );
  XNOR U26677 ( .A(n26450), .B(n26823), .Z(n26825) );
  XOR U26678 ( .A(n26831), .B(n26832), .Z(n26450) );
  AND U26679 ( .A(n404), .B(n26833), .Z(n26832) );
  XOR U26680 ( .A(n26834), .B(n26831), .Z(n26833) );
  XOR U26681 ( .A(n26835), .B(n26836), .Z(n26823) );
  AND U26682 ( .A(n26837), .B(n26838), .Z(n26836) );
  XOR U26683 ( .A(n26835), .B(n26465), .Z(n26838) );
  XOR U26684 ( .A(n26839), .B(n26840), .Z(n26465) );
  AND U26685 ( .A(n406), .B(n26841), .Z(n26840) );
  XOR U26686 ( .A(n26842), .B(n26839), .Z(n26841) );
  XNOR U26687 ( .A(n26462), .B(n26835), .Z(n26837) );
  XOR U26688 ( .A(n26843), .B(n26844), .Z(n26462) );
  AND U26689 ( .A(n404), .B(n26845), .Z(n26844) );
  XOR U26690 ( .A(n26846), .B(n26843), .Z(n26845) );
  XOR U26691 ( .A(n26847), .B(n26848), .Z(n26835) );
  AND U26692 ( .A(n26849), .B(n26850), .Z(n26848) );
  XOR U26693 ( .A(n26847), .B(n26477), .Z(n26850) );
  XOR U26694 ( .A(n26851), .B(n26852), .Z(n26477) );
  AND U26695 ( .A(n406), .B(n26853), .Z(n26852) );
  XOR U26696 ( .A(n26854), .B(n26851), .Z(n26853) );
  XNOR U26697 ( .A(n26474), .B(n26847), .Z(n26849) );
  XOR U26698 ( .A(n26855), .B(n26856), .Z(n26474) );
  AND U26699 ( .A(n404), .B(n26857), .Z(n26856) );
  XOR U26700 ( .A(n26858), .B(n26855), .Z(n26857) );
  XOR U26701 ( .A(n26859), .B(n26860), .Z(n26847) );
  AND U26702 ( .A(n26861), .B(n26862), .Z(n26860) );
  XOR U26703 ( .A(n26859), .B(n26489), .Z(n26862) );
  XOR U26704 ( .A(n26863), .B(n26864), .Z(n26489) );
  AND U26705 ( .A(n406), .B(n26865), .Z(n26864) );
  XOR U26706 ( .A(n26866), .B(n26863), .Z(n26865) );
  XNOR U26707 ( .A(n26486), .B(n26859), .Z(n26861) );
  XOR U26708 ( .A(n26867), .B(n26868), .Z(n26486) );
  AND U26709 ( .A(n404), .B(n26869), .Z(n26868) );
  XOR U26710 ( .A(n26870), .B(n26867), .Z(n26869) );
  XOR U26711 ( .A(n26871), .B(n26872), .Z(n26859) );
  AND U26712 ( .A(n26873), .B(n26874), .Z(n26872) );
  XOR U26713 ( .A(n26501), .B(n26871), .Z(n26874) );
  XOR U26714 ( .A(n26875), .B(n26876), .Z(n26501) );
  AND U26715 ( .A(n406), .B(n26877), .Z(n26876) );
  XOR U26716 ( .A(n26875), .B(n26878), .Z(n26877) );
  XNOR U26717 ( .A(n26871), .B(n26498), .Z(n26873) );
  XOR U26718 ( .A(n26879), .B(n26880), .Z(n26498) );
  AND U26719 ( .A(n404), .B(n26881), .Z(n26880) );
  XOR U26720 ( .A(n26879), .B(n26882), .Z(n26881) );
  XOR U26721 ( .A(n26883), .B(n26884), .Z(n26871) );
  AND U26722 ( .A(n26885), .B(n26886), .Z(n26884) );
  XNOR U26723 ( .A(n26887), .B(n26514), .Z(n26886) );
  XOR U26724 ( .A(n26888), .B(n26889), .Z(n26514) );
  AND U26725 ( .A(n406), .B(n26890), .Z(n26889) );
  XOR U26726 ( .A(n26891), .B(n26888), .Z(n26890) );
  XNOR U26727 ( .A(n26511), .B(n26883), .Z(n26885) );
  XOR U26728 ( .A(n26892), .B(n26893), .Z(n26511) );
  AND U26729 ( .A(n404), .B(n26894), .Z(n26893) );
  XOR U26730 ( .A(n26895), .B(n26892), .Z(n26894) );
  IV U26731 ( .A(n26887), .Z(n26883) );
  AND U26732 ( .A(n26519), .B(n26522), .Z(n26887) );
  XNOR U26733 ( .A(n26896), .B(n26897), .Z(n26522) );
  AND U26734 ( .A(n406), .B(n26898), .Z(n26897) );
  XNOR U26735 ( .A(n26899), .B(n26896), .Z(n26898) );
  XOR U26736 ( .A(n26900), .B(n26901), .Z(n406) );
  AND U26737 ( .A(n26902), .B(n26903), .Z(n26901) );
  XOR U26738 ( .A(n26530), .B(n26900), .Z(n26903) );
  IV U26739 ( .A(n26904), .Z(n26530) );
  AND U26740 ( .A(p_input[511]), .B(p_input[479]), .Z(n26904) );
  XOR U26741 ( .A(n26900), .B(n26527), .Z(n26902) );
  AND U26742 ( .A(p_input[415]), .B(p_input[447]), .Z(n26527) );
  XOR U26743 ( .A(n26905), .B(n26906), .Z(n26900) );
  AND U26744 ( .A(n26907), .B(n26908), .Z(n26906) );
  XOR U26745 ( .A(n26905), .B(n26542), .Z(n26908) );
  XNOR U26746 ( .A(p_input[478]), .B(n26909), .Z(n26542) );
  AND U26747 ( .A(n606), .B(n26910), .Z(n26909) );
  XOR U26748 ( .A(p_input[510]), .B(p_input[478]), .Z(n26910) );
  XNOR U26749 ( .A(n26539), .B(n26905), .Z(n26907) );
  XOR U26750 ( .A(n26911), .B(n26912), .Z(n26539) );
  AND U26751 ( .A(n604), .B(n26913), .Z(n26912) );
  XOR U26752 ( .A(p_input[446]), .B(p_input[414]), .Z(n26913) );
  XOR U26753 ( .A(n26914), .B(n26915), .Z(n26905) );
  AND U26754 ( .A(n26916), .B(n26917), .Z(n26915) );
  XOR U26755 ( .A(n26914), .B(n26554), .Z(n26917) );
  XNOR U26756 ( .A(p_input[477]), .B(n26918), .Z(n26554) );
  AND U26757 ( .A(n606), .B(n26919), .Z(n26918) );
  XOR U26758 ( .A(p_input[509]), .B(p_input[477]), .Z(n26919) );
  XNOR U26759 ( .A(n26551), .B(n26914), .Z(n26916) );
  XOR U26760 ( .A(n26920), .B(n26921), .Z(n26551) );
  AND U26761 ( .A(n604), .B(n26922), .Z(n26921) );
  XOR U26762 ( .A(p_input[445]), .B(p_input[413]), .Z(n26922) );
  XOR U26763 ( .A(n26923), .B(n26924), .Z(n26914) );
  AND U26764 ( .A(n26925), .B(n26926), .Z(n26924) );
  XOR U26765 ( .A(n26923), .B(n26566), .Z(n26926) );
  XNOR U26766 ( .A(p_input[476]), .B(n26927), .Z(n26566) );
  AND U26767 ( .A(n606), .B(n26928), .Z(n26927) );
  XOR U26768 ( .A(p_input[508]), .B(p_input[476]), .Z(n26928) );
  XNOR U26769 ( .A(n26563), .B(n26923), .Z(n26925) );
  XOR U26770 ( .A(n26929), .B(n26930), .Z(n26563) );
  AND U26771 ( .A(n604), .B(n26931), .Z(n26930) );
  XOR U26772 ( .A(p_input[444]), .B(p_input[412]), .Z(n26931) );
  XOR U26773 ( .A(n26932), .B(n26933), .Z(n26923) );
  AND U26774 ( .A(n26934), .B(n26935), .Z(n26933) );
  XOR U26775 ( .A(n26932), .B(n26578), .Z(n26935) );
  XNOR U26776 ( .A(p_input[475]), .B(n26936), .Z(n26578) );
  AND U26777 ( .A(n606), .B(n26937), .Z(n26936) );
  XOR U26778 ( .A(p_input[507]), .B(p_input[475]), .Z(n26937) );
  XNOR U26779 ( .A(n26575), .B(n26932), .Z(n26934) );
  XOR U26780 ( .A(n26938), .B(n26939), .Z(n26575) );
  AND U26781 ( .A(n604), .B(n26940), .Z(n26939) );
  XOR U26782 ( .A(p_input[443]), .B(p_input[411]), .Z(n26940) );
  XOR U26783 ( .A(n26941), .B(n26942), .Z(n26932) );
  AND U26784 ( .A(n26943), .B(n26944), .Z(n26942) );
  XOR U26785 ( .A(n26941), .B(n26590), .Z(n26944) );
  XNOR U26786 ( .A(p_input[474]), .B(n26945), .Z(n26590) );
  AND U26787 ( .A(n606), .B(n26946), .Z(n26945) );
  XOR U26788 ( .A(p_input[506]), .B(p_input[474]), .Z(n26946) );
  XNOR U26789 ( .A(n26587), .B(n26941), .Z(n26943) );
  XOR U26790 ( .A(n26947), .B(n26948), .Z(n26587) );
  AND U26791 ( .A(n604), .B(n26949), .Z(n26948) );
  XOR U26792 ( .A(p_input[442]), .B(p_input[410]), .Z(n26949) );
  XOR U26793 ( .A(n26950), .B(n26951), .Z(n26941) );
  AND U26794 ( .A(n26952), .B(n26953), .Z(n26951) );
  XOR U26795 ( .A(n26950), .B(n26602), .Z(n26953) );
  XNOR U26796 ( .A(p_input[473]), .B(n26954), .Z(n26602) );
  AND U26797 ( .A(n606), .B(n26955), .Z(n26954) );
  XOR U26798 ( .A(p_input[505]), .B(p_input[473]), .Z(n26955) );
  XNOR U26799 ( .A(n26599), .B(n26950), .Z(n26952) );
  XOR U26800 ( .A(n26956), .B(n26957), .Z(n26599) );
  AND U26801 ( .A(n604), .B(n26958), .Z(n26957) );
  XOR U26802 ( .A(p_input[441]), .B(p_input[409]), .Z(n26958) );
  XOR U26803 ( .A(n26959), .B(n26960), .Z(n26950) );
  AND U26804 ( .A(n26961), .B(n26962), .Z(n26960) );
  XOR U26805 ( .A(n26959), .B(n26614), .Z(n26962) );
  XNOR U26806 ( .A(p_input[472]), .B(n26963), .Z(n26614) );
  AND U26807 ( .A(n606), .B(n26964), .Z(n26963) );
  XOR U26808 ( .A(p_input[504]), .B(p_input[472]), .Z(n26964) );
  XNOR U26809 ( .A(n26611), .B(n26959), .Z(n26961) );
  XOR U26810 ( .A(n26965), .B(n26966), .Z(n26611) );
  AND U26811 ( .A(n604), .B(n26967), .Z(n26966) );
  XOR U26812 ( .A(p_input[440]), .B(p_input[408]), .Z(n26967) );
  XOR U26813 ( .A(n26968), .B(n26969), .Z(n26959) );
  AND U26814 ( .A(n26970), .B(n26971), .Z(n26969) );
  XOR U26815 ( .A(n26968), .B(n26626), .Z(n26971) );
  XNOR U26816 ( .A(p_input[471]), .B(n26972), .Z(n26626) );
  AND U26817 ( .A(n606), .B(n26973), .Z(n26972) );
  XOR U26818 ( .A(p_input[503]), .B(p_input[471]), .Z(n26973) );
  XNOR U26819 ( .A(n26623), .B(n26968), .Z(n26970) );
  XOR U26820 ( .A(n26974), .B(n26975), .Z(n26623) );
  AND U26821 ( .A(n604), .B(n26976), .Z(n26975) );
  XOR U26822 ( .A(p_input[439]), .B(p_input[407]), .Z(n26976) );
  XOR U26823 ( .A(n26977), .B(n26978), .Z(n26968) );
  AND U26824 ( .A(n26979), .B(n26980), .Z(n26978) );
  XOR U26825 ( .A(n26977), .B(n26638), .Z(n26980) );
  XNOR U26826 ( .A(p_input[470]), .B(n26981), .Z(n26638) );
  AND U26827 ( .A(n606), .B(n26982), .Z(n26981) );
  XOR U26828 ( .A(p_input[502]), .B(p_input[470]), .Z(n26982) );
  XNOR U26829 ( .A(n26635), .B(n26977), .Z(n26979) );
  XOR U26830 ( .A(n26983), .B(n26984), .Z(n26635) );
  AND U26831 ( .A(n604), .B(n26985), .Z(n26984) );
  XOR U26832 ( .A(p_input[438]), .B(p_input[406]), .Z(n26985) );
  XOR U26833 ( .A(n26986), .B(n26987), .Z(n26977) );
  AND U26834 ( .A(n26988), .B(n26989), .Z(n26987) );
  XOR U26835 ( .A(n26986), .B(n26650), .Z(n26989) );
  XNOR U26836 ( .A(p_input[469]), .B(n26990), .Z(n26650) );
  AND U26837 ( .A(n606), .B(n26991), .Z(n26990) );
  XOR U26838 ( .A(p_input[501]), .B(p_input[469]), .Z(n26991) );
  XNOR U26839 ( .A(n26647), .B(n26986), .Z(n26988) );
  XOR U26840 ( .A(n26992), .B(n26993), .Z(n26647) );
  AND U26841 ( .A(n604), .B(n26994), .Z(n26993) );
  XOR U26842 ( .A(p_input[437]), .B(p_input[405]), .Z(n26994) );
  XOR U26843 ( .A(n26995), .B(n26996), .Z(n26986) );
  AND U26844 ( .A(n26997), .B(n26998), .Z(n26996) );
  XOR U26845 ( .A(n26995), .B(n26662), .Z(n26998) );
  XNOR U26846 ( .A(p_input[468]), .B(n26999), .Z(n26662) );
  AND U26847 ( .A(n606), .B(n27000), .Z(n26999) );
  XOR U26848 ( .A(p_input[500]), .B(p_input[468]), .Z(n27000) );
  XNOR U26849 ( .A(n26659), .B(n26995), .Z(n26997) );
  XOR U26850 ( .A(n27001), .B(n27002), .Z(n26659) );
  AND U26851 ( .A(n604), .B(n27003), .Z(n27002) );
  XOR U26852 ( .A(p_input[436]), .B(p_input[404]), .Z(n27003) );
  XOR U26853 ( .A(n27004), .B(n27005), .Z(n26995) );
  AND U26854 ( .A(n27006), .B(n27007), .Z(n27005) );
  XOR U26855 ( .A(n27004), .B(n26674), .Z(n27007) );
  XNOR U26856 ( .A(p_input[467]), .B(n27008), .Z(n26674) );
  AND U26857 ( .A(n606), .B(n27009), .Z(n27008) );
  XOR U26858 ( .A(p_input[499]), .B(p_input[467]), .Z(n27009) );
  XNOR U26859 ( .A(n26671), .B(n27004), .Z(n27006) );
  XOR U26860 ( .A(n27010), .B(n27011), .Z(n26671) );
  AND U26861 ( .A(n604), .B(n27012), .Z(n27011) );
  XOR U26862 ( .A(p_input[435]), .B(p_input[403]), .Z(n27012) );
  XOR U26863 ( .A(n27013), .B(n27014), .Z(n27004) );
  AND U26864 ( .A(n27015), .B(n27016), .Z(n27014) );
  XOR U26865 ( .A(n27013), .B(n26686), .Z(n27016) );
  XNOR U26866 ( .A(p_input[466]), .B(n27017), .Z(n26686) );
  AND U26867 ( .A(n606), .B(n27018), .Z(n27017) );
  XOR U26868 ( .A(p_input[498]), .B(p_input[466]), .Z(n27018) );
  XNOR U26869 ( .A(n26683), .B(n27013), .Z(n27015) );
  XOR U26870 ( .A(n27019), .B(n27020), .Z(n26683) );
  AND U26871 ( .A(n604), .B(n27021), .Z(n27020) );
  XOR U26872 ( .A(p_input[434]), .B(p_input[402]), .Z(n27021) );
  XOR U26873 ( .A(n27022), .B(n27023), .Z(n27013) );
  AND U26874 ( .A(n27024), .B(n27025), .Z(n27023) );
  XOR U26875 ( .A(n27022), .B(n26698), .Z(n27025) );
  XNOR U26876 ( .A(p_input[465]), .B(n27026), .Z(n26698) );
  AND U26877 ( .A(n606), .B(n27027), .Z(n27026) );
  XOR U26878 ( .A(p_input[497]), .B(p_input[465]), .Z(n27027) );
  XNOR U26879 ( .A(n26695), .B(n27022), .Z(n27024) );
  XOR U26880 ( .A(n27028), .B(n27029), .Z(n26695) );
  AND U26881 ( .A(n604), .B(n27030), .Z(n27029) );
  XOR U26882 ( .A(p_input[433]), .B(p_input[401]), .Z(n27030) );
  XOR U26883 ( .A(n27031), .B(n27032), .Z(n27022) );
  AND U26884 ( .A(n27033), .B(n27034), .Z(n27032) );
  XOR U26885 ( .A(n27031), .B(n26710), .Z(n27034) );
  XNOR U26886 ( .A(p_input[464]), .B(n27035), .Z(n26710) );
  AND U26887 ( .A(n606), .B(n27036), .Z(n27035) );
  XOR U26888 ( .A(p_input[496]), .B(p_input[464]), .Z(n27036) );
  XNOR U26889 ( .A(n26707), .B(n27031), .Z(n27033) );
  XOR U26890 ( .A(n27037), .B(n27038), .Z(n26707) );
  AND U26891 ( .A(n604), .B(n27039), .Z(n27038) );
  XOR U26892 ( .A(p_input[432]), .B(p_input[400]), .Z(n27039) );
  XOR U26893 ( .A(n27040), .B(n27041), .Z(n27031) );
  AND U26894 ( .A(n27042), .B(n27043), .Z(n27041) );
  XOR U26895 ( .A(n27040), .B(n26722), .Z(n27043) );
  XNOR U26896 ( .A(p_input[463]), .B(n27044), .Z(n26722) );
  AND U26897 ( .A(n606), .B(n27045), .Z(n27044) );
  XOR U26898 ( .A(p_input[495]), .B(p_input[463]), .Z(n27045) );
  XNOR U26899 ( .A(n26719), .B(n27040), .Z(n27042) );
  XOR U26900 ( .A(n27046), .B(n27047), .Z(n26719) );
  AND U26901 ( .A(n604), .B(n27048), .Z(n27047) );
  XOR U26902 ( .A(p_input[431]), .B(p_input[399]), .Z(n27048) );
  XOR U26903 ( .A(n27049), .B(n27050), .Z(n27040) );
  AND U26904 ( .A(n27051), .B(n27052), .Z(n27050) );
  XOR U26905 ( .A(n27049), .B(n26734), .Z(n27052) );
  XNOR U26906 ( .A(p_input[462]), .B(n27053), .Z(n26734) );
  AND U26907 ( .A(n606), .B(n27054), .Z(n27053) );
  XOR U26908 ( .A(p_input[494]), .B(p_input[462]), .Z(n27054) );
  XNOR U26909 ( .A(n26731), .B(n27049), .Z(n27051) );
  XOR U26910 ( .A(n27055), .B(n27056), .Z(n26731) );
  AND U26911 ( .A(n604), .B(n27057), .Z(n27056) );
  XOR U26912 ( .A(p_input[430]), .B(p_input[398]), .Z(n27057) );
  XOR U26913 ( .A(n27058), .B(n27059), .Z(n27049) );
  AND U26914 ( .A(n27060), .B(n27061), .Z(n27059) );
  XOR U26915 ( .A(n27058), .B(n26746), .Z(n27061) );
  XNOR U26916 ( .A(p_input[461]), .B(n27062), .Z(n26746) );
  AND U26917 ( .A(n606), .B(n27063), .Z(n27062) );
  XOR U26918 ( .A(p_input[493]), .B(p_input[461]), .Z(n27063) );
  XNOR U26919 ( .A(n26743), .B(n27058), .Z(n27060) );
  XOR U26920 ( .A(n27064), .B(n27065), .Z(n26743) );
  AND U26921 ( .A(n604), .B(n27066), .Z(n27065) );
  XOR U26922 ( .A(p_input[429]), .B(p_input[397]), .Z(n27066) );
  XOR U26923 ( .A(n27067), .B(n27068), .Z(n27058) );
  AND U26924 ( .A(n27069), .B(n27070), .Z(n27068) );
  XOR U26925 ( .A(n27067), .B(n26758), .Z(n27070) );
  XNOR U26926 ( .A(p_input[460]), .B(n27071), .Z(n26758) );
  AND U26927 ( .A(n606), .B(n27072), .Z(n27071) );
  XOR U26928 ( .A(p_input[492]), .B(p_input[460]), .Z(n27072) );
  XNOR U26929 ( .A(n26755), .B(n27067), .Z(n27069) );
  XOR U26930 ( .A(n27073), .B(n27074), .Z(n26755) );
  AND U26931 ( .A(n604), .B(n27075), .Z(n27074) );
  XOR U26932 ( .A(p_input[428]), .B(p_input[396]), .Z(n27075) );
  XOR U26933 ( .A(n27076), .B(n27077), .Z(n27067) );
  AND U26934 ( .A(n27078), .B(n27079), .Z(n27077) );
  XOR U26935 ( .A(n27076), .B(n26770), .Z(n27079) );
  XNOR U26936 ( .A(p_input[459]), .B(n27080), .Z(n26770) );
  AND U26937 ( .A(n606), .B(n27081), .Z(n27080) );
  XOR U26938 ( .A(p_input[491]), .B(p_input[459]), .Z(n27081) );
  XNOR U26939 ( .A(n26767), .B(n27076), .Z(n27078) );
  XOR U26940 ( .A(n27082), .B(n27083), .Z(n26767) );
  AND U26941 ( .A(n604), .B(n27084), .Z(n27083) );
  XOR U26942 ( .A(p_input[427]), .B(p_input[395]), .Z(n27084) );
  XOR U26943 ( .A(n27085), .B(n27086), .Z(n27076) );
  AND U26944 ( .A(n27087), .B(n27088), .Z(n27086) );
  XOR U26945 ( .A(n27085), .B(n26782), .Z(n27088) );
  XNOR U26946 ( .A(p_input[458]), .B(n27089), .Z(n26782) );
  AND U26947 ( .A(n606), .B(n27090), .Z(n27089) );
  XOR U26948 ( .A(p_input[490]), .B(p_input[458]), .Z(n27090) );
  XNOR U26949 ( .A(n26779), .B(n27085), .Z(n27087) );
  XOR U26950 ( .A(n27091), .B(n27092), .Z(n26779) );
  AND U26951 ( .A(n604), .B(n27093), .Z(n27092) );
  XOR U26952 ( .A(p_input[426]), .B(p_input[394]), .Z(n27093) );
  XOR U26953 ( .A(n27094), .B(n27095), .Z(n27085) );
  AND U26954 ( .A(n27096), .B(n27097), .Z(n27095) );
  XOR U26955 ( .A(n27094), .B(n26794), .Z(n27097) );
  XNOR U26956 ( .A(p_input[457]), .B(n27098), .Z(n26794) );
  AND U26957 ( .A(n606), .B(n27099), .Z(n27098) );
  XOR U26958 ( .A(p_input[489]), .B(p_input[457]), .Z(n27099) );
  XNOR U26959 ( .A(n26791), .B(n27094), .Z(n27096) );
  XOR U26960 ( .A(n27100), .B(n27101), .Z(n26791) );
  AND U26961 ( .A(n604), .B(n27102), .Z(n27101) );
  XOR U26962 ( .A(p_input[425]), .B(p_input[393]), .Z(n27102) );
  XOR U26963 ( .A(n27103), .B(n27104), .Z(n27094) );
  AND U26964 ( .A(n27105), .B(n27106), .Z(n27104) );
  XOR U26965 ( .A(n27103), .B(n26806), .Z(n27106) );
  XNOR U26966 ( .A(p_input[456]), .B(n27107), .Z(n26806) );
  AND U26967 ( .A(n606), .B(n27108), .Z(n27107) );
  XOR U26968 ( .A(p_input[488]), .B(p_input[456]), .Z(n27108) );
  XNOR U26969 ( .A(n26803), .B(n27103), .Z(n27105) );
  XOR U26970 ( .A(n27109), .B(n27110), .Z(n26803) );
  AND U26971 ( .A(n604), .B(n27111), .Z(n27110) );
  XOR U26972 ( .A(p_input[424]), .B(p_input[392]), .Z(n27111) );
  XOR U26973 ( .A(n27112), .B(n27113), .Z(n27103) );
  AND U26974 ( .A(n27114), .B(n27115), .Z(n27113) );
  XOR U26975 ( .A(n27112), .B(n26818), .Z(n27115) );
  XNOR U26976 ( .A(p_input[455]), .B(n27116), .Z(n26818) );
  AND U26977 ( .A(n606), .B(n27117), .Z(n27116) );
  XOR U26978 ( .A(p_input[487]), .B(p_input[455]), .Z(n27117) );
  XNOR U26979 ( .A(n26815), .B(n27112), .Z(n27114) );
  XOR U26980 ( .A(n27118), .B(n27119), .Z(n26815) );
  AND U26981 ( .A(n604), .B(n27120), .Z(n27119) );
  XOR U26982 ( .A(p_input[423]), .B(p_input[391]), .Z(n27120) );
  XOR U26983 ( .A(n27121), .B(n27122), .Z(n27112) );
  AND U26984 ( .A(n27123), .B(n27124), .Z(n27122) );
  XOR U26985 ( .A(n27121), .B(n26830), .Z(n27124) );
  XNOR U26986 ( .A(p_input[454]), .B(n27125), .Z(n26830) );
  AND U26987 ( .A(n606), .B(n27126), .Z(n27125) );
  XOR U26988 ( .A(p_input[486]), .B(p_input[454]), .Z(n27126) );
  XNOR U26989 ( .A(n26827), .B(n27121), .Z(n27123) );
  XOR U26990 ( .A(n27127), .B(n27128), .Z(n26827) );
  AND U26991 ( .A(n604), .B(n27129), .Z(n27128) );
  XOR U26992 ( .A(p_input[422]), .B(p_input[390]), .Z(n27129) );
  XOR U26993 ( .A(n27130), .B(n27131), .Z(n27121) );
  AND U26994 ( .A(n27132), .B(n27133), .Z(n27131) );
  XOR U26995 ( .A(n27130), .B(n26842), .Z(n27133) );
  XNOR U26996 ( .A(p_input[453]), .B(n27134), .Z(n26842) );
  AND U26997 ( .A(n606), .B(n27135), .Z(n27134) );
  XOR U26998 ( .A(p_input[485]), .B(p_input[453]), .Z(n27135) );
  XNOR U26999 ( .A(n26839), .B(n27130), .Z(n27132) );
  XOR U27000 ( .A(n27136), .B(n27137), .Z(n26839) );
  AND U27001 ( .A(n604), .B(n27138), .Z(n27137) );
  XOR U27002 ( .A(p_input[421]), .B(p_input[389]), .Z(n27138) );
  XOR U27003 ( .A(n27139), .B(n27140), .Z(n27130) );
  AND U27004 ( .A(n27141), .B(n27142), .Z(n27140) );
  XOR U27005 ( .A(n27139), .B(n26854), .Z(n27142) );
  XNOR U27006 ( .A(p_input[452]), .B(n27143), .Z(n26854) );
  AND U27007 ( .A(n606), .B(n27144), .Z(n27143) );
  XOR U27008 ( .A(p_input[484]), .B(p_input[452]), .Z(n27144) );
  XNOR U27009 ( .A(n26851), .B(n27139), .Z(n27141) );
  XOR U27010 ( .A(n27145), .B(n27146), .Z(n26851) );
  AND U27011 ( .A(n604), .B(n27147), .Z(n27146) );
  XOR U27012 ( .A(p_input[420]), .B(p_input[388]), .Z(n27147) );
  XOR U27013 ( .A(n27148), .B(n27149), .Z(n27139) );
  AND U27014 ( .A(n27150), .B(n27151), .Z(n27149) );
  XOR U27015 ( .A(n27148), .B(n26866), .Z(n27151) );
  XNOR U27016 ( .A(p_input[451]), .B(n27152), .Z(n26866) );
  AND U27017 ( .A(n606), .B(n27153), .Z(n27152) );
  XOR U27018 ( .A(p_input[483]), .B(p_input[451]), .Z(n27153) );
  XNOR U27019 ( .A(n26863), .B(n27148), .Z(n27150) );
  XOR U27020 ( .A(n27154), .B(n27155), .Z(n26863) );
  AND U27021 ( .A(n604), .B(n27156), .Z(n27155) );
  XOR U27022 ( .A(p_input[419]), .B(p_input[387]), .Z(n27156) );
  XOR U27023 ( .A(n27157), .B(n27158), .Z(n27148) );
  AND U27024 ( .A(n27159), .B(n27160), .Z(n27158) );
  XOR U27025 ( .A(n26878), .B(n27157), .Z(n27160) );
  XNOR U27026 ( .A(p_input[450]), .B(n27161), .Z(n26878) );
  AND U27027 ( .A(n606), .B(n27162), .Z(n27161) );
  XOR U27028 ( .A(p_input[482]), .B(p_input[450]), .Z(n27162) );
  XNOR U27029 ( .A(n27157), .B(n26875), .Z(n27159) );
  XOR U27030 ( .A(n27163), .B(n27164), .Z(n26875) );
  AND U27031 ( .A(n604), .B(n27165), .Z(n27164) );
  XOR U27032 ( .A(p_input[418]), .B(p_input[386]), .Z(n27165) );
  XOR U27033 ( .A(n27166), .B(n27167), .Z(n27157) );
  AND U27034 ( .A(n27168), .B(n27169), .Z(n27167) );
  XNOR U27035 ( .A(n27170), .B(n26891), .Z(n27169) );
  XNOR U27036 ( .A(p_input[449]), .B(n27171), .Z(n26891) );
  AND U27037 ( .A(n606), .B(n27172), .Z(n27171) );
  XNOR U27038 ( .A(p_input[481]), .B(n27173), .Z(n27172) );
  IV U27039 ( .A(p_input[449]), .Z(n27173) );
  XNOR U27040 ( .A(n26888), .B(n27166), .Z(n27168) );
  XNOR U27041 ( .A(p_input[385]), .B(n27174), .Z(n26888) );
  AND U27042 ( .A(n604), .B(n27175), .Z(n27174) );
  XOR U27043 ( .A(p_input[417]), .B(p_input[385]), .Z(n27175) );
  IV U27044 ( .A(n27170), .Z(n27166) );
  AND U27045 ( .A(n26896), .B(n26899), .Z(n27170) );
  XOR U27046 ( .A(p_input[448]), .B(n27176), .Z(n26899) );
  AND U27047 ( .A(n606), .B(n27177), .Z(n27176) );
  XOR U27048 ( .A(p_input[480]), .B(p_input[448]), .Z(n27177) );
  XOR U27049 ( .A(n27178), .B(n27179), .Z(n606) );
  AND U27050 ( .A(n27180), .B(n27181), .Z(n27179) );
  XNOR U27051 ( .A(p_input[511]), .B(n27178), .Z(n27181) );
  XOR U27052 ( .A(n27178), .B(p_input[479]), .Z(n27180) );
  XOR U27053 ( .A(n27182), .B(n27183), .Z(n27178) );
  AND U27054 ( .A(n27184), .B(n27185), .Z(n27183) );
  XNOR U27055 ( .A(p_input[510]), .B(n27182), .Z(n27185) );
  XOR U27056 ( .A(n27182), .B(p_input[478]), .Z(n27184) );
  XOR U27057 ( .A(n27186), .B(n27187), .Z(n27182) );
  AND U27058 ( .A(n27188), .B(n27189), .Z(n27187) );
  XNOR U27059 ( .A(p_input[509]), .B(n27186), .Z(n27189) );
  XOR U27060 ( .A(n27186), .B(p_input[477]), .Z(n27188) );
  XOR U27061 ( .A(n27190), .B(n27191), .Z(n27186) );
  AND U27062 ( .A(n27192), .B(n27193), .Z(n27191) );
  XNOR U27063 ( .A(p_input[508]), .B(n27190), .Z(n27193) );
  XOR U27064 ( .A(n27190), .B(p_input[476]), .Z(n27192) );
  XOR U27065 ( .A(n27194), .B(n27195), .Z(n27190) );
  AND U27066 ( .A(n27196), .B(n27197), .Z(n27195) );
  XNOR U27067 ( .A(p_input[507]), .B(n27194), .Z(n27197) );
  XOR U27068 ( .A(n27194), .B(p_input[475]), .Z(n27196) );
  XOR U27069 ( .A(n27198), .B(n27199), .Z(n27194) );
  AND U27070 ( .A(n27200), .B(n27201), .Z(n27199) );
  XNOR U27071 ( .A(p_input[506]), .B(n27198), .Z(n27201) );
  XOR U27072 ( .A(n27198), .B(p_input[474]), .Z(n27200) );
  XOR U27073 ( .A(n27202), .B(n27203), .Z(n27198) );
  AND U27074 ( .A(n27204), .B(n27205), .Z(n27203) );
  XNOR U27075 ( .A(p_input[505]), .B(n27202), .Z(n27205) );
  XOR U27076 ( .A(n27202), .B(p_input[473]), .Z(n27204) );
  XOR U27077 ( .A(n27206), .B(n27207), .Z(n27202) );
  AND U27078 ( .A(n27208), .B(n27209), .Z(n27207) );
  XNOR U27079 ( .A(p_input[504]), .B(n27206), .Z(n27209) );
  XOR U27080 ( .A(n27206), .B(p_input[472]), .Z(n27208) );
  XOR U27081 ( .A(n27210), .B(n27211), .Z(n27206) );
  AND U27082 ( .A(n27212), .B(n27213), .Z(n27211) );
  XNOR U27083 ( .A(p_input[503]), .B(n27210), .Z(n27213) );
  XOR U27084 ( .A(n27210), .B(p_input[471]), .Z(n27212) );
  XOR U27085 ( .A(n27214), .B(n27215), .Z(n27210) );
  AND U27086 ( .A(n27216), .B(n27217), .Z(n27215) );
  XNOR U27087 ( .A(p_input[502]), .B(n27214), .Z(n27217) );
  XOR U27088 ( .A(n27214), .B(p_input[470]), .Z(n27216) );
  XOR U27089 ( .A(n27218), .B(n27219), .Z(n27214) );
  AND U27090 ( .A(n27220), .B(n27221), .Z(n27219) );
  XNOR U27091 ( .A(p_input[501]), .B(n27218), .Z(n27221) );
  XOR U27092 ( .A(n27218), .B(p_input[469]), .Z(n27220) );
  XOR U27093 ( .A(n27222), .B(n27223), .Z(n27218) );
  AND U27094 ( .A(n27224), .B(n27225), .Z(n27223) );
  XNOR U27095 ( .A(p_input[500]), .B(n27222), .Z(n27225) );
  XOR U27096 ( .A(n27222), .B(p_input[468]), .Z(n27224) );
  XOR U27097 ( .A(n27226), .B(n27227), .Z(n27222) );
  AND U27098 ( .A(n27228), .B(n27229), .Z(n27227) );
  XNOR U27099 ( .A(p_input[499]), .B(n27226), .Z(n27229) );
  XOR U27100 ( .A(n27226), .B(p_input[467]), .Z(n27228) );
  XOR U27101 ( .A(n27230), .B(n27231), .Z(n27226) );
  AND U27102 ( .A(n27232), .B(n27233), .Z(n27231) );
  XNOR U27103 ( .A(p_input[498]), .B(n27230), .Z(n27233) );
  XOR U27104 ( .A(n27230), .B(p_input[466]), .Z(n27232) );
  XOR U27105 ( .A(n27234), .B(n27235), .Z(n27230) );
  AND U27106 ( .A(n27236), .B(n27237), .Z(n27235) );
  XNOR U27107 ( .A(p_input[497]), .B(n27234), .Z(n27237) );
  XOR U27108 ( .A(n27234), .B(p_input[465]), .Z(n27236) );
  XOR U27109 ( .A(n27238), .B(n27239), .Z(n27234) );
  AND U27110 ( .A(n27240), .B(n27241), .Z(n27239) );
  XNOR U27111 ( .A(p_input[496]), .B(n27238), .Z(n27241) );
  XOR U27112 ( .A(n27238), .B(p_input[464]), .Z(n27240) );
  XOR U27113 ( .A(n27242), .B(n27243), .Z(n27238) );
  AND U27114 ( .A(n27244), .B(n27245), .Z(n27243) );
  XNOR U27115 ( .A(p_input[495]), .B(n27242), .Z(n27245) );
  XOR U27116 ( .A(n27242), .B(p_input[463]), .Z(n27244) );
  XOR U27117 ( .A(n27246), .B(n27247), .Z(n27242) );
  AND U27118 ( .A(n27248), .B(n27249), .Z(n27247) );
  XNOR U27119 ( .A(p_input[494]), .B(n27246), .Z(n27249) );
  XOR U27120 ( .A(n27246), .B(p_input[462]), .Z(n27248) );
  XOR U27121 ( .A(n27250), .B(n27251), .Z(n27246) );
  AND U27122 ( .A(n27252), .B(n27253), .Z(n27251) );
  XNOR U27123 ( .A(p_input[493]), .B(n27250), .Z(n27253) );
  XOR U27124 ( .A(n27250), .B(p_input[461]), .Z(n27252) );
  XOR U27125 ( .A(n27254), .B(n27255), .Z(n27250) );
  AND U27126 ( .A(n27256), .B(n27257), .Z(n27255) );
  XNOR U27127 ( .A(p_input[492]), .B(n27254), .Z(n27257) );
  XOR U27128 ( .A(n27254), .B(p_input[460]), .Z(n27256) );
  XOR U27129 ( .A(n27258), .B(n27259), .Z(n27254) );
  AND U27130 ( .A(n27260), .B(n27261), .Z(n27259) );
  XNOR U27131 ( .A(p_input[491]), .B(n27258), .Z(n27261) );
  XOR U27132 ( .A(n27258), .B(p_input[459]), .Z(n27260) );
  XOR U27133 ( .A(n27262), .B(n27263), .Z(n27258) );
  AND U27134 ( .A(n27264), .B(n27265), .Z(n27263) );
  XNOR U27135 ( .A(p_input[490]), .B(n27262), .Z(n27265) );
  XOR U27136 ( .A(n27262), .B(p_input[458]), .Z(n27264) );
  XOR U27137 ( .A(n27266), .B(n27267), .Z(n27262) );
  AND U27138 ( .A(n27268), .B(n27269), .Z(n27267) );
  XNOR U27139 ( .A(p_input[489]), .B(n27266), .Z(n27269) );
  XOR U27140 ( .A(n27266), .B(p_input[457]), .Z(n27268) );
  XOR U27141 ( .A(n27270), .B(n27271), .Z(n27266) );
  AND U27142 ( .A(n27272), .B(n27273), .Z(n27271) );
  XNOR U27143 ( .A(p_input[488]), .B(n27270), .Z(n27273) );
  XOR U27144 ( .A(n27270), .B(p_input[456]), .Z(n27272) );
  XOR U27145 ( .A(n27274), .B(n27275), .Z(n27270) );
  AND U27146 ( .A(n27276), .B(n27277), .Z(n27275) );
  XNOR U27147 ( .A(p_input[487]), .B(n27274), .Z(n27277) );
  XOR U27148 ( .A(n27274), .B(p_input[455]), .Z(n27276) );
  XOR U27149 ( .A(n27278), .B(n27279), .Z(n27274) );
  AND U27150 ( .A(n27280), .B(n27281), .Z(n27279) );
  XNOR U27151 ( .A(p_input[486]), .B(n27278), .Z(n27281) );
  XOR U27152 ( .A(n27278), .B(p_input[454]), .Z(n27280) );
  XOR U27153 ( .A(n27282), .B(n27283), .Z(n27278) );
  AND U27154 ( .A(n27284), .B(n27285), .Z(n27283) );
  XNOR U27155 ( .A(p_input[485]), .B(n27282), .Z(n27285) );
  XOR U27156 ( .A(n27282), .B(p_input[453]), .Z(n27284) );
  XOR U27157 ( .A(n27286), .B(n27287), .Z(n27282) );
  AND U27158 ( .A(n27288), .B(n27289), .Z(n27287) );
  XNOR U27159 ( .A(p_input[484]), .B(n27286), .Z(n27289) );
  XOR U27160 ( .A(n27286), .B(p_input[452]), .Z(n27288) );
  XOR U27161 ( .A(n27290), .B(n27291), .Z(n27286) );
  AND U27162 ( .A(n27292), .B(n27293), .Z(n27291) );
  XNOR U27163 ( .A(p_input[483]), .B(n27290), .Z(n27293) );
  XOR U27164 ( .A(n27290), .B(p_input[451]), .Z(n27292) );
  XOR U27165 ( .A(n27294), .B(n27295), .Z(n27290) );
  AND U27166 ( .A(n27296), .B(n27297), .Z(n27295) );
  XNOR U27167 ( .A(p_input[482]), .B(n27294), .Z(n27297) );
  XOR U27168 ( .A(n27294), .B(p_input[450]), .Z(n27296) );
  XNOR U27169 ( .A(n27298), .B(n27299), .Z(n27294) );
  AND U27170 ( .A(n27300), .B(n27301), .Z(n27299) );
  XOR U27171 ( .A(p_input[481]), .B(n27298), .Z(n27301) );
  XNOR U27172 ( .A(p_input[449]), .B(n27298), .Z(n27300) );
  AND U27173 ( .A(p_input[480]), .B(n27302), .Z(n27298) );
  IV U27174 ( .A(p_input[448]), .Z(n27302) );
  XNOR U27175 ( .A(p_input[384]), .B(n27303), .Z(n26896) );
  AND U27176 ( .A(n604), .B(n27304), .Z(n27303) );
  XOR U27177 ( .A(p_input[416]), .B(p_input[384]), .Z(n27304) );
  XOR U27178 ( .A(n27305), .B(n27306), .Z(n604) );
  AND U27179 ( .A(n27307), .B(n27308), .Z(n27306) );
  XNOR U27180 ( .A(p_input[447]), .B(n27305), .Z(n27308) );
  XOR U27181 ( .A(n27305), .B(p_input[415]), .Z(n27307) );
  XOR U27182 ( .A(n27309), .B(n27310), .Z(n27305) );
  AND U27183 ( .A(n27311), .B(n27312), .Z(n27310) );
  XNOR U27184 ( .A(p_input[446]), .B(n27309), .Z(n27312) );
  XNOR U27185 ( .A(n27309), .B(n26911), .Z(n27311) );
  IV U27186 ( .A(p_input[414]), .Z(n26911) );
  XOR U27187 ( .A(n27313), .B(n27314), .Z(n27309) );
  AND U27188 ( .A(n27315), .B(n27316), .Z(n27314) );
  XNOR U27189 ( .A(p_input[445]), .B(n27313), .Z(n27316) );
  XNOR U27190 ( .A(n27313), .B(n26920), .Z(n27315) );
  IV U27191 ( .A(p_input[413]), .Z(n26920) );
  XOR U27192 ( .A(n27317), .B(n27318), .Z(n27313) );
  AND U27193 ( .A(n27319), .B(n27320), .Z(n27318) );
  XNOR U27194 ( .A(p_input[444]), .B(n27317), .Z(n27320) );
  XNOR U27195 ( .A(n27317), .B(n26929), .Z(n27319) );
  IV U27196 ( .A(p_input[412]), .Z(n26929) );
  XOR U27197 ( .A(n27321), .B(n27322), .Z(n27317) );
  AND U27198 ( .A(n27323), .B(n27324), .Z(n27322) );
  XNOR U27199 ( .A(p_input[443]), .B(n27321), .Z(n27324) );
  XNOR U27200 ( .A(n27321), .B(n26938), .Z(n27323) );
  IV U27201 ( .A(p_input[411]), .Z(n26938) );
  XOR U27202 ( .A(n27325), .B(n27326), .Z(n27321) );
  AND U27203 ( .A(n27327), .B(n27328), .Z(n27326) );
  XNOR U27204 ( .A(p_input[442]), .B(n27325), .Z(n27328) );
  XNOR U27205 ( .A(n27325), .B(n26947), .Z(n27327) );
  IV U27206 ( .A(p_input[410]), .Z(n26947) );
  XOR U27207 ( .A(n27329), .B(n27330), .Z(n27325) );
  AND U27208 ( .A(n27331), .B(n27332), .Z(n27330) );
  XNOR U27209 ( .A(p_input[441]), .B(n27329), .Z(n27332) );
  XNOR U27210 ( .A(n27329), .B(n26956), .Z(n27331) );
  IV U27211 ( .A(p_input[409]), .Z(n26956) );
  XOR U27212 ( .A(n27333), .B(n27334), .Z(n27329) );
  AND U27213 ( .A(n27335), .B(n27336), .Z(n27334) );
  XNOR U27214 ( .A(p_input[440]), .B(n27333), .Z(n27336) );
  XNOR U27215 ( .A(n27333), .B(n26965), .Z(n27335) );
  IV U27216 ( .A(p_input[408]), .Z(n26965) );
  XOR U27217 ( .A(n27337), .B(n27338), .Z(n27333) );
  AND U27218 ( .A(n27339), .B(n27340), .Z(n27338) );
  XNOR U27219 ( .A(p_input[439]), .B(n27337), .Z(n27340) );
  XNOR U27220 ( .A(n27337), .B(n26974), .Z(n27339) );
  IV U27221 ( .A(p_input[407]), .Z(n26974) );
  XOR U27222 ( .A(n27341), .B(n27342), .Z(n27337) );
  AND U27223 ( .A(n27343), .B(n27344), .Z(n27342) );
  XNOR U27224 ( .A(p_input[438]), .B(n27341), .Z(n27344) );
  XNOR U27225 ( .A(n27341), .B(n26983), .Z(n27343) );
  IV U27226 ( .A(p_input[406]), .Z(n26983) );
  XOR U27227 ( .A(n27345), .B(n27346), .Z(n27341) );
  AND U27228 ( .A(n27347), .B(n27348), .Z(n27346) );
  XNOR U27229 ( .A(p_input[437]), .B(n27345), .Z(n27348) );
  XNOR U27230 ( .A(n27345), .B(n26992), .Z(n27347) );
  IV U27231 ( .A(p_input[405]), .Z(n26992) );
  XOR U27232 ( .A(n27349), .B(n27350), .Z(n27345) );
  AND U27233 ( .A(n27351), .B(n27352), .Z(n27350) );
  XNOR U27234 ( .A(p_input[436]), .B(n27349), .Z(n27352) );
  XNOR U27235 ( .A(n27349), .B(n27001), .Z(n27351) );
  IV U27236 ( .A(p_input[404]), .Z(n27001) );
  XOR U27237 ( .A(n27353), .B(n27354), .Z(n27349) );
  AND U27238 ( .A(n27355), .B(n27356), .Z(n27354) );
  XNOR U27239 ( .A(p_input[435]), .B(n27353), .Z(n27356) );
  XNOR U27240 ( .A(n27353), .B(n27010), .Z(n27355) );
  IV U27241 ( .A(p_input[403]), .Z(n27010) );
  XOR U27242 ( .A(n27357), .B(n27358), .Z(n27353) );
  AND U27243 ( .A(n27359), .B(n27360), .Z(n27358) );
  XNOR U27244 ( .A(p_input[434]), .B(n27357), .Z(n27360) );
  XNOR U27245 ( .A(n27357), .B(n27019), .Z(n27359) );
  IV U27246 ( .A(p_input[402]), .Z(n27019) );
  XOR U27247 ( .A(n27361), .B(n27362), .Z(n27357) );
  AND U27248 ( .A(n27363), .B(n27364), .Z(n27362) );
  XNOR U27249 ( .A(p_input[433]), .B(n27361), .Z(n27364) );
  XNOR U27250 ( .A(n27361), .B(n27028), .Z(n27363) );
  IV U27251 ( .A(p_input[401]), .Z(n27028) );
  XOR U27252 ( .A(n27365), .B(n27366), .Z(n27361) );
  AND U27253 ( .A(n27367), .B(n27368), .Z(n27366) );
  XNOR U27254 ( .A(p_input[432]), .B(n27365), .Z(n27368) );
  XNOR U27255 ( .A(n27365), .B(n27037), .Z(n27367) );
  IV U27256 ( .A(p_input[400]), .Z(n27037) );
  XOR U27257 ( .A(n27369), .B(n27370), .Z(n27365) );
  AND U27258 ( .A(n27371), .B(n27372), .Z(n27370) );
  XNOR U27259 ( .A(p_input[431]), .B(n27369), .Z(n27372) );
  XNOR U27260 ( .A(n27369), .B(n27046), .Z(n27371) );
  IV U27261 ( .A(p_input[399]), .Z(n27046) );
  XOR U27262 ( .A(n27373), .B(n27374), .Z(n27369) );
  AND U27263 ( .A(n27375), .B(n27376), .Z(n27374) );
  XNOR U27264 ( .A(p_input[430]), .B(n27373), .Z(n27376) );
  XNOR U27265 ( .A(n27373), .B(n27055), .Z(n27375) );
  IV U27266 ( .A(p_input[398]), .Z(n27055) );
  XOR U27267 ( .A(n27377), .B(n27378), .Z(n27373) );
  AND U27268 ( .A(n27379), .B(n27380), .Z(n27378) );
  XNOR U27269 ( .A(p_input[429]), .B(n27377), .Z(n27380) );
  XNOR U27270 ( .A(n27377), .B(n27064), .Z(n27379) );
  IV U27271 ( .A(p_input[397]), .Z(n27064) );
  XOR U27272 ( .A(n27381), .B(n27382), .Z(n27377) );
  AND U27273 ( .A(n27383), .B(n27384), .Z(n27382) );
  XNOR U27274 ( .A(p_input[428]), .B(n27381), .Z(n27384) );
  XNOR U27275 ( .A(n27381), .B(n27073), .Z(n27383) );
  IV U27276 ( .A(p_input[396]), .Z(n27073) );
  XOR U27277 ( .A(n27385), .B(n27386), .Z(n27381) );
  AND U27278 ( .A(n27387), .B(n27388), .Z(n27386) );
  XNOR U27279 ( .A(p_input[427]), .B(n27385), .Z(n27388) );
  XNOR U27280 ( .A(n27385), .B(n27082), .Z(n27387) );
  IV U27281 ( .A(p_input[395]), .Z(n27082) );
  XOR U27282 ( .A(n27389), .B(n27390), .Z(n27385) );
  AND U27283 ( .A(n27391), .B(n27392), .Z(n27390) );
  XNOR U27284 ( .A(p_input[426]), .B(n27389), .Z(n27392) );
  XNOR U27285 ( .A(n27389), .B(n27091), .Z(n27391) );
  IV U27286 ( .A(p_input[394]), .Z(n27091) );
  XOR U27287 ( .A(n27393), .B(n27394), .Z(n27389) );
  AND U27288 ( .A(n27395), .B(n27396), .Z(n27394) );
  XNOR U27289 ( .A(p_input[425]), .B(n27393), .Z(n27396) );
  XNOR U27290 ( .A(n27393), .B(n27100), .Z(n27395) );
  IV U27291 ( .A(p_input[393]), .Z(n27100) );
  XOR U27292 ( .A(n27397), .B(n27398), .Z(n27393) );
  AND U27293 ( .A(n27399), .B(n27400), .Z(n27398) );
  XNOR U27294 ( .A(p_input[424]), .B(n27397), .Z(n27400) );
  XNOR U27295 ( .A(n27397), .B(n27109), .Z(n27399) );
  IV U27296 ( .A(p_input[392]), .Z(n27109) );
  XOR U27297 ( .A(n27401), .B(n27402), .Z(n27397) );
  AND U27298 ( .A(n27403), .B(n27404), .Z(n27402) );
  XNOR U27299 ( .A(p_input[423]), .B(n27401), .Z(n27404) );
  XNOR U27300 ( .A(n27401), .B(n27118), .Z(n27403) );
  IV U27301 ( .A(p_input[391]), .Z(n27118) );
  XOR U27302 ( .A(n27405), .B(n27406), .Z(n27401) );
  AND U27303 ( .A(n27407), .B(n27408), .Z(n27406) );
  XNOR U27304 ( .A(p_input[422]), .B(n27405), .Z(n27408) );
  XNOR U27305 ( .A(n27405), .B(n27127), .Z(n27407) );
  IV U27306 ( .A(p_input[390]), .Z(n27127) );
  XOR U27307 ( .A(n27409), .B(n27410), .Z(n27405) );
  AND U27308 ( .A(n27411), .B(n27412), .Z(n27410) );
  XNOR U27309 ( .A(p_input[421]), .B(n27409), .Z(n27412) );
  XNOR U27310 ( .A(n27409), .B(n27136), .Z(n27411) );
  IV U27311 ( .A(p_input[389]), .Z(n27136) );
  XOR U27312 ( .A(n27413), .B(n27414), .Z(n27409) );
  AND U27313 ( .A(n27415), .B(n27416), .Z(n27414) );
  XNOR U27314 ( .A(p_input[420]), .B(n27413), .Z(n27416) );
  XNOR U27315 ( .A(n27413), .B(n27145), .Z(n27415) );
  IV U27316 ( .A(p_input[388]), .Z(n27145) );
  XOR U27317 ( .A(n27417), .B(n27418), .Z(n27413) );
  AND U27318 ( .A(n27419), .B(n27420), .Z(n27418) );
  XNOR U27319 ( .A(p_input[419]), .B(n27417), .Z(n27420) );
  XNOR U27320 ( .A(n27417), .B(n27154), .Z(n27419) );
  IV U27321 ( .A(p_input[387]), .Z(n27154) );
  XOR U27322 ( .A(n27421), .B(n27422), .Z(n27417) );
  AND U27323 ( .A(n27423), .B(n27424), .Z(n27422) );
  XNOR U27324 ( .A(p_input[418]), .B(n27421), .Z(n27424) );
  XNOR U27325 ( .A(n27421), .B(n27163), .Z(n27423) );
  IV U27326 ( .A(p_input[386]), .Z(n27163) );
  XNOR U27327 ( .A(n27425), .B(n27426), .Z(n27421) );
  AND U27328 ( .A(n27427), .B(n27428), .Z(n27426) );
  XOR U27329 ( .A(p_input[417]), .B(n27425), .Z(n27428) );
  XNOR U27330 ( .A(p_input[385]), .B(n27425), .Z(n27427) );
  AND U27331 ( .A(p_input[416]), .B(n27429), .Z(n27425) );
  IV U27332 ( .A(p_input[384]), .Z(n27429) );
  XOR U27333 ( .A(n27430), .B(n27431), .Z(n26519) );
  AND U27334 ( .A(n404), .B(n27432), .Z(n27431) );
  XNOR U27335 ( .A(n27433), .B(n27430), .Z(n27432) );
  XOR U27336 ( .A(n27434), .B(n27435), .Z(n404) );
  AND U27337 ( .A(n27436), .B(n27437), .Z(n27435) );
  XNOR U27338 ( .A(n26534), .B(n27434), .Z(n27437) );
  AND U27339 ( .A(p_input[383]), .B(p_input[351]), .Z(n26534) );
  XNOR U27340 ( .A(n27434), .B(n26531), .Z(n27436) );
  IV U27341 ( .A(n27438), .Z(n26531) );
  AND U27342 ( .A(p_input[287]), .B(p_input[319]), .Z(n27438) );
  XOR U27343 ( .A(n27439), .B(n27440), .Z(n27434) );
  AND U27344 ( .A(n27441), .B(n27442), .Z(n27440) );
  XOR U27345 ( .A(n27439), .B(n26546), .Z(n27442) );
  XNOR U27346 ( .A(p_input[350]), .B(n27443), .Z(n26546) );
  AND U27347 ( .A(n610), .B(n27444), .Z(n27443) );
  XOR U27348 ( .A(p_input[382]), .B(p_input[350]), .Z(n27444) );
  XNOR U27349 ( .A(n26543), .B(n27439), .Z(n27441) );
  XOR U27350 ( .A(n27445), .B(n27446), .Z(n26543) );
  AND U27351 ( .A(n607), .B(n27447), .Z(n27446) );
  XOR U27352 ( .A(p_input[318]), .B(p_input[286]), .Z(n27447) );
  XOR U27353 ( .A(n27448), .B(n27449), .Z(n27439) );
  AND U27354 ( .A(n27450), .B(n27451), .Z(n27449) );
  XOR U27355 ( .A(n27448), .B(n26558), .Z(n27451) );
  XNOR U27356 ( .A(p_input[349]), .B(n27452), .Z(n26558) );
  AND U27357 ( .A(n610), .B(n27453), .Z(n27452) );
  XOR U27358 ( .A(p_input[381]), .B(p_input[349]), .Z(n27453) );
  XNOR U27359 ( .A(n26555), .B(n27448), .Z(n27450) );
  XOR U27360 ( .A(n27454), .B(n27455), .Z(n26555) );
  AND U27361 ( .A(n607), .B(n27456), .Z(n27455) );
  XOR U27362 ( .A(p_input[317]), .B(p_input[285]), .Z(n27456) );
  XOR U27363 ( .A(n27457), .B(n27458), .Z(n27448) );
  AND U27364 ( .A(n27459), .B(n27460), .Z(n27458) );
  XOR U27365 ( .A(n27457), .B(n26570), .Z(n27460) );
  XNOR U27366 ( .A(p_input[348]), .B(n27461), .Z(n26570) );
  AND U27367 ( .A(n610), .B(n27462), .Z(n27461) );
  XOR U27368 ( .A(p_input[380]), .B(p_input[348]), .Z(n27462) );
  XNOR U27369 ( .A(n26567), .B(n27457), .Z(n27459) );
  XOR U27370 ( .A(n27463), .B(n27464), .Z(n26567) );
  AND U27371 ( .A(n607), .B(n27465), .Z(n27464) );
  XOR U27372 ( .A(p_input[316]), .B(p_input[284]), .Z(n27465) );
  XOR U27373 ( .A(n27466), .B(n27467), .Z(n27457) );
  AND U27374 ( .A(n27468), .B(n27469), .Z(n27467) );
  XOR U27375 ( .A(n27466), .B(n26582), .Z(n27469) );
  XNOR U27376 ( .A(p_input[347]), .B(n27470), .Z(n26582) );
  AND U27377 ( .A(n610), .B(n27471), .Z(n27470) );
  XOR U27378 ( .A(p_input[379]), .B(p_input[347]), .Z(n27471) );
  XNOR U27379 ( .A(n26579), .B(n27466), .Z(n27468) );
  XOR U27380 ( .A(n27472), .B(n27473), .Z(n26579) );
  AND U27381 ( .A(n607), .B(n27474), .Z(n27473) );
  XOR U27382 ( .A(p_input[315]), .B(p_input[283]), .Z(n27474) );
  XOR U27383 ( .A(n27475), .B(n27476), .Z(n27466) );
  AND U27384 ( .A(n27477), .B(n27478), .Z(n27476) );
  XOR U27385 ( .A(n27475), .B(n26594), .Z(n27478) );
  XNOR U27386 ( .A(p_input[346]), .B(n27479), .Z(n26594) );
  AND U27387 ( .A(n610), .B(n27480), .Z(n27479) );
  XOR U27388 ( .A(p_input[378]), .B(p_input[346]), .Z(n27480) );
  XNOR U27389 ( .A(n26591), .B(n27475), .Z(n27477) );
  XOR U27390 ( .A(n27481), .B(n27482), .Z(n26591) );
  AND U27391 ( .A(n607), .B(n27483), .Z(n27482) );
  XOR U27392 ( .A(p_input[314]), .B(p_input[282]), .Z(n27483) );
  XOR U27393 ( .A(n27484), .B(n27485), .Z(n27475) );
  AND U27394 ( .A(n27486), .B(n27487), .Z(n27485) );
  XOR U27395 ( .A(n27484), .B(n26606), .Z(n27487) );
  XNOR U27396 ( .A(p_input[345]), .B(n27488), .Z(n26606) );
  AND U27397 ( .A(n610), .B(n27489), .Z(n27488) );
  XOR U27398 ( .A(p_input[377]), .B(p_input[345]), .Z(n27489) );
  XNOR U27399 ( .A(n26603), .B(n27484), .Z(n27486) );
  XOR U27400 ( .A(n27490), .B(n27491), .Z(n26603) );
  AND U27401 ( .A(n607), .B(n27492), .Z(n27491) );
  XOR U27402 ( .A(p_input[313]), .B(p_input[281]), .Z(n27492) );
  XOR U27403 ( .A(n27493), .B(n27494), .Z(n27484) );
  AND U27404 ( .A(n27495), .B(n27496), .Z(n27494) );
  XOR U27405 ( .A(n27493), .B(n26618), .Z(n27496) );
  XNOR U27406 ( .A(p_input[344]), .B(n27497), .Z(n26618) );
  AND U27407 ( .A(n610), .B(n27498), .Z(n27497) );
  XOR U27408 ( .A(p_input[376]), .B(p_input[344]), .Z(n27498) );
  XNOR U27409 ( .A(n26615), .B(n27493), .Z(n27495) );
  XOR U27410 ( .A(n27499), .B(n27500), .Z(n26615) );
  AND U27411 ( .A(n607), .B(n27501), .Z(n27500) );
  XOR U27412 ( .A(p_input[312]), .B(p_input[280]), .Z(n27501) );
  XOR U27413 ( .A(n27502), .B(n27503), .Z(n27493) );
  AND U27414 ( .A(n27504), .B(n27505), .Z(n27503) );
  XOR U27415 ( .A(n27502), .B(n26630), .Z(n27505) );
  XNOR U27416 ( .A(p_input[343]), .B(n27506), .Z(n26630) );
  AND U27417 ( .A(n610), .B(n27507), .Z(n27506) );
  XOR U27418 ( .A(p_input[375]), .B(p_input[343]), .Z(n27507) );
  XNOR U27419 ( .A(n26627), .B(n27502), .Z(n27504) );
  XOR U27420 ( .A(n27508), .B(n27509), .Z(n26627) );
  AND U27421 ( .A(n607), .B(n27510), .Z(n27509) );
  XOR U27422 ( .A(p_input[311]), .B(p_input[279]), .Z(n27510) );
  XOR U27423 ( .A(n27511), .B(n27512), .Z(n27502) );
  AND U27424 ( .A(n27513), .B(n27514), .Z(n27512) );
  XOR U27425 ( .A(n27511), .B(n26642), .Z(n27514) );
  XNOR U27426 ( .A(p_input[342]), .B(n27515), .Z(n26642) );
  AND U27427 ( .A(n610), .B(n27516), .Z(n27515) );
  XOR U27428 ( .A(p_input[374]), .B(p_input[342]), .Z(n27516) );
  XNOR U27429 ( .A(n26639), .B(n27511), .Z(n27513) );
  XOR U27430 ( .A(n27517), .B(n27518), .Z(n26639) );
  AND U27431 ( .A(n607), .B(n27519), .Z(n27518) );
  XOR U27432 ( .A(p_input[310]), .B(p_input[278]), .Z(n27519) );
  XOR U27433 ( .A(n27520), .B(n27521), .Z(n27511) );
  AND U27434 ( .A(n27522), .B(n27523), .Z(n27521) );
  XOR U27435 ( .A(n27520), .B(n26654), .Z(n27523) );
  XNOR U27436 ( .A(p_input[341]), .B(n27524), .Z(n26654) );
  AND U27437 ( .A(n610), .B(n27525), .Z(n27524) );
  XOR U27438 ( .A(p_input[373]), .B(p_input[341]), .Z(n27525) );
  XNOR U27439 ( .A(n26651), .B(n27520), .Z(n27522) );
  XOR U27440 ( .A(n27526), .B(n27527), .Z(n26651) );
  AND U27441 ( .A(n607), .B(n27528), .Z(n27527) );
  XOR U27442 ( .A(p_input[309]), .B(p_input[277]), .Z(n27528) );
  XOR U27443 ( .A(n27529), .B(n27530), .Z(n27520) );
  AND U27444 ( .A(n27531), .B(n27532), .Z(n27530) );
  XOR U27445 ( .A(n27529), .B(n26666), .Z(n27532) );
  XNOR U27446 ( .A(p_input[340]), .B(n27533), .Z(n26666) );
  AND U27447 ( .A(n610), .B(n27534), .Z(n27533) );
  XOR U27448 ( .A(p_input[372]), .B(p_input[340]), .Z(n27534) );
  XNOR U27449 ( .A(n26663), .B(n27529), .Z(n27531) );
  XOR U27450 ( .A(n27535), .B(n27536), .Z(n26663) );
  AND U27451 ( .A(n607), .B(n27537), .Z(n27536) );
  XOR U27452 ( .A(p_input[308]), .B(p_input[276]), .Z(n27537) );
  XOR U27453 ( .A(n27538), .B(n27539), .Z(n27529) );
  AND U27454 ( .A(n27540), .B(n27541), .Z(n27539) );
  XOR U27455 ( .A(n27538), .B(n26678), .Z(n27541) );
  XNOR U27456 ( .A(p_input[339]), .B(n27542), .Z(n26678) );
  AND U27457 ( .A(n610), .B(n27543), .Z(n27542) );
  XOR U27458 ( .A(p_input[371]), .B(p_input[339]), .Z(n27543) );
  XNOR U27459 ( .A(n26675), .B(n27538), .Z(n27540) );
  XOR U27460 ( .A(n27544), .B(n27545), .Z(n26675) );
  AND U27461 ( .A(n607), .B(n27546), .Z(n27545) );
  XOR U27462 ( .A(p_input[307]), .B(p_input[275]), .Z(n27546) );
  XOR U27463 ( .A(n27547), .B(n27548), .Z(n27538) );
  AND U27464 ( .A(n27549), .B(n27550), .Z(n27548) );
  XOR U27465 ( .A(n27547), .B(n26690), .Z(n27550) );
  XNOR U27466 ( .A(p_input[338]), .B(n27551), .Z(n26690) );
  AND U27467 ( .A(n610), .B(n27552), .Z(n27551) );
  XOR U27468 ( .A(p_input[370]), .B(p_input[338]), .Z(n27552) );
  XNOR U27469 ( .A(n26687), .B(n27547), .Z(n27549) );
  XOR U27470 ( .A(n27553), .B(n27554), .Z(n26687) );
  AND U27471 ( .A(n607), .B(n27555), .Z(n27554) );
  XOR U27472 ( .A(p_input[306]), .B(p_input[274]), .Z(n27555) );
  XOR U27473 ( .A(n27556), .B(n27557), .Z(n27547) );
  AND U27474 ( .A(n27558), .B(n27559), .Z(n27557) );
  XOR U27475 ( .A(n27556), .B(n26702), .Z(n27559) );
  XNOR U27476 ( .A(p_input[337]), .B(n27560), .Z(n26702) );
  AND U27477 ( .A(n610), .B(n27561), .Z(n27560) );
  XOR U27478 ( .A(p_input[369]), .B(p_input[337]), .Z(n27561) );
  XNOR U27479 ( .A(n26699), .B(n27556), .Z(n27558) );
  XOR U27480 ( .A(n27562), .B(n27563), .Z(n26699) );
  AND U27481 ( .A(n607), .B(n27564), .Z(n27563) );
  XOR U27482 ( .A(p_input[305]), .B(p_input[273]), .Z(n27564) );
  XOR U27483 ( .A(n27565), .B(n27566), .Z(n27556) );
  AND U27484 ( .A(n27567), .B(n27568), .Z(n27566) );
  XOR U27485 ( .A(n27565), .B(n26714), .Z(n27568) );
  XNOR U27486 ( .A(p_input[336]), .B(n27569), .Z(n26714) );
  AND U27487 ( .A(n610), .B(n27570), .Z(n27569) );
  XOR U27488 ( .A(p_input[368]), .B(p_input[336]), .Z(n27570) );
  XNOR U27489 ( .A(n26711), .B(n27565), .Z(n27567) );
  XOR U27490 ( .A(n27571), .B(n27572), .Z(n26711) );
  AND U27491 ( .A(n607), .B(n27573), .Z(n27572) );
  XOR U27492 ( .A(p_input[304]), .B(p_input[272]), .Z(n27573) );
  XOR U27493 ( .A(n27574), .B(n27575), .Z(n27565) );
  AND U27494 ( .A(n27576), .B(n27577), .Z(n27575) );
  XOR U27495 ( .A(n27574), .B(n26726), .Z(n27577) );
  XNOR U27496 ( .A(p_input[335]), .B(n27578), .Z(n26726) );
  AND U27497 ( .A(n610), .B(n27579), .Z(n27578) );
  XOR U27498 ( .A(p_input[367]), .B(p_input[335]), .Z(n27579) );
  XNOR U27499 ( .A(n26723), .B(n27574), .Z(n27576) );
  XOR U27500 ( .A(n27580), .B(n27581), .Z(n26723) );
  AND U27501 ( .A(n607), .B(n27582), .Z(n27581) );
  XOR U27502 ( .A(p_input[303]), .B(p_input[271]), .Z(n27582) );
  XOR U27503 ( .A(n27583), .B(n27584), .Z(n27574) );
  AND U27504 ( .A(n27585), .B(n27586), .Z(n27584) );
  XOR U27505 ( .A(n27583), .B(n26738), .Z(n27586) );
  XNOR U27506 ( .A(p_input[334]), .B(n27587), .Z(n26738) );
  AND U27507 ( .A(n610), .B(n27588), .Z(n27587) );
  XOR U27508 ( .A(p_input[366]), .B(p_input[334]), .Z(n27588) );
  XNOR U27509 ( .A(n26735), .B(n27583), .Z(n27585) );
  XOR U27510 ( .A(n27589), .B(n27590), .Z(n26735) );
  AND U27511 ( .A(n607), .B(n27591), .Z(n27590) );
  XOR U27512 ( .A(p_input[302]), .B(p_input[270]), .Z(n27591) );
  XOR U27513 ( .A(n27592), .B(n27593), .Z(n27583) );
  AND U27514 ( .A(n27594), .B(n27595), .Z(n27593) );
  XOR U27515 ( .A(n27592), .B(n26750), .Z(n27595) );
  XNOR U27516 ( .A(p_input[333]), .B(n27596), .Z(n26750) );
  AND U27517 ( .A(n610), .B(n27597), .Z(n27596) );
  XOR U27518 ( .A(p_input[365]), .B(p_input[333]), .Z(n27597) );
  XNOR U27519 ( .A(n26747), .B(n27592), .Z(n27594) );
  XOR U27520 ( .A(n27598), .B(n27599), .Z(n26747) );
  AND U27521 ( .A(n607), .B(n27600), .Z(n27599) );
  XOR U27522 ( .A(p_input[301]), .B(p_input[269]), .Z(n27600) );
  XOR U27523 ( .A(n27601), .B(n27602), .Z(n27592) );
  AND U27524 ( .A(n27603), .B(n27604), .Z(n27602) );
  XOR U27525 ( .A(n27601), .B(n26762), .Z(n27604) );
  XNOR U27526 ( .A(p_input[332]), .B(n27605), .Z(n26762) );
  AND U27527 ( .A(n610), .B(n27606), .Z(n27605) );
  XOR U27528 ( .A(p_input[364]), .B(p_input[332]), .Z(n27606) );
  XNOR U27529 ( .A(n26759), .B(n27601), .Z(n27603) );
  XOR U27530 ( .A(n27607), .B(n27608), .Z(n26759) );
  AND U27531 ( .A(n607), .B(n27609), .Z(n27608) );
  XOR U27532 ( .A(p_input[300]), .B(p_input[268]), .Z(n27609) );
  XOR U27533 ( .A(n27610), .B(n27611), .Z(n27601) );
  AND U27534 ( .A(n27612), .B(n27613), .Z(n27611) );
  XOR U27535 ( .A(n27610), .B(n26774), .Z(n27613) );
  XNOR U27536 ( .A(p_input[331]), .B(n27614), .Z(n26774) );
  AND U27537 ( .A(n610), .B(n27615), .Z(n27614) );
  XOR U27538 ( .A(p_input[363]), .B(p_input[331]), .Z(n27615) );
  XNOR U27539 ( .A(n26771), .B(n27610), .Z(n27612) );
  XOR U27540 ( .A(n27616), .B(n27617), .Z(n26771) );
  AND U27541 ( .A(n607), .B(n27618), .Z(n27617) );
  XOR U27542 ( .A(p_input[299]), .B(p_input[267]), .Z(n27618) );
  XOR U27543 ( .A(n27619), .B(n27620), .Z(n27610) );
  AND U27544 ( .A(n27621), .B(n27622), .Z(n27620) );
  XOR U27545 ( .A(n27619), .B(n26786), .Z(n27622) );
  XNOR U27546 ( .A(p_input[330]), .B(n27623), .Z(n26786) );
  AND U27547 ( .A(n610), .B(n27624), .Z(n27623) );
  XOR U27548 ( .A(p_input[362]), .B(p_input[330]), .Z(n27624) );
  XNOR U27549 ( .A(n26783), .B(n27619), .Z(n27621) );
  XOR U27550 ( .A(n27625), .B(n27626), .Z(n26783) );
  AND U27551 ( .A(n607), .B(n27627), .Z(n27626) );
  XOR U27552 ( .A(p_input[298]), .B(p_input[266]), .Z(n27627) );
  XOR U27553 ( .A(n27628), .B(n27629), .Z(n27619) );
  AND U27554 ( .A(n27630), .B(n27631), .Z(n27629) );
  XOR U27555 ( .A(n27628), .B(n26798), .Z(n27631) );
  XNOR U27556 ( .A(p_input[329]), .B(n27632), .Z(n26798) );
  AND U27557 ( .A(n610), .B(n27633), .Z(n27632) );
  XOR U27558 ( .A(p_input[361]), .B(p_input[329]), .Z(n27633) );
  XNOR U27559 ( .A(n26795), .B(n27628), .Z(n27630) );
  XOR U27560 ( .A(n27634), .B(n27635), .Z(n26795) );
  AND U27561 ( .A(n607), .B(n27636), .Z(n27635) );
  XOR U27562 ( .A(p_input[297]), .B(p_input[265]), .Z(n27636) );
  XOR U27563 ( .A(n27637), .B(n27638), .Z(n27628) );
  AND U27564 ( .A(n27639), .B(n27640), .Z(n27638) );
  XOR U27565 ( .A(n27637), .B(n26810), .Z(n27640) );
  XNOR U27566 ( .A(p_input[328]), .B(n27641), .Z(n26810) );
  AND U27567 ( .A(n610), .B(n27642), .Z(n27641) );
  XOR U27568 ( .A(p_input[360]), .B(p_input[328]), .Z(n27642) );
  XNOR U27569 ( .A(n26807), .B(n27637), .Z(n27639) );
  XOR U27570 ( .A(n27643), .B(n27644), .Z(n26807) );
  AND U27571 ( .A(n607), .B(n27645), .Z(n27644) );
  XOR U27572 ( .A(p_input[296]), .B(p_input[264]), .Z(n27645) );
  XOR U27573 ( .A(n27646), .B(n27647), .Z(n27637) );
  AND U27574 ( .A(n27648), .B(n27649), .Z(n27647) );
  XOR U27575 ( .A(n27646), .B(n26822), .Z(n27649) );
  XNOR U27576 ( .A(p_input[327]), .B(n27650), .Z(n26822) );
  AND U27577 ( .A(n610), .B(n27651), .Z(n27650) );
  XOR U27578 ( .A(p_input[359]), .B(p_input[327]), .Z(n27651) );
  XNOR U27579 ( .A(n26819), .B(n27646), .Z(n27648) );
  XOR U27580 ( .A(n27652), .B(n27653), .Z(n26819) );
  AND U27581 ( .A(n607), .B(n27654), .Z(n27653) );
  XOR U27582 ( .A(p_input[295]), .B(p_input[263]), .Z(n27654) );
  XOR U27583 ( .A(n27655), .B(n27656), .Z(n27646) );
  AND U27584 ( .A(n27657), .B(n27658), .Z(n27656) );
  XOR U27585 ( .A(n27655), .B(n26834), .Z(n27658) );
  XNOR U27586 ( .A(p_input[326]), .B(n27659), .Z(n26834) );
  AND U27587 ( .A(n610), .B(n27660), .Z(n27659) );
  XOR U27588 ( .A(p_input[358]), .B(p_input[326]), .Z(n27660) );
  XNOR U27589 ( .A(n26831), .B(n27655), .Z(n27657) );
  XOR U27590 ( .A(n27661), .B(n27662), .Z(n26831) );
  AND U27591 ( .A(n607), .B(n27663), .Z(n27662) );
  XOR U27592 ( .A(p_input[294]), .B(p_input[262]), .Z(n27663) );
  XOR U27593 ( .A(n27664), .B(n27665), .Z(n27655) );
  AND U27594 ( .A(n27666), .B(n27667), .Z(n27665) );
  XOR U27595 ( .A(n27664), .B(n26846), .Z(n27667) );
  XNOR U27596 ( .A(p_input[325]), .B(n27668), .Z(n26846) );
  AND U27597 ( .A(n610), .B(n27669), .Z(n27668) );
  XOR U27598 ( .A(p_input[357]), .B(p_input[325]), .Z(n27669) );
  XNOR U27599 ( .A(n26843), .B(n27664), .Z(n27666) );
  XOR U27600 ( .A(n27670), .B(n27671), .Z(n26843) );
  AND U27601 ( .A(n607), .B(n27672), .Z(n27671) );
  XOR U27602 ( .A(p_input[293]), .B(p_input[261]), .Z(n27672) );
  XOR U27603 ( .A(n27673), .B(n27674), .Z(n27664) );
  AND U27604 ( .A(n27675), .B(n27676), .Z(n27674) );
  XOR U27605 ( .A(n27673), .B(n26858), .Z(n27676) );
  XNOR U27606 ( .A(p_input[324]), .B(n27677), .Z(n26858) );
  AND U27607 ( .A(n610), .B(n27678), .Z(n27677) );
  XOR U27608 ( .A(p_input[356]), .B(p_input[324]), .Z(n27678) );
  XNOR U27609 ( .A(n26855), .B(n27673), .Z(n27675) );
  XOR U27610 ( .A(n27679), .B(n27680), .Z(n26855) );
  AND U27611 ( .A(n607), .B(n27681), .Z(n27680) );
  XOR U27612 ( .A(p_input[292]), .B(p_input[260]), .Z(n27681) );
  XOR U27613 ( .A(n27682), .B(n27683), .Z(n27673) );
  AND U27614 ( .A(n27684), .B(n27685), .Z(n27683) );
  XOR U27615 ( .A(n27682), .B(n26870), .Z(n27685) );
  XNOR U27616 ( .A(p_input[323]), .B(n27686), .Z(n26870) );
  AND U27617 ( .A(n610), .B(n27687), .Z(n27686) );
  XOR U27618 ( .A(p_input[355]), .B(p_input[323]), .Z(n27687) );
  XNOR U27619 ( .A(n26867), .B(n27682), .Z(n27684) );
  XOR U27620 ( .A(n27688), .B(n27689), .Z(n26867) );
  AND U27621 ( .A(n607), .B(n27690), .Z(n27689) );
  XOR U27622 ( .A(p_input[291]), .B(p_input[259]), .Z(n27690) );
  XOR U27623 ( .A(n27691), .B(n27692), .Z(n27682) );
  AND U27624 ( .A(n27693), .B(n27694), .Z(n27692) );
  XOR U27625 ( .A(n26882), .B(n27691), .Z(n27694) );
  XNOR U27626 ( .A(p_input[322]), .B(n27695), .Z(n26882) );
  AND U27627 ( .A(n610), .B(n27696), .Z(n27695) );
  XOR U27628 ( .A(p_input[354]), .B(p_input[322]), .Z(n27696) );
  XNOR U27629 ( .A(n27691), .B(n26879), .Z(n27693) );
  XOR U27630 ( .A(n27697), .B(n27698), .Z(n26879) );
  AND U27631 ( .A(n607), .B(n27699), .Z(n27698) );
  XOR U27632 ( .A(p_input[290]), .B(p_input[258]), .Z(n27699) );
  XOR U27633 ( .A(n27700), .B(n27701), .Z(n27691) );
  AND U27634 ( .A(n27702), .B(n27703), .Z(n27701) );
  XNOR U27635 ( .A(n27704), .B(n26895), .Z(n27703) );
  XNOR U27636 ( .A(p_input[321]), .B(n27705), .Z(n26895) );
  AND U27637 ( .A(n610), .B(n27706), .Z(n27705) );
  XNOR U27638 ( .A(p_input[353]), .B(n27707), .Z(n27706) );
  IV U27639 ( .A(p_input[321]), .Z(n27707) );
  XNOR U27640 ( .A(n26892), .B(n27700), .Z(n27702) );
  XNOR U27641 ( .A(p_input[257]), .B(n27708), .Z(n26892) );
  AND U27642 ( .A(n607), .B(n27709), .Z(n27708) );
  XOR U27643 ( .A(p_input[289]), .B(p_input[257]), .Z(n27709) );
  IV U27644 ( .A(n27704), .Z(n27700) );
  AND U27645 ( .A(n27430), .B(n27433), .Z(n27704) );
  XOR U27646 ( .A(p_input[320]), .B(n27710), .Z(n27433) );
  AND U27647 ( .A(n610), .B(n27711), .Z(n27710) );
  XOR U27648 ( .A(p_input[352]), .B(p_input[320]), .Z(n27711) );
  XOR U27649 ( .A(n27712), .B(n27713), .Z(n610) );
  AND U27650 ( .A(n27714), .B(n27715), .Z(n27713) );
  XNOR U27651 ( .A(p_input[383]), .B(n27712), .Z(n27715) );
  XOR U27652 ( .A(n27712), .B(p_input[351]), .Z(n27714) );
  XOR U27653 ( .A(n27716), .B(n27717), .Z(n27712) );
  AND U27654 ( .A(n27718), .B(n27719), .Z(n27717) );
  XNOR U27655 ( .A(p_input[382]), .B(n27716), .Z(n27719) );
  XOR U27656 ( .A(n27716), .B(p_input[350]), .Z(n27718) );
  XOR U27657 ( .A(n27720), .B(n27721), .Z(n27716) );
  AND U27658 ( .A(n27722), .B(n27723), .Z(n27721) );
  XNOR U27659 ( .A(p_input[381]), .B(n27720), .Z(n27723) );
  XOR U27660 ( .A(n27720), .B(p_input[349]), .Z(n27722) );
  XOR U27661 ( .A(n27724), .B(n27725), .Z(n27720) );
  AND U27662 ( .A(n27726), .B(n27727), .Z(n27725) );
  XNOR U27663 ( .A(p_input[380]), .B(n27724), .Z(n27727) );
  XOR U27664 ( .A(n27724), .B(p_input[348]), .Z(n27726) );
  XOR U27665 ( .A(n27728), .B(n27729), .Z(n27724) );
  AND U27666 ( .A(n27730), .B(n27731), .Z(n27729) );
  XNOR U27667 ( .A(p_input[379]), .B(n27728), .Z(n27731) );
  XOR U27668 ( .A(n27728), .B(p_input[347]), .Z(n27730) );
  XOR U27669 ( .A(n27732), .B(n27733), .Z(n27728) );
  AND U27670 ( .A(n27734), .B(n27735), .Z(n27733) );
  XNOR U27671 ( .A(p_input[378]), .B(n27732), .Z(n27735) );
  XOR U27672 ( .A(n27732), .B(p_input[346]), .Z(n27734) );
  XOR U27673 ( .A(n27736), .B(n27737), .Z(n27732) );
  AND U27674 ( .A(n27738), .B(n27739), .Z(n27737) );
  XNOR U27675 ( .A(p_input[377]), .B(n27736), .Z(n27739) );
  XOR U27676 ( .A(n27736), .B(p_input[345]), .Z(n27738) );
  XOR U27677 ( .A(n27740), .B(n27741), .Z(n27736) );
  AND U27678 ( .A(n27742), .B(n27743), .Z(n27741) );
  XNOR U27679 ( .A(p_input[376]), .B(n27740), .Z(n27743) );
  XOR U27680 ( .A(n27740), .B(p_input[344]), .Z(n27742) );
  XOR U27681 ( .A(n27744), .B(n27745), .Z(n27740) );
  AND U27682 ( .A(n27746), .B(n27747), .Z(n27745) );
  XNOR U27683 ( .A(p_input[375]), .B(n27744), .Z(n27747) );
  XOR U27684 ( .A(n27744), .B(p_input[343]), .Z(n27746) );
  XOR U27685 ( .A(n27748), .B(n27749), .Z(n27744) );
  AND U27686 ( .A(n27750), .B(n27751), .Z(n27749) );
  XNOR U27687 ( .A(p_input[374]), .B(n27748), .Z(n27751) );
  XOR U27688 ( .A(n27748), .B(p_input[342]), .Z(n27750) );
  XOR U27689 ( .A(n27752), .B(n27753), .Z(n27748) );
  AND U27690 ( .A(n27754), .B(n27755), .Z(n27753) );
  XNOR U27691 ( .A(p_input[373]), .B(n27752), .Z(n27755) );
  XOR U27692 ( .A(n27752), .B(p_input[341]), .Z(n27754) );
  XOR U27693 ( .A(n27756), .B(n27757), .Z(n27752) );
  AND U27694 ( .A(n27758), .B(n27759), .Z(n27757) );
  XNOR U27695 ( .A(p_input[372]), .B(n27756), .Z(n27759) );
  XOR U27696 ( .A(n27756), .B(p_input[340]), .Z(n27758) );
  XOR U27697 ( .A(n27760), .B(n27761), .Z(n27756) );
  AND U27698 ( .A(n27762), .B(n27763), .Z(n27761) );
  XNOR U27699 ( .A(p_input[371]), .B(n27760), .Z(n27763) );
  XOR U27700 ( .A(n27760), .B(p_input[339]), .Z(n27762) );
  XOR U27701 ( .A(n27764), .B(n27765), .Z(n27760) );
  AND U27702 ( .A(n27766), .B(n27767), .Z(n27765) );
  XNOR U27703 ( .A(p_input[370]), .B(n27764), .Z(n27767) );
  XOR U27704 ( .A(n27764), .B(p_input[338]), .Z(n27766) );
  XOR U27705 ( .A(n27768), .B(n27769), .Z(n27764) );
  AND U27706 ( .A(n27770), .B(n27771), .Z(n27769) );
  XNOR U27707 ( .A(p_input[369]), .B(n27768), .Z(n27771) );
  XOR U27708 ( .A(n27768), .B(p_input[337]), .Z(n27770) );
  XOR U27709 ( .A(n27772), .B(n27773), .Z(n27768) );
  AND U27710 ( .A(n27774), .B(n27775), .Z(n27773) );
  XNOR U27711 ( .A(p_input[368]), .B(n27772), .Z(n27775) );
  XOR U27712 ( .A(n27772), .B(p_input[336]), .Z(n27774) );
  XOR U27713 ( .A(n27776), .B(n27777), .Z(n27772) );
  AND U27714 ( .A(n27778), .B(n27779), .Z(n27777) );
  XNOR U27715 ( .A(p_input[367]), .B(n27776), .Z(n27779) );
  XOR U27716 ( .A(n27776), .B(p_input[335]), .Z(n27778) );
  XOR U27717 ( .A(n27780), .B(n27781), .Z(n27776) );
  AND U27718 ( .A(n27782), .B(n27783), .Z(n27781) );
  XNOR U27719 ( .A(p_input[366]), .B(n27780), .Z(n27783) );
  XOR U27720 ( .A(n27780), .B(p_input[334]), .Z(n27782) );
  XOR U27721 ( .A(n27784), .B(n27785), .Z(n27780) );
  AND U27722 ( .A(n27786), .B(n27787), .Z(n27785) );
  XNOR U27723 ( .A(p_input[365]), .B(n27784), .Z(n27787) );
  XOR U27724 ( .A(n27784), .B(p_input[333]), .Z(n27786) );
  XOR U27725 ( .A(n27788), .B(n27789), .Z(n27784) );
  AND U27726 ( .A(n27790), .B(n27791), .Z(n27789) );
  XNOR U27727 ( .A(p_input[364]), .B(n27788), .Z(n27791) );
  XOR U27728 ( .A(n27788), .B(p_input[332]), .Z(n27790) );
  XOR U27729 ( .A(n27792), .B(n27793), .Z(n27788) );
  AND U27730 ( .A(n27794), .B(n27795), .Z(n27793) );
  XNOR U27731 ( .A(p_input[363]), .B(n27792), .Z(n27795) );
  XOR U27732 ( .A(n27792), .B(p_input[331]), .Z(n27794) );
  XOR U27733 ( .A(n27796), .B(n27797), .Z(n27792) );
  AND U27734 ( .A(n27798), .B(n27799), .Z(n27797) );
  XNOR U27735 ( .A(p_input[362]), .B(n27796), .Z(n27799) );
  XOR U27736 ( .A(n27796), .B(p_input[330]), .Z(n27798) );
  XOR U27737 ( .A(n27800), .B(n27801), .Z(n27796) );
  AND U27738 ( .A(n27802), .B(n27803), .Z(n27801) );
  XNOR U27739 ( .A(p_input[361]), .B(n27800), .Z(n27803) );
  XOR U27740 ( .A(n27800), .B(p_input[329]), .Z(n27802) );
  XOR U27741 ( .A(n27804), .B(n27805), .Z(n27800) );
  AND U27742 ( .A(n27806), .B(n27807), .Z(n27805) );
  XNOR U27743 ( .A(p_input[360]), .B(n27804), .Z(n27807) );
  XOR U27744 ( .A(n27804), .B(p_input[328]), .Z(n27806) );
  XOR U27745 ( .A(n27808), .B(n27809), .Z(n27804) );
  AND U27746 ( .A(n27810), .B(n27811), .Z(n27809) );
  XNOR U27747 ( .A(p_input[359]), .B(n27808), .Z(n27811) );
  XOR U27748 ( .A(n27808), .B(p_input[327]), .Z(n27810) );
  XOR U27749 ( .A(n27812), .B(n27813), .Z(n27808) );
  AND U27750 ( .A(n27814), .B(n27815), .Z(n27813) );
  XNOR U27751 ( .A(p_input[358]), .B(n27812), .Z(n27815) );
  XOR U27752 ( .A(n27812), .B(p_input[326]), .Z(n27814) );
  XOR U27753 ( .A(n27816), .B(n27817), .Z(n27812) );
  AND U27754 ( .A(n27818), .B(n27819), .Z(n27817) );
  XNOR U27755 ( .A(p_input[357]), .B(n27816), .Z(n27819) );
  XOR U27756 ( .A(n27816), .B(p_input[325]), .Z(n27818) );
  XOR U27757 ( .A(n27820), .B(n27821), .Z(n27816) );
  AND U27758 ( .A(n27822), .B(n27823), .Z(n27821) );
  XNOR U27759 ( .A(p_input[356]), .B(n27820), .Z(n27823) );
  XOR U27760 ( .A(n27820), .B(p_input[324]), .Z(n27822) );
  XOR U27761 ( .A(n27824), .B(n27825), .Z(n27820) );
  AND U27762 ( .A(n27826), .B(n27827), .Z(n27825) );
  XNOR U27763 ( .A(p_input[355]), .B(n27824), .Z(n27827) );
  XOR U27764 ( .A(n27824), .B(p_input[323]), .Z(n27826) );
  XOR U27765 ( .A(n27828), .B(n27829), .Z(n27824) );
  AND U27766 ( .A(n27830), .B(n27831), .Z(n27829) );
  XNOR U27767 ( .A(p_input[354]), .B(n27828), .Z(n27831) );
  XOR U27768 ( .A(n27828), .B(p_input[322]), .Z(n27830) );
  XNOR U27769 ( .A(n27832), .B(n27833), .Z(n27828) );
  AND U27770 ( .A(n27834), .B(n27835), .Z(n27833) );
  XOR U27771 ( .A(p_input[353]), .B(n27832), .Z(n27835) );
  XNOR U27772 ( .A(p_input[321]), .B(n27832), .Z(n27834) );
  AND U27773 ( .A(p_input[352]), .B(n27836), .Z(n27832) );
  IV U27774 ( .A(p_input[320]), .Z(n27836) );
  XNOR U27775 ( .A(p_input[256]), .B(n27837), .Z(n27430) );
  AND U27776 ( .A(n607), .B(n27838), .Z(n27837) );
  XOR U27777 ( .A(p_input[288]), .B(p_input[256]), .Z(n27838) );
  XOR U27778 ( .A(n27839), .B(n27840), .Z(n607) );
  AND U27779 ( .A(n27841), .B(n27842), .Z(n27840) );
  XNOR U27780 ( .A(p_input[319]), .B(n27839), .Z(n27842) );
  XOR U27781 ( .A(n27839), .B(p_input[287]), .Z(n27841) );
  XOR U27782 ( .A(n27843), .B(n27844), .Z(n27839) );
  AND U27783 ( .A(n27845), .B(n27846), .Z(n27844) );
  XNOR U27784 ( .A(p_input[318]), .B(n27843), .Z(n27846) );
  XNOR U27785 ( .A(n27843), .B(n27445), .Z(n27845) );
  IV U27786 ( .A(p_input[286]), .Z(n27445) );
  XOR U27787 ( .A(n27847), .B(n27848), .Z(n27843) );
  AND U27788 ( .A(n27849), .B(n27850), .Z(n27848) );
  XNOR U27789 ( .A(p_input[317]), .B(n27847), .Z(n27850) );
  XNOR U27790 ( .A(n27847), .B(n27454), .Z(n27849) );
  IV U27791 ( .A(p_input[285]), .Z(n27454) );
  XOR U27792 ( .A(n27851), .B(n27852), .Z(n27847) );
  AND U27793 ( .A(n27853), .B(n27854), .Z(n27852) );
  XNOR U27794 ( .A(p_input[316]), .B(n27851), .Z(n27854) );
  XNOR U27795 ( .A(n27851), .B(n27463), .Z(n27853) );
  IV U27796 ( .A(p_input[284]), .Z(n27463) );
  XOR U27797 ( .A(n27855), .B(n27856), .Z(n27851) );
  AND U27798 ( .A(n27857), .B(n27858), .Z(n27856) );
  XNOR U27799 ( .A(p_input[315]), .B(n27855), .Z(n27858) );
  XNOR U27800 ( .A(n27855), .B(n27472), .Z(n27857) );
  IV U27801 ( .A(p_input[283]), .Z(n27472) );
  XOR U27802 ( .A(n27859), .B(n27860), .Z(n27855) );
  AND U27803 ( .A(n27861), .B(n27862), .Z(n27860) );
  XNOR U27804 ( .A(p_input[314]), .B(n27859), .Z(n27862) );
  XNOR U27805 ( .A(n27859), .B(n27481), .Z(n27861) );
  IV U27806 ( .A(p_input[282]), .Z(n27481) );
  XOR U27807 ( .A(n27863), .B(n27864), .Z(n27859) );
  AND U27808 ( .A(n27865), .B(n27866), .Z(n27864) );
  XNOR U27809 ( .A(p_input[313]), .B(n27863), .Z(n27866) );
  XNOR U27810 ( .A(n27863), .B(n27490), .Z(n27865) );
  IV U27811 ( .A(p_input[281]), .Z(n27490) );
  XOR U27812 ( .A(n27867), .B(n27868), .Z(n27863) );
  AND U27813 ( .A(n27869), .B(n27870), .Z(n27868) );
  XNOR U27814 ( .A(p_input[312]), .B(n27867), .Z(n27870) );
  XNOR U27815 ( .A(n27867), .B(n27499), .Z(n27869) );
  IV U27816 ( .A(p_input[280]), .Z(n27499) );
  XOR U27817 ( .A(n27871), .B(n27872), .Z(n27867) );
  AND U27818 ( .A(n27873), .B(n27874), .Z(n27872) );
  XNOR U27819 ( .A(p_input[311]), .B(n27871), .Z(n27874) );
  XNOR U27820 ( .A(n27871), .B(n27508), .Z(n27873) );
  IV U27821 ( .A(p_input[279]), .Z(n27508) );
  XOR U27822 ( .A(n27875), .B(n27876), .Z(n27871) );
  AND U27823 ( .A(n27877), .B(n27878), .Z(n27876) );
  XNOR U27824 ( .A(p_input[310]), .B(n27875), .Z(n27878) );
  XNOR U27825 ( .A(n27875), .B(n27517), .Z(n27877) );
  IV U27826 ( .A(p_input[278]), .Z(n27517) );
  XOR U27827 ( .A(n27879), .B(n27880), .Z(n27875) );
  AND U27828 ( .A(n27881), .B(n27882), .Z(n27880) );
  XNOR U27829 ( .A(p_input[309]), .B(n27879), .Z(n27882) );
  XNOR U27830 ( .A(n27879), .B(n27526), .Z(n27881) );
  IV U27831 ( .A(p_input[277]), .Z(n27526) );
  XOR U27832 ( .A(n27883), .B(n27884), .Z(n27879) );
  AND U27833 ( .A(n27885), .B(n27886), .Z(n27884) );
  XNOR U27834 ( .A(p_input[308]), .B(n27883), .Z(n27886) );
  XNOR U27835 ( .A(n27883), .B(n27535), .Z(n27885) );
  IV U27836 ( .A(p_input[276]), .Z(n27535) );
  XOR U27837 ( .A(n27887), .B(n27888), .Z(n27883) );
  AND U27838 ( .A(n27889), .B(n27890), .Z(n27888) );
  XNOR U27839 ( .A(p_input[307]), .B(n27887), .Z(n27890) );
  XNOR U27840 ( .A(n27887), .B(n27544), .Z(n27889) );
  IV U27841 ( .A(p_input[275]), .Z(n27544) );
  XOR U27842 ( .A(n27891), .B(n27892), .Z(n27887) );
  AND U27843 ( .A(n27893), .B(n27894), .Z(n27892) );
  XNOR U27844 ( .A(p_input[306]), .B(n27891), .Z(n27894) );
  XNOR U27845 ( .A(n27891), .B(n27553), .Z(n27893) );
  IV U27846 ( .A(p_input[274]), .Z(n27553) );
  XOR U27847 ( .A(n27895), .B(n27896), .Z(n27891) );
  AND U27848 ( .A(n27897), .B(n27898), .Z(n27896) );
  XNOR U27849 ( .A(p_input[305]), .B(n27895), .Z(n27898) );
  XNOR U27850 ( .A(n27895), .B(n27562), .Z(n27897) );
  IV U27851 ( .A(p_input[273]), .Z(n27562) );
  XOR U27852 ( .A(n27899), .B(n27900), .Z(n27895) );
  AND U27853 ( .A(n27901), .B(n27902), .Z(n27900) );
  XNOR U27854 ( .A(p_input[304]), .B(n27899), .Z(n27902) );
  XNOR U27855 ( .A(n27899), .B(n27571), .Z(n27901) );
  IV U27856 ( .A(p_input[272]), .Z(n27571) );
  XOR U27857 ( .A(n27903), .B(n27904), .Z(n27899) );
  AND U27858 ( .A(n27905), .B(n27906), .Z(n27904) );
  XNOR U27859 ( .A(p_input[303]), .B(n27903), .Z(n27906) );
  XNOR U27860 ( .A(n27903), .B(n27580), .Z(n27905) );
  IV U27861 ( .A(p_input[271]), .Z(n27580) );
  XOR U27862 ( .A(n27907), .B(n27908), .Z(n27903) );
  AND U27863 ( .A(n27909), .B(n27910), .Z(n27908) );
  XNOR U27864 ( .A(p_input[302]), .B(n27907), .Z(n27910) );
  XNOR U27865 ( .A(n27907), .B(n27589), .Z(n27909) );
  IV U27866 ( .A(p_input[270]), .Z(n27589) );
  XOR U27867 ( .A(n27911), .B(n27912), .Z(n27907) );
  AND U27868 ( .A(n27913), .B(n27914), .Z(n27912) );
  XNOR U27869 ( .A(p_input[301]), .B(n27911), .Z(n27914) );
  XNOR U27870 ( .A(n27911), .B(n27598), .Z(n27913) );
  IV U27871 ( .A(p_input[269]), .Z(n27598) );
  XOR U27872 ( .A(n27915), .B(n27916), .Z(n27911) );
  AND U27873 ( .A(n27917), .B(n27918), .Z(n27916) );
  XNOR U27874 ( .A(p_input[300]), .B(n27915), .Z(n27918) );
  XNOR U27875 ( .A(n27915), .B(n27607), .Z(n27917) );
  IV U27876 ( .A(p_input[268]), .Z(n27607) );
  XOR U27877 ( .A(n27919), .B(n27920), .Z(n27915) );
  AND U27878 ( .A(n27921), .B(n27922), .Z(n27920) );
  XNOR U27879 ( .A(p_input[299]), .B(n27919), .Z(n27922) );
  XNOR U27880 ( .A(n27919), .B(n27616), .Z(n27921) );
  IV U27881 ( .A(p_input[267]), .Z(n27616) );
  XOR U27882 ( .A(n27923), .B(n27924), .Z(n27919) );
  AND U27883 ( .A(n27925), .B(n27926), .Z(n27924) );
  XNOR U27884 ( .A(p_input[298]), .B(n27923), .Z(n27926) );
  XNOR U27885 ( .A(n27923), .B(n27625), .Z(n27925) );
  IV U27886 ( .A(p_input[266]), .Z(n27625) );
  XOR U27887 ( .A(n27927), .B(n27928), .Z(n27923) );
  AND U27888 ( .A(n27929), .B(n27930), .Z(n27928) );
  XNOR U27889 ( .A(p_input[297]), .B(n27927), .Z(n27930) );
  XNOR U27890 ( .A(n27927), .B(n27634), .Z(n27929) );
  IV U27891 ( .A(p_input[265]), .Z(n27634) );
  XOR U27892 ( .A(n27931), .B(n27932), .Z(n27927) );
  AND U27893 ( .A(n27933), .B(n27934), .Z(n27932) );
  XNOR U27894 ( .A(p_input[296]), .B(n27931), .Z(n27934) );
  XNOR U27895 ( .A(n27931), .B(n27643), .Z(n27933) );
  IV U27896 ( .A(p_input[264]), .Z(n27643) );
  XOR U27897 ( .A(n27935), .B(n27936), .Z(n27931) );
  AND U27898 ( .A(n27937), .B(n27938), .Z(n27936) );
  XNOR U27899 ( .A(p_input[295]), .B(n27935), .Z(n27938) );
  XNOR U27900 ( .A(n27935), .B(n27652), .Z(n27937) );
  IV U27901 ( .A(p_input[263]), .Z(n27652) );
  XOR U27902 ( .A(n27939), .B(n27940), .Z(n27935) );
  AND U27903 ( .A(n27941), .B(n27942), .Z(n27940) );
  XNOR U27904 ( .A(p_input[294]), .B(n27939), .Z(n27942) );
  XNOR U27905 ( .A(n27939), .B(n27661), .Z(n27941) );
  IV U27906 ( .A(p_input[262]), .Z(n27661) );
  XOR U27907 ( .A(n27943), .B(n27944), .Z(n27939) );
  AND U27908 ( .A(n27945), .B(n27946), .Z(n27944) );
  XNOR U27909 ( .A(p_input[293]), .B(n27943), .Z(n27946) );
  XNOR U27910 ( .A(n27943), .B(n27670), .Z(n27945) );
  IV U27911 ( .A(p_input[261]), .Z(n27670) );
  XOR U27912 ( .A(n27947), .B(n27948), .Z(n27943) );
  AND U27913 ( .A(n27949), .B(n27950), .Z(n27948) );
  XNOR U27914 ( .A(p_input[292]), .B(n27947), .Z(n27950) );
  XNOR U27915 ( .A(n27947), .B(n27679), .Z(n27949) );
  IV U27916 ( .A(p_input[260]), .Z(n27679) );
  XOR U27917 ( .A(n27951), .B(n27952), .Z(n27947) );
  AND U27918 ( .A(n27953), .B(n27954), .Z(n27952) );
  XNOR U27919 ( .A(p_input[291]), .B(n27951), .Z(n27954) );
  XNOR U27920 ( .A(n27951), .B(n27688), .Z(n27953) );
  IV U27921 ( .A(p_input[259]), .Z(n27688) );
  XOR U27922 ( .A(n27955), .B(n27956), .Z(n27951) );
  AND U27923 ( .A(n27957), .B(n27958), .Z(n27956) );
  XNOR U27924 ( .A(p_input[290]), .B(n27955), .Z(n27958) );
  XNOR U27925 ( .A(n27955), .B(n27697), .Z(n27957) );
  IV U27926 ( .A(p_input[258]), .Z(n27697) );
  XNOR U27927 ( .A(n27959), .B(n27960), .Z(n27955) );
  AND U27928 ( .A(n27961), .B(n27962), .Z(n27960) );
  XOR U27929 ( .A(p_input[289]), .B(n27959), .Z(n27962) );
  XNOR U27930 ( .A(p_input[257]), .B(n27959), .Z(n27961) );
  AND U27931 ( .A(p_input[288]), .B(n27963), .Z(n27959) );
  IV U27932 ( .A(p_input[256]), .Z(n27963) );
  XOR U27933 ( .A(n27964), .B(n27965), .Z(n26142) );
  AND U27934 ( .A(n531), .B(n27966), .Z(n27965) );
  XNOR U27935 ( .A(n27967), .B(n27964), .Z(n27966) );
  XOR U27936 ( .A(n27968), .B(n27969), .Z(n531) );
  AND U27937 ( .A(n27970), .B(n27971), .Z(n27969) );
  XOR U27938 ( .A(n27968), .B(n26157), .Z(n27971) );
  XNOR U27939 ( .A(n27972), .B(n27973), .Z(n26157) );
  AND U27940 ( .A(n27974), .B(n410), .Z(n27973) );
  AND U27941 ( .A(n27972), .B(n27975), .Z(n27974) );
  XNOR U27942 ( .A(n26154), .B(n27968), .Z(n27970) );
  XOR U27943 ( .A(n27976), .B(n27977), .Z(n26154) );
  AND U27944 ( .A(n27978), .B(n407), .Z(n27977) );
  NOR U27945 ( .A(n27976), .B(n27979), .Z(n27978) );
  XOR U27946 ( .A(n27980), .B(n27981), .Z(n27968) );
  AND U27947 ( .A(n27982), .B(n27983), .Z(n27981) );
  XOR U27948 ( .A(n27980), .B(n26169), .Z(n27983) );
  XOR U27949 ( .A(n27984), .B(n27985), .Z(n26169) );
  AND U27950 ( .A(n410), .B(n27986), .Z(n27985) );
  XOR U27951 ( .A(n27987), .B(n27984), .Z(n27986) );
  XNOR U27952 ( .A(n26166), .B(n27980), .Z(n27982) );
  XOR U27953 ( .A(n27988), .B(n27989), .Z(n26166) );
  AND U27954 ( .A(n407), .B(n27990), .Z(n27989) );
  XOR U27955 ( .A(n27991), .B(n27988), .Z(n27990) );
  XOR U27956 ( .A(n27992), .B(n27993), .Z(n27980) );
  AND U27957 ( .A(n27994), .B(n27995), .Z(n27993) );
  XOR U27958 ( .A(n27992), .B(n26181), .Z(n27995) );
  XOR U27959 ( .A(n27996), .B(n27997), .Z(n26181) );
  AND U27960 ( .A(n410), .B(n27998), .Z(n27997) );
  XOR U27961 ( .A(n27999), .B(n27996), .Z(n27998) );
  XNOR U27962 ( .A(n26178), .B(n27992), .Z(n27994) );
  XOR U27963 ( .A(n28000), .B(n28001), .Z(n26178) );
  AND U27964 ( .A(n407), .B(n28002), .Z(n28001) );
  XOR U27965 ( .A(n28003), .B(n28000), .Z(n28002) );
  XOR U27966 ( .A(n28004), .B(n28005), .Z(n27992) );
  AND U27967 ( .A(n28006), .B(n28007), .Z(n28005) );
  XOR U27968 ( .A(n28004), .B(n26193), .Z(n28007) );
  XOR U27969 ( .A(n28008), .B(n28009), .Z(n26193) );
  AND U27970 ( .A(n410), .B(n28010), .Z(n28009) );
  XOR U27971 ( .A(n28011), .B(n28008), .Z(n28010) );
  XNOR U27972 ( .A(n26190), .B(n28004), .Z(n28006) );
  XOR U27973 ( .A(n28012), .B(n28013), .Z(n26190) );
  AND U27974 ( .A(n407), .B(n28014), .Z(n28013) );
  XOR U27975 ( .A(n28015), .B(n28012), .Z(n28014) );
  XOR U27976 ( .A(n28016), .B(n28017), .Z(n28004) );
  AND U27977 ( .A(n28018), .B(n28019), .Z(n28017) );
  XOR U27978 ( .A(n28016), .B(n26205), .Z(n28019) );
  XOR U27979 ( .A(n28020), .B(n28021), .Z(n26205) );
  AND U27980 ( .A(n410), .B(n28022), .Z(n28021) );
  XOR U27981 ( .A(n28023), .B(n28020), .Z(n28022) );
  XNOR U27982 ( .A(n26202), .B(n28016), .Z(n28018) );
  XOR U27983 ( .A(n28024), .B(n28025), .Z(n26202) );
  AND U27984 ( .A(n407), .B(n28026), .Z(n28025) );
  XOR U27985 ( .A(n28027), .B(n28024), .Z(n28026) );
  XOR U27986 ( .A(n28028), .B(n28029), .Z(n28016) );
  AND U27987 ( .A(n28030), .B(n28031), .Z(n28029) );
  XOR U27988 ( .A(n28028), .B(n26217), .Z(n28031) );
  XOR U27989 ( .A(n28032), .B(n28033), .Z(n26217) );
  AND U27990 ( .A(n410), .B(n28034), .Z(n28033) );
  XOR U27991 ( .A(n28035), .B(n28032), .Z(n28034) );
  XNOR U27992 ( .A(n26214), .B(n28028), .Z(n28030) );
  XOR U27993 ( .A(n28036), .B(n28037), .Z(n26214) );
  AND U27994 ( .A(n407), .B(n28038), .Z(n28037) );
  XOR U27995 ( .A(n28039), .B(n28036), .Z(n28038) );
  XOR U27996 ( .A(n28040), .B(n28041), .Z(n28028) );
  AND U27997 ( .A(n28042), .B(n28043), .Z(n28041) );
  XOR U27998 ( .A(n28040), .B(n26229), .Z(n28043) );
  XOR U27999 ( .A(n28044), .B(n28045), .Z(n26229) );
  AND U28000 ( .A(n410), .B(n28046), .Z(n28045) );
  XOR U28001 ( .A(n28047), .B(n28044), .Z(n28046) );
  XNOR U28002 ( .A(n26226), .B(n28040), .Z(n28042) );
  XOR U28003 ( .A(n28048), .B(n28049), .Z(n26226) );
  AND U28004 ( .A(n407), .B(n28050), .Z(n28049) );
  XOR U28005 ( .A(n28051), .B(n28048), .Z(n28050) );
  XOR U28006 ( .A(n28052), .B(n28053), .Z(n28040) );
  AND U28007 ( .A(n28054), .B(n28055), .Z(n28053) );
  XOR U28008 ( .A(n28052), .B(n26241), .Z(n28055) );
  XOR U28009 ( .A(n28056), .B(n28057), .Z(n26241) );
  AND U28010 ( .A(n410), .B(n28058), .Z(n28057) );
  XOR U28011 ( .A(n28059), .B(n28056), .Z(n28058) );
  XNOR U28012 ( .A(n26238), .B(n28052), .Z(n28054) );
  XOR U28013 ( .A(n28060), .B(n28061), .Z(n26238) );
  AND U28014 ( .A(n407), .B(n28062), .Z(n28061) );
  XOR U28015 ( .A(n28063), .B(n28060), .Z(n28062) );
  XOR U28016 ( .A(n28064), .B(n28065), .Z(n28052) );
  AND U28017 ( .A(n28066), .B(n28067), .Z(n28065) );
  XOR U28018 ( .A(n28064), .B(n26253), .Z(n28067) );
  XOR U28019 ( .A(n28068), .B(n28069), .Z(n26253) );
  AND U28020 ( .A(n410), .B(n28070), .Z(n28069) );
  XOR U28021 ( .A(n28071), .B(n28068), .Z(n28070) );
  XNOR U28022 ( .A(n26250), .B(n28064), .Z(n28066) );
  XOR U28023 ( .A(n28072), .B(n28073), .Z(n26250) );
  AND U28024 ( .A(n407), .B(n28074), .Z(n28073) );
  XOR U28025 ( .A(n28075), .B(n28072), .Z(n28074) );
  XOR U28026 ( .A(n28076), .B(n28077), .Z(n28064) );
  AND U28027 ( .A(n28078), .B(n28079), .Z(n28077) );
  XOR U28028 ( .A(n28076), .B(n26265), .Z(n28079) );
  XOR U28029 ( .A(n28080), .B(n28081), .Z(n26265) );
  AND U28030 ( .A(n410), .B(n28082), .Z(n28081) );
  XOR U28031 ( .A(n28083), .B(n28080), .Z(n28082) );
  XNOR U28032 ( .A(n26262), .B(n28076), .Z(n28078) );
  XOR U28033 ( .A(n28084), .B(n28085), .Z(n26262) );
  AND U28034 ( .A(n407), .B(n28086), .Z(n28085) );
  XOR U28035 ( .A(n28087), .B(n28084), .Z(n28086) );
  XOR U28036 ( .A(n28088), .B(n28089), .Z(n28076) );
  AND U28037 ( .A(n28090), .B(n28091), .Z(n28089) );
  XOR U28038 ( .A(n28088), .B(n26277), .Z(n28091) );
  XOR U28039 ( .A(n28092), .B(n28093), .Z(n26277) );
  AND U28040 ( .A(n410), .B(n28094), .Z(n28093) );
  XOR U28041 ( .A(n28095), .B(n28092), .Z(n28094) );
  XNOR U28042 ( .A(n26274), .B(n28088), .Z(n28090) );
  XOR U28043 ( .A(n28096), .B(n28097), .Z(n26274) );
  AND U28044 ( .A(n407), .B(n28098), .Z(n28097) );
  XOR U28045 ( .A(n28099), .B(n28096), .Z(n28098) );
  XOR U28046 ( .A(n28100), .B(n28101), .Z(n28088) );
  AND U28047 ( .A(n28102), .B(n28103), .Z(n28101) );
  XOR U28048 ( .A(n28100), .B(n26289), .Z(n28103) );
  XOR U28049 ( .A(n28104), .B(n28105), .Z(n26289) );
  AND U28050 ( .A(n410), .B(n28106), .Z(n28105) );
  XOR U28051 ( .A(n28107), .B(n28104), .Z(n28106) );
  XNOR U28052 ( .A(n26286), .B(n28100), .Z(n28102) );
  XOR U28053 ( .A(n28108), .B(n28109), .Z(n26286) );
  AND U28054 ( .A(n407), .B(n28110), .Z(n28109) );
  XOR U28055 ( .A(n28111), .B(n28108), .Z(n28110) );
  XOR U28056 ( .A(n28112), .B(n28113), .Z(n28100) );
  AND U28057 ( .A(n28114), .B(n28115), .Z(n28113) );
  XOR U28058 ( .A(n28112), .B(n26301), .Z(n28115) );
  XOR U28059 ( .A(n28116), .B(n28117), .Z(n26301) );
  AND U28060 ( .A(n410), .B(n28118), .Z(n28117) );
  XOR U28061 ( .A(n28119), .B(n28116), .Z(n28118) );
  XNOR U28062 ( .A(n26298), .B(n28112), .Z(n28114) );
  XOR U28063 ( .A(n28120), .B(n28121), .Z(n26298) );
  AND U28064 ( .A(n407), .B(n28122), .Z(n28121) );
  XOR U28065 ( .A(n28123), .B(n28120), .Z(n28122) );
  XOR U28066 ( .A(n28124), .B(n28125), .Z(n28112) );
  AND U28067 ( .A(n28126), .B(n28127), .Z(n28125) );
  XOR U28068 ( .A(n28124), .B(n26313), .Z(n28127) );
  XOR U28069 ( .A(n28128), .B(n28129), .Z(n26313) );
  AND U28070 ( .A(n410), .B(n28130), .Z(n28129) );
  XOR U28071 ( .A(n28131), .B(n28128), .Z(n28130) );
  XNOR U28072 ( .A(n26310), .B(n28124), .Z(n28126) );
  XOR U28073 ( .A(n28132), .B(n28133), .Z(n26310) );
  AND U28074 ( .A(n407), .B(n28134), .Z(n28133) );
  XOR U28075 ( .A(n28135), .B(n28132), .Z(n28134) );
  XOR U28076 ( .A(n28136), .B(n28137), .Z(n28124) );
  AND U28077 ( .A(n28138), .B(n28139), .Z(n28137) );
  XOR U28078 ( .A(n28136), .B(n26325), .Z(n28139) );
  XOR U28079 ( .A(n28140), .B(n28141), .Z(n26325) );
  AND U28080 ( .A(n410), .B(n28142), .Z(n28141) );
  XOR U28081 ( .A(n28143), .B(n28140), .Z(n28142) );
  XNOR U28082 ( .A(n26322), .B(n28136), .Z(n28138) );
  XOR U28083 ( .A(n28144), .B(n28145), .Z(n26322) );
  AND U28084 ( .A(n407), .B(n28146), .Z(n28145) );
  XOR U28085 ( .A(n28147), .B(n28144), .Z(n28146) );
  XOR U28086 ( .A(n28148), .B(n28149), .Z(n28136) );
  AND U28087 ( .A(n28150), .B(n28151), .Z(n28149) );
  XOR U28088 ( .A(n28148), .B(n26337), .Z(n28151) );
  XOR U28089 ( .A(n28152), .B(n28153), .Z(n26337) );
  AND U28090 ( .A(n410), .B(n28154), .Z(n28153) );
  XOR U28091 ( .A(n28155), .B(n28152), .Z(n28154) );
  XNOR U28092 ( .A(n26334), .B(n28148), .Z(n28150) );
  XOR U28093 ( .A(n28156), .B(n28157), .Z(n26334) );
  AND U28094 ( .A(n407), .B(n28158), .Z(n28157) );
  XOR U28095 ( .A(n28159), .B(n28156), .Z(n28158) );
  XOR U28096 ( .A(n28160), .B(n28161), .Z(n28148) );
  AND U28097 ( .A(n28162), .B(n28163), .Z(n28161) );
  XOR U28098 ( .A(n28160), .B(n26349), .Z(n28163) );
  XOR U28099 ( .A(n28164), .B(n28165), .Z(n26349) );
  AND U28100 ( .A(n410), .B(n28166), .Z(n28165) );
  XOR U28101 ( .A(n28167), .B(n28164), .Z(n28166) );
  XNOR U28102 ( .A(n26346), .B(n28160), .Z(n28162) );
  XOR U28103 ( .A(n28168), .B(n28169), .Z(n26346) );
  AND U28104 ( .A(n407), .B(n28170), .Z(n28169) );
  XOR U28105 ( .A(n28171), .B(n28168), .Z(n28170) );
  XOR U28106 ( .A(n28172), .B(n28173), .Z(n28160) );
  AND U28107 ( .A(n28174), .B(n28175), .Z(n28173) );
  XOR U28108 ( .A(n28172), .B(n26361), .Z(n28175) );
  XOR U28109 ( .A(n28176), .B(n28177), .Z(n26361) );
  AND U28110 ( .A(n410), .B(n28178), .Z(n28177) );
  XOR U28111 ( .A(n28179), .B(n28176), .Z(n28178) );
  XNOR U28112 ( .A(n26358), .B(n28172), .Z(n28174) );
  XOR U28113 ( .A(n28180), .B(n28181), .Z(n26358) );
  AND U28114 ( .A(n407), .B(n28182), .Z(n28181) );
  XOR U28115 ( .A(n28183), .B(n28180), .Z(n28182) );
  XOR U28116 ( .A(n28184), .B(n28185), .Z(n28172) );
  AND U28117 ( .A(n28186), .B(n28187), .Z(n28185) );
  XOR U28118 ( .A(n28184), .B(n26373), .Z(n28187) );
  XOR U28119 ( .A(n28188), .B(n28189), .Z(n26373) );
  AND U28120 ( .A(n410), .B(n28190), .Z(n28189) );
  XOR U28121 ( .A(n28191), .B(n28188), .Z(n28190) );
  XNOR U28122 ( .A(n26370), .B(n28184), .Z(n28186) );
  XOR U28123 ( .A(n28192), .B(n28193), .Z(n26370) );
  AND U28124 ( .A(n407), .B(n28194), .Z(n28193) );
  XOR U28125 ( .A(n28195), .B(n28192), .Z(n28194) );
  XOR U28126 ( .A(n28196), .B(n28197), .Z(n28184) );
  AND U28127 ( .A(n28198), .B(n28199), .Z(n28197) );
  XOR U28128 ( .A(n28196), .B(n26385), .Z(n28199) );
  XOR U28129 ( .A(n28200), .B(n28201), .Z(n26385) );
  AND U28130 ( .A(n410), .B(n28202), .Z(n28201) );
  XOR U28131 ( .A(n28203), .B(n28200), .Z(n28202) );
  XNOR U28132 ( .A(n26382), .B(n28196), .Z(n28198) );
  XOR U28133 ( .A(n28204), .B(n28205), .Z(n26382) );
  AND U28134 ( .A(n407), .B(n28206), .Z(n28205) );
  XOR U28135 ( .A(n28207), .B(n28204), .Z(n28206) );
  XOR U28136 ( .A(n28208), .B(n28209), .Z(n28196) );
  AND U28137 ( .A(n28210), .B(n28211), .Z(n28209) );
  XOR U28138 ( .A(n28208), .B(n26397), .Z(n28211) );
  XOR U28139 ( .A(n28212), .B(n28213), .Z(n26397) );
  AND U28140 ( .A(n410), .B(n28214), .Z(n28213) );
  XOR U28141 ( .A(n28215), .B(n28212), .Z(n28214) );
  XNOR U28142 ( .A(n26394), .B(n28208), .Z(n28210) );
  XOR U28143 ( .A(n28216), .B(n28217), .Z(n26394) );
  AND U28144 ( .A(n407), .B(n28218), .Z(n28217) );
  XOR U28145 ( .A(n28219), .B(n28216), .Z(n28218) );
  XOR U28146 ( .A(n28220), .B(n28221), .Z(n28208) );
  AND U28147 ( .A(n28222), .B(n28223), .Z(n28221) );
  XOR U28148 ( .A(n28220), .B(n26409), .Z(n28223) );
  XOR U28149 ( .A(n28224), .B(n28225), .Z(n26409) );
  AND U28150 ( .A(n410), .B(n28226), .Z(n28225) );
  XOR U28151 ( .A(n28227), .B(n28224), .Z(n28226) );
  XNOR U28152 ( .A(n26406), .B(n28220), .Z(n28222) );
  XOR U28153 ( .A(n28228), .B(n28229), .Z(n26406) );
  AND U28154 ( .A(n407), .B(n28230), .Z(n28229) );
  XOR U28155 ( .A(n28231), .B(n28228), .Z(n28230) );
  XOR U28156 ( .A(n28232), .B(n28233), .Z(n28220) );
  AND U28157 ( .A(n28234), .B(n28235), .Z(n28233) );
  XOR U28158 ( .A(n28232), .B(n26421), .Z(n28235) );
  XOR U28159 ( .A(n28236), .B(n28237), .Z(n26421) );
  AND U28160 ( .A(n410), .B(n28238), .Z(n28237) );
  XOR U28161 ( .A(n28239), .B(n28236), .Z(n28238) );
  XNOR U28162 ( .A(n26418), .B(n28232), .Z(n28234) );
  XOR U28163 ( .A(n28240), .B(n28241), .Z(n26418) );
  AND U28164 ( .A(n407), .B(n28242), .Z(n28241) );
  XOR U28165 ( .A(n28243), .B(n28240), .Z(n28242) );
  XOR U28166 ( .A(n28244), .B(n28245), .Z(n28232) );
  AND U28167 ( .A(n28246), .B(n28247), .Z(n28245) );
  XOR U28168 ( .A(n28244), .B(n26433), .Z(n28247) );
  XOR U28169 ( .A(n28248), .B(n28249), .Z(n26433) );
  AND U28170 ( .A(n410), .B(n28250), .Z(n28249) );
  XOR U28171 ( .A(n28251), .B(n28248), .Z(n28250) );
  XNOR U28172 ( .A(n26430), .B(n28244), .Z(n28246) );
  XOR U28173 ( .A(n28252), .B(n28253), .Z(n26430) );
  AND U28174 ( .A(n407), .B(n28254), .Z(n28253) );
  XOR U28175 ( .A(n28255), .B(n28252), .Z(n28254) );
  XOR U28176 ( .A(n28256), .B(n28257), .Z(n28244) );
  AND U28177 ( .A(n28258), .B(n28259), .Z(n28257) );
  XOR U28178 ( .A(n28256), .B(n26445), .Z(n28259) );
  XOR U28179 ( .A(n28260), .B(n28261), .Z(n26445) );
  AND U28180 ( .A(n410), .B(n28262), .Z(n28261) );
  XOR U28181 ( .A(n28263), .B(n28260), .Z(n28262) );
  XNOR U28182 ( .A(n26442), .B(n28256), .Z(n28258) );
  XOR U28183 ( .A(n28264), .B(n28265), .Z(n26442) );
  AND U28184 ( .A(n407), .B(n28266), .Z(n28265) );
  XOR U28185 ( .A(n28267), .B(n28264), .Z(n28266) );
  XOR U28186 ( .A(n28268), .B(n28269), .Z(n28256) );
  AND U28187 ( .A(n28270), .B(n28271), .Z(n28269) );
  XOR U28188 ( .A(n28268), .B(n26457), .Z(n28271) );
  XOR U28189 ( .A(n28272), .B(n28273), .Z(n26457) );
  AND U28190 ( .A(n410), .B(n28274), .Z(n28273) );
  XOR U28191 ( .A(n28275), .B(n28272), .Z(n28274) );
  XNOR U28192 ( .A(n26454), .B(n28268), .Z(n28270) );
  XOR U28193 ( .A(n28276), .B(n28277), .Z(n26454) );
  AND U28194 ( .A(n407), .B(n28278), .Z(n28277) );
  XOR U28195 ( .A(n28279), .B(n28276), .Z(n28278) );
  XOR U28196 ( .A(n28280), .B(n28281), .Z(n28268) );
  AND U28197 ( .A(n28282), .B(n28283), .Z(n28281) );
  XOR U28198 ( .A(n28280), .B(n26469), .Z(n28283) );
  XOR U28199 ( .A(n28284), .B(n28285), .Z(n26469) );
  AND U28200 ( .A(n410), .B(n28286), .Z(n28285) );
  XOR U28201 ( .A(n28287), .B(n28284), .Z(n28286) );
  XNOR U28202 ( .A(n26466), .B(n28280), .Z(n28282) );
  XOR U28203 ( .A(n28288), .B(n28289), .Z(n26466) );
  AND U28204 ( .A(n407), .B(n28290), .Z(n28289) );
  XOR U28205 ( .A(n28291), .B(n28288), .Z(n28290) );
  XOR U28206 ( .A(n28292), .B(n28293), .Z(n28280) );
  AND U28207 ( .A(n28294), .B(n28295), .Z(n28293) );
  XOR U28208 ( .A(n28292), .B(n26481), .Z(n28295) );
  XOR U28209 ( .A(n28296), .B(n28297), .Z(n26481) );
  AND U28210 ( .A(n410), .B(n28298), .Z(n28297) );
  XOR U28211 ( .A(n28299), .B(n28296), .Z(n28298) );
  XNOR U28212 ( .A(n26478), .B(n28292), .Z(n28294) );
  XOR U28213 ( .A(n28300), .B(n28301), .Z(n26478) );
  AND U28214 ( .A(n407), .B(n28302), .Z(n28301) );
  XOR U28215 ( .A(n28303), .B(n28300), .Z(n28302) );
  XOR U28216 ( .A(n28304), .B(n28305), .Z(n28292) );
  AND U28217 ( .A(n28306), .B(n28307), .Z(n28305) );
  XOR U28218 ( .A(n28304), .B(n26493), .Z(n28307) );
  XOR U28219 ( .A(n28308), .B(n28309), .Z(n26493) );
  AND U28220 ( .A(n410), .B(n28310), .Z(n28309) );
  XOR U28221 ( .A(n28311), .B(n28308), .Z(n28310) );
  XNOR U28222 ( .A(n26490), .B(n28304), .Z(n28306) );
  XOR U28223 ( .A(n28312), .B(n28313), .Z(n26490) );
  AND U28224 ( .A(n407), .B(n28314), .Z(n28313) );
  XOR U28225 ( .A(n28315), .B(n28312), .Z(n28314) );
  XOR U28226 ( .A(n28316), .B(n28317), .Z(n28304) );
  AND U28227 ( .A(n28318), .B(n28319), .Z(n28317) );
  XOR U28228 ( .A(n26505), .B(n28316), .Z(n28319) );
  XOR U28229 ( .A(n28320), .B(n28321), .Z(n26505) );
  AND U28230 ( .A(n410), .B(n28322), .Z(n28321) );
  XOR U28231 ( .A(n28320), .B(n28323), .Z(n28322) );
  XNOR U28232 ( .A(n28316), .B(n26502), .Z(n28318) );
  XOR U28233 ( .A(n28324), .B(n28325), .Z(n26502) );
  AND U28234 ( .A(n407), .B(n28326), .Z(n28325) );
  XOR U28235 ( .A(n28324), .B(n28327), .Z(n28326) );
  XOR U28236 ( .A(n28328), .B(n28329), .Z(n28316) );
  AND U28237 ( .A(n28330), .B(n28331), .Z(n28329) );
  XNOR U28238 ( .A(n28332), .B(n26518), .Z(n28331) );
  XOR U28239 ( .A(n28333), .B(n28334), .Z(n26518) );
  AND U28240 ( .A(n410), .B(n28335), .Z(n28334) );
  XOR U28241 ( .A(n28336), .B(n28333), .Z(n28335) );
  XNOR U28242 ( .A(n26515), .B(n28328), .Z(n28330) );
  XOR U28243 ( .A(n28337), .B(n28338), .Z(n26515) );
  AND U28244 ( .A(n407), .B(n28339), .Z(n28338) );
  XOR U28245 ( .A(n28340), .B(n28337), .Z(n28339) );
  IV U28246 ( .A(n28332), .Z(n28328) );
  AND U28247 ( .A(n27964), .B(n27967), .Z(n28332) );
  XNOR U28248 ( .A(n28341), .B(n28342), .Z(n27967) );
  AND U28249 ( .A(n410), .B(n28343), .Z(n28342) );
  XNOR U28250 ( .A(n28344), .B(n28341), .Z(n28343) );
  XOR U28251 ( .A(n28345), .B(n28346), .Z(n410) );
  AND U28252 ( .A(n28347), .B(n28348), .Z(n28346) );
  XOR U28253 ( .A(n27975), .B(n28345), .Z(n28348) );
  IV U28254 ( .A(n28349), .Z(n27975) );
  AND U28255 ( .A(p_input[255]), .B(p_input[223]), .Z(n28349) );
  XOR U28256 ( .A(n28345), .B(n27972), .Z(n28347) );
  AND U28257 ( .A(p_input[159]), .B(p_input[191]), .Z(n27972) );
  XOR U28258 ( .A(n28350), .B(n28351), .Z(n28345) );
  AND U28259 ( .A(n28352), .B(n28353), .Z(n28351) );
  XOR U28260 ( .A(n28350), .B(n27987), .Z(n28353) );
  XNOR U28261 ( .A(p_input[222]), .B(n28354), .Z(n27987) );
  AND U28262 ( .A(n630), .B(n28355), .Z(n28354) );
  XOR U28263 ( .A(p_input[254]), .B(p_input[222]), .Z(n28355) );
  XNOR U28264 ( .A(n27984), .B(n28350), .Z(n28352) );
  XOR U28265 ( .A(n28356), .B(n28357), .Z(n27984) );
  AND U28266 ( .A(n628), .B(n28358), .Z(n28357) );
  XOR U28267 ( .A(p_input[190]), .B(p_input[158]), .Z(n28358) );
  XOR U28268 ( .A(n28359), .B(n28360), .Z(n28350) );
  AND U28269 ( .A(n28361), .B(n28362), .Z(n28360) );
  XOR U28270 ( .A(n28359), .B(n27999), .Z(n28362) );
  XNOR U28271 ( .A(p_input[221]), .B(n28363), .Z(n27999) );
  AND U28272 ( .A(n630), .B(n28364), .Z(n28363) );
  XOR U28273 ( .A(p_input[253]), .B(p_input[221]), .Z(n28364) );
  XNOR U28274 ( .A(n27996), .B(n28359), .Z(n28361) );
  XOR U28275 ( .A(n28365), .B(n28366), .Z(n27996) );
  AND U28276 ( .A(n628), .B(n28367), .Z(n28366) );
  XOR U28277 ( .A(p_input[189]), .B(p_input[157]), .Z(n28367) );
  XOR U28278 ( .A(n28368), .B(n28369), .Z(n28359) );
  AND U28279 ( .A(n28370), .B(n28371), .Z(n28369) );
  XOR U28280 ( .A(n28368), .B(n28011), .Z(n28371) );
  XNOR U28281 ( .A(p_input[220]), .B(n28372), .Z(n28011) );
  AND U28282 ( .A(n630), .B(n28373), .Z(n28372) );
  XOR U28283 ( .A(p_input[252]), .B(p_input[220]), .Z(n28373) );
  XNOR U28284 ( .A(n28008), .B(n28368), .Z(n28370) );
  XOR U28285 ( .A(n28374), .B(n28375), .Z(n28008) );
  AND U28286 ( .A(n628), .B(n28376), .Z(n28375) );
  XOR U28287 ( .A(p_input[188]), .B(p_input[156]), .Z(n28376) );
  XOR U28288 ( .A(n28377), .B(n28378), .Z(n28368) );
  AND U28289 ( .A(n28379), .B(n28380), .Z(n28378) );
  XOR U28290 ( .A(n28377), .B(n28023), .Z(n28380) );
  XNOR U28291 ( .A(p_input[219]), .B(n28381), .Z(n28023) );
  AND U28292 ( .A(n630), .B(n28382), .Z(n28381) );
  XOR U28293 ( .A(p_input[251]), .B(p_input[219]), .Z(n28382) );
  XNOR U28294 ( .A(n28020), .B(n28377), .Z(n28379) );
  XOR U28295 ( .A(n28383), .B(n28384), .Z(n28020) );
  AND U28296 ( .A(n628), .B(n28385), .Z(n28384) );
  XOR U28297 ( .A(p_input[187]), .B(p_input[155]), .Z(n28385) );
  XOR U28298 ( .A(n28386), .B(n28387), .Z(n28377) );
  AND U28299 ( .A(n28388), .B(n28389), .Z(n28387) );
  XOR U28300 ( .A(n28386), .B(n28035), .Z(n28389) );
  XNOR U28301 ( .A(p_input[218]), .B(n28390), .Z(n28035) );
  AND U28302 ( .A(n630), .B(n28391), .Z(n28390) );
  XOR U28303 ( .A(p_input[250]), .B(p_input[218]), .Z(n28391) );
  XNOR U28304 ( .A(n28032), .B(n28386), .Z(n28388) );
  XOR U28305 ( .A(n28392), .B(n28393), .Z(n28032) );
  AND U28306 ( .A(n628), .B(n28394), .Z(n28393) );
  XOR U28307 ( .A(p_input[186]), .B(p_input[154]), .Z(n28394) );
  XOR U28308 ( .A(n28395), .B(n28396), .Z(n28386) );
  AND U28309 ( .A(n28397), .B(n28398), .Z(n28396) );
  XOR U28310 ( .A(n28395), .B(n28047), .Z(n28398) );
  XNOR U28311 ( .A(p_input[217]), .B(n28399), .Z(n28047) );
  AND U28312 ( .A(n630), .B(n28400), .Z(n28399) );
  XOR U28313 ( .A(p_input[249]), .B(p_input[217]), .Z(n28400) );
  XNOR U28314 ( .A(n28044), .B(n28395), .Z(n28397) );
  XOR U28315 ( .A(n28401), .B(n28402), .Z(n28044) );
  AND U28316 ( .A(n628), .B(n28403), .Z(n28402) );
  XOR U28317 ( .A(p_input[185]), .B(p_input[153]), .Z(n28403) );
  XOR U28318 ( .A(n28404), .B(n28405), .Z(n28395) );
  AND U28319 ( .A(n28406), .B(n28407), .Z(n28405) );
  XOR U28320 ( .A(n28404), .B(n28059), .Z(n28407) );
  XNOR U28321 ( .A(p_input[216]), .B(n28408), .Z(n28059) );
  AND U28322 ( .A(n630), .B(n28409), .Z(n28408) );
  XOR U28323 ( .A(p_input[248]), .B(p_input[216]), .Z(n28409) );
  XNOR U28324 ( .A(n28056), .B(n28404), .Z(n28406) );
  XOR U28325 ( .A(n28410), .B(n28411), .Z(n28056) );
  AND U28326 ( .A(n628), .B(n28412), .Z(n28411) );
  XOR U28327 ( .A(p_input[184]), .B(p_input[152]), .Z(n28412) );
  XOR U28328 ( .A(n28413), .B(n28414), .Z(n28404) );
  AND U28329 ( .A(n28415), .B(n28416), .Z(n28414) );
  XOR U28330 ( .A(n28413), .B(n28071), .Z(n28416) );
  XNOR U28331 ( .A(p_input[215]), .B(n28417), .Z(n28071) );
  AND U28332 ( .A(n630), .B(n28418), .Z(n28417) );
  XOR U28333 ( .A(p_input[247]), .B(p_input[215]), .Z(n28418) );
  XNOR U28334 ( .A(n28068), .B(n28413), .Z(n28415) );
  XOR U28335 ( .A(n28419), .B(n28420), .Z(n28068) );
  AND U28336 ( .A(n628), .B(n28421), .Z(n28420) );
  XOR U28337 ( .A(p_input[183]), .B(p_input[151]), .Z(n28421) );
  XOR U28338 ( .A(n28422), .B(n28423), .Z(n28413) );
  AND U28339 ( .A(n28424), .B(n28425), .Z(n28423) );
  XOR U28340 ( .A(n28422), .B(n28083), .Z(n28425) );
  XNOR U28341 ( .A(p_input[214]), .B(n28426), .Z(n28083) );
  AND U28342 ( .A(n630), .B(n28427), .Z(n28426) );
  XOR U28343 ( .A(p_input[246]), .B(p_input[214]), .Z(n28427) );
  XNOR U28344 ( .A(n28080), .B(n28422), .Z(n28424) );
  XOR U28345 ( .A(n28428), .B(n28429), .Z(n28080) );
  AND U28346 ( .A(n628), .B(n28430), .Z(n28429) );
  XOR U28347 ( .A(p_input[182]), .B(p_input[150]), .Z(n28430) );
  XOR U28348 ( .A(n28431), .B(n28432), .Z(n28422) );
  AND U28349 ( .A(n28433), .B(n28434), .Z(n28432) );
  XOR U28350 ( .A(n28431), .B(n28095), .Z(n28434) );
  XNOR U28351 ( .A(p_input[213]), .B(n28435), .Z(n28095) );
  AND U28352 ( .A(n630), .B(n28436), .Z(n28435) );
  XOR U28353 ( .A(p_input[245]), .B(p_input[213]), .Z(n28436) );
  XNOR U28354 ( .A(n28092), .B(n28431), .Z(n28433) );
  XOR U28355 ( .A(n28437), .B(n28438), .Z(n28092) );
  AND U28356 ( .A(n628), .B(n28439), .Z(n28438) );
  XOR U28357 ( .A(p_input[181]), .B(p_input[149]), .Z(n28439) );
  XOR U28358 ( .A(n28440), .B(n28441), .Z(n28431) );
  AND U28359 ( .A(n28442), .B(n28443), .Z(n28441) );
  XOR U28360 ( .A(n28440), .B(n28107), .Z(n28443) );
  XNOR U28361 ( .A(p_input[212]), .B(n28444), .Z(n28107) );
  AND U28362 ( .A(n630), .B(n28445), .Z(n28444) );
  XOR U28363 ( .A(p_input[244]), .B(p_input[212]), .Z(n28445) );
  XNOR U28364 ( .A(n28104), .B(n28440), .Z(n28442) );
  XOR U28365 ( .A(n28446), .B(n28447), .Z(n28104) );
  AND U28366 ( .A(n628), .B(n28448), .Z(n28447) );
  XOR U28367 ( .A(p_input[180]), .B(p_input[148]), .Z(n28448) );
  XOR U28368 ( .A(n28449), .B(n28450), .Z(n28440) );
  AND U28369 ( .A(n28451), .B(n28452), .Z(n28450) );
  XOR U28370 ( .A(n28449), .B(n28119), .Z(n28452) );
  XNOR U28371 ( .A(p_input[211]), .B(n28453), .Z(n28119) );
  AND U28372 ( .A(n630), .B(n28454), .Z(n28453) );
  XOR U28373 ( .A(p_input[243]), .B(p_input[211]), .Z(n28454) );
  XNOR U28374 ( .A(n28116), .B(n28449), .Z(n28451) );
  XOR U28375 ( .A(n28455), .B(n28456), .Z(n28116) );
  AND U28376 ( .A(n628), .B(n28457), .Z(n28456) );
  XOR U28377 ( .A(p_input[179]), .B(p_input[147]), .Z(n28457) );
  XOR U28378 ( .A(n28458), .B(n28459), .Z(n28449) );
  AND U28379 ( .A(n28460), .B(n28461), .Z(n28459) );
  XOR U28380 ( .A(n28458), .B(n28131), .Z(n28461) );
  XNOR U28381 ( .A(p_input[210]), .B(n28462), .Z(n28131) );
  AND U28382 ( .A(n630), .B(n28463), .Z(n28462) );
  XOR U28383 ( .A(p_input[242]), .B(p_input[210]), .Z(n28463) );
  XNOR U28384 ( .A(n28128), .B(n28458), .Z(n28460) );
  XOR U28385 ( .A(n28464), .B(n28465), .Z(n28128) );
  AND U28386 ( .A(n628), .B(n28466), .Z(n28465) );
  XOR U28387 ( .A(p_input[178]), .B(p_input[146]), .Z(n28466) );
  XOR U28388 ( .A(n28467), .B(n28468), .Z(n28458) );
  AND U28389 ( .A(n28469), .B(n28470), .Z(n28468) );
  XOR U28390 ( .A(n28467), .B(n28143), .Z(n28470) );
  XNOR U28391 ( .A(p_input[209]), .B(n28471), .Z(n28143) );
  AND U28392 ( .A(n630), .B(n28472), .Z(n28471) );
  XOR U28393 ( .A(p_input[241]), .B(p_input[209]), .Z(n28472) );
  XNOR U28394 ( .A(n28140), .B(n28467), .Z(n28469) );
  XOR U28395 ( .A(n28473), .B(n28474), .Z(n28140) );
  AND U28396 ( .A(n628), .B(n28475), .Z(n28474) );
  XOR U28397 ( .A(p_input[177]), .B(p_input[145]), .Z(n28475) );
  XOR U28398 ( .A(n28476), .B(n28477), .Z(n28467) );
  AND U28399 ( .A(n28478), .B(n28479), .Z(n28477) );
  XOR U28400 ( .A(n28476), .B(n28155), .Z(n28479) );
  XNOR U28401 ( .A(p_input[208]), .B(n28480), .Z(n28155) );
  AND U28402 ( .A(n630), .B(n28481), .Z(n28480) );
  XOR U28403 ( .A(p_input[240]), .B(p_input[208]), .Z(n28481) );
  XNOR U28404 ( .A(n28152), .B(n28476), .Z(n28478) );
  XOR U28405 ( .A(n28482), .B(n28483), .Z(n28152) );
  AND U28406 ( .A(n628), .B(n28484), .Z(n28483) );
  XOR U28407 ( .A(p_input[176]), .B(p_input[144]), .Z(n28484) );
  XOR U28408 ( .A(n28485), .B(n28486), .Z(n28476) );
  AND U28409 ( .A(n28487), .B(n28488), .Z(n28486) );
  XOR U28410 ( .A(n28485), .B(n28167), .Z(n28488) );
  XNOR U28411 ( .A(p_input[207]), .B(n28489), .Z(n28167) );
  AND U28412 ( .A(n630), .B(n28490), .Z(n28489) );
  XOR U28413 ( .A(p_input[239]), .B(p_input[207]), .Z(n28490) );
  XNOR U28414 ( .A(n28164), .B(n28485), .Z(n28487) );
  XOR U28415 ( .A(n28491), .B(n28492), .Z(n28164) );
  AND U28416 ( .A(n628), .B(n28493), .Z(n28492) );
  XOR U28417 ( .A(p_input[175]), .B(p_input[143]), .Z(n28493) );
  XOR U28418 ( .A(n28494), .B(n28495), .Z(n28485) );
  AND U28419 ( .A(n28496), .B(n28497), .Z(n28495) );
  XOR U28420 ( .A(n28494), .B(n28179), .Z(n28497) );
  XNOR U28421 ( .A(p_input[206]), .B(n28498), .Z(n28179) );
  AND U28422 ( .A(n630), .B(n28499), .Z(n28498) );
  XOR U28423 ( .A(p_input[238]), .B(p_input[206]), .Z(n28499) );
  XNOR U28424 ( .A(n28176), .B(n28494), .Z(n28496) );
  XOR U28425 ( .A(n28500), .B(n28501), .Z(n28176) );
  AND U28426 ( .A(n628), .B(n28502), .Z(n28501) );
  XOR U28427 ( .A(p_input[174]), .B(p_input[142]), .Z(n28502) );
  XOR U28428 ( .A(n28503), .B(n28504), .Z(n28494) );
  AND U28429 ( .A(n28505), .B(n28506), .Z(n28504) );
  XOR U28430 ( .A(n28503), .B(n28191), .Z(n28506) );
  XNOR U28431 ( .A(p_input[205]), .B(n28507), .Z(n28191) );
  AND U28432 ( .A(n630), .B(n28508), .Z(n28507) );
  XOR U28433 ( .A(p_input[237]), .B(p_input[205]), .Z(n28508) );
  XNOR U28434 ( .A(n28188), .B(n28503), .Z(n28505) );
  XOR U28435 ( .A(n28509), .B(n28510), .Z(n28188) );
  AND U28436 ( .A(n628), .B(n28511), .Z(n28510) );
  XOR U28437 ( .A(p_input[173]), .B(p_input[141]), .Z(n28511) );
  XOR U28438 ( .A(n28512), .B(n28513), .Z(n28503) );
  AND U28439 ( .A(n28514), .B(n28515), .Z(n28513) );
  XOR U28440 ( .A(n28512), .B(n28203), .Z(n28515) );
  XNOR U28441 ( .A(p_input[204]), .B(n28516), .Z(n28203) );
  AND U28442 ( .A(n630), .B(n28517), .Z(n28516) );
  XOR U28443 ( .A(p_input[236]), .B(p_input[204]), .Z(n28517) );
  XNOR U28444 ( .A(n28200), .B(n28512), .Z(n28514) );
  XOR U28445 ( .A(n28518), .B(n28519), .Z(n28200) );
  AND U28446 ( .A(n628), .B(n28520), .Z(n28519) );
  XOR U28447 ( .A(p_input[172]), .B(p_input[140]), .Z(n28520) );
  XOR U28448 ( .A(n28521), .B(n28522), .Z(n28512) );
  AND U28449 ( .A(n28523), .B(n28524), .Z(n28522) );
  XOR U28450 ( .A(n28521), .B(n28215), .Z(n28524) );
  XNOR U28451 ( .A(p_input[203]), .B(n28525), .Z(n28215) );
  AND U28452 ( .A(n630), .B(n28526), .Z(n28525) );
  XOR U28453 ( .A(p_input[235]), .B(p_input[203]), .Z(n28526) );
  XNOR U28454 ( .A(n28212), .B(n28521), .Z(n28523) );
  XOR U28455 ( .A(n28527), .B(n28528), .Z(n28212) );
  AND U28456 ( .A(n628), .B(n28529), .Z(n28528) );
  XOR U28457 ( .A(p_input[171]), .B(p_input[139]), .Z(n28529) );
  XOR U28458 ( .A(n28530), .B(n28531), .Z(n28521) );
  AND U28459 ( .A(n28532), .B(n28533), .Z(n28531) );
  XOR U28460 ( .A(n28530), .B(n28227), .Z(n28533) );
  XNOR U28461 ( .A(p_input[202]), .B(n28534), .Z(n28227) );
  AND U28462 ( .A(n630), .B(n28535), .Z(n28534) );
  XOR U28463 ( .A(p_input[234]), .B(p_input[202]), .Z(n28535) );
  XNOR U28464 ( .A(n28224), .B(n28530), .Z(n28532) );
  XOR U28465 ( .A(n28536), .B(n28537), .Z(n28224) );
  AND U28466 ( .A(n628), .B(n28538), .Z(n28537) );
  XOR U28467 ( .A(p_input[170]), .B(p_input[138]), .Z(n28538) );
  XOR U28468 ( .A(n28539), .B(n28540), .Z(n28530) );
  AND U28469 ( .A(n28541), .B(n28542), .Z(n28540) );
  XOR U28470 ( .A(n28539), .B(n28239), .Z(n28542) );
  XNOR U28471 ( .A(p_input[201]), .B(n28543), .Z(n28239) );
  AND U28472 ( .A(n630), .B(n28544), .Z(n28543) );
  XOR U28473 ( .A(p_input[233]), .B(p_input[201]), .Z(n28544) );
  XNOR U28474 ( .A(n28236), .B(n28539), .Z(n28541) );
  XOR U28475 ( .A(n28545), .B(n28546), .Z(n28236) );
  AND U28476 ( .A(n628), .B(n28547), .Z(n28546) );
  XOR U28477 ( .A(p_input[169]), .B(p_input[137]), .Z(n28547) );
  XOR U28478 ( .A(n28548), .B(n28549), .Z(n28539) );
  AND U28479 ( .A(n28550), .B(n28551), .Z(n28549) );
  XOR U28480 ( .A(n28548), .B(n28251), .Z(n28551) );
  XNOR U28481 ( .A(p_input[200]), .B(n28552), .Z(n28251) );
  AND U28482 ( .A(n630), .B(n28553), .Z(n28552) );
  XOR U28483 ( .A(p_input[232]), .B(p_input[200]), .Z(n28553) );
  XNOR U28484 ( .A(n28248), .B(n28548), .Z(n28550) );
  XOR U28485 ( .A(n28554), .B(n28555), .Z(n28248) );
  AND U28486 ( .A(n628), .B(n28556), .Z(n28555) );
  XOR U28487 ( .A(p_input[168]), .B(p_input[136]), .Z(n28556) );
  XOR U28488 ( .A(n28557), .B(n28558), .Z(n28548) );
  AND U28489 ( .A(n28559), .B(n28560), .Z(n28558) );
  XOR U28490 ( .A(n28557), .B(n28263), .Z(n28560) );
  XNOR U28491 ( .A(p_input[199]), .B(n28561), .Z(n28263) );
  AND U28492 ( .A(n630), .B(n28562), .Z(n28561) );
  XOR U28493 ( .A(p_input[231]), .B(p_input[199]), .Z(n28562) );
  XNOR U28494 ( .A(n28260), .B(n28557), .Z(n28559) );
  XOR U28495 ( .A(n28563), .B(n28564), .Z(n28260) );
  AND U28496 ( .A(n628), .B(n28565), .Z(n28564) );
  XOR U28497 ( .A(p_input[167]), .B(p_input[135]), .Z(n28565) );
  XOR U28498 ( .A(n28566), .B(n28567), .Z(n28557) );
  AND U28499 ( .A(n28568), .B(n28569), .Z(n28567) );
  XOR U28500 ( .A(n28566), .B(n28275), .Z(n28569) );
  XNOR U28501 ( .A(p_input[198]), .B(n28570), .Z(n28275) );
  AND U28502 ( .A(n630), .B(n28571), .Z(n28570) );
  XOR U28503 ( .A(p_input[230]), .B(p_input[198]), .Z(n28571) );
  XNOR U28504 ( .A(n28272), .B(n28566), .Z(n28568) );
  XOR U28505 ( .A(n28572), .B(n28573), .Z(n28272) );
  AND U28506 ( .A(n628), .B(n28574), .Z(n28573) );
  XOR U28507 ( .A(p_input[166]), .B(p_input[134]), .Z(n28574) );
  XOR U28508 ( .A(n28575), .B(n28576), .Z(n28566) );
  AND U28509 ( .A(n28577), .B(n28578), .Z(n28576) );
  XOR U28510 ( .A(n28575), .B(n28287), .Z(n28578) );
  XNOR U28511 ( .A(p_input[197]), .B(n28579), .Z(n28287) );
  AND U28512 ( .A(n630), .B(n28580), .Z(n28579) );
  XOR U28513 ( .A(p_input[229]), .B(p_input[197]), .Z(n28580) );
  XNOR U28514 ( .A(n28284), .B(n28575), .Z(n28577) );
  XOR U28515 ( .A(n28581), .B(n28582), .Z(n28284) );
  AND U28516 ( .A(n628), .B(n28583), .Z(n28582) );
  XOR U28517 ( .A(p_input[165]), .B(p_input[133]), .Z(n28583) );
  XOR U28518 ( .A(n28584), .B(n28585), .Z(n28575) );
  AND U28519 ( .A(n28586), .B(n28587), .Z(n28585) );
  XOR U28520 ( .A(n28584), .B(n28299), .Z(n28587) );
  XNOR U28521 ( .A(p_input[196]), .B(n28588), .Z(n28299) );
  AND U28522 ( .A(n630), .B(n28589), .Z(n28588) );
  XOR U28523 ( .A(p_input[228]), .B(p_input[196]), .Z(n28589) );
  XNOR U28524 ( .A(n28296), .B(n28584), .Z(n28586) );
  XOR U28525 ( .A(n28590), .B(n28591), .Z(n28296) );
  AND U28526 ( .A(n628), .B(n28592), .Z(n28591) );
  XOR U28527 ( .A(p_input[164]), .B(p_input[132]), .Z(n28592) );
  XOR U28528 ( .A(n28593), .B(n28594), .Z(n28584) );
  AND U28529 ( .A(n28595), .B(n28596), .Z(n28594) );
  XOR U28530 ( .A(n28593), .B(n28311), .Z(n28596) );
  XNOR U28531 ( .A(p_input[195]), .B(n28597), .Z(n28311) );
  AND U28532 ( .A(n630), .B(n28598), .Z(n28597) );
  XOR U28533 ( .A(p_input[227]), .B(p_input[195]), .Z(n28598) );
  XNOR U28534 ( .A(n28308), .B(n28593), .Z(n28595) );
  XOR U28535 ( .A(n28599), .B(n28600), .Z(n28308) );
  AND U28536 ( .A(n628), .B(n28601), .Z(n28600) );
  XOR U28537 ( .A(p_input[163]), .B(p_input[131]), .Z(n28601) );
  XOR U28538 ( .A(n28602), .B(n28603), .Z(n28593) );
  AND U28539 ( .A(n28604), .B(n28605), .Z(n28603) );
  XOR U28540 ( .A(n28323), .B(n28602), .Z(n28605) );
  XNOR U28541 ( .A(p_input[194]), .B(n28606), .Z(n28323) );
  AND U28542 ( .A(n630), .B(n28607), .Z(n28606) );
  XOR U28543 ( .A(p_input[226]), .B(p_input[194]), .Z(n28607) );
  XNOR U28544 ( .A(n28602), .B(n28320), .Z(n28604) );
  XOR U28545 ( .A(n28608), .B(n28609), .Z(n28320) );
  AND U28546 ( .A(n628), .B(n28610), .Z(n28609) );
  XOR U28547 ( .A(p_input[162]), .B(p_input[130]), .Z(n28610) );
  XOR U28548 ( .A(n28611), .B(n28612), .Z(n28602) );
  AND U28549 ( .A(n28613), .B(n28614), .Z(n28612) );
  XNOR U28550 ( .A(n28615), .B(n28336), .Z(n28614) );
  XNOR U28551 ( .A(p_input[193]), .B(n28616), .Z(n28336) );
  AND U28552 ( .A(n630), .B(n28617), .Z(n28616) );
  XNOR U28553 ( .A(p_input[225]), .B(n28618), .Z(n28617) );
  IV U28554 ( .A(p_input[193]), .Z(n28618) );
  XNOR U28555 ( .A(n28333), .B(n28611), .Z(n28613) );
  XNOR U28556 ( .A(p_input[129]), .B(n28619), .Z(n28333) );
  AND U28557 ( .A(n628), .B(n28620), .Z(n28619) );
  XOR U28558 ( .A(p_input[161]), .B(p_input[129]), .Z(n28620) );
  IV U28559 ( .A(n28615), .Z(n28611) );
  AND U28560 ( .A(n28341), .B(n28344), .Z(n28615) );
  XOR U28561 ( .A(p_input[192]), .B(n28621), .Z(n28344) );
  AND U28562 ( .A(n630), .B(n28622), .Z(n28621) );
  XOR U28563 ( .A(p_input[224]), .B(p_input[192]), .Z(n28622) );
  XOR U28564 ( .A(n28623), .B(n28624), .Z(n630) );
  AND U28565 ( .A(n28625), .B(n28626), .Z(n28624) );
  XNOR U28566 ( .A(p_input[255]), .B(n28623), .Z(n28626) );
  XOR U28567 ( .A(n28623), .B(p_input[223]), .Z(n28625) );
  XOR U28568 ( .A(n28627), .B(n28628), .Z(n28623) );
  AND U28569 ( .A(n28629), .B(n28630), .Z(n28628) );
  XNOR U28570 ( .A(p_input[254]), .B(n28627), .Z(n28630) );
  XOR U28571 ( .A(n28627), .B(p_input[222]), .Z(n28629) );
  XOR U28572 ( .A(n28631), .B(n28632), .Z(n28627) );
  AND U28573 ( .A(n28633), .B(n28634), .Z(n28632) );
  XNOR U28574 ( .A(p_input[253]), .B(n28631), .Z(n28634) );
  XOR U28575 ( .A(n28631), .B(p_input[221]), .Z(n28633) );
  XOR U28576 ( .A(n28635), .B(n28636), .Z(n28631) );
  AND U28577 ( .A(n28637), .B(n28638), .Z(n28636) );
  XNOR U28578 ( .A(p_input[252]), .B(n28635), .Z(n28638) );
  XOR U28579 ( .A(n28635), .B(p_input[220]), .Z(n28637) );
  XOR U28580 ( .A(n28639), .B(n28640), .Z(n28635) );
  AND U28581 ( .A(n28641), .B(n28642), .Z(n28640) );
  XNOR U28582 ( .A(p_input[251]), .B(n28639), .Z(n28642) );
  XOR U28583 ( .A(n28639), .B(p_input[219]), .Z(n28641) );
  XOR U28584 ( .A(n28643), .B(n28644), .Z(n28639) );
  AND U28585 ( .A(n28645), .B(n28646), .Z(n28644) );
  XNOR U28586 ( .A(p_input[250]), .B(n28643), .Z(n28646) );
  XOR U28587 ( .A(n28643), .B(p_input[218]), .Z(n28645) );
  XOR U28588 ( .A(n28647), .B(n28648), .Z(n28643) );
  AND U28589 ( .A(n28649), .B(n28650), .Z(n28648) );
  XNOR U28590 ( .A(p_input[249]), .B(n28647), .Z(n28650) );
  XOR U28591 ( .A(n28647), .B(p_input[217]), .Z(n28649) );
  XOR U28592 ( .A(n28651), .B(n28652), .Z(n28647) );
  AND U28593 ( .A(n28653), .B(n28654), .Z(n28652) );
  XNOR U28594 ( .A(p_input[248]), .B(n28651), .Z(n28654) );
  XOR U28595 ( .A(n28651), .B(p_input[216]), .Z(n28653) );
  XOR U28596 ( .A(n28655), .B(n28656), .Z(n28651) );
  AND U28597 ( .A(n28657), .B(n28658), .Z(n28656) );
  XNOR U28598 ( .A(p_input[247]), .B(n28655), .Z(n28658) );
  XOR U28599 ( .A(n28655), .B(p_input[215]), .Z(n28657) );
  XOR U28600 ( .A(n28659), .B(n28660), .Z(n28655) );
  AND U28601 ( .A(n28661), .B(n28662), .Z(n28660) );
  XNOR U28602 ( .A(p_input[246]), .B(n28659), .Z(n28662) );
  XOR U28603 ( .A(n28659), .B(p_input[214]), .Z(n28661) );
  XOR U28604 ( .A(n28663), .B(n28664), .Z(n28659) );
  AND U28605 ( .A(n28665), .B(n28666), .Z(n28664) );
  XNOR U28606 ( .A(p_input[245]), .B(n28663), .Z(n28666) );
  XOR U28607 ( .A(n28663), .B(p_input[213]), .Z(n28665) );
  XOR U28608 ( .A(n28667), .B(n28668), .Z(n28663) );
  AND U28609 ( .A(n28669), .B(n28670), .Z(n28668) );
  XNOR U28610 ( .A(p_input[244]), .B(n28667), .Z(n28670) );
  XOR U28611 ( .A(n28667), .B(p_input[212]), .Z(n28669) );
  XOR U28612 ( .A(n28671), .B(n28672), .Z(n28667) );
  AND U28613 ( .A(n28673), .B(n28674), .Z(n28672) );
  XNOR U28614 ( .A(p_input[243]), .B(n28671), .Z(n28674) );
  XOR U28615 ( .A(n28671), .B(p_input[211]), .Z(n28673) );
  XOR U28616 ( .A(n28675), .B(n28676), .Z(n28671) );
  AND U28617 ( .A(n28677), .B(n28678), .Z(n28676) );
  XNOR U28618 ( .A(p_input[242]), .B(n28675), .Z(n28678) );
  XOR U28619 ( .A(n28675), .B(p_input[210]), .Z(n28677) );
  XOR U28620 ( .A(n28679), .B(n28680), .Z(n28675) );
  AND U28621 ( .A(n28681), .B(n28682), .Z(n28680) );
  XNOR U28622 ( .A(p_input[241]), .B(n28679), .Z(n28682) );
  XOR U28623 ( .A(n28679), .B(p_input[209]), .Z(n28681) );
  XOR U28624 ( .A(n28683), .B(n28684), .Z(n28679) );
  AND U28625 ( .A(n28685), .B(n28686), .Z(n28684) );
  XNOR U28626 ( .A(p_input[240]), .B(n28683), .Z(n28686) );
  XOR U28627 ( .A(n28683), .B(p_input[208]), .Z(n28685) );
  XOR U28628 ( .A(n28687), .B(n28688), .Z(n28683) );
  AND U28629 ( .A(n28689), .B(n28690), .Z(n28688) );
  XNOR U28630 ( .A(p_input[239]), .B(n28687), .Z(n28690) );
  XOR U28631 ( .A(n28687), .B(p_input[207]), .Z(n28689) );
  XOR U28632 ( .A(n28691), .B(n28692), .Z(n28687) );
  AND U28633 ( .A(n28693), .B(n28694), .Z(n28692) );
  XNOR U28634 ( .A(p_input[238]), .B(n28691), .Z(n28694) );
  XOR U28635 ( .A(n28691), .B(p_input[206]), .Z(n28693) );
  XOR U28636 ( .A(n28695), .B(n28696), .Z(n28691) );
  AND U28637 ( .A(n28697), .B(n28698), .Z(n28696) );
  XNOR U28638 ( .A(p_input[237]), .B(n28695), .Z(n28698) );
  XOR U28639 ( .A(n28695), .B(p_input[205]), .Z(n28697) );
  XOR U28640 ( .A(n28699), .B(n28700), .Z(n28695) );
  AND U28641 ( .A(n28701), .B(n28702), .Z(n28700) );
  XNOR U28642 ( .A(p_input[236]), .B(n28699), .Z(n28702) );
  XOR U28643 ( .A(n28699), .B(p_input[204]), .Z(n28701) );
  XOR U28644 ( .A(n28703), .B(n28704), .Z(n28699) );
  AND U28645 ( .A(n28705), .B(n28706), .Z(n28704) );
  XNOR U28646 ( .A(p_input[235]), .B(n28703), .Z(n28706) );
  XOR U28647 ( .A(n28703), .B(p_input[203]), .Z(n28705) );
  XOR U28648 ( .A(n28707), .B(n28708), .Z(n28703) );
  AND U28649 ( .A(n28709), .B(n28710), .Z(n28708) );
  XNOR U28650 ( .A(p_input[234]), .B(n28707), .Z(n28710) );
  XOR U28651 ( .A(n28707), .B(p_input[202]), .Z(n28709) );
  XOR U28652 ( .A(n28711), .B(n28712), .Z(n28707) );
  AND U28653 ( .A(n28713), .B(n28714), .Z(n28712) );
  XNOR U28654 ( .A(p_input[233]), .B(n28711), .Z(n28714) );
  XOR U28655 ( .A(n28711), .B(p_input[201]), .Z(n28713) );
  XOR U28656 ( .A(n28715), .B(n28716), .Z(n28711) );
  AND U28657 ( .A(n28717), .B(n28718), .Z(n28716) );
  XNOR U28658 ( .A(p_input[232]), .B(n28715), .Z(n28718) );
  XOR U28659 ( .A(n28715), .B(p_input[200]), .Z(n28717) );
  XOR U28660 ( .A(n28719), .B(n28720), .Z(n28715) );
  AND U28661 ( .A(n28721), .B(n28722), .Z(n28720) );
  XNOR U28662 ( .A(p_input[231]), .B(n28719), .Z(n28722) );
  XOR U28663 ( .A(n28719), .B(p_input[199]), .Z(n28721) );
  XOR U28664 ( .A(n28723), .B(n28724), .Z(n28719) );
  AND U28665 ( .A(n28725), .B(n28726), .Z(n28724) );
  XNOR U28666 ( .A(p_input[230]), .B(n28723), .Z(n28726) );
  XOR U28667 ( .A(n28723), .B(p_input[198]), .Z(n28725) );
  XOR U28668 ( .A(n28727), .B(n28728), .Z(n28723) );
  AND U28669 ( .A(n28729), .B(n28730), .Z(n28728) );
  XNOR U28670 ( .A(p_input[229]), .B(n28727), .Z(n28730) );
  XOR U28671 ( .A(n28727), .B(p_input[197]), .Z(n28729) );
  XOR U28672 ( .A(n28731), .B(n28732), .Z(n28727) );
  AND U28673 ( .A(n28733), .B(n28734), .Z(n28732) );
  XNOR U28674 ( .A(p_input[228]), .B(n28731), .Z(n28734) );
  XOR U28675 ( .A(n28731), .B(p_input[196]), .Z(n28733) );
  XOR U28676 ( .A(n28735), .B(n28736), .Z(n28731) );
  AND U28677 ( .A(n28737), .B(n28738), .Z(n28736) );
  XNOR U28678 ( .A(p_input[227]), .B(n28735), .Z(n28738) );
  XOR U28679 ( .A(n28735), .B(p_input[195]), .Z(n28737) );
  XOR U28680 ( .A(n28739), .B(n28740), .Z(n28735) );
  AND U28681 ( .A(n28741), .B(n28742), .Z(n28740) );
  XNOR U28682 ( .A(p_input[226]), .B(n28739), .Z(n28742) );
  XOR U28683 ( .A(n28739), .B(p_input[194]), .Z(n28741) );
  XNOR U28684 ( .A(n28743), .B(n28744), .Z(n28739) );
  AND U28685 ( .A(n28745), .B(n28746), .Z(n28744) );
  XOR U28686 ( .A(p_input[225]), .B(n28743), .Z(n28746) );
  XNOR U28687 ( .A(p_input[193]), .B(n28743), .Z(n28745) );
  AND U28688 ( .A(p_input[224]), .B(n28747), .Z(n28743) );
  IV U28689 ( .A(p_input[192]), .Z(n28747) );
  XNOR U28690 ( .A(p_input[128]), .B(n28748), .Z(n28341) );
  AND U28691 ( .A(n628), .B(n28749), .Z(n28748) );
  XOR U28692 ( .A(p_input[160]), .B(p_input[128]), .Z(n28749) );
  XOR U28693 ( .A(n28750), .B(n28751), .Z(n628) );
  AND U28694 ( .A(n28752), .B(n28753), .Z(n28751) );
  XNOR U28695 ( .A(p_input[191]), .B(n28750), .Z(n28753) );
  XOR U28696 ( .A(n28750), .B(p_input[159]), .Z(n28752) );
  XOR U28697 ( .A(n28754), .B(n28755), .Z(n28750) );
  AND U28698 ( .A(n28756), .B(n28757), .Z(n28755) );
  XNOR U28699 ( .A(p_input[190]), .B(n28754), .Z(n28757) );
  XNOR U28700 ( .A(n28754), .B(n28356), .Z(n28756) );
  IV U28701 ( .A(p_input[158]), .Z(n28356) );
  XOR U28702 ( .A(n28758), .B(n28759), .Z(n28754) );
  AND U28703 ( .A(n28760), .B(n28761), .Z(n28759) );
  XNOR U28704 ( .A(p_input[189]), .B(n28758), .Z(n28761) );
  XNOR U28705 ( .A(n28758), .B(n28365), .Z(n28760) );
  IV U28706 ( .A(p_input[157]), .Z(n28365) );
  XOR U28707 ( .A(n28762), .B(n28763), .Z(n28758) );
  AND U28708 ( .A(n28764), .B(n28765), .Z(n28763) );
  XNOR U28709 ( .A(p_input[188]), .B(n28762), .Z(n28765) );
  XNOR U28710 ( .A(n28762), .B(n28374), .Z(n28764) );
  IV U28711 ( .A(p_input[156]), .Z(n28374) );
  XOR U28712 ( .A(n28766), .B(n28767), .Z(n28762) );
  AND U28713 ( .A(n28768), .B(n28769), .Z(n28767) );
  XNOR U28714 ( .A(p_input[187]), .B(n28766), .Z(n28769) );
  XNOR U28715 ( .A(n28766), .B(n28383), .Z(n28768) );
  IV U28716 ( .A(p_input[155]), .Z(n28383) );
  XOR U28717 ( .A(n28770), .B(n28771), .Z(n28766) );
  AND U28718 ( .A(n28772), .B(n28773), .Z(n28771) );
  XNOR U28719 ( .A(p_input[186]), .B(n28770), .Z(n28773) );
  XNOR U28720 ( .A(n28770), .B(n28392), .Z(n28772) );
  IV U28721 ( .A(p_input[154]), .Z(n28392) );
  XOR U28722 ( .A(n28774), .B(n28775), .Z(n28770) );
  AND U28723 ( .A(n28776), .B(n28777), .Z(n28775) );
  XNOR U28724 ( .A(p_input[185]), .B(n28774), .Z(n28777) );
  XNOR U28725 ( .A(n28774), .B(n28401), .Z(n28776) );
  IV U28726 ( .A(p_input[153]), .Z(n28401) );
  XOR U28727 ( .A(n28778), .B(n28779), .Z(n28774) );
  AND U28728 ( .A(n28780), .B(n28781), .Z(n28779) );
  XNOR U28729 ( .A(p_input[184]), .B(n28778), .Z(n28781) );
  XNOR U28730 ( .A(n28778), .B(n28410), .Z(n28780) );
  IV U28731 ( .A(p_input[152]), .Z(n28410) );
  XOR U28732 ( .A(n28782), .B(n28783), .Z(n28778) );
  AND U28733 ( .A(n28784), .B(n28785), .Z(n28783) );
  XNOR U28734 ( .A(p_input[183]), .B(n28782), .Z(n28785) );
  XNOR U28735 ( .A(n28782), .B(n28419), .Z(n28784) );
  IV U28736 ( .A(p_input[151]), .Z(n28419) );
  XOR U28737 ( .A(n28786), .B(n28787), .Z(n28782) );
  AND U28738 ( .A(n28788), .B(n28789), .Z(n28787) );
  XNOR U28739 ( .A(p_input[182]), .B(n28786), .Z(n28789) );
  XNOR U28740 ( .A(n28786), .B(n28428), .Z(n28788) );
  IV U28741 ( .A(p_input[150]), .Z(n28428) );
  XOR U28742 ( .A(n28790), .B(n28791), .Z(n28786) );
  AND U28743 ( .A(n28792), .B(n28793), .Z(n28791) );
  XNOR U28744 ( .A(p_input[181]), .B(n28790), .Z(n28793) );
  XNOR U28745 ( .A(n28790), .B(n28437), .Z(n28792) );
  IV U28746 ( .A(p_input[149]), .Z(n28437) );
  XOR U28747 ( .A(n28794), .B(n28795), .Z(n28790) );
  AND U28748 ( .A(n28796), .B(n28797), .Z(n28795) );
  XNOR U28749 ( .A(p_input[180]), .B(n28794), .Z(n28797) );
  XNOR U28750 ( .A(n28794), .B(n28446), .Z(n28796) );
  IV U28751 ( .A(p_input[148]), .Z(n28446) );
  XOR U28752 ( .A(n28798), .B(n28799), .Z(n28794) );
  AND U28753 ( .A(n28800), .B(n28801), .Z(n28799) );
  XNOR U28754 ( .A(p_input[179]), .B(n28798), .Z(n28801) );
  XNOR U28755 ( .A(n28798), .B(n28455), .Z(n28800) );
  IV U28756 ( .A(p_input[147]), .Z(n28455) );
  XOR U28757 ( .A(n28802), .B(n28803), .Z(n28798) );
  AND U28758 ( .A(n28804), .B(n28805), .Z(n28803) );
  XNOR U28759 ( .A(p_input[178]), .B(n28802), .Z(n28805) );
  XNOR U28760 ( .A(n28802), .B(n28464), .Z(n28804) );
  IV U28761 ( .A(p_input[146]), .Z(n28464) );
  XOR U28762 ( .A(n28806), .B(n28807), .Z(n28802) );
  AND U28763 ( .A(n28808), .B(n28809), .Z(n28807) );
  XNOR U28764 ( .A(p_input[177]), .B(n28806), .Z(n28809) );
  XNOR U28765 ( .A(n28806), .B(n28473), .Z(n28808) );
  IV U28766 ( .A(p_input[145]), .Z(n28473) );
  XOR U28767 ( .A(n28810), .B(n28811), .Z(n28806) );
  AND U28768 ( .A(n28812), .B(n28813), .Z(n28811) );
  XNOR U28769 ( .A(p_input[176]), .B(n28810), .Z(n28813) );
  XNOR U28770 ( .A(n28810), .B(n28482), .Z(n28812) );
  IV U28771 ( .A(p_input[144]), .Z(n28482) );
  XOR U28772 ( .A(n28814), .B(n28815), .Z(n28810) );
  AND U28773 ( .A(n28816), .B(n28817), .Z(n28815) );
  XNOR U28774 ( .A(p_input[175]), .B(n28814), .Z(n28817) );
  XNOR U28775 ( .A(n28814), .B(n28491), .Z(n28816) );
  IV U28776 ( .A(p_input[143]), .Z(n28491) );
  XOR U28777 ( .A(n28818), .B(n28819), .Z(n28814) );
  AND U28778 ( .A(n28820), .B(n28821), .Z(n28819) );
  XNOR U28779 ( .A(p_input[174]), .B(n28818), .Z(n28821) );
  XNOR U28780 ( .A(n28818), .B(n28500), .Z(n28820) );
  IV U28781 ( .A(p_input[142]), .Z(n28500) );
  XOR U28782 ( .A(n28822), .B(n28823), .Z(n28818) );
  AND U28783 ( .A(n28824), .B(n28825), .Z(n28823) );
  XNOR U28784 ( .A(p_input[173]), .B(n28822), .Z(n28825) );
  XNOR U28785 ( .A(n28822), .B(n28509), .Z(n28824) );
  IV U28786 ( .A(p_input[141]), .Z(n28509) );
  XOR U28787 ( .A(n28826), .B(n28827), .Z(n28822) );
  AND U28788 ( .A(n28828), .B(n28829), .Z(n28827) );
  XNOR U28789 ( .A(p_input[172]), .B(n28826), .Z(n28829) );
  XNOR U28790 ( .A(n28826), .B(n28518), .Z(n28828) );
  IV U28791 ( .A(p_input[140]), .Z(n28518) );
  XOR U28792 ( .A(n28830), .B(n28831), .Z(n28826) );
  AND U28793 ( .A(n28832), .B(n28833), .Z(n28831) );
  XNOR U28794 ( .A(p_input[171]), .B(n28830), .Z(n28833) );
  XNOR U28795 ( .A(n28830), .B(n28527), .Z(n28832) );
  IV U28796 ( .A(p_input[139]), .Z(n28527) );
  XOR U28797 ( .A(n28834), .B(n28835), .Z(n28830) );
  AND U28798 ( .A(n28836), .B(n28837), .Z(n28835) );
  XNOR U28799 ( .A(p_input[170]), .B(n28834), .Z(n28837) );
  XNOR U28800 ( .A(n28834), .B(n28536), .Z(n28836) );
  IV U28801 ( .A(p_input[138]), .Z(n28536) );
  XOR U28802 ( .A(n28838), .B(n28839), .Z(n28834) );
  AND U28803 ( .A(n28840), .B(n28841), .Z(n28839) );
  XNOR U28804 ( .A(p_input[169]), .B(n28838), .Z(n28841) );
  XNOR U28805 ( .A(n28838), .B(n28545), .Z(n28840) );
  IV U28806 ( .A(p_input[137]), .Z(n28545) );
  XOR U28807 ( .A(n28842), .B(n28843), .Z(n28838) );
  AND U28808 ( .A(n28844), .B(n28845), .Z(n28843) );
  XNOR U28809 ( .A(p_input[168]), .B(n28842), .Z(n28845) );
  XNOR U28810 ( .A(n28842), .B(n28554), .Z(n28844) );
  IV U28811 ( .A(p_input[136]), .Z(n28554) );
  XOR U28812 ( .A(n28846), .B(n28847), .Z(n28842) );
  AND U28813 ( .A(n28848), .B(n28849), .Z(n28847) );
  XNOR U28814 ( .A(p_input[167]), .B(n28846), .Z(n28849) );
  XNOR U28815 ( .A(n28846), .B(n28563), .Z(n28848) );
  IV U28816 ( .A(p_input[135]), .Z(n28563) );
  XOR U28817 ( .A(n28850), .B(n28851), .Z(n28846) );
  AND U28818 ( .A(n28852), .B(n28853), .Z(n28851) );
  XNOR U28819 ( .A(p_input[166]), .B(n28850), .Z(n28853) );
  XNOR U28820 ( .A(n28850), .B(n28572), .Z(n28852) );
  IV U28821 ( .A(p_input[134]), .Z(n28572) );
  XOR U28822 ( .A(n28854), .B(n28855), .Z(n28850) );
  AND U28823 ( .A(n28856), .B(n28857), .Z(n28855) );
  XNOR U28824 ( .A(p_input[165]), .B(n28854), .Z(n28857) );
  XNOR U28825 ( .A(n28854), .B(n28581), .Z(n28856) );
  IV U28826 ( .A(p_input[133]), .Z(n28581) );
  XOR U28827 ( .A(n28858), .B(n28859), .Z(n28854) );
  AND U28828 ( .A(n28860), .B(n28861), .Z(n28859) );
  XNOR U28829 ( .A(p_input[164]), .B(n28858), .Z(n28861) );
  XNOR U28830 ( .A(n28858), .B(n28590), .Z(n28860) );
  IV U28831 ( .A(p_input[132]), .Z(n28590) );
  XOR U28832 ( .A(n28862), .B(n28863), .Z(n28858) );
  AND U28833 ( .A(n28864), .B(n28865), .Z(n28863) );
  XNOR U28834 ( .A(p_input[163]), .B(n28862), .Z(n28865) );
  XNOR U28835 ( .A(n28862), .B(n28599), .Z(n28864) );
  IV U28836 ( .A(p_input[131]), .Z(n28599) );
  XOR U28837 ( .A(n28866), .B(n28867), .Z(n28862) );
  AND U28838 ( .A(n28868), .B(n28869), .Z(n28867) );
  XNOR U28839 ( .A(p_input[162]), .B(n28866), .Z(n28869) );
  XNOR U28840 ( .A(n28866), .B(n28608), .Z(n28868) );
  IV U28841 ( .A(p_input[130]), .Z(n28608) );
  XNOR U28842 ( .A(n28870), .B(n28871), .Z(n28866) );
  AND U28843 ( .A(n28872), .B(n28873), .Z(n28871) );
  XOR U28844 ( .A(p_input[161]), .B(n28870), .Z(n28873) );
  XNOR U28845 ( .A(p_input[129]), .B(n28870), .Z(n28872) );
  AND U28846 ( .A(p_input[160]), .B(n28874), .Z(n28870) );
  IV U28847 ( .A(p_input[128]), .Z(n28874) );
  XOR U28848 ( .A(n28875), .B(n28876), .Z(n27964) );
  AND U28849 ( .A(n407), .B(n28877), .Z(n28876) );
  XNOR U28850 ( .A(n28878), .B(n28875), .Z(n28877) );
  XOR U28851 ( .A(n28879), .B(n28880), .Z(n407) );
  AND U28852 ( .A(n28881), .B(n28882), .Z(n28880) );
  XNOR U28853 ( .A(n27979), .B(n28879), .Z(n28882) );
  AND U28854 ( .A(p_input[95]), .B(p_input[127]), .Z(n27979) );
  XNOR U28855 ( .A(n28879), .B(n27976), .Z(n28881) );
  IV U28856 ( .A(n28883), .Z(n27976) );
  AND U28857 ( .A(p_input[31]), .B(p_input[63]), .Z(n28883) );
  XOR U28858 ( .A(n28884), .B(n28885), .Z(n28879) );
  AND U28859 ( .A(n28886), .B(n28887), .Z(n28885) );
  XOR U28860 ( .A(n28884), .B(n27991), .Z(n28887) );
  XNOR U28861 ( .A(p_input[94]), .B(n28888), .Z(n27991) );
  AND U28862 ( .A(n638), .B(n28889), .Z(n28888) );
  XOR U28863 ( .A(p_input[94]), .B(p_input[126]), .Z(n28889) );
  XNOR U28864 ( .A(n27988), .B(n28884), .Z(n28886) );
  XOR U28865 ( .A(n28890), .B(n28891), .Z(n27988) );
  AND U28866 ( .A(n635), .B(n28892), .Z(n28891) );
  XOR U28867 ( .A(p_input[62]), .B(p_input[30]), .Z(n28892) );
  XOR U28868 ( .A(n28893), .B(n28894), .Z(n28884) );
  AND U28869 ( .A(n28895), .B(n28896), .Z(n28894) );
  XOR U28870 ( .A(n28893), .B(n28003), .Z(n28896) );
  XNOR U28871 ( .A(p_input[93]), .B(n28897), .Z(n28003) );
  AND U28872 ( .A(n638), .B(n28898), .Z(n28897) );
  XOR U28873 ( .A(p_input[93]), .B(p_input[125]), .Z(n28898) );
  XNOR U28874 ( .A(n28000), .B(n28893), .Z(n28895) );
  XOR U28875 ( .A(n28899), .B(n28900), .Z(n28000) );
  AND U28876 ( .A(n635), .B(n28901), .Z(n28900) );
  XOR U28877 ( .A(p_input[61]), .B(p_input[29]), .Z(n28901) );
  XOR U28878 ( .A(n28902), .B(n28903), .Z(n28893) );
  AND U28879 ( .A(n28904), .B(n28905), .Z(n28903) );
  XOR U28880 ( .A(n28902), .B(n28015), .Z(n28905) );
  XNOR U28881 ( .A(p_input[92]), .B(n28906), .Z(n28015) );
  AND U28882 ( .A(n638), .B(n28907), .Z(n28906) );
  XOR U28883 ( .A(p_input[92]), .B(p_input[124]), .Z(n28907) );
  XNOR U28884 ( .A(n28012), .B(n28902), .Z(n28904) );
  XOR U28885 ( .A(n28908), .B(n28909), .Z(n28012) );
  AND U28886 ( .A(n635), .B(n28910), .Z(n28909) );
  XOR U28887 ( .A(p_input[60]), .B(p_input[28]), .Z(n28910) );
  XOR U28888 ( .A(n28911), .B(n28912), .Z(n28902) );
  AND U28889 ( .A(n28913), .B(n28914), .Z(n28912) );
  XOR U28890 ( .A(n28911), .B(n28027), .Z(n28914) );
  XNOR U28891 ( .A(p_input[91]), .B(n28915), .Z(n28027) );
  AND U28892 ( .A(n638), .B(n28916), .Z(n28915) );
  XOR U28893 ( .A(p_input[91]), .B(p_input[123]), .Z(n28916) );
  XNOR U28894 ( .A(n28024), .B(n28911), .Z(n28913) );
  XOR U28895 ( .A(n28917), .B(n28918), .Z(n28024) );
  AND U28896 ( .A(n635), .B(n28919), .Z(n28918) );
  XOR U28897 ( .A(p_input[59]), .B(p_input[27]), .Z(n28919) );
  XOR U28898 ( .A(n28920), .B(n28921), .Z(n28911) );
  AND U28899 ( .A(n28922), .B(n28923), .Z(n28921) );
  XOR U28900 ( .A(n28920), .B(n28039), .Z(n28923) );
  XNOR U28901 ( .A(p_input[90]), .B(n28924), .Z(n28039) );
  AND U28902 ( .A(n638), .B(n28925), .Z(n28924) );
  XOR U28903 ( .A(p_input[90]), .B(p_input[122]), .Z(n28925) );
  XNOR U28904 ( .A(n28036), .B(n28920), .Z(n28922) );
  XOR U28905 ( .A(n28926), .B(n28927), .Z(n28036) );
  AND U28906 ( .A(n635), .B(n28928), .Z(n28927) );
  XOR U28907 ( .A(p_input[58]), .B(p_input[26]), .Z(n28928) );
  XOR U28908 ( .A(n28929), .B(n28930), .Z(n28920) );
  AND U28909 ( .A(n28931), .B(n28932), .Z(n28930) );
  XOR U28910 ( .A(n28929), .B(n28051), .Z(n28932) );
  XNOR U28911 ( .A(p_input[89]), .B(n28933), .Z(n28051) );
  AND U28912 ( .A(n638), .B(n28934), .Z(n28933) );
  XOR U28913 ( .A(p_input[89]), .B(p_input[121]), .Z(n28934) );
  XNOR U28914 ( .A(n28048), .B(n28929), .Z(n28931) );
  XOR U28915 ( .A(n28935), .B(n28936), .Z(n28048) );
  AND U28916 ( .A(n635), .B(n28937), .Z(n28936) );
  XOR U28917 ( .A(p_input[57]), .B(p_input[25]), .Z(n28937) );
  XOR U28918 ( .A(n28938), .B(n28939), .Z(n28929) );
  AND U28919 ( .A(n28940), .B(n28941), .Z(n28939) );
  XOR U28920 ( .A(n28938), .B(n28063), .Z(n28941) );
  XNOR U28921 ( .A(p_input[88]), .B(n28942), .Z(n28063) );
  AND U28922 ( .A(n638), .B(n28943), .Z(n28942) );
  XOR U28923 ( .A(p_input[88]), .B(p_input[120]), .Z(n28943) );
  XNOR U28924 ( .A(n28060), .B(n28938), .Z(n28940) );
  XOR U28925 ( .A(n28944), .B(n28945), .Z(n28060) );
  AND U28926 ( .A(n635), .B(n28946), .Z(n28945) );
  XOR U28927 ( .A(p_input[56]), .B(p_input[24]), .Z(n28946) );
  XOR U28928 ( .A(n28947), .B(n28948), .Z(n28938) );
  AND U28929 ( .A(n28949), .B(n28950), .Z(n28948) );
  XOR U28930 ( .A(n28947), .B(n28075), .Z(n28950) );
  XNOR U28931 ( .A(p_input[87]), .B(n28951), .Z(n28075) );
  AND U28932 ( .A(n638), .B(n28952), .Z(n28951) );
  XOR U28933 ( .A(p_input[87]), .B(p_input[119]), .Z(n28952) );
  XNOR U28934 ( .A(n28072), .B(n28947), .Z(n28949) );
  XOR U28935 ( .A(n28953), .B(n28954), .Z(n28072) );
  AND U28936 ( .A(n635), .B(n28955), .Z(n28954) );
  XOR U28937 ( .A(p_input[55]), .B(p_input[23]), .Z(n28955) );
  XOR U28938 ( .A(n28956), .B(n28957), .Z(n28947) );
  AND U28939 ( .A(n28958), .B(n28959), .Z(n28957) );
  XOR U28940 ( .A(n28956), .B(n28087), .Z(n28959) );
  XNOR U28941 ( .A(p_input[86]), .B(n28960), .Z(n28087) );
  AND U28942 ( .A(n638), .B(n28961), .Z(n28960) );
  XOR U28943 ( .A(p_input[86]), .B(p_input[118]), .Z(n28961) );
  XNOR U28944 ( .A(n28084), .B(n28956), .Z(n28958) );
  XOR U28945 ( .A(n28962), .B(n28963), .Z(n28084) );
  AND U28946 ( .A(n635), .B(n28964), .Z(n28963) );
  XOR U28947 ( .A(p_input[54]), .B(p_input[22]), .Z(n28964) );
  XOR U28948 ( .A(n28965), .B(n28966), .Z(n28956) );
  AND U28949 ( .A(n28967), .B(n28968), .Z(n28966) );
  XOR U28950 ( .A(n28965), .B(n28099), .Z(n28968) );
  XNOR U28951 ( .A(p_input[85]), .B(n28969), .Z(n28099) );
  AND U28952 ( .A(n638), .B(n28970), .Z(n28969) );
  XOR U28953 ( .A(p_input[85]), .B(p_input[117]), .Z(n28970) );
  XNOR U28954 ( .A(n28096), .B(n28965), .Z(n28967) );
  XOR U28955 ( .A(n28971), .B(n28972), .Z(n28096) );
  AND U28956 ( .A(n635), .B(n28973), .Z(n28972) );
  XOR U28957 ( .A(p_input[53]), .B(p_input[21]), .Z(n28973) );
  XOR U28958 ( .A(n28974), .B(n28975), .Z(n28965) );
  AND U28959 ( .A(n28976), .B(n28977), .Z(n28975) );
  XOR U28960 ( .A(n28974), .B(n28111), .Z(n28977) );
  XNOR U28961 ( .A(p_input[84]), .B(n28978), .Z(n28111) );
  AND U28962 ( .A(n638), .B(n28979), .Z(n28978) );
  XOR U28963 ( .A(p_input[84]), .B(p_input[116]), .Z(n28979) );
  XNOR U28964 ( .A(n28108), .B(n28974), .Z(n28976) );
  XOR U28965 ( .A(n28980), .B(n28981), .Z(n28108) );
  AND U28966 ( .A(n635), .B(n28982), .Z(n28981) );
  XOR U28967 ( .A(p_input[52]), .B(p_input[20]), .Z(n28982) );
  XOR U28968 ( .A(n28983), .B(n28984), .Z(n28974) );
  AND U28969 ( .A(n28985), .B(n28986), .Z(n28984) );
  XOR U28970 ( .A(n28983), .B(n28123), .Z(n28986) );
  XNOR U28971 ( .A(p_input[83]), .B(n28987), .Z(n28123) );
  AND U28972 ( .A(n638), .B(n28988), .Z(n28987) );
  XOR U28973 ( .A(p_input[83]), .B(p_input[115]), .Z(n28988) );
  XNOR U28974 ( .A(n28120), .B(n28983), .Z(n28985) );
  XOR U28975 ( .A(n28989), .B(n28990), .Z(n28120) );
  AND U28976 ( .A(n635), .B(n28991), .Z(n28990) );
  XOR U28977 ( .A(p_input[51]), .B(p_input[19]), .Z(n28991) );
  XOR U28978 ( .A(n28992), .B(n28993), .Z(n28983) );
  AND U28979 ( .A(n28994), .B(n28995), .Z(n28993) );
  XOR U28980 ( .A(n28992), .B(n28135), .Z(n28995) );
  XNOR U28981 ( .A(p_input[82]), .B(n28996), .Z(n28135) );
  AND U28982 ( .A(n638), .B(n28997), .Z(n28996) );
  XOR U28983 ( .A(p_input[82]), .B(p_input[114]), .Z(n28997) );
  XNOR U28984 ( .A(n28132), .B(n28992), .Z(n28994) );
  XOR U28985 ( .A(n28998), .B(n28999), .Z(n28132) );
  AND U28986 ( .A(n635), .B(n29000), .Z(n28999) );
  XOR U28987 ( .A(p_input[50]), .B(p_input[18]), .Z(n29000) );
  XOR U28988 ( .A(n29001), .B(n29002), .Z(n28992) );
  AND U28989 ( .A(n29003), .B(n29004), .Z(n29002) );
  XOR U28990 ( .A(n29001), .B(n28147), .Z(n29004) );
  XNOR U28991 ( .A(p_input[81]), .B(n29005), .Z(n28147) );
  AND U28992 ( .A(n638), .B(n29006), .Z(n29005) );
  XOR U28993 ( .A(p_input[81]), .B(p_input[113]), .Z(n29006) );
  XNOR U28994 ( .A(n28144), .B(n29001), .Z(n29003) );
  XOR U28995 ( .A(n29007), .B(n29008), .Z(n28144) );
  AND U28996 ( .A(n635), .B(n29009), .Z(n29008) );
  XOR U28997 ( .A(p_input[49]), .B(p_input[17]), .Z(n29009) );
  XOR U28998 ( .A(n29010), .B(n29011), .Z(n29001) );
  AND U28999 ( .A(n29012), .B(n29013), .Z(n29011) );
  XOR U29000 ( .A(n29010), .B(n28159), .Z(n29013) );
  XNOR U29001 ( .A(p_input[80]), .B(n29014), .Z(n28159) );
  AND U29002 ( .A(n638), .B(n29015), .Z(n29014) );
  XOR U29003 ( .A(p_input[80]), .B(p_input[112]), .Z(n29015) );
  XNOR U29004 ( .A(n28156), .B(n29010), .Z(n29012) );
  XOR U29005 ( .A(n29016), .B(n29017), .Z(n28156) );
  AND U29006 ( .A(n635), .B(n29018), .Z(n29017) );
  XOR U29007 ( .A(p_input[48]), .B(p_input[16]), .Z(n29018) );
  XOR U29008 ( .A(n29019), .B(n29020), .Z(n29010) );
  AND U29009 ( .A(n29021), .B(n29022), .Z(n29020) );
  XOR U29010 ( .A(n29019), .B(n28171), .Z(n29022) );
  XNOR U29011 ( .A(p_input[79]), .B(n29023), .Z(n28171) );
  AND U29012 ( .A(n638), .B(n29024), .Z(n29023) );
  XOR U29013 ( .A(p_input[79]), .B(p_input[111]), .Z(n29024) );
  XNOR U29014 ( .A(n28168), .B(n29019), .Z(n29021) );
  XOR U29015 ( .A(n29025), .B(n29026), .Z(n28168) );
  AND U29016 ( .A(n635), .B(n29027), .Z(n29026) );
  XOR U29017 ( .A(p_input[47]), .B(p_input[15]), .Z(n29027) );
  XOR U29018 ( .A(n29028), .B(n29029), .Z(n29019) );
  AND U29019 ( .A(n29030), .B(n29031), .Z(n29029) );
  XOR U29020 ( .A(n29028), .B(n28183), .Z(n29031) );
  XNOR U29021 ( .A(p_input[78]), .B(n29032), .Z(n28183) );
  AND U29022 ( .A(n638), .B(n29033), .Z(n29032) );
  XOR U29023 ( .A(p_input[78]), .B(p_input[110]), .Z(n29033) );
  XNOR U29024 ( .A(n28180), .B(n29028), .Z(n29030) );
  XOR U29025 ( .A(n29034), .B(n29035), .Z(n28180) );
  AND U29026 ( .A(n635), .B(n29036), .Z(n29035) );
  XOR U29027 ( .A(p_input[46]), .B(p_input[14]), .Z(n29036) );
  XOR U29028 ( .A(n29037), .B(n29038), .Z(n29028) );
  AND U29029 ( .A(n29039), .B(n29040), .Z(n29038) );
  XOR U29030 ( .A(n29037), .B(n28195), .Z(n29040) );
  XNOR U29031 ( .A(p_input[77]), .B(n29041), .Z(n28195) );
  AND U29032 ( .A(n638), .B(n29042), .Z(n29041) );
  XOR U29033 ( .A(p_input[77]), .B(p_input[109]), .Z(n29042) );
  XNOR U29034 ( .A(n28192), .B(n29037), .Z(n29039) );
  XOR U29035 ( .A(n29043), .B(n29044), .Z(n28192) );
  AND U29036 ( .A(n635), .B(n29045), .Z(n29044) );
  XOR U29037 ( .A(p_input[45]), .B(p_input[13]), .Z(n29045) );
  XOR U29038 ( .A(n29046), .B(n29047), .Z(n29037) );
  AND U29039 ( .A(n29048), .B(n29049), .Z(n29047) );
  XOR U29040 ( .A(n29046), .B(n28207), .Z(n29049) );
  XNOR U29041 ( .A(p_input[76]), .B(n29050), .Z(n28207) );
  AND U29042 ( .A(n638), .B(n29051), .Z(n29050) );
  XOR U29043 ( .A(p_input[76]), .B(p_input[108]), .Z(n29051) );
  XNOR U29044 ( .A(n28204), .B(n29046), .Z(n29048) );
  XOR U29045 ( .A(n29052), .B(n29053), .Z(n28204) );
  AND U29046 ( .A(n635), .B(n29054), .Z(n29053) );
  XOR U29047 ( .A(p_input[44]), .B(p_input[12]), .Z(n29054) );
  XOR U29048 ( .A(n29055), .B(n29056), .Z(n29046) );
  AND U29049 ( .A(n29057), .B(n29058), .Z(n29056) );
  XOR U29050 ( .A(n29055), .B(n28219), .Z(n29058) );
  XNOR U29051 ( .A(p_input[75]), .B(n29059), .Z(n28219) );
  AND U29052 ( .A(n638), .B(n29060), .Z(n29059) );
  XOR U29053 ( .A(p_input[75]), .B(p_input[107]), .Z(n29060) );
  XNOR U29054 ( .A(n28216), .B(n29055), .Z(n29057) );
  XOR U29055 ( .A(n29061), .B(n29062), .Z(n28216) );
  AND U29056 ( .A(n635), .B(n29063), .Z(n29062) );
  XOR U29057 ( .A(p_input[43]), .B(p_input[11]), .Z(n29063) );
  XOR U29058 ( .A(n29064), .B(n29065), .Z(n29055) );
  AND U29059 ( .A(n29066), .B(n29067), .Z(n29065) );
  XOR U29060 ( .A(n29064), .B(n28231), .Z(n29067) );
  XNOR U29061 ( .A(p_input[74]), .B(n29068), .Z(n28231) );
  AND U29062 ( .A(n638), .B(n29069), .Z(n29068) );
  XOR U29063 ( .A(p_input[74]), .B(p_input[106]), .Z(n29069) );
  XNOR U29064 ( .A(n28228), .B(n29064), .Z(n29066) );
  XOR U29065 ( .A(n29070), .B(n29071), .Z(n28228) );
  AND U29066 ( .A(n635), .B(n29072), .Z(n29071) );
  XOR U29067 ( .A(p_input[42]), .B(p_input[10]), .Z(n29072) );
  XOR U29068 ( .A(n29073), .B(n29074), .Z(n29064) );
  AND U29069 ( .A(n29075), .B(n29076), .Z(n29074) );
  XOR U29070 ( .A(n29073), .B(n28243), .Z(n29076) );
  XNOR U29071 ( .A(p_input[73]), .B(n29077), .Z(n28243) );
  AND U29072 ( .A(n638), .B(n29078), .Z(n29077) );
  XOR U29073 ( .A(p_input[73]), .B(p_input[105]), .Z(n29078) );
  XNOR U29074 ( .A(n28240), .B(n29073), .Z(n29075) );
  XOR U29075 ( .A(n29079), .B(n29080), .Z(n28240) );
  AND U29076 ( .A(n635), .B(n29081), .Z(n29080) );
  XOR U29077 ( .A(p_input[9]), .B(p_input[41]), .Z(n29081) );
  XOR U29078 ( .A(n29082), .B(n29083), .Z(n29073) );
  AND U29079 ( .A(n29084), .B(n29085), .Z(n29083) );
  XOR U29080 ( .A(n29082), .B(n28255), .Z(n29085) );
  XNOR U29081 ( .A(p_input[72]), .B(n29086), .Z(n28255) );
  AND U29082 ( .A(n638), .B(n29087), .Z(n29086) );
  XOR U29083 ( .A(p_input[72]), .B(p_input[104]), .Z(n29087) );
  XNOR U29084 ( .A(n28252), .B(n29082), .Z(n29084) );
  XOR U29085 ( .A(n29088), .B(n29089), .Z(n28252) );
  AND U29086 ( .A(n635), .B(n29090), .Z(n29089) );
  XOR U29087 ( .A(p_input[8]), .B(p_input[40]), .Z(n29090) );
  XOR U29088 ( .A(n29091), .B(n29092), .Z(n29082) );
  AND U29089 ( .A(n29093), .B(n29094), .Z(n29092) );
  XOR U29090 ( .A(n29091), .B(n28267), .Z(n29094) );
  XNOR U29091 ( .A(p_input[71]), .B(n29095), .Z(n28267) );
  AND U29092 ( .A(n638), .B(n29096), .Z(n29095) );
  XOR U29093 ( .A(p_input[71]), .B(p_input[103]), .Z(n29096) );
  XNOR U29094 ( .A(n28264), .B(n29091), .Z(n29093) );
  XOR U29095 ( .A(n29097), .B(n29098), .Z(n28264) );
  AND U29096 ( .A(n635), .B(n29099), .Z(n29098) );
  XOR U29097 ( .A(p_input[7]), .B(p_input[39]), .Z(n29099) );
  XOR U29098 ( .A(n29100), .B(n29101), .Z(n29091) );
  AND U29099 ( .A(n29102), .B(n29103), .Z(n29101) );
  XOR U29100 ( .A(n29100), .B(n28279), .Z(n29103) );
  XNOR U29101 ( .A(p_input[70]), .B(n29104), .Z(n28279) );
  AND U29102 ( .A(n638), .B(n29105), .Z(n29104) );
  XOR U29103 ( .A(p_input[70]), .B(p_input[102]), .Z(n29105) );
  XNOR U29104 ( .A(n28276), .B(n29100), .Z(n29102) );
  XOR U29105 ( .A(n29106), .B(n29107), .Z(n28276) );
  AND U29106 ( .A(n635), .B(n29108), .Z(n29107) );
  XOR U29107 ( .A(p_input[6]), .B(p_input[38]), .Z(n29108) );
  XOR U29108 ( .A(n29109), .B(n29110), .Z(n29100) );
  AND U29109 ( .A(n29111), .B(n29112), .Z(n29110) );
  XOR U29110 ( .A(n29109), .B(n28291), .Z(n29112) );
  XNOR U29111 ( .A(p_input[69]), .B(n29113), .Z(n28291) );
  AND U29112 ( .A(n638), .B(n29114), .Z(n29113) );
  XOR U29113 ( .A(p_input[69]), .B(p_input[101]), .Z(n29114) );
  XNOR U29114 ( .A(n28288), .B(n29109), .Z(n29111) );
  XOR U29115 ( .A(n29115), .B(n29116), .Z(n28288) );
  AND U29116 ( .A(n635), .B(n29117), .Z(n29116) );
  XOR U29117 ( .A(p_input[5]), .B(p_input[37]), .Z(n29117) );
  XOR U29118 ( .A(n29118), .B(n29119), .Z(n29109) );
  AND U29119 ( .A(n29120), .B(n29121), .Z(n29119) );
  XOR U29120 ( .A(n29118), .B(n28303), .Z(n29121) );
  XNOR U29121 ( .A(p_input[68]), .B(n29122), .Z(n28303) );
  AND U29122 ( .A(n638), .B(n29123), .Z(n29122) );
  XOR U29123 ( .A(p_input[68]), .B(p_input[100]), .Z(n29123) );
  XNOR U29124 ( .A(n28300), .B(n29118), .Z(n29120) );
  XOR U29125 ( .A(n29124), .B(n29125), .Z(n28300) );
  AND U29126 ( .A(n635), .B(n29126), .Z(n29125) );
  XOR U29127 ( .A(p_input[4]), .B(p_input[36]), .Z(n29126) );
  XOR U29128 ( .A(n29127), .B(n29128), .Z(n29118) );
  AND U29129 ( .A(n29129), .B(n29130), .Z(n29128) );
  XOR U29130 ( .A(n29127), .B(n28315), .Z(n29130) );
  XNOR U29131 ( .A(p_input[67]), .B(n29131), .Z(n28315) );
  AND U29132 ( .A(n638), .B(n29132), .Z(n29131) );
  XOR U29133 ( .A(p_input[99]), .B(p_input[67]), .Z(n29132) );
  XNOR U29134 ( .A(n28312), .B(n29127), .Z(n29129) );
  XOR U29135 ( .A(n29133), .B(n29134), .Z(n28312) );
  AND U29136 ( .A(n635), .B(n29135), .Z(n29134) );
  XOR U29137 ( .A(p_input[3]), .B(p_input[35]), .Z(n29135) );
  XOR U29138 ( .A(n29136), .B(n29137), .Z(n29127) );
  AND U29139 ( .A(n29138), .B(n29139), .Z(n29137) );
  XOR U29140 ( .A(n28327), .B(n29136), .Z(n29139) );
  XNOR U29141 ( .A(p_input[66]), .B(n29140), .Z(n28327) );
  AND U29142 ( .A(n638), .B(n29141), .Z(n29140) );
  XOR U29143 ( .A(p_input[98]), .B(p_input[66]), .Z(n29141) );
  XNOR U29144 ( .A(n29136), .B(n28324), .Z(n29138) );
  XOR U29145 ( .A(n29142), .B(n29143), .Z(n28324) );
  AND U29146 ( .A(n635), .B(n29144), .Z(n29143) );
  XOR U29147 ( .A(p_input[34]), .B(p_input[2]), .Z(n29144) );
  XOR U29148 ( .A(n29145), .B(n29146), .Z(n29136) );
  AND U29149 ( .A(n29147), .B(n29148), .Z(n29146) );
  XNOR U29150 ( .A(n29149), .B(n28340), .Z(n29148) );
  XNOR U29151 ( .A(p_input[65]), .B(n29150), .Z(n28340) );
  AND U29152 ( .A(n638), .B(n29151), .Z(n29150) );
  XNOR U29153 ( .A(p_input[97]), .B(n29152), .Z(n29151) );
  IV U29154 ( .A(p_input[65]), .Z(n29152) );
  XNOR U29155 ( .A(n28337), .B(n29145), .Z(n29147) );
  XNOR U29156 ( .A(p_input[1]), .B(n29153), .Z(n28337) );
  AND U29157 ( .A(n635), .B(n29154), .Z(n29153) );
  XOR U29158 ( .A(p_input[33]), .B(p_input[1]), .Z(n29154) );
  IV U29159 ( .A(n29149), .Z(n29145) );
  AND U29160 ( .A(n28875), .B(n28878), .Z(n29149) );
  XOR U29161 ( .A(p_input[64]), .B(n29155), .Z(n28878) );
  AND U29162 ( .A(n638), .B(n29156), .Z(n29155) );
  XOR U29163 ( .A(p_input[96]), .B(p_input[64]), .Z(n29156) );
  XOR U29164 ( .A(n29157), .B(n29158), .Z(n638) );
  AND U29165 ( .A(n29159), .B(n29160), .Z(n29158) );
  XNOR U29166 ( .A(p_input[127]), .B(n29157), .Z(n29160) );
  XOR U29167 ( .A(n29157), .B(p_input[95]), .Z(n29159) );
  XOR U29168 ( .A(n29161), .B(n29162), .Z(n29157) );
  AND U29169 ( .A(n29163), .B(n29164), .Z(n29162) );
  XNOR U29170 ( .A(p_input[126]), .B(n29161), .Z(n29164) );
  XOR U29171 ( .A(n29161), .B(p_input[94]), .Z(n29163) );
  XOR U29172 ( .A(n29165), .B(n29166), .Z(n29161) );
  AND U29173 ( .A(n29167), .B(n29168), .Z(n29166) );
  XNOR U29174 ( .A(p_input[125]), .B(n29165), .Z(n29168) );
  XOR U29175 ( .A(n29165), .B(p_input[93]), .Z(n29167) );
  XOR U29176 ( .A(n29169), .B(n29170), .Z(n29165) );
  AND U29177 ( .A(n29171), .B(n29172), .Z(n29170) );
  XNOR U29178 ( .A(p_input[124]), .B(n29169), .Z(n29172) );
  XOR U29179 ( .A(n29169), .B(p_input[92]), .Z(n29171) );
  XOR U29180 ( .A(n29173), .B(n29174), .Z(n29169) );
  AND U29181 ( .A(n29175), .B(n29176), .Z(n29174) );
  XNOR U29182 ( .A(p_input[123]), .B(n29173), .Z(n29176) );
  XOR U29183 ( .A(n29173), .B(p_input[91]), .Z(n29175) );
  XOR U29184 ( .A(n29177), .B(n29178), .Z(n29173) );
  AND U29185 ( .A(n29179), .B(n29180), .Z(n29178) );
  XNOR U29186 ( .A(p_input[122]), .B(n29177), .Z(n29180) );
  XOR U29187 ( .A(n29177), .B(p_input[90]), .Z(n29179) );
  XOR U29188 ( .A(n29181), .B(n29182), .Z(n29177) );
  AND U29189 ( .A(n29183), .B(n29184), .Z(n29182) );
  XNOR U29190 ( .A(p_input[121]), .B(n29181), .Z(n29184) );
  XOR U29191 ( .A(n29181), .B(p_input[89]), .Z(n29183) );
  XOR U29192 ( .A(n29185), .B(n29186), .Z(n29181) );
  AND U29193 ( .A(n29187), .B(n29188), .Z(n29186) );
  XNOR U29194 ( .A(p_input[120]), .B(n29185), .Z(n29188) );
  XOR U29195 ( .A(n29185), .B(p_input[88]), .Z(n29187) );
  XOR U29196 ( .A(n29189), .B(n29190), .Z(n29185) );
  AND U29197 ( .A(n29191), .B(n29192), .Z(n29190) );
  XNOR U29198 ( .A(p_input[119]), .B(n29189), .Z(n29192) );
  XOR U29199 ( .A(n29189), .B(p_input[87]), .Z(n29191) );
  XOR U29200 ( .A(n29193), .B(n29194), .Z(n29189) );
  AND U29201 ( .A(n29195), .B(n29196), .Z(n29194) );
  XNOR U29202 ( .A(p_input[118]), .B(n29193), .Z(n29196) );
  XOR U29203 ( .A(n29193), .B(p_input[86]), .Z(n29195) );
  XOR U29204 ( .A(n29197), .B(n29198), .Z(n29193) );
  AND U29205 ( .A(n29199), .B(n29200), .Z(n29198) );
  XNOR U29206 ( .A(p_input[117]), .B(n29197), .Z(n29200) );
  XOR U29207 ( .A(n29197), .B(p_input[85]), .Z(n29199) );
  XOR U29208 ( .A(n29201), .B(n29202), .Z(n29197) );
  AND U29209 ( .A(n29203), .B(n29204), .Z(n29202) );
  XNOR U29210 ( .A(p_input[116]), .B(n29201), .Z(n29204) );
  XOR U29211 ( .A(n29201), .B(p_input[84]), .Z(n29203) );
  XOR U29212 ( .A(n29205), .B(n29206), .Z(n29201) );
  AND U29213 ( .A(n29207), .B(n29208), .Z(n29206) );
  XNOR U29214 ( .A(p_input[115]), .B(n29205), .Z(n29208) );
  XOR U29215 ( .A(n29205), .B(p_input[83]), .Z(n29207) );
  XOR U29216 ( .A(n29209), .B(n29210), .Z(n29205) );
  AND U29217 ( .A(n29211), .B(n29212), .Z(n29210) );
  XNOR U29218 ( .A(p_input[114]), .B(n29209), .Z(n29212) );
  XOR U29219 ( .A(n29209), .B(p_input[82]), .Z(n29211) );
  XOR U29220 ( .A(n29213), .B(n29214), .Z(n29209) );
  AND U29221 ( .A(n29215), .B(n29216), .Z(n29214) );
  XNOR U29222 ( .A(p_input[113]), .B(n29213), .Z(n29216) );
  XOR U29223 ( .A(n29213), .B(p_input[81]), .Z(n29215) );
  XOR U29224 ( .A(n29217), .B(n29218), .Z(n29213) );
  AND U29225 ( .A(n29219), .B(n29220), .Z(n29218) );
  XNOR U29226 ( .A(p_input[112]), .B(n29217), .Z(n29220) );
  XOR U29227 ( .A(n29217), .B(p_input[80]), .Z(n29219) );
  XOR U29228 ( .A(n29221), .B(n29222), .Z(n29217) );
  AND U29229 ( .A(n29223), .B(n29224), .Z(n29222) );
  XNOR U29230 ( .A(p_input[111]), .B(n29221), .Z(n29224) );
  XOR U29231 ( .A(n29221), .B(p_input[79]), .Z(n29223) );
  XOR U29232 ( .A(n29225), .B(n29226), .Z(n29221) );
  AND U29233 ( .A(n29227), .B(n29228), .Z(n29226) );
  XNOR U29234 ( .A(p_input[110]), .B(n29225), .Z(n29228) );
  XOR U29235 ( .A(n29225), .B(p_input[78]), .Z(n29227) );
  XOR U29236 ( .A(n29229), .B(n29230), .Z(n29225) );
  AND U29237 ( .A(n29231), .B(n29232), .Z(n29230) );
  XNOR U29238 ( .A(p_input[109]), .B(n29229), .Z(n29232) );
  XOR U29239 ( .A(n29229), .B(p_input[77]), .Z(n29231) );
  XOR U29240 ( .A(n29233), .B(n29234), .Z(n29229) );
  AND U29241 ( .A(n29235), .B(n29236), .Z(n29234) );
  XNOR U29242 ( .A(p_input[108]), .B(n29233), .Z(n29236) );
  XOR U29243 ( .A(n29233), .B(p_input[76]), .Z(n29235) );
  XOR U29244 ( .A(n29237), .B(n29238), .Z(n29233) );
  AND U29245 ( .A(n29239), .B(n29240), .Z(n29238) );
  XNOR U29246 ( .A(p_input[107]), .B(n29237), .Z(n29240) );
  XOR U29247 ( .A(n29237), .B(p_input[75]), .Z(n29239) );
  XOR U29248 ( .A(n29241), .B(n29242), .Z(n29237) );
  AND U29249 ( .A(n29243), .B(n29244), .Z(n29242) );
  XNOR U29250 ( .A(p_input[106]), .B(n29241), .Z(n29244) );
  XOR U29251 ( .A(n29241), .B(p_input[74]), .Z(n29243) );
  XOR U29252 ( .A(n29245), .B(n29246), .Z(n29241) );
  AND U29253 ( .A(n29247), .B(n29248), .Z(n29246) );
  XNOR U29254 ( .A(p_input[105]), .B(n29245), .Z(n29248) );
  XOR U29255 ( .A(n29245), .B(p_input[73]), .Z(n29247) );
  XOR U29256 ( .A(n29249), .B(n29250), .Z(n29245) );
  AND U29257 ( .A(n29251), .B(n29252), .Z(n29250) );
  XNOR U29258 ( .A(p_input[104]), .B(n29249), .Z(n29252) );
  XOR U29259 ( .A(n29249), .B(p_input[72]), .Z(n29251) );
  XOR U29260 ( .A(n29253), .B(n29254), .Z(n29249) );
  AND U29261 ( .A(n29255), .B(n29256), .Z(n29254) );
  XNOR U29262 ( .A(p_input[103]), .B(n29253), .Z(n29256) );
  XOR U29263 ( .A(n29253), .B(p_input[71]), .Z(n29255) );
  XOR U29264 ( .A(n29257), .B(n29258), .Z(n29253) );
  AND U29265 ( .A(n29259), .B(n29260), .Z(n29258) );
  XNOR U29266 ( .A(p_input[102]), .B(n29257), .Z(n29260) );
  XOR U29267 ( .A(n29257), .B(p_input[70]), .Z(n29259) );
  XOR U29268 ( .A(n29261), .B(n29262), .Z(n29257) );
  AND U29269 ( .A(n29263), .B(n29264), .Z(n29262) );
  XNOR U29270 ( .A(p_input[101]), .B(n29261), .Z(n29264) );
  XOR U29271 ( .A(n29261), .B(p_input[69]), .Z(n29263) );
  XOR U29272 ( .A(n29265), .B(n29266), .Z(n29261) );
  AND U29273 ( .A(n29267), .B(n29268), .Z(n29266) );
  XNOR U29274 ( .A(p_input[100]), .B(n29265), .Z(n29268) );
  XOR U29275 ( .A(n29265), .B(p_input[68]), .Z(n29267) );
  XOR U29276 ( .A(n29269), .B(n29270), .Z(n29265) );
  AND U29277 ( .A(n29271), .B(n29272), .Z(n29270) );
  XNOR U29278 ( .A(p_input[99]), .B(n29269), .Z(n29272) );
  XOR U29279 ( .A(n29269), .B(p_input[67]), .Z(n29271) );
  XOR U29280 ( .A(n29273), .B(n29274), .Z(n29269) );
  AND U29281 ( .A(n29275), .B(n29276), .Z(n29274) );
  XNOR U29282 ( .A(p_input[98]), .B(n29273), .Z(n29276) );
  XOR U29283 ( .A(n29273), .B(p_input[66]), .Z(n29275) );
  XNOR U29284 ( .A(n29277), .B(n29278), .Z(n29273) );
  AND U29285 ( .A(n29279), .B(n29280), .Z(n29278) );
  XOR U29286 ( .A(p_input[97]), .B(n29277), .Z(n29280) );
  XNOR U29287 ( .A(p_input[65]), .B(n29277), .Z(n29279) );
  AND U29288 ( .A(p_input[96]), .B(n29281), .Z(n29277) );
  IV U29289 ( .A(p_input[64]), .Z(n29281) );
  XNOR U29290 ( .A(p_input[0]), .B(n29282), .Z(n28875) );
  AND U29291 ( .A(n635), .B(n29283), .Z(n29282) );
  XOR U29292 ( .A(p_input[32]), .B(p_input[0]), .Z(n29283) );
  XOR U29293 ( .A(n29284), .B(n29285), .Z(n635) );
  AND U29294 ( .A(n29286), .B(n29287), .Z(n29285) );
  XNOR U29295 ( .A(p_input[63]), .B(n29284), .Z(n29287) );
  XOR U29296 ( .A(n29284), .B(p_input[31]), .Z(n29286) );
  XOR U29297 ( .A(n29288), .B(n29289), .Z(n29284) );
  AND U29298 ( .A(n29290), .B(n29291), .Z(n29289) );
  XNOR U29299 ( .A(p_input[62]), .B(n29288), .Z(n29291) );
  XNOR U29300 ( .A(n29288), .B(n28890), .Z(n29290) );
  IV U29301 ( .A(p_input[30]), .Z(n28890) );
  XOR U29302 ( .A(n29292), .B(n29293), .Z(n29288) );
  AND U29303 ( .A(n29294), .B(n29295), .Z(n29293) );
  XNOR U29304 ( .A(p_input[61]), .B(n29292), .Z(n29295) );
  XNOR U29305 ( .A(n29292), .B(n28899), .Z(n29294) );
  IV U29306 ( .A(p_input[29]), .Z(n28899) );
  XOR U29307 ( .A(n29296), .B(n29297), .Z(n29292) );
  AND U29308 ( .A(n29298), .B(n29299), .Z(n29297) );
  XNOR U29309 ( .A(p_input[60]), .B(n29296), .Z(n29299) );
  XNOR U29310 ( .A(n29296), .B(n28908), .Z(n29298) );
  IV U29311 ( .A(p_input[28]), .Z(n28908) );
  XOR U29312 ( .A(n29300), .B(n29301), .Z(n29296) );
  AND U29313 ( .A(n29302), .B(n29303), .Z(n29301) );
  XNOR U29314 ( .A(p_input[59]), .B(n29300), .Z(n29303) );
  XNOR U29315 ( .A(n29300), .B(n28917), .Z(n29302) );
  IV U29316 ( .A(p_input[27]), .Z(n28917) );
  XOR U29317 ( .A(n29304), .B(n29305), .Z(n29300) );
  AND U29318 ( .A(n29306), .B(n29307), .Z(n29305) );
  XNOR U29319 ( .A(p_input[58]), .B(n29304), .Z(n29307) );
  XNOR U29320 ( .A(n29304), .B(n28926), .Z(n29306) );
  IV U29321 ( .A(p_input[26]), .Z(n28926) );
  XOR U29322 ( .A(n29308), .B(n29309), .Z(n29304) );
  AND U29323 ( .A(n29310), .B(n29311), .Z(n29309) );
  XNOR U29324 ( .A(p_input[57]), .B(n29308), .Z(n29311) );
  XNOR U29325 ( .A(n29308), .B(n28935), .Z(n29310) );
  IV U29326 ( .A(p_input[25]), .Z(n28935) );
  XOR U29327 ( .A(n29312), .B(n29313), .Z(n29308) );
  AND U29328 ( .A(n29314), .B(n29315), .Z(n29313) );
  XNOR U29329 ( .A(p_input[56]), .B(n29312), .Z(n29315) );
  XNOR U29330 ( .A(n29312), .B(n28944), .Z(n29314) );
  IV U29331 ( .A(p_input[24]), .Z(n28944) );
  XOR U29332 ( .A(n29316), .B(n29317), .Z(n29312) );
  AND U29333 ( .A(n29318), .B(n29319), .Z(n29317) );
  XNOR U29334 ( .A(p_input[55]), .B(n29316), .Z(n29319) );
  XNOR U29335 ( .A(n29316), .B(n28953), .Z(n29318) );
  IV U29336 ( .A(p_input[23]), .Z(n28953) );
  XOR U29337 ( .A(n29320), .B(n29321), .Z(n29316) );
  AND U29338 ( .A(n29322), .B(n29323), .Z(n29321) );
  XNOR U29339 ( .A(p_input[54]), .B(n29320), .Z(n29323) );
  XNOR U29340 ( .A(n29320), .B(n28962), .Z(n29322) );
  IV U29341 ( .A(p_input[22]), .Z(n28962) );
  XOR U29342 ( .A(n29324), .B(n29325), .Z(n29320) );
  AND U29343 ( .A(n29326), .B(n29327), .Z(n29325) );
  XNOR U29344 ( .A(p_input[53]), .B(n29324), .Z(n29327) );
  XNOR U29345 ( .A(n29324), .B(n28971), .Z(n29326) );
  IV U29346 ( .A(p_input[21]), .Z(n28971) );
  XOR U29347 ( .A(n29328), .B(n29329), .Z(n29324) );
  AND U29348 ( .A(n29330), .B(n29331), .Z(n29329) );
  XNOR U29349 ( .A(p_input[52]), .B(n29328), .Z(n29331) );
  XNOR U29350 ( .A(n29328), .B(n28980), .Z(n29330) );
  IV U29351 ( .A(p_input[20]), .Z(n28980) );
  XOR U29352 ( .A(n29332), .B(n29333), .Z(n29328) );
  AND U29353 ( .A(n29334), .B(n29335), .Z(n29333) );
  XNOR U29354 ( .A(p_input[51]), .B(n29332), .Z(n29335) );
  XNOR U29355 ( .A(n29332), .B(n28989), .Z(n29334) );
  IV U29356 ( .A(p_input[19]), .Z(n28989) );
  XOR U29357 ( .A(n29336), .B(n29337), .Z(n29332) );
  AND U29358 ( .A(n29338), .B(n29339), .Z(n29337) );
  XNOR U29359 ( .A(p_input[50]), .B(n29336), .Z(n29339) );
  XNOR U29360 ( .A(n29336), .B(n28998), .Z(n29338) );
  IV U29361 ( .A(p_input[18]), .Z(n28998) );
  XOR U29362 ( .A(n29340), .B(n29341), .Z(n29336) );
  AND U29363 ( .A(n29342), .B(n29343), .Z(n29341) );
  XNOR U29364 ( .A(p_input[49]), .B(n29340), .Z(n29343) );
  XNOR U29365 ( .A(n29340), .B(n29007), .Z(n29342) );
  IV U29366 ( .A(p_input[17]), .Z(n29007) );
  XOR U29367 ( .A(n29344), .B(n29345), .Z(n29340) );
  AND U29368 ( .A(n29346), .B(n29347), .Z(n29345) );
  XNOR U29369 ( .A(p_input[48]), .B(n29344), .Z(n29347) );
  XNOR U29370 ( .A(n29344), .B(n29016), .Z(n29346) );
  IV U29371 ( .A(p_input[16]), .Z(n29016) );
  XOR U29372 ( .A(n29348), .B(n29349), .Z(n29344) );
  AND U29373 ( .A(n29350), .B(n29351), .Z(n29349) );
  XNOR U29374 ( .A(p_input[47]), .B(n29348), .Z(n29351) );
  XNOR U29375 ( .A(n29348), .B(n29025), .Z(n29350) );
  IV U29376 ( .A(p_input[15]), .Z(n29025) );
  XOR U29377 ( .A(n29352), .B(n29353), .Z(n29348) );
  AND U29378 ( .A(n29354), .B(n29355), .Z(n29353) );
  XNOR U29379 ( .A(p_input[46]), .B(n29352), .Z(n29355) );
  XNOR U29380 ( .A(n29352), .B(n29034), .Z(n29354) );
  IV U29381 ( .A(p_input[14]), .Z(n29034) );
  XOR U29382 ( .A(n29356), .B(n29357), .Z(n29352) );
  AND U29383 ( .A(n29358), .B(n29359), .Z(n29357) );
  XNOR U29384 ( .A(p_input[45]), .B(n29356), .Z(n29359) );
  XNOR U29385 ( .A(n29356), .B(n29043), .Z(n29358) );
  IV U29386 ( .A(p_input[13]), .Z(n29043) );
  XOR U29387 ( .A(n29360), .B(n29361), .Z(n29356) );
  AND U29388 ( .A(n29362), .B(n29363), .Z(n29361) );
  XNOR U29389 ( .A(p_input[44]), .B(n29360), .Z(n29363) );
  XNOR U29390 ( .A(n29360), .B(n29052), .Z(n29362) );
  IV U29391 ( .A(p_input[12]), .Z(n29052) );
  XOR U29392 ( .A(n29364), .B(n29365), .Z(n29360) );
  AND U29393 ( .A(n29366), .B(n29367), .Z(n29365) );
  XNOR U29394 ( .A(p_input[43]), .B(n29364), .Z(n29367) );
  XNOR U29395 ( .A(n29364), .B(n29061), .Z(n29366) );
  IV U29396 ( .A(p_input[11]), .Z(n29061) );
  XOR U29397 ( .A(n29368), .B(n29369), .Z(n29364) );
  AND U29398 ( .A(n29370), .B(n29371), .Z(n29369) );
  XNOR U29399 ( .A(p_input[42]), .B(n29368), .Z(n29371) );
  XNOR U29400 ( .A(n29368), .B(n29070), .Z(n29370) );
  IV U29401 ( .A(p_input[10]), .Z(n29070) );
  XOR U29402 ( .A(n29372), .B(n29373), .Z(n29368) );
  AND U29403 ( .A(n29374), .B(n29375), .Z(n29373) );
  XNOR U29404 ( .A(p_input[41]), .B(n29372), .Z(n29375) );
  XNOR U29405 ( .A(n29372), .B(n29079), .Z(n29374) );
  IV U29406 ( .A(p_input[9]), .Z(n29079) );
  XOR U29407 ( .A(n29376), .B(n29377), .Z(n29372) );
  AND U29408 ( .A(n29378), .B(n29379), .Z(n29377) );
  XNOR U29409 ( .A(p_input[40]), .B(n29376), .Z(n29379) );
  XNOR U29410 ( .A(n29376), .B(n29088), .Z(n29378) );
  IV U29411 ( .A(p_input[8]), .Z(n29088) );
  XOR U29412 ( .A(n29380), .B(n29381), .Z(n29376) );
  AND U29413 ( .A(n29382), .B(n29383), .Z(n29381) );
  XNOR U29414 ( .A(p_input[39]), .B(n29380), .Z(n29383) );
  XNOR U29415 ( .A(n29380), .B(n29097), .Z(n29382) );
  IV U29416 ( .A(p_input[7]), .Z(n29097) );
  XOR U29417 ( .A(n29384), .B(n29385), .Z(n29380) );
  AND U29418 ( .A(n29386), .B(n29387), .Z(n29385) );
  XNOR U29419 ( .A(p_input[38]), .B(n29384), .Z(n29387) );
  XNOR U29420 ( .A(n29384), .B(n29106), .Z(n29386) );
  IV U29421 ( .A(p_input[6]), .Z(n29106) );
  XOR U29422 ( .A(n29388), .B(n29389), .Z(n29384) );
  AND U29423 ( .A(n29390), .B(n29391), .Z(n29389) );
  XNOR U29424 ( .A(p_input[37]), .B(n29388), .Z(n29391) );
  XNOR U29425 ( .A(n29388), .B(n29115), .Z(n29390) );
  IV U29426 ( .A(p_input[5]), .Z(n29115) );
  XOR U29427 ( .A(n29392), .B(n29393), .Z(n29388) );
  AND U29428 ( .A(n29394), .B(n29395), .Z(n29393) );
  XNOR U29429 ( .A(p_input[36]), .B(n29392), .Z(n29395) );
  XNOR U29430 ( .A(n29392), .B(n29124), .Z(n29394) );
  IV U29431 ( .A(p_input[4]), .Z(n29124) );
  XOR U29432 ( .A(n29396), .B(n29397), .Z(n29392) );
  AND U29433 ( .A(n29398), .B(n29399), .Z(n29397) );
  XNOR U29434 ( .A(p_input[35]), .B(n29396), .Z(n29399) );
  XNOR U29435 ( .A(n29396), .B(n29133), .Z(n29398) );
  IV U29436 ( .A(p_input[3]), .Z(n29133) );
  XOR U29437 ( .A(n29400), .B(n29401), .Z(n29396) );
  AND U29438 ( .A(n29402), .B(n29403), .Z(n29401) );
  XNOR U29439 ( .A(p_input[34]), .B(n29400), .Z(n29403) );
  XNOR U29440 ( .A(n29400), .B(n29142), .Z(n29402) );
  IV U29441 ( .A(p_input[2]), .Z(n29142) );
  XNOR U29442 ( .A(n29404), .B(n29405), .Z(n29400) );
  AND U29443 ( .A(n29406), .B(n29407), .Z(n29405) );
  XOR U29444 ( .A(p_input[33]), .B(n29404), .Z(n29407) );
  XNOR U29445 ( .A(p_input[1]), .B(n29404), .Z(n29406) );
  AND U29446 ( .A(p_input[32]), .B(n29408), .Z(n29404) );
  IV U29447 ( .A(p_input[0]), .Z(n29408) );
endmodule

