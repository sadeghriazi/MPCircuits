
module voting_N2_M9 ( p_input, o );
  input [1023:0] p_input;
  output [1:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641,
         n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
         n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
         n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
         n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
         n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
         n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
         n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
         n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785,
         n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
         n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
         n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
         n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849,
         n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857,
         n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
         n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
         n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
         n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897,
         n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
         n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
         n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921,
         n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929,
         n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
         n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945,
         n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
         n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
         n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969,
         n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
         n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985,
         n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993,
         n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001,
         n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
         n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017,
         n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
         n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033,
         n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041,
         n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
         n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057,
         n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065,
         n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073,
         n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
         n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089,
         n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
         n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
         n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113,
         n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
         n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129,
         n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137,
         n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145,
         n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
         n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161,
         n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
         n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
         n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185,
         n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193,
         n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
         n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209,
         n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217,
         n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
         n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233,
         n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
         n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249,
         n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257,
         n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265,
         n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
         n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281,
         n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289,
         n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
         n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305,
         n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
         n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321,
         n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329,
         n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
         n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
         n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353,
         n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361,
         n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
         n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377,
         n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
         n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393,
         n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401,
         n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
         n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417,
         n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425,
         n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433,
         n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
         n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449,
         n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
         n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
         n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
         n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
         n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
         n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497,
         n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
         n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
         n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521,
         n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
         n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
         n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
         n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553,
         n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561,
         n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569,
         n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577,
         n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
         n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593,
         n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
         n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
         n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617,
         n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
         n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633,
         n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641,
         n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649,
         n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
         n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665,
         n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
         n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
         n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689,
         n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
         n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705,
         n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713,
         n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
         n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
         n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
         n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
         n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
         n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761,
         n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769,
         n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777,
         n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785,
         n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793,
         n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
         n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
         n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
         n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
         n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833,
         n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841,
         n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849,
         n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857,
         n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865,
         n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
         n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881,
         n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
         n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
         n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905,
         n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913,
         n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921,
         n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929,
         n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
         n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
         n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953,
         n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
         n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969,
         n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977,
         n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985,
         n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993,
         n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
         n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009,
         n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
         n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025,
         n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
         n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041,
         n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
         n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057,
         n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
         n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
         n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081,
         n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
         n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097,
         n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
         n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113,
         n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121,
         n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129,
         n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137,
         n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
         n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153,
         n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
         n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169,
         n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
         n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185,
         n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193,
         n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201,
         n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
         n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217,
         n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225,
         n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
         n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241,
         n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
         n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257,
         n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
         n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273,
         n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
         n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289,
         n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297,
         n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305,
         n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313,
         n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
         n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
         n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337,
         n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345,
         n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353,
         n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361,
         n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369,
         n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377,
         n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385,
         n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
         n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401,
         n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409,
         n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417,
         n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425,
         n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433,
         n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441,
         n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
         n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
         n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465,
         n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473,
         n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481,
         n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489,
         n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497,
         n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505,
         n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513,
         n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
         n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529,
         n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537,
         n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545,
         n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553,
         n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561,
         n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569,
         n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577,
         n38578, n38579, n38580, n38581, n38582, n38583, n38584, n38585,
         n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593,
         n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601,
         n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609,
         n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617,
         n38618, n38619, n38620, n38621, n38622, n38623, n38624, n38625,
         n38626, n38627, n38628, n38629, n38630, n38631, n38632, n38633,
         n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641,
         n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649,
         n38650, n38651, n38652, n38653, n38654, n38655, n38656, n38657,
         n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665,
         n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673,
         n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681,
         n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689,
         n38690, n38691, n38692, n38693, n38694, n38695, n38696, n38697,
         n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705,
         n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713,
         n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721,
         n38722, n38723, n38724, n38725, n38726, n38727, n38728, n38729,
         n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737,
         n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745,
         n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753,
         n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761,
         n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769,
         n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777,
         n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785,
         n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793,
         n38794, n38795, n38796, n38797, n38798, n38799, n38800, n38801,
         n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809,
         n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817,
         n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825,
         n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833,
         n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841,
         n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849,
         n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857,
         n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865,
         n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873,
         n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881,
         n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889,
         n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897,
         n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905,
         n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913,
         n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921,
         n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929,
         n38930, n38931, n38932, n38933, n38934, n38935, n38936, n38937,
         n38938, n38939, n38940, n38941, n38942, n38943, n38944, n38945,
         n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953,
         n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961,
         n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969,
         n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977,
         n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985,
         n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993,
         n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001,
         n39002, n39003, n39004, n39005, n39006, n39007, n39008, n39009,
         n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017,
         n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025,
         n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033,
         n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041,
         n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049,
         n39050, n39051, n39052, n39053, n39054, n39055, n39056, n39057,
         n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065,
         n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073,
         n39074, n39075, n39076, n39077, n39078, n39079, n39080, n39081,
         n39082, n39083, n39084, n39085, n39086, n39087, n39088, n39089,
         n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097,
         n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105,
         n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113,
         n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121,
         n39122, n39123, n39124, n39125, n39126, n39127, n39128, n39129,
         n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137,
         n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145,
         n39146, n39147, n39148, n39149, n39150, n39151, n39152, n39153,
         n39154, n39155, n39156, n39157, n39158, n39159, n39160, n39161,
         n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169,
         n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177,
         n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185,
         n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193,
         n39194, n39195, n39196, n39197, n39198, n39199, n39200, n39201,
         n39202, n39203, n39204, n39205, n39206, n39207, n39208, n39209,
         n39210, n39211, n39212, n39213, n39214, n39215, n39216, n39217,
         n39218, n39219, n39220, n39221, n39222, n39223, n39224, n39225,
         n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233,
         n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241,
         n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249,
         n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257,
         n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265,
         n39266, n39267, n39268, n39269, n39270, n39271, n39272, n39273,
         n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281,
         n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289,
         n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297,
         n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305,
         n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313,
         n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321,
         n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329,
         n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337,
         n39338, n39339, n39340, n39341, n39342, n39343, n39344, n39345,
         n39346, n39347, n39348, n39349, n39350, n39351, n39352, n39353,
         n39354, n39355, n39356, n39357, n39358, n39359, n39360, n39361,
         n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369,
         n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377,
         n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385,
         n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393,
         n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401,
         n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409,
         n39410, n39411, n39412, n39413, n39414, n39415, n39416, n39417,
         n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425,
         n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433,
         n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441,
         n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449,
         n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457,
         n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465,
         n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473,
         n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481,
         n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489,
         n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497,
         n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505,
         n39506, n39507, n39508, n39509, n39510, n39511, n39512, n39513,
         n39514, n39515, n39516, n39517, n39518, n39519, n39520, n39521,
         n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529,
         n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537,
         n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545,
         n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553,
         n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561,
         n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569,
         n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577,
         n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585,
         n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593,
         n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601,
         n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609,
         n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617,
         n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625,
         n39626, n39627, n39628, n39629, n39630, n39631, n39632, n39633,
         n39634, n39635, n39636, n39637, n39638, n39639, n39640, n39641,
         n39642, n39643, n39644, n39645, n39646, n39647, n39648, n39649,
         n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657,
         n39658, n39659, n39660, n39661, n39662, n39663, n39664, n39665,
         n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673,
         n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681,
         n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689,
         n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697,
         n39698, n39699, n39700, n39701, n39702, n39703, n39704, n39705,
         n39706, n39707, n39708, n39709, n39710, n39711, n39712, n39713,
         n39714, n39715, n39716, n39717, n39718, n39719, n39720, n39721,
         n39722, n39723, n39724, n39725, n39726, n39727, n39728, n39729,
         n39730, n39731, n39732, n39733, n39734, n39735, n39736, n39737,
         n39738, n39739, n39740, n39741, n39742, n39743, n39744, n39745,
         n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753,
         n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761,
         n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769,
         n39770, n39771, n39772, n39773, n39774, n39775, n39776, n39777,
         n39778, n39779, n39780, n39781, n39782, n39783, n39784, n39785,
         n39786, n39787, n39788, n39789, n39790, n39791, n39792, n39793,
         n39794, n39795, n39796, n39797, n39798, n39799, n39800, n39801,
         n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809,
         n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817,
         n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825,
         n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833,
         n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841,
         n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849,
         n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857,
         n39858, n39859, n39860, n39861, n39862, n39863, n39864, n39865,
         n39866, n39867, n39868, n39869, n39870, n39871, n39872, n39873,
         n39874, n39875, n39876, n39877, n39878, n39879, n39880, n39881,
         n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889,
         n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897,
         n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905,
         n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913,
         n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921,
         n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929,
         n39930, n39931, n39932, n39933, n39934, n39935, n39936, n39937,
         n39938, n39939, n39940, n39941, n39942, n39943, n39944, n39945,
         n39946, n39947, n39948, n39949, n39950, n39951, n39952, n39953,
         n39954, n39955, n39956, n39957, n39958, n39959, n39960, n39961,
         n39962, n39963, n39964, n39965, n39966, n39967, n39968, n39969,
         n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977,
         n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985,
         n39986, n39987, n39988, n39989, n39990, n39991, n39992, n39993,
         n39994, n39995, n39996, n39997, n39998, n39999, n40000, n40001,
         n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009,
         n40010, n40011, n40012, n40013, n40014, n40015, n40016, n40017,
         n40018, n40019, n40020, n40021, n40022, n40023, n40024, n40025,
         n40026, n40027, n40028, n40029, n40030, n40031, n40032, n40033,
         n40034, n40035, n40036, n40037, n40038, n40039, n40040, n40041,
         n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049,
         n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057,
         n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065,
         n40066, n40067, n40068, n40069, n40070, n40071, n40072, n40073,
         n40074, n40075, n40076, n40077, n40078, n40079, n40080, n40081,
         n40082, n40083, n40084, n40085, n40086, n40087, n40088, n40089,
         n40090, n40091, n40092, n40093, n40094, n40095, n40096, n40097,
         n40098, n40099, n40100, n40101, n40102, n40103, n40104, n40105,
         n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113,
         n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121,
         n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129,
         n40130, n40131, n40132, n40133, n40134, n40135, n40136, n40137,
         n40138, n40139, n40140, n40141, n40142, n40143, n40144, n40145,
         n40146, n40147, n40148, n40149, n40150, n40151, n40152, n40153,
         n40154, n40155, n40156, n40157, n40158, n40159, n40160, n40161,
         n40162, n40163, n40164, n40165, n40166, n40167, n40168, n40169,
         n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177,
         n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185,
         n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193,
         n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201,
         n40202, n40203, n40204, n40205, n40206, n40207, n40208, n40209,
         n40210, n40211, n40212, n40213, n40214, n40215, n40216, n40217,
         n40218, n40219, n40220, n40221, n40222, n40223, n40224, n40225,
         n40226, n40227, n40228, n40229, n40230, n40231, n40232, n40233,
         n40234, n40235, n40236, n40237, n40238, n40239, n40240, n40241,
         n40242, n40243, n40244, n40245, n40246, n40247, n40248, n40249,
         n40250, n40251, n40252, n40253, n40254, n40255, n40256, n40257,
         n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265,
         n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273,
         n40274, n40275, n40276, n40277, n40278, n40279, n40280, n40281,
         n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289,
         n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297,
         n40298, n40299, n40300, n40301, n40302, n40303, n40304, n40305,
         n40306, n40307, n40308, n40309, n40310, n40311, n40312, n40313,
         n40314, n40315, n40316, n40317, n40318, n40319, n40320, n40321,
         n40322, n40323, n40324, n40325, n40326, n40327, n40328, n40329,
         n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337,
         n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345,
         n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353,
         n40354, n40355, n40356, n40357, n40358, n40359, n40360, n40361,
         n40362, n40363, n40364, n40365, n40366, n40367, n40368, n40369,
         n40370, n40371, n40372, n40373, n40374, n40375, n40376, n40377,
         n40378, n40379, n40380, n40381, n40382, n40383, n40384, n40385,
         n40386, n40387, n40388, n40389, n40390, n40391, n40392, n40393,
         n40394, n40395, n40396, n40397, n40398, n40399, n40400, n40401,
         n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409,
         n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417,
         n40418, n40419, n40420, n40421, n40422, n40423, n40424, n40425,
         n40426, n40427, n40428, n40429, n40430, n40431, n40432, n40433,
         n40434, n40435, n40436, n40437, n40438, n40439, n40440, n40441,
         n40442, n40443, n40444, n40445, n40446, n40447, n40448, n40449,
         n40450, n40451, n40452, n40453, n40454, n40455, n40456, n40457,
         n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465,
         n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473,
         n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481,
         n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489,
         n40490, n40491, n40492, n40493, n40494, n40495, n40496, n40497,
         n40498, n40499, n40500, n40501, n40502, n40503, n40504, n40505,
         n40506, n40507, n40508, n40509, n40510, n40511, n40512, n40513,
         n40514, n40515, n40516, n40517, n40518, n40519, n40520, n40521,
         n40522, n40523, n40524, n40525, n40526, n40527, n40528, n40529,
         n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537,
         n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545,
         n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553,
         n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561,
         n40562, n40563, n40564, n40565, n40566, n40567, n40568, n40569,
         n40570, n40571, n40572, n40573, n40574, n40575, n40576, n40577,
         n40578, n40579, n40580, n40581, n40582, n40583, n40584, n40585,
         n40586, n40587, n40588, n40589, n40590, n40591, n40592, n40593,
         n40594, n40595, n40596, n40597, n40598, n40599, n40600, n40601,
         n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609,
         n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617,
         n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625,
         n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633,
         n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641,
         n40642, n40643, n40644, n40645, n40646, n40647, n40648, n40649,
         n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657,
         n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665,
         n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673,
         n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681,
         n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689,
         n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697,
         n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705,
         n40706, n40707, n40708, n40709, n40710, n40711, n40712, n40713,
         n40714, n40715, n40716, n40717, n40718, n40719, n40720, n40721,
         n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729,
         n40730, n40731, n40732, n40733, n40734, n40735, n40736, n40737,
         n40738, n40739, n40740, n40741, n40742, n40743, n40744, n40745,
         n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753,
         n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761,
         n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769,
         n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777,
         n40778, n40779, n40780, n40781, n40782, n40783, n40784, n40785,
         n40786, n40787, n40788, n40789, n40790, n40791, n40792, n40793,
         n40794, n40795, n40796, n40797, n40798, n40799, n40800, n40801,
         n40802, n40803, n40804, n40805, n40806, n40807, n40808, n40809,
         n40810, n40811, n40812, n40813, n40814, n40815, n40816, n40817,
         n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825,
         n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833,
         n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841,
         n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849,
         n40850, n40851, n40852, n40853, n40854, n40855, n40856, n40857,
         n40858, n40859, n40860, n40861, n40862, n40863, n40864, n40865,
         n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873,
         n40874, n40875, n40876, n40877, n40878, n40879, n40880, n40881,
         n40882, n40883, n40884, n40885, n40886, n40887, n40888, n40889,
         n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897,
         n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905,
         n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913,
         n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921,
         n40922, n40923, n40924, n40925, n40926, n40927, n40928, n40929,
         n40930, n40931, n40932, n40933, n40934, n40935, n40936, n40937,
         n40938, n40939, n40940, n40941, n40942, n40943, n40944, n40945,
         n40946, n40947, n40948, n40949, n40950, n40951, n40952, n40953,
         n40954, n40955, n40956, n40957, n40958, n40959, n40960, n40961,
         n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969,
         n40970, n40971, n40972, n40973, n40974, n40975, n40976, n40977,
         n40978, n40979, n40980, n40981, n40982, n40983, n40984, n40985,
         n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993,
         n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001,
         n41002, n41003, n41004, n41005, n41006, n41007, n41008, n41009,
         n41010, n41011, n41012, n41013, n41014, n41015, n41016, n41017,
         n41018, n41019, n41020, n41021, n41022, n41023, n41024, n41025,
         n41026, n41027, n41028, n41029, n41030, n41031, n41032, n41033,
         n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041,
         n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049,
         n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057,
         n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065,
         n41066, n41067, n41068, n41069, n41070, n41071, n41072, n41073,
         n41074, n41075, n41076, n41077, n41078, n41079, n41080, n41081,
         n41082, n41083, n41084, n41085, n41086, n41087, n41088, n41089,
         n41090, n41091, n41092, n41093, n41094, n41095, n41096, n41097,
         n41098, n41099, n41100, n41101, n41102, n41103, n41104, n41105,
         n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113,
         n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121,
         n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129,
         n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137,
         n41138, n41139, n41140, n41141, n41142, n41143, n41144, n41145,
         n41146, n41147, n41148, n41149, n41150, n41151, n41152, n41153,
         n41154, n41155, n41156, n41157, n41158, n41159, n41160, n41161,
         n41162, n41163, n41164, n41165, n41166, n41167, n41168, n41169,
         n41170, n41171, n41172, n41173, n41174, n41175, n41176, n41177,
         n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185,
         n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193,
         n41194, n41195, n41196, n41197, n41198, n41199, n41200, n41201,
         n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209,
         n41210, n41211, n41212, n41213, n41214, n41215, n41216, n41217,
         n41218, n41219, n41220, n41221, n41222, n41223, n41224, n41225,
         n41226, n41227, n41228, n41229, n41230, n41231, n41232, n41233,
         n41234, n41235, n41236, n41237, n41238, n41239, n41240, n41241,
         n41242, n41243, n41244, n41245, n41246, n41247, n41248, n41249,
         n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257,
         n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265,
         n41266, n41267, n41268, n41269, n41270, n41271, n41272, n41273,
         n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281,
         n41282, n41283, n41284, n41285, n41286, n41287, n41288, n41289,
         n41290, n41291, n41292, n41293, n41294, n41295, n41296, n41297,
         n41298, n41299, n41300, n41301, n41302, n41303, n41304, n41305,
         n41306, n41307, n41308, n41309, n41310, n41311, n41312, n41313,
         n41314, n41315, n41316, n41317, n41318, n41319, n41320, n41321,
         n41322, n41323, n41324, n41325, n41326, n41327, n41328, n41329,
         n41330, n41331, n41332, n41333, n41334, n41335, n41336, n41337,
         n41338, n41339, n41340, n41341, n41342, n41343, n41344, n41345,
         n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353,
         n41354, n41355, n41356, n41357, n41358, n41359, n41360, n41361,
         n41362, n41363, n41364, n41365, n41366, n41367, n41368, n41369,
         n41370, n41371, n41372, n41373, n41374, n41375, n41376, n41377,
         n41378, n41379, n41380, n41381, n41382, n41383, n41384, n41385,
         n41386, n41387, n41388, n41389, n41390, n41391, n41392, n41393,
         n41394, n41395, n41396, n41397, n41398, n41399, n41400, n41401,
         n41402, n41403, n41404, n41405, n41406, n41407, n41408, n41409,
         n41410, n41411, n41412, n41413, n41414, n41415, n41416, n41417,
         n41418, n41419, n41420, n41421, n41422, n41423, n41424, n41425,
         n41426, n41427, n41428, n41429, n41430, n41431, n41432, n41433,
         n41434, n41435, n41436, n41437, n41438, n41439, n41440, n41441,
         n41442, n41443, n41444, n41445, n41446, n41447, n41448, n41449,
         n41450, n41451, n41452, n41453, n41454, n41455, n41456, n41457,
         n41458, n41459, n41460, n41461, n41462, n41463, n41464, n41465,
         n41466, n41467, n41468, n41469, n41470, n41471, n41472, n41473,
         n41474, n41475, n41476, n41477, n41478, n41479, n41480, n41481,
         n41482, n41483, n41484, n41485, n41486, n41487, n41488, n41489,
         n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497,
         n41498, n41499, n41500, n41501, n41502, n41503, n41504, n41505,
         n41506, n41507, n41508, n41509, n41510, n41511, n41512, n41513,
         n41514, n41515, n41516, n41517, n41518, n41519, n41520, n41521,
         n41522, n41523, n41524, n41525, n41526, n41527, n41528, n41529,
         n41530, n41531, n41532, n41533, n41534, n41535, n41536, n41537,
         n41538, n41539, n41540, n41541, n41542, n41543, n41544, n41545,
         n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553,
         n41554, n41555, n41556, n41557, n41558, n41559, n41560, n41561,
         n41562, n41563, n41564, n41565, n41566, n41567, n41568, n41569,
         n41570, n41571, n41572, n41573, n41574, n41575, n41576, n41577,
         n41578, n41579, n41580, n41581, n41582, n41583, n41584, n41585,
         n41586, n41587, n41588, n41589, n41590, n41591, n41592, n41593,
         n41594, n41595, n41596, n41597, n41598, n41599, n41600, n41601,
         n41602, n41603, n41604, n41605, n41606, n41607, n41608, n41609,
         n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617,
         n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625,
         n41626, n41627, n41628, n41629, n41630, n41631, n41632, n41633,
         n41634, n41635, n41636, n41637, n41638, n41639, n41640, n41641,
         n41642, n41643, n41644, n41645, n41646, n41647, n41648, n41649,
         n41650, n41651, n41652, n41653, n41654, n41655, n41656, n41657,
         n41658, n41659, n41660, n41661, n41662, n41663, n41664, n41665,
         n41666, n41667, n41668, n41669, n41670, n41671, n41672, n41673,
         n41674, n41675, n41676, n41677, n41678, n41679, n41680, n41681,
         n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41689,
         n41690, n41691, n41692, n41693, n41694, n41695, n41696, n41697,
         n41698, n41699, n41700, n41701, n41702, n41703, n41704, n41705,
         n41706, n41707, n41708, n41709, n41710, n41711, n41712, n41713,
         n41714, n41715, n41716, n41717, n41718, n41719, n41720, n41721,
         n41722, n41723, n41724, n41725, n41726, n41727, n41728, n41729,
         n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737,
         n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745,
         n41746, n41747, n41748, n41749, n41750, n41751, n41752, n41753,
         n41754, n41755, n41756, n41757, n41758, n41759, n41760, n41761,
         n41762, n41763, n41764, n41765, n41766, n41767, n41768, n41769,
         n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777,
         n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785,
         n41786, n41787, n41788, n41789, n41790, n41791, n41792, n41793,
         n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801,
         n41802, n41803, n41804, n41805, n41806, n41807, n41808, n41809,
         n41810, n41811, n41812, n41813, n41814, n41815, n41816, n41817,
         n41818, n41819, n41820, n41821, n41822, n41823, n41824, n41825,
         n41826, n41827, n41828, n41829, n41830, n41831, n41832, n41833,
         n41834, n41835, n41836, n41837, n41838, n41839, n41840, n41841,
         n41842, n41843, n41844, n41845, n41846, n41847, n41848, n41849,
         n41850, n41851, n41852, n41853, n41854, n41855, n41856, n41857,
         n41858, n41859, n41860, n41861, n41862, n41863, n41864, n41865,
         n41866, n41867, n41868, n41869, n41870, n41871, n41872, n41873,
         n41874, n41875, n41876, n41877, n41878, n41879, n41880, n41881,
         n41882, n41883, n41884, n41885, n41886, n41887, n41888, n41889,
         n41890, n41891, n41892, n41893, n41894, n41895, n41896, n41897,
         n41898, n41899, n41900, n41901, n41902, n41903, n41904, n41905,
         n41906, n41907, n41908, n41909, n41910, n41911, n41912, n41913,
         n41914, n41915, n41916, n41917, n41918, n41919, n41920, n41921,
         n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929,
         n41930, n41931, n41932, n41933, n41934, n41935, n41936, n41937,
         n41938, n41939, n41940, n41941, n41942, n41943, n41944, n41945,
         n41946, n41947, n41948, n41949, n41950, n41951, n41952, n41953,
         n41954, n41955, n41956, n41957, n41958, n41959, n41960, n41961,
         n41962, n41963, n41964, n41965, n41966, n41967, n41968, n41969,
         n41970, n41971, n41972, n41973, n41974, n41975, n41976, n41977,
         n41978, n41979, n41980, n41981, n41982, n41983, n41984, n41985,
         n41986, n41987, n41988, n41989, n41990, n41991, n41992, n41993,
         n41994, n41995, n41996, n41997, n41998, n41999, n42000, n42001,
         n42002, n42003, n42004, n42005, n42006, n42007, n42008, n42009,
         n42010, n42011, n42012, n42013, n42014, n42015, n42016, n42017,
         n42018, n42019, n42020, n42021, n42022, n42023, n42024, n42025,
         n42026, n42027, n42028, n42029, n42030, n42031, n42032, n42033,
         n42034, n42035, n42036, n42037, n42038, n42039, n42040, n42041,
         n42042, n42043, n42044, n42045, n42046, n42047, n42048, n42049,
         n42050, n42051, n42052, n42053, n42054, n42055, n42056, n42057,
         n42058, n42059, n42060, n42061, n42062, n42063, n42064, n42065,
         n42066, n42067, n42068, n42069, n42070, n42071, n42072, n42073,
         n42074, n42075, n42076, n42077, n42078, n42079, n42080, n42081,
         n42082, n42083, n42084, n42085, n42086, n42087, n42088, n42089,
         n42090, n42091, n42092, n42093, n42094, n42095, n42096, n42097,
         n42098, n42099, n42100, n42101, n42102, n42103, n42104, n42105,
         n42106, n42107, n42108, n42109, n42110, n42111, n42112, n42113,
         n42114, n42115, n42116, n42117, n42118, n42119, n42120, n42121,
         n42122, n42123, n42124, n42125, n42126, n42127, n42128, n42129,
         n42130, n42131, n42132, n42133, n42134, n42135, n42136, n42137,
         n42138, n42139, n42140, n42141, n42142, n42143, n42144, n42145,
         n42146, n42147, n42148, n42149, n42150, n42151, n42152, n42153,
         n42154, n42155, n42156, n42157, n42158, n42159, n42160, n42161,
         n42162, n42163, n42164, n42165, n42166, n42167, n42168, n42169,
         n42170, n42171, n42172, n42173, n42174, n42175, n42176, n42177,
         n42178, n42179, n42180, n42181, n42182, n42183, n42184, n42185,
         n42186, n42187, n42188, n42189, n42190, n42191, n42192, n42193,
         n42194, n42195, n42196, n42197, n42198, n42199, n42200, n42201,
         n42202, n42203, n42204, n42205, n42206, n42207, n42208, n42209,
         n42210, n42211, n42212, n42213, n42214, n42215, n42216, n42217,
         n42218, n42219, n42220, n42221, n42222, n42223, n42224, n42225,
         n42226, n42227, n42228, n42229, n42230, n42231, n42232, n42233,
         n42234, n42235, n42236, n42237, n42238, n42239, n42240, n42241,
         n42242, n42243, n42244, n42245, n42246, n42247, n42248, n42249,
         n42250, n42251, n42252, n42253, n42254, n42255, n42256, n42257,
         n42258, n42259, n42260, n42261, n42262, n42263, n42264, n42265,
         n42266, n42267, n42268, n42269, n42270, n42271, n42272, n42273,
         n42274, n42275, n42276, n42277, n42278, n42279, n42280, n42281,
         n42282, n42283, n42284, n42285, n42286, n42287, n42288, n42289,
         n42290, n42291, n42292, n42293, n42294, n42295, n42296, n42297,
         n42298, n42299, n42300, n42301, n42302, n42303, n42304, n42305,
         n42306, n42307, n42308, n42309, n42310, n42311, n42312, n42313,
         n42314, n42315, n42316, n42317, n42318, n42319, n42320, n42321,
         n42322, n42323, n42324, n42325, n42326, n42327, n42328, n42329,
         n42330, n42331, n42332, n42333, n42334, n42335, n42336, n42337,
         n42338, n42339, n42340, n42341, n42342, n42343, n42344, n42345,
         n42346, n42347, n42348, n42349, n42350, n42351, n42352, n42353,
         n42354, n42355, n42356, n42357, n42358, n42359, n42360, n42361,
         n42362, n42363, n42364, n42365, n42366, n42367, n42368, n42369,
         n42370, n42371, n42372, n42373, n42374, n42375, n42376, n42377,
         n42378, n42379, n42380, n42381, n42382, n42383, n42384, n42385,
         n42386, n42387, n42388, n42389, n42390, n42391, n42392, n42393,
         n42394, n42395, n42396, n42397, n42398, n42399, n42400, n42401,
         n42402, n42403, n42404, n42405, n42406, n42407, n42408, n42409,
         n42410, n42411, n42412, n42413, n42414, n42415, n42416, n42417,
         n42418, n42419, n42420, n42421, n42422, n42423, n42424, n42425,
         n42426, n42427, n42428, n42429, n42430, n42431, n42432, n42433,
         n42434, n42435, n42436, n42437, n42438, n42439, n42440, n42441,
         n42442, n42443, n42444, n42445, n42446, n42447, n42448, n42449,
         n42450, n42451, n42452, n42453, n42454, n42455, n42456, n42457,
         n42458, n42459, n42460, n42461, n42462, n42463, n42464, n42465,
         n42466, n42467, n42468, n42469, n42470, n42471, n42472, n42473,
         n42474, n42475, n42476, n42477, n42478, n42479, n42480, n42481,
         n42482, n42483, n42484, n42485, n42486, n42487, n42488, n42489,
         n42490, n42491, n42492, n42493, n42494, n42495, n42496, n42497,
         n42498, n42499, n42500, n42501, n42502, n42503, n42504, n42505,
         n42506, n42507, n42508, n42509, n42510, n42511, n42512, n42513,
         n42514, n42515, n42516, n42517, n42518, n42519, n42520, n42521,
         n42522, n42523, n42524, n42525, n42526, n42527, n42528, n42529,
         n42530, n42531, n42532, n42533, n42534, n42535, n42536, n42537,
         n42538, n42539, n42540, n42541, n42542, n42543, n42544, n42545,
         n42546, n42547, n42548, n42549, n42550, n42551, n42552, n42553,
         n42554, n42555, n42556, n42557, n42558, n42559, n42560, n42561,
         n42562, n42563, n42564, n42565, n42566, n42567, n42568, n42569,
         n42570, n42571, n42572, n42573, n42574, n42575, n42576, n42577,
         n42578, n42579, n42580, n42581, n42582, n42583, n42584, n42585,
         n42586, n42587, n42588, n42589, n42590, n42591, n42592, n42593,
         n42594, n42595, n42596, n42597, n42598, n42599, n42600, n42601,
         n42602, n42603, n42604, n42605, n42606, n42607, n42608, n42609,
         n42610, n42611, n42612, n42613, n42614, n42615, n42616, n42617,
         n42618, n42619, n42620, n42621, n42622, n42623, n42624, n42625,
         n42626, n42627, n42628, n42629, n42630, n42631, n42632, n42633,
         n42634, n42635, n42636, n42637, n42638, n42639, n42640, n42641,
         n42642, n42643, n42644, n42645, n42646, n42647, n42648, n42649,
         n42650, n42651, n42652, n42653, n42654, n42655, n42656, n42657,
         n42658, n42659, n42660, n42661, n42662, n42663, n42664, n42665,
         n42666, n42667, n42668, n42669, n42670, n42671, n42672, n42673,
         n42674, n42675, n42676, n42677, n42678, n42679, n42680, n42681,
         n42682, n42683, n42684, n42685, n42686, n42687, n42688, n42689,
         n42690, n42691, n42692, n42693, n42694, n42695, n42696, n42697,
         n42698, n42699, n42700, n42701, n42702, n42703, n42704, n42705,
         n42706, n42707, n42708, n42709, n42710, n42711, n42712, n42713,
         n42714, n42715, n42716, n42717, n42718, n42719, n42720, n42721,
         n42722, n42723, n42724, n42725, n42726, n42727, n42728, n42729,
         n42730, n42731, n42732, n42733, n42734, n42735, n42736, n42737,
         n42738, n42739, n42740, n42741, n42742, n42743, n42744, n42745,
         n42746, n42747, n42748, n42749, n42750, n42751, n42752, n42753,
         n42754, n42755, n42756, n42757, n42758, n42759, n42760, n42761,
         n42762, n42763, n42764, n42765, n42766, n42767, n42768, n42769,
         n42770, n42771, n42772, n42773, n42774, n42775, n42776, n42777,
         n42778, n42779, n42780, n42781, n42782, n42783, n42784, n42785,
         n42786, n42787, n42788, n42789, n42790, n42791, n42792, n42793,
         n42794, n42795, n42796, n42797, n42798, n42799, n42800, n42801,
         n42802, n42803, n42804, n42805, n42806, n42807, n42808, n42809,
         n42810, n42811, n42812, n42813, n42814, n42815, n42816, n42817,
         n42818, n42819, n42820, n42821, n42822, n42823, n42824, n42825,
         n42826, n42827, n42828, n42829, n42830, n42831, n42832, n42833,
         n42834, n42835, n42836, n42837, n42838, n42839, n42840, n42841,
         n42842, n42843, n42844, n42845, n42846, n42847, n42848, n42849,
         n42850, n42851, n42852, n42853, n42854, n42855, n42856, n42857,
         n42858, n42859, n42860, n42861, n42862, n42863, n42864, n42865,
         n42866, n42867, n42868, n42869, n42870, n42871, n42872, n42873,
         n42874, n42875, n42876, n42877, n42878, n42879, n42880, n42881,
         n42882, n42883, n42884, n42885, n42886, n42887, n42888, n42889,
         n42890, n42891, n42892, n42893, n42894, n42895, n42896, n42897,
         n42898, n42899, n42900, n42901, n42902, n42903, n42904, n42905,
         n42906, n42907, n42908, n42909, n42910, n42911, n42912, n42913,
         n42914, n42915, n42916, n42917, n42918, n42919, n42920, n42921,
         n42922, n42923, n42924, n42925, n42926, n42927, n42928, n42929,
         n42930, n42931, n42932, n42933, n42934, n42935, n42936, n42937,
         n42938, n42939, n42940, n42941, n42942, n42943, n42944, n42945,
         n42946, n42947, n42948, n42949, n42950, n42951, n42952, n42953,
         n42954, n42955, n42956, n42957, n42958, n42959, n42960, n42961,
         n42962, n42963, n42964, n42965, n42966, n42967, n42968, n42969,
         n42970, n42971, n42972, n42973, n42974, n42975, n42976, n42977,
         n42978, n42979, n42980, n42981, n42982, n42983, n42984, n42985,
         n42986, n42987, n42988, n42989, n42990, n42991, n42992, n42993,
         n42994, n42995, n42996, n42997, n42998, n42999, n43000, n43001,
         n43002, n43003, n43004, n43005, n43006, n43007, n43008, n43009,
         n43010, n43011, n43012, n43013, n43014, n43015, n43016, n43017,
         n43018, n43019, n43020, n43021, n43022, n43023, n43024, n43025,
         n43026, n43027, n43028, n43029, n43030, n43031, n43032, n43033,
         n43034, n43035, n43036, n43037, n43038, n43039, n43040, n43041,
         n43042, n43043, n43044, n43045, n43046, n43047, n43048, n43049,
         n43050, n43051, n43052, n43053, n43054, n43055, n43056, n43057,
         n43058, n43059, n43060, n43061, n43062, n43063, n43064, n43065,
         n43066, n43067, n43068, n43069, n43070, n43071, n43072, n43073,
         n43074, n43075, n43076, n43077, n43078, n43079, n43080, n43081,
         n43082, n43083, n43084, n43085, n43086, n43087, n43088, n43089,
         n43090, n43091, n43092, n43093, n43094, n43095, n43096, n43097,
         n43098, n43099, n43100, n43101, n43102, n43103, n43104, n43105,
         n43106, n43107, n43108, n43109, n43110, n43111, n43112, n43113,
         n43114, n43115, n43116, n43117, n43118, n43119, n43120, n43121,
         n43122, n43123, n43124, n43125, n43126, n43127, n43128, n43129,
         n43130, n43131, n43132, n43133, n43134, n43135, n43136, n43137,
         n43138, n43139, n43140, n43141, n43142, n43143, n43144, n43145,
         n43146, n43147, n43148, n43149, n43150, n43151, n43152, n43153,
         n43154, n43155, n43156, n43157, n43158, n43159, n43160, n43161,
         n43162, n43163, n43164, n43165, n43166, n43167, n43168, n43169,
         n43170, n43171, n43172, n43173, n43174, n43175, n43176, n43177,
         n43178, n43179, n43180, n43181, n43182, n43183, n43184, n43185,
         n43186, n43187, n43188, n43189, n43190, n43191, n43192, n43193,
         n43194, n43195, n43196, n43197, n43198, n43199, n43200, n43201,
         n43202, n43203, n43204, n43205, n43206, n43207, n43208, n43209,
         n43210, n43211, n43212, n43213, n43214, n43215, n43216, n43217,
         n43218, n43219, n43220, n43221, n43222, n43223, n43224, n43225,
         n43226, n43227, n43228, n43229, n43230, n43231, n43232, n43233,
         n43234, n43235, n43236, n43237, n43238, n43239, n43240, n43241,
         n43242, n43243, n43244, n43245, n43246, n43247, n43248, n43249,
         n43250, n43251, n43252, n43253, n43254, n43255, n43256, n43257,
         n43258, n43259, n43260, n43261, n43262, n43263, n43264, n43265,
         n43266, n43267, n43268, n43269, n43270, n43271, n43272, n43273,
         n43274, n43275, n43276, n43277, n43278, n43279, n43280, n43281,
         n43282, n43283, n43284, n43285, n43286, n43287, n43288, n43289,
         n43290, n43291, n43292, n43293, n43294, n43295, n43296, n43297,
         n43298, n43299, n43300, n43301, n43302, n43303, n43304, n43305,
         n43306, n43307, n43308, n43309, n43310, n43311, n43312, n43313,
         n43314, n43315, n43316, n43317, n43318, n43319, n43320, n43321,
         n43322, n43323, n43324, n43325, n43326, n43327, n43328, n43329,
         n43330, n43331, n43332, n43333, n43334, n43335, n43336, n43337,
         n43338, n43339, n43340, n43341, n43342, n43343, n43344, n43345,
         n43346, n43347, n43348, n43349, n43350, n43351, n43352, n43353,
         n43354, n43355, n43356, n43357, n43358, n43359, n43360, n43361,
         n43362, n43363, n43364, n43365, n43366, n43367, n43368, n43369,
         n43370, n43371, n43372, n43373, n43374, n43375, n43376, n43377,
         n43378, n43379, n43380, n43381, n43382, n43383, n43384, n43385,
         n43386, n43387, n43388, n43389, n43390, n43391, n43392, n43393,
         n43394, n43395, n43396, n43397, n43398, n43399, n43400, n43401,
         n43402, n43403, n43404, n43405, n43406, n43407, n43408, n43409,
         n43410, n43411, n43412, n43413, n43414, n43415, n43416, n43417,
         n43418, n43419, n43420, n43421, n43422, n43423, n43424, n43425,
         n43426, n43427, n43428, n43429, n43430, n43431, n43432, n43433,
         n43434, n43435, n43436, n43437, n43438, n43439, n43440, n43441,
         n43442, n43443, n43444, n43445, n43446, n43447, n43448, n43449,
         n43450, n43451, n43452, n43453, n43454, n43455, n43456, n43457,
         n43458, n43459, n43460, n43461, n43462, n43463, n43464, n43465,
         n43466, n43467, n43468, n43469, n43470, n43471, n43472, n43473,
         n43474, n43475, n43476, n43477, n43478, n43479, n43480, n43481,
         n43482, n43483, n43484, n43485, n43486, n43487, n43488, n43489,
         n43490, n43491, n43492, n43493, n43494, n43495, n43496, n43497,
         n43498, n43499, n43500, n43501, n43502, n43503, n43504, n43505,
         n43506, n43507, n43508, n43509, n43510, n43511, n43512, n43513,
         n43514, n43515, n43516, n43517, n43518, n43519, n43520, n43521,
         n43522, n43523, n43524, n43525, n43526, n43527, n43528, n43529,
         n43530, n43531, n43532, n43533, n43534, n43535, n43536, n43537,
         n43538, n43539, n43540, n43541, n43542, n43543, n43544, n43545,
         n43546, n43547, n43548, n43549, n43550, n43551, n43552, n43553,
         n43554, n43555, n43556, n43557, n43558, n43559, n43560, n43561,
         n43562, n43563, n43564, n43565, n43566, n43567, n43568, n43569,
         n43570, n43571, n43572, n43573, n43574, n43575, n43576, n43577,
         n43578, n43579, n43580, n43581, n43582, n43583, n43584, n43585,
         n43586, n43587, n43588, n43589, n43590, n43591, n43592, n43593,
         n43594, n43595, n43596, n43597, n43598, n43599, n43600, n43601,
         n43602, n43603, n43604, n43605, n43606, n43607, n43608, n43609,
         n43610, n43611, n43612, n43613, n43614, n43615, n43616, n43617,
         n43618, n43619, n43620, n43621, n43622, n43623, n43624, n43625,
         n43626, n43627, n43628, n43629, n43630, n43631, n43632, n43633,
         n43634, n43635, n43636, n43637, n43638, n43639, n43640, n43641,
         n43642, n43643, n43644, n43645, n43646, n43647, n43648, n43649,
         n43650, n43651, n43652, n43653, n43654, n43655, n43656, n43657,
         n43658, n43659, n43660, n43661, n43662, n43663, n43664, n43665,
         n43666, n43667, n43668, n43669, n43670, n43671, n43672, n43673,
         n43674, n43675, n43676, n43677, n43678, n43679, n43680, n43681,
         n43682, n43683, n43684, n43685, n43686, n43687, n43688, n43689,
         n43690, n43691, n43692, n43693, n43694, n43695, n43696, n43697,
         n43698, n43699, n43700, n43701, n43702, n43703, n43704, n43705,
         n43706, n43707, n43708, n43709, n43710, n43711, n43712, n43713,
         n43714, n43715, n43716, n43717, n43718, n43719, n43720, n43721,
         n43722, n43723, n43724, n43725, n43726, n43727, n43728, n43729,
         n43730, n43731, n43732, n43733, n43734, n43735, n43736, n43737,
         n43738, n43739, n43740, n43741, n43742, n43743, n43744, n43745,
         n43746, n43747, n43748, n43749, n43750, n43751, n43752, n43753,
         n43754, n43755, n43756, n43757, n43758, n43759, n43760, n43761,
         n43762, n43763, n43764, n43765, n43766, n43767, n43768, n43769,
         n43770, n43771, n43772, n43773, n43774, n43775, n43776, n43777,
         n43778, n43779, n43780, n43781, n43782, n43783, n43784, n43785,
         n43786, n43787, n43788, n43789, n43790, n43791, n43792, n43793,
         n43794, n43795, n43796, n43797, n43798, n43799, n43800, n43801,
         n43802, n43803, n43804, n43805, n43806, n43807, n43808, n43809,
         n43810, n43811, n43812, n43813, n43814, n43815, n43816, n43817,
         n43818, n43819, n43820, n43821, n43822, n43823, n43824, n43825,
         n43826, n43827, n43828, n43829, n43830, n43831, n43832, n43833,
         n43834, n43835, n43836, n43837, n43838, n43839, n43840, n43841,
         n43842, n43843, n43844, n43845, n43846, n43847, n43848, n43849,
         n43850, n43851, n43852, n43853, n43854, n43855, n43856, n43857,
         n43858, n43859, n43860, n43861, n43862, n43863, n43864, n43865,
         n43866, n43867, n43868, n43869, n43870, n43871, n43872, n43873,
         n43874, n43875, n43876, n43877, n43878, n43879, n43880, n43881,
         n43882, n43883, n43884, n43885, n43886, n43887, n43888, n43889,
         n43890, n43891, n43892, n43893, n43894, n43895, n43896, n43897,
         n43898, n43899, n43900, n43901, n43902, n43903, n43904, n43905,
         n43906, n43907, n43908, n43909, n43910, n43911, n43912, n43913,
         n43914, n43915, n43916, n43917, n43918, n43919, n43920, n43921,
         n43922, n43923, n43924, n43925, n43926, n43927, n43928, n43929,
         n43930, n43931, n43932, n43933, n43934, n43935, n43936, n43937,
         n43938, n43939, n43940, n43941, n43942, n43943, n43944, n43945,
         n43946, n43947, n43948, n43949, n43950, n43951, n43952, n43953,
         n43954, n43955, n43956, n43957, n43958, n43959, n43960, n43961,
         n43962, n43963, n43964, n43965, n43966, n43967, n43968, n43969,
         n43970, n43971, n43972, n43973, n43974, n43975, n43976, n43977,
         n43978, n43979, n43980, n43981, n43982, n43983, n43984, n43985,
         n43986, n43987, n43988, n43989, n43990, n43991, n43992, n43993,
         n43994, n43995, n43996, n43997, n43998, n43999, n44000, n44001,
         n44002, n44003, n44004, n44005, n44006, n44007, n44008, n44009,
         n44010, n44011, n44012, n44013, n44014, n44015, n44016, n44017,
         n44018, n44019, n44020, n44021, n44022, n44023, n44024, n44025,
         n44026, n44027, n44028, n44029, n44030, n44031, n44032, n44033,
         n44034, n44035, n44036, n44037, n44038, n44039, n44040, n44041,
         n44042, n44043, n44044, n44045, n44046, n44047, n44048, n44049,
         n44050, n44051, n44052, n44053, n44054, n44055, n44056, n44057,
         n44058, n44059, n44060, n44061, n44062, n44063, n44064, n44065,
         n44066, n44067, n44068, n44069, n44070, n44071, n44072, n44073,
         n44074, n44075, n44076, n44077, n44078, n44079, n44080, n44081,
         n44082, n44083, n44084, n44085, n44086, n44087, n44088, n44089,
         n44090, n44091, n44092, n44093, n44094, n44095, n44096, n44097,
         n44098, n44099, n44100, n44101, n44102, n44103, n44104, n44105,
         n44106, n44107, n44108, n44109, n44110, n44111, n44112, n44113,
         n44114, n44115, n44116, n44117, n44118, n44119, n44120, n44121,
         n44122, n44123, n44124, n44125, n44126, n44127, n44128, n44129,
         n44130, n44131, n44132, n44133, n44134, n44135, n44136, n44137,
         n44138, n44139, n44140, n44141, n44142, n44143, n44144, n44145,
         n44146, n44147, n44148, n44149, n44150, n44151, n44152, n44153,
         n44154, n44155, n44156, n44157, n44158, n44159, n44160, n44161,
         n44162, n44163, n44164, n44165, n44166, n44167, n44168, n44169,
         n44170, n44171, n44172, n44173, n44174, n44175, n44176, n44177,
         n44178, n44179, n44180, n44181, n44182, n44183, n44184, n44185,
         n44186, n44187, n44188, n44189, n44190, n44191, n44192, n44193,
         n44194, n44195, n44196, n44197, n44198, n44199, n44200, n44201,
         n44202, n44203, n44204, n44205, n44206, n44207, n44208, n44209,
         n44210, n44211, n44212, n44213, n44214, n44215, n44216, n44217,
         n44218, n44219, n44220, n44221, n44222, n44223, n44224, n44225,
         n44226, n44227, n44228, n44229, n44230, n44231, n44232, n44233,
         n44234, n44235, n44236, n44237, n44238, n44239, n44240, n44241,
         n44242, n44243, n44244, n44245, n44246, n44247, n44248, n44249,
         n44250, n44251, n44252, n44253, n44254, n44255, n44256, n44257,
         n44258, n44259, n44260, n44261, n44262, n44263, n44264, n44265,
         n44266, n44267, n44268, n44269, n44270, n44271, n44272, n44273,
         n44274, n44275, n44276, n44277, n44278, n44279, n44280, n44281,
         n44282, n44283, n44284, n44285, n44286, n44287, n44288, n44289,
         n44290, n44291, n44292, n44293, n44294, n44295, n44296, n44297,
         n44298, n44299, n44300, n44301, n44302, n44303, n44304, n44305,
         n44306, n44307, n44308, n44309, n44310, n44311, n44312, n44313,
         n44314, n44315, n44316, n44317, n44318, n44319, n44320, n44321,
         n44322, n44323, n44324, n44325, n44326, n44327, n44328, n44329,
         n44330, n44331, n44332, n44333, n44334, n44335, n44336, n44337,
         n44338, n44339, n44340, n44341, n44342, n44343, n44344, n44345,
         n44346, n44347, n44348, n44349, n44350, n44351, n44352, n44353,
         n44354, n44355, n44356, n44357, n44358, n44359, n44360, n44361,
         n44362, n44363, n44364, n44365, n44366, n44367, n44368, n44369,
         n44370, n44371, n44372, n44373, n44374, n44375, n44376, n44377,
         n44378, n44379, n44380, n44381, n44382, n44383, n44384, n44385,
         n44386, n44387, n44388, n44389, n44390, n44391, n44392, n44393,
         n44394, n44395, n44396, n44397, n44398, n44399, n44400, n44401,
         n44402, n44403, n44404, n44405, n44406, n44407, n44408, n44409,
         n44410, n44411, n44412, n44413, n44414, n44415, n44416, n44417,
         n44418, n44419, n44420, n44421, n44422, n44423, n44424, n44425,
         n44426, n44427, n44428, n44429, n44430, n44431, n44432, n44433,
         n44434, n44435, n44436, n44437, n44438, n44439, n44440, n44441,
         n44442, n44443, n44444, n44445, n44446, n44447, n44448, n44449,
         n44450, n44451, n44452, n44453, n44454, n44455, n44456, n44457,
         n44458, n44459, n44460, n44461, n44462, n44463, n44464, n44465,
         n44466, n44467, n44468, n44469, n44470, n44471, n44472, n44473,
         n44474, n44475, n44476, n44477, n44478, n44479, n44480, n44481,
         n44482, n44483, n44484, n44485, n44486, n44487, n44488, n44489,
         n44490, n44491, n44492, n44493, n44494, n44495, n44496, n44497,
         n44498, n44499, n44500, n44501, n44502, n44503, n44504, n44505,
         n44506, n44507, n44508, n44509, n44510, n44511, n44512, n44513,
         n44514, n44515, n44516, n44517, n44518, n44519, n44520, n44521,
         n44522, n44523, n44524, n44525, n44526, n44527, n44528, n44529,
         n44530, n44531, n44532, n44533, n44534, n44535, n44536, n44537,
         n44538, n44539, n44540, n44541, n44542, n44543, n44544, n44545,
         n44546, n44547, n44548, n44549, n44550, n44551, n44552, n44553,
         n44554, n44555, n44556, n44557, n44558, n44559, n44560, n44561,
         n44562, n44563, n44564, n44565, n44566, n44567, n44568, n44569,
         n44570, n44571, n44572, n44573, n44574, n44575, n44576, n44577,
         n44578, n44579, n44580, n44581, n44582, n44583, n44584, n44585,
         n44586, n44587, n44588, n44589, n44590, n44591, n44592, n44593,
         n44594, n44595, n44596, n44597, n44598, n44599, n44600, n44601,
         n44602, n44603, n44604, n44605, n44606, n44607, n44608, n44609,
         n44610, n44611, n44612, n44613, n44614, n44615, n44616, n44617,
         n44618, n44619, n44620, n44621, n44622, n44623, n44624, n44625,
         n44626, n44627, n44628, n44629, n44630, n44631, n44632, n44633,
         n44634, n44635, n44636, n44637, n44638, n44639, n44640, n44641,
         n44642, n44643, n44644, n44645, n44646, n44647, n44648, n44649,
         n44650, n44651, n44652, n44653, n44654, n44655, n44656, n44657,
         n44658, n44659, n44660, n44661, n44662, n44663, n44664, n44665,
         n44666, n44667, n44668, n44669, n44670, n44671, n44672, n44673,
         n44674, n44675, n44676, n44677, n44678, n44679, n44680, n44681,
         n44682, n44683, n44684, n44685, n44686, n44687, n44688, n44689,
         n44690, n44691, n44692, n44693, n44694, n44695, n44696, n44697,
         n44698, n44699, n44700, n44701, n44702, n44703, n44704, n44705,
         n44706, n44707, n44708, n44709, n44710;

  XOR U2 ( .A(n1), .B(n2), .Z(o[0]) );
  AND U3 ( .A(o[1]), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(n5), .Z(n3) );
  IV U5 ( .A(n1), .Z(n5) );
  XNOR U6 ( .A(n6), .B(n7), .Z(o[1]) );
  AND U7 ( .A(n8), .B(n9), .Z(n7) );
  XOR U8 ( .A(n6), .B(n10), .Z(n9) );
  XOR U9 ( .A(n11), .B(n12), .Z(n10) );
  AND U10 ( .A(n4), .B(n13), .Z(n11) );
  XNOR U11 ( .A(n14), .B(n12), .Z(n13) );
  XOR U12 ( .A(n15), .B(n6), .Z(n8) );
  XOR U13 ( .A(n16), .B(n17), .Z(n15) );
  AND U14 ( .A(n1), .B(n18), .Z(n17) );
  XNOR U15 ( .A(n19), .B(n20), .Z(n18) );
  XOR U16 ( .A(n21), .B(n22), .Z(n6) );
  AND U17 ( .A(n23), .B(n24), .Z(n22) );
  XOR U18 ( .A(n21), .B(n25), .Z(n24) );
  XNOR U19 ( .A(n26), .B(n27), .Z(n25) );
  AND U20 ( .A(n4), .B(n28), .Z(n26) );
  XNOR U21 ( .A(n29), .B(n27), .Z(n28) );
  XOR U22 ( .A(n30), .B(n21), .Z(n23) );
  XOR U23 ( .A(n31), .B(n32), .Z(n30) );
  AND U24 ( .A(n1), .B(n33), .Z(n32) );
  XOR U25 ( .A(n34), .B(n35), .Z(n33) );
  XOR U26 ( .A(n36), .B(n37), .Z(n21) );
  AND U27 ( .A(n38), .B(n39), .Z(n37) );
  XOR U28 ( .A(n36), .B(n40), .Z(n39) );
  XNOR U29 ( .A(n41), .B(n42), .Z(n40) );
  AND U30 ( .A(n4), .B(n43), .Z(n41) );
  XNOR U31 ( .A(n44), .B(n45), .Z(n43) );
  XOR U32 ( .A(n46), .B(n36), .Z(n38) );
  XNOR U33 ( .A(n47), .B(n48), .Z(n46) );
  AND U34 ( .A(n1), .B(n49), .Z(n48) );
  XNOR U35 ( .A(n50), .B(n47), .Z(n49) );
  XOR U36 ( .A(n51), .B(n52), .Z(n36) );
  AND U37 ( .A(n53), .B(n54), .Z(n52) );
  XOR U38 ( .A(n55), .B(n51), .Z(n54) );
  XNOR U39 ( .A(n56), .B(n57), .Z(n55) );
  AND U40 ( .A(n4), .B(n58), .Z(n57) );
  XOR U41 ( .A(n59), .B(n60), .Z(n58) );
  XOR U42 ( .A(n51), .B(n61), .Z(n53) );
  XNOR U43 ( .A(n62), .B(n63), .Z(n61) );
  AND U44 ( .A(n1), .B(n64), .Z(n62) );
  XOR U45 ( .A(n63), .B(n65), .Z(n64) );
  XOR U46 ( .A(n66), .B(n67), .Z(n51) );
  AND U47 ( .A(n68), .B(n69), .Z(n67) );
  XOR U48 ( .A(n66), .B(n70), .Z(n69) );
  XNOR U49 ( .A(n71), .B(n72), .Z(n70) );
  AND U50 ( .A(n4), .B(n73), .Z(n71) );
  XNOR U51 ( .A(n74), .B(n72), .Z(n73) );
  XOR U52 ( .A(n75), .B(n66), .Z(n68) );
  XOR U53 ( .A(n76), .B(n77), .Z(n75) );
  AND U54 ( .A(n1), .B(n78), .Z(n77) );
  XOR U55 ( .A(n79), .B(n80), .Z(n78) );
  IV U56 ( .A(n76), .Z(n80) );
  XOR U57 ( .A(n81), .B(n82), .Z(n66) );
  AND U58 ( .A(n83), .B(n84), .Z(n82) );
  XOR U59 ( .A(n81), .B(n85), .Z(n84) );
  XNOR U60 ( .A(n86), .B(n87), .Z(n85) );
  AND U61 ( .A(n4), .B(n88), .Z(n86) );
  XNOR U62 ( .A(n89), .B(n87), .Z(n88) );
  XOR U63 ( .A(n90), .B(n81), .Z(n83) );
  XOR U64 ( .A(n91), .B(n92), .Z(n90) );
  AND U65 ( .A(n1), .B(n93), .Z(n92) );
  XOR U66 ( .A(n94), .B(n95), .Z(n93) );
  IV U67 ( .A(n91), .Z(n95) );
  XOR U68 ( .A(n96), .B(n97), .Z(n81) );
  AND U69 ( .A(n98), .B(n99), .Z(n97) );
  XOR U70 ( .A(n96), .B(n100), .Z(n99) );
  XNOR U71 ( .A(n101), .B(n102), .Z(n100) );
  AND U72 ( .A(n4), .B(n103), .Z(n101) );
  XNOR U73 ( .A(n104), .B(n102), .Z(n103) );
  XOR U74 ( .A(n105), .B(n96), .Z(n98) );
  XOR U75 ( .A(n106), .B(n107), .Z(n105) );
  AND U76 ( .A(n1), .B(n108), .Z(n107) );
  XOR U77 ( .A(n109), .B(n110), .Z(n108) );
  IV U78 ( .A(n106), .Z(n110) );
  XOR U79 ( .A(n111), .B(n112), .Z(n96) );
  AND U80 ( .A(n113), .B(n114), .Z(n112) );
  XOR U81 ( .A(n111), .B(n115), .Z(n114) );
  XNOR U82 ( .A(n116), .B(n117), .Z(n115) );
  AND U83 ( .A(n4), .B(n118), .Z(n116) );
  XNOR U84 ( .A(n119), .B(n117), .Z(n118) );
  XOR U85 ( .A(n120), .B(n111), .Z(n113) );
  XOR U86 ( .A(n121), .B(n122), .Z(n120) );
  AND U87 ( .A(n1), .B(n123), .Z(n122) );
  XOR U88 ( .A(n124), .B(n125), .Z(n123) );
  IV U89 ( .A(n121), .Z(n125) );
  XOR U90 ( .A(n126), .B(n127), .Z(n111) );
  AND U91 ( .A(n128), .B(n129), .Z(n127) );
  XOR U92 ( .A(n130), .B(n131), .Z(n129) );
  XOR U93 ( .A(n126), .B(n132), .Z(n131) );
  AND U94 ( .A(n4), .B(n133), .Z(n132) );
  XOR U95 ( .A(n130), .B(n134), .Z(n133) );
  XNOR U96 ( .A(n135), .B(n136), .Z(n128) );
  XOR U97 ( .A(n126), .B(n137), .Z(n136) );
  AND U98 ( .A(n1), .B(n138), .Z(n137) );
  XOR U99 ( .A(n139), .B(n135), .Z(n138) );
  AND U100 ( .A(n140), .B(n141), .Z(n126) );
  XNOR U101 ( .A(n142), .B(n143), .Z(n141) );
  AND U102 ( .A(n4), .B(n144), .Z(n142) );
  XNOR U103 ( .A(n145), .B(n143), .Z(n144) );
  XNOR U104 ( .A(n146), .B(n147), .Z(n4) );
  AND U105 ( .A(n148), .B(n149), .Z(n147) );
  XNOR U106 ( .A(n146), .B(n14), .Z(n149) );
  XNOR U107 ( .A(n150), .B(n151), .Z(n14) );
  AND U108 ( .A(n152), .B(n153), .Z(n151) );
  XOR U109 ( .A(n29), .B(n150), .Z(n152) );
  XOR U110 ( .A(n154), .B(n155), .Z(n150) );
  AND U111 ( .A(n29), .B(n154), .Z(n155) );
  XNOR U112 ( .A(n12), .B(n146), .Z(n148) );
  XOR U113 ( .A(n156), .B(n157), .Z(n12) );
  AND U114 ( .A(n158), .B(n159), .Z(n157) );
  XOR U115 ( .A(n160), .B(n156), .Z(n158) );
  XOR U116 ( .A(n161), .B(n162), .Z(n156) );
  NOR U117 ( .A(n27), .B(n163), .Z(n162) );
  IV U118 ( .A(n161), .Z(n163) );
  IV U119 ( .A(n160), .Z(n27) );
  XOR U120 ( .A(n164), .B(n165), .Z(n146) );
  AND U121 ( .A(n166), .B(n167), .Z(n165) );
  XOR U122 ( .A(n164), .B(n29), .Z(n167) );
  XOR U123 ( .A(n154), .B(n153), .Z(n29) );
  XNOR U124 ( .A(n168), .B(n169), .Z(n153) );
  XOR U125 ( .A(n170), .B(n171), .Z(n169) );
  XOR U126 ( .A(n172), .B(n173), .Z(n171) );
  NOR U127 ( .A(n174), .B(n175), .Z(n172) );
  XOR U128 ( .A(n176), .B(n177), .Z(n170) );
  NOR U129 ( .A(n178), .B(n179), .Z(n177) );
  NOR U130 ( .A(n180), .B(n181), .Z(n176) );
  XOR U131 ( .A(n182), .B(n183), .Z(n168) );
  XOR U132 ( .A(n175), .B(n179), .Z(n183) );
  XNOR U133 ( .A(n184), .B(n181), .Z(n182) );
  XOR U134 ( .A(n185), .B(n186), .Z(n184) );
  XOR U135 ( .A(n187), .B(n188), .Z(n186) );
  XOR U136 ( .A(n189), .B(n190), .Z(n188) );
  XOR U137 ( .A(n191), .B(n192), .Z(n187) );
  NOR U138 ( .A(n193), .B(n194), .Z(n192) );
  AND U139 ( .A(n195), .B(n173), .Z(n191) );
  XOR U140 ( .A(n196), .B(n197), .Z(n185) );
  XOR U141 ( .A(n198), .B(n199), .Z(n197) );
  XOR U142 ( .A(n200), .B(n201), .Z(n199) );
  XOR U143 ( .A(n202), .B(n203), .Z(n201) );
  XOR U144 ( .A(n204), .B(n205), .Z(n203) );
  XOR U145 ( .A(n206), .B(n207), .Z(n205) );
  XNOR U146 ( .A(n208), .B(n209), .Z(n204) );
  XNOR U147 ( .A(n210), .B(n211), .Z(n209) );
  NOR U148 ( .A(n212), .B(n207), .Z(n210) );
  XOR U149 ( .A(n213), .B(n214), .Z(n202) );
  XOR U150 ( .A(n215), .B(n216), .Z(n214) );
  XNOR U151 ( .A(n217), .B(n218), .Z(n216) );
  XOR U152 ( .A(n219), .B(n220), .Z(n218) );
  XOR U153 ( .A(n221), .B(n222), .Z(n220) );
  XOR U154 ( .A(n223), .B(n224), .Z(n222) );
  XOR U155 ( .A(n225), .B(n226), .Z(n221) );
  XOR U156 ( .A(n227), .B(n228), .Z(n226) );
  XOR U157 ( .A(n229), .B(n230), .Z(n228) );
  XOR U158 ( .A(n231), .B(n232), .Z(n230) );
  XOR U159 ( .A(n233), .B(n234), .Z(n232) );
  XNOR U160 ( .A(n235), .B(n236), .Z(n231) );
  XNOR U161 ( .A(n237), .B(n238), .Z(n236) );
  NOR U162 ( .A(n239), .B(n234), .Z(n237) );
  XOR U163 ( .A(n240), .B(n241), .Z(n229) );
  XOR U164 ( .A(n242), .B(n243), .Z(n241) );
  XNOR U165 ( .A(n244), .B(n245), .Z(n243) );
  XOR U166 ( .A(n246), .B(n247), .Z(n245) );
  XOR U167 ( .A(n248), .B(n249), .Z(n247) );
  XOR U168 ( .A(n250), .B(n251), .Z(n249) );
  XOR U169 ( .A(n252), .B(n253), .Z(n248) );
  XOR U170 ( .A(n254), .B(n255), .Z(n253) );
  XOR U171 ( .A(n256), .B(n257), .Z(n255) );
  XOR U172 ( .A(n258), .B(n259), .Z(n257) );
  XOR U173 ( .A(n260), .B(n261), .Z(n259) );
  XNOR U174 ( .A(n262), .B(n263), .Z(n258) );
  XNOR U175 ( .A(n264), .B(n265), .Z(n263) );
  NOR U176 ( .A(n266), .B(n261), .Z(n264) );
  XOR U177 ( .A(n267), .B(n268), .Z(n256) );
  XOR U178 ( .A(n269), .B(n270), .Z(n268) );
  XNOR U179 ( .A(n271), .B(n272), .Z(n270) );
  XOR U180 ( .A(n273), .B(n274), .Z(n272) );
  XOR U181 ( .A(n275), .B(n276), .Z(n274) );
  XOR U182 ( .A(n277), .B(n278), .Z(n276) );
  XOR U183 ( .A(n279), .B(n280), .Z(n275) );
  XOR U184 ( .A(n281), .B(n282), .Z(n280) );
  XOR U185 ( .A(n283), .B(n284), .Z(n282) );
  XOR U186 ( .A(n285), .B(n286), .Z(n284) );
  XOR U187 ( .A(n287), .B(n288), .Z(n286) );
  XNOR U188 ( .A(n289), .B(n290), .Z(n285) );
  XNOR U189 ( .A(n291), .B(n292), .Z(n290) );
  NOR U190 ( .A(n293), .B(n288), .Z(n291) );
  XOR U191 ( .A(n294), .B(n295), .Z(n283) );
  XOR U192 ( .A(n296), .B(n297), .Z(n295) );
  XNOR U193 ( .A(n298), .B(n299), .Z(n297) );
  XOR U194 ( .A(n300), .B(n301), .Z(n299) );
  XOR U195 ( .A(n302), .B(n303), .Z(n301) );
  XOR U196 ( .A(n304), .B(n305), .Z(n303) );
  XOR U197 ( .A(n306), .B(n307), .Z(n302) );
  XOR U198 ( .A(n308), .B(n309), .Z(n307) );
  XOR U199 ( .A(n310), .B(n311), .Z(n309) );
  XOR U200 ( .A(n312), .B(n313), .Z(n311) );
  XOR U201 ( .A(n314), .B(n315), .Z(n313) );
  XNOR U202 ( .A(n316), .B(n317), .Z(n312) );
  XNOR U203 ( .A(n318), .B(n319), .Z(n317) );
  NOR U204 ( .A(n320), .B(n315), .Z(n318) );
  XOR U205 ( .A(n321), .B(n322), .Z(n310) );
  XOR U206 ( .A(n323), .B(n324), .Z(n322) );
  XNOR U207 ( .A(n325), .B(n326), .Z(n324) );
  XOR U208 ( .A(n327), .B(n328), .Z(n326) );
  XOR U209 ( .A(n329), .B(n330), .Z(n328) );
  XOR U210 ( .A(n331), .B(n332), .Z(n330) );
  XOR U211 ( .A(n333), .B(n334), .Z(n329) );
  XOR U212 ( .A(n335), .B(n336), .Z(n334) );
  XOR U213 ( .A(n337), .B(n338), .Z(n336) );
  XOR U214 ( .A(n339), .B(n340), .Z(n338) );
  XOR U215 ( .A(n341), .B(n342), .Z(n340) );
  XNOR U216 ( .A(n343), .B(n344), .Z(n339) );
  XNOR U217 ( .A(n345), .B(n346), .Z(n344) );
  NOR U218 ( .A(n347), .B(n342), .Z(n345) );
  XOR U219 ( .A(n348), .B(n349), .Z(n337) );
  XOR U220 ( .A(n350), .B(n351), .Z(n349) );
  XNOR U221 ( .A(n352), .B(n353), .Z(n351) );
  XOR U222 ( .A(n354), .B(n355), .Z(n353) );
  XOR U223 ( .A(n356), .B(n357), .Z(n355) );
  XOR U224 ( .A(n358), .B(n359), .Z(n357) );
  XOR U225 ( .A(n360), .B(n361), .Z(n356) );
  XOR U226 ( .A(n362), .B(n363), .Z(n361) );
  XOR U227 ( .A(n364), .B(n365), .Z(n363) );
  XOR U228 ( .A(n366), .B(n367), .Z(n365) );
  XOR U229 ( .A(n368), .B(n369), .Z(n367) );
  XNOR U230 ( .A(n370), .B(n371), .Z(n366) );
  XNOR U231 ( .A(n372), .B(n373), .Z(n371) );
  NOR U232 ( .A(n374), .B(n369), .Z(n372) );
  XOR U233 ( .A(n375), .B(n376), .Z(n364) );
  XOR U234 ( .A(n377), .B(n378), .Z(n376) );
  XNOR U235 ( .A(n379), .B(n380), .Z(n378) );
  XOR U236 ( .A(n381), .B(n382), .Z(n380) );
  XOR U237 ( .A(n383), .B(n384), .Z(n382) );
  XOR U238 ( .A(n385), .B(n386), .Z(n384) );
  XOR U239 ( .A(n387), .B(n388), .Z(n383) );
  XOR U240 ( .A(n389), .B(n390), .Z(n388) );
  XOR U241 ( .A(n391), .B(n392), .Z(n390) );
  XOR U242 ( .A(n393), .B(n394), .Z(n392) );
  XOR U243 ( .A(n395), .B(n396), .Z(n394) );
  XNOR U244 ( .A(n397), .B(n398), .Z(n393) );
  XNOR U245 ( .A(n399), .B(n400), .Z(n398) );
  NOR U246 ( .A(n401), .B(n396), .Z(n399) );
  XOR U247 ( .A(n402), .B(n403), .Z(n391) );
  XOR U248 ( .A(n404), .B(n405), .Z(n403) );
  XNOR U249 ( .A(n406), .B(n407), .Z(n405) );
  XOR U250 ( .A(n408), .B(n409), .Z(n407) );
  XOR U251 ( .A(n410), .B(n411), .Z(n409) );
  XOR U252 ( .A(n412), .B(n413), .Z(n411) );
  XOR U253 ( .A(n414), .B(n415), .Z(n410) );
  XOR U254 ( .A(n416), .B(n417), .Z(n415) );
  XOR U255 ( .A(n418), .B(n419), .Z(n417) );
  XOR U256 ( .A(n420), .B(n421), .Z(n419) );
  XOR U257 ( .A(n422), .B(n423), .Z(n421) );
  XNOR U258 ( .A(n424), .B(n425), .Z(n420) );
  XNOR U259 ( .A(n426), .B(n427), .Z(n425) );
  NOR U260 ( .A(n428), .B(n423), .Z(n426) );
  XOR U261 ( .A(n429), .B(n430), .Z(n418) );
  XOR U262 ( .A(n431), .B(n432), .Z(n430) );
  XNOR U263 ( .A(n433), .B(n434), .Z(n432) );
  XOR U264 ( .A(n435), .B(n436), .Z(n434) );
  XOR U265 ( .A(n437), .B(n438), .Z(n436) );
  XOR U266 ( .A(n439), .B(n440), .Z(n438) );
  XOR U267 ( .A(n441), .B(n442), .Z(n437) );
  XOR U268 ( .A(n443), .B(n444), .Z(n442) );
  XOR U269 ( .A(n445), .B(n446), .Z(n444) );
  XOR U270 ( .A(n447), .B(n448), .Z(n446) );
  XOR U271 ( .A(n449), .B(n450), .Z(n448) );
  XNOR U272 ( .A(n451), .B(n452), .Z(n447) );
  XNOR U273 ( .A(n453), .B(n454), .Z(n452) );
  NOR U274 ( .A(n455), .B(n450), .Z(n453) );
  XOR U275 ( .A(n456), .B(n457), .Z(n445) );
  XOR U276 ( .A(n458), .B(n459), .Z(n457) );
  XNOR U277 ( .A(n460), .B(n461), .Z(n459) );
  XOR U278 ( .A(n462), .B(n463), .Z(n461) );
  XOR U279 ( .A(n464), .B(n465), .Z(n463) );
  XOR U280 ( .A(n466), .B(n467), .Z(n465) );
  XOR U281 ( .A(n468), .B(n469), .Z(n464) );
  XOR U282 ( .A(n470), .B(n471), .Z(n469) );
  XOR U283 ( .A(n472), .B(n473), .Z(n471) );
  XOR U284 ( .A(n474), .B(n475), .Z(n473) );
  XOR U285 ( .A(n476), .B(n477), .Z(n475) );
  XNOR U286 ( .A(n478), .B(n479), .Z(n474) );
  XNOR U287 ( .A(n480), .B(n481), .Z(n479) );
  NOR U288 ( .A(n482), .B(n477), .Z(n480) );
  XOR U289 ( .A(n483), .B(n484), .Z(n472) );
  XOR U290 ( .A(n485), .B(n486), .Z(n484) );
  XNOR U291 ( .A(n487), .B(n488), .Z(n486) );
  XOR U292 ( .A(n489), .B(n490), .Z(n488) );
  XOR U293 ( .A(n491), .B(n492), .Z(n490) );
  XOR U294 ( .A(n493), .B(n494), .Z(n492) );
  XOR U295 ( .A(n495), .B(n496), .Z(n491) );
  XOR U296 ( .A(n497), .B(n498), .Z(n496) );
  XOR U297 ( .A(n499), .B(n500), .Z(n498) );
  XOR U298 ( .A(n501), .B(n502), .Z(n500) );
  XOR U299 ( .A(n503), .B(n504), .Z(n502) );
  XNOR U300 ( .A(n505), .B(n506), .Z(n501) );
  XNOR U301 ( .A(n507), .B(n508), .Z(n506) );
  NOR U302 ( .A(n509), .B(n504), .Z(n507) );
  XOR U303 ( .A(n510), .B(n511), .Z(n499) );
  XOR U304 ( .A(n512), .B(n513), .Z(n511) );
  XNOR U305 ( .A(n514), .B(n515), .Z(n513) );
  XOR U306 ( .A(n516), .B(n517), .Z(n515) );
  XOR U307 ( .A(n518), .B(n519), .Z(n517) );
  XOR U308 ( .A(n520), .B(n521), .Z(n519) );
  XOR U309 ( .A(n522), .B(n523), .Z(n518) );
  XOR U310 ( .A(n524), .B(n525), .Z(n523) );
  XOR U311 ( .A(n526), .B(n527), .Z(n525) );
  XOR U312 ( .A(n528), .B(n529), .Z(n527) );
  XOR U313 ( .A(n530), .B(n531), .Z(n529) );
  XNOR U314 ( .A(n532), .B(n533), .Z(n528) );
  XNOR U315 ( .A(n534), .B(n535), .Z(n533) );
  NOR U316 ( .A(n536), .B(n531), .Z(n534) );
  XOR U317 ( .A(n537), .B(n538), .Z(n526) );
  XOR U318 ( .A(n539), .B(n540), .Z(n538) );
  XNOR U319 ( .A(n541), .B(n542), .Z(n540) );
  XOR U320 ( .A(n543), .B(n544), .Z(n542) );
  XOR U321 ( .A(n545), .B(n546), .Z(n544) );
  XOR U322 ( .A(n547), .B(n548), .Z(n546) );
  XOR U323 ( .A(n549), .B(n550), .Z(n545) );
  XOR U324 ( .A(n551), .B(n552), .Z(n550) );
  XOR U325 ( .A(n553), .B(n554), .Z(n552) );
  XOR U326 ( .A(n555), .B(n556), .Z(n554) );
  XOR U327 ( .A(n557), .B(n558), .Z(n556) );
  XNOR U328 ( .A(n559), .B(n560), .Z(n555) );
  XNOR U329 ( .A(n561), .B(n562), .Z(n560) );
  NOR U330 ( .A(n563), .B(n558), .Z(n561) );
  XOR U331 ( .A(n564), .B(n565), .Z(n553) );
  XOR U332 ( .A(n566), .B(n567), .Z(n565) );
  XNOR U333 ( .A(n568), .B(n569), .Z(n567) );
  XOR U334 ( .A(n570), .B(n571), .Z(n569) );
  XOR U335 ( .A(n572), .B(n573), .Z(n571) );
  XOR U336 ( .A(n574), .B(n575), .Z(n573) );
  XOR U337 ( .A(n576), .B(n577), .Z(n572) );
  XOR U338 ( .A(n578), .B(n579), .Z(n577) );
  XOR U339 ( .A(n580), .B(n581), .Z(n579) );
  XOR U340 ( .A(n582), .B(n583), .Z(n581) );
  XOR U341 ( .A(n584), .B(n585), .Z(n583) );
  XNOR U342 ( .A(n586), .B(n587), .Z(n582) );
  XNOR U343 ( .A(n588), .B(n589), .Z(n587) );
  NOR U344 ( .A(n590), .B(n585), .Z(n588) );
  XOR U345 ( .A(n591), .B(n592), .Z(n580) );
  XOR U346 ( .A(n593), .B(n594), .Z(n592) );
  XNOR U347 ( .A(n595), .B(n596), .Z(n594) );
  XOR U348 ( .A(n597), .B(n598), .Z(n596) );
  XOR U349 ( .A(n599), .B(n600), .Z(n598) );
  XOR U350 ( .A(n601), .B(n602), .Z(n600) );
  XOR U351 ( .A(n603), .B(n604), .Z(n599) );
  XOR U352 ( .A(n605), .B(n606), .Z(n604) );
  XOR U353 ( .A(n607), .B(n608), .Z(n606) );
  XOR U354 ( .A(n609), .B(n610), .Z(n608) );
  XOR U355 ( .A(n611), .B(n612), .Z(n610) );
  XNOR U356 ( .A(n613), .B(n614), .Z(n609) );
  XNOR U357 ( .A(n615), .B(n616), .Z(n614) );
  NOR U358 ( .A(n617), .B(n612), .Z(n615) );
  XOR U359 ( .A(n618), .B(n619), .Z(n607) );
  XOR U360 ( .A(n620), .B(n621), .Z(n619) );
  XNOR U361 ( .A(n622), .B(n623), .Z(n621) );
  XOR U362 ( .A(n624), .B(n625), .Z(n623) );
  XOR U363 ( .A(n626), .B(n627), .Z(n625) );
  XOR U364 ( .A(n628), .B(n629), .Z(n627) );
  XOR U365 ( .A(n630), .B(n631), .Z(n626) );
  XOR U366 ( .A(n632), .B(n633), .Z(n631) );
  XOR U367 ( .A(n634), .B(n635), .Z(n633) );
  XOR U368 ( .A(n636), .B(n637), .Z(n635) );
  XOR U369 ( .A(n638), .B(n639), .Z(n637) );
  XNOR U370 ( .A(n640), .B(n641), .Z(n636) );
  XNOR U371 ( .A(n642), .B(n643), .Z(n641) );
  NOR U372 ( .A(n644), .B(n639), .Z(n642) );
  XOR U373 ( .A(n645), .B(n646), .Z(n634) );
  XOR U374 ( .A(n647), .B(n648), .Z(n646) );
  XNOR U375 ( .A(n649), .B(n650), .Z(n648) );
  XOR U376 ( .A(n651), .B(n652), .Z(n650) );
  XOR U377 ( .A(n653), .B(n654), .Z(n652) );
  XOR U378 ( .A(n655), .B(n656), .Z(n654) );
  XOR U379 ( .A(n657), .B(n658), .Z(n653) );
  XOR U380 ( .A(n659), .B(n660), .Z(n658) );
  XOR U381 ( .A(n661), .B(n662), .Z(n660) );
  XOR U382 ( .A(n663), .B(n664), .Z(n662) );
  XOR U383 ( .A(n665), .B(n666), .Z(n664) );
  XNOR U384 ( .A(n667), .B(n668), .Z(n663) );
  XNOR U385 ( .A(n669), .B(n670), .Z(n668) );
  NOR U386 ( .A(n671), .B(n666), .Z(n669) );
  XOR U387 ( .A(n672), .B(n673), .Z(n661) );
  XOR U388 ( .A(n674), .B(n675), .Z(n673) );
  XNOR U389 ( .A(n676), .B(n677), .Z(n675) );
  XOR U390 ( .A(n678), .B(n679), .Z(n677) );
  XOR U391 ( .A(n680), .B(n681), .Z(n679) );
  XOR U392 ( .A(n682), .B(n683), .Z(n681) );
  XOR U393 ( .A(n684), .B(n685), .Z(n680) );
  XOR U394 ( .A(n686), .B(n687), .Z(n685) );
  XOR U395 ( .A(n688), .B(n689), .Z(n687) );
  XOR U396 ( .A(n690), .B(n691), .Z(n689) );
  XOR U397 ( .A(n692), .B(n693), .Z(n691) );
  XNOR U398 ( .A(n694), .B(n695), .Z(n690) );
  XNOR U399 ( .A(n696), .B(n697), .Z(n695) );
  NOR U400 ( .A(n698), .B(n693), .Z(n696) );
  XOR U401 ( .A(n699), .B(n700), .Z(n688) );
  XOR U402 ( .A(n701), .B(n702), .Z(n700) );
  XNOR U403 ( .A(n703), .B(n704), .Z(n702) );
  XOR U404 ( .A(n705), .B(n706), .Z(n704) );
  XOR U405 ( .A(n707), .B(n708), .Z(n706) );
  XOR U406 ( .A(n709), .B(n710), .Z(n708) );
  XOR U407 ( .A(n711), .B(n712), .Z(n707) );
  XOR U408 ( .A(n713), .B(n714), .Z(n712) );
  XOR U409 ( .A(n715), .B(n716), .Z(n714) );
  XOR U410 ( .A(n717), .B(n718), .Z(n716) );
  XOR U411 ( .A(n719), .B(n720), .Z(n718) );
  XNOR U412 ( .A(n721), .B(n722), .Z(n717) );
  XNOR U413 ( .A(n723), .B(n724), .Z(n722) );
  NOR U414 ( .A(n725), .B(n720), .Z(n723) );
  XOR U415 ( .A(n726), .B(n727), .Z(n715) );
  XOR U416 ( .A(n728), .B(n729), .Z(n727) );
  XNOR U417 ( .A(n730), .B(n731), .Z(n729) );
  XOR U418 ( .A(n732), .B(n733), .Z(n731) );
  XOR U419 ( .A(n734), .B(n735), .Z(n733) );
  XOR U420 ( .A(n736), .B(n737), .Z(n735) );
  XOR U421 ( .A(n738), .B(n739), .Z(n734) );
  XOR U422 ( .A(n740), .B(n741), .Z(n739) );
  XOR U423 ( .A(n742), .B(n743), .Z(n741) );
  XOR U424 ( .A(n744), .B(n745), .Z(n743) );
  XOR U425 ( .A(n746), .B(n747), .Z(n745) );
  XNOR U426 ( .A(n748), .B(n749), .Z(n744) );
  XNOR U427 ( .A(n750), .B(n751), .Z(n749) );
  NOR U428 ( .A(n752), .B(n747), .Z(n750) );
  XOR U429 ( .A(n753), .B(n754), .Z(n742) );
  XOR U430 ( .A(n755), .B(n756), .Z(n754) );
  XOR U431 ( .A(n757), .B(n758), .Z(n756) );
  XOR U432 ( .A(n759), .B(n760), .Z(n755) );
  XOR U433 ( .A(n761), .B(n762), .Z(n753) );
  XOR U434 ( .A(n763), .B(n764), .Z(n762) );
  AND U435 ( .A(n765), .B(n766), .Z(n764) );
  XOR U436 ( .A(n767), .B(n758), .Z(n765) );
  XOR U437 ( .A(n768), .B(n769), .Z(n758) );
  NOR U438 ( .A(n767), .B(n768), .Z(n769) );
  NOR U439 ( .A(n770), .B(n759), .Z(n763) );
  XOR U440 ( .A(n771), .B(n772), .Z(n761) );
  NOR U441 ( .A(n773), .B(n760), .Z(n772) );
  NOR U442 ( .A(n774), .B(n757), .Z(n771) );
  XOR U443 ( .A(n775), .B(n776), .Z(n740) );
  NOR U444 ( .A(n777), .B(n751), .Z(n776) );
  NOR U445 ( .A(n778), .B(n748), .Z(n775) );
  XOR U446 ( .A(n779), .B(n780), .Z(n738) );
  XOR U447 ( .A(n781), .B(n782), .Z(n780) );
  NOR U448 ( .A(n783), .B(n746), .Z(n782) );
  NOR U449 ( .A(n784), .B(n785), .Z(n781) );
  XOR U450 ( .A(n786), .B(n787), .Z(n779) );
  NOR U451 ( .A(n788), .B(n789), .Z(n787) );
  NOR U452 ( .A(n790), .B(n736), .Z(n786) );
  XOR U453 ( .A(n791), .B(n792), .Z(n732) );
  XOR U454 ( .A(n785), .B(n789), .Z(n792) );
  XOR U455 ( .A(n793), .B(n794), .Z(n791) );
  NOR U456 ( .A(n795), .B(n737), .Z(n794) );
  NOR U457 ( .A(n796), .B(n797), .Z(n793) );
  XOR U458 ( .A(n798), .B(n799), .Z(n728) );
  XOR U459 ( .A(n800), .B(n801), .Z(n726) );
  XNOR U460 ( .A(n802), .B(n797), .Z(n801) );
  NOR U461 ( .A(n803), .B(n798), .Z(n802) );
  XOR U462 ( .A(n804), .B(n805), .Z(n800) );
  NOR U463 ( .A(n806), .B(n799), .Z(n805) );
  NOR U464 ( .A(n807), .B(n730), .Z(n804) );
  XOR U465 ( .A(n808), .B(n809), .Z(n713) );
  NOR U466 ( .A(n810), .B(n724), .Z(n809) );
  NOR U467 ( .A(n811), .B(n721), .Z(n808) );
  XOR U468 ( .A(n812), .B(n813), .Z(n711) );
  XOR U469 ( .A(n814), .B(n815), .Z(n813) );
  NOR U470 ( .A(n816), .B(n719), .Z(n815) );
  NOR U471 ( .A(n817), .B(n818), .Z(n814) );
  XOR U472 ( .A(n819), .B(n820), .Z(n812) );
  NOR U473 ( .A(n821), .B(n822), .Z(n820) );
  NOR U474 ( .A(n823), .B(n709), .Z(n819) );
  XOR U475 ( .A(n824), .B(n825), .Z(n705) );
  XOR U476 ( .A(n818), .B(n822), .Z(n825) );
  XOR U477 ( .A(n826), .B(n827), .Z(n824) );
  NOR U478 ( .A(n828), .B(n710), .Z(n827) );
  NOR U479 ( .A(n829), .B(n830), .Z(n826) );
  XOR U480 ( .A(n831), .B(n832), .Z(n701) );
  XOR U481 ( .A(n833), .B(n834), .Z(n699) );
  XNOR U482 ( .A(n835), .B(n830), .Z(n834) );
  NOR U483 ( .A(n836), .B(n831), .Z(n835) );
  XOR U484 ( .A(n837), .B(n838), .Z(n833) );
  NOR U485 ( .A(n839), .B(n832), .Z(n838) );
  NOR U486 ( .A(n840), .B(n703), .Z(n837) );
  XOR U487 ( .A(n841), .B(n842), .Z(n686) );
  NOR U488 ( .A(n843), .B(n697), .Z(n842) );
  NOR U489 ( .A(n844), .B(n694), .Z(n841) );
  XOR U490 ( .A(n845), .B(n846), .Z(n684) );
  XOR U491 ( .A(n847), .B(n848), .Z(n846) );
  NOR U492 ( .A(n849), .B(n692), .Z(n848) );
  NOR U493 ( .A(n850), .B(n851), .Z(n847) );
  XOR U494 ( .A(n852), .B(n853), .Z(n845) );
  NOR U495 ( .A(n854), .B(n855), .Z(n853) );
  NOR U496 ( .A(n856), .B(n682), .Z(n852) );
  XOR U497 ( .A(n857), .B(n858), .Z(n678) );
  XOR U498 ( .A(n851), .B(n855), .Z(n858) );
  XOR U499 ( .A(n859), .B(n860), .Z(n857) );
  NOR U500 ( .A(n861), .B(n683), .Z(n860) );
  NOR U501 ( .A(n862), .B(n863), .Z(n859) );
  XOR U502 ( .A(n864), .B(n865), .Z(n674) );
  XOR U503 ( .A(n866), .B(n867), .Z(n672) );
  XNOR U504 ( .A(n868), .B(n863), .Z(n867) );
  NOR U505 ( .A(n869), .B(n864), .Z(n868) );
  XOR U506 ( .A(n870), .B(n871), .Z(n866) );
  NOR U507 ( .A(n872), .B(n865), .Z(n871) );
  NOR U508 ( .A(n873), .B(n676), .Z(n870) );
  XOR U509 ( .A(n874), .B(n875), .Z(n659) );
  NOR U510 ( .A(n876), .B(n670), .Z(n875) );
  NOR U511 ( .A(n877), .B(n667), .Z(n874) );
  XOR U512 ( .A(n878), .B(n879), .Z(n657) );
  XOR U513 ( .A(n880), .B(n881), .Z(n879) );
  NOR U514 ( .A(n882), .B(n665), .Z(n881) );
  NOR U515 ( .A(n883), .B(n884), .Z(n880) );
  XOR U516 ( .A(n885), .B(n886), .Z(n878) );
  NOR U517 ( .A(n887), .B(n888), .Z(n886) );
  NOR U518 ( .A(n889), .B(n655), .Z(n885) );
  XOR U519 ( .A(n890), .B(n891), .Z(n651) );
  XOR U520 ( .A(n884), .B(n888), .Z(n891) );
  XOR U521 ( .A(n892), .B(n893), .Z(n890) );
  NOR U522 ( .A(n894), .B(n656), .Z(n893) );
  NOR U523 ( .A(n895), .B(n896), .Z(n892) );
  XOR U524 ( .A(n897), .B(n898), .Z(n647) );
  XOR U525 ( .A(n899), .B(n900), .Z(n645) );
  XNOR U526 ( .A(n901), .B(n896), .Z(n900) );
  NOR U527 ( .A(n902), .B(n897), .Z(n901) );
  XOR U528 ( .A(n903), .B(n904), .Z(n899) );
  NOR U529 ( .A(n905), .B(n898), .Z(n904) );
  NOR U530 ( .A(n906), .B(n649), .Z(n903) );
  XOR U531 ( .A(n907), .B(n908), .Z(n632) );
  NOR U532 ( .A(n909), .B(n643), .Z(n908) );
  NOR U533 ( .A(n910), .B(n640), .Z(n907) );
  XOR U534 ( .A(n911), .B(n912), .Z(n630) );
  XOR U535 ( .A(n913), .B(n914), .Z(n912) );
  NOR U536 ( .A(n915), .B(n638), .Z(n914) );
  NOR U537 ( .A(n916), .B(n917), .Z(n913) );
  XOR U538 ( .A(n918), .B(n919), .Z(n911) );
  NOR U539 ( .A(n920), .B(n921), .Z(n919) );
  NOR U540 ( .A(n922), .B(n628), .Z(n918) );
  XOR U541 ( .A(n923), .B(n924), .Z(n624) );
  XOR U542 ( .A(n917), .B(n921), .Z(n924) );
  XOR U543 ( .A(n925), .B(n926), .Z(n923) );
  NOR U544 ( .A(n927), .B(n629), .Z(n926) );
  NOR U545 ( .A(n928), .B(n929), .Z(n925) );
  XOR U546 ( .A(n930), .B(n931), .Z(n620) );
  XOR U547 ( .A(n932), .B(n933), .Z(n618) );
  XNOR U548 ( .A(n934), .B(n929), .Z(n933) );
  NOR U549 ( .A(n935), .B(n930), .Z(n934) );
  XOR U550 ( .A(n936), .B(n937), .Z(n932) );
  NOR U551 ( .A(n938), .B(n931), .Z(n937) );
  NOR U552 ( .A(n939), .B(n622), .Z(n936) );
  XOR U553 ( .A(n940), .B(n941), .Z(n605) );
  NOR U554 ( .A(n942), .B(n616), .Z(n941) );
  NOR U555 ( .A(n943), .B(n613), .Z(n940) );
  XOR U556 ( .A(n944), .B(n945), .Z(n603) );
  XOR U557 ( .A(n946), .B(n947), .Z(n945) );
  NOR U558 ( .A(n948), .B(n611), .Z(n947) );
  NOR U559 ( .A(n949), .B(n950), .Z(n946) );
  XOR U560 ( .A(n951), .B(n952), .Z(n944) );
  NOR U561 ( .A(n953), .B(n954), .Z(n952) );
  NOR U562 ( .A(n955), .B(n601), .Z(n951) );
  XOR U563 ( .A(n956), .B(n957), .Z(n597) );
  XOR U564 ( .A(n950), .B(n954), .Z(n957) );
  XOR U565 ( .A(n958), .B(n959), .Z(n956) );
  NOR U566 ( .A(n960), .B(n602), .Z(n959) );
  NOR U567 ( .A(n961), .B(n962), .Z(n958) );
  XOR U568 ( .A(n963), .B(n964), .Z(n593) );
  XOR U569 ( .A(n965), .B(n966), .Z(n591) );
  XNOR U570 ( .A(n967), .B(n962), .Z(n966) );
  NOR U571 ( .A(n968), .B(n963), .Z(n967) );
  XOR U572 ( .A(n969), .B(n970), .Z(n965) );
  NOR U573 ( .A(n971), .B(n964), .Z(n970) );
  NOR U574 ( .A(n972), .B(n595), .Z(n969) );
  XOR U575 ( .A(n973), .B(n974), .Z(n578) );
  NOR U576 ( .A(n975), .B(n589), .Z(n974) );
  NOR U577 ( .A(n976), .B(n586), .Z(n973) );
  XOR U578 ( .A(n977), .B(n978), .Z(n576) );
  XOR U579 ( .A(n979), .B(n980), .Z(n978) );
  NOR U580 ( .A(n981), .B(n584), .Z(n980) );
  NOR U581 ( .A(n982), .B(n983), .Z(n979) );
  XOR U582 ( .A(n984), .B(n985), .Z(n977) );
  NOR U583 ( .A(n986), .B(n987), .Z(n985) );
  NOR U584 ( .A(n988), .B(n574), .Z(n984) );
  XOR U585 ( .A(n989), .B(n990), .Z(n570) );
  XOR U586 ( .A(n983), .B(n987), .Z(n990) );
  XOR U587 ( .A(n991), .B(n992), .Z(n989) );
  NOR U588 ( .A(n993), .B(n575), .Z(n992) );
  NOR U589 ( .A(n994), .B(n995), .Z(n991) );
  XOR U590 ( .A(n996), .B(n997), .Z(n566) );
  XOR U591 ( .A(n998), .B(n999), .Z(n564) );
  XNOR U592 ( .A(n1000), .B(n995), .Z(n999) );
  NOR U593 ( .A(n1001), .B(n996), .Z(n1000) );
  XOR U594 ( .A(n1002), .B(n1003), .Z(n998) );
  NOR U595 ( .A(n1004), .B(n997), .Z(n1003) );
  NOR U596 ( .A(n1005), .B(n568), .Z(n1002) );
  XOR U597 ( .A(n1006), .B(n1007), .Z(n551) );
  NOR U598 ( .A(n1008), .B(n562), .Z(n1007) );
  NOR U599 ( .A(n1009), .B(n559), .Z(n1006) );
  XOR U600 ( .A(n1010), .B(n1011), .Z(n549) );
  XOR U601 ( .A(n1012), .B(n1013), .Z(n1011) );
  NOR U602 ( .A(n1014), .B(n557), .Z(n1013) );
  NOR U603 ( .A(n1015), .B(n1016), .Z(n1012) );
  XOR U604 ( .A(n1017), .B(n1018), .Z(n1010) );
  NOR U605 ( .A(n1019), .B(n1020), .Z(n1018) );
  NOR U606 ( .A(n1021), .B(n547), .Z(n1017) );
  XOR U607 ( .A(n1022), .B(n1023), .Z(n543) );
  XOR U608 ( .A(n1016), .B(n1020), .Z(n1023) );
  XOR U609 ( .A(n1024), .B(n1025), .Z(n1022) );
  NOR U610 ( .A(n1026), .B(n548), .Z(n1025) );
  NOR U611 ( .A(n1027), .B(n1028), .Z(n1024) );
  XOR U612 ( .A(n1029), .B(n1030), .Z(n539) );
  XOR U613 ( .A(n1031), .B(n1032), .Z(n537) );
  XNOR U614 ( .A(n1033), .B(n1028), .Z(n1032) );
  NOR U615 ( .A(n1034), .B(n1029), .Z(n1033) );
  XOR U616 ( .A(n1035), .B(n1036), .Z(n1031) );
  NOR U617 ( .A(n1037), .B(n1030), .Z(n1036) );
  NOR U618 ( .A(n1038), .B(n541), .Z(n1035) );
  XOR U619 ( .A(n1039), .B(n1040), .Z(n524) );
  NOR U620 ( .A(n1041), .B(n535), .Z(n1040) );
  NOR U621 ( .A(n1042), .B(n532), .Z(n1039) );
  XOR U622 ( .A(n1043), .B(n1044), .Z(n522) );
  XOR U623 ( .A(n1045), .B(n1046), .Z(n1044) );
  NOR U624 ( .A(n1047), .B(n530), .Z(n1046) );
  NOR U625 ( .A(n1048), .B(n1049), .Z(n1045) );
  XOR U626 ( .A(n1050), .B(n1051), .Z(n1043) );
  NOR U627 ( .A(n1052), .B(n1053), .Z(n1051) );
  NOR U628 ( .A(n1054), .B(n520), .Z(n1050) );
  XOR U629 ( .A(n1055), .B(n1056), .Z(n516) );
  XOR U630 ( .A(n1049), .B(n1053), .Z(n1056) );
  XOR U631 ( .A(n1057), .B(n1058), .Z(n1055) );
  NOR U632 ( .A(n1059), .B(n521), .Z(n1058) );
  NOR U633 ( .A(n1060), .B(n1061), .Z(n1057) );
  XOR U634 ( .A(n1062), .B(n1063), .Z(n512) );
  XOR U635 ( .A(n1064), .B(n1065), .Z(n510) );
  XNOR U636 ( .A(n1066), .B(n1061), .Z(n1065) );
  NOR U637 ( .A(n1067), .B(n1062), .Z(n1066) );
  XOR U638 ( .A(n1068), .B(n1069), .Z(n1064) );
  NOR U639 ( .A(n1070), .B(n1063), .Z(n1069) );
  NOR U640 ( .A(n1071), .B(n514), .Z(n1068) );
  XOR U641 ( .A(n1072), .B(n1073), .Z(n497) );
  NOR U642 ( .A(n1074), .B(n508), .Z(n1073) );
  NOR U643 ( .A(n1075), .B(n505), .Z(n1072) );
  XOR U644 ( .A(n1076), .B(n1077), .Z(n495) );
  XOR U645 ( .A(n1078), .B(n1079), .Z(n1077) );
  NOR U646 ( .A(n1080), .B(n503), .Z(n1079) );
  NOR U647 ( .A(n1081), .B(n1082), .Z(n1078) );
  XOR U648 ( .A(n1083), .B(n1084), .Z(n1076) );
  NOR U649 ( .A(n1085), .B(n1086), .Z(n1084) );
  NOR U650 ( .A(n1087), .B(n493), .Z(n1083) );
  XOR U651 ( .A(n1088), .B(n1089), .Z(n489) );
  XOR U652 ( .A(n1082), .B(n1086), .Z(n1089) );
  XOR U653 ( .A(n1090), .B(n1091), .Z(n1088) );
  NOR U654 ( .A(n1092), .B(n494), .Z(n1091) );
  NOR U655 ( .A(n1093), .B(n1094), .Z(n1090) );
  XOR U656 ( .A(n1095), .B(n1096), .Z(n485) );
  XOR U657 ( .A(n1097), .B(n1098), .Z(n483) );
  XNOR U658 ( .A(n1099), .B(n1094), .Z(n1098) );
  NOR U659 ( .A(n1100), .B(n1095), .Z(n1099) );
  XOR U660 ( .A(n1101), .B(n1102), .Z(n1097) );
  NOR U661 ( .A(n1103), .B(n1096), .Z(n1102) );
  NOR U662 ( .A(n1104), .B(n487), .Z(n1101) );
  XOR U663 ( .A(n1105), .B(n1106), .Z(n470) );
  NOR U664 ( .A(n1107), .B(n481), .Z(n1106) );
  NOR U665 ( .A(n1108), .B(n478), .Z(n1105) );
  XOR U666 ( .A(n1109), .B(n1110), .Z(n468) );
  XOR U667 ( .A(n1111), .B(n1112), .Z(n1110) );
  NOR U668 ( .A(n1113), .B(n476), .Z(n1112) );
  NOR U669 ( .A(n1114), .B(n1115), .Z(n1111) );
  XOR U670 ( .A(n1116), .B(n1117), .Z(n1109) );
  NOR U671 ( .A(n1118), .B(n1119), .Z(n1117) );
  NOR U672 ( .A(n1120), .B(n466), .Z(n1116) );
  XOR U673 ( .A(n1121), .B(n1122), .Z(n462) );
  XOR U674 ( .A(n1115), .B(n1119), .Z(n1122) );
  XOR U675 ( .A(n1123), .B(n1124), .Z(n1121) );
  NOR U676 ( .A(n1125), .B(n467), .Z(n1124) );
  NOR U677 ( .A(n1126), .B(n1127), .Z(n1123) );
  XOR U678 ( .A(n1128), .B(n1129), .Z(n458) );
  XOR U679 ( .A(n1130), .B(n1131), .Z(n456) );
  XNOR U680 ( .A(n1132), .B(n1127), .Z(n1131) );
  NOR U681 ( .A(n1133), .B(n1128), .Z(n1132) );
  XOR U682 ( .A(n1134), .B(n1135), .Z(n1130) );
  NOR U683 ( .A(n1136), .B(n1129), .Z(n1135) );
  NOR U684 ( .A(n1137), .B(n460), .Z(n1134) );
  XOR U685 ( .A(n1138), .B(n1139), .Z(n443) );
  NOR U686 ( .A(n1140), .B(n454), .Z(n1139) );
  NOR U687 ( .A(n1141), .B(n451), .Z(n1138) );
  XOR U688 ( .A(n1142), .B(n1143), .Z(n441) );
  XOR U689 ( .A(n1144), .B(n1145), .Z(n1143) );
  NOR U690 ( .A(n1146), .B(n449), .Z(n1145) );
  NOR U691 ( .A(n1147), .B(n1148), .Z(n1144) );
  XOR U692 ( .A(n1149), .B(n1150), .Z(n1142) );
  NOR U693 ( .A(n1151), .B(n1152), .Z(n1150) );
  NOR U694 ( .A(n1153), .B(n439), .Z(n1149) );
  XOR U695 ( .A(n1154), .B(n1155), .Z(n435) );
  XOR U696 ( .A(n1148), .B(n1152), .Z(n1155) );
  XOR U697 ( .A(n1156), .B(n1157), .Z(n1154) );
  NOR U698 ( .A(n1158), .B(n440), .Z(n1157) );
  NOR U699 ( .A(n1159), .B(n1160), .Z(n1156) );
  XOR U700 ( .A(n1161), .B(n1162), .Z(n431) );
  XOR U701 ( .A(n1163), .B(n1164), .Z(n429) );
  XNOR U702 ( .A(n1165), .B(n1160), .Z(n1164) );
  NOR U703 ( .A(n1166), .B(n1161), .Z(n1165) );
  XOR U704 ( .A(n1167), .B(n1168), .Z(n1163) );
  NOR U705 ( .A(n1169), .B(n1162), .Z(n1168) );
  NOR U706 ( .A(n1170), .B(n433), .Z(n1167) );
  XOR U707 ( .A(n1171), .B(n1172), .Z(n416) );
  NOR U708 ( .A(n1173), .B(n427), .Z(n1172) );
  NOR U709 ( .A(n1174), .B(n424), .Z(n1171) );
  XOR U710 ( .A(n1175), .B(n1176), .Z(n414) );
  XOR U711 ( .A(n1177), .B(n1178), .Z(n1176) );
  NOR U712 ( .A(n1179), .B(n422), .Z(n1178) );
  NOR U713 ( .A(n1180), .B(n1181), .Z(n1177) );
  XOR U714 ( .A(n1182), .B(n1183), .Z(n1175) );
  NOR U715 ( .A(n1184), .B(n1185), .Z(n1183) );
  NOR U716 ( .A(n1186), .B(n412), .Z(n1182) );
  XOR U717 ( .A(n1187), .B(n1188), .Z(n408) );
  XOR U718 ( .A(n1181), .B(n1185), .Z(n1188) );
  XOR U719 ( .A(n1189), .B(n1190), .Z(n1187) );
  NOR U720 ( .A(n1191), .B(n413), .Z(n1190) );
  NOR U721 ( .A(n1192), .B(n1193), .Z(n1189) );
  XOR U722 ( .A(n1194), .B(n1195), .Z(n404) );
  XOR U723 ( .A(n1196), .B(n1197), .Z(n402) );
  XNOR U724 ( .A(n1198), .B(n1193), .Z(n1197) );
  NOR U725 ( .A(n1199), .B(n1194), .Z(n1198) );
  XOR U726 ( .A(n1200), .B(n1201), .Z(n1196) );
  NOR U727 ( .A(n1202), .B(n1195), .Z(n1201) );
  NOR U728 ( .A(n1203), .B(n406), .Z(n1200) );
  XOR U729 ( .A(n1204), .B(n1205), .Z(n389) );
  NOR U730 ( .A(n1206), .B(n400), .Z(n1205) );
  NOR U731 ( .A(n1207), .B(n397), .Z(n1204) );
  XOR U732 ( .A(n1208), .B(n1209), .Z(n387) );
  XOR U733 ( .A(n1210), .B(n1211), .Z(n1209) );
  NOR U734 ( .A(n1212), .B(n395), .Z(n1211) );
  NOR U735 ( .A(n1213), .B(n1214), .Z(n1210) );
  XOR U736 ( .A(n1215), .B(n1216), .Z(n1208) );
  NOR U737 ( .A(n1217), .B(n1218), .Z(n1216) );
  NOR U738 ( .A(n1219), .B(n385), .Z(n1215) );
  XOR U739 ( .A(n1220), .B(n1221), .Z(n381) );
  XOR U740 ( .A(n1214), .B(n1218), .Z(n1221) );
  XOR U741 ( .A(n1222), .B(n1223), .Z(n1220) );
  NOR U742 ( .A(n1224), .B(n386), .Z(n1223) );
  NOR U743 ( .A(n1225), .B(n1226), .Z(n1222) );
  XOR U744 ( .A(n1227), .B(n1228), .Z(n377) );
  XOR U745 ( .A(n1229), .B(n1230), .Z(n375) );
  XNOR U746 ( .A(n1231), .B(n1226), .Z(n1230) );
  NOR U747 ( .A(n1232), .B(n1227), .Z(n1231) );
  XOR U748 ( .A(n1233), .B(n1234), .Z(n1229) );
  NOR U749 ( .A(n1235), .B(n1228), .Z(n1234) );
  NOR U750 ( .A(n1236), .B(n379), .Z(n1233) );
  XOR U751 ( .A(n1237), .B(n1238), .Z(n362) );
  NOR U752 ( .A(n1239), .B(n373), .Z(n1238) );
  NOR U753 ( .A(n1240), .B(n370), .Z(n1237) );
  XOR U754 ( .A(n1241), .B(n1242), .Z(n360) );
  XOR U755 ( .A(n1243), .B(n1244), .Z(n1242) );
  NOR U756 ( .A(n1245), .B(n368), .Z(n1244) );
  NOR U757 ( .A(n1246), .B(n1247), .Z(n1243) );
  XOR U758 ( .A(n1248), .B(n1249), .Z(n1241) );
  NOR U759 ( .A(n1250), .B(n1251), .Z(n1249) );
  NOR U760 ( .A(n1252), .B(n358), .Z(n1248) );
  XOR U761 ( .A(n1253), .B(n1254), .Z(n354) );
  XOR U762 ( .A(n1247), .B(n1251), .Z(n1254) );
  XOR U763 ( .A(n1255), .B(n1256), .Z(n1253) );
  NOR U764 ( .A(n1257), .B(n359), .Z(n1256) );
  NOR U765 ( .A(n1258), .B(n1259), .Z(n1255) );
  XOR U766 ( .A(n1260), .B(n1261), .Z(n350) );
  XOR U767 ( .A(n1262), .B(n1263), .Z(n348) );
  XNOR U768 ( .A(n1264), .B(n1259), .Z(n1263) );
  NOR U769 ( .A(n1265), .B(n1260), .Z(n1264) );
  XOR U770 ( .A(n1266), .B(n1267), .Z(n1262) );
  NOR U771 ( .A(n1268), .B(n1261), .Z(n1267) );
  NOR U772 ( .A(n1269), .B(n352), .Z(n1266) );
  XOR U773 ( .A(n1270), .B(n1271), .Z(n335) );
  NOR U774 ( .A(n1272), .B(n346), .Z(n1271) );
  NOR U775 ( .A(n1273), .B(n343), .Z(n1270) );
  XOR U776 ( .A(n1274), .B(n1275), .Z(n333) );
  XOR U777 ( .A(n1276), .B(n1277), .Z(n1275) );
  NOR U778 ( .A(n1278), .B(n341), .Z(n1277) );
  NOR U779 ( .A(n1279), .B(n1280), .Z(n1276) );
  XOR U780 ( .A(n1281), .B(n1282), .Z(n1274) );
  NOR U781 ( .A(n1283), .B(n1284), .Z(n1282) );
  NOR U782 ( .A(n1285), .B(n331), .Z(n1281) );
  XOR U783 ( .A(n1286), .B(n1287), .Z(n327) );
  XOR U784 ( .A(n1280), .B(n1284), .Z(n1287) );
  XOR U785 ( .A(n1288), .B(n1289), .Z(n1286) );
  NOR U786 ( .A(n1290), .B(n332), .Z(n1289) );
  NOR U787 ( .A(n1291), .B(n1292), .Z(n1288) );
  XOR U788 ( .A(n1293), .B(n1294), .Z(n323) );
  XOR U789 ( .A(n1295), .B(n1296), .Z(n321) );
  XNOR U790 ( .A(n1297), .B(n1292), .Z(n1296) );
  NOR U791 ( .A(n1298), .B(n1293), .Z(n1297) );
  XOR U792 ( .A(n1299), .B(n1300), .Z(n1295) );
  NOR U793 ( .A(n1301), .B(n1294), .Z(n1300) );
  NOR U794 ( .A(n1302), .B(n325), .Z(n1299) );
  XOR U795 ( .A(n1303), .B(n1304), .Z(n308) );
  NOR U796 ( .A(n1305), .B(n319), .Z(n1304) );
  NOR U797 ( .A(n1306), .B(n316), .Z(n1303) );
  XOR U798 ( .A(n1307), .B(n1308), .Z(n306) );
  XOR U799 ( .A(n1309), .B(n1310), .Z(n1308) );
  NOR U800 ( .A(n1311), .B(n314), .Z(n1310) );
  NOR U801 ( .A(n1312), .B(n1313), .Z(n1309) );
  XOR U802 ( .A(n1314), .B(n1315), .Z(n1307) );
  NOR U803 ( .A(n1316), .B(n1317), .Z(n1315) );
  NOR U804 ( .A(n1318), .B(n304), .Z(n1314) );
  XOR U805 ( .A(n1319), .B(n1320), .Z(n300) );
  XOR U806 ( .A(n1313), .B(n1317), .Z(n1320) );
  XOR U807 ( .A(n1321), .B(n1322), .Z(n1319) );
  NOR U808 ( .A(n1323), .B(n305), .Z(n1322) );
  NOR U809 ( .A(n1324), .B(n1325), .Z(n1321) );
  XOR U810 ( .A(n1326), .B(n1327), .Z(n296) );
  XOR U811 ( .A(n1328), .B(n1329), .Z(n294) );
  XNOR U812 ( .A(n1330), .B(n1325), .Z(n1329) );
  NOR U813 ( .A(n1331), .B(n1326), .Z(n1330) );
  XOR U814 ( .A(n1332), .B(n1333), .Z(n1328) );
  NOR U815 ( .A(n1334), .B(n1327), .Z(n1333) );
  NOR U816 ( .A(n1335), .B(n298), .Z(n1332) );
  XOR U817 ( .A(n1336), .B(n1337), .Z(n281) );
  NOR U818 ( .A(n1338), .B(n292), .Z(n1337) );
  NOR U819 ( .A(n1339), .B(n289), .Z(n1336) );
  XOR U820 ( .A(n1340), .B(n1341), .Z(n279) );
  XOR U821 ( .A(n1342), .B(n1343), .Z(n1341) );
  NOR U822 ( .A(n1344), .B(n287), .Z(n1343) );
  NOR U823 ( .A(n1345), .B(n1346), .Z(n1342) );
  XOR U824 ( .A(n1347), .B(n1348), .Z(n1340) );
  NOR U825 ( .A(n1349), .B(n1350), .Z(n1348) );
  NOR U826 ( .A(n1351), .B(n277), .Z(n1347) );
  XOR U827 ( .A(n1352), .B(n1353), .Z(n273) );
  XOR U828 ( .A(n1346), .B(n1350), .Z(n1353) );
  XOR U829 ( .A(n1354), .B(n1355), .Z(n1352) );
  NOR U830 ( .A(n1356), .B(n278), .Z(n1355) );
  NOR U831 ( .A(n1357), .B(n1358), .Z(n1354) );
  XOR U832 ( .A(n1359), .B(n1360), .Z(n269) );
  XOR U833 ( .A(n1361), .B(n1362), .Z(n267) );
  XNOR U834 ( .A(n1363), .B(n1358), .Z(n1362) );
  NOR U835 ( .A(n1364), .B(n1359), .Z(n1363) );
  XOR U836 ( .A(n1365), .B(n1366), .Z(n1361) );
  NOR U837 ( .A(n1367), .B(n1360), .Z(n1366) );
  NOR U838 ( .A(n1368), .B(n271), .Z(n1365) );
  XOR U839 ( .A(n1369), .B(n1370), .Z(n254) );
  NOR U840 ( .A(n1371), .B(n265), .Z(n1370) );
  NOR U841 ( .A(n1372), .B(n262), .Z(n1369) );
  XOR U842 ( .A(n1373), .B(n1374), .Z(n252) );
  XOR U843 ( .A(n1375), .B(n1376), .Z(n1374) );
  NOR U844 ( .A(n1377), .B(n260), .Z(n1376) );
  NOR U845 ( .A(n1378), .B(n1379), .Z(n1375) );
  XOR U846 ( .A(n1380), .B(n1381), .Z(n1373) );
  NOR U847 ( .A(n1382), .B(n1383), .Z(n1381) );
  NOR U848 ( .A(n1384), .B(n250), .Z(n1380) );
  XOR U849 ( .A(n1385), .B(n1386), .Z(n246) );
  XOR U850 ( .A(n1379), .B(n1383), .Z(n1386) );
  XOR U851 ( .A(n1387), .B(n1388), .Z(n1385) );
  NOR U852 ( .A(n1389), .B(n251), .Z(n1388) );
  NOR U853 ( .A(n1390), .B(n1391), .Z(n1387) );
  XOR U854 ( .A(n1392), .B(n1393), .Z(n242) );
  XOR U855 ( .A(n1394), .B(n1395), .Z(n240) );
  XNOR U856 ( .A(n1396), .B(n1391), .Z(n1395) );
  NOR U857 ( .A(n1397), .B(n1392), .Z(n1396) );
  XOR U858 ( .A(n1398), .B(n1399), .Z(n1394) );
  NOR U859 ( .A(n1400), .B(n1393), .Z(n1399) );
  NOR U860 ( .A(n1401), .B(n244), .Z(n1398) );
  XOR U861 ( .A(n1402), .B(n1403), .Z(n227) );
  NOR U862 ( .A(n1404), .B(n238), .Z(n1403) );
  NOR U863 ( .A(n1405), .B(n235), .Z(n1402) );
  XOR U864 ( .A(n1406), .B(n1407), .Z(n225) );
  XOR U865 ( .A(n1408), .B(n1409), .Z(n1407) );
  NOR U866 ( .A(n1410), .B(n233), .Z(n1409) );
  NOR U867 ( .A(n1411), .B(n1412), .Z(n1408) );
  XOR U868 ( .A(n1413), .B(n1414), .Z(n1406) );
  NOR U869 ( .A(n1415), .B(n1416), .Z(n1414) );
  NOR U870 ( .A(n1417), .B(n223), .Z(n1413) );
  XOR U871 ( .A(n1418), .B(n1419), .Z(n219) );
  XOR U872 ( .A(n1412), .B(n1416), .Z(n1419) );
  XOR U873 ( .A(n1420), .B(n1421), .Z(n1418) );
  NOR U874 ( .A(n1422), .B(n224), .Z(n1421) );
  NOR U875 ( .A(n1423), .B(n1424), .Z(n1420) );
  XOR U876 ( .A(n1425), .B(n1426), .Z(n215) );
  XOR U877 ( .A(n1427), .B(n1428), .Z(n213) );
  XNOR U878 ( .A(n1429), .B(n1424), .Z(n1428) );
  NOR U879 ( .A(n1430), .B(n1425), .Z(n1429) );
  XOR U880 ( .A(n1431), .B(n1432), .Z(n1427) );
  NOR U881 ( .A(n1433), .B(n1426), .Z(n1432) );
  NOR U882 ( .A(n1434), .B(n217), .Z(n1431) );
  XOR U883 ( .A(n1435), .B(n1436), .Z(n200) );
  NOR U884 ( .A(n1437), .B(n211), .Z(n1436) );
  NOR U885 ( .A(n1438), .B(n208), .Z(n1435) );
  XOR U886 ( .A(n1439), .B(n1440), .Z(n198) );
  XOR U887 ( .A(n1441), .B(n1442), .Z(n1440) );
  NOR U888 ( .A(n1443), .B(n206), .Z(n1442) );
  NOR U889 ( .A(n1444), .B(n189), .Z(n1441) );
  XOR U890 ( .A(n1445), .B(n1446), .Z(n1439) );
  NOR U891 ( .A(n1447), .B(n190), .Z(n1446) );
  NOR U892 ( .A(n1448), .B(n1449), .Z(n1445) );
  XNOR U893 ( .A(n194), .B(n1449), .Z(n196) );
  XNOR U894 ( .A(n1450), .B(n1451), .Z(n154) );
  NOR U895 ( .A(n44), .B(n1450), .Z(n1451) );
  XNOR U896 ( .A(n160), .B(n164), .Z(n166) );
  XOR U897 ( .A(n161), .B(n159), .Z(n160) );
  XNOR U898 ( .A(n1452), .B(n1453), .Z(n159) );
  XOR U899 ( .A(n1454), .B(n1455), .Z(n1453) );
  XOR U900 ( .A(n1456), .B(n1457), .Z(n1455) );
  AND U901 ( .A(n1458), .B(n1457), .Z(n1456) );
  XOR U902 ( .A(n1459), .B(n1460), .Z(n1454) );
  AND U903 ( .A(n1461), .B(n1462), .Z(n1460) );
  NOR U904 ( .A(n1463), .B(n1464), .Z(n1459) );
  XOR U905 ( .A(n1465), .B(n1466), .Z(n1452) );
  XOR U906 ( .A(n1467), .B(n1468), .Z(n1466) );
  XOR U907 ( .A(n1469), .B(n1470), .Z(n1468) );
  XOR U908 ( .A(n1471), .B(n1472), .Z(n1470) );
  XOR U909 ( .A(n1473), .B(n1474), .Z(n1472) );
  AND U910 ( .A(n1475), .B(n1474), .Z(n1473) );
  XOR U911 ( .A(n1476), .B(n1477), .Z(n1471) );
  XOR U912 ( .A(n1478), .B(n1479), .Z(n1477) );
  XOR U913 ( .A(n1480), .B(n1481), .Z(n1479) );
  XNOR U914 ( .A(n1482), .B(n1483), .Z(n1481) );
  NOR U915 ( .A(n1484), .B(n1483), .Z(n1482) );
  XOR U916 ( .A(n1485), .B(n1486), .Z(n1480) );
  XOR U917 ( .A(n1487), .B(n1488), .Z(n1486) );
  XOR U918 ( .A(n1489), .B(n1490), .Z(n1488) );
  XNOR U919 ( .A(n1491), .B(n1492), .Z(n1490) );
  NOR U920 ( .A(n1493), .B(n1492), .Z(n1491) );
  XOR U921 ( .A(n1494), .B(n1495), .Z(n1489) );
  XOR U922 ( .A(n1496), .B(n1497), .Z(n1495) );
  XOR U923 ( .A(n1498), .B(n1499), .Z(n1497) );
  XNOR U924 ( .A(n1500), .B(n1501), .Z(n1499) );
  NOR U925 ( .A(n1502), .B(n1501), .Z(n1500) );
  XOR U926 ( .A(n1503), .B(n1504), .Z(n1498) );
  XOR U927 ( .A(n1505), .B(n1506), .Z(n1504) );
  XOR U928 ( .A(n1507), .B(n1508), .Z(n1506) );
  XNOR U929 ( .A(n1509), .B(n1510), .Z(n1508) );
  NOR U930 ( .A(n1511), .B(n1510), .Z(n1509) );
  XOR U931 ( .A(n1512), .B(n1513), .Z(n1507) );
  XOR U932 ( .A(n1514), .B(n1515), .Z(n1513) );
  XOR U933 ( .A(n1516), .B(n1517), .Z(n1515) );
  XNOR U934 ( .A(n1518), .B(n1519), .Z(n1517) );
  NOR U935 ( .A(n1520), .B(n1519), .Z(n1518) );
  XOR U936 ( .A(n1521), .B(n1522), .Z(n1516) );
  XOR U937 ( .A(n1523), .B(n1524), .Z(n1522) );
  XOR U938 ( .A(n1525), .B(n1526), .Z(n1524) );
  XNOR U939 ( .A(n1527), .B(n1528), .Z(n1526) );
  NOR U940 ( .A(n1529), .B(n1528), .Z(n1527) );
  XOR U941 ( .A(n1530), .B(n1531), .Z(n1525) );
  XOR U942 ( .A(n1532), .B(n1533), .Z(n1531) );
  XOR U943 ( .A(n1534), .B(n1535), .Z(n1533) );
  XNOR U944 ( .A(n1536), .B(n1537), .Z(n1535) );
  NOR U945 ( .A(n1538), .B(n1537), .Z(n1536) );
  XOR U946 ( .A(n1539), .B(n1540), .Z(n1534) );
  XOR U947 ( .A(n1541), .B(n1542), .Z(n1540) );
  XOR U948 ( .A(n1543), .B(n1544), .Z(n1542) );
  XNOR U949 ( .A(n1545), .B(n1546), .Z(n1544) );
  NOR U950 ( .A(n1547), .B(n1546), .Z(n1545) );
  XOR U951 ( .A(n1548), .B(n1549), .Z(n1543) );
  XOR U952 ( .A(n1550), .B(n1551), .Z(n1549) );
  XOR U953 ( .A(n1552), .B(n1553), .Z(n1551) );
  XNOR U954 ( .A(n1554), .B(n1555), .Z(n1553) );
  NOR U955 ( .A(n1556), .B(n1555), .Z(n1554) );
  XOR U956 ( .A(n1557), .B(n1558), .Z(n1552) );
  XOR U957 ( .A(n1559), .B(n1560), .Z(n1558) );
  XOR U958 ( .A(n1561), .B(n1562), .Z(n1560) );
  XNOR U959 ( .A(n1563), .B(n1564), .Z(n1562) );
  NOR U960 ( .A(n1565), .B(n1564), .Z(n1563) );
  XOR U961 ( .A(n1566), .B(n1567), .Z(n1561) );
  XOR U962 ( .A(n1568), .B(n1569), .Z(n1567) );
  XOR U963 ( .A(n1570), .B(n1571), .Z(n1569) );
  XNOR U964 ( .A(n1572), .B(n1573), .Z(n1571) );
  NOR U965 ( .A(n1574), .B(n1573), .Z(n1572) );
  XOR U966 ( .A(n1575), .B(n1576), .Z(n1570) );
  XOR U967 ( .A(n1577), .B(n1578), .Z(n1576) );
  XOR U968 ( .A(n1579), .B(n1580), .Z(n1578) );
  XNOR U969 ( .A(n1581), .B(n1582), .Z(n1580) );
  NOR U970 ( .A(n1583), .B(n1582), .Z(n1581) );
  XOR U971 ( .A(n1584), .B(n1585), .Z(n1579) );
  XOR U972 ( .A(n1586), .B(n1587), .Z(n1585) );
  XOR U973 ( .A(n1588), .B(n1589), .Z(n1587) );
  XNOR U974 ( .A(n1590), .B(n1591), .Z(n1589) );
  NOR U975 ( .A(n1592), .B(n1591), .Z(n1590) );
  XOR U976 ( .A(n1593), .B(n1594), .Z(n1588) );
  XOR U977 ( .A(n1595), .B(n1596), .Z(n1594) );
  XOR U978 ( .A(n1597), .B(n1598), .Z(n1596) );
  XNOR U979 ( .A(n1599), .B(n1600), .Z(n1598) );
  NOR U980 ( .A(n1601), .B(n1600), .Z(n1599) );
  XOR U981 ( .A(n1602), .B(n1603), .Z(n1597) );
  XOR U982 ( .A(n1604), .B(n1605), .Z(n1603) );
  XOR U983 ( .A(n1606), .B(n1607), .Z(n1605) );
  XNOR U984 ( .A(n1608), .B(n1609), .Z(n1607) );
  NOR U985 ( .A(n1610), .B(n1609), .Z(n1608) );
  XOR U986 ( .A(n1611), .B(n1612), .Z(n1606) );
  XOR U987 ( .A(n1613), .B(n1614), .Z(n1612) );
  XOR U988 ( .A(n1615), .B(n1616), .Z(n1614) );
  XNOR U989 ( .A(n1617), .B(n1618), .Z(n1616) );
  NOR U990 ( .A(n1619), .B(n1618), .Z(n1617) );
  XOR U991 ( .A(n1620), .B(n1621), .Z(n1615) );
  XOR U992 ( .A(n1622), .B(n1623), .Z(n1621) );
  XOR U993 ( .A(n1624), .B(n1625), .Z(n1623) );
  XNOR U994 ( .A(n1626), .B(n1627), .Z(n1625) );
  NOR U995 ( .A(n1628), .B(n1627), .Z(n1626) );
  XOR U996 ( .A(n1629), .B(n1630), .Z(n1624) );
  XOR U997 ( .A(n1631), .B(n1632), .Z(n1630) );
  XOR U998 ( .A(n1633), .B(n1634), .Z(n1632) );
  XNOR U999 ( .A(n1635), .B(n1636), .Z(n1634) );
  NOR U1000 ( .A(n1637), .B(n1636), .Z(n1635) );
  XOR U1001 ( .A(n1638), .B(n1639), .Z(n1633) );
  XOR U1002 ( .A(n1640), .B(n1641), .Z(n1639) );
  XOR U1003 ( .A(n1642), .B(n1643), .Z(n1641) );
  XNOR U1004 ( .A(n1644), .B(n1645), .Z(n1643) );
  NOR U1005 ( .A(n1646), .B(n1645), .Z(n1644) );
  XOR U1006 ( .A(n1647), .B(n1648), .Z(n1642) );
  XOR U1007 ( .A(n1649), .B(n1650), .Z(n1648) );
  XOR U1008 ( .A(n1651), .B(n1652), .Z(n1650) );
  XNOR U1009 ( .A(n1653), .B(n1654), .Z(n1652) );
  NOR U1010 ( .A(n1655), .B(n1654), .Z(n1653) );
  XOR U1011 ( .A(n1656), .B(n1657), .Z(n1651) );
  XOR U1012 ( .A(n1658), .B(n1659), .Z(n1657) );
  XOR U1013 ( .A(n1660), .B(n1661), .Z(n1659) );
  XNOR U1014 ( .A(n1662), .B(n1663), .Z(n1661) );
  NOR U1015 ( .A(n1664), .B(n1663), .Z(n1662) );
  XOR U1016 ( .A(n1665), .B(n1666), .Z(n1660) );
  XOR U1017 ( .A(n1667), .B(n1668), .Z(n1666) );
  XOR U1018 ( .A(n1669), .B(n1670), .Z(n1668) );
  XNOR U1019 ( .A(n1671), .B(n1672), .Z(n1670) );
  NOR U1020 ( .A(n1673), .B(n1672), .Z(n1671) );
  XOR U1021 ( .A(n1674), .B(n1675), .Z(n1669) );
  XOR U1022 ( .A(n1676), .B(n1677), .Z(n1675) );
  XOR U1023 ( .A(n1678), .B(n1679), .Z(n1677) );
  XNOR U1024 ( .A(n1680), .B(n1681), .Z(n1679) );
  NOR U1025 ( .A(n1682), .B(n1681), .Z(n1680) );
  XOR U1026 ( .A(n1683), .B(n1684), .Z(n1678) );
  XOR U1027 ( .A(n1685), .B(n1686), .Z(n1684) );
  XOR U1028 ( .A(n1687), .B(n1688), .Z(n1686) );
  XNOR U1029 ( .A(n1689), .B(n1690), .Z(n1688) );
  NOR U1030 ( .A(n1691), .B(n1690), .Z(n1689) );
  XOR U1031 ( .A(n1692), .B(n1693), .Z(n1687) );
  XOR U1032 ( .A(n1694), .B(n1695), .Z(n1693) );
  XOR U1033 ( .A(n1696), .B(n1697), .Z(n1695) );
  XNOR U1034 ( .A(n1698), .B(n1699), .Z(n1697) );
  NOR U1035 ( .A(n1700), .B(n1699), .Z(n1698) );
  XOR U1036 ( .A(n1701), .B(n1702), .Z(n1696) );
  XOR U1037 ( .A(n1703), .B(n1704), .Z(n1702) );
  XOR U1038 ( .A(n1705), .B(n1706), .Z(n1704) );
  XNOR U1039 ( .A(n1707), .B(n1708), .Z(n1706) );
  NOR U1040 ( .A(n1709), .B(n1708), .Z(n1707) );
  XOR U1041 ( .A(n1710), .B(n1711), .Z(n1705) );
  XOR U1042 ( .A(n1712), .B(n1713), .Z(n1711) );
  XOR U1043 ( .A(n1714), .B(n1715), .Z(n1713) );
  XNOR U1044 ( .A(n1716), .B(n1717), .Z(n1715) );
  NOR U1045 ( .A(n1718), .B(n1717), .Z(n1716) );
  XOR U1046 ( .A(n1719), .B(n1720), .Z(n1714) );
  XOR U1047 ( .A(n1721), .B(n1722), .Z(n1720) );
  XOR U1048 ( .A(n1723), .B(n1724), .Z(n1722) );
  XNOR U1049 ( .A(n1725), .B(n1726), .Z(n1724) );
  NOR U1050 ( .A(n1727), .B(n1726), .Z(n1725) );
  XOR U1051 ( .A(n1728), .B(n1729), .Z(n1723) );
  XOR U1052 ( .A(n1730), .B(n1731), .Z(n1729) );
  XOR U1053 ( .A(n1732), .B(n1733), .Z(n1731) );
  XNOR U1054 ( .A(n1734), .B(n1735), .Z(n1733) );
  NOR U1055 ( .A(n1736), .B(n1735), .Z(n1734) );
  XOR U1056 ( .A(n1737), .B(n1738), .Z(n1732) );
  XOR U1057 ( .A(n1739), .B(n1740), .Z(n1738) );
  XOR U1058 ( .A(n1741), .B(n1742), .Z(n1740) );
  XNOR U1059 ( .A(n1743), .B(n1744), .Z(n1742) );
  NOR U1060 ( .A(n1745), .B(n1744), .Z(n1743) );
  XOR U1061 ( .A(n1746), .B(n1747), .Z(n1741) );
  XOR U1062 ( .A(n1748), .B(n1749), .Z(n1747) );
  XOR U1063 ( .A(n1750), .B(n1751), .Z(n1749) );
  XNOR U1064 ( .A(n1752), .B(n1753), .Z(n1751) );
  NOR U1065 ( .A(n1754), .B(n1753), .Z(n1752) );
  XOR U1066 ( .A(n1755), .B(n1756), .Z(n1750) );
  XOR U1067 ( .A(n1757), .B(n1758), .Z(n1756) );
  XOR U1068 ( .A(n1759), .B(n1760), .Z(n1758) );
  XNOR U1069 ( .A(n1761), .B(n1762), .Z(n1760) );
  NOR U1070 ( .A(n1763), .B(n1762), .Z(n1761) );
  XOR U1071 ( .A(n1764), .B(n1765), .Z(n1759) );
  XOR U1072 ( .A(n1766), .B(n1767), .Z(n1765) );
  XOR U1073 ( .A(n1768), .B(n1769), .Z(n1767) );
  XNOR U1074 ( .A(n1770), .B(n1771), .Z(n1769) );
  NOR U1075 ( .A(n1772), .B(n1771), .Z(n1770) );
  XOR U1076 ( .A(n1773), .B(n1774), .Z(n1768) );
  XOR U1077 ( .A(n1775), .B(n1776), .Z(n1774) );
  XOR U1078 ( .A(n1777), .B(n1778), .Z(n1776) );
  XNOR U1079 ( .A(n1779), .B(n1780), .Z(n1778) );
  NOR U1080 ( .A(n1781), .B(n1780), .Z(n1779) );
  XOR U1081 ( .A(n1782), .B(n1783), .Z(n1777) );
  XOR U1082 ( .A(n1784), .B(n1785), .Z(n1783) );
  XOR U1083 ( .A(n1786), .B(n1787), .Z(n1785) );
  XNOR U1084 ( .A(n1788), .B(n1789), .Z(n1787) );
  NOR U1085 ( .A(n1790), .B(n1789), .Z(n1788) );
  XOR U1086 ( .A(n1791), .B(n1792), .Z(n1786) );
  XOR U1087 ( .A(n1793), .B(n1794), .Z(n1792) );
  XOR U1088 ( .A(n1795), .B(n1796), .Z(n1794) );
  XNOR U1089 ( .A(n1797), .B(n1798), .Z(n1796) );
  NOR U1090 ( .A(n1799), .B(n1798), .Z(n1797) );
  XOR U1091 ( .A(n1800), .B(n1801), .Z(n1795) );
  XOR U1092 ( .A(n1802), .B(n1803), .Z(n1801) );
  XOR U1093 ( .A(n1804), .B(n1805), .Z(n1803) );
  XNOR U1094 ( .A(n1806), .B(n1807), .Z(n1805) );
  NOR U1095 ( .A(n1808), .B(n1807), .Z(n1806) );
  XOR U1096 ( .A(n1809), .B(n1810), .Z(n1804) );
  XOR U1097 ( .A(n1811), .B(n1812), .Z(n1810) );
  XOR U1098 ( .A(n1813), .B(n1814), .Z(n1812) );
  XNOR U1099 ( .A(n1815), .B(n1816), .Z(n1814) );
  NOR U1100 ( .A(n1817), .B(n1816), .Z(n1815) );
  XOR U1101 ( .A(n1818), .B(n1819), .Z(n1813) );
  XOR U1102 ( .A(n1820), .B(n1821), .Z(n1819) );
  XOR U1103 ( .A(n1822), .B(n1823), .Z(n1821) );
  XNOR U1104 ( .A(n1824), .B(n1825), .Z(n1823) );
  NOR U1105 ( .A(n1826), .B(n1825), .Z(n1824) );
  XOR U1106 ( .A(n1827), .B(n1828), .Z(n1822) );
  XOR U1107 ( .A(n1829), .B(n1830), .Z(n1828) );
  XOR U1108 ( .A(n1831), .B(n1832), .Z(n1830) );
  XNOR U1109 ( .A(n1833), .B(n1834), .Z(n1832) );
  NOR U1110 ( .A(n1835), .B(n1834), .Z(n1833) );
  XOR U1111 ( .A(n1836), .B(n1837), .Z(n1831) );
  XOR U1112 ( .A(n1838), .B(n1839), .Z(n1837) );
  XOR U1113 ( .A(n1840), .B(n1841), .Z(n1839) );
  XNOR U1114 ( .A(n1842), .B(n1843), .Z(n1841) );
  NOR U1115 ( .A(n1844), .B(n1843), .Z(n1842) );
  XOR U1116 ( .A(n1845), .B(n1846), .Z(n1840) );
  XOR U1117 ( .A(n1847), .B(n1848), .Z(n1846) );
  XOR U1118 ( .A(n1849), .B(n1850), .Z(n1848) );
  XNOR U1119 ( .A(n1851), .B(n1852), .Z(n1850) );
  NOR U1120 ( .A(n1853), .B(n1852), .Z(n1851) );
  XOR U1121 ( .A(n1854), .B(n1855), .Z(n1849) );
  XOR U1122 ( .A(n1856), .B(n1857), .Z(n1855) );
  XOR U1123 ( .A(n1858), .B(n1859), .Z(n1857) );
  XNOR U1124 ( .A(n1860), .B(n1861), .Z(n1859) );
  NOR U1125 ( .A(n1862), .B(n1861), .Z(n1860) );
  XOR U1126 ( .A(n1863), .B(n1864), .Z(n1858) );
  XOR U1127 ( .A(n1865), .B(n1866), .Z(n1864) );
  XOR U1128 ( .A(n1867), .B(n1868), .Z(n1866) );
  XNOR U1129 ( .A(n1869), .B(n1870), .Z(n1868) );
  NOR U1130 ( .A(n1871), .B(n1870), .Z(n1869) );
  XOR U1131 ( .A(n1872), .B(n1873), .Z(n1867) );
  XOR U1132 ( .A(n1874), .B(n1875), .Z(n1873) );
  XOR U1133 ( .A(n1876), .B(n1877), .Z(n1875) );
  XNOR U1134 ( .A(n1878), .B(n1879), .Z(n1877) );
  NOR U1135 ( .A(n1880), .B(n1879), .Z(n1878) );
  XOR U1136 ( .A(n1881), .B(n1882), .Z(n1876) );
  XOR U1137 ( .A(n1883), .B(n1884), .Z(n1882) );
  XOR U1138 ( .A(n1885), .B(n1886), .Z(n1884) );
  XNOR U1139 ( .A(n1887), .B(n1888), .Z(n1886) );
  NOR U1140 ( .A(n1889), .B(n1888), .Z(n1887) );
  XOR U1141 ( .A(n1890), .B(n1891), .Z(n1885) );
  XOR U1142 ( .A(n1892), .B(n1893), .Z(n1891) );
  XOR U1143 ( .A(n1894), .B(n1895), .Z(n1893) );
  XNOR U1144 ( .A(n1896), .B(n1897), .Z(n1895) );
  NOR U1145 ( .A(n1898), .B(n1897), .Z(n1896) );
  XOR U1146 ( .A(n1899), .B(n1900), .Z(n1894) );
  XOR U1147 ( .A(n1901), .B(n1902), .Z(n1900) );
  XOR U1148 ( .A(n1903), .B(n1904), .Z(n1902) );
  XNOR U1149 ( .A(n1905), .B(n1906), .Z(n1904) );
  NOR U1150 ( .A(n1907), .B(n1906), .Z(n1905) );
  XOR U1151 ( .A(n1908), .B(n1909), .Z(n1903) );
  XOR U1152 ( .A(n1910), .B(n1911), .Z(n1909) );
  XOR U1153 ( .A(n1912), .B(n1913), .Z(n1911) );
  XNOR U1154 ( .A(n1914), .B(n1915), .Z(n1913) );
  NOR U1155 ( .A(n1916), .B(n1915), .Z(n1914) );
  XOR U1156 ( .A(n1917), .B(n1918), .Z(n1912) );
  XOR U1157 ( .A(n1919), .B(n1920), .Z(n1918) );
  XOR U1158 ( .A(n1921), .B(n1922), .Z(n1920) );
  XNOR U1159 ( .A(n1923), .B(n1924), .Z(n1922) );
  NOR U1160 ( .A(n1925), .B(n1924), .Z(n1923) );
  XOR U1161 ( .A(n1926), .B(n1927), .Z(n1921) );
  XOR U1162 ( .A(n1928), .B(n1929), .Z(n1927) );
  XOR U1163 ( .A(n1930), .B(n1931), .Z(n1929) );
  XNOR U1164 ( .A(n1932), .B(n1933), .Z(n1931) );
  NOR U1165 ( .A(n1934), .B(n1933), .Z(n1932) );
  XOR U1166 ( .A(n1935), .B(n1936), .Z(n1930) );
  XOR U1167 ( .A(n1937), .B(n1938), .Z(n1936) );
  XOR U1168 ( .A(n1939), .B(n1940), .Z(n1938) );
  XNOR U1169 ( .A(n1941), .B(n1942), .Z(n1940) );
  NOR U1170 ( .A(n1943), .B(n1942), .Z(n1941) );
  XOR U1171 ( .A(n1944), .B(n1945), .Z(n1939) );
  XOR U1172 ( .A(n1946), .B(n1947), .Z(n1945) );
  XOR U1173 ( .A(n1948), .B(n1949), .Z(n1947) );
  XNOR U1174 ( .A(n1950), .B(n1951), .Z(n1949) );
  NOR U1175 ( .A(n1952), .B(n1951), .Z(n1950) );
  XOR U1176 ( .A(n1953), .B(n1954), .Z(n1948) );
  XOR U1177 ( .A(n1955), .B(n1956), .Z(n1954) );
  XOR U1178 ( .A(n1957), .B(n1958), .Z(n1956) );
  XNOR U1179 ( .A(n1959), .B(n1960), .Z(n1958) );
  NOR U1180 ( .A(n1961), .B(n1960), .Z(n1959) );
  XOR U1181 ( .A(n1962), .B(n1963), .Z(n1957) );
  XOR U1182 ( .A(n1964), .B(n1965), .Z(n1963) );
  XOR U1183 ( .A(n1966), .B(n1967), .Z(n1965) );
  XNOR U1184 ( .A(n1968), .B(n1969), .Z(n1967) );
  NOR U1185 ( .A(n1970), .B(n1969), .Z(n1968) );
  XOR U1186 ( .A(n1971), .B(n1972), .Z(n1966) );
  XOR U1187 ( .A(n1973), .B(n1974), .Z(n1972) );
  XOR U1188 ( .A(n1975), .B(n1976), .Z(n1974) );
  XNOR U1189 ( .A(n1977), .B(n1978), .Z(n1976) );
  NOR U1190 ( .A(n1979), .B(n1978), .Z(n1977) );
  XOR U1191 ( .A(n1980), .B(n1981), .Z(n1975) );
  XOR U1192 ( .A(n1982), .B(n1983), .Z(n1981) );
  XOR U1193 ( .A(n1984), .B(n1985), .Z(n1983) );
  XNOR U1194 ( .A(n1986), .B(n1987), .Z(n1985) );
  NOR U1195 ( .A(n1988), .B(n1987), .Z(n1986) );
  XOR U1196 ( .A(n1989), .B(n1990), .Z(n1984) );
  XOR U1197 ( .A(n1991), .B(n1992), .Z(n1990) );
  XOR U1198 ( .A(n1993), .B(n1994), .Z(n1992) );
  XNOR U1199 ( .A(n1995), .B(n1996), .Z(n1994) );
  NOR U1200 ( .A(n1997), .B(n1996), .Z(n1995) );
  XOR U1201 ( .A(n1998), .B(n1999), .Z(n1993) );
  XOR U1202 ( .A(n2000), .B(n2001), .Z(n1999) );
  XOR U1203 ( .A(n2002), .B(n2003), .Z(n2001) );
  XNOR U1204 ( .A(n2004), .B(n2005), .Z(n2003) );
  NOR U1205 ( .A(n2006), .B(n2005), .Z(n2004) );
  XOR U1206 ( .A(n2007), .B(n2008), .Z(n2002) );
  XOR U1207 ( .A(n2009), .B(n2010), .Z(n2008) );
  XOR U1208 ( .A(n2011), .B(n2012), .Z(n2010) );
  XNOR U1209 ( .A(n2013), .B(n2014), .Z(n2012) );
  NOR U1210 ( .A(n2015), .B(n2014), .Z(n2013) );
  XOR U1211 ( .A(n2016), .B(n2017), .Z(n2011) );
  XOR U1212 ( .A(n2018), .B(n2019), .Z(n2017) );
  XOR U1213 ( .A(n2020), .B(n2021), .Z(n2019) );
  XOR U1214 ( .A(n2022), .B(n2023), .Z(n2018) );
  XNOR U1215 ( .A(n2024), .B(n2025), .Z(n2023) );
  XOR U1216 ( .A(n2026), .B(n2027), .Z(n2025) );
  XOR U1217 ( .A(n2028), .B(n2029), .Z(n2027) );
  XOR U1218 ( .A(n2030), .B(n2031), .Z(n2029) );
  XOR U1219 ( .A(n2032), .B(n2033), .Z(n2028) );
  XOR U1220 ( .A(n2034), .B(n2035), .Z(n2026) );
  XOR U1221 ( .A(n2036), .B(n2037), .Z(n2035) );
  AND U1222 ( .A(n2038), .B(n2039), .Z(n2037) );
  XNOR U1223 ( .A(n2040), .B(n2031), .Z(n2038) );
  XNOR U1224 ( .A(n2041), .B(n2042), .Z(n2031) );
  AND U1225 ( .A(n2040), .B(n2041), .Z(n2042) );
  NOR U1226 ( .A(n2043), .B(n2032), .Z(n2036) );
  XOR U1227 ( .A(n2044), .B(n2045), .Z(n2034) );
  NOR U1228 ( .A(n2046), .B(n2033), .Z(n2045) );
  NOR U1229 ( .A(n2047), .B(n2030), .Z(n2044) );
  XNOR U1230 ( .A(n2048), .B(n2049), .Z(n2022) );
  XNOR U1231 ( .A(n2050), .B(n2051), .Z(n2049) );
  NOR U1232 ( .A(n2052), .B(n2024), .Z(n2050) );
  XOR U1233 ( .A(n2053), .B(n2054), .Z(n2016) );
  XOR U1234 ( .A(n2055), .B(n2056), .Z(n2054) );
  NOR U1235 ( .A(n2057), .B(n2020), .Z(n2056) );
  NOR U1236 ( .A(n2058), .B(n2051), .Z(n2055) );
  XOR U1237 ( .A(n2059), .B(n2060), .Z(n2053) );
  NOR U1238 ( .A(n2061), .B(n2048), .Z(n2060) );
  NOR U1239 ( .A(n2062), .B(n2021), .Z(n2059) );
  XOR U1240 ( .A(n2063), .B(n2064), .Z(n2009) );
  XOR U1241 ( .A(n2065), .B(n2066), .Z(n2007) );
  XNOR U1242 ( .A(n2067), .B(n2068), .Z(n2066) );
  NOR U1243 ( .A(n2069), .B(n2068), .Z(n2067) );
  XOR U1244 ( .A(n2070), .B(n2071), .Z(n2065) );
  NOR U1245 ( .A(n2072), .B(n2063), .Z(n2071) );
  NOR U1246 ( .A(n2073), .B(n2064), .Z(n2070) );
  XOR U1247 ( .A(n2074), .B(n2075), .Z(n2000) );
  XOR U1248 ( .A(n2076), .B(n2077), .Z(n1998) );
  XNOR U1249 ( .A(n2078), .B(n2079), .Z(n2077) );
  NOR U1250 ( .A(n2080), .B(n2079), .Z(n2078) );
  XOR U1251 ( .A(n2081), .B(n2082), .Z(n2076) );
  NOR U1252 ( .A(n2083), .B(n2074), .Z(n2082) );
  NOR U1253 ( .A(n2084), .B(n2075), .Z(n2081) );
  XOR U1254 ( .A(n2085), .B(n2086), .Z(n1991) );
  XOR U1255 ( .A(n2087), .B(n2088), .Z(n1989) );
  XNOR U1256 ( .A(n2089), .B(n2090), .Z(n2088) );
  NOR U1257 ( .A(n2091), .B(n2090), .Z(n2089) );
  XOR U1258 ( .A(n2092), .B(n2093), .Z(n2087) );
  NOR U1259 ( .A(n2094), .B(n2085), .Z(n2093) );
  NOR U1260 ( .A(n2095), .B(n2086), .Z(n2092) );
  XOR U1261 ( .A(n2096), .B(n2097), .Z(n1982) );
  XOR U1262 ( .A(n2098), .B(n2099), .Z(n1980) );
  XNOR U1263 ( .A(n2100), .B(n2101), .Z(n2099) );
  NOR U1264 ( .A(n2102), .B(n2101), .Z(n2100) );
  XOR U1265 ( .A(n2103), .B(n2104), .Z(n2098) );
  NOR U1266 ( .A(n2105), .B(n2096), .Z(n2104) );
  NOR U1267 ( .A(n2106), .B(n2097), .Z(n2103) );
  XOR U1268 ( .A(n2107), .B(n2108), .Z(n1973) );
  XOR U1269 ( .A(n2109), .B(n2110), .Z(n1971) );
  XNOR U1270 ( .A(n2111), .B(n2112), .Z(n2110) );
  NOR U1271 ( .A(n2113), .B(n2112), .Z(n2111) );
  XOR U1272 ( .A(n2114), .B(n2115), .Z(n2109) );
  NOR U1273 ( .A(n2116), .B(n2107), .Z(n2115) );
  NOR U1274 ( .A(n2117), .B(n2108), .Z(n2114) );
  XOR U1275 ( .A(n2118), .B(n2119), .Z(n1964) );
  XOR U1276 ( .A(n2120), .B(n2121), .Z(n1962) );
  XNOR U1277 ( .A(n2122), .B(n2123), .Z(n2121) );
  NOR U1278 ( .A(n2124), .B(n2123), .Z(n2122) );
  XOR U1279 ( .A(n2125), .B(n2126), .Z(n2120) );
  NOR U1280 ( .A(n2127), .B(n2118), .Z(n2126) );
  NOR U1281 ( .A(n2128), .B(n2119), .Z(n2125) );
  XOR U1282 ( .A(n2129), .B(n2130), .Z(n1955) );
  XOR U1283 ( .A(n2131), .B(n2132), .Z(n1953) );
  XNOR U1284 ( .A(n2133), .B(n2134), .Z(n2132) );
  NOR U1285 ( .A(n2135), .B(n2134), .Z(n2133) );
  XOR U1286 ( .A(n2136), .B(n2137), .Z(n2131) );
  NOR U1287 ( .A(n2138), .B(n2129), .Z(n2137) );
  NOR U1288 ( .A(n2139), .B(n2130), .Z(n2136) );
  XOR U1289 ( .A(n2140), .B(n2141), .Z(n1946) );
  XOR U1290 ( .A(n2142), .B(n2143), .Z(n1944) );
  XNOR U1291 ( .A(n2144), .B(n2145), .Z(n2143) );
  NOR U1292 ( .A(n2146), .B(n2145), .Z(n2144) );
  XOR U1293 ( .A(n2147), .B(n2148), .Z(n2142) );
  NOR U1294 ( .A(n2149), .B(n2140), .Z(n2148) );
  NOR U1295 ( .A(n2150), .B(n2141), .Z(n2147) );
  XOR U1296 ( .A(n2151), .B(n2152), .Z(n1937) );
  XOR U1297 ( .A(n2153), .B(n2154), .Z(n1935) );
  XNOR U1298 ( .A(n2155), .B(n2156), .Z(n2154) );
  NOR U1299 ( .A(n2157), .B(n2156), .Z(n2155) );
  XOR U1300 ( .A(n2158), .B(n2159), .Z(n2153) );
  NOR U1301 ( .A(n2160), .B(n2151), .Z(n2159) );
  NOR U1302 ( .A(n2161), .B(n2152), .Z(n2158) );
  XOR U1303 ( .A(n2162), .B(n2163), .Z(n1928) );
  XOR U1304 ( .A(n2164), .B(n2165), .Z(n1926) );
  XNOR U1305 ( .A(n2166), .B(n2167), .Z(n2165) );
  NOR U1306 ( .A(n2168), .B(n2167), .Z(n2166) );
  XOR U1307 ( .A(n2169), .B(n2170), .Z(n2164) );
  NOR U1308 ( .A(n2171), .B(n2162), .Z(n2170) );
  NOR U1309 ( .A(n2172), .B(n2163), .Z(n2169) );
  XOR U1310 ( .A(n2173), .B(n2174), .Z(n1919) );
  XOR U1311 ( .A(n2175), .B(n2176), .Z(n1917) );
  XNOR U1312 ( .A(n2177), .B(n2178), .Z(n2176) );
  NOR U1313 ( .A(n2179), .B(n2178), .Z(n2177) );
  XOR U1314 ( .A(n2180), .B(n2181), .Z(n2175) );
  NOR U1315 ( .A(n2182), .B(n2173), .Z(n2181) );
  NOR U1316 ( .A(n2183), .B(n2174), .Z(n2180) );
  XOR U1317 ( .A(n2184), .B(n2185), .Z(n1910) );
  XOR U1318 ( .A(n2186), .B(n2187), .Z(n1908) );
  XNOR U1319 ( .A(n2188), .B(n2189), .Z(n2187) );
  NOR U1320 ( .A(n2190), .B(n2189), .Z(n2188) );
  XOR U1321 ( .A(n2191), .B(n2192), .Z(n2186) );
  NOR U1322 ( .A(n2193), .B(n2184), .Z(n2192) );
  NOR U1323 ( .A(n2194), .B(n2185), .Z(n2191) );
  XOR U1324 ( .A(n2195), .B(n2196), .Z(n1901) );
  XOR U1325 ( .A(n2197), .B(n2198), .Z(n1899) );
  XNOR U1326 ( .A(n2199), .B(n2200), .Z(n2198) );
  NOR U1327 ( .A(n2201), .B(n2200), .Z(n2199) );
  XOR U1328 ( .A(n2202), .B(n2203), .Z(n2197) );
  NOR U1329 ( .A(n2204), .B(n2195), .Z(n2203) );
  NOR U1330 ( .A(n2205), .B(n2196), .Z(n2202) );
  XOR U1331 ( .A(n2206), .B(n2207), .Z(n1892) );
  XOR U1332 ( .A(n2208), .B(n2209), .Z(n1890) );
  XNOR U1333 ( .A(n2210), .B(n2211), .Z(n2209) );
  NOR U1334 ( .A(n2212), .B(n2211), .Z(n2210) );
  XOR U1335 ( .A(n2213), .B(n2214), .Z(n2208) );
  NOR U1336 ( .A(n2215), .B(n2206), .Z(n2214) );
  NOR U1337 ( .A(n2216), .B(n2207), .Z(n2213) );
  XOR U1338 ( .A(n2217), .B(n2218), .Z(n1883) );
  XOR U1339 ( .A(n2219), .B(n2220), .Z(n1881) );
  XNOR U1340 ( .A(n2221), .B(n2222), .Z(n2220) );
  NOR U1341 ( .A(n2223), .B(n2222), .Z(n2221) );
  XOR U1342 ( .A(n2224), .B(n2225), .Z(n2219) );
  NOR U1343 ( .A(n2226), .B(n2217), .Z(n2225) );
  NOR U1344 ( .A(n2227), .B(n2218), .Z(n2224) );
  XOR U1345 ( .A(n2228), .B(n2229), .Z(n1874) );
  XOR U1346 ( .A(n2230), .B(n2231), .Z(n1872) );
  XNOR U1347 ( .A(n2232), .B(n2233), .Z(n2231) );
  NOR U1348 ( .A(n2234), .B(n2233), .Z(n2232) );
  XOR U1349 ( .A(n2235), .B(n2236), .Z(n2230) );
  NOR U1350 ( .A(n2237), .B(n2228), .Z(n2236) );
  NOR U1351 ( .A(n2238), .B(n2229), .Z(n2235) );
  XOR U1352 ( .A(n2239), .B(n2240), .Z(n1865) );
  XOR U1353 ( .A(n2241), .B(n2242), .Z(n1863) );
  XNOR U1354 ( .A(n2243), .B(n2244), .Z(n2242) );
  NOR U1355 ( .A(n2245), .B(n2244), .Z(n2243) );
  XOR U1356 ( .A(n2246), .B(n2247), .Z(n2241) );
  NOR U1357 ( .A(n2248), .B(n2239), .Z(n2247) );
  NOR U1358 ( .A(n2249), .B(n2240), .Z(n2246) );
  XOR U1359 ( .A(n2250), .B(n2251), .Z(n1856) );
  XOR U1360 ( .A(n2252), .B(n2253), .Z(n1854) );
  XNOR U1361 ( .A(n2254), .B(n2255), .Z(n2253) );
  NOR U1362 ( .A(n2256), .B(n2255), .Z(n2254) );
  XOR U1363 ( .A(n2257), .B(n2258), .Z(n2252) );
  NOR U1364 ( .A(n2259), .B(n2250), .Z(n2258) );
  NOR U1365 ( .A(n2260), .B(n2251), .Z(n2257) );
  XOR U1366 ( .A(n2261), .B(n2262), .Z(n1847) );
  XOR U1367 ( .A(n2263), .B(n2264), .Z(n1845) );
  XNOR U1368 ( .A(n2265), .B(n2266), .Z(n2264) );
  NOR U1369 ( .A(n2267), .B(n2266), .Z(n2265) );
  XOR U1370 ( .A(n2268), .B(n2269), .Z(n2263) );
  NOR U1371 ( .A(n2270), .B(n2261), .Z(n2269) );
  NOR U1372 ( .A(n2271), .B(n2262), .Z(n2268) );
  XOR U1373 ( .A(n2272), .B(n2273), .Z(n1838) );
  XOR U1374 ( .A(n2274), .B(n2275), .Z(n1836) );
  XNOR U1375 ( .A(n2276), .B(n2277), .Z(n2275) );
  NOR U1376 ( .A(n2278), .B(n2277), .Z(n2276) );
  XOR U1377 ( .A(n2279), .B(n2280), .Z(n2274) );
  NOR U1378 ( .A(n2281), .B(n2272), .Z(n2280) );
  NOR U1379 ( .A(n2282), .B(n2273), .Z(n2279) );
  XOR U1380 ( .A(n2283), .B(n2284), .Z(n1829) );
  XOR U1381 ( .A(n2285), .B(n2286), .Z(n1827) );
  XNOR U1382 ( .A(n2287), .B(n2288), .Z(n2286) );
  NOR U1383 ( .A(n2289), .B(n2288), .Z(n2287) );
  XOR U1384 ( .A(n2290), .B(n2291), .Z(n2285) );
  NOR U1385 ( .A(n2292), .B(n2283), .Z(n2291) );
  NOR U1386 ( .A(n2293), .B(n2284), .Z(n2290) );
  XOR U1387 ( .A(n2294), .B(n2295), .Z(n1820) );
  XOR U1388 ( .A(n2296), .B(n2297), .Z(n1818) );
  XNOR U1389 ( .A(n2298), .B(n2299), .Z(n2297) );
  NOR U1390 ( .A(n2300), .B(n2299), .Z(n2298) );
  XOR U1391 ( .A(n2301), .B(n2302), .Z(n2296) );
  NOR U1392 ( .A(n2303), .B(n2294), .Z(n2302) );
  NOR U1393 ( .A(n2304), .B(n2295), .Z(n2301) );
  XOR U1394 ( .A(n2305), .B(n2306), .Z(n1811) );
  XOR U1395 ( .A(n2307), .B(n2308), .Z(n1809) );
  XNOR U1396 ( .A(n2309), .B(n2310), .Z(n2308) );
  NOR U1397 ( .A(n2311), .B(n2310), .Z(n2309) );
  XOR U1398 ( .A(n2312), .B(n2313), .Z(n2307) );
  NOR U1399 ( .A(n2314), .B(n2305), .Z(n2313) );
  NOR U1400 ( .A(n2315), .B(n2306), .Z(n2312) );
  XOR U1401 ( .A(n2316), .B(n2317), .Z(n1802) );
  XOR U1402 ( .A(n2318), .B(n2319), .Z(n1800) );
  XNOR U1403 ( .A(n2320), .B(n2321), .Z(n2319) );
  NOR U1404 ( .A(n2322), .B(n2321), .Z(n2320) );
  XOR U1405 ( .A(n2323), .B(n2324), .Z(n2318) );
  NOR U1406 ( .A(n2325), .B(n2316), .Z(n2324) );
  NOR U1407 ( .A(n2326), .B(n2317), .Z(n2323) );
  XOR U1408 ( .A(n2327), .B(n2328), .Z(n1793) );
  XOR U1409 ( .A(n2329), .B(n2330), .Z(n1791) );
  XNOR U1410 ( .A(n2331), .B(n2332), .Z(n2330) );
  NOR U1411 ( .A(n2333), .B(n2332), .Z(n2331) );
  XOR U1412 ( .A(n2334), .B(n2335), .Z(n2329) );
  NOR U1413 ( .A(n2336), .B(n2327), .Z(n2335) );
  NOR U1414 ( .A(n2337), .B(n2328), .Z(n2334) );
  XOR U1415 ( .A(n2338), .B(n2339), .Z(n1784) );
  XOR U1416 ( .A(n2340), .B(n2341), .Z(n1782) );
  XNOR U1417 ( .A(n2342), .B(n2343), .Z(n2341) );
  NOR U1418 ( .A(n2344), .B(n2343), .Z(n2342) );
  XOR U1419 ( .A(n2345), .B(n2346), .Z(n2340) );
  NOR U1420 ( .A(n2347), .B(n2338), .Z(n2346) );
  NOR U1421 ( .A(n2348), .B(n2339), .Z(n2345) );
  XOR U1422 ( .A(n2349), .B(n2350), .Z(n1775) );
  XOR U1423 ( .A(n2351), .B(n2352), .Z(n1773) );
  XNOR U1424 ( .A(n2353), .B(n2354), .Z(n2352) );
  NOR U1425 ( .A(n2355), .B(n2354), .Z(n2353) );
  XOR U1426 ( .A(n2356), .B(n2357), .Z(n2351) );
  NOR U1427 ( .A(n2358), .B(n2349), .Z(n2357) );
  NOR U1428 ( .A(n2359), .B(n2350), .Z(n2356) );
  XOR U1429 ( .A(n2360), .B(n2361), .Z(n1766) );
  XOR U1430 ( .A(n2362), .B(n2363), .Z(n1764) );
  XNOR U1431 ( .A(n2364), .B(n2365), .Z(n2363) );
  NOR U1432 ( .A(n2366), .B(n2365), .Z(n2364) );
  XOR U1433 ( .A(n2367), .B(n2368), .Z(n2362) );
  NOR U1434 ( .A(n2369), .B(n2360), .Z(n2368) );
  NOR U1435 ( .A(n2370), .B(n2361), .Z(n2367) );
  XOR U1436 ( .A(n2371), .B(n2372), .Z(n1757) );
  XOR U1437 ( .A(n2373), .B(n2374), .Z(n1755) );
  XNOR U1438 ( .A(n2375), .B(n2376), .Z(n2374) );
  NOR U1439 ( .A(n2377), .B(n2376), .Z(n2375) );
  XOR U1440 ( .A(n2378), .B(n2379), .Z(n2373) );
  NOR U1441 ( .A(n2380), .B(n2371), .Z(n2379) );
  NOR U1442 ( .A(n2381), .B(n2372), .Z(n2378) );
  XOR U1443 ( .A(n2382), .B(n2383), .Z(n1748) );
  XOR U1444 ( .A(n2384), .B(n2385), .Z(n1746) );
  XNOR U1445 ( .A(n2386), .B(n2387), .Z(n2385) );
  NOR U1446 ( .A(n2388), .B(n2387), .Z(n2386) );
  XOR U1447 ( .A(n2389), .B(n2390), .Z(n2384) );
  NOR U1448 ( .A(n2391), .B(n2382), .Z(n2390) );
  NOR U1449 ( .A(n2392), .B(n2383), .Z(n2389) );
  XOR U1450 ( .A(n2393), .B(n2394), .Z(n1739) );
  XOR U1451 ( .A(n2395), .B(n2396), .Z(n1737) );
  XNOR U1452 ( .A(n2397), .B(n2398), .Z(n2396) );
  NOR U1453 ( .A(n2399), .B(n2398), .Z(n2397) );
  XOR U1454 ( .A(n2400), .B(n2401), .Z(n2395) );
  NOR U1455 ( .A(n2402), .B(n2393), .Z(n2401) );
  NOR U1456 ( .A(n2403), .B(n2394), .Z(n2400) );
  XOR U1457 ( .A(n2404), .B(n2405), .Z(n1730) );
  XOR U1458 ( .A(n2406), .B(n2407), .Z(n1728) );
  XNOR U1459 ( .A(n2408), .B(n2409), .Z(n2407) );
  NOR U1460 ( .A(n2410), .B(n2409), .Z(n2408) );
  XOR U1461 ( .A(n2411), .B(n2412), .Z(n2406) );
  NOR U1462 ( .A(n2413), .B(n2404), .Z(n2412) );
  NOR U1463 ( .A(n2414), .B(n2405), .Z(n2411) );
  XOR U1464 ( .A(n2415), .B(n2416), .Z(n1721) );
  XOR U1465 ( .A(n2417), .B(n2418), .Z(n1719) );
  XNOR U1466 ( .A(n2419), .B(n2420), .Z(n2418) );
  NOR U1467 ( .A(n2421), .B(n2420), .Z(n2419) );
  XOR U1468 ( .A(n2422), .B(n2423), .Z(n2417) );
  NOR U1469 ( .A(n2424), .B(n2415), .Z(n2423) );
  NOR U1470 ( .A(n2425), .B(n2416), .Z(n2422) );
  XOR U1471 ( .A(n2426), .B(n2427), .Z(n1712) );
  XOR U1472 ( .A(n2428), .B(n2429), .Z(n1710) );
  XNOR U1473 ( .A(n2430), .B(n2431), .Z(n2429) );
  NOR U1474 ( .A(n2432), .B(n2431), .Z(n2430) );
  XOR U1475 ( .A(n2433), .B(n2434), .Z(n2428) );
  NOR U1476 ( .A(n2435), .B(n2426), .Z(n2434) );
  NOR U1477 ( .A(n2436), .B(n2427), .Z(n2433) );
  XOR U1478 ( .A(n2437), .B(n2438), .Z(n1703) );
  XOR U1479 ( .A(n2439), .B(n2440), .Z(n1701) );
  XNOR U1480 ( .A(n2441), .B(n2442), .Z(n2440) );
  NOR U1481 ( .A(n2443), .B(n2442), .Z(n2441) );
  XOR U1482 ( .A(n2444), .B(n2445), .Z(n2439) );
  NOR U1483 ( .A(n2446), .B(n2437), .Z(n2445) );
  NOR U1484 ( .A(n2447), .B(n2438), .Z(n2444) );
  XOR U1485 ( .A(n2448), .B(n2449), .Z(n1694) );
  XOR U1486 ( .A(n2450), .B(n2451), .Z(n1692) );
  XNOR U1487 ( .A(n2452), .B(n2453), .Z(n2451) );
  NOR U1488 ( .A(n2454), .B(n2453), .Z(n2452) );
  XOR U1489 ( .A(n2455), .B(n2456), .Z(n2450) );
  NOR U1490 ( .A(n2457), .B(n2448), .Z(n2456) );
  NOR U1491 ( .A(n2458), .B(n2449), .Z(n2455) );
  XOR U1492 ( .A(n2459), .B(n2460), .Z(n1685) );
  XOR U1493 ( .A(n2461), .B(n2462), .Z(n1683) );
  XNOR U1494 ( .A(n2463), .B(n2464), .Z(n2462) );
  NOR U1495 ( .A(n2465), .B(n2464), .Z(n2463) );
  XOR U1496 ( .A(n2466), .B(n2467), .Z(n2461) );
  NOR U1497 ( .A(n2468), .B(n2459), .Z(n2467) );
  NOR U1498 ( .A(n2469), .B(n2460), .Z(n2466) );
  XOR U1499 ( .A(n2470), .B(n2471), .Z(n1676) );
  XOR U1500 ( .A(n2472), .B(n2473), .Z(n1674) );
  XNOR U1501 ( .A(n2474), .B(n2475), .Z(n2473) );
  NOR U1502 ( .A(n2476), .B(n2475), .Z(n2474) );
  XOR U1503 ( .A(n2477), .B(n2478), .Z(n2472) );
  NOR U1504 ( .A(n2479), .B(n2470), .Z(n2478) );
  NOR U1505 ( .A(n2480), .B(n2471), .Z(n2477) );
  XOR U1506 ( .A(n2481), .B(n2482), .Z(n1667) );
  XOR U1507 ( .A(n2483), .B(n2484), .Z(n1665) );
  XNOR U1508 ( .A(n2485), .B(n2486), .Z(n2484) );
  NOR U1509 ( .A(n2487), .B(n2486), .Z(n2485) );
  XOR U1510 ( .A(n2488), .B(n2489), .Z(n2483) );
  NOR U1511 ( .A(n2490), .B(n2481), .Z(n2489) );
  NOR U1512 ( .A(n2491), .B(n2482), .Z(n2488) );
  XOR U1513 ( .A(n2492), .B(n2493), .Z(n1658) );
  XOR U1514 ( .A(n2494), .B(n2495), .Z(n1656) );
  XNOR U1515 ( .A(n2496), .B(n2497), .Z(n2495) );
  NOR U1516 ( .A(n2498), .B(n2497), .Z(n2496) );
  XOR U1517 ( .A(n2499), .B(n2500), .Z(n2494) );
  NOR U1518 ( .A(n2501), .B(n2492), .Z(n2500) );
  NOR U1519 ( .A(n2502), .B(n2493), .Z(n2499) );
  XOR U1520 ( .A(n2503), .B(n2504), .Z(n1649) );
  XOR U1521 ( .A(n2505), .B(n2506), .Z(n1647) );
  XNOR U1522 ( .A(n2507), .B(n2508), .Z(n2506) );
  NOR U1523 ( .A(n2509), .B(n2508), .Z(n2507) );
  XOR U1524 ( .A(n2510), .B(n2511), .Z(n2505) );
  NOR U1525 ( .A(n2512), .B(n2503), .Z(n2511) );
  NOR U1526 ( .A(n2513), .B(n2504), .Z(n2510) );
  XOR U1527 ( .A(n2514), .B(n2515), .Z(n1640) );
  XOR U1528 ( .A(n2516), .B(n2517), .Z(n1638) );
  XNOR U1529 ( .A(n2518), .B(n2519), .Z(n2517) );
  NOR U1530 ( .A(n2520), .B(n2519), .Z(n2518) );
  XOR U1531 ( .A(n2521), .B(n2522), .Z(n2516) );
  NOR U1532 ( .A(n2523), .B(n2514), .Z(n2522) );
  NOR U1533 ( .A(n2524), .B(n2515), .Z(n2521) );
  XOR U1534 ( .A(n2525), .B(n2526), .Z(n1631) );
  XOR U1535 ( .A(n2527), .B(n2528), .Z(n1629) );
  XNOR U1536 ( .A(n2529), .B(n2530), .Z(n2528) );
  NOR U1537 ( .A(n2531), .B(n2530), .Z(n2529) );
  XOR U1538 ( .A(n2532), .B(n2533), .Z(n2527) );
  NOR U1539 ( .A(n2534), .B(n2525), .Z(n2533) );
  NOR U1540 ( .A(n2535), .B(n2526), .Z(n2532) );
  XOR U1541 ( .A(n2536), .B(n2537), .Z(n1622) );
  XOR U1542 ( .A(n2538), .B(n2539), .Z(n1620) );
  XNOR U1543 ( .A(n2540), .B(n2541), .Z(n2539) );
  NOR U1544 ( .A(n2542), .B(n2541), .Z(n2540) );
  XOR U1545 ( .A(n2543), .B(n2544), .Z(n2538) );
  NOR U1546 ( .A(n2545), .B(n2536), .Z(n2544) );
  NOR U1547 ( .A(n2546), .B(n2537), .Z(n2543) );
  XOR U1548 ( .A(n2547), .B(n2548), .Z(n1613) );
  XOR U1549 ( .A(n2549), .B(n2550), .Z(n1611) );
  XNOR U1550 ( .A(n2551), .B(n2552), .Z(n2550) );
  NOR U1551 ( .A(n2553), .B(n2552), .Z(n2551) );
  XOR U1552 ( .A(n2554), .B(n2555), .Z(n2549) );
  NOR U1553 ( .A(n2556), .B(n2547), .Z(n2555) );
  NOR U1554 ( .A(n2557), .B(n2548), .Z(n2554) );
  XOR U1555 ( .A(n2558), .B(n2559), .Z(n1604) );
  XOR U1556 ( .A(n2560), .B(n2561), .Z(n1602) );
  XNOR U1557 ( .A(n2562), .B(n2563), .Z(n2561) );
  NOR U1558 ( .A(n2564), .B(n2563), .Z(n2562) );
  XOR U1559 ( .A(n2565), .B(n2566), .Z(n2560) );
  NOR U1560 ( .A(n2567), .B(n2558), .Z(n2566) );
  NOR U1561 ( .A(n2568), .B(n2559), .Z(n2565) );
  XOR U1562 ( .A(n2569), .B(n2570), .Z(n1595) );
  XOR U1563 ( .A(n2571), .B(n2572), .Z(n1593) );
  XNOR U1564 ( .A(n2573), .B(n2574), .Z(n2572) );
  NOR U1565 ( .A(n2575), .B(n2574), .Z(n2573) );
  XOR U1566 ( .A(n2576), .B(n2577), .Z(n2571) );
  NOR U1567 ( .A(n2578), .B(n2569), .Z(n2577) );
  NOR U1568 ( .A(n2579), .B(n2570), .Z(n2576) );
  XOR U1569 ( .A(n2580), .B(n2581), .Z(n1586) );
  XOR U1570 ( .A(n2582), .B(n2583), .Z(n1584) );
  XNOR U1571 ( .A(n2584), .B(n2585), .Z(n2583) );
  NOR U1572 ( .A(n2586), .B(n2585), .Z(n2584) );
  XOR U1573 ( .A(n2587), .B(n2588), .Z(n2582) );
  NOR U1574 ( .A(n2589), .B(n2580), .Z(n2588) );
  NOR U1575 ( .A(n2590), .B(n2581), .Z(n2587) );
  XOR U1576 ( .A(n2591), .B(n2592), .Z(n1577) );
  XOR U1577 ( .A(n2593), .B(n2594), .Z(n1575) );
  XNOR U1578 ( .A(n2595), .B(n2596), .Z(n2594) );
  NOR U1579 ( .A(n2597), .B(n2596), .Z(n2595) );
  XOR U1580 ( .A(n2598), .B(n2599), .Z(n2593) );
  NOR U1581 ( .A(n2600), .B(n2591), .Z(n2599) );
  NOR U1582 ( .A(n2601), .B(n2592), .Z(n2598) );
  XOR U1583 ( .A(n2602), .B(n2603), .Z(n1568) );
  XOR U1584 ( .A(n2604), .B(n2605), .Z(n1566) );
  XNOR U1585 ( .A(n2606), .B(n2607), .Z(n2605) );
  NOR U1586 ( .A(n2608), .B(n2607), .Z(n2606) );
  XOR U1587 ( .A(n2609), .B(n2610), .Z(n2604) );
  NOR U1588 ( .A(n2611), .B(n2602), .Z(n2610) );
  NOR U1589 ( .A(n2612), .B(n2603), .Z(n2609) );
  XOR U1590 ( .A(n2613), .B(n2614), .Z(n1559) );
  XOR U1591 ( .A(n2615), .B(n2616), .Z(n1557) );
  XNOR U1592 ( .A(n2617), .B(n2618), .Z(n2616) );
  NOR U1593 ( .A(n2619), .B(n2618), .Z(n2617) );
  XOR U1594 ( .A(n2620), .B(n2621), .Z(n2615) );
  NOR U1595 ( .A(n2622), .B(n2613), .Z(n2621) );
  NOR U1596 ( .A(n2623), .B(n2614), .Z(n2620) );
  XOR U1597 ( .A(n2624), .B(n2625), .Z(n1550) );
  XOR U1598 ( .A(n2626), .B(n2627), .Z(n1548) );
  XNOR U1599 ( .A(n2628), .B(n2629), .Z(n2627) );
  NOR U1600 ( .A(n2630), .B(n2629), .Z(n2628) );
  XOR U1601 ( .A(n2631), .B(n2632), .Z(n2626) );
  NOR U1602 ( .A(n2633), .B(n2624), .Z(n2632) );
  NOR U1603 ( .A(n2634), .B(n2625), .Z(n2631) );
  XOR U1604 ( .A(n2635), .B(n2636), .Z(n1541) );
  XOR U1605 ( .A(n2637), .B(n2638), .Z(n1539) );
  XNOR U1606 ( .A(n2639), .B(n2640), .Z(n2638) );
  NOR U1607 ( .A(n2641), .B(n2640), .Z(n2639) );
  XOR U1608 ( .A(n2642), .B(n2643), .Z(n2637) );
  NOR U1609 ( .A(n2644), .B(n2635), .Z(n2643) );
  NOR U1610 ( .A(n2645), .B(n2636), .Z(n2642) );
  XOR U1611 ( .A(n2646), .B(n2647), .Z(n1532) );
  XOR U1612 ( .A(n2648), .B(n2649), .Z(n1530) );
  XNOR U1613 ( .A(n2650), .B(n2651), .Z(n2649) );
  NOR U1614 ( .A(n2652), .B(n2651), .Z(n2650) );
  XOR U1615 ( .A(n2653), .B(n2654), .Z(n2648) );
  NOR U1616 ( .A(n2655), .B(n2646), .Z(n2654) );
  NOR U1617 ( .A(n2656), .B(n2647), .Z(n2653) );
  XOR U1618 ( .A(n2657), .B(n2658), .Z(n1523) );
  XOR U1619 ( .A(n2659), .B(n2660), .Z(n1521) );
  XNOR U1620 ( .A(n2661), .B(n2662), .Z(n2660) );
  NOR U1621 ( .A(n2663), .B(n2662), .Z(n2661) );
  XOR U1622 ( .A(n2664), .B(n2665), .Z(n2659) );
  NOR U1623 ( .A(n2666), .B(n2657), .Z(n2665) );
  NOR U1624 ( .A(n2667), .B(n2658), .Z(n2664) );
  XOR U1625 ( .A(n2668), .B(n2669), .Z(n1514) );
  XOR U1626 ( .A(n2670), .B(n2671), .Z(n1512) );
  XNOR U1627 ( .A(n2672), .B(n2673), .Z(n2671) );
  NOR U1628 ( .A(n2674), .B(n2673), .Z(n2672) );
  XOR U1629 ( .A(n2675), .B(n2676), .Z(n2670) );
  NOR U1630 ( .A(n2677), .B(n2668), .Z(n2676) );
  NOR U1631 ( .A(n2678), .B(n2669), .Z(n2675) );
  XOR U1632 ( .A(n2679), .B(n2680), .Z(n1505) );
  XOR U1633 ( .A(n2681), .B(n2682), .Z(n1503) );
  XNOR U1634 ( .A(n2683), .B(n2684), .Z(n2682) );
  NOR U1635 ( .A(n2685), .B(n2684), .Z(n2683) );
  XOR U1636 ( .A(n2686), .B(n2687), .Z(n2681) );
  NOR U1637 ( .A(n2688), .B(n2679), .Z(n2687) );
  NOR U1638 ( .A(n2689), .B(n2680), .Z(n2686) );
  XOR U1639 ( .A(n2690), .B(n2691), .Z(n1496) );
  XOR U1640 ( .A(n2692), .B(n2693), .Z(n1494) );
  XNOR U1641 ( .A(n2694), .B(n2695), .Z(n2693) );
  NOR U1642 ( .A(n2696), .B(n2695), .Z(n2694) );
  XOR U1643 ( .A(n2697), .B(n2698), .Z(n2692) );
  NOR U1644 ( .A(n2699), .B(n2690), .Z(n2698) );
  NOR U1645 ( .A(n2700), .B(n2691), .Z(n2697) );
  XOR U1646 ( .A(n2701), .B(n2702), .Z(n1487) );
  XOR U1647 ( .A(n2703), .B(n2704), .Z(n1485) );
  XNOR U1648 ( .A(n2705), .B(n2706), .Z(n2704) );
  NOR U1649 ( .A(n2707), .B(n2706), .Z(n2705) );
  XOR U1650 ( .A(n2708), .B(n2709), .Z(n2703) );
  NOR U1651 ( .A(n2710), .B(n2701), .Z(n2709) );
  NOR U1652 ( .A(n2711), .B(n2702), .Z(n2708) );
  XOR U1653 ( .A(n2712), .B(n2713), .Z(n1478) );
  XOR U1654 ( .A(n2714), .B(n2715), .Z(n1476) );
  XNOR U1655 ( .A(n2716), .B(n2717), .Z(n2715) );
  NOR U1656 ( .A(n2718), .B(n2717), .Z(n2716) );
  XOR U1657 ( .A(n2719), .B(n2720), .Z(n2714) );
  NOR U1658 ( .A(n2721), .B(n2712), .Z(n2720) );
  NOR U1659 ( .A(n2722), .B(n2713), .Z(n2719) );
  XOR U1660 ( .A(n2723), .B(n2724), .Z(n1469) );
  XOR U1661 ( .A(n2725), .B(n2726), .Z(n1467) );
  XNOR U1662 ( .A(n2727), .B(n2728), .Z(n2726) );
  NOR U1663 ( .A(n2729), .B(n2728), .Z(n2727) );
  XOR U1664 ( .A(n2730), .B(n2731), .Z(n2725) );
  NOR U1665 ( .A(n2732), .B(n2723), .Z(n2731) );
  NOR U1666 ( .A(n2733), .B(n2724), .Z(n2730) );
  XOR U1667 ( .A(n1464), .B(n1462), .Z(n1465) );
  XOR U1668 ( .A(n2734), .B(n2735), .Z(n161) );
  NOR U1669 ( .A(n42), .B(n2736), .Z(n2735) );
  IV U1670 ( .A(n2734), .Z(n2736) );
  IV U1671 ( .A(n45), .Z(n42) );
  XOR U1672 ( .A(n2737), .B(n2738), .Z(n164) );
  AND U1673 ( .A(n2739), .B(n2740), .Z(n2738) );
  XNOR U1674 ( .A(n2737), .B(n44), .Z(n2740) );
  XNOR U1675 ( .A(n1450), .B(n180), .Z(n44) );
  XNOR U1676 ( .A(n181), .B(n178), .Z(n180) );
  XNOR U1677 ( .A(n179), .B(n174), .Z(n178) );
  XOR U1678 ( .A(n175), .B(n195), .Z(n174) );
  XOR U1679 ( .A(n2741), .B(n193), .Z(n195) );
  XNOR U1680 ( .A(n194), .B(n1448), .Z(n193) );
  XNOR U1681 ( .A(n1449), .B(n1447), .Z(n1448) );
  XNOR U1682 ( .A(n190), .B(n1444), .Z(n1447) );
  XNOR U1683 ( .A(n189), .B(n212), .Z(n1444) );
  XNOR U1684 ( .A(n207), .B(n1443), .Z(n212) );
  XNOR U1685 ( .A(n206), .B(n1438), .Z(n1443) );
  XNOR U1686 ( .A(n208), .B(n1437), .Z(n1438) );
  XNOR U1687 ( .A(n211), .B(n1434), .Z(n1437) );
  XNOR U1688 ( .A(n217), .B(n1433), .Z(n1434) );
  XNOR U1689 ( .A(n1426), .B(n1430), .Z(n1433) );
  XNOR U1690 ( .A(n1425), .B(n1423), .Z(n1430) );
  XNOR U1691 ( .A(n1424), .B(n1422), .Z(n1423) );
  XNOR U1692 ( .A(n224), .B(n1417), .Z(n1422) );
  XNOR U1693 ( .A(n223), .B(n1415), .Z(n1417) );
  XNOR U1694 ( .A(n1416), .B(n1411), .Z(n1415) );
  XNOR U1695 ( .A(n1412), .B(n239), .Z(n1411) );
  XNOR U1696 ( .A(n234), .B(n1410), .Z(n239) );
  XNOR U1697 ( .A(n233), .B(n1405), .Z(n1410) );
  XNOR U1698 ( .A(n235), .B(n1404), .Z(n1405) );
  XNOR U1699 ( .A(n238), .B(n1401), .Z(n1404) );
  XNOR U1700 ( .A(n244), .B(n1400), .Z(n1401) );
  XNOR U1701 ( .A(n1393), .B(n1397), .Z(n1400) );
  XNOR U1702 ( .A(n1392), .B(n1390), .Z(n1397) );
  XNOR U1703 ( .A(n1391), .B(n1389), .Z(n1390) );
  XNOR U1704 ( .A(n251), .B(n1384), .Z(n1389) );
  XNOR U1705 ( .A(n250), .B(n1382), .Z(n1384) );
  XNOR U1706 ( .A(n1383), .B(n1378), .Z(n1382) );
  XNOR U1707 ( .A(n1379), .B(n266), .Z(n1378) );
  XNOR U1708 ( .A(n261), .B(n1377), .Z(n266) );
  XNOR U1709 ( .A(n260), .B(n1372), .Z(n1377) );
  XNOR U1710 ( .A(n262), .B(n1371), .Z(n1372) );
  XNOR U1711 ( .A(n265), .B(n1368), .Z(n1371) );
  XNOR U1712 ( .A(n271), .B(n1367), .Z(n1368) );
  XNOR U1713 ( .A(n1360), .B(n1364), .Z(n1367) );
  XNOR U1714 ( .A(n1359), .B(n1357), .Z(n1364) );
  XNOR U1715 ( .A(n1358), .B(n1356), .Z(n1357) );
  XNOR U1716 ( .A(n278), .B(n1351), .Z(n1356) );
  XNOR U1717 ( .A(n277), .B(n1349), .Z(n1351) );
  XNOR U1718 ( .A(n1350), .B(n1345), .Z(n1349) );
  XNOR U1719 ( .A(n1346), .B(n293), .Z(n1345) );
  XNOR U1720 ( .A(n288), .B(n1344), .Z(n293) );
  XNOR U1721 ( .A(n287), .B(n1339), .Z(n1344) );
  XNOR U1722 ( .A(n289), .B(n1338), .Z(n1339) );
  XNOR U1723 ( .A(n292), .B(n1335), .Z(n1338) );
  XNOR U1724 ( .A(n298), .B(n1334), .Z(n1335) );
  XNOR U1725 ( .A(n1327), .B(n1331), .Z(n1334) );
  XNOR U1726 ( .A(n1326), .B(n1324), .Z(n1331) );
  XNOR U1727 ( .A(n1325), .B(n1323), .Z(n1324) );
  XNOR U1728 ( .A(n305), .B(n1318), .Z(n1323) );
  XNOR U1729 ( .A(n304), .B(n1316), .Z(n1318) );
  XNOR U1730 ( .A(n1317), .B(n1312), .Z(n1316) );
  XNOR U1731 ( .A(n1313), .B(n320), .Z(n1312) );
  XNOR U1732 ( .A(n315), .B(n1311), .Z(n320) );
  XNOR U1733 ( .A(n314), .B(n1306), .Z(n1311) );
  XNOR U1734 ( .A(n316), .B(n1305), .Z(n1306) );
  XNOR U1735 ( .A(n319), .B(n1302), .Z(n1305) );
  XNOR U1736 ( .A(n325), .B(n1301), .Z(n1302) );
  XNOR U1737 ( .A(n1294), .B(n1298), .Z(n1301) );
  XNOR U1738 ( .A(n1293), .B(n1291), .Z(n1298) );
  XNOR U1739 ( .A(n1292), .B(n1290), .Z(n1291) );
  XNOR U1740 ( .A(n332), .B(n1285), .Z(n1290) );
  XNOR U1741 ( .A(n331), .B(n1283), .Z(n1285) );
  XNOR U1742 ( .A(n1284), .B(n1279), .Z(n1283) );
  XNOR U1743 ( .A(n1280), .B(n347), .Z(n1279) );
  XNOR U1744 ( .A(n342), .B(n1278), .Z(n347) );
  XNOR U1745 ( .A(n341), .B(n1273), .Z(n1278) );
  XNOR U1746 ( .A(n343), .B(n1272), .Z(n1273) );
  XNOR U1747 ( .A(n346), .B(n1269), .Z(n1272) );
  XNOR U1748 ( .A(n352), .B(n1268), .Z(n1269) );
  XNOR U1749 ( .A(n1261), .B(n1265), .Z(n1268) );
  XNOR U1750 ( .A(n1260), .B(n1258), .Z(n1265) );
  XNOR U1751 ( .A(n1259), .B(n1257), .Z(n1258) );
  XNOR U1752 ( .A(n359), .B(n1252), .Z(n1257) );
  XNOR U1753 ( .A(n358), .B(n1250), .Z(n1252) );
  XNOR U1754 ( .A(n1251), .B(n1246), .Z(n1250) );
  XNOR U1755 ( .A(n1247), .B(n374), .Z(n1246) );
  XNOR U1756 ( .A(n369), .B(n1245), .Z(n374) );
  XNOR U1757 ( .A(n368), .B(n1240), .Z(n1245) );
  XNOR U1758 ( .A(n370), .B(n1239), .Z(n1240) );
  XNOR U1759 ( .A(n373), .B(n1236), .Z(n1239) );
  XNOR U1760 ( .A(n379), .B(n1235), .Z(n1236) );
  XNOR U1761 ( .A(n1228), .B(n1232), .Z(n1235) );
  XNOR U1762 ( .A(n1227), .B(n1225), .Z(n1232) );
  XNOR U1763 ( .A(n1226), .B(n1224), .Z(n1225) );
  XNOR U1764 ( .A(n386), .B(n1219), .Z(n1224) );
  XNOR U1765 ( .A(n385), .B(n1217), .Z(n1219) );
  XNOR U1766 ( .A(n1218), .B(n1213), .Z(n1217) );
  XNOR U1767 ( .A(n1214), .B(n401), .Z(n1213) );
  XNOR U1768 ( .A(n396), .B(n1212), .Z(n401) );
  XNOR U1769 ( .A(n395), .B(n1207), .Z(n1212) );
  XNOR U1770 ( .A(n397), .B(n1206), .Z(n1207) );
  XNOR U1771 ( .A(n400), .B(n1203), .Z(n1206) );
  XNOR U1772 ( .A(n406), .B(n1202), .Z(n1203) );
  XNOR U1773 ( .A(n1195), .B(n1199), .Z(n1202) );
  XNOR U1774 ( .A(n1194), .B(n1192), .Z(n1199) );
  XNOR U1775 ( .A(n1193), .B(n1191), .Z(n1192) );
  XNOR U1776 ( .A(n413), .B(n1186), .Z(n1191) );
  XNOR U1777 ( .A(n412), .B(n1184), .Z(n1186) );
  XNOR U1778 ( .A(n1185), .B(n1180), .Z(n1184) );
  XNOR U1779 ( .A(n1181), .B(n428), .Z(n1180) );
  XNOR U1780 ( .A(n423), .B(n1179), .Z(n428) );
  XNOR U1781 ( .A(n422), .B(n1174), .Z(n1179) );
  XNOR U1782 ( .A(n424), .B(n1173), .Z(n1174) );
  XNOR U1783 ( .A(n427), .B(n1170), .Z(n1173) );
  XNOR U1784 ( .A(n433), .B(n1169), .Z(n1170) );
  XNOR U1785 ( .A(n1162), .B(n1166), .Z(n1169) );
  XNOR U1786 ( .A(n1161), .B(n1159), .Z(n1166) );
  XNOR U1787 ( .A(n1160), .B(n1158), .Z(n1159) );
  XNOR U1788 ( .A(n440), .B(n1153), .Z(n1158) );
  XNOR U1789 ( .A(n439), .B(n1151), .Z(n1153) );
  XNOR U1790 ( .A(n1152), .B(n1147), .Z(n1151) );
  XNOR U1791 ( .A(n1148), .B(n455), .Z(n1147) );
  XNOR U1792 ( .A(n450), .B(n1146), .Z(n455) );
  XNOR U1793 ( .A(n449), .B(n1141), .Z(n1146) );
  XNOR U1794 ( .A(n451), .B(n1140), .Z(n1141) );
  XNOR U1795 ( .A(n454), .B(n1137), .Z(n1140) );
  XNOR U1796 ( .A(n460), .B(n1136), .Z(n1137) );
  XNOR U1797 ( .A(n1129), .B(n1133), .Z(n1136) );
  XNOR U1798 ( .A(n1128), .B(n1126), .Z(n1133) );
  XNOR U1799 ( .A(n1127), .B(n1125), .Z(n1126) );
  XNOR U1800 ( .A(n467), .B(n1120), .Z(n1125) );
  XNOR U1801 ( .A(n466), .B(n1118), .Z(n1120) );
  XNOR U1802 ( .A(n1119), .B(n1114), .Z(n1118) );
  XNOR U1803 ( .A(n1115), .B(n482), .Z(n1114) );
  XNOR U1804 ( .A(n477), .B(n1113), .Z(n482) );
  XNOR U1805 ( .A(n476), .B(n1108), .Z(n1113) );
  XNOR U1806 ( .A(n478), .B(n1107), .Z(n1108) );
  XNOR U1807 ( .A(n481), .B(n1104), .Z(n1107) );
  XNOR U1808 ( .A(n487), .B(n1103), .Z(n1104) );
  XNOR U1809 ( .A(n1096), .B(n1100), .Z(n1103) );
  XNOR U1810 ( .A(n1095), .B(n1093), .Z(n1100) );
  XNOR U1811 ( .A(n1094), .B(n1092), .Z(n1093) );
  XNOR U1812 ( .A(n494), .B(n1087), .Z(n1092) );
  XNOR U1813 ( .A(n493), .B(n1085), .Z(n1087) );
  XNOR U1814 ( .A(n1086), .B(n1081), .Z(n1085) );
  XNOR U1815 ( .A(n1082), .B(n509), .Z(n1081) );
  XNOR U1816 ( .A(n504), .B(n1080), .Z(n509) );
  XNOR U1817 ( .A(n503), .B(n1075), .Z(n1080) );
  XNOR U1818 ( .A(n505), .B(n1074), .Z(n1075) );
  XNOR U1819 ( .A(n508), .B(n1071), .Z(n1074) );
  XNOR U1820 ( .A(n514), .B(n1070), .Z(n1071) );
  XNOR U1821 ( .A(n1063), .B(n1067), .Z(n1070) );
  XNOR U1822 ( .A(n1062), .B(n1060), .Z(n1067) );
  XNOR U1823 ( .A(n1061), .B(n1059), .Z(n1060) );
  XNOR U1824 ( .A(n521), .B(n1054), .Z(n1059) );
  XNOR U1825 ( .A(n520), .B(n1052), .Z(n1054) );
  XNOR U1826 ( .A(n1053), .B(n1048), .Z(n1052) );
  XNOR U1827 ( .A(n1049), .B(n536), .Z(n1048) );
  XNOR U1828 ( .A(n531), .B(n1047), .Z(n536) );
  XNOR U1829 ( .A(n530), .B(n1042), .Z(n1047) );
  XNOR U1830 ( .A(n532), .B(n1041), .Z(n1042) );
  XNOR U1831 ( .A(n535), .B(n1038), .Z(n1041) );
  XNOR U1832 ( .A(n541), .B(n1037), .Z(n1038) );
  XNOR U1833 ( .A(n1030), .B(n1034), .Z(n1037) );
  XNOR U1834 ( .A(n1029), .B(n1027), .Z(n1034) );
  XNOR U1835 ( .A(n1028), .B(n1026), .Z(n1027) );
  XNOR U1836 ( .A(n548), .B(n1021), .Z(n1026) );
  XNOR U1837 ( .A(n547), .B(n1019), .Z(n1021) );
  XNOR U1838 ( .A(n1020), .B(n1015), .Z(n1019) );
  XNOR U1839 ( .A(n1016), .B(n563), .Z(n1015) );
  XNOR U1840 ( .A(n558), .B(n1014), .Z(n563) );
  XNOR U1841 ( .A(n557), .B(n1009), .Z(n1014) );
  XNOR U1842 ( .A(n559), .B(n1008), .Z(n1009) );
  XNOR U1843 ( .A(n562), .B(n1005), .Z(n1008) );
  XNOR U1844 ( .A(n568), .B(n1004), .Z(n1005) );
  XNOR U1845 ( .A(n997), .B(n1001), .Z(n1004) );
  XNOR U1846 ( .A(n996), .B(n994), .Z(n1001) );
  XNOR U1847 ( .A(n995), .B(n993), .Z(n994) );
  XNOR U1848 ( .A(n575), .B(n988), .Z(n993) );
  XNOR U1849 ( .A(n574), .B(n986), .Z(n988) );
  XNOR U1850 ( .A(n987), .B(n982), .Z(n986) );
  XNOR U1851 ( .A(n983), .B(n590), .Z(n982) );
  XNOR U1852 ( .A(n585), .B(n981), .Z(n590) );
  XNOR U1853 ( .A(n584), .B(n976), .Z(n981) );
  XNOR U1854 ( .A(n586), .B(n975), .Z(n976) );
  XNOR U1855 ( .A(n589), .B(n972), .Z(n975) );
  XNOR U1856 ( .A(n595), .B(n971), .Z(n972) );
  XNOR U1857 ( .A(n964), .B(n968), .Z(n971) );
  XNOR U1858 ( .A(n963), .B(n961), .Z(n968) );
  XNOR U1859 ( .A(n962), .B(n960), .Z(n961) );
  XNOR U1860 ( .A(n602), .B(n955), .Z(n960) );
  XNOR U1861 ( .A(n601), .B(n953), .Z(n955) );
  XNOR U1862 ( .A(n954), .B(n949), .Z(n953) );
  XNOR U1863 ( .A(n950), .B(n617), .Z(n949) );
  XNOR U1864 ( .A(n612), .B(n948), .Z(n617) );
  XNOR U1865 ( .A(n611), .B(n943), .Z(n948) );
  XNOR U1866 ( .A(n613), .B(n942), .Z(n943) );
  XNOR U1867 ( .A(n616), .B(n939), .Z(n942) );
  XNOR U1868 ( .A(n622), .B(n938), .Z(n939) );
  XNOR U1869 ( .A(n931), .B(n935), .Z(n938) );
  XNOR U1870 ( .A(n930), .B(n928), .Z(n935) );
  XNOR U1871 ( .A(n929), .B(n927), .Z(n928) );
  XNOR U1872 ( .A(n629), .B(n922), .Z(n927) );
  XNOR U1873 ( .A(n628), .B(n920), .Z(n922) );
  XNOR U1874 ( .A(n921), .B(n916), .Z(n920) );
  XNOR U1875 ( .A(n917), .B(n644), .Z(n916) );
  XNOR U1876 ( .A(n639), .B(n915), .Z(n644) );
  XNOR U1877 ( .A(n638), .B(n910), .Z(n915) );
  XNOR U1878 ( .A(n640), .B(n909), .Z(n910) );
  XNOR U1879 ( .A(n643), .B(n906), .Z(n909) );
  XNOR U1880 ( .A(n649), .B(n905), .Z(n906) );
  XNOR U1881 ( .A(n898), .B(n902), .Z(n905) );
  XNOR U1882 ( .A(n897), .B(n895), .Z(n902) );
  XNOR U1883 ( .A(n896), .B(n894), .Z(n895) );
  XNOR U1884 ( .A(n656), .B(n889), .Z(n894) );
  XNOR U1885 ( .A(n655), .B(n887), .Z(n889) );
  XNOR U1886 ( .A(n888), .B(n883), .Z(n887) );
  XNOR U1887 ( .A(n884), .B(n671), .Z(n883) );
  XNOR U1888 ( .A(n666), .B(n882), .Z(n671) );
  XNOR U1889 ( .A(n665), .B(n877), .Z(n882) );
  XNOR U1890 ( .A(n667), .B(n876), .Z(n877) );
  XNOR U1891 ( .A(n670), .B(n873), .Z(n876) );
  XNOR U1892 ( .A(n676), .B(n872), .Z(n873) );
  XNOR U1893 ( .A(n865), .B(n869), .Z(n872) );
  XNOR U1894 ( .A(n864), .B(n862), .Z(n869) );
  XNOR U1895 ( .A(n863), .B(n861), .Z(n862) );
  XNOR U1896 ( .A(n683), .B(n856), .Z(n861) );
  XNOR U1897 ( .A(n682), .B(n854), .Z(n856) );
  XNOR U1898 ( .A(n855), .B(n850), .Z(n854) );
  XNOR U1899 ( .A(n851), .B(n698), .Z(n850) );
  XNOR U1900 ( .A(n693), .B(n849), .Z(n698) );
  XNOR U1901 ( .A(n692), .B(n844), .Z(n849) );
  XNOR U1902 ( .A(n694), .B(n843), .Z(n844) );
  XNOR U1903 ( .A(n697), .B(n840), .Z(n843) );
  XNOR U1904 ( .A(n703), .B(n839), .Z(n840) );
  XNOR U1905 ( .A(n832), .B(n836), .Z(n839) );
  XNOR U1906 ( .A(n831), .B(n829), .Z(n836) );
  XNOR U1907 ( .A(n830), .B(n828), .Z(n829) );
  XNOR U1908 ( .A(n710), .B(n823), .Z(n828) );
  XNOR U1909 ( .A(n709), .B(n821), .Z(n823) );
  XNOR U1910 ( .A(n822), .B(n817), .Z(n821) );
  XNOR U1911 ( .A(n818), .B(n725), .Z(n817) );
  XNOR U1912 ( .A(n720), .B(n816), .Z(n725) );
  XNOR U1913 ( .A(n719), .B(n811), .Z(n816) );
  XNOR U1914 ( .A(n721), .B(n810), .Z(n811) );
  XNOR U1915 ( .A(n724), .B(n807), .Z(n810) );
  XNOR U1916 ( .A(n730), .B(n806), .Z(n807) );
  XNOR U1917 ( .A(n799), .B(n803), .Z(n806) );
  XNOR U1918 ( .A(n798), .B(n796), .Z(n803) );
  XNOR U1919 ( .A(n797), .B(n795), .Z(n796) );
  XNOR U1920 ( .A(n737), .B(n790), .Z(n795) );
  XNOR U1921 ( .A(n736), .B(n788), .Z(n790) );
  XNOR U1922 ( .A(n789), .B(n784), .Z(n788) );
  XNOR U1923 ( .A(n785), .B(n752), .Z(n784) );
  XNOR U1924 ( .A(n747), .B(n783), .Z(n752) );
  XNOR U1925 ( .A(n746), .B(n778), .Z(n783) );
  XNOR U1926 ( .A(n748), .B(n777), .Z(n778) );
  XNOR U1927 ( .A(n751), .B(n774), .Z(n777) );
  XNOR U1928 ( .A(n757), .B(n773), .Z(n774) );
  XNOR U1929 ( .A(n760), .B(n770), .Z(n773) );
  XNOR U1930 ( .A(n759), .B(n767), .Z(n770) );
  XOR U1931 ( .A(n768), .B(n766), .Z(n767) );
  XNOR U1932 ( .A(n2742), .B(n2743), .Z(n766) );
  XOR U1933 ( .A(n2744), .B(n2745), .Z(n2743) );
  XOR U1934 ( .A(n2746), .B(n2747), .Z(n2745) );
  NOR U1935 ( .A(n2748), .B(n2749), .Z(n2747) );
  NOR U1936 ( .A(n2750), .B(n2751), .Z(n2746) );
  NOR U1937 ( .A(n2752), .B(n2753), .Z(n2744) );
  XOR U1938 ( .A(n2754), .B(n2755), .Z(n2742) );
  XOR U1939 ( .A(n2756), .B(n2757), .Z(n2755) );
  XOR U1940 ( .A(n2758), .B(n2759), .Z(n2757) );
  XNOR U1941 ( .A(n2760), .B(n2761), .Z(n2759) );
  XOR U1942 ( .A(n2762), .B(n2763), .Z(n2761) );
  XOR U1943 ( .A(n2764), .B(n2765), .Z(n2763) );
  XOR U1944 ( .A(n2766), .B(n2767), .Z(n2765) );
  XOR U1945 ( .A(n2768), .B(n2769), .Z(n2764) );
  XOR U1946 ( .A(n2770), .B(n2771), .Z(n2769) );
  XOR U1947 ( .A(n2772), .B(n2773), .Z(n2771) );
  XOR U1948 ( .A(n2774), .B(n2775), .Z(n2773) );
  XOR U1949 ( .A(n2776), .B(n2777), .Z(n2775) );
  XNOR U1950 ( .A(n2778), .B(n2779), .Z(n2774) );
  XNOR U1951 ( .A(n2780), .B(n2781), .Z(n2779) );
  NOR U1952 ( .A(n2782), .B(n2777), .Z(n2780) );
  XOR U1953 ( .A(n2783), .B(n2784), .Z(n2772) );
  XOR U1954 ( .A(n2785), .B(n2786), .Z(n2784) );
  XNOR U1955 ( .A(n2787), .B(n2788), .Z(n2786) );
  XOR U1956 ( .A(n2789), .B(n2790), .Z(n2788) );
  XOR U1957 ( .A(n2791), .B(n2792), .Z(n2790) );
  XOR U1958 ( .A(n2793), .B(n2794), .Z(n2792) );
  XOR U1959 ( .A(n2795), .B(n2796), .Z(n2791) );
  XOR U1960 ( .A(n2797), .B(n2798), .Z(n2796) );
  XOR U1961 ( .A(n2799), .B(n2800), .Z(n2798) );
  XOR U1962 ( .A(n2801), .B(n2802), .Z(n2800) );
  XOR U1963 ( .A(n2803), .B(n2804), .Z(n2802) );
  XNOR U1964 ( .A(n2805), .B(n2806), .Z(n2801) );
  XNOR U1965 ( .A(n2807), .B(n2808), .Z(n2806) );
  NOR U1966 ( .A(n2809), .B(n2804), .Z(n2807) );
  XOR U1967 ( .A(n2810), .B(n2811), .Z(n2799) );
  XOR U1968 ( .A(n2812), .B(n2813), .Z(n2811) );
  XNOR U1969 ( .A(n2814), .B(n2815), .Z(n2813) );
  XOR U1970 ( .A(n2816), .B(n2817), .Z(n2815) );
  XOR U1971 ( .A(n2818), .B(n2819), .Z(n2817) );
  XOR U1972 ( .A(n2820), .B(n2821), .Z(n2819) );
  XOR U1973 ( .A(n2822), .B(n2823), .Z(n2818) );
  XOR U1974 ( .A(n2824), .B(n2825), .Z(n2823) );
  XOR U1975 ( .A(n2826), .B(n2827), .Z(n2825) );
  XOR U1976 ( .A(n2828), .B(n2829), .Z(n2827) );
  XOR U1977 ( .A(n2830), .B(n2831), .Z(n2829) );
  XNOR U1978 ( .A(n2832), .B(n2833), .Z(n2828) );
  XNOR U1979 ( .A(n2834), .B(n2835), .Z(n2833) );
  NOR U1980 ( .A(n2836), .B(n2831), .Z(n2834) );
  XOR U1981 ( .A(n2837), .B(n2838), .Z(n2826) );
  XOR U1982 ( .A(n2839), .B(n2840), .Z(n2838) );
  XNOR U1983 ( .A(n2841), .B(n2842), .Z(n2840) );
  XOR U1984 ( .A(n2843), .B(n2844), .Z(n2842) );
  XOR U1985 ( .A(n2845), .B(n2846), .Z(n2844) );
  XOR U1986 ( .A(n2847), .B(n2848), .Z(n2846) );
  XOR U1987 ( .A(n2849), .B(n2850), .Z(n2845) );
  XOR U1988 ( .A(n2851), .B(n2852), .Z(n2850) );
  XOR U1989 ( .A(n2853), .B(n2854), .Z(n2852) );
  XOR U1990 ( .A(n2855), .B(n2856), .Z(n2854) );
  XOR U1991 ( .A(n2857), .B(n2858), .Z(n2856) );
  XNOR U1992 ( .A(n2859), .B(n2860), .Z(n2855) );
  XNOR U1993 ( .A(n2861), .B(n2862), .Z(n2860) );
  NOR U1994 ( .A(n2863), .B(n2858), .Z(n2861) );
  XOR U1995 ( .A(n2864), .B(n2865), .Z(n2853) );
  XOR U1996 ( .A(n2866), .B(n2867), .Z(n2865) );
  XNOR U1997 ( .A(n2868), .B(n2869), .Z(n2867) );
  XOR U1998 ( .A(n2870), .B(n2871), .Z(n2869) );
  XOR U1999 ( .A(n2872), .B(n2873), .Z(n2871) );
  XOR U2000 ( .A(n2874), .B(n2875), .Z(n2873) );
  XOR U2001 ( .A(n2876), .B(n2877), .Z(n2872) );
  XOR U2002 ( .A(n2878), .B(n2879), .Z(n2877) );
  XOR U2003 ( .A(n2880), .B(n2881), .Z(n2879) );
  XOR U2004 ( .A(n2882), .B(n2883), .Z(n2881) );
  XOR U2005 ( .A(n2884), .B(n2885), .Z(n2883) );
  XNOR U2006 ( .A(n2886), .B(n2887), .Z(n2882) );
  XNOR U2007 ( .A(n2888), .B(n2889), .Z(n2887) );
  NOR U2008 ( .A(n2890), .B(n2885), .Z(n2888) );
  XOR U2009 ( .A(n2891), .B(n2892), .Z(n2880) );
  XOR U2010 ( .A(n2893), .B(n2894), .Z(n2892) );
  XNOR U2011 ( .A(n2895), .B(n2896), .Z(n2894) );
  XOR U2012 ( .A(n2897), .B(n2898), .Z(n2896) );
  XOR U2013 ( .A(n2899), .B(n2900), .Z(n2898) );
  XOR U2014 ( .A(n2901), .B(n2902), .Z(n2900) );
  XOR U2015 ( .A(n2903), .B(n2904), .Z(n2899) );
  XOR U2016 ( .A(n2905), .B(n2906), .Z(n2904) );
  XOR U2017 ( .A(n2907), .B(n2908), .Z(n2906) );
  XOR U2018 ( .A(n2909), .B(n2910), .Z(n2908) );
  XOR U2019 ( .A(n2911), .B(n2912), .Z(n2910) );
  XNOR U2020 ( .A(n2913), .B(n2914), .Z(n2909) );
  XNOR U2021 ( .A(n2915), .B(n2916), .Z(n2914) );
  NOR U2022 ( .A(n2917), .B(n2912), .Z(n2915) );
  XOR U2023 ( .A(n2918), .B(n2919), .Z(n2907) );
  XOR U2024 ( .A(n2920), .B(n2921), .Z(n2919) );
  XNOR U2025 ( .A(n2922), .B(n2923), .Z(n2921) );
  XOR U2026 ( .A(n2924), .B(n2925), .Z(n2923) );
  XOR U2027 ( .A(n2926), .B(n2927), .Z(n2925) );
  XOR U2028 ( .A(n2928), .B(n2929), .Z(n2927) );
  XOR U2029 ( .A(n2930), .B(n2931), .Z(n2926) );
  XOR U2030 ( .A(n2932), .B(n2933), .Z(n2931) );
  XOR U2031 ( .A(n2934), .B(n2935), .Z(n2933) );
  XOR U2032 ( .A(n2936), .B(n2937), .Z(n2935) );
  XOR U2033 ( .A(n2938), .B(n2939), .Z(n2937) );
  XNOR U2034 ( .A(n2940), .B(n2941), .Z(n2936) );
  XNOR U2035 ( .A(n2942), .B(n2943), .Z(n2941) );
  NOR U2036 ( .A(n2944), .B(n2939), .Z(n2942) );
  XOR U2037 ( .A(n2945), .B(n2946), .Z(n2934) );
  XOR U2038 ( .A(n2947), .B(n2948), .Z(n2946) );
  XNOR U2039 ( .A(n2949), .B(n2950), .Z(n2948) );
  XOR U2040 ( .A(n2951), .B(n2952), .Z(n2950) );
  XOR U2041 ( .A(n2953), .B(n2954), .Z(n2952) );
  XOR U2042 ( .A(n2955), .B(n2956), .Z(n2954) );
  XOR U2043 ( .A(n2957), .B(n2958), .Z(n2953) );
  XOR U2044 ( .A(n2959), .B(n2960), .Z(n2958) );
  XOR U2045 ( .A(n2961), .B(n2962), .Z(n2960) );
  XOR U2046 ( .A(n2963), .B(n2964), .Z(n2962) );
  XOR U2047 ( .A(n2965), .B(n2966), .Z(n2964) );
  XNOR U2048 ( .A(n2967), .B(n2968), .Z(n2963) );
  XNOR U2049 ( .A(n2969), .B(n2970), .Z(n2968) );
  NOR U2050 ( .A(n2971), .B(n2966), .Z(n2969) );
  XOR U2051 ( .A(n2972), .B(n2973), .Z(n2961) );
  XOR U2052 ( .A(n2974), .B(n2975), .Z(n2973) );
  XNOR U2053 ( .A(n2976), .B(n2977), .Z(n2975) );
  XOR U2054 ( .A(n2978), .B(n2979), .Z(n2977) );
  XOR U2055 ( .A(n2980), .B(n2981), .Z(n2979) );
  XOR U2056 ( .A(n2982), .B(n2983), .Z(n2981) );
  XOR U2057 ( .A(n2984), .B(n2985), .Z(n2980) );
  XOR U2058 ( .A(n2986), .B(n2987), .Z(n2985) );
  XOR U2059 ( .A(n2988), .B(n2989), .Z(n2987) );
  XOR U2060 ( .A(n2990), .B(n2991), .Z(n2989) );
  XOR U2061 ( .A(n2992), .B(n2993), .Z(n2991) );
  XNOR U2062 ( .A(n2994), .B(n2995), .Z(n2990) );
  XNOR U2063 ( .A(n2996), .B(n2997), .Z(n2995) );
  NOR U2064 ( .A(n2998), .B(n2993), .Z(n2996) );
  XOR U2065 ( .A(n2999), .B(n3000), .Z(n2988) );
  XOR U2066 ( .A(n3001), .B(n3002), .Z(n3000) );
  XNOR U2067 ( .A(n3003), .B(n3004), .Z(n3002) );
  XOR U2068 ( .A(n3005), .B(n3006), .Z(n3004) );
  XOR U2069 ( .A(n3007), .B(n3008), .Z(n3006) );
  XOR U2070 ( .A(n3009), .B(n3010), .Z(n3008) );
  XOR U2071 ( .A(n3011), .B(n3012), .Z(n3007) );
  XOR U2072 ( .A(n3013), .B(n3014), .Z(n3012) );
  XOR U2073 ( .A(n3015), .B(n3016), .Z(n3014) );
  XOR U2074 ( .A(n3017), .B(n3018), .Z(n3016) );
  XOR U2075 ( .A(n3019), .B(n3020), .Z(n3018) );
  XNOR U2076 ( .A(n3021), .B(n3022), .Z(n3017) );
  XNOR U2077 ( .A(n3023), .B(n3024), .Z(n3022) );
  NOR U2078 ( .A(n3025), .B(n3020), .Z(n3023) );
  XOR U2079 ( .A(n3026), .B(n3027), .Z(n3015) );
  XOR U2080 ( .A(n3028), .B(n3029), .Z(n3027) );
  XOR U2081 ( .A(n3030), .B(n3031), .Z(n3029) );
  XOR U2082 ( .A(n3032), .B(n3033), .Z(n3028) );
  XOR U2083 ( .A(n3034), .B(n3035), .Z(n3026) );
  XOR U2084 ( .A(n3036), .B(n3037), .Z(n3035) );
  AND U2085 ( .A(n3038), .B(n3039), .Z(n3037) );
  XOR U2086 ( .A(n3040), .B(n3031), .Z(n3038) );
  XOR U2087 ( .A(n3041), .B(n3042), .Z(n3031) );
  NOR U2088 ( .A(n3040), .B(n3041), .Z(n3042) );
  NOR U2089 ( .A(n3043), .B(n3032), .Z(n3036) );
  XOR U2090 ( .A(n3044), .B(n3045), .Z(n3034) );
  NOR U2091 ( .A(n3046), .B(n3033), .Z(n3045) );
  NOR U2092 ( .A(n3047), .B(n3030), .Z(n3044) );
  XOR U2093 ( .A(n3048), .B(n3049), .Z(n3013) );
  NOR U2094 ( .A(n3050), .B(n3024), .Z(n3049) );
  NOR U2095 ( .A(n3051), .B(n3021), .Z(n3048) );
  XOR U2096 ( .A(n3052), .B(n3053), .Z(n3011) );
  XOR U2097 ( .A(n3054), .B(n3055), .Z(n3053) );
  NOR U2098 ( .A(n3056), .B(n3019), .Z(n3055) );
  NOR U2099 ( .A(n3057), .B(n3058), .Z(n3054) );
  XOR U2100 ( .A(n3059), .B(n3060), .Z(n3052) );
  NOR U2101 ( .A(n3061), .B(n3062), .Z(n3060) );
  NOR U2102 ( .A(n3063), .B(n3009), .Z(n3059) );
  XOR U2103 ( .A(n3064), .B(n3065), .Z(n3005) );
  XOR U2104 ( .A(n3058), .B(n3062), .Z(n3065) );
  XOR U2105 ( .A(n3066), .B(n3067), .Z(n3064) );
  NOR U2106 ( .A(n3068), .B(n3010), .Z(n3067) );
  NOR U2107 ( .A(n3069), .B(n3070), .Z(n3066) );
  XOR U2108 ( .A(n3071), .B(n3072), .Z(n3001) );
  XOR U2109 ( .A(n3073), .B(n3074), .Z(n2999) );
  XNOR U2110 ( .A(n3075), .B(n3070), .Z(n3074) );
  NOR U2111 ( .A(n3076), .B(n3071), .Z(n3075) );
  XOR U2112 ( .A(n3077), .B(n3078), .Z(n3073) );
  NOR U2113 ( .A(n3079), .B(n3072), .Z(n3078) );
  NOR U2114 ( .A(n3080), .B(n3003), .Z(n3077) );
  XOR U2115 ( .A(n3081), .B(n3082), .Z(n2986) );
  NOR U2116 ( .A(n3083), .B(n2997), .Z(n3082) );
  NOR U2117 ( .A(n3084), .B(n2994), .Z(n3081) );
  XOR U2118 ( .A(n3085), .B(n3086), .Z(n2984) );
  XOR U2119 ( .A(n3087), .B(n3088), .Z(n3086) );
  NOR U2120 ( .A(n3089), .B(n2992), .Z(n3088) );
  NOR U2121 ( .A(n3090), .B(n3091), .Z(n3087) );
  XOR U2122 ( .A(n3092), .B(n3093), .Z(n3085) );
  NOR U2123 ( .A(n3094), .B(n3095), .Z(n3093) );
  NOR U2124 ( .A(n3096), .B(n2982), .Z(n3092) );
  XOR U2125 ( .A(n3097), .B(n3098), .Z(n2978) );
  XOR U2126 ( .A(n3091), .B(n3095), .Z(n3098) );
  XOR U2127 ( .A(n3099), .B(n3100), .Z(n3097) );
  NOR U2128 ( .A(n3101), .B(n2983), .Z(n3100) );
  NOR U2129 ( .A(n3102), .B(n3103), .Z(n3099) );
  XOR U2130 ( .A(n3104), .B(n3105), .Z(n2974) );
  XOR U2131 ( .A(n3106), .B(n3107), .Z(n2972) );
  XNOR U2132 ( .A(n3108), .B(n3103), .Z(n3107) );
  NOR U2133 ( .A(n3109), .B(n3104), .Z(n3108) );
  XOR U2134 ( .A(n3110), .B(n3111), .Z(n3106) );
  NOR U2135 ( .A(n3112), .B(n3105), .Z(n3111) );
  NOR U2136 ( .A(n3113), .B(n2976), .Z(n3110) );
  XOR U2137 ( .A(n3114), .B(n3115), .Z(n2959) );
  NOR U2138 ( .A(n3116), .B(n2970), .Z(n3115) );
  NOR U2139 ( .A(n3117), .B(n2967), .Z(n3114) );
  XOR U2140 ( .A(n3118), .B(n3119), .Z(n2957) );
  XOR U2141 ( .A(n3120), .B(n3121), .Z(n3119) );
  NOR U2142 ( .A(n3122), .B(n2965), .Z(n3121) );
  NOR U2143 ( .A(n3123), .B(n3124), .Z(n3120) );
  XOR U2144 ( .A(n3125), .B(n3126), .Z(n3118) );
  NOR U2145 ( .A(n3127), .B(n3128), .Z(n3126) );
  NOR U2146 ( .A(n3129), .B(n2955), .Z(n3125) );
  XOR U2147 ( .A(n3130), .B(n3131), .Z(n2951) );
  XOR U2148 ( .A(n3124), .B(n3128), .Z(n3131) );
  XOR U2149 ( .A(n3132), .B(n3133), .Z(n3130) );
  NOR U2150 ( .A(n3134), .B(n2956), .Z(n3133) );
  NOR U2151 ( .A(n3135), .B(n3136), .Z(n3132) );
  XOR U2152 ( .A(n3137), .B(n3138), .Z(n2947) );
  XOR U2153 ( .A(n3139), .B(n3140), .Z(n2945) );
  XNOR U2154 ( .A(n3141), .B(n3136), .Z(n3140) );
  NOR U2155 ( .A(n3142), .B(n3137), .Z(n3141) );
  XOR U2156 ( .A(n3143), .B(n3144), .Z(n3139) );
  NOR U2157 ( .A(n3145), .B(n3138), .Z(n3144) );
  NOR U2158 ( .A(n3146), .B(n2949), .Z(n3143) );
  XOR U2159 ( .A(n3147), .B(n3148), .Z(n2932) );
  NOR U2160 ( .A(n3149), .B(n2943), .Z(n3148) );
  NOR U2161 ( .A(n3150), .B(n2940), .Z(n3147) );
  XOR U2162 ( .A(n3151), .B(n3152), .Z(n2930) );
  XOR U2163 ( .A(n3153), .B(n3154), .Z(n3152) );
  NOR U2164 ( .A(n3155), .B(n2938), .Z(n3154) );
  NOR U2165 ( .A(n3156), .B(n3157), .Z(n3153) );
  XOR U2166 ( .A(n3158), .B(n3159), .Z(n3151) );
  NOR U2167 ( .A(n3160), .B(n3161), .Z(n3159) );
  NOR U2168 ( .A(n3162), .B(n2928), .Z(n3158) );
  XOR U2169 ( .A(n3163), .B(n3164), .Z(n2924) );
  XOR U2170 ( .A(n3157), .B(n3161), .Z(n3164) );
  XOR U2171 ( .A(n3165), .B(n3166), .Z(n3163) );
  NOR U2172 ( .A(n3167), .B(n2929), .Z(n3166) );
  NOR U2173 ( .A(n3168), .B(n3169), .Z(n3165) );
  XOR U2174 ( .A(n3170), .B(n3171), .Z(n2920) );
  XOR U2175 ( .A(n3172), .B(n3173), .Z(n2918) );
  XNOR U2176 ( .A(n3174), .B(n3169), .Z(n3173) );
  NOR U2177 ( .A(n3175), .B(n3170), .Z(n3174) );
  XOR U2178 ( .A(n3176), .B(n3177), .Z(n3172) );
  NOR U2179 ( .A(n3178), .B(n3171), .Z(n3177) );
  NOR U2180 ( .A(n3179), .B(n2922), .Z(n3176) );
  XOR U2181 ( .A(n3180), .B(n3181), .Z(n2905) );
  NOR U2182 ( .A(n3182), .B(n2916), .Z(n3181) );
  NOR U2183 ( .A(n3183), .B(n2913), .Z(n3180) );
  XOR U2184 ( .A(n3184), .B(n3185), .Z(n2903) );
  XOR U2185 ( .A(n3186), .B(n3187), .Z(n3185) );
  NOR U2186 ( .A(n3188), .B(n2911), .Z(n3187) );
  NOR U2187 ( .A(n3189), .B(n3190), .Z(n3186) );
  XOR U2188 ( .A(n3191), .B(n3192), .Z(n3184) );
  NOR U2189 ( .A(n3193), .B(n3194), .Z(n3192) );
  NOR U2190 ( .A(n3195), .B(n2901), .Z(n3191) );
  XOR U2191 ( .A(n3196), .B(n3197), .Z(n2897) );
  XOR U2192 ( .A(n3190), .B(n3194), .Z(n3197) );
  XOR U2193 ( .A(n3198), .B(n3199), .Z(n3196) );
  NOR U2194 ( .A(n3200), .B(n2902), .Z(n3199) );
  NOR U2195 ( .A(n3201), .B(n3202), .Z(n3198) );
  XOR U2196 ( .A(n3203), .B(n3204), .Z(n2893) );
  XOR U2197 ( .A(n3205), .B(n3206), .Z(n2891) );
  XNOR U2198 ( .A(n3207), .B(n3202), .Z(n3206) );
  NOR U2199 ( .A(n3208), .B(n3203), .Z(n3207) );
  XOR U2200 ( .A(n3209), .B(n3210), .Z(n3205) );
  NOR U2201 ( .A(n3211), .B(n3204), .Z(n3210) );
  NOR U2202 ( .A(n3212), .B(n2895), .Z(n3209) );
  XOR U2203 ( .A(n3213), .B(n3214), .Z(n2878) );
  NOR U2204 ( .A(n3215), .B(n2889), .Z(n3214) );
  NOR U2205 ( .A(n3216), .B(n2886), .Z(n3213) );
  XOR U2206 ( .A(n3217), .B(n3218), .Z(n2876) );
  XOR U2207 ( .A(n3219), .B(n3220), .Z(n3218) );
  NOR U2208 ( .A(n3221), .B(n2884), .Z(n3220) );
  NOR U2209 ( .A(n3222), .B(n3223), .Z(n3219) );
  XOR U2210 ( .A(n3224), .B(n3225), .Z(n3217) );
  NOR U2211 ( .A(n3226), .B(n3227), .Z(n3225) );
  NOR U2212 ( .A(n3228), .B(n2874), .Z(n3224) );
  XOR U2213 ( .A(n3229), .B(n3230), .Z(n2870) );
  XOR U2214 ( .A(n3223), .B(n3227), .Z(n3230) );
  XOR U2215 ( .A(n3231), .B(n3232), .Z(n3229) );
  NOR U2216 ( .A(n3233), .B(n2875), .Z(n3232) );
  NOR U2217 ( .A(n3234), .B(n3235), .Z(n3231) );
  XOR U2218 ( .A(n3236), .B(n3237), .Z(n2866) );
  XOR U2219 ( .A(n3238), .B(n3239), .Z(n2864) );
  XNOR U2220 ( .A(n3240), .B(n3235), .Z(n3239) );
  NOR U2221 ( .A(n3241), .B(n3236), .Z(n3240) );
  XOR U2222 ( .A(n3242), .B(n3243), .Z(n3238) );
  NOR U2223 ( .A(n3244), .B(n3237), .Z(n3243) );
  NOR U2224 ( .A(n3245), .B(n2868), .Z(n3242) );
  XOR U2225 ( .A(n3246), .B(n3247), .Z(n2851) );
  NOR U2226 ( .A(n3248), .B(n2862), .Z(n3247) );
  NOR U2227 ( .A(n3249), .B(n2859), .Z(n3246) );
  XOR U2228 ( .A(n3250), .B(n3251), .Z(n2849) );
  XOR U2229 ( .A(n3252), .B(n3253), .Z(n3251) );
  NOR U2230 ( .A(n3254), .B(n2857), .Z(n3253) );
  NOR U2231 ( .A(n3255), .B(n3256), .Z(n3252) );
  XOR U2232 ( .A(n3257), .B(n3258), .Z(n3250) );
  NOR U2233 ( .A(n3259), .B(n3260), .Z(n3258) );
  NOR U2234 ( .A(n3261), .B(n2847), .Z(n3257) );
  XOR U2235 ( .A(n3262), .B(n3263), .Z(n2843) );
  XOR U2236 ( .A(n3256), .B(n3260), .Z(n3263) );
  XOR U2237 ( .A(n3264), .B(n3265), .Z(n3262) );
  NOR U2238 ( .A(n3266), .B(n2848), .Z(n3265) );
  NOR U2239 ( .A(n3267), .B(n3268), .Z(n3264) );
  XOR U2240 ( .A(n3269), .B(n3270), .Z(n2839) );
  XOR U2241 ( .A(n3271), .B(n3272), .Z(n2837) );
  XNOR U2242 ( .A(n3273), .B(n3268), .Z(n3272) );
  NOR U2243 ( .A(n3274), .B(n3269), .Z(n3273) );
  XOR U2244 ( .A(n3275), .B(n3276), .Z(n3271) );
  NOR U2245 ( .A(n3277), .B(n3270), .Z(n3276) );
  NOR U2246 ( .A(n3278), .B(n2841), .Z(n3275) );
  XOR U2247 ( .A(n3279), .B(n3280), .Z(n2824) );
  NOR U2248 ( .A(n3281), .B(n2835), .Z(n3280) );
  NOR U2249 ( .A(n3282), .B(n2832), .Z(n3279) );
  XOR U2250 ( .A(n3283), .B(n3284), .Z(n2822) );
  XOR U2251 ( .A(n3285), .B(n3286), .Z(n3284) );
  NOR U2252 ( .A(n3287), .B(n2830), .Z(n3286) );
  NOR U2253 ( .A(n3288), .B(n3289), .Z(n3285) );
  XOR U2254 ( .A(n3290), .B(n3291), .Z(n3283) );
  NOR U2255 ( .A(n3292), .B(n3293), .Z(n3291) );
  NOR U2256 ( .A(n3294), .B(n2820), .Z(n3290) );
  XOR U2257 ( .A(n3295), .B(n3296), .Z(n2816) );
  XOR U2258 ( .A(n3289), .B(n3293), .Z(n3296) );
  XOR U2259 ( .A(n3297), .B(n3298), .Z(n3295) );
  NOR U2260 ( .A(n3299), .B(n2821), .Z(n3298) );
  NOR U2261 ( .A(n3300), .B(n3301), .Z(n3297) );
  XOR U2262 ( .A(n3302), .B(n3303), .Z(n2812) );
  XOR U2263 ( .A(n3304), .B(n3305), .Z(n2810) );
  XNOR U2264 ( .A(n3306), .B(n3301), .Z(n3305) );
  NOR U2265 ( .A(n3307), .B(n3302), .Z(n3306) );
  XOR U2266 ( .A(n3308), .B(n3309), .Z(n3304) );
  NOR U2267 ( .A(n3310), .B(n3303), .Z(n3309) );
  NOR U2268 ( .A(n3311), .B(n2814), .Z(n3308) );
  XOR U2269 ( .A(n3312), .B(n3313), .Z(n2797) );
  NOR U2270 ( .A(n3314), .B(n2808), .Z(n3313) );
  NOR U2271 ( .A(n3315), .B(n2805), .Z(n3312) );
  XOR U2272 ( .A(n3316), .B(n3317), .Z(n2795) );
  XOR U2273 ( .A(n3318), .B(n3319), .Z(n3317) );
  NOR U2274 ( .A(n3320), .B(n2803), .Z(n3319) );
  NOR U2275 ( .A(n3321), .B(n3322), .Z(n3318) );
  XOR U2276 ( .A(n3323), .B(n3324), .Z(n3316) );
  NOR U2277 ( .A(n3325), .B(n3326), .Z(n3324) );
  NOR U2278 ( .A(n3327), .B(n2793), .Z(n3323) );
  XOR U2279 ( .A(n3328), .B(n3329), .Z(n2789) );
  XOR U2280 ( .A(n3322), .B(n3326), .Z(n3329) );
  XOR U2281 ( .A(n3330), .B(n3331), .Z(n3328) );
  NOR U2282 ( .A(n3332), .B(n2794), .Z(n3331) );
  NOR U2283 ( .A(n3333), .B(n3334), .Z(n3330) );
  XOR U2284 ( .A(n3335), .B(n3336), .Z(n2785) );
  XOR U2285 ( .A(n3337), .B(n3338), .Z(n2783) );
  XNOR U2286 ( .A(n3339), .B(n3334), .Z(n3338) );
  NOR U2287 ( .A(n3340), .B(n3335), .Z(n3339) );
  XOR U2288 ( .A(n3341), .B(n3342), .Z(n3337) );
  NOR U2289 ( .A(n3343), .B(n3336), .Z(n3342) );
  NOR U2290 ( .A(n3344), .B(n2787), .Z(n3341) );
  XOR U2291 ( .A(n3345), .B(n3346), .Z(n2770) );
  NOR U2292 ( .A(n3347), .B(n2781), .Z(n3346) );
  NOR U2293 ( .A(n3348), .B(n2778), .Z(n3345) );
  XOR U2294 ( .A(n3349), .B(n3350), .Z(n2768) );
  XOR U2295 ( .A(n3351), .B(n3352), .Z(n3350) );
  NOR U2296 ( .A(n3353), .B(n2776), .Z(n3352) );
  NOR U2297 ( .A(n3354), .B(n3355), .Z(n3351) );
  XOR U2298 ( .A(n3356), .B(n3357), .Z(n3349) );
  NOR U2299 ( .A(n3358), .B(n3359), .Z(n3357) );
  NOR U2300 ( .A(n3360), .B(n2766), .Z(n3356) );
  XOR U2301 ( .A(n3361), .B(n3362), .Z(n2762) );
  XOR U2302 ( .A(n3355), .B(n3359), .Z(n3362) );
  XOR U2303 ( .A(n3363), .B(n3364), .Z(n3361) );
  NOR U2304 ( .A(n3365), .B(n2767), .Z(n3364) );
  NOR U2305 ( .A(n3366), .B(n3367), .Z(n3363) );
  XOR U2306 ( .A(n3368), .B(n3369), .Z(n2758) );
  XOR U2307 ( .A(n3370), .B(n3371), .Z(n2756) );
  XNOR U2308 ( .A(n3372), .B(n3367), .Z(n3371) );
  NOR U2309 ( .A(n3373), .B(n3368), .Z(n3372) );
  XOR U2310 ( .A(n3374), .B(n3375), .Z(n3370) );
  NOR U2311 ( .A(n3376), .B(n3369), .Z(n3375) );
  NOR U2312 ( .A(n3377), .B(n2760), .Z(n3374) );
  XOR U2313 ( .A(n3378), .B(n3379), .Z(n2754) );
  XNOR U2314 ( .A(n2749), .B(n3380), .Z(n3379) );
  XNOR U2315 ( .A(n3381), .B(n2753), .Z(n3380) );
  NOR U2316 ( .A(n3382), .B(n3383), .Z(n3381) );
  XNOR U2317 ( .A(n3383), .B(n2751), .Z(n3378) );
  XOR U2318 ( .A(n3384), .B(n3385), .Z(n768) );
  NOR U2319 ( .A(n3386), .B(n3384), .Z(n3385) );
  XOR U2320 ( .A(n3387), .B(n3388), .Z(n759) );
  NOR U2321 ( .A(n3389), .B(n3387), .Z(n3388) );
  XOR U2322 ( .A(n3390), .B(n3391), .Z(n760) );
  NOR U2323 ( .A(n3392), .B(n3390), .Z(n3391) );
  XOR U2324 ( .A(n3393), .B(n3394), .Z(n757) );
  NOR U2325 ( .A(n3395), .B(n3393), .Z(n3394) );
  XOR U2326 ( .A(n3396), .B(n3397), .Z(n751) );
  NOR U2327 ( .A(n3398), .B(n3396), .Z(n3397) );
  XOR U2328 ( .A(n3399), .B(n3400), .Z(n748) );
  NOR U2329 ( .A(n3401), .B(n3399), .Z(n3400) );
  XOR U2330 ( .A(n3402), .B(n3403), .Z(n746) );
  NOR U2331 ( .A(n3404), .B(n3402), .Z(n3403) );
  XOR U2332 ( .A(n3405), .B(n3406), .Z(n747) );
  NOR U2333 ( .A(n3407), .B(n3405), .Z(n3406) );
  XOR U2334 ( .A(n3408), .B(n3409), .Z(n785) );
  NOR U2335 ( .A(n3410), .B(n3408), .Z(n3409) );
  XOR U2336 ( .A(n3411), .B(n3412), .Z(n789) );
  NOR U2337 ( .A(n3413), .B(n3411), .Z(n3412) );
  XOR U2338 ( .A(n3414), .B(n3415), .Z(n736) );
  NOR U2339 ( .A(n3416), .B(n3414), .Z(n3415) );
  XOR U2340 ( .A(n3417), .B(n3418), .Z(n737) );
  NOR U2341 ( .A(n3419), .B(n3417), .Z(n3418) );
  XOR U2342 ( .A(n3420), .B(n3421), .Z(n797) );
  NOR U2343 ( .A(n3422), .B(n3420), .Z(n3421) );
  XOR U2344 ( .A(n3423), .B(n3424), .Z(n798) );
  NOR U2345 ( .A(n3425), .B(n3423), .Z(n3424) );
  XOR U2346 ( .A(n3426), .B(n3427), .Z(n799) );
  NOR U2347 ( .A(n3428), .B(n3426), .Z(n3427) );
  XOR U2348 ( .A(n3429), .B(n3430), .Z(n730) );
  NOR U2349 ( .A(n3431), .B(n3429), .Z(n3430) );
  XOR U2350 ( .A(n3432), .B(n3433), .Z(n724) );
  NOR U2351 ( .A(n3434), .B(n3432), .Z(n3433) );
  XOR U2352 ( .A(n3435), .B(n3436), .Z(n721) );
  NOR U2353 ( .A(n3437), .B(n3435), .Z(n3436) );
  XOR U2354 ( .A(n3438), .B(n3439), .Z(n719) );
  NOR U2355 ( .A(n3440), .B(n3438), .Z(n3439) );
  XOR U2356 ( .A(n3441), .B(n3442), .Z(n720) );
  NOR U2357 ( .A(n3443), .B(n3441), .Z(n3442) );
  XOR U2358 ( .A(n3444), .B(n3445), .Z(n818) );
  NOR U2359 ( .A(n3446), .B(n3444), .Z(n3445) );
  XOR U2360 ( .A(n3447), .B(n3448), .Z(n822) );
  NOR U2361 ( .A(n3449), .B(n3447), .Z(n3448) );
  XOR U2362 ( .A(n3450), .B(n3451), .Z(n709) );
  NOR U2363 ( .A(n3452), .B(n3450), .Z(n3451) );
  XOR U2364 ( .A(n3453), .B(n3454), .Z(n710) );
  NOR U2365 ( .A(n3455), .B(n3453), .Z(n3454) );
  XOR U2366 ( .A(n3456), .B(n3457), .Z(n830) );
  NOR U2367 ( .A(n3458), .B(n3456), .Z(n3457) );
  XOR U2368 ( .A(n3459), .B(n3460), .Z(n831) );
  NOR U2369 ( .A(n3461), .B(n3459), .Z(n3460) );
  XOR U2370 ( .A(n3462), .B(n3463), .Z(n832) );
  NOR U2371 ( .A(n3464), .B(n3462), .Z(n3463) );
  XOR U2372 ( .A(n3465), .B(n3466), .Z(n703) );
  NOR U2373 ( .A(n3467), .B(n3465), .Z(n3466) );
  XOR U2374 ( .A(n3468), .B(n3469), .Z(n697) );
  NOR U2375 ( .A(n3470), .B(n3468), .Z(n3469) );
  XOR U2376 ( .A(n3471), .B(n3472), .Z(n694) );
  NOR U2377 ( .A(n3473), .B(n3471), .Z(n3472) );
  XOR U2378 ( .A(n3474), .B(n3475), .Z(n692) );
  NOR U2379 ( .A(n3476), .B(n3474), .Z(n3475) );
  XOR U2380 ( .A(n3477), .B(n3478), .Z(n693) );
  NOR U2381 ( .A(n3479), .B(n3477), .Z(n3478) );
  XOR U2382 ( .A(n3480), .B(n3481), .Z(n851) );
  NOR U2383 ( .A(n3482), .B(n3480), .Z(n3481) );
  XOR U2384 ( .A(n3483), .B(n3484), .Z(n855) );
  NOR U2385 ( .A(n3485), .B(n3483), .Z(n3484) );
  XOR U2386 ( .A(n3486), .B(n3487), .Z(n682) );
  NOR U2387 ( .A(n3488), .B(n3486), .Z(n3487) );
  XOR U2388 ( .A(n3489), .B(n3490), .Z(n683) );
  NOR U2389 ( .A(n3491), .B(n3489), .Z(n3490) );
  XOR U2390 ( .A(n3492), .B(n3493), .Z(n863) );
  NOR U2391 ( .A(n3494), .B(n3492), .Z(n3493) );
  XOR U2392 ( .A(n3495), .B(n3496), .Z(n864) );
  NOR U2393 ( .A(n3497), .B(n3495), .Z(n3496) );
  XOR U2394 ( .A(n3498), .B(n3499), .Z(n865) );
  NOR U2395 ( .A(n3500), .B(n3498), .Z(n3499) );
  XOR U2396 ( .A(n3501), .B(n3502), .Z(n676) );
  NOR U2397 ( .A(n3503), .B(n3501), .Z(n3502) );
  XOR U2398 ( .A(n3504), .B(n3505), .Z(n670) );
  NOR U2399 ( .A(n3506), .B(n3504), .Z(n3505) );
  XOR U2400 ( .A(n3507), .B(n3508), .Z(n667) );
  NOR U2401 ( .A(n3509), .B(n3507), .Z(n3508) );
  XOR U2402 ( .A(n3510), .B(n3511), .Z(n665) );
  NOR U2403 ( .A(n3512), .B(n3510), .Z(n3511) );
  XOR U2404 ( .A(n3513), .B(n3514), .Z(n666) );
  NOR U2405 ( .A(n3515), .B(n3513), .Z(n3514) );
  XOR U2406 ( .A(n3516), .B(n3517), .Z(n884) );
  NOR U2407 ( .A(n3518), .B(n3516), .Z(n3517) );
  XOR U2408 ( .A(n3519), .B(n3520), .Z(n888) );
  NOR U2409 ( .A(n3521), .B(n3519), .Z(n3520) );
  XOR U2410 ( .A(n3522), .B(n3523), .Z(n655) );
  NOR U2411 ( .A(n3524), .B(n3522), .Z(n3523) );
  XOR U2412 ( .A(n3525), .B(n3526), .Z(n656) );
  NOR U2413 ( .A(n3527), .B(n3525), .Z(n3526) );
  XOR U2414 ( .A(n3528), .B(n3529), .Z(n896) );
  NOR U2415 ( .A(n3530), .B(n3528), .Z(n3529) );
  XOR U2416 ( .A(n3531), .B(n3532), .Z(n897) );
  NOR U2417 ( .A(n3533), .B(n3531), .Z(n3532) );
  XOR U2418 ( .A(n3534), .B(n3535), .Z(n898) );
  NOR U2419 ( .A(n3536), .B(n3534), .Z(n3535) );
  XOR U2420 ( .A(n3537), .B(n3538), .Z(n649) );
  NOR U2421 ( .A(n3539), .B(n3537), .Z(n3538) );
  XOR U2422 ( .A(n3540), .B(n3541), .Z(n643) );
  NOR U2423 ( .A(n3542), .B(n3540), .Z(n3541) );
  XOR U2424 ( .A(n3543), .B(n3544), .Z(n640) );
  NOR U2425 ( .A(n3545), .B(n3543), .Z(n3544) );
  XOR U2426 ( .A(n3546), .B(n3547), .Z(n638) );
  NOR U2427 ( .A(n3548), .B(n3546), .Z(n3547) );
  XOR U2428 ( .A(n3549), .B(n3550), .Z(n639) );
  NOR U2429 ( .A(n3551), .B(n3549), .Z(n3550) );
  XOR U2430 ( .A(n3552), .B(n3553), .Z(n917) );
  NOR U2431 ( .A(n3554), .B(n3552), .Z(n3553) );
  XOR U2432 ( .A(n3555), .B(n3556), .Z(n921) );
  NOR U2433 ( .A(n3557), .B(n3555), .Z(n3556) );
  XOR U2434 ( .A(n3558), .B(n3559), .Z(n628) );
  NOR U2435 ( .A(n3560), .B(n3558), .Z(n3559) );
  XOR U2436 ( .A(n3561), .B(n3562), .Z(n629) );
  NOR U2437 ( .A(n3563), .B(n3561), .Z(n3562) );
  XOR U2438 ( .A(n3564), .B(n3565), .Z(n929) );
  NOR U2439 ( .A(n3566), .B(n3564), .Z(n3565) );
  XOR U2440 ( .A(n3567), .B(n3568), .Z(n930) );
  NOR U2441 ( .A(n3569), .B(n3567), .Z(n3568) );
  XOR U2442 ( .A(n3570), .B(n3571), .Z(n931) );
  NOR U2443 ( .A(n3572), .B(n3570), .Z(n3571) );
  XOR U2444 ( .A(n3573), .B(n3574), .Z(n622) );
  NOR U2445 ( .A(n3575), .B(n3573), .Z(n3574) );
  XOR U2446 ( .A(n3576), .B(n3577), .Z(n616) );
  NOR U2447 ( .A(n3578), .B(n3576), .Z(n3577) );
  XOR U2448 ( .A(n3579), .B(n3580), .Z(n613) );
  NOR U2449 ( .A(n3581), .B(n3579), .Z(n3580) );
  XOR U2450 ( .A(n3582), .B(n3583), .Z(n611) );
  NOR U2451 ( .A(n3584), .B(n3582), .Z(n3583) );
  XOR U2452 ( .A(n3585), .B(n3586), .Z(n612) );
  NOR U2453 ( .A(n3587), .B(n3585), .Z(n3586) );
  XOR U2454 ( .A(n3588), .B(n3589), .Z(n950) );
  NOR U2455 ( .A(n3590), .B(n3588), .Z(n3589) );
  XOR U2456 ( .A(n3591), .B(n3592), .Z(n954) );
  NOR U2457 ( .A(n3593), .B(n3591), .Z(n3592) );
  XOR U2458 ( .A(n3594), .B(n3595), .Z(n601) );
  NOR U2459 ( .A(n3596), .B(n3594), .Z(n3595) );
  XOR U2460 ( .A(n3597), .B(n3598), .Z(n602) );
  NOR U2461 ( .A(n3599), .B(n3597), .Z(n3598) );
  XOR U2462 ( .A(n3600), .B(n3601), .Z(n962) );
  NOR U2463 ( .A(n3602), .B(n3600), .Z(n3601) );
  XOR U2464 ( .A(n3603), .B(n3604), .Z(n963) );
  NOR U2465 ( .A(n3605), .B(n3603), .Z(n3604) );
  XOR U2466 ( .A(n3606), .B(n3607), .Z(n964) );
  NOR U2467 ( .A(n3608), .B(n3606), .Z(n3607) );
  XOR U2468 ( .A(n3609), .B(n3610), .Z(n595) );
  NOR U2469 ( .A(n3611), .B(n3609), .Z(n3610) );
  XOR U2470 ( .A(n3612), .B(n3613), .Z(n589) );
  NOR U2471 ( .A(n3614), .B(n3612), .Z(n3613) );
  XOR U2472 ( .A(n3615), .B(n3616), .Z(n586) );
  NOR U2473 ( .A(n3617), .B(n3615), .Z(n3616) );
  XOR U2474 ( .A(n3618), .B(n3619), .Z(n584) );
  NOR U2475 ( .A(n3620), .B(n3618), .Z(n3619) );
  XOR U2476 ( .A(n3621), .B(n3622), .Z(n585) );
  NOR U2477 ( .A(n3623), .B(n3621), .Z(n3622) );
  XOR U2478 ( .A(n3624), .B(n3625), .Z(n983) );
  NOR U2479 ( .A(n3626), .B(n3624), .Z(n3625) );
  XOR U2480 ( .A(n3627), .B(n3628), .Z(n987) );
  NOR U2481 ( .A(n3629), .B(n3627), .Z(n3628) );
  XOR U2482 ( .A(n3630), .B(n3631), .Z(n574) );
  NOR U2483 ( .A(n3632), .B(n3630), .Z(n3631) );
  XOR U2484 ( .A(n3633), .B(n3634), .Z(n575) );
  NOR U2485 ( .A(n3635), .B(n3633), .Z(n3634) );
  XOR U2486 ( .A(n3636), .B(n3637), .Z(n995) );
  NOR U2487 ( .A(n3638), .B(n3636), .Z(n3637) );
  XOR U2488 ( .A(n3639), .B(n3640), .Z(n996) );
  NOR U2489 ( .A(n3641), .B(n3639), .Z(n3640) );
  XOR U2490 ( .A(n3642), .B(n3643), .Z(n997) );
  NOR U2491 ( .A(n3644), .B(n3642), .Z(n3643) );
  XOR U2492 ( .A(n3645), .B(n3646), .Z(n568) );
  NOR U2493 ( .A(n3647), .B(n3645), .Z(n3646) );
  XOR U2494 ( .A(n3648), .B(n3649), .Z(n562) );
  NOR U2495 ( .A(n3650), .B(n3648), .Z(n3649) );
  XOR U2496 ( .A(n3651), .B(n3652), .Z(n559) );
  NOR U2497 ( .A(n3653), .B(n3651), .Z(n3652) );
  XOR U2498 ( .A(n3654), .B(n3655), .Z(n557) );
  NOR U2499 ( .A(n3656), .B(n3654), .Z(n3655) );
  XOR U2500 ( .A(n3657), .B(n3658), .Z(n558) );
  NOR U2501 ( .A(n3659), .B(n3657), .Z(n3658) );
  XOR U2502 ( .A(n3660), .B(n3661), .Z(n1016) );
  NOR U2503 ( .A(n3662), .B(n3660), .Z(n3661) );
  XOR U2504 ( .A(n3663), .B(n3664), .Z(n1020) );
  NOR U2505 ( .A(n3665), .B(n3663), .Z(n3664) );
  XOR U2506 ( .A(n3666), .B(n3667), .Z(n547) );
  NOR U2507 ( .A(n3668), .B(n3666), .Z(n3667) );
  XOR U2508 ( .A(n3669), .B(n3670), .Z(n548) );
  NOR U2509 ( .A(n3671), .B(n3669), .Z(n3670) );
  XOR U2510 ( .A(n3672), .B(n3673), .Z(n1028) );
  NOR U2511 ( .A(n3674), .B(n3672), .Z(n3673) );
  XOR U2512 ( .A(n3675), .B(n3676), .Z(n1029) );
  NOR U2513 ( .A(n3677), .B(n3675), .Z(n3676) );
  XOR U2514 ( .A(n3678), .B(n3679), .Z(n1030) );
  NOR U2515 ( .A(n3680), .B(n3678), .Z(n3679) );
  XOR U2516 ( .A(n3681), .B(n3682), .Z(n541) );
  NOR U2517 ( .A(n3683), .B(n3681), .Z(n3682) );
  XOR U2518 ( .A(n3684), .B(n3685), .Z(n535) );
  NOR U2519 ( .A(n3686), .B(n3684), .Z(n3685) );
  XOR U2520 ( .A(n3687), .B(n3688), .Z(n532) );
  NOR U2521 ( .A(n3689), .B(n3687), .Z(n3688) );
  XOR U2522 ( .A(n3690), .B(n3691), .Z(n530) );
  NOR U2523 ( .A(n3692), .B(n3690), .Z(n3691) );
  XOR U2524 ( .A(n3693), .B(n3694), .Z(n531) );
  NOR U2525 ( .A(n3695), .B(n3693), .Z(n3694) );
  XOR U2526 ( .A(n3696), .B(n3697), .Z(n1049) );
  NOR U2527 ( .A(n3698), .B(n3696), .Z(n3697) );
  XOR U2528 ( .A(n3699), .B(n3700), .Z(n1053) );
  NOR U2529 ( .A(n3701), .B(n3699), .Z(n3700) );
  XOR U2530 ( .A(n3702), .B(n3703), .Z(n520) );
  NOR U2531 ( .A(n3704), .B(n3702), .Z(n3703) );
  XOR U2532 ( .A(n3705), .B(n3706), .Z(n521) );
  NOR U2533 ( .A(n3707), .B(n3705), .Z(n3706) );
  XOR U2534 ( .A(n3708), .B(n3709), .Z(n1061) );
  NOR U2535 ( .A(n3710), .B(n3708), .Z(n3709) );
  XOR U2536 ( .A(n3711), .B(n3712), .Z(n1062) );
  NOR U2537 ( .A(n3713), .B(n3711), .Z(n3712) );
  XOR U2538 ( .A(n3714), .B(n3715), .Z(n1063) );
  NOR U2539 ( .A(n3716), .B(n3714), .Z(n3715) );
  XOR U2540 ( .A(n3717), .B(n3718), .Z(n514) );
  NOR U2541 ( .A(n3719), .B(n3717), .Z(n3718) );
  XOR U2542 ( .A(n3720), .B(n3721), .Z(n508) );
  NOR U2543 ( .A(n3722), .B(n3720), .Z(n3721) );
  XOR U2544 ( .A(n3723), .B(n3724), .Z(n505) );
  NOR U2545 ( .A(n3725), .B(n3723), .Z(n3724) );
  XOR U2546 ( .A(n3726), .B(n3727), .Z(n503) );
  NOR U2547 ( .A(n3728), .B(n3726), .Z(n3727) );
  XOR U2548 ( .A(n3729), .B(n3730), .Z(n504) );
  NOR U2549 ( .A(n3731), .B(n3729), .Z(n3730) );
  XOR U2550 ( .A(n3732), .B(n3733), .Z(n1082) );
  NOR U2551 ( .A(n3734), .B(n3732), .Z(n3733) );
  XOR U2552 ( .A(n3735), .B(n3736), .Z(n1086) );
  NOR U2553 ( .A(n3737), .B(n3735), .Z(n3736) );
  XOR U2554 ( .A(n3738), .B(n3739), .Z(n493) );
  NOR U2555 ( .A(n3740), .B(n3738), .Z(n3739) );
  XOR U2556 ( .A(n3741), .B(n3742), .Z(n494) );
  NOR U2557 ( .A(n3743), .B(n3741), .Z(n3742) );
  XOR U2558 ( .A(n3744), .B(n3745), .Z(n1094) );
  NOR U2559 ( .A(n3746), .B(n3744), .Z(n3745) );
  XOR U2560 ( .A(n3747), .B(n3748), .Z(n1095) );
  NOR U2561 ( .A(n3749), .B(n3747), .Z(n3748) );
  XOR U2562 ( .A(n3750), .B(n3751), .Z(n1096) );
  NOR U2563 ( .A(n3752), .B(n3750), .Z(n3751) );
  XOR U2564 ( .A(n3753), .B(n3754), .Z(n487) );
  NOR U2565 ( .A(n3755), .B(n3753), .Z(n3754) );
  XOR U2566 ( .A(n3756), .B(n3757), .Z(n481) );
  NOR U2567 ( .A(n3758), .B(n3756), .Z(n3757) );
  XOR U2568 ( .A(n3759), .B(n3760), .Z(n478) );
  NOR U2569 ( .A(n3761), .B(n3759), .Z(n3760) );
  XOR U2570 ( .A(n3762), .B(n3763), .Z(n476) );
  NOR U2571 ( .A(n3764), .B(n3762), .Z(n3763) );
  XOR U2572 ( .A(n3765), .B(n3766), .Z(n477) );
  NOR U2573 ( .A(n3767), .B(n3765), .Z(n3766) );
  XOR U2574 ( .A(n3768), .B(n3769), .Z(n1115) );
  NOR U2575 ( .A(n3770), .B(n3768), .Z(n3769) );
  XOR U2576 ( .A(n3771), .B(n3772), .Z(n1119) );
  NOR U2577 ( .A(n3773), .B(n3771), .Z(n3772) );
  XOR U2578 ( .A(n3774), .B(n3775), .Z(n466) );
  NOR U2579 ( .A(n3776), .B(n3774), .Z(n3775) );
  XOR U2580 ( .A(n3777), .B(n3778), .Z(n467) );
  NOR U2581 ( .A(n3779), .B(n3777), .Z(n3778) );
  XOR U2582 ( .A(n3780), .B(n3781), .Z(n1127) );
  NOR U2583 ( .A(n3782), .B(n3780), .Z(n3781) );
  XOR U2584 ( .A(n3783), .B(n3784), .Z(n1128) );
  NOR U2585 ( .A(n3785), .B(n3783), .Z(n3784) );
  XOR U2586 ( .A(n3786), .B(n3787), .Z(n1129) );
  NOR U2587 ( .A(n3788), .B(n3786), .Z(n3787) );
  XOR U2588 ( .A(n3789), .B(n3790), .Z(n460) );
  NOR U2589 ( .A(n3791), .B(n3789), .Z(n3790) );
  XOR U2590 ( .A(n3792), .B(n3793), .Z(n454) );
  NOR U2591 ( .A(n3794), .B(n3792), .Z(n3793) );
  XOR U2592 ( .A(n3795), .B(n3796), .Z(n451) );
  NOR U2593 ( .A(n3797), .B(n3795), .Z(n3796) );
  XOR U2594 ( .A(n3798), .B(n3799), .Z(n449) );
  NOR U2595 ( .A(n3800), .B(n3798), .Z(n3799) );
  XOR U2596 ( .A(n3801), .B(n3802), .Z(n450) );
  NOR U2597 ( .A(n3803), .B(n3801), .Z(n3802) );
  XOR U2598 ( .A(n3804), .B(n3805), .Z(n1148) );
  NOR U2599 ( .A(n3806), .B(n3804), .Z(n3805) );
  XOR U2600 ( .A(n3807), .B(n3808), .Z(n1152) );
  NOR U2601 ( .A(n3809), .B(n3807), .Z(n3808) );
  XOR U2602 ( .A(n3810), .B(n3811), .Z(n439) );
  NOR U2603 ( .A(n3812), .B(n3810), .Z(n3811) );
  XOR U2604 ( .A(n3813), .B(n3814), .Z(n440) );
  NOR U2605 ( .A(n3815), .B(n3813), .Z(n3814) );
  XOR U2606 ( .A(n3816), .B(n3817), .Z(n1160) );
  NOR U2607 ( .A(n3818), .B(n3816), .Z(n3817) );
  XOR U2608 ( .A(n3819), .B(n3820), .Z(n1161) );
  NOR U2609 ( .A(n3821), .B(n3819), .Z(n3820) );
  XOR U2610 ( .A(n3822), .B(n3823), .Z(n1162) );
  NOR U2611 ( .A(n3824), .B(n3822), .Z(n3823) );
  XOR U2612 ( .A(n3825), .B(n3826), .Z(n433) );
  NOR U2613 ( .A(n3827), .B(n3825), .Z(n3826) );
  XOR U2614 ( .A(n3828), .B(n3829), .Z(n427) );
  NOR U2615 ( .A(n3830), .B(n3828), .Z(n3829) );
  XOR U2616 ( .A(n3831), .B(n3832), .Z(n424) );
  NOR U2617 ( .A(n3833), .B(n3831), .Z(n3832) );
  XOR U2618 ( .A(n3834), .B(n3835), .Z(n422) );
  NOR U2619 ( .A(n3836), .B(n3834), .Z(n3835) );
  XOR U2620 ( .A(n3837), .B(n3838), .Z(n423) );
  NOR U2621 ( .A(n3839), .B(n3837), .Z(n3838) );
  XOR U2622 ( .A(n3840), .B(n3841), .Z(n1181) );
  NOR U2623 ( .A(n3842), .B(n3840), .Z(n3841) );
  XOR U2624 ( .A(n3843), .B(n3844), .Z(n1185) );
  NOR U2625 ( .A(n3845), .B(n3843), .Z(n3844) );
  XOR U2626 ( .A(n3846), .B(n3847), .Z(n412) );
  NOR U2627 ( .A(n3848), .B(n3846), .Z(n3847) );
  XOR U2628 ( .A(n3849), .B(n3850), .Z(n413) );
  NOR U2629 ( .A(n3851), .B(n3849), .Z(n3850) );
  XOR U2630 ( .A(n3852), .B(n3853), .Z(n1193) );
  NOR U2631 ( .A(n3854), .B(n3852), .Z(n3853) );
  XOR U2632 ( .A(n3855), .B(n3856), .Z(n1194) );
  NOR U2633 ( .A(n3857), .B(n3855), .Z(n3856) );
  XOR U2634 ( .A(n3858), .B(n3859), .Z(n1195) );
  NOR U2635 ( .A(n3860), .B(n3858), .Z(n3859) );
  XOR U2636 ( .A(n3861), .B(n3862), .Z(n406) );
  NOR U2637 ( .A(n3863), .B(n3861), .Z(n3862) );
  XOR U2638 ( .A(n3864), .B(n3865), .Z(n400) );
  NOR U2639 ( .A(n3866), .B(n3864), .Z(n3865) );
  XOR U2640 ( .A(n3867), .B(n3868), .Z(n397) );
  NOR U2641 ( .A(n3869), .B(n3867), .Z(n3868) );
  XOR U2642 ( .A(n3870), .B(n3871), .Z(n395) );
  NOR U2643 ( .A(n3872), .B(n3870), .Z(n3871) );
  XOR U2644 ( .A(n3873), .B(n3874), .Z(n396) );
  NOR U2645 ( .A(n3875), .B(n3873), .Z(n3874) );
  XOR U2646 ( .A(n3876), .B(n3877), .Z(n1214) );
  NOR U2647 ( .A(n3878), .B(n3876), .Z(n3877) );
  XOR U2648 ( .A(n3879), .B(n3880), .Z(n1218) );
  NOR U2649 ( .A(n3881), .B(n3879), .Z(n3880) );
  XOR U2650 ( .A(n3882), .B(n3883), .Z(n385) );
  NOR U2651 ( .A(n3884), .B(n3882), .Z(n3883) );
  XOR U2652 ( .A(n3885), .B(n3886), .Z(n386) );
  NOR U2653 ( .A(n3887), .B(n3885), .Z(n3886) );
  XOR U2654 ( .A(n3888), .B(n3889), .Z(n1226) );
  NOR U2655 ( .A(n3890), .B(n3888), .Z(n3889) );
  XOR U2656 ( .A(n3891), .B(n3892), .Z(n1227) );
  NOR U2657 ( .A(n3893), .B(n3891), .Z(n3892) );
  XOR U2658 ( .A(n3894), .B(n3895), .Z(n1228) );
  NOR U2659 ( .A(n3896), .B(n3894), .Z(n3895) );
  XOR U2660 ( .A(n3897), .B(n3898), .Z(n379) );
  NOR U2661 ( .A(n3899), .B(n3897), .Z(n3898) );
  XOR U2662 ( .A(n3900), .B(n3901), .Z(n373) );
  NOR U2663 ( .A(n3902), .B(n3900), .Z(n3901) );
  XOR U2664 ( .A(n3903), .B(n3904), .Z(n370) );
  NOR U2665 ( .A(n3905), .B(n3903), .Z(n3904) );
  XOR U2666 ( .A(n3906), .B(n3907), .Z(n368) );
  NOR U2667 ( .A(n3908), .B(n3906), .Z(n3907) );
  XOR U2668 ( .A(n3909), .B(n3910), .Z(n369) );
  NOR U2669 ( .A(n3911), .B(n3909), .Z(n3910) );
  XOR U2670 ( .A(n3912), .B(n3913), .Z(n1247) );
  NOR U2671 ( .A(n3914), .B(n3912), .Z(n3913) );
  XOR U2672 ( .A(n3915), .B(n3916), .Z(n1251) );
  NOR U2673 ( .A(n3917), .B(n3915), .Z(n3916) );
  XOR U2674 ( .A(n3918), .B(n3919), .Z(n358) );
  NOR U2675 ( .A(n3920), .B(n3918), .Z(n3919) );
  XOR U2676 ( .A(n3921), .B(n3922), .Z(n359) );
  NOR U2677 ( .A(n3923), .B(n3921), .Z(n3922) );
  XOR U2678 ( .A(n3924), .B(n3925), .Z(n1259) );
  NOR U2679 ( .A(n3926), .B(n3924), .Z(n3925) );
  XOR U2680 ( .A(n3927), .B(n3928), .Z(n1260) );
  NOR U2681 ( .A(n3929), .B(n3927), .Z(n3928) );
  XOR U2682 ( .A(n3930), .B(n3931), .Z(n1261) );
  NOR U2683 ( .A(n3932), .B(n3930), .Z(n3931) );
  XOR U2684 ( .A(n3933), .B(n3934), .Z(n352) );
  NOR U2685 ( .A(n3935), .B(n3933), .Z(n3934) );
  XOR U2686 ( .A(n3936), .B(n3937), .Z(n346) );
  NOR U2687 ( .A(n3938), .B(n3936), .Z(n3937) );
  XOR U2688 ( .A(n3939), .B(n3940), .Z(n343) );
  NOR U2689 ( .A(n3941), .B(n3939), .Z(n3940) );
  XOR U2690 ( .A(n3942), .B(n3943), .Z(n341) );
  NOR U2691 ( .A(n3944), .B(n3942), .Z(n3943) );
  XOR U2692 ( .A(n3945), .B(n3946), .Z(n342) );
  NOR U2693 ( .A(n3947), .B(n3945), .Z(n3946) );
  XOR U2694 ( .A(n3948), .B(n3949), .Z(n1280) );
  NOR U2695 ( .A(n3950), .B(n3948), .Z(n3949) );
  XOR U2696 ( .A(n3951), .B(n3952), .Z(n1284) );
  NOR U2697 ( .A(n3953), .B(n3951), .Z(n3952) );
  XOR U2698 ( .A(n3954), .B(n3955), .Z(n331) );
  NOR U2699 ( .A(n3956), .B(n3954), .Z(n3955) );
  XOR U2700 ( .A(n3957), .B(n3958), .Z(n332) );
  NOR U2701 ( .A(n3959), .B(n3957), .Z(n3958) );
  XOR U2702 ( .A(n3960), .B(n3961), .Z(n1292) );
  NOR U2703 ( .A(n3962), .B(n3960), .Z(n3961) );
  XOR U2704 ( .A(n3963), .B(n3964), .Z(n1293) );
  NOR U2705 ( .A(n3965), .B(n3963), .Z(n3964) );
  XOR U2706 ( .A(n3966), .B(n3967), .Z(n1294) );
  NOR U2707 ( .A(n3968), .B(n3966), .Z(n3967) );
  XOR U2708 ( .A(n3969), .B(n3970), .Z(n325) );
  NOR U2709 ( .A(n3971), .B(n3969), .Z(n3970) );
  XOR U2710 ( .A(n3972), .B(n3973), .Z(n319) );
  NOR U2711 ( .A(n3974), .B(n3972), .Z(n3973) );
  XOR U2712 ( .A(n3975), .B(n3976), .Z(n316) );
  NOR U2713 ( .A(n3977), .B(n3975), .Z(n3976) );
  XOR U2714 ( .A(n3978), .B(n3979), .Z(n314) );
  NOR U2715 ( .A(n3980), .B(n3978), .Z(n3979) );
  XOR U2716 ( .A(n3981), .B(n3982), .Z(n315) );
  NOR U2717 ( .A(n3983), .B(n3981), .Z(n3982) );
  XOR U2718 ( .A(n3984), .B(n3985), .Z(n1313) );
  NOR U2719 ( .A(n3986), .B(n3984), .Z(n3985) );
  XOR U2720 ( .A(n3987), .B(n3988), .Z(n1317) );
  NOR U2721 ( .A(n3989), .B(n3987), .Z(n3988) );
  XOR U2722 ( .A(n3990), .B(n3991), .Z(n304) );
  NOR U2723 ( .A(n3992), .B(n3990), .Z(n3991) );
  XOR U2724 ( .A(n3993), .B(n3994), .Z(n305) );
  NOR U2725 ( .A(n3995), .B(n3993), .Z(n3994) );
  XOR U2726 ( .A(n3996), .B(n3997), .Z(n1325) );
  NOR U2727 ( .A(n3998), .B(n3996), .Z(n3997) );
  XOR U2728 ( .A(n3999), .B(n4000), .Z(n1326) );
  NOR U2729 ( .A(n4001), .B(n3999), .Z(n4000) );
  XOR U2730 ( .A(n4002), .B(n4003), .Z(n1327) );
  NOR U2731 ( .A(n4004), .B(n4002), .Z(n4003) );
  XOR U2732 ( .A(n4005), .B(n4006), .Z(n298) );
  NOR U2733 ( .A(n4007), .B(n4005), .Z(n4006) );
  XOR U2734 ( .A(n4008), .B(n4009), .Z(n292) );
  NOR U2735 ( .A(n4010), .B(n4008), .Z(n4009) );
  XOR U2736 ( .A(n4011), .B(n4012), .Z(n289) );
  NOR U2737 ( .A(n4013), .B(n4011), .Z(n4012) );
  XOR U2738 ( .A(n4014), .B(n4015), .Z(n287) );
  NOR U2739 ( .A(n4016), .B(n4014), .Z(n4015) );
  XOR U2740 ( .A(n4017), .B(n4018), .Z(n288) );
  NOR U2741 ( .A(n4019), .B(n4017), .Z(n4018) );
  XOR U2742 ( .A(n4020), .B(n4021), .Z(n1346) );
  NOR U2743 ( .A(n4022), .B(n4020), .Z(n4021) );
  XOR U2744 ( .A(n4023), .B(n4024), .Z(n1350) );
  NOR U2745 ( .A(n4025), .B(n4023), .Z(n4024) );
  XOR U2746 ( .A(n4026), .B(n4027), .Z(n277) );
  NOR U2747 ( .A(n4028), .B(n4026), .Z(n4027) );
  XOR U2748 ( .A(n4029), .B(n4030), .Z(n278) );
  NOR U2749 ( .A(n4031), .B(n4029), .Z(n4030) );
  XOR U2750 ( .A(n4032), .B(n4033), .Z(n1358) );
  NOR U2751 ( .A(n4034), .B(n4032), .Z(n4033) );
  XOR U2752 ( .A(n4035), .B(n4036), .Z(n1359) );
  NOR U2753 ( .A(n4037), .B(n4035), .Z(n4036) );
  XOR U2754 ( .A(n4038), .B(n4039), .Z(n1360) );
  NOR U2755 ( .A(n4040), .B(n4038), .Z(n4039) );
  XOR U2756 ( .A(n4041), .B(n4042), .Z(n271) );
  NOR U2757 ( .A(n4043), .B(n4041), .Z(n4042) );
  XOR U2758 ( .A(n4044), .B(n4045), .Z(n265) );
  NOR U2759 ( .A(n4046), .B(n4044), .Z(n4045) );
  XOR U2760 ( .A(n4047), .B(n4048), .Z(n262) );
  NOR U2761 ( .A(n4049), .B(n4047), .Z(n4048) );
  XOR U2762 ( .A(n4050), .B(n4051), .Z(n260) );
  NOR U2763 ( .A(n4052), .B(n4050), .Z(n4051) );
  XOR U2764 ( .A(n4053), .B(n4054), .Z(n261) );
  NOR U2765 ( .A(n4055), .B(n4053), .Z(n4054) );
  XOR U2766 ( .A(n4056), .B(n4057), .Z(n1379) );
  NOR U2767 ( .A(n4058), .B(n4056), .Z(n4057) );
  XOR U2768 ( .A(n4059), .B(n4060), .Z(n1383) );
  NOR U2769 ( .A(n4061), .B(n4059), .Z(n4060) );
  XOR U2770 ( .A(n4062), .B(n4063), .Z(n250) );
  NOR U2771 ( .A(n4064), .B(n4062), .Z(n4063) );
  XOR U2772 ( .A(n4065), .B(n4066), .Z(n251) );
  NOR U2773 ( .A(n4067), .B(n4065), .Z(n4066) );
  XOR U2774 ( .A(n4068), .B(n4069), .Z(n1391) );
  NOR U2775 ( .A(n4070), .B(n4068), .Z(n4069) );
  XOR U2776 ( .A(n4071), .B(n4072), .Z(n1392) );
  NOR U2777 ( .A(n4073), .B(n4071), .Z(n4072) );
  XOR U2778 ( .A(n4074), .B(n4075), .Z(n1393) );
  NOR U2779 ( .A(n4076), .B(n4074), .Z(n4075) );
  XOR U2780 ( .A(n4077), .B(n4078), .Z(n244) );
  NOR U2781 ( .A(n4079), .B(n4077), .Z(n4078) );
  XOR U2782 ( .A(n4080), .B(n4081), .Z(n238) );
  NOR U2783 ( .A(n4082), .B(n4080), .Z(n4081) );
  XOR U2784 ( .A(n4083), .B(n4084), .Z(n235) );
  NOR U2785 ( .A(n4085), .B(n4083), .Z(n4084) );
  XOR U2786 ( .A(n4086), .B(n4087), .Z(n233) );
  NOR U2787 ( .A(n4088), .B(n4086), .Z(n4087) );
  XOR U2788 ( .A(n4089), .B(n4090), .Z(n234) );
  NOR U2789 ( .A(n4091), .B(n4089), .Z(n4090) );
  XOR U2790 ( .A(n4092), .B(n4093), .Z(n1412) );
  NOR U2791 ( .A(n4094), .B(n4092), .Z(n4093) );
  XOR U2792 ( .A(n4095), .B(n4096), .Z(n1416) );
  NOR U2793 ( .A(n4097), .B(n4095), .Z(n4096) );
  XOR U2794 ( .A(n4098), .B(n4099), .Z(n223) );
  NOR U2795 ( .A(n4100), .B(n4098), .Z(n4099) );
  XOR U2796 ( .A(n4101), .B(n4102), .Z(n224) );
  NOR U2797 ( .A(n4103), .B(n4101), .Z(n4102) );
  XOR U2798 ( .A(n4104), .B(n4105), .Z(n1424) );
  NOR U2799 ( .A(n4106), .B(n4104), .Z(n4105) );
  XOR U2800 ( .A(n4107), .B(n4108), .Z(n1425) );
  NOR U2801 ( .A(n4109), .B(n4107), .Z(n4108) );
  XOR U2802 ( .A(n4110), .B(n4111), .Z(n1426) );
  NOR U2803 ( .A(n4112), .B(n4110), .Z(n4111) );
  XOR U2804 ( .A(n4113), .B(n4114), .Z(n217) );
  NOR U2805 ( .A(n4115), .B(n4113), .Z(n4114) );
  XOR U2806 ( .A(n4116), .B(n4117), .Z(n211) );
  NOR U2807 ( .A(n4118), .B(n4116), .Z(n4117) );
  XOR U2808 ( .A(n4119), .B(n4120), .Z(n208) );
  NOR U2809 ( .A(n4121), .B(n4119), .Z(n4120) );
  XOR U2810 ( .A(n4122), .B(n4123), .Z(n206) );
  NOR U2811 ( .A(n4124), .B(n4122), .Z(n4123) );
  XOR U2812 ( .A(n4125), .B(n4126), .Z(n207) );
  NOR U2813 ( .A(n4127), .B(n4125), .Z(n4126) );
  XOR U2814 ( .A(n4128), .B(n4129), .Z(n189) );
  NOR U2815 ( .A(n4130), .B(n4128), .Z(n4129) );
  XOR U2816 ( .A(n4131), .B(n4132), .Z(n190) );
  NOR U2817 ( .A(n4133), .B(n4131), .Z(n4132) );
  XOR U2818 ( .A(n4134), .B(n4135), .Z(n1449) );
  NOR U2819 ( .A(n4136), .B(n4134), .Z(n4135) );
  XOR U2820 ( .A(n4137), .B(n4138), .Z(n194) );
  NOR U2821 ( .A(n4139), .B(n4137), .Z(n4138) );
  IV U2822 ( .A(n173), .Z(n2741) );
  XNOR U2823 ( .A(n4140), .B(n4141), .Z(n173) );
  NOR U2824 ( .A(n4142), .B(n4140), .Z(n4141) );
  XOR U2825 ( .A(n4143), .B(n4144), .Z(n175) );
  NOR U2826 ( .A(n4145), .B(n4143), .Z(n4144) );
  XOR U2827 ( .A(n4146), .B(n4147), .Z(n179) );
  NOR U2828 ( .A(n4148), .B(n4146), .Z(n4147) );
  XNOR U2829 ( .A(n4149), .B(n4150), .Z(n181) );
  AND U2830 ( .A(n4151), .B(n4149), .Z(n4150) );
  XNOR U2831 ( .A(n4152), .B(n4153), .Z(n1450) );
  AND U2832 ( .A(n60), .B(n4152), .Z(n4153) );
  XNOR U2833 ( .A(n45), .B(n2737), .Z(n2739) );
  XOR U2834 ( .A(n2734), .B(n1475), .Z(n45) );
  XOR U2835 ( .A(n4154), .B(n1463), .Z(n1475) );
  XOR U2836 ( .A(n1464), .B(n1461), .Z(n1463) );
  XOR U2837 ( .A(n1462), .B(n1458), .Z(n1461) );
  XNOR U2838 ( .A(n1457), .B(n1484), .Z(n1458) );
  XNOR U2839 ( .A(n1483), .B(n2733), .Z(n1484) );
  XNOR U2840 ( .A(n2724), .B(n2732), .Z(n2733) );
  XNOR U2841 ( .A(n2723), .B(n2729), .Z(n2732) );
  XNOR U2842 ( .A(n2728), .B(n1493), .Z(n2729) );
  XNOR U2843 ( .A(n1492), .B(n2722), .Z(n1493) );
  XNOR U2844 ( .A(n2713), .B(n2721), .Z(n2722) );
  XNOR U2845 ( .A(n2712), .B(n2718), .Z(n2721) );
  XNOR U2846 ( .A(n2717), .B(n1502), .Z(n2718) );
  XNOR U2847 ( .A(n1501), .B(n2711), .Z(n1502) );
  XNOR U2848 ( .A(n2702), .B(n2710), .Z(n2711) );
  XNOR U2849 ( .A(n2701), .B(n2707), .Z(n2710) );
  XNOR U2850 ( .A(n2706), .B(n1511), .Z(n2707) );
  XNOR U2851 ( .A(n1510), .B(n2700), .Z(n1511) );
  XNOR U2852 ( .A(n2691), .B(n2699), .Z(n2700) );
  XNOR U2853 ( .A(n2690), .B(n2696), .Z(n2699) );
  XNOR U2854 ( .A(n2695), .B(n1520), .Z(n2696) );
  XNOR U2855 ( .A(n1519), .B(n2689), .Z(n1520) );
  XNOR U2856 ( .A(n2680), .B(n2688), .Z(n2689) );
  XNOR U2857 ( .A(n2679), .B(n2685), .Z(n2688) );
  XNOR U2858 ( .A(n2684), .B(n1529), .Z(n2685) );
  XNOR U2859 ( .A(n1528), .B(n2678), .Z(n1529) );
  XNOR U2860 ( .A(n2669), .B(n2677), .Z(n2678) );
  XNOR U2861 ( .A(n2668), .B(n2674), .Z(n2677) );
  XNOR U2862 ( .A(n2673), .B(n1538), .Z(n2674) );
  XNOR U2863 ( .A(n1537), .B(n2667), .Z(n1538) );
  XNOR U2864 ( .A(n2658), .B(n2666), .Z(n2667) );
  XNOR U2865 ( .A(n2657), .B(n2663), .Z(n2666) );
  XNOR U2866 ( .A(n2662), .B(n1547), .Z(n2663) );
  XNOR U2867 ( .A(n1546), .B(n2656), .Z(n1547) );
  XNOR U2868 ( .A(n2647), .B(n2655), .Z(n2656) );
  XNOR U2869 ( .A(n2646), .B(n2652), .Z(n2655) );
  XNOR U2870 ( .A(n2651), .B(n1556), .Z(n2652) );
  XNOR U2871 ( .A(n1555), .B(n2645), .Z(n1556) );
  XNOR U2872 ( .A(n2636), .B(n2644), .Z(n2645) );
  XNOR U2873 ( .A(n2635), .B(n2641), .Z(n2644) );
  XNOR U2874 ( .A(n2640), .B(n1565), .Z(n2641) );
  XNOR U2875 ( .A(n1564), .B(n2634), .Z(n1565) );
  XNOR U2876 ( .A(n2625), .B(n2633), .Z(n2634) );
  XNOR U2877 ( .A(n2624), .B(n2630), .Z(n2633) );
  XNOR U2878 ( .A(n2629), .B(n1574), .Z(n2630) );
  XNOR U2879 ( .A(n1573), .B(n2623), .Z(n1574) );
  XNOR U2880 ( .A(n2614), .B(n2622), .Z(n2623) );
  XNOR U2881 ( .A(n2613), .B(n2619), .Z(n2622) );
  XNOR U2882 ( .A(n2618), .B(n1583), .Z(n2619) );
  XNOR U2883 ( .A(n1582), .B(n2612), .Z(n1583) );
  XNOR U2884 ( .A(n2603), .B(n2611), .Z(n2612) );
  XNOR U2885 ( .A(n2602), .B(n2608), .Z(n2611) );
  XNOR U2886 ( .A(n2607), .B(n1592), .Z(n2608) );
  XNOR U2887 ( .A(n1591), .B(n2601), .Z(n1592) );
  XNOR U2888 ( .A(n2592), .B(n2600), .Z(n2601) );
  XNOR U2889 ( .A(n2591), .B(n2597), .Z(n2600) );
  XNOR U2890 ( .A(n2596), .B(n1601), .Z(n2597) );
  XNOR U2891 ( .A(n1600), .B(n2590), .Z(n1601) );
  XNOR U2892 ( .A(n2581), .B(n2589), .Z(n2590) );
  XNOR U2893 ( .A(n2580), .B(n2586), .Z(n2589) );
  XNOR U2894 ( .A(n2585), .B(n1610), .Z(n2586) );
  XNOR U2895 ( .A(n1609), .B(n2579), .Z(n1610) );
  XNOR U2896 ( .A(n2570), .B(n2578), .Z(n2579) );
  XNOR U2897 ( .A(n2569), .B(n2575), .Z(n2578) );
  XNOR U2898 ( .A(n2574), .B(n1619), .Z(n2575) );
  XNOR U2899 ( .A(n1618), .B(n2568), .Z(n1619) );
  XNOR U2900 ( .A(n2559), .B(n2567), .Z(n2568) );
  XNOR U2901 ( .A(n2558), .B(n2564), .Z(n2567) );
  XNOR U2902 ( .A(n2563), .B(n1628), .Z(n2564) );
  XNOR U2903 ( .A(n1627), .B(n2557), .Z(n1628) );
  XNOR U2904 ( .A(n2548), .B(n2556), .Z(n2557) );
  XNOR U2905 ( .A(n2547), .B(n2553), .Z(n2556) );
  XNOR U2906 ( .A(n2552), .B(n1637), .Z(n2553) );
  XNOR U2907 ( .A(n1636), .B(n2546), .Z(n1637) );
  XNOR U2908 ( .A(n2537), .B(n2545), .Z(n2546) );
  XNOR U2909 ( .A(n2536), .B(n2542), .Z(n2545) );
  XNOR U2910 ( .A(n2541), .B(n1646), .Z(n2542) );
  XNOR U2911 ( .A(n1645), .B(n2535), .Z(n1646) );
  XNOR U2912 ( .A(n2526), .B(n2534), .Z(n2535) );
  XNOR U2913 ( .A(n2525), .B(n2531), .Z(n2534) );
  XNOR U2914 ( .A(n2530), .B(n1655), .Z(n2531) );
  XNOR U2915 ( .A(n1654), .B(n2524), .Z(n1655) );
  XNOR U2916 ( .A(n2515), .B(n2523), .Z(n2524) );
  XNOR U2917 ( .A(n2514), .B(n2520), .Z(n2523) );
  XNOR U2918 ( .A(n2519), .B(n1664), .Z(n2520) );
  XNOR U2919 ( .A(n1663), .B(n2513), .Z(n1664) );
  XNOR U2920 ( .A(n2504), .B(n2512), .Z(n2513) );
  XNOR U2921 ( .A(n2503), .B(n2509), .Z(n2512) );
  XNOR U2922 ( .A(n2508), .B(n1673), .Z(n2509) );
  XNOR U2923 ( .A(n1672), .B(n2502), .Z(n1673) );
  XNOR U2924 ( .A(n2493), .B(n2501), .Z(n2502) );
  XNOR U2925 ( .A(n2492), .B(n2498), .Z(n2501) );
  XNOR U2926 ( .A(n2497), .B(n1682), .Z(n2498) );
  XNOR U2927 ( .A(n1681), .B(n2491), .Z(n1682) );
  XNOR U2928 ( .A(n2482), .B(n2490), .Z(n2491) );
  XNOR U2929 ( .A(n2481), .B(n2487), .Z(n2490) );
  XNOR U2930 ( .A(n2486), .B(n1691), .Z(n2487) );
  XNOR U2931 ( .A(n1690), .B(n2480), .Z(n1691) );
  XNOR U2932 ( .A(n2471), .B(n2479), .Z(n2480) );
  XNOR U2933 ( .A(n2470), .B(n2476), .Z(n2479) );
  XNOR U2934 ( .A(n2475), .B(n1700), .Z(n2476) );
  XNOR U2935 ( .A(n1699), .B(n2469), .Z(n1700) );
  XNOR U2936 ( .A(n2460), .B(n2468), .Z(n2469) );
  XNOR U2937 ( .A(n2459), .B(n2465), .Z(n2468) );
  XNOR U2938 ( .A(n2464), .B(n1709), .Z(n2465) );
  XNOR U2939 ( .A(n1708), .B(n2458), .Z(n1709) );
  XNOR U2940 ( .A(n2449), .B(n2457), .Z(n2458) );
  XNOR U2941 ( .A(n2448), .B(n2454), .Z(n2457) );
  XNOR U2942 ( .A(n2453), .B(n1718), .Z(n2454) );
  XNOR U2943 ( .A(n1717), .B(n2447), .Z(n1718) );
  XNOR U2944 ( .A(n2438), .B(n2446), .Z(n2447) );
  XNOR U2945 ( .A(n2437), .B(n2443), .Z(n2446) );
  XNOR U2946 ( .A(n2442), .B(n1727), .Z(n2443) );
  XNOR U2947 ( .A(n1726), .B(n2436), .Z(n1727) );
  XNOR U2948 ( .A(n2427), .B(n2435), .Z(n2436) );
  XNOR U2949 ( .A(n2426), .B(n2432), .Z(n2435) );
  XNOR U2950 ( .A(n2431), .B(n1736), .Z(n2432) );
  XNOR U2951 ( .A(n1735), .B(n2425), .Z(n1736) );
  XNOR U2952 ( .A(n2416), .B(n2424), .Z(n2425) );
  XNOR U2953 ( .A(n2415), .B(n2421), .Z(n2424) );
  XNOR U2954 ( .A(n2420), .B(n1745), .Z(n2421) );
  XNOR U2955 ( .A(n1744), .B(n2414), .Z(n1745) );
  XNOR U2956 ( .A(n2405), .B(n2413), .Z(n2414) );
  XNOR U2957 ( .A(n2404), .B(n2410), .Z(n2413) );
  XNOR U2958 ( .A(n2409), .B(n1754), .Z(n2410) );
  XNOR U2959 ( .A(n1753), .B(n2403), .Z(n1754) );
  XNOR U2960 ( .A(n2394), .B(n2402), .Z(n2403) );
  XNOR U2961 ( .A(n2393), .B(n2399), .Z(n2402) );
  XNOR U2962 ( .A(n2398), .B(n1763), .Z(n2399) );
  XNOR U2963 ( .A(n1762), .B(n2392), .Z(n1763) );
  XNOR U2964 ( .A(n2383), .B(n2391), .Z(n2392) );
  XNOR U2965 ( .A(n2382), .B(n2388), .Z(n2391) );
  XNOR U2966 ( .A(n2387), .B(n1772), .Z(n2388) );
  XNOR U2967 ( .A(n1771), .B(n2381), .Z(n1772) );
  XNOR U2968 ( .A(n2372), .B(n2380), .Z(n2381) );
  XNOR U2969 ( .A(n2371), .B(n2377), .Z(n2380) );
  XNOR U2970 ( .A(n2376), .B(n1781), .Z(n2377) );
  XNOR U2971 ( .A(n1780), .B(n2370), .Z(n1781) );
  XNOR U2972 ( .A(n2361), .B(n2369), .Z(n2370) );
  XNOR U2973 ( .A(n2360), .B(n2366), .Z(n2369) );
  XNOR U2974 ( .A(n2365), .B(n1790), .Z(n2366) );
  XNOR U2975 ( .A(n1789), .B(n2359), .Z(n1790) );
  XNOR U2976 ( .A(n2350), .B(n2358), .Z(n2359) );
  XNOR U2977 ( .A(n2349), .B(n2355), .Z(n2358) );
  XNOR U2978 ( .A(n2354), .B(n1799), .Z(n2355) );
  XNOR U2979 ( .A(n1798), .B(n2348), .Z(n1799) );
  XNOR U2980 ( .A(n2339), .B(n2347), .Z(n2348) );
  XNOR U2981 ( .A(n2338), .B(n2344), .Z(n2347) );
  XNOR U2982 ( .A(n2343), .B(n1808), .Z(n2344) );
  XNOR U2983 ( .A(n1807), .B(n2337), .Z(n1808) );
  XNOR U2984 ( .A(n2328), .B(n2336), .Z(n2337) );
  XNOR U2985 ( .A(n2327), .B(n2333), .Z(n2336) );
  XNOR U2986 ( .A(n2332), .B(n1817), .Z(n2333) );
  XNOR U2987 ( .A(n1816), .B(n2326), .Z(n1817) );
  XNOR U2988 ( .A(n2317), .B(n2325), .Z(n2326) );
  XNOR U2989 ( .A(n2316), .B(n2322), .Z(n2325) );
  XNOR U2990 ( .A(n2321), .B(n1826), .Z(n2322) );
  XNOR U2991 ( .A(n1825), .B(n2315), .Z(n1826) );
  XNOR U2992 ( .A(n2306), .B(n2314), .Z(n2315) );
  XNOR U2993 ( .A(n2305), .B(n2311), .Z(n2314) );
  XNOR U2994 ( .A(n2310), .B(n1835), .Z(n2311) );
  XNOR U2995 ( .A(n1834), .B(n2304), .Z(n1835) );
  XNOR U2996 ( .A(n2295), .B(n2303), .Z(n2304) );
  XNOR U2997 ( .A(n2294), .B(n2300), .Z(n2303) );
  XNOR U2998 ( .A(n2299), .B(n1844), .Z(n2300) );
  XNOR U2999 ( .A(n1843), .B(n2293), .Z(n1844) );
  XNOR U3000 ( .A(n2284), .B(n2292), .Z(n2293) );
  XNOR U3001 ( .A(n2283), .B(n2289), .Z(n2292) );
  XNOR U3002 ( .A(n2288), .B(n1853), .Z(n2289) );
  XNOR U3003 ( .A(n1852), .B(n2282), .Z(n1853) );
  XNOR U3004 ( .A(n2273), .B(n2281), .Z(n2282) );
  XNOR U3005 ( .A(n2272), .B(n2278), .Z(n2281) );
  XNOR U3006 ( .A(n2277), .B(n1862), .Z(n2278) );
  XNOR U3007 ( .A(n1861), .B(n2271), .Z(n1862) );
  XNOR U3008 ( .A(n2262), .B(n2270), .Z(n2271) );
  XNOR U3009 ( .A(n2261), .B(n2267), .Z(n2270) );
  XNOR U3010 ( .A(n2266), .B(n1871), .Z(n2267) );
  XNOR U3011 ( .A(n1870), .B(n2260), .Z(n1871) );
  XNOR U3012 ( .A(n2251), .B(n2259), .Z(n2260) );
  XNOR U3013 ( .A(n2250), .B(n2256), .Z(n2259) );
  XNOR U3014 ( .A(n2255), .B(n1880), .Z(n2256) );
  XNOR U3015 ( .A(n1879), .B(n2249), .Z(n1880) );
  XNOR U3016 ( .A(n2240), .B(n2248), .Z(n2249) );
  XNOR U3017 ( .A(n2239), .B(n2245), .Z(n2248) );
  XNOR U3018 ( .A(n2244), .B(n1889), .Z(n2245) );
  XNOR U3019 ( .A(n1888), .B(n2238), .Z(n1889) );
  XNOR U3020 ( .A(n2229), .B(n2237), .Z(n2238) );
  XNOR U3021 ( .A(n2228), .B(n2234), .Z(n2237) );
  XNOR U3022 ( .A(n2233), .B(n1898), .Z(n2234) );
  XNOR U3023 ( .A(n1897), .B(n2227), .Z(n1898) );
  XNOR U3024 ( .A(n2218), .B(n2226), .Z(n2227) );
  XNOR U3025 ( .A(n2217), .B(n2223), .Z(n2226) );
  XNOR U3026 ( .A(n2222), .B(n1907), .Z(n2223) );
  XNOR U3027 ( .A(n1906), .B(n2216), .Z(n1907) );
  XNOR U3028 ( .A(n2207), .B(n2215), .Z(n2216) );
  XNOR U3029 ( .A(n2206), .B(n2212), .Z(n2215) );
  XNOR U3030 ( .A(n2211), .B(n1916), .Z(n2212) );
  XNOR U3031 ( .A(n1915), .B(n2205), .Z(n1916) );
  XNOR U3032 ( .A(n2196), .B(n2204), .Z(n2205) );
  XNOR U3033 ( .A(n2195), .B(n2201), .Z(n2204) );
  XNOR U3034 ( .A(n2200), .B(n1925), .Z(n2201) );
  XNOR U3035 ( .A(n1924), .B(n2194), .Z(n1925) );
  XNOR U3036 ( .A(n2185), .B(n2193), .Z(n2194) );
  XNOR U3037 ( .A(n2184), .B(n2190), .Z(n2193) );
  XNOR U3038 ( .A(n2189), .B(n1934), .Z(n2190) );
  XNOR U3039 ( .A(n1933), .B(n2183), .Z(n1934) );
  XNOR U3040 ( .A(n2174), .B(n2182), .Z(n2183) );
  XNOR U3041 ( .A(n2173), .B(n2179), .Z(n2182) );
  XNOR U3042 ( .A(n2178), .B(n1943), .Z(n2179) );
  XNOR U3043 ( .A(n1942), .B(n2172), .Z(n1943) );
  XNOR U3044 ( .A(n2163), .B(n2171), .Z(n2172) );
  XNOR U3045 ( .A(n2162), .B(n2168), .Z(n2171) );
  XNOR U3046 ( .A(n2167), .B(n1952), .Z(n2168) );
  XNOR U3047 ( .A(n1951), .B(n2161), .Z(n1952) );
  XNOR U3048 ( .A(n2152), .B(n2160), .Z(n2161) );
  XNOR U3049 ( .A(n2151), .B(n2157), .Z(n2160) );
  XNOR U3050 ( .A(n2156), .B(n1961), .Z(n2157) );
  XNOR U3051 ( .A(n1960), .B(n2150), .Z(n1961) );
  XNOR U3052 ( .A(n2141), .B(n2149), .Z(n2150) );
  XNOR U3053 ( .A(n2140), .B(n2146), .Z(n2149) );
  XNOR U3054 ( .A(n2145), .B(n1970), .Z(n2146) );
  XNOR U3055 ( .A(n1969), .B(n2139), .Z(n1970) );
  XNOR U3056 ( .A(n2130), .B(n2138), .Z(n2139) );
  XNOR U3057 ( .A(n2129), .B(n2135), .Z(n2138) );
  XNOR U3058 ( .A(n2134), .B(n1979), .Z(n2135) );
  XNOR U3059 ( .A(n1978), .B(n2128), .Z(n1979) );
  XNOR U3060 ( .A(n2119), .B(n2127), .Z(n2128) );
  XNOR U3061 ( .A(n2118), .B(n2124), .Z(n2127) );
  XNOR U3062 ( .A(n2123), .B(n1988), .Z(n2124) );
  XNOR U3063 ( .A(n1987), .B(n2117), .Z(n1988) );
  XNOR U3064 ( .A(n2108), .B(n2116), .Z(n2117) );
  XNOR U3065 ( .A(n2107), .B(n2113), .Z(n2116) );
  XNOR U3066 ( .A(n2112), .B(n1997), .Z(n2113) );
  XNOR U3067 ( .A(n1996), .B(n2106), .Z(n1997) );
  XNOR U3068 ( .A(n2097), .B(n2105), .Z(n2106) );
  XNOR U3069 ( .A(n2096), .B(n2102), .Z(n2105) );
  XNOR U3070 ( .A(n2101), .B(n2006), .Z(n2102) );
  XNOR U3071 ( .A(n2005), .B(n2095), .Z(n2006) );
  XNOR U3072 ( .A(n2086), .B(n2094), .Z(n2095) );
  XNOR U3073 ( .A(n2085), .B(n2091), .Z(n2094) );
  XNOR U3074 ( .A(n2090), .B(n2015), .Z(n2091) );
  XNOR U3075 ( .A(n2014), .B(n2084), .Z(n2015) );
  XNOR U3076 ( .A(n2075), .B(n2083), .Z(n2084) );
  XNOR U3077 ( .A(n2074), .B(n2080), .Z(n2083) );
  XNOR U3078 ( .A(n2079), .B(n2062), .Z(n2080) );
  XNOR U3079 ( .A(n2021), .B(n2073), .Z(n2062) );
  XNOR U3080 ( .A(n2064), .B(n2072), .Z(n2073) );
  XNOR U3081 ( .A(n2063), .B(n2069), .Z(n2072) );
  XNOR U3082 ( .A(n2068), .B(n2052), .Z(n2069) );
  XNOR U3083 ( .A(n2024), .B(n2061), .Z(n2052) );
  XNOR U3084 ( .A(n2048), .B(n2058), .Z(n2061) );
  XNOR U3085 ( .A(n2051), .B(n2057), .Z(n2058) );
  XNOR U3086 ( .A(n2020), .B(n2047), .Z(n2057) );
  XNOR U3087 ( .A(n2030), .B(n2046), .Z(n2047) );
  XNOR U3088 ( .A(n2033), .B(n2043), .Z(n2046) );
  XOR U3089 ( .A(n2032), .B(n2040), .Z(n2043) );
  XOR U3090 ( .A(n2041), .B(n2039), .Z(n2040) );
  XNOR U3091 ( .A(n4155), .B(n4156), .Z(n2039) );
  XOR U3092 ( .A(n4157), .B(n4158), .Z(n4156) );
  XNOR U3093 ( .A(n4159), .B(n4160), .Z(n4158) );
  NOR U3094 ( .A(n4161), .B(n4160), .Z(n4159) );
  XOR U3095 ( .A(n4162), .B(n4163), .Z(n4157) );
  NOR U3096 ( .A(n4164), .B(n4165), .Z(n4163) );
  AND U3097 ( .A(n4166), .B(n4167), .Z(n4162) );
  XOR U3098 ( .A(n4168), .B(n4169), .Z(n4155) );
  XOR U3099 ( .A(n4170), .B(n4171), .Z(n4169) );
  XOR U3100 ( .A(n4172), .B(n4173), .Z(n4171) );
  XOR U3101 ( .A(n4174), .B(n4175), .Z(n4173) );
  XNOR U3102 ( .A(n4176), .B(n4177), .Z(n4175) );
  NOR U3103 ( .A(n4178), .B(n4177), .Z(n4176) );
  XOR U3104 ( .A(n4179), .B(n4180), .Z(n4174) );
  XOR U3105 ( .A(n4181), .B(n4182), .Z(n4180) );
  XOR U3106 ( .A(n4183), .B(n4184), .Z(n4182) );
  XNOR U3107 ( .A(n4185), .B(n4186), .Z(n4184) );
  NOR U3108 ( .A(n4187), .B(n4186), .Z(n4185) );
  XOR U3109 ( .A(n4188), .B(n4189), .Z(n4183) );
  XOR U3110 ( .A(n4190), .B(n4191), .Z(n4189) );
  XOR U3111 ( .A(n4192), .B(n4193), .Z(n4191) );
  XNOR U3112 ( .A(n4194), .B(n4195), .Z(n4193) );
  NOR U3113 ( .A(n4196), .B(n4195), .Z(n4194) );
  XOR U3114 ( .A(n4197), .B(n4198), .Z(n4192) );
  XOR U3115 ( .A(n4199), .B(n4200), .Z(n4198) );
  XOR U3116 ( .A(n4201), .B(n4202), .Z(n4200) );
  XNOR U3117 ( .A(n4203), .B(n4204), .Z(n4202) );
  NOR U3118 ( .A(n4205), .B(n4204), .Z(n4203) );
  XOR U3119 ( .A(n4206), .B(n4207), .Z(n4201) );
  XOR U3120 ( .A(n4208), .B(n4209), .Z(n4207) );
  XOR U3121 ( .A(n4210), .B(n4211), .Z(n4209) );
  XNOR U3122 ( .A(n4212), .B(n4213), .Z(n4211) );
  NOR U3123 ( .A(n4214), .B(n4213), .Z(n4212) );
  XOR U3124 ( .A(n4215), .B(n4216), .Z(n4210) );
  XOR U3125 ( .A(n4217), .B(n4218), .Z(n4216) );
  XOR U3126 ( .A(n4219), .B(n4220), .Z(n4218) );
  XNOR U3127 ( .A(n4221), .B(n4222), .Z(n4220) );
  NOR U3128 ( .A(n4223), .B(n4222), .Z(n4221) );
  XOR U3129 ( .A(n4224), .B(n4225), .Z(n4219) );
  XOR U3130 ( .A(n4226), .B(n4227), .Z(n4225) );
  XOR U3131 ( .A(n4228), .B(n4229), .Z(n4227) );
  XNOR U3132 ( .A(n4230), .B(n4231), .Z(n4229) );
  NOR U3133 ( .A(n4232), .B(n4231), .Z(n4230) );
  XOR U3134 ( .A(n4233), .B(n4234), .Z(n4228) );
  XOR U3135 ( .A(n4235), .B(n4236), .Z(n4234) );
  XOR U3136 ( .A(n4237), .B(n4238), .Z(n4236) );
  XNOR U3137 ( .A(n4239), .B(n4240), .Z(n4238) );
  NOR U3138 ( .A(n4241), .B(n4240), .Z(n4239) );
  XOR U3139 ( .A(n4242), .B(n4243), .Z(n4237) );
  XOR U3140 ( .A(n4244), .B(n4245), .Z(n4243) );
  XOR U3141 ( .A(n4246), .B(n4247), .Z(n4245) );
  XNOR U3142 ( .A(n4248), .B(n4249), .Z(n4247) );
  NOR U3143 ( .A(n4250), .B(n4249), .Z(n4248) );
  XOR U3144 ( .A(n4251), .B(n4252), .Z(n4246) );
  XOR U3145 ( .A(n4253), .B(n4254), .Z(n4252) );
  XOR U3146 ( .A(n4255), .B(n4256), .Z(n4254) );
  XNOR U3147 ( .A(n4257), .B(n4258), .Z(n4256) );
  NOR U3148 ( .A(n4259), .B(n4258), .Z(n4257) );
  XOR U3149 ( .A(n4260), .B(n4261), .Z(n4255) );
  XOR U3150 ( .A(n4262), .B(n4263), .Z(n4261) );
  XOR U3151 ( .A(n4264), .B(n4265), .Z(n4263) );
  XNOR U3152 ( .A(n4266), .B(n4267), .Z(n4265) );
  NOR U3153 ( .A(n4268), .B(n4267), .Z(n4266) );
  XOR U3154 ( .A(n4269), .B(n4270), .Z(n4264) );
  XOR U3155 ( .A(n4271), .B(n4272), .Z(n4270) );
  XOR U3156 ( .A(n4273), .B(n4274), .Z(n4272) );
  XNOR U3157 ( .A(n4275), .B(n4276), .Z(n4274) );
  NOR U3158 ( .A(n4277), .B(n4276), .Z(n4275) );
  XOR U3159 ( .A(n4278), .B(n4279), .Z(n4273) );
  XOR U3160 ( .A(n4280), .B(n4281), .Z(n4279) );
  XOR U3161 ( .A(n4282), .B(n4283), .Z(n4281) );
  XNOR U3162 ( .A(n4284), .B(n4285), .Z(n4283) );
  NOR U3163 ( .A(n4286), .B(n4285), .Z(n4284) );
  XOR U3164 ( .A(n4287), .B(n4288), .Z(n4282) );
  XOR U3165 ( .A(n4289), .B(n4290), .Z(n4288) );
  XOR U3166 ( .A(n4291), .B(n4292), .Z(n4290) );
  XNOR U3167 ( .A(n4293), .B(n4294), .Z(n4292) );
  NOR U3168 ( .A(n4295), .B(n4294), .Z(n4293) );
  XOR U3169 ( .A(n4296), .B(n4297), .Z(n4291) );
  XOR U3170 ( .A(n4298), .B(n4299), .Z(n4297) );
  XOR U3171 ( .A(n4300), .B(n4301), .Z(n4299) );
  XNOR U3172 ( .A(n4302), .B(n4303), .Z(n4301) );
  NOR U3173 ( .A(n4304), .B(n4303), .Z(n4302) );
  XOR U3174 ( .A(n4305), .B(n4306), .Z(n4300) );
  XOR U3175 ( .A(n4307), .B(n4308), .Z(n4306) );
  XOR U3176 ( .A(n4309), .B(n4310), .Z(n4308) );
  XNOR U3177 ( .A(n4311), .B(n4312), .Z(n4310) );
  NOR U3178 ( .A(n4313), .B(n4312), .Z(n4311) );
  XOR U3179 ( .A(n4314), .B(n4315), .Z(n4309) );
  XOR U3180 ( .A(n4316), .B(n4317), .Z(n4315) );
  XOR U3181 ( .A(n4318), .B(n4319), .Z(n4317) );
  XNOR U3182 ( .A(n4320), .B(n4321), .Z(n4319) );
  NOR U3183 ( .A(n4322), .B(n4321), .Z(n4320) );
  XOR U3184 ( .A(n4323), .B(n4324), .Z(n4318) );
  XOR U3185 ( .A(n4325), .B(n4326), .Z(n4324) );
  XOR U3186 ( .A(n4327), .B(n4328), .Z(n4326) );
  XNOR U3187 ( .A(n4329), .B(n4330), .Z(n4328) );
  NOR U3188 ( .A(n4331), .B(n4330), .Z(n4329) );
  XOR U3189 ( .A(n4332), .B(n4333), .Z(n4327) );
  XOR U3190 ( .A(n4334), .B(n4335), .Z(n4333) );
  XOR U3191 ( .A(n4336), .B(n4337), .Z(n4335) );
  XNOR U3192 ( .A(n4338), .B(n4339), .Z(n4337) );
  NOR U3193 ( .A(n4340), .B(n4339), .Z(n4338) );
  XOR U3194 ( .A(n4341), .B(n4342), .Z(n4336) );
  XOR U3195 ( .A(n4343), .B(n4344), .Z(n4342) );
  XOR U3196 ( .A(n4345), .B(n4346), .Z(n4344) );
  XNOR U3197 ( .A(n4347), .B(n4348), .Z(n4346) );
  NOR U3198 ( .A(n4349), .B(n4348), .Z(n4347) );
  XOR U3199 ( .A(n4350), .B(n4351), .Z(n4345) );
  XOR U3200 ( .A(n4352), .B(n4353), .Z(n4351) );
  XOR U3201 ( .A(n4354), .B(n4355), .Z(n4353) );
  XNOR U3202 ( .A(n4356), .B(n4357), .Z(n4355) );
  NOR U3203 ( .A(n4358), .B(n4357), .Z(n4356) );
  XOR U3204 ( .A(n4359), .B(n4360), .Z(n4354) );
  XOR U3205 ( .A(n4361), .B(n4362), .Z(n4360) );
  XOR U3206 ( .A(n4363), .B(n4364), .Z(n4362) );
  XNOR U3207 ( .A(n4365), .B(n4366), .Z(n4364) );
  NOR U3208 ( .A(n4367), .B(n4366), .Z(n4365) );
  XOR U3209 ( .A(n4368), .B(n4369), .Z(n4363) );
  XOR U3210 ( .A(n4370), .B(n4371), .Z(n4369) );
  XOR U3211 ( .A(n4372), .B(n4373), .Z(n4371) );
  XNOR U3212 ( .A(n4374), .B(n4375), .Z(n4373) );
  NOR U3213 ( .A(n4376), .B(n4375), .Z(n4374) );
  XOR U3214 ( .A(n4377), .B(n4378), .Z(n4372) );
  XOR U3215 ( .A(n4379), .B(n4380), .Z(n4378) );
  XOR U3216 ( .A(n4381), .B(n4382), .Z(n4380) );
  XNOR U3217 ( .A(n4383), .B(n4384), .Z(n4382) );
  NOR U3218 ( .A(n4385), .B(n4384), .Z(n4383) );
  XOR U3219 ( .A(n4386), .B(n4387), .Z(n4381) );
  XOR U3220 ( .A(n4388), .B(n4389), .Z(n4387) );
  XOR U3221 ( .A(n4390), .B(n4391), .Z(n4389) );
  XNOR U3222 ( .A(n4392), .B(n4393), .Z(n4391) );
  NOR U3223 ( .A(n4394), .B(n4393), .Z(n4392) );
  XOR U3224 ( .A(n4395), .B(n4396), .Z(n4390) );
  XOR U3225 ( .A(n4397), .B(n4398), .Z(n4396) );
  XOR U3226 ( .A(n4399), .B(n4400), .Z(n4398) );
  XNOR U3227 ( .A(n4401), .B(n4402), .Z(n4400) );
  NOR U3228 ( .A(n4403), .B(n4402), .Z(n4401) );
  XOR U3229 ( .A(n4404), .B(n4405), .Z(n4399) );
  XOR U3230 ( .A(n4406), .B(n4407), .Z(n4405) );
  XOR U3231 ( .A(n4408), .B(n4409), .Z(n4407) );
  XNOR U3232 ( .A(n4410), .B(n4411), .Z(n4409) );
  NOR U3233 ( .A(n4412), .B(n4411), .Z(n4410) );
  XOR U3234 ( .A(n4413), .B(n4414), .Z(n4408) );
  XOR U3235 ( .A(n4415), .B(n4416), .Z(n4414) );
  XOR U3236 ( .A(n4417), .B(n4418), .Z(n4416) );
  XNOR U3237 ( .A(n4419), .B(n4420), .Z(n4418) );
  NOR U3238 ( .A(n4421), .B(n4420), .Z(n4419) );
  XOR U3239 ( .A(n4422), .B(n4423), .Z(n4417) );
  XOR U3240 ( .A(n4424), .B(n4425), .Z(n4423) );
  XOR U3241 ( .A(n4426), .B(n4427), .Z(n4425) );
  XNOR U3242 ( .A(n4428), .B(n4429), .Z(n4427) );
  NOR U3243 ( .A(n4430), .B(n4429), .Z(n4428) );
  XOR U3244 ( .A(n4431), .B(n4432), .Z(n4426) );
  XOR U3245 ( .A(n4433), .B(n4434), .Z(n4432) );
  XOR U3246 ( .A(n4435), .B(n4436), .Z(n4434) );
  XOR U3247 ( .A(n4437), .B(n4438), .Z(n4433) );
  XNOR U3248 ( .A(n4439), .B(n4440), .Z(n4438) );
  XOR U3249 ( .A(n4441), .B(n4442), .Z(n4440) );
  XOR U3250 ( .A(n4443), .B(n4444), .Z(n4442) );
  XNOR U3251 ( .A(n4445), .B(n4446), .Z(n4444) );
  XOR U3252 ( .A(n4447), .B(n4448), .Z(n4443) );
  XOR U3253 ( .A(n4449), .B(n4450), .Z(n4441) );
  XOR U3254 ( .A(n4451), .B(n4452), .Z(n4450) );
  AND U3255 ( .A(n4453), .B(n4454), .Z(n4452) );
  XOR U3256 ( .A(n4446), .B(n4455), .Z(n4453) );
  XOR U3257 ( .A(n4456), .B(n4457), .Z(n4446) );
  AND U3258 ( .A(n4455), .B(n4456), .Z(n4457) );
  NOR U3259 ( .A(n4458), .B(n4447), .Z(n4451) );
  XOR U3260 ( .A(n4459), .B(n4460), .Z(n4449) );
  NOR U3261 ( .A(n4461), .B(n4448), .Z(n4460) );
  NOR U3262 ( .A(n4462), .B(n4445), .Z(n4459) );
  XNOR U3263 ( .A(n4463), .B(n4464), .Z(n4437) );
  XNOR U3264 ( .A(n4465), .B(n4466), .Z(n4464) );
  NOR U3265 ( .A(n4467), .B(n4439), .Z(n4465) );
  XOR U3266 ( .A(n4468), .B(n4469), .Z(n4431) );
  XOR U3267 ( .A(n4470), .B(n4471), .Z(n4469) );
  NOR U3268 ( .A(n4472), .B(n4435), .Z(n4471) );
  NOR U3269 ( .A(n4473), .B(n4466), .Z(n4470) );
  XOR U3270 ( .A(n4474), .B(n4475), .Z(n4468) );
  NOR U3271 ( .A(n4476), .B(n4463), .Z(n4475) );
  NOR U3272 ( .A(n4477), .B(n4436), .Z(n4474) );
  XOR U3273 ( .A(n4478), .B(n4479), .Z(n4424) );
  XOR U3274 ( .A(n4480), .B(n4481), .Z(n4422) );
  XNOR U3275 ( .A(n4482), .B(n4483), .Z(n4481) );
  NOR U3276 ( .A(n4484), .B(n4483), .Z(n4482) );
  XOR U3277 ( .A(n4485), .B(n4486), .Z(n4480) );
  NOR U3278 ( .A(n4487), .B(n4478), .Z(n4486) );
  NOR U3279 ( .A(n4488), .B(n4479), .Z(n4485) );
  XOR U3280 ( .A(n4489), .B(n4490), .Z(n4415) );
  XOR U3281 ( .A(n4491), .B(n4492), .Z(n4413) );
  XNOR U3282 ( .A(n4493), .B(n4494), .Z(n4492) );
  NOR U3283 ( .A(n4495), .B(n4494), .Z(n4493) );
  XOR U3284 ( .A(n4496), .B(n4497), .Z(n4491) );
  NOR U3285 ( .A(n4498), .B(n4489), .Z(n4497) );
  NOR U3286 ( .A(n4499), .B(n4490), .Z(n4496) );
  XOR U3287 ( .A(n4500), .B(n4501), .Z(n4406) );
  XOR U3288 ( .A(n4502), .B(n4503), .Z(n4404) );
  XNOR U3289 ( .A(n4504), .B(n4505), .Z(n4503) );
  NOR U3290 ( .A(n4506), .B(n4505), .Z(n4504) );
  XOR U3291 ( .A(n4507), .B(n4508), .Z(n4502) );
  NOR U3292 ( .A(n4509), .B(n4500), .Z(n4508) );
  NOR U3293 ( .A(n4510), .B(n4501), .Z(n4507) );
  XOR U3294 ( .A(n4511), .B(n4512), .Z(n4397) );
  XOR U3295 ( .A(n4513), .B(n4514), .Z(n4395) );
  XNOR U3296 ( .A(n4515), .B(n4516), .Z(n4514) );
  NOR U3297 ( .A(n4517), .B(n4516), .Z(n4515) );
  XOR U3298 ( .A(n4518), .B(n4519), .Z(n4513) );
  NOR U3299 ( .A(n4520), .B(n4511), .Z(n4519) );
  NOR U3300 ( .A(n4521), .B(n4512), .Z(n4518) );
  XOR U3301 ( .A(n4522), .B(n4523), .Z(n4388) );
  XOR U3302 ( .A(n4524), .B(n4525), .Z(n4386) );
  XNOR U3303 ( .A(n4526), .B(n4527), .Z(n4525) );
  NOR U3304 ( .A(n4528), .B(n4527), .Z(n4526) );
  XOR U3305 ( .A(n4529), .B(n4530), .Z(n4524) );
  NOR U3306 ( .A(n4531), .B(n4522), .Z(n4530) );
  NOR U3307 ( .A(n4532), .B(n4523), .Z(n4529) );
  XOR U3308 ( .A(n4533), .B(n4534), .Z(n4379) );
  XOR U3309 ( .A(n4535), .B(n4536), .Z(n4377) );
  XNOR U3310 ( .A(n4537), .B(n4538), .Z(n4536) );
  NOR U3311 ( .A(n4539), .B(n4538), .Z(n4537) );
  XOR U3312 ( .A(n4540), .B(n4541), .Z(n4535) );
  NOR U3313 ( .A(n4542), .B(n4533), .Z(n4541) );
  NOR U3314 ( .A(n4543), .B(n4534), .Z(n4540) );
  XOR U3315 ( .A(n4544), .B(n4545), .Z(n4370) );
  XOR U3316 ( .A(n4546), .B(n4547), .Z(n4368) );
  XNOR U3317 ( .A(n4548), .B(n4549), .Z(n4547) );
  NOR U3318 ( .A(n4550), .B(n4549), .Z(n4548) );
  XOR U3319 ( .A(n4551), .B(n4552), .Z(n4546) );
  NOR U3320 ( .A(n4553), .B(n4544), .Z(n4552) );
  NOR U3321 ( .A(n4554), .B(n4545), .Z(n4551) );
  XOR U3322 ( .A(n4555), .B(n4556), .Z(n4361) );
  XOR U3323 ( .A(n4557), .B(n4558), .Z(n4359) );
  XNOR U3324 ( .A(n4559), .B(n4560), .Z(n4558) );
  NOR U3325 ( .A(n4561), .B(n4560), .Z(n4559) );
  XOR U3326 ( .A(n4562), .B(n4563), .Z(n4557) );
  NOR U3327 ( .A(n4564), .B(n4555), .Z(n4563) );
  NOR U3328 ( .A(n4565), .B(n4556), .Z(n4562) );
  XOR U3329 ( .A(n4566), .B(n4567), .Z(n4352) );
  XOR U3330 ( .A(n4568), .B(n4569), .Z(n4350) );
  XNOR U3331 ( .A(n4570), .B(n4571), .Z(n4569) );
  NOR U3332 ( .A(n4572), .B(n4571), .Z(n4570) );
  XOR U3333 ( .A(n4573), .B(n4574), .Z(n4568) );
  NOR U3334 ( .A(n4575), .B(n4566), .Z(n4574) );
  NOR U3335 ( .A(n4576), .B(n4567), .Z(n4573) );
  XOR U3336 ( .A(n4577), .B(n4578), .Z(n4343) );
  XOR U3337 ( .A(n4579), .B(n4580), .Z(n4341) );
  XNOR U3338 ( .A(n4581), .B(n4582), .Z(n4580) );
  NOR U3339 ( .A(n4583), .B(n4582), .Z(n4581) );
  XOR U3340 ( .A(n4584), .B(n4585), .Z(n4579) );
  NOR U3341 ( .A(n4586), .B(n4577), .Z(n4585) );
  NOR U3342 ( .A(n4587), .B(n4578), .Z(n4584) );
  XOR U3343 ( .A(n4588), .B(n4589), .Z(n4334) );
  XOR U3344 ( .A(n4590), .B(n4591), .Z(n4332) );
  XNOR U3345 ( .A(n4592), .B(n4593), .Z(n4591) );
  NOR U3346 ( .A(n4594), .B(n4593), .Z(n4592) );
  XOR U3347 ( .A(n4595), .B(n4596), .Z(n4590) );
  NOR U3348 ( .A(n4597), .B(n4588), .Z(n4596) );
  NOR U3349 ( .A(n4598), .B(n4589), .Z(n4595) );
  XOR U3350 ( .A(n4599), .B(n4600), .Z(n4325) );
  XOR U3351 ( .A(n4601), .B(n4602), .Z(n4323) );
  XNOR U3352 ( .A(n4603), .B(n4604), .Z(n4602) );
  NOR U3353 ( .A(n4605), .B(n4604), .Z(n4603) );
  XOR U3354 ( .A(n4606), .B(n4607), .Z(n4601) );
  NOR U3355 ( .A(n4608), .B(n4599), .Z(n4607) );
  NOR U3356 ( .A(n4609), .B(n4600), .Z(n4606) );
  XOR U3357 ( .A(n4610), .B(n4611), .Z(n4316) );
  XOR U3358 ( .A(n4612), .B(n4613), .Z(n4314) );
  XNOR U3359 ( .A(n4614), .B(n4615), .Z(n4613) );
  NOR U3360 ( .A(n4616), .B(n4615), .Z(n4614) );
  XOR U3361 ( .A(n4617), .B(n4618), .Z(n4612) );
  NOR U3362 ( .A(n4619), .B(n4610), .Z(n4618) );
  NOR U3363 ( .A(n4620), .B(n4611), .Z(n4617) );
  XOR U3364 ( .A(n4621), .B(n4622), .Z(n4307) );
  XOR U3365 ( .A(n4623), .B(n4624), .Z(n4305) );
  XNOR U3366 ( .A(n4625), .B(n4626), .Z(n4624) );
  NOR U3367 ( .A(n4627), .B(n4626), .Z(n4625) );
  XOR U3368 ( .A(n4628), .B(n4629), .Z(n4623) );
  NOR U3369 ( .A(n4630), .B(n4621), .Z(n4629) );
  NOR U3370 ( .A(n4631), .B(n4622), .Z(n4628) );
  XOR U3371 ( .A(n4632), .B(n4633), .Z(n4298) );
  XOR U3372 ( .A(n4634), .B(n4635), .Z(n4296) );
  XNOR U3373 ( .A(n4636), .B(n4637), .Z(n4635) );
  NOR U3374 ( .A(n4638), .B(n4637), .Z(n4636) );
  XOR U3375 ( .A(n4639), .B(n4640), .Z(n4634) );
  NOR U3376 ( .A(n4641), .B(n4632), .Z(n4640) );
  NOR U3377 ( .A(n4642), .B(n4633), .Z(n4639) );
  XOR U3378 ( .A(n4643), .B(n4644), .Z(n4289) );
  XOR U3379 ( .A(n4645), .B(n4646), .Z(n4287) );
  XNOR U3380 ( .A(n4647), .B(n4648), .Z(n4646) );
  NOR U3381 ( .A(n4649), .B(n4648), .Z(n4647) );
  XOR U3382 ( .A(n4650), .B(n4651), .Z(n4645) );
  NOR U3383 ( .A(n4652), .B(n4643), .Z(n4651) );
  NOR U3384 ( .A(n4653), .B(n4644), .Z(n4650) );
  XOR U3385 ( .A(n4654), .B(n4655), .Z(n4280) );
  XOR U3386 ( .A(n4656), .B(n4657), .Z(n4278) );
  XNOR U3387 ( .A(n4658), .B(n4659), .Z(n4657) );
  NOR U3388 ( .A(n4660), .B(n4659), .Z(n4658) );
  XOR U3389 ( .A(n4661), .B(n4662), .Z(n4656) );
  NOR U3390 ( .A(n4663), .B(n4654), .Z(n4662) );
  NOR U3391 ( .A(n4664), .B(n4655), .Z(n4661) );
  XOR U3392 ( .A(n4665), .B(n4666), .Z(n4271) );
  XOR U3393 ( .A(n4667), .B(n4668), .Z(n4269) );
  XNOR U3394 ( .A(n4669), .B(n4670), .Z(n4668) );
  NOR U3395 ( .A(n4671), .B(n4670), .Z(n4669) );
  XOR U3396 ( .A(n4672), .B(n4673), .Z(n4667) );
  NOR U3397 ( .A(n4674), .B(n4665), .Z(n4673) );
  NOR U3398 ( .A(n4675), .B(n4666), .Z(n4672) );
  XOR U3399 ( .A(n4676), .B(n4677), .Z(n4262) );
  XOR U3400 ( .A(n4678), .B(n4679), .Z(n4260) );
  XNOR U3401 ( .A(n4680), .B(n4681), .Z(n4679) );
  NOR U3402 ( .A(n4682), .B(n4681), .Z(n4680) );
  XOR U3403 ( .A(n4683), .B(n4684), .Z(n4678) );
  NOR U3404 ( .A(n4685), .B(n4676), .Z(n4684) );
  NOR U3405 ( .A(n4686), .B(n4677), .Z(n4683) );
  XOR U3406 ( .A(n4687), .B(n4688), .Z(n4253) );
  XOR U3407 ( .A(n4689), .B(n4690), .Z(n4251) );
  XNOR U3408 ( .A(n4691), .B(n4692), .Z(n4690) );
  NOR U3409 ( .A(n4693), .B(n4692), .Z(n4691) );
  XOR U3410 ( .A(n4694), .B(n4695), .Z(n4689) );
  NOR U3411 ( .A(n4696), .B(n4687), .Z(n4695) );
  NOR U3412 ( .A(n4697), .B(n4688), .Z(n4694) );
  XOR U3413 ( .A(n4698), .B(n4699), .Z(n4244) );
  XOR U3414 ( .A(n4700), .B(n4701), .Z(n4242) );
  XNOR U3415 ( .A(n4702), .B(n4703), .Z(n4701) );
  NOR U3416 ( .A(n4704), .B(n4703), .Z(n4702) );
  XOR U3417 ( .A(n4705), .B(n4706), .Z(n4700) );
  NOR U3418 ( .A(n4707), .B(n4698), .Z(n4706) );
  NOR U3419 ( .A(n4708), .B(n4699), .Z(n4705) );
  XOR U3420 ( .A(n4709), .B(n4710), .Z(n4235) );
  XOR U3421 ( .A(n4711), .B(n4712), .Z(n4233) );
  XNOR U3422 ( .A(n4713), .B(n4714), .Z(n4712) );
  NOR U3423 ( .A(n4715), .B(n4714), .Z(n4713) );
  XOR U3424 ( .A(n4716), .B(n4717), .Z(n4711) );
  NOR U3425 ( .A(n4718), .B(n4709), .Z(n4717) );
  NOR U3426 ( .A(n4719), .B(n4710), .Z(n4716) );
  XOR U3427 ( .A(n4720), .B(n4721), .Z(n4226) );
  XOR U3428 ( .A(n4722), .B(n4723), .Z(n4224) );
  XNOR U3429 ( .A(n4724), .B(n4725), .Z(n4723) );
  NOR U3430 ( .A(n4726), .B(n4725), .Z(n4724) );
  XOR U3431 ( .A(n4727), .B(n4728), .Z(n4722) );
  NOR U3432 ( .A(n4729), .B(n4720), .Z(n4728) );
  NOR U3433 ( .A(n4730), .B(n4721), .Z(n4727) );
  XOR U3434 ( .A(n4731), .B(n4732), .Z(n4217) );
  XOR U3435 ( .A(n4733), .B(n4734), .Z(n4215) );
  XNOR U3436 ( .A(n4735), .B(n4736), .Z(n4734) );
  NOR U3437 ( .A(n4737), .B(n4736), .Z(n4735) );
  XOR U3438 ( .A(n4738), .B(n4739), .Z(n4733) );
  NOR U3439 ( .A(n4740), .B(n4731), .Z(n4739) );
  NOR U3440 ( .A(n4741), .B(n4732), .Z(n4738) );
  XOR U3441 ( .A(n4742), .B(n4743), .Z(n4208) );
  XOR U3442 ( .A(n4744), .B(n4745), .Z(n4206) );
  XNOR U3443 ( .A(n4746), .B(n4747), .Z(n4745) );
  NOR U3444 ( .A(n4748), .B(n4747), .Z(n4746) );
  XOR U3445 ( .A(n4749), .B(n4750), .Z(n4744) );
  NOR U3446 ( .A(n4751), .B(n4742), .Z(n4750) );
  NOR U3447 ( .A(n4752), .B(n4743), .Z(n4749) );
  XOR U3448 ( .A(n4753), .B(n4754), .Z(n4199) );
  XOR U3449 ( .A(n4755), .B(n4756), .Z(n4197) );
  XNOR U3450 ( .A(n4757), .B(n4758), .Z(n4756) );
  NOR U3451 ( .A(n4759), .B(n4758), .Z(n4757) );
  XOR U3452 ( .A(n4760), .B(n4761), .Z(n4755) );
  NOR U3453 ( .A(n4762), .B(n4753), .Z(n4761) );
  NOR U3454 ( .A(n4763), .B(n4754), .Z(n4760) );
  XOR U3455 ( .A(n4764), .B(n4765), .Z(n4190) );
  XOR U3456 ( .A(n4766), .B(n4767), .Z(n4188) );
  XNOR U3457 ( .A(n4768), .B(n4769), .Z(n4767) );
  NOR U3458 ( .A(n4770), .B(n4769), .Z(n4768) );
  XOR U3459 ( .A(n4771), .B(n4772), .Z(n4766) );
  NOR U3460 ( .A(n4773), .B(n4764), .Z(n4772) );
  NOR U3461 ( .A(n4774), .B(n4765), .Z(n4771) );
  XOR U3462 ( .A(n4775), .B(n4776), .Z(n4181) );
  XOR U3463 ( .A(n4777), .B(n4778), .Z(n4179) );
  XNOR U3464 ( .A(n4779), .B(n4780), .Z(n4778) );
  NOR U3465 ( .A(n4781), .B(n4780), .Z(n4779) );
  XOR U3466 ( .A(n4782), .B(n4783), .Z(n4777) );
  NOR U3467 ( .A(n4784), .B(n4775), .Z(n4783) );
  NOR U3468 ( .A(n4785), .B(n4776), .Z(n4782) );
  XOR U3469 ( .A(n4786), .B(n4787), .Z(n4172) );
  XOR U3470 ( .A(n4788), .B(n4789), .Z(n4170) );
  XNOR U3471 ( .A(n4790), .B(n4791), .Z(n4789) );
  NOR U3472 ( .A(n4792), .B(n4791), .Z(n4790) );
  XOR U3473 ( .A(n4793), .B(n4794), .Z(n4788) );
  NOR U3474 ( .A(n4795), .B(n4786), .Z(n4794) );
  NOR U3475 ( .A(n4796), .B(n4787), .Z(n4793) );
  XOR U3476 ( .A(n4167), .B(n4165), .Z(n4168) );
  XNOR U3477 ( .A(n4797), .B(n4798), .Z(n2041) );
  NOR U3478 ( .A(n4799), .B(n4797), .Z(n4798) );
  XOR U3479 ( .A(n4800), .B(n4801), .Z(n2032) );
  NOR U3480 ( .A(n4802), .B(n4800), .Z(n4801) );
  XOR U3481 ( .A(n4803), .B(n4804), .Z(n2033) );
  NOR U3482 ( .A(n4805), .B(n4803), .Z(n4804) );
  XOR U3483 ( .A(n4806), .B(n4807), .Z(n2030) );
  NOR U3484 ( .A(n4808), .B(n4806), .Z(n4807) );
  XOR U3485 ( .A(n4809), .B(n4810), .Z(n2020) );
  NOR U3486 ( .A(n4811), .B(n4809), .Z(n4810) );
  XOR U3487 ( .A(n4812), .B(n4813), .Z(n2051) );
  NOR U3488 ( .A(n4814), .B(n4812), .Z(n4813) );
  XOR U3489 ( .A(n4815), .B(n4816), .Z(n2048) );
  NOR U3490 ( .A(n4817), .B(n4815), .Z(n4816) );
  XOR U3491 ( .A(n4818), .B(n4819), .Z(n2024) );
  NOR U3492 ( .A(n4820), .B(n4818), .Z(n4819) );
  XOR U3493 ( .A(n4821), .B(n4822), .Z(n2068) );
  NOR U3494 ( .A(n4823), .B(n4821), .Z(n4822) );
  XOR U3495 ( .A(n4824), .B(n4825), .Z(n2063) );
  NOR U3496 ( .A(n4826), .B(n4824), .Z(n4825) );
  XOR U3497 ( .A(n4827), .B(n4828), .Z(n2064) );
  NOR U3498 ( .A(n4829), .B(n4827), .Z(n4828) );
  XOR U3499 ( .A(n4830), .B(n4831), .Z(n2021) );
  NOR U3500 ( .A(n4832), .B(n4830), .Z(n4831) );
  XOR U3501 ( .A(n4833), .B(n4834), .Z(n2079) );
  NOR U3502 ( .A(n4835), .B(n4833), .Z(n4834) );
  XOR U3503 ( .A(n4836), .B(n4837), .Z(n2074) );
  NOR U3504 ( .A(n4838), .B(n4836), .Z(n4837) );
  XOR U3505 ( .A(n4839), .B(n4840), .Z(n2075) );
  NOR U3506 ( .A(n4841), .B(n4839), .Z(n4840) );
  XOR U3507 ( .A(n4842), .B(n4843), .Z(n2014) );
  NOR U3508 ( .A(n4844), .B(n4842), .Z(n4843) );
  XOR U3509 ( .A(n4845), .B(n4846), .Z(n2090) );
  NOR U3510 ( .A(n4847), .B(n4845), .Z(n4846) );
  XOR U3511 ( .A(n4848), .B(n4849), .Z(n2085) );
  NOR U3512 ( .A(n4850), .B(n4848), .Z(n4849) );
  XOR U3513 ( .A(n4851), .B(n4852), .Z(n2086) );
  NOR U3514 ( .A(n4853), .B(n4851), .Z(n4852) );
  XOR U3515 ( .A(n4854), .B(n4855), .Z(n2005) );
  NOR U3516 ( .A(n4856), .B(n4854), .Z(n4855) );
  XOR U3517 ( .A(n4857), .B(n4858), .Z(n2101) );
  NOR U3518 ( .A(n4859), .B(n4857), .Z(n4858) );
  XOR U3519 ( .A(n4860), .B(n4861), .Z(n2096) );
  NOR U3520 ( .A(n4862), .B(n4860), .Z(n4861) );
  XOR U3521 ( .A(n4863), .B(n4864), .Z(n2097) );
  NOR U3522 ( .A(n4865), .B(n4863), .Z(n4864) );
  XOR U3523 ( .A(n4866), .B(n4867), .Z(n1996) );
  NOR U3524 ( .A(n4868), .B(n4866), .Z(n4867) );
  XOR U3525 ( .A(n4869), .B(n4870), .Z(n2112) );
  NOR U3526 ( .A(n4871), .B(n4869), .Z(n4870) );
  XOR U3527 ( .A(n4872), .B(n4873), .Z(n2107) );
  NOR U3528 ( .A(n4874), .B(n4872), .Z(n4873) );
  XOR U3529 ( .A(n4875), .B(n4876), .Z(n2108) );
  NOR U3530 ( .A(n4877), .B(n4875), .Z(n4876) );
  XOR U3531 ( .A(n4878), .B(n4879), .Z(n1987) );
  NOR U3532 ( .A(n4880), .B(n4878), .Z(n4879) );
  XOR U3533 ( .A(n4881), .B(n4882), .Z(n2123) );
  NOR U3534 ( .A(n4883), .B(n4881), .Z(n4882) );
  XOR U3535 ( .A(n4884), .B(n4885), .Z(n2118) );
  NOR U3536 ( .A(n4886), .B(n4884), .Z(n4885) );
  XOR U3537 ( .A(n4887), .B(n4888), .Z(n2119) );
  NOR U3538 ( .A(n4889), .B(n4887), .Z(n4888) );
  XOR U3539 ( .A(n4890), .B(n4891), .Z(n1978) );
  NOR U3540 ( .A(n4892), .B(n4890), .Z(n4891) );
  XOR U3541 ( .A(n4893), .B(n4894), .Z(n2134) );
  NOR U3542 ( .A(n4895), .B(n4893), .Z(n4894) );
  XOR U3543 ( .A(n4896), .B(n4897), .Z(n2129) );
  NOR U3544 ( .A(n4898), .B(n4896), .Z(n4897) );
  XOR U3545 ( .A(n4899), .B(n4900), .Z(n2130) );
  NOR U3546 ( .A(n4901), .B(n4899), .Z(n4900) );
  XOR U3547 ( .A(n4902), .B(n4903), .Z(n1969) );
  NOR U3548 ( .A(n4904), .B(n4902), .Z(n4903) );
  XOR U3549 ( .A(n4905), .B(n4906), .Z(n2145) );
  NOR U3550 ( .A(n4907), .B(n4905), .Z(n4906) );
  XOR U3551 ( .A(n4908), .B(n4909), .Z(n2140) );
  NOR U3552 ( .A(n4910), .B(n4908), .Z(n4909) );
  XOR U3553 ( .A(n4911), .B(n4912), .Z(n2141) );
  NOR U3554 ( .A(n4913), .B(n4911), .Z(n4912) );
  XOR U3555 ( .A(n4914), .B(n4915), .Z(n1960) );
  NOR U3556 ( .A(n4916), .B(n4914), .Z(n4915) );
  XOR U3557 ( .A(n4917), .B(n4918), .Z(n2156) );
  NOR U3558 ( .A(n4919), .B(n4917), .Z(n4918) );
  XOR U3559 ( .A(n4920), .B(n4921), .Z(n2151) );
  NOR U3560 ( .A(n4922), .B(n4920), .Z(n4921) );
  XOR U3561 ( .A(n4923), .B(n4924), .Z(n2152) );
  NOR U3562 ( .A(n4925), .B(n4923), .Z(n4924) );
  XOR U3563 ( .A(n4926), .B(n4927), .Z(n1951) );
  NOR U3564 ( .A(n4928), .B(n4926), .Z(n4927) );
  XOR U3565 ( .A(n4929), .B(n4930), .Z(n2167) );
  NOR U3566 ( .A(n4931), .B(n4929), .Z(n4930) );
  XOR U3567 ( .A(n4932), .B(n4933), .Z(n2162) );
  NOR U3568 ( .A(n4934), .B(n4932), .Z(n4933) );
  XOR U3569 ( .A(n4935), .B(n4936), .Z(n2163) );
  NOR U3570 ( .A(n4937), .B(n4935), .Z(n4936) );
  XOR U3571 ( .A(n4938), .B(n4939), .Z(n1942) );
  NOR U3572 ( .A(n4940), .B(n4938), .Z(n4939) );
  XOR U3573 ( .A(n4941), .B(n4942), .Z(n2178) );
  NOR U3574 ( .A(n4943), .B(n4941), .Z(n4942) );
  XOR U3575 ( .A(n4944), .B(n4945), .Z(n2173) );
  NOR U3576 ( .A(n4946), .B(n4944), .Z(n4945) );
  XOR U3577 ( .A(n4947), .B(n4948), .Z(n2174) );
  NOR U3578 ( .A(n4949), .B(n4947), .Z(n4948) );
  XOR U3579 ( .A(n4950), .B(n4951), .Z(n1933) );
  NOR U3580 ( .A(n4952), .B(n4950), .Z(n4951) );
  XOR U3581 ( .A(n4953), .B(n4954), .Z(n2189) );
  NOR U3582 ( .A(n4955), .B(n4953), .Z(n4954) );
  XOR U3583 ( .A(n4956), .B(n4957), .Z(n2184) );
  NOR U3584 ( .A(n4958), .B(n4956), .Z(n4957) );
  XOR U3585 ( .A(n4959), .B(n4960), .Z(n2185) );
  NOR U3586 ( .A(n4961), .B(n4959), .Z(n4960) );
  XOR U3587 ( .A(n4962), .B(n4963), .Z(n1924) );
  NOR U3588 ( .A(n4964), .B(n4962), .Z(n4963) );
  XOR U3589 ( .A(n4965), .B(n4966), .Z(n2200) );
  NOR U3590 ( .A(n4967), .B(n4965), .Z(n4966) );
  XOR U3591 ( .A(n4968), .B(n4969), .Z(n2195) );
  NOR U3592 ( .A(n4970), .B(n4968), .Z(n4969) );
  XOR U3593 ( .A(n4971), .B(n4972), .Z(n2196) );
  NOR U3594 ( .A(n4973), .B(n4971), .Z(n4972) );
  XOR U3595 ( .A(n4974), .B(n4975), .Z(n1915) );
  NOR U3596 ( .A(n4976), .B(n4974), .Z(n4975) );
  XOR U3597 ( .A(n4977), .B(n4978), .Z(n2211) );
  NOR U3598 ( .A(n4979), .B(n4977), .Z(n4978) );
  XOR U3599 ( .A(n4980), .B(n4981), .Z(n2206) );
  NOR U3600 ( .A(n4982), .B(n4980), .Z(n4981) );
  XOR U3601 ( .A(n4983), .B(n4984), .Z(n2207) );
  NOR U3602 ( .A(n4985), .B(n4983), .Z(n4984) );
  XOR U3603 ( .A(n4986), .B(n4987), .Z(n1906) );
  NOR U3604 ( .A(n4988), .B(n4986), .Z(n4987) );
  XOR U3605 ( .A(n4989), .B(n4990), .Z(n2222) );
  NOR U3606 ( .A(n4991), .B(n4989), .Z(n4990) );
  XOR U3607 ( .A(n4992), .B(n4993), .Z(n2217) );
  NOR U3608 ( .A(n4994), .B(n4992), .Z(n4993) );
  XOR U3609 ( .A(n4995), .B(n4996), .Z(n2218) );
  NOR U3610 ( .A(n4997), .B(n4995), .Z(n4996) );
  XOR U3611 ( .A(n4998), .B(n4999), .Z(n1897) );
  NOR U3612 ( .A(n5000), .B(n4998), .Z(n4999) );
  XOR U3613 ( .A(n5001), .B(n5002), .Z(n2233) );
  NOR U3614 ( .A(n5003), .B(n5001), .Z(n5002) );
  XOR U3615 ( .A(n5004), .B(n5005), .Z(n2228) );
  NOR U3616 ( .A(n5006), .B(n5004), .Z(n5005) );
  XOR U3617 ( .A(n5007), .B(n5008), .Z(n2229) );
  NOR U3618 ( .A(n5009), .B(n5007), .Z(n5008) );
  XOR U3619 ( .A(n5010), .B(n5011), .Z(n1888) );
  NOR U3620 ( .A(n5012), .B(n5010), .Z(n5011) );
  XOR U3621 ( .A(n5013), .B(n5014), .Z(n2244) );
  NOR U3622 ( .A(n5015), .B(n5013), .Z(n5014) );
  XOR U3623 ( .A(n5016), .B(n5017), .Z(n2239) );
  NOR U3624 ( .A(n5018), .B(n5016), .Z(n5017) );
  XOR U3625 ( .A(n5019), .B(n5020), .Z(n2240) );
  NOR U3626 ( .A(n5021), .B(n5019), .Z(n5020) );
  XOR U3627 ( .A(n5022), .B(n5023), .Z(n1879) );
  NOR U3628 ( .A(n5024), .B(n5022), .Z(n5023) );
  XOR U3629 ( .A(n5025), .B(n5026), .Z(n2255) );
  NOR U3630 ( .A(n5027), .B(n5025), .Z(n5026) );
  XOR U3631 ( .A(n5028), .B(n5029), .Z(n2250) );
  NOR U3632 ( .A(n5030), .B(n5028), .Z(n5029) );
  XOR U3633 ( .A(n5031), .B(n5032), .Z(n2251) );
  NOR U3634 ( .A(n5033), .B(n5031), .Z(n5032) );
  XOR U3635 ( .A(n5034), .B(n5035), .Z(n1870) );
  NOR U3636 ( .A(n5036), .B(n5034), .Z(n5035) );
  XOR U3637 ( .A(n5037), .B(n5038), .Z(n2266) );
  NOR U3638 ( .A(n5039), .B(n5037), .Z(n5038) );
  XOR U3639 ( .A(n5040), .B(n5041), .Z(n2261) );
  NOR U3640 ( .A(n5042), .B(n5040), .Z(n5041) );
  XOR U3641 ( .A(n5043), .B(n5044), .Z(n2262) );
  NOR U3642 ( .A(n5045), .B(n5043), .Z(n5044) );
  XOR U3643 ( .A(n5046), .B(n5047), .Z(n1861) );
  NOR U3644 ( .A(n5048), .B(n5046), .Z(n5047) );
  XOR U3645 ( .A(n5049), .B(n5050), .Z(n2277) );
  NOR U3646 ( .A(n5051), .B(n5049), .Z(n5050) );
  XOR U3647 ( .A(n5052), .B(n5053), .Z(n2272) );
  NOR U3648 ( .A(n5054), .B(n5052), .Z(n5053) );
  XOR U3649 ( .A(n5055), .B(n5056), .Z(n2273) );
  NOR U3650 ( .A(n5057), .B(n5055), .Z(n5056) );
  XOR U3651 ( .A(n5058), .B(n5059), .Z(n1852) );
  NOR U3652 ( .A(n5060), .B(n5058), .Z(n5059) );
  XOR U3653 ( .A(n5061), .B(n5062), .Z(n2288) );
  NOR U3654 ( .A(n5063), .B(n5061), .Z(n5062) );
  XOR U3655 ( .A(n5064), .B(n5065), .Z(n2283) );
  NOR U3656 ( .A(n5066), .B(n5064), .Z(n5065) );
  XOR U3657 ( .A(n5067), .B(n5068), .Z(n2284) );
  NOR U3658 ( .A(n5069), .B(n5067), .Z(n5068) );
  XOR U3659 ( .A(n5070), .B(n5071), .Z(n1843) );
  NOR U3660 ( .A(n5072), .B(n5070), .Z(n5071) );
  XOR U3661 ( .A(n5073), .B(n5074), .Z(n2299) );
  NOR U3662 ( .A(n5075), .B(n5073), .Z(n5074) );
  XOR U3663 ( .A(n5076), .B(n5077), .Z(n2294) );
  NOR U3664 ( .A(n5078), .B(n5076), .Z(n5077) );
  XOR U3665 ( .A(n5079), .B(n5080), .Z(n2295) );
  NOR U3666 ( .A(n5081), .B(n5079), .Z(n5080) );
  XOR U3667 ( .A(n5082), .B(n5083), .Z(n1834) );
  NOR U3668 ( .A(n5084), .B(n5082), .Z(n5083) );
  XOR U3669 ( .A(n5085), .B(n5086), .Z(n2310) );
  NOR U3670 ( .A(n5087), .B(n5085), .Z(n5086) );
  XOR U3671 ( .A(n5088), .B(n5089), .Z(n2305) );
  NOR U3672 ( .A(n5090), .B(n5088), .Z(n5089) );
  XOR U3673 ( .A(n5091), .B(n5092), .Z(n2306) );
  NOR U3674 ( .A(n5093), .B(n5091), .Z(n5092) );
  XOR U3675 ( .A(n5094), .B(n5095), .Z(n1825) );
  NOR U3676 ( .A(n5096), .B(n5094), .Z(n5095) );
  XOR U3677 ( .A(n5097), .B(n5098), .Z(n2321) );
  NOR U3678 ( .A(n5099), .B(n5097), .Z(n5098) );
  XOR U3679 ( .A(n5100), .B(n5101), .Z(n2316) );
  NOR U3680 ( .A(n5102), .B(n5100), .Z(n5101) );
  XOR U3681 ( .A(n5103), .B(n5104), .Z(n2317) );
  NOR U3682 ( .A(n5105), .B(n5103), .Z(n5104) );
  XOR U3683 ( .A(n5106), .B(n5107), .Z(n1816) );
  NOR U3684 ( .A(n5108), .B(n5106), .Z(n5107) );
  XOR U3685 ( .A(n5109), .B(n5110), .Z(n2332) );
  NOR U3686 ( .A(n5111), .B(n5109), .Z(n5110) );
  XOR U3687 ( .A(n5112), .B(n5113), .Z(n2327) );
  NOR U3688 ( .A(n5114), .B(n5112), .Z(n5113) );
  XOR U3689 ( .A(n5115), .B(n5116), .Z(n2328) );
  NOR U3690 ( .A(n5117), .B(n5115), .Z(n5116) );
  XOR U3691 ( .A(n5118), .B(n5119), .Z(n1807) );
  NOR U3692 ( .A(n5120), .B(n5118), .Z(n5119) );
  XOR U3693 ( .A(n5121), .B(n5122), .Z(n2343) );
  NOR U3694 ( .A(n5123), .B(n5121), .Z(n5122) );
  XOR U3695 ( .A(n5124), .B(n5125), .Z(n2338) );
  NOR U3696 ( .A(n5126), .B(n5124), .Z(n5125) );
  XOR U3697 ( .A(n5127), .B(n5128), .Z(n2339) );
  NOR U3698 ( .A(n5129), .B(n5127), .Z(n5128) );
  XOR U3699 ( .A(n5130), .B(n5131), .Z(n1798) );
  NOR U3700 ( .A(n5132), .B(n5130), .Z(n5131) );
  XOR U3701 ( .A(n5133), .B(n5134), .Z(n2354) );
  NOR U3702 ( .A(n5135), .B(n5133), .Z(n5134) );
  XOR U3703 ( .A(n5136), .B(n5137), .Z(n2349) );
  NOR U3704 ( .A(n5138), .B(n5136), .Z(n5137) );
  XOR U3705 ( .A(n5139), .B(n5140), .Z(n2350) );
  NOR U3706 ( .A(n5141), .B(n5139), .Z(n5140) );
  XOR U3707 ( .A(n5142), .B(n5143), .Z(n1789) );
  NOR U3708 ( .A(n5144), .B(n5142), .Z(n5143) );
  XOR U3709 ( .A(n5145), .B(n5146), .Z(n2365) );
  NOR U3710 ( .A(n5147), .B(n5145), .Z(n5146) );
  XOR U3711 ( .A(n5148), .B(n5149), .Z(n2360) );
  NOR U3712 ( .A(n5150), .B(n5148), .Z(n5149) );
  XOR U3713 ( .A(n5151), .B(n5152), .Z(n2361) );
  NOR U3714 ( .A(n5153), .B(n5151), .Z(n5152) );
  XOR U3715 ( .A(n5154), .B(n5155), .Z(n1780) );
  NOR U3716 ( .A(n5156), .B(n5154), .Z(n5155) );
  XOR U3717 ( .A(n5157), .B(n5158), .Z(n2376) );
  NOR U3718 ( .A(n5159), .B(n5157), .Z(n5158) );
  XOR U3719 ( .A(n5160), .B(n5161), .Z(n2371) );
  NOR U3720 ( .A(n5162), .B(n5160), .Z(n5161) );
  XOR U3721 ( .A(n5163), .B(n5164), .Z(n2372) );
  NOR U3722 ( .A(n5165), .B(n5163), .Z(n5164) );
  XOR U3723 ( .A(n5166), .B(n5167), .Z(n1771) );
  NOR U3724 ( .A(n5168), .B(n5166), .Z(n5167) );
  XOR U3725 ( .A(n5169), .B(n5170), .Z(n2387) );
  NOR U3726 ( .A(n5171), .B(n5169), .Z(n5170) );
  XOR U3727 ( .A(n5172), .B(n5173), .Z(n2382) );
  NOR U3728 ( .A(n5174), .B(n5172), .Z(n5173) );
  XOR U3729 ( .A(n5175), .B(n5176), .Z(n2383) );
  NOR U3730 ( .A(n5177), .B(n5175), .Z(n5176) );
  XOR U3731 ( .A(n5178), .B(n5179), .Z(n1762) );
  NOR U3732 ( .A(n5180), .B(n5178), .Z(n5179) );
  XOR U3733 ( .A(n5181), .B(n5182), .Z(n2398) );
  NOR U3734 ( .A(n5183), .B(n5181), .Z(n5182) );
  XOR U3735 ( .A(n5184), .B(n5185), .Z(n2393) );
  NOR U3736 ( .A(n5186), .B(n5184), .Z(n5185) );
  XOR U3737 ( .A(n5187), .B(n5188), .Z(n2394) );
  NOR U3738 ( .A(n5189), .B(n5187), .Z(n5188) );
  XOR U3739 ( .A(n5190), .B(n5191), .Z(n1753) );
  NOR U3740 ( .A(n5192), .B(n5190), .Z(n5191) );
  XOR U3741 ( .A(n5193), .B(n5194), .Z(n2409) );
  NOR U3742 ( .A(n5195), .B(n5193), .Z(n5194) );
  XOR U3743 ( .A(n5196), .B(n5197), .Z(n2404) );
  NOR U3744 ( .A(n5198), .B(n5196), .Z(n5197) );
  XOR U3745 ( .A(n5199), .B(n5200), .Z(n2405) );
  NOR U3746 ( .A(n5201), .B(n5199), .Z(n5200) );
  XOR U3747 ( .A(n5202), .B(n5203), .Z(n1744) );
  NOR U3748 ( .A(n5204), .B(n5202), .Z(n5203) );
  XOR U3749 ( .A(n5205), .B(n5206), .Z(n2420) );
  NOR U3750 ( .A(n5207), .B(n5205), .Z(n5206) );
  XOR U3751 ( .A(n5208), .B(n5209), .Z(n2415) );
  NOR U3752 ( .A(n5210), .B(n5208), .Z(n5209) );
  XOR U3753 ( .A(n5211), .B(n5212), .Z(n2416) );
  NOR U3754 ( .A(n5213), .B(n5211), .Z(n5212) );
  XOR U3755 ( .A(n5214), .B(n5215), .Z(n1735) );
  NOR U3756 ( .A(n5216), .B(n5214), .Z(n5215) );
  XOR U3757 ( .A(n5217), .B(n5218), .Z(n2431) );
  NOR U3758 ( .A(n5219), .B(n5217), .Z(n5218) );
  XOR U3759 ( .A(n5220), .B(n5221), .Z(n2426) );
  NOR U3760 ( .A(n5222), .B(n5220), .Z(n5221) );
  XOR U3761 ( .A(n5223), .B(n5224), .Z(n2427) );
  NOR U3762 ( .A(n5225), .B(n5223), .Z(n5224) );
  XOR U3763 ( .A(n5226), .B(n5227), .Z(n1726) );
  NOR U3764 ( .A(n5228), .B(n5226), .Z(n5227) );
  XOR U3765 ( .A(n5229), .B(n5230), .Z(n2442) );
  NOR U3766 ( .A(n5231), .B(n5229), .Z(n5230) );
  XOR U3767 ( .A(n5232), .B(n5233), .Z(n2437) );
  NOR U3768 ( .A(n5234), .B(n5232), .Z(n5233) );
  XOR U3769 ( .A(n5235), .B(n5236), .Z(n2438) );
  NOR U3770 ( .A(n5237), .B(n5235), .Z(n5236) );
  XOR U3771 ( .A(n5238), .B(n5239), .Z(n1717) );
  NOR U3772 ( .A(n5240), .B(n5238), .Z(n5239) );
  XOR U3773 ( .A(n5241), .B(n5242), .Z(n2453) );
  NOR U3774 ( .A(n5243), .B(n5241), .Z(n5242) );
  XOR U3775 ( .A(n5244), .B(n5245), .Z(n2448) );
  NOR U3776 ( .A(n5246), .B(n5244), .Z(n5245) );
  XOR U3777 ( .A(n5247), .B(n5248), .Z(n2449) );
  NOR U3778 ( .A(n5249), .B(n5247), .Z(n5248) );
  XOR U3779 ( .A(n5250), .B(n5251), .Z(n1708) );
  NOR U3780 ( .A(n5252), .B(n5250), .Z(n5251) );
  XOR U3781 ( .A(n5253), .B(n5254), .Z(n2464) );
  NOR U3782 ( .A(n5255), .B(n5253), .Z(n5254) );
  XOR U3783 ( .A(n5256), .B(n5257), .Z(n2459) );
  NOR U3784 ( .A(n5258), .B(n5256), .Z(n5257) );
  XOR U3785 ( .A(n5259), .B(n5260), .Z(n2460) );
  NOR U3786 ( .A(n5261), .B(n5259), .Z(n5260) );
  XOR U3787 ( .A(n5262), .B(n5263), .Z(n1699) );
  NOR U3788 ( .A(n5264), .B(n5262), .Z(n5263) );
  XOR U3789 ( .A(n5265), .B(n5266), .Z(n2475) );
  NOR U3790 ( .A(n5267), .B(n5265), .Z(n5266) );
  XOR U3791 ( .A(n5268), .B(n5269), .Z(n2470) );
  NOR U3792 ( .A(n5270), .B(n5268), .Z(n5269) );
  XOR U3793 ( .A(n5271), .B(n5272), .Z(n2471) );
  NOR U3794 ( .A(n5273), .B(n5271), .Z(n5272) );
  XOR U3795 ( .A(n5274), .B(n5275), .Z(n1690) );
  NOR U3796 ( .A(n5276), .B(n5274), .Z(n5275) );
  XOR U3797 ( .A(n5277), .B(n5278), .Z(n2486) );
  NOR U3798 ( .A(n5279), .B(n5277), .Z(n5278) );
  XOR U3799 ( .A(n5280), .B(n5281), .Z(n2481) );
  NOR U3800 ( .A(n5282), .B(n5280), .Z(n5281) );
  XOR U3801 ( .A(n5283), .B(n5284), .Z(n2482) );
  NOR U3802 ( .A(n5285), .B(n5283), .Z(n5284) );
  XOR U3803 ( .A(n5286), .B(n5287), .Z(n1681) );
  NOR U3804 ( .A(n5288), .B(n5286), .Z(n5287) );
  XOR U3805 ( .A(n5289), .B(n5290), .Z(n2497) );
  NOR U3806 ( .A(n5291), .B(n5289), .Z(n5290) );
  XOR U3807 ( .A(n5292), .B(n5293), .Z(n2492) );
  NOR U3808 ( .A(n5294), .B(n5292), .Z(n5293) );
  XOR U3809 ( .A(n5295), .B(n5296), .Z(n2493) );
  NOR U3810 ( .A(n5297), .B(n5295), .Z(n5296) );
  XOR U3811 ( .A(n5298), .B(n5299), .Z(n1672) );
  NOR U3812 ( .A(n5300), .B(n5298), .Z(n5299) );
  XOR U3813 ( .A(n5301), .B(n5302), .Z(n2508) );
  NOR U3814 ( .A(n5303), .B(n5301), .Z(n5302) );
  XOR U3815 ( .A(n5304), .B(n5305), .Z(n2503) );
  NOR U3816 ( .A(n5306), .B(n5304), .Z(n5305) );
  XOR U3817 ( .A(n5307), .B(n5308), .Z(n2504) );
  NOR U3818 ( .A(n5309), .B(n5307), .Z(n5308) );
  XOR U3819 ( .A(n5310), .B(n5311), .Z(n1663) );
  NOR U3820 ( .A(n5312), .B(n5310), .Z(n5311) );
  XOR U3821 ( .A(n5313), .B(n5314), .Z(n2519) );
  NOR U3822 ( .A(n5315), .B(n5313), .Z(n5314) );
  XOR U3823 ( .A(n5316), .B(n5317), .Z(n2514) );
  NOR U3824 ( .A(n5318), .B(n5316), .Z(n5317) );
  XOR U3825 ( .A(n5319), .B(n5320), .Z(n2515) );
  NOR U3826 ( .A(n5321), .B(n5319), .Z(n5320) );
  XOR U3827 ( .A(n5322), .B(n5323), .Z(n1654) );
  NOR U3828 ( .A(n5324), .B(n5322), .Z(n5323) );
  XOR U3829 ( .A(n5325), .B(n5326), .Z(n2530) );
  NOR U3830 ( .A(n5327), .B(n5325), .Z(n5326) );
  XOR U3831 ( .A(n5328), .B(n5329), .Z(n2525) );
  NOR U3832 ( .A(n5330), .B(n5328), .Z(n5329) );
  XOR U3833 ( .A(n5331), .B(n5332), .Z(n2526) );
  NOR U3834 ( .A(n5333), .B(n5331), .Z(n5332) );
  XOR U3835 ( .A(n5334), .B(n5335), .Z(n1645) );
  NOR U3836 ( .A(n5336), .B(n5334), .Z(n5335) );
  XOR U3837 ( .A(n5337), .B(n5338), .Z(n2541) );
  NOR U3838 ( .A(n5339), .B(n5337), .Z(n5338) );
  XOR U3839 ( .A(n5340), .B(n5341), .Z(n2536) );
  NOR U3840 ( .A(n5342), .B(n5340), .Z(n5341) );
  XOR U3841 ( .A(n5343), .B(n5344), .Z(n2537) );
  NOR U3842 ( .A(n5345), .B(n5343), .Z(n5344) );
  XOR U3843 ( .A(n5346), .B(n5347), .Z(n1636) );
  NOR U3844 ( .A(n5348), .B(n5346), .Z(n5347) );
  XOR U3845 ( .A(n5349), .B(n5350), .Z(n2552) );
  NOR U3846 ( .A(n5351), .B(n5349), .Z(n5350) );
  XOR U3847 ( .A(n5352), .B(n5353), .Z(n2547) );
  NOR U3848 ( .A(n5354), .B(n5352), .Z(n5353) );
  XOR U3849 ( .A(n5355), .B(n5356), .Z(n2548) );
  NOR U3850 ( .A(n5357), .B(n5355), .Z(n5356) );
  XOR U3851 ( .A(n5358), .B(n5359), .Z(n1627) );
  NOR U3852 ( .A(n5360), .B(n5358), .Z(n5359) );
  XOR U3853 ( .A(n5361), .B(n5362), .Z(n2563) );
  NOR U3854 ( .A(n5363), .B(n5361), .Z(n5362) );
  XOR U3855 ( .A(n5364), .B(n5365), .Z(n2558) );
  NOR U3856 ( .A(n5366), .B(n5364), .Z(n5365) );
  XOR U3857 ( .A(n5367), .B(n5368), .Z(n2559) );
  NOR U3858 ( .A(n5369), .B(n5367), .Z(n5368) );
  XOR U3859 ( .A(n5370), .B(n5371), .Z(n1618) );
  NOR U3860 ( .A(n5372), .B(n5370), .Z(n5371) );
  XOR U3861 ( .A(n5373), .B(n5374), .Z(n2574) );
  NOR U3862 ( .A(n5375), .B(n5373), .Z(n5374) );
  XOR U3863 ( .A(n5376), .B(n5377), .Z(n2569) );
  NOR U3864 ( .A(n5378), .B(n5376), .Z(n5377) );
  XOR U3865 ( .A(n5379), .B(n5380), .Z(n2570) );
  NOR U3866 ( .A(n5381), .B(n5379), .Z(n5380) );
  XOR U3867 ( .A(n5382), .B(n5383), .Z(n1609) );
  NOR U3868 ( .A(n5384), .B(n5382), .Z(n5383) );
  XOR U3869 ( .A(n5385), .B(n5386), .Z(n2585) );
  NOR U3870 ( .A(n5387), .B(n5385), .Z(n5386) );
  XOR U3871 ( .A(n5388), .B(n5389), .Z(n2580) );
  NOR U3872 ( .A(n5390), .B(n5388), .Z(n5389) );
  XOR U3873 ( .A(n5391), .B(n5392), .Z(n2581) );
  NOR U3874 ( .A(n5393), .B(n5391), .Z(n5392) );
  XOR U3875 ( .A(n5394), .B(n5395), .Z(n1600) );
  NOR U3876 ( .A(n5396), .B(n5394), .Z(n5395) );
  XOR U3877 ( .A(n5397), .B(n5398), .Z(n2596) );
  NOR U3878 ( .A(n5399), .B(n5397), .Z(n5398) );
  XOR U3879 ( .A(n5400), .B(n5401), .Z(n2591) );
  NOR U3880 ( .A(n5402), .B(n5400), .Z(n5401) );
  XOR U3881 ( .A(n5403), .B(n5404), .Z(n2592) );
  NOR U3882 ( .A(n5405), .B(n5403), .Z(n5404) );
  XOR U3883 ( .A(n5406), .B(n5407), .Z(n1591) );
  NOR U3884 ( .A(n5408), .B(n5406), .Z(n5407) );
  XOR U3885 ( .A(n5409), .B(n5410), .Z(n2607) );
  NOR U3886 ( .A(n5411), .B(n5409), .Z(n5410) );
  XOR U3887 ( .A(n5412), .B(n5413), .Z(n2602) );
  NOR U3888 ( .A(n5414), .B(n5412), .Z(n5413) );
  XOR U3889 ( .A(n5415), .B(n5416), .Z(n2603) );
  NOR U3890 ( .A(n5417), .B(n5415), .Z(n5416) );
  XOR U3891 ( .A(n5418), .B(n5419), .Z(n1582) );
  NOR U3892 ( .A(n5420), .B(n5418), .Z(n5419) );
  XOR U3893 ( .A(n5421), .B(n5422), .Z(n2618) );
  NOR U3894 ( .A(n5423), .B(n5421), .Z(n5422) );
  XOR U3895 ( .A(n5424), .B(n5425), .Z(n2613) );
  NOR U3896 ( .A(n5426), .B(n5424), .Z(n5425) );
  XOR U3897 ( .A(n5427), .B(n5428), .Z(n2614) );
  NOR U3898 ( .A(n5429), .B(n5427), .Z(n5428) );
  XOR U3899 ( .A(n5430), .B(n5431), .Z(n1573) );
  NOR U3900 ( .A(n5432), .B(n5430), .Z(n5431) );
  XOR U3901 ( .A(n5433), .B(n5434), .Z(n2629) );
  NOR U3902 ( .A(n5435), .B(n5433), .Z(n5434) );
  XOR U3903 ( .A(n5436), .B(n5437), .Z(n2624) );
  NOR U3904 ( .A(n5438), .B(n5436), .Z(n5437) );
  XOR U3905 ( .A(n5439), .B(n5440), .Z(n2625) );
  NOR U3906 ( .A(n5441), .B(n5439), .Z(n5440) );
  XOR U3907 ( .A(n5442), .B(n5443), .Z(n1564) );
  NOR U3908 ( .A(n5444), .B(n5442), .Z(n5443) );
  XOR U3909 ( .A(n5445), .B(n5446), .Z(n2640) );
  NOR U3910 ( .A(n5447), .B(n5445), .Z(n5446) );
  XOR U3911 ( .A(n5448), .B(n5449), .Z(n2635) );
  NOR U3912 ( .A(n5450), .B(n5448), .Z(n5449) );
  XOR U3913 ( .A(n5451), .B(n5452), .Z(n2636) );
  NOR U3914 ( .A(n5453), .B(n5451), .Z(n5452) );
  XOR U3915 ( .A(n5454), .B(n5455), .Z(n1555) );
  NOR U3916 ( .A(n5456), .B(n5454), .Z(n5455) );
  XOR U3917 ( .A(n5457), .B(n5458), .Z(n2651) );
  NOR U3918 ( .A(n5459), .B(n5457), .Z(n5458) );
  XOR U3919 ( .A(n5460), .B(n5461), .Z(n2646) );
  NOR U3920 ( .A(n5462), .B(n5460), .Z(n5461) );
  XOR U3921 ( .A(n5463), .B(n5464), .Z(n2647) );
  NOR U3922 ( .A(n5465), .B(n5463), .Z(n5464) );
  XOR U3923 ( .A(n5466), .B(n5467), .Z(n1546) );
  NOR U3924 ( .A(n5468), .B(n5466), .Z(n5467) );
  XOR U3925 ( .A(n5469), .B(n5470), .Z(n2662) );
  NOR U3926 ( .A(n5471), .B(n5469), .Z(n5470) );
  XOR U3927 ( .A(n5472), .B(n5473), .Z(n2657) );
  NOR U3928 ( .A(n5474), .B(n5472), .Z(n5473) );
  XOR U3929 ( .A(n5475), .B(n5476), .Z(n2658) );
  NOR U3930 ( .A(n5477), .B(n5475), .Z(n5476) );
  XOR U3931 ( .A(n5478), .B(n5479), .Z(n1537) );
  NOR U3932 ( .A(n5480), .B(n5478), .Z(n5479) );
  XOR U3933 ( .A(n5481), .B(n5482), .Z(n2673) );
  NOR U3934 ( .A(n5483), .B(n5481), .Z(n5482) );
  XOR U3935 ( .A(n5484), .B(n5485), .Z(n2668) );
  NOR U3936 ( .A(n5486), .B(n5484), .Z(n5485) );
  XOR U3937 ( .A(n5487), .B(n5488), .Z(n2669) );
  NOR U3938 ( .A(n5489), .B(n5487), .Z(n5488) );
  XOR U3939 ( .A(n5490), .B(n5491), .Z(n1528) );
  NOR U3940 ( .A(n5492), .B(n5490), .Z(n5491) );
  XOR U3941 ( .A(n5493), .B(n5494), .Z(n2684) );
  NOR U3942 ( .A(n5495), .B(n5493), .Z(n5494) );
  XOR U3943 ( .A(n5496), .B(n5497), .Z(n2679) );
  NOR U3944 ( .A(n5498), .B(n5496), .Z(n5497) );
  XOR U3945 ( .A(n5499), .B(n5500), .Z(n2680) );
  NOR U3946 ( .A(n5501), .B(n5499), .Z(n5500) );
  XOR U3947 ( .A(n5502), .B(n5503), .Z(n1519) );
  NOR U3948 ( .A(n5504), .B(n5502), .Z(n5503) );
  XOR U3949 ( .A(n5505), .B(n5506), .Z(n2695) );
  NOR U3950 ( .A(n5507), .B(n5505), .Z(n5506) );
  XOR U3951 ( .A(n5508), .B(n5509), .Z(n2690) );
  NOR U3952 ( .A(n5510), .B(n5508), .Z(n5509) );
  XOR U3953 ( .A(n5511), .B(n5512), .Z(n2691) );
  NOR U3954 ( .A(n5513), .B(n5511), .Z(n5512) );
  XOR U3955 ( .A(n5514), .B(n5515), .Z(n1510) );
  NOR U3956 ( .A(n5516), .B(n5514), .Z(n5515) );
  XOR U3957 ( .A(n5517), .B(n5518), .Z(n2706) );
  NOR U3958 ( .A(n5519), .B(n5517), .Z(n5518) );
  XOR U3959 ( .A(n5520), .B(n5521), .Z(n2701) );
  NOR U3960 ( .A(n5522), .B(n5520), .Z(n5521) );
  XOR U3961 ( .A(n5523), .B(n5524), .Z(n2702) );
  NOR U3962 ( .A(n5525), .B(n5523), .Z(n5524) );
  XOR U3963 ( .A(n5526), .B(n5527), .Z(n1501) );
  NOR U3964 ( .A(n5528), .B(n5526), .Z(n5527) );
  XOR U3965 ( .A(n5529), .B(n5530), .Z(n2717) );
  NOR U3966 ( .A(n5531), .B(n5529), .Z(n5530) );
  XOR U3967 ( .A(n5532), .B(n5533), .Z(n2712) );
  NOR U3968 ( .A(n5534), .B(n5532), .Z(n5533) );
  XOR U3969 ( .A(n5535), .B(n5536), .Z(n2713) );
  NOR U3970 ( .A(n5537), .B(n5535), .Z(n5536) );
  XOR U3971 ( .A(n5538), .B(n5539), .Z(n1492) );
  NOR U3972 ( .A(n5540), .B(n5538), .Z(n5539) );
  XOR U3973 ( .A(n5541), .B(n5542), .Z(n2728) );
  NOR U3974 ( .A(n5543), .B(n5541), .Z(n5542) );
  XOR U3975 ( .A(n5544), .B(n5545), .Z(n2723) );
  NOR U3976 ( .A(n5546), .B(n5544), .Z(n5545) );
  XOR U3977 ( .A(n5547), .B(n5548), .Z(n2724) );
  NOR U3978 ( .A(n5549), .B(n5547), .Z(n5548) );
  XOR U3979 ( .A(n5550), .B(n5551), .Z(n1483) );
  NOR U3980 ( .A(n5552), .B(n5550), .Z(n5551) );
  XNOR U3981 ( .A(n5553), .B(n5554), .Z(n1457) );
  NOR U3982 ( .A(n5555), .B(n5553), .Z(n5554) );
  XNOR U3983 ( .A(n5556), .B(n5557), .Z(n1462) );
  NOR U3984 ( .A(n5558), .B(n5556), .Z(n5557) );
  XOR U3985 ( .A(n5559), .B(n5560), .Z(n1464) );
  NOR U3986 ( .A(n5561), .B(n5559), .Z(n5560) );
  IV U3987 ( .A(n1474), .Z(n4154) );
  XNOR U3988 ( .A(n5562), .B(n5563), .Z(n1474) );
  NOR U3989 ( .A(n5564), .B(n5562), .Z(n5563) );
  XOR U3990 ( .A(n5565), .B(n5566), .Z(n2734) );
  NOR U3991 ( .A(n56), .B(n5567), .Z(n5566) );
  IV U3992 ( .A(n5565), .Z(n5567) );
  XOR U3993 ( .A(n5568), .B(n5569), .Z(n2737) );
  AND U3994 ( .A(n5570), .B(n5571), .Z(n5569) );
  XOR U3995 ( .A(n5568), .B(n60), .Z(n5571) );
  XOR U3996 ( .A(n4152), .B(n4151), .Z(n60) );
  XNOR U3997 ( .A(n4149), .B(n4148), .Z(n4151) );
  XNOR U3998 ( .A(n4146), .B(n4145), .Z(n4148) );
  XNOR U3999 ( .A(n4143), .B(n4142), .Z(n4145) );
  XNOR U4000 ( .A(n4140), .B(n4139), .Z(n4142) );
  XNOR U4001 ( .A(n4137), .B(n4136), .Z(n4139) );
  XNOR U4002 ( .A(n4134), .B(n4133), .Z(n4136) );
  XNOR U4003 ( .A(n4131), .B(n4130), .Z(n4133) );
  XNOR U4004 ( .A(n4128), .B(n4127), .Z(n4130) );
  XNOR U4005 ( .A(n4125), .B(n4124), .Z(n4127) );
  XNOR U4006 ( .A(n4122), .B(n4121), .Z(n4124) );
  XNOR U4007 ( .A(n4119), .B(n4118), .Z(n4121) );
  XNOR U4008 ( .A(n4116), .B(n4115), .Z(n4118) );
  XNOR U4009 ( .A(n4113), .B(n4112), .Z(n4115) );
  XNOR U4010 ( .A(n4110), .B(n4109), .Z(n4112) );
  XNOR U4011 ( .A(n4107), .B(n4106), .Z(n4109) );
  XNOR U4012 ( .A(n4104), .B(n4103), .Z(n4106) );
  XNOR U4013 ( .A(n4101), .B(n4100), .Z(n4103) );
  XNOR U4014 ( .A(n4098), .B(n4097), .Z(n4100) );
  XNOR U4015 ( .A(n4095), .B(n4094), .Z(n4097) );
  XNOR U4016 ( .A(n4092), .B(n4091), .Z(n4094) );
  XNOR U4017 ( .A(n4089), .B(n4088), .Z(n4091) );
  XNOR U4018 ( .A(n4086), .B(n4085), .Z(n4088) );
  XNOR U4019 ( .A(n4083), .B(n4082), .Z(n4085) );
  XNOR U4020 ( .A(n4080), .B(n4079), .Z(n4082) );
  XNOR U4021 ( .A(n4077), .B(n4076), .Z(n4079) );
  XNOR U4022 ( .A(n4074), .B(n4073), .Z(n4076) );
  XNOR U4023 ( .A(n4071), .B(n4070), .Z(n4073) );
  XNOR U4024 ( .A(n4068), .B(n4067), .Z(n4070) );
  XNOR U4025 ( .A(n4065), .B(n4064), .Z(n4067) );
  XNOR U4026 ( .A(n4062), .B(n4061), .Z(n4064) );
  XNOR U4027 ( .A(n4059), .B(n4058), .Z(n4061) );
  XNOR U4028 ( .A(n4056), .B(n4055), .Z(n4058) );
  XNOR U4029 ( .A(n4053), .B(n4052), .Z(n4055) );
  XNOR U4030 ( .A(n4050), .B(n4049), .Z(n4052) );
  XNOR U4031 ( .A(n4047), .B(n4046), .Z(n4049) );
  XNOR U4032 ( .A(n4044), .B(n4043), .Z(n4046) );
  XNOR U4033 ( .A(n4041), .B(n4040), .Z(n4043) );
  XNOR U4034 ( .A(n4038), .B(n4037), .Z(n4040) );
  XNOR U4035 ( .A(n4035), .B(n4034), .Z(n4037) );
  XNOR U4036 ( .A(n4032), .B(n4031), .Z(n4034) );
  XNOR U4037 ( .A(n4029), .B(n4028), .Z(n4031) );
  XNOR U4038 ( .A(n4026), .B(n4025), .Z(n4028) );
  XNOR U4039 ( .A(n4023), .B(n4022), .Z(n4025) );
  XNOR U4040 ( .A(n4020), .B(n4019), .Z(n4022) );
  XNOR U4041 ( .A(n4017), .B(n4016), .Z(n4019) );
  XNOR U4042 ( .A(n4014), .B(n4013), .Z(n4016) );
  XNOR U4043 ( .A(n4011), .B(n4010), .Z(n4013) );
  XNOR U4044 ( .A(n4008), .B(n4007), .Z(n4010) );
  XNOR U4045 ( .A(n4005), .B(n4004), .Z(n4007) );
  XNOR U4046 ( .A(n4002), .B(n4001), .Z(n4004) );
  XNOR U4047 ( .A(n3999), .B(n3998), .Z(n4001) );
  XNOR U4048 ( .A(n3996), .B(n3995), .Z(n3998) );
  XNOR U4049 ( .A(n3993), .B(n3992), .Z(n3995) );
  XNOR U4050 ( .A(n3990), .B(n3989), .Z(n3992) );
  XNOR U4051 ( .A(n3987), .B(n3986), .Z(n3989) );
  XNOR U4052 ( .A(n3984), .B(n3983), .Z(n3986) );
  XNOR U4053 ( .A(n3981), .B(n3980), .Z(n3983) );
  XNOR U4054 ( .A(n3978), .B(n3977), .Z(n3980) );
  XNOR U4055 ( .A(n3975), .B(n3974), .Z(n3977) );
  XNOR U4056 ( .A(n3972), .B(n3971), .Z(n3974) );
  XNOR U4057 ( .A(n3969), .B(n3968), .Z(n3971) );
  XNOR U4058 ( .A(n3966), .B(n3965), .Z(n3968) );
  XNOR U4059 ( .A(n3963), .B(n3962), .Z(n3965) );
  XNOR U4060 ( .A(n3960), .B(n3959), .Z(n3962) );
  XNOR U4061 ( .A(n3957), .B(n3956), .Z(n3959) );
  XNOR U4062 ( .A(n3954), .B(n3953), .Z(n3956) );
  XNOR U4063 ( .A(n3951), .B(n3950), .Z(n3953) );
  XNOR U4064 ( .A(n3948), .B(n3947), .Z(n3950) );
  XNOR U4065 ( .A(n3945), .B(n3944), .Z(n3947) );
  XNOR U4066 ( .A(n3942), .B(n3941), .Z(n3944) );
  XNOR U4067 ( .A(n3939), .B(n3938), .Z(n3941) );
  XNOR U4068 ( .A(n3936), .B(n3935), .Z(n3938) );
  XNOR U4069 ( .A(n3933), .B(n3932), .Z(n3935) );
  XNOR U4070 ( .A(n3930), .B(n3929), .Z(n3932) );
  XNOR U4071 ( .A(n3927), .B(n3926), .Z(n3929) );
  XNOR U4072 ( .A(n3924), .B(n3923), .Z(n3926) );
  XNOR U4073 ( .A(n3921), .B(n3920), .Z(n3923) );
  XNOR U4074 ( .A(n3918), .B(n3917), .Z(n3920) );
  XNOR U4075 ( .A(n3915), .B(n3914), .Z(n3917) );
  XNOR U4076 ( .A(n3912), .B(n3911), .Z(n3914) );
  XNOR U4077 ( .A(n3909), .B(n3908), .Z(n3911) );
  XNOR U4078 ( .A(n3906), .B(n3905), .Z(n3908) );
  XNOR U4079 ( .A(n3903), .B(n3902), .Z(n3905) );
  XNOR U4080 ( .A(n3900), .B(n3899), .Z(n3902) );
  XNOR U4081 ( .A(n3897), .B(n3896), .Z(n3899) );
  XNOR U4082 ( .A(n3894), .B(n3893), .Z(n3896) );
  XNOR U4083 ( .A(n3891), .B(n3890), .Z(n3893) );
  XNOR U4084 ( .A(n3888), .B(n3887), .Z(n3890) );
  XNOR U4085 ( .A(n3885), .B(n3884), .Z(n3887) );
  XNOR U4086 ( .A(n3882), .B(n3881), .Z(n3884) );
  XNOR U4087 ( .A(n3879), .B(n3878), .Z(n3881) );
  XNOR U4088 ( .A(n3876), .B(n3875), .Z(n3878) );
  XNOR U4089 ( .A(n3873), .B(n3872), .Z(n3875) );
  XNOR U4090 ( .A(n3870), .B(n3869), .Z(n3872) );
  XNOR U4091 ( .A(n3867), .B(n3866), .Z(n3869) );
  XNOR U4092 ( .A(n3864), .B(n3863), .Z(n3866) );
  XNOR U4093 ( .A(n3861), .B(n3860), .Z(n3863) );
  XNOR U4094 ( .A(n3858), .B(n3857), .Z(n3860) );
  XNOR U4095 ( .A(n3855), .B(n3854), .Z(n3857) );
  XNOR U4096 ( .A(n3852), .B(n3851), .Z(n3854) );
  XNOR U4097 ( .A(n3849), .B(n3848), .Z(n3851) );
  XNOR U4098 ( .A(n3846), .B(n3845), .Z(n3848) );
  XNOR U4099 ( .A(n3843), .B(n3842), .Z(n3845) );
  XNOR U4100 ( .A(n3840), .B(n3839), .Z(n3842) );
  XNOR U4101 ( .A(n3837), .B(n3836), .Z(n3839) );
  XNOR U4102 ( .A(n3834), .B(n3833), .Z(n3836) );
  XNOR U4103 ( .A(n3831), .B(n3830), .Z(n3833) );
  XNOR U4104 ( .A(n3828), .B(n3827), .Z(n3830) );
  XNOR U4105 ( .A(n3825), .B(n3824), .Z(n3827) );
  XNOR U4106 ( .A(n3822), .B(n3821), .Z(n3824) );
  XNOR U4107 ( .A(n3819), .B(n3818), .Z(n3821) );
  XNOR U4108 ( .A(n3816), .B(n3815), .Z(n3818) );
  XNOR U4109 ( .A(n3813), .B(n3812), .Z(n3815) );
  XNOR U4110 ( .A(n3810), .B(n3809), .Z(n3812) );
  XNOR U4111 ( .A(n3807), .B(n3806), .Z(n3809) );
  XNOR U4112 ( .A(n3804), .B(n3803), .Z(n3806) );
  XNOR U4113 ( .A(n3801), .B(n3800), .Z(n3803) );
  XNOR U4114 ( .A(n3798), .B(n3797), .Z(n3800) );
  XNOR U4115 ( .A(n3795), .B(n3794), .Z(n3797) );
  XNOR U4116 ( .A(n3792), .B(n3791), .Z(n3794) );
  XNOR U4117 ( .A(n3789), .B(n3788), .Z(n3791) );
  XNOR U4118 ( .A(n3786), .B(n3785), .Z(n3788) );
  XNOR U4119 ( .A(n3783), .B(n3782), .Z(n3785) );
  XNOR U4120 ( .A(n3780), .B(n3779), .Z(n3782) );
  XNOR U4121 ( .A(n3777), .B(n3776), .Z(n3779) );
  XNOR U4122 ( .A(n3774), .B(n3773), .Z(n3776) );
  XNOR U4123 ( .A(n3771), .B(n3770), .Z(n3773) );
  XNOR U4124 ( .A(n3768), .B(n3767), .Z(n3770) );
  XNOR U4125 ( .A(n3765), .B(n3764), .Z(n3767) );
  XNOR U4126 ( .A(n3762), .B(n3761), .Z(n3764) );
  XNOR U4127 ( .A(n3759), .B(n3758), .Z(n3761) );
  XNOR U4128 ( .A(n3756), .B(n3755), .Z(n3758) );
  XNOR U4129 ( .A(n3753), .B(n3752), .Z(n3755) );
  XNOR U4130 ( .A(n3750), .B(n3749), .Z(n3752) );
  XNOR U4131 ( .A(n3747), .B(n3746), .Z(n3749) );
  XNOR U4132 ( .A(n3744), .B(n3743), .Z(n3746) );
  XNOR U4133 ( .A(n3741), .B(n3740), .Z(n3743) );
  XNOR U4134 ( .A(n3738), .B(n3737), .Z(n3740) );
  XNOR U4135 ( .A(n3735), .B(n3734), .Z(n3737) );
  XNOR U4136 ( .A(n3732), .B(n3731), .Z(n3734) );
  XNOR U4137 ( .A(n3729), .B(n3728), .Z(n3731) );
  XNOR U4138 ( .A(n3726), .B(n3725), .Z(n3728) );
  XNOR U4139 ( .A(n3723), .B(n3722), .Z(n3725) );
  XNOR U4140 ( .A(n3720), .B(n3719), .Z(n3722) );
  XNOR U4141 ( .A(n3717), .B(n3716), .Z(n3719) );
  XNOR U4142 ( .A(n3714), .B(n3713), .Z(n3716) );
  XNOR U4143 ( .A(n3711), .B(n3710), .Z(n3713) );
  XNOR U4144 ( .A(n3708), .B(n3707), .Z(n3710) );
  XNOR U4145 ( .A(n3705), .B(n3704), .Z(n3707) );
  XNOR U4146 ( .A(n3702), .B(n3701), .Z(n3704) );
  XNOR U4147 ( .A(n3699), .B(n3698), .Z(n3701) );
  XNOR U4148 ( .A(n3696), .B(n3695), .Z(n3698) );
  XNOR U4149 ( .A(n3693), .B(n3692), .Z(n3695) );
  XNOR U4150 ( .A(n3690), .B(n3689), .Z(n3692) );
  XNOR U4151 ( .A(n3687), .B(n3686), .Z(n3689) );
  XNOR U4152 ( .A(n3684), .B(n3683), .Z(n3686) );
  XNOR U4153 ( .A(n3681), .B(n3680), .Z(n3683) );
  XNOR U4154 ( .A(n3678), .B(n3677), .Z(n3680) );
  XNOR U4155 ( .A(n3675), .B(n3674), .Z(n3677) );
  XNOR U4156 ( .A(n3672), .B(n3671), .Z(n3674) );
  XNOR U4157 ( .A(n3669), .B(n3668), .Z(n3671) );
  XNOR U4158 ( .A(n3666), .B(n3665), .Z(n3668) );
  XNOR U4159 ( .A(n3663), .B(n3662), .Z(n3665) );
  XNOR U4160 ( .A(n3660), .B(n3659), .Z(n3662) );
  XNOR U4161 ( .A(n3657), .B(n3656), .Z(n3659) );
  XNOR U4162 ( .A(n3654), .B(n3653), .Z(n3656) );
  XNOR U4163 ( .A(n3651), .B(n3650), .Z(n3653) );
  XNOR U4164 ( .A(n3648), .B(n3647), .Z(n3650) );
  XNOR U4165 ( .A(n3645), .B(n3644), .Z(n3647) );
  XNOR U4166 ( .A(n3642), .B(n3641), .Z(n3644) );
  XNOR U4167 ( .A(n3639), .B(n3638), .Z(n3641) );
  XNOR U4168 ( .A(n3636), .B(n3635), .Z(n3638) );
  XNOR U4169 ( .A(n3633), .B(n3632), .Z(n3635) );
  XNOR U4170 ( .A(n3630), .B(n3629), .Z(n3632) );
  XNOR U4171 ( .A(n3627), .B(n3626), .Z(n3629) );
  XNOR U4172 ( .A(n3624), .B(n3623), .Z(n3626) );
  XNOR U4173 ( .A(n3621), .B(n3620), .Z(n3623) );
  XNOR U4174 ( .A(n3618), .B(n3617), .Z(n3620) );
  XNOR U4175 ( .A(n3615), .B(n3614), .Z(n3617) );
  XNOR U4176 ( .A(n3612), .B(n3611), .Z(n3614) );
  XNOR U4177 ( .A(n3609), .B(n3608), .Z(n3611) );
  XNOR U4178 ( .A(n3606), .B(n3605), .Z(n3608) );
  XNOR U4179 ( .A(n3603), .B(n3602), .Z(n3605) );
  XNOR U4180 ( .A(n3600), .B(n3599), .Z(n3602) );
  XNOR U4181 ( .A(n3597), .B(n3596), .Z(n3599) );
  XNOR U4182 ( .A(n3594), .B(n3593), .Z(n3596) );
  XNOR U4183 ( .A(n3591), .B(n3590), .Z(n3593) );
  XNOR U4184 ( .A(n3588), .B(n3587), .Z(n3590) );
  XNOR U4185 ( .A(n3585), .B(n3584), .Z(n3587) );
  XNOR U4186 ( .A(n3582), .B(n3581), .Z(n3584) );
  XNOR U4187 ( .A(n3579), .B(n3578), .Z(n3581) );
  XNOR U4188 ( .A(n3576), .B(n3575), .Z(n3578) );
  XNOR U4189 ( .A(n3573), .B(n3572), .Z(n3575) );
  XNOR U4190 ( .A(n3570), .B(n3569), .Z(n3572) );
  XNOR U4191 ( .A(n3567), .B(n3566), .Z(n3569) );
  XNOR U4192 ( .A(n3564), .B(n3563), .Z(n3566) );
  XNOR U4193 ( .A(n3561), .B(n3560), .Z(n3563) );
  XNOR U4194 ( .A(n3558), .B(n3557), .Z(n3560) );
  XNOR U4195 ( .A(n3555), .B(n3554), .Z(n3557) );
  XNOR U4196 ( .A(n3552), .B(n3551), .Z(n3554) );
  XNOR U4197 ( .A(n3549), .B(n3548), .Z(n3551) );
  XNOR U4198 ( .A(n3546), .B(n3545), .Z(n3548) );
  XNOR U4199 ( .A(n3543), .B(n3542), .Z(n3545) );
  XNOR U4200 ( .A(n3540), .B(n3539), .Z(n3542) );
  XNOR U4201 ( .A(n3537), .B(n3536), .Z(n3539) );
  XNOR U4202 ( .A(n3534), .B(n3533), .Z(n3536) );
  XNOR U4203 ( .A(n3531), .B(n3530), .Z(n3533) );
  XNOR U4204 ( .A(n3528), .B(n3527), .Z(n3530) );
  XNOR U4205 ( .A(n3525), .B(n3524), .Z(n3527) );
  XNOR U4206 ( .A(n3522), .B(n3521), .Z(n3524) );
  XNOR U4207 ( .A(n3519), .B(n3518), .Z(n3521) );
  XNOR U4208 ( .A(n3516), .B(n3515), .Z(n3518) );
  XNOR U4209 ( .A(n3513), .B(n3512), .Z(n3515) );
  XNOR U4210 ( .A(n3510), .B(n3509), .Z(n3512) );
  XNOR U4211 ( .A(n3507), .B(n3506), .Z(n3509) );
  XNOR U4212 ( .A(n3504), .B(n3503), .Z(n3506) );
  XNOR U4213 ( .A(n3501), .B(n3500), .Z(n3503) );
  XNOR U4214 ( .A(n3498), .B(n3497), .Z(n3500) );
  XNOR U4215 ( .A(n3495), .B(n3494), .Z(n3497) );
  XNOR U4216 ( .A(n3492), .B(n3491), .Z(n3494) );
  XNOR U4217 ( .A(n3489), .B(n3488), .Z(n3491) );
  XNOR U4218 ( .A(n3486), .B(n3485), .Z(n3488) );
  XNOR U4219 ( .A(n3483), .B(n3482), .Z(n3485) );
  XNOR U4220 ( .A(n3480), .B(n3479), .Z(n3482) );
  XNOR U4221 ( .A(n3477), .B(n3476), .Z(n3479) );
  XNOR U4222 ( .A(n3474), .B(n3473), .Z(n3476) );
  XNOR U4223 ( .A(n3471), .B(n3470), .Z(n3473) );
  XNOR U4224 ( .A(n3468), .B(n3467), .Z(n3470) );
  XNOR U4225 ( .A(n3465), .B(n3464), .Z(n3467) );
  XNOR U4226 ( .A(n3462), .B(n3461), .Z(n3464) );
  XNOR U4227 ( .A(n3459), .B(n3458), .Z(n3461) );
  XNOR U4228 ( .A(n3456), .B(n3455), .Z(n3458) );
  XNOR U4229 ( .A(n3453), .B(n3452), .Z(n3455) );
  XNOR U4230 ( .A(n3450), .B(n3449), .Z(n3452) );
  XNOR U4231 ( .A(n3447), .B(n3446), .Z(n3449) );
  XNOR U4232 ( .A(n3444), .B(n3443), .Z(n3446) );
  XNOR U4233 ( .A(n3441), .B(n3440), .Z(n3443) );
  XNOR U4234 ( .A(n3438), .B(n3437), .Z(n3440) );
  XNOR U4235 ( .A(n3435), .B(n3434), .Z(n3437) );
  XNOR U4236 ( .A(n3432), .B(n3431), .Z(n3434) );
  XNOR U4237 ( .A(n3429), .B(n3428), .Z(n3431) );
  XNOR U4238 ( .A(n3426), .B(n3425), .Z(n3428) );
  XNOR U4239 ( .A(n3423), .B(n3422), .Z(n3425) );
  XNOR U4240 ( .A(n3420), .B(n3419), .Z(n3422) );
  XNOR U4241 ( .A(n3417), .B(n3416), .Z(n3419) );
  XNOR U4242 ( .A(n3414), .B(n3413), .Z(n3416) );
  XNOR U4243 ( .A(n3411), .B(n3410), .Z(n3413) );
  XNOR U4244 ( .A(n3408), .B(n3407), .Z(n3410) );
  XNOR U4245 ( .A(n3405), .B(n3404), .Z(n3407) );
  XNOR U4246 ( .A(n3402), .B(n3401), .Z(n3404) );
  XNOR U4247 ( .A(n3399), .B(n3398), .Z(n3401) );
  XNOR U4248 ( .A(n3396), .B(n3395), .Z(n3398) );
  XNOR U4249 ( .A(n3393), .B(n3392), .Z(n3395) );
  XNOR U4250 ( .A(n3390), .B(n3389), .Z(n3392) );
  XNOR U4251 ( .A(n3387), .B(n3386), .Z(n3389) );
  XNOR U4252 ( .A(n3384), .B(n3382), .Z(n3386) );
  XNOR U4253 ( .A(n3383), .B(n2750), .Z(n3382) );
  XNOR U4254 ( .A(n2751), .B(n2748), .Z(n2750) );
  XNOR U4255 ( .A(n2749), .B(n2752), .Z(n2748) );
  XNOR U4256 ( .A(n2753), .B(n3377), .Z(n2752) );
  XNOR U4257 ( .A(n2760), .B(n3376), .Z(n3377) );
  XNOR U4258 ( .A(n3369), .B(n3373), .Z(n3376) );
  XNOR U4259 ( .A(n3368), .B(n3366), .Z(n3373) );
  XNOR U4260 ( .A(n3367), .B(n3365), .Z(n3366) );
  XNOR U4261 ( .A(n2767), .B(n3360), .Z(n3365) );
  XNOR U4262 ( .A(n2766), .B(n3358), .Z(n3360) );
  XNOR U4263 ( .A(n3359), .B(n3354), .Z(n3358) );
  XNOR U4264 ( .A(n3355), .B(n2782), .Z(n3354) );
  XNOR U4265 ( .A(n2777), .B(n3353), .Z(n2782) );
  XNOR U4266 ( .A(n2776), .B(n3348), .Z(n3353) );
  XNOR U4267 ( .A(n2778), .B(n3347), .Z(n3348) );
  XNOR U4268 ( .A(n2781), .B(n3344), .Z(n3347) );
  XNOR U4269 ( .A(n2787), .B(n3343), .Z(n3344) );
  XNOR U4270 ( .A(n3336), .B(n3340), .Z(n3343) );
  XNOR U4271 ( .A(n3335), .B(n3333), .Z(n3340) );
  XNOR U4272 ( .A(n3334), .B(n3332), .Z(n3333) );
  XNOR U4273 ( .A(n2794), .B(n3327), .Z(n3332) );
  XNOR U4274 ( .A(n2793), .B(n3325), .Z(n3327) );
  XNOR U4275 ( .A(n3326), .B(n3321), .Z(n3325) );
  XNOR U4276 ( .A(n3322), .B(n2809), .Z(n3321) );
  XNOR U4277 ( .A(n2804), .B(n3320), .Z(n2809) );
  XNOR U4278 ( .A(n2803), .B(n3315), .Z(n3320) );
  XNOR U4279 ( .A(n2805), .B(n3314), .Z(n3315) );
  XNOR U4280 ( .A(n2808), .B(n3311), .Z(n3314) );
  XNOR U4281 ( .A(n2814), .B(n3310), .Z(n3311) );
  XNOR U4282 ( .A(n3303), .B(n3307), .Z(n3310) );
  XNOR U4283 ( .A(n3302), .B(n3300), .Z(n3307) );
  XNOR U4284 ( .A(n3301), .B(n3299), .Z(n3300) );
  XNOR U4285 ( .A(n2821), .B(n3294), .Z(n3299) );
  XNOR U4286 ( .A(n2820), .B(n3292), .Z(n3294) );
  XNOR U4287 ( .A(n3293), .B(n3288), .Z(n3292) );
  XNOR U4288 ( .A(n3289), .B(n2836), .Z(n3288) );
  XNOR U4289 ( .A(n2831), .B(n3287), .Z(n2836) );
  XNOR U4290 ( .A(n2830), .B(n3282), .Z(n3287) );
  XNOR U4291 ( .A(n2832), .B(n3281), .Z(n3282) );
  XNOR U4292 ( .A(n2835), .B(n3278), .Z(n3281) );
  XNOR U4293 ( .A(n2841), .B(n3277), .Z(n3278) );
  XNOR U4294 ( .A(n3270), .B(n3274), .Z(n3277) );
  XNOR U4295 ( .A(n3269), .B(n3267), .Z(n3274) );
  XNOR U4296 ( .A(n3268), .B(n3266), .Z(n3267) );
  XNOR U4297 ( .A(n2848), .B(n3261), .Z(n3266) );
  XNOR U4298 ( .A(n2847), .B(n3259), .Z(n3261) );
  XNOR U4299 ( .A(n3260), .B(n3255), .Z(n3259) );
  XNOR U4300 ( .A(n3256), .B(n2863), .Z(n3255) );
  XNOR U4301 ( .A(n2858), .B(n3254), .Z(n2863) );
  XNOR U4302 ( .A(n2857), .B(n3249), .Z(n3254) );
  XNOR U4303 ( .A(n2859), .B(n3248), .Z(n3249) );
  XNOR U4304 ( .A(n2862), .B(n3245), .Z(n3248) );
  XNOR U4305 ( .A(n2868), .B(n3244), .Z(n3245) );
  XNOR U4306 ( .A(n3237), .B(n3241), .Z(n3244) );
  XNOR U4307 ( .A(n3236), .B(n3234), .Z(n3241) );
  XNOR U4308 ( .A(n3235), .B(n3233), .Z(n3234) );
  XNOR U4309 ( .A(n2875), .B(n3228), .Z(n3233) );
  XNOR U4310 ( .A(n2874), .B(n3226), .Z(n3228) );
  XNOR U4311 ( .A(n3227), .B(n3222), .Z(n3226) );
  XNOR U4312 ( .A(n3223), .B(n2890), .Z(n3222) );
  XNOR U4313 ( .A(n2885), .B(n3221), .Z(n2890) );
  XNOR U4314 ( .A(n2884), .B(n3216), .Z(n3221) );
  XNOR U4315 ( .A(n2886), .B(n3215), .Z(n3216) );
  XNOR U4316 ( .A(n2889), .B(n3212), .Z(n3215) );
  XNOR U4317 ( .A(n2895), .B(n3211), .Z(n3212) );
  XNOR U4318 ( .A(n3204), .B(n3208), .Z(n3211) );
  XNOR U4319 ( .A(n3203), .B(n3201), .Z(n3208) );
  XNOR U4320 ( .A(n3202), .B(n3200), .Z(n3201) );
  XNOR U4321 ( .A(n2902), .B(n3195), .Z(n3200) );
  XNOR U4322 ( .A(n2901), .B(n3193), .Z(n3195) );
  XNOR U4323 ( .A(n3194), .B(n3189), .Z(n3193) );
  XNOR U4324 ( .A(n3190), .B(n2917), .Z(n3189) );
  XNOR U4325 ( .A(n2912), .B(n3188), .Z(n2917) );
  XNOR U4326 ( .A(n2911), .B(n3183), .Z(n3188) );
  XNOR U4327 ( .A(n2913), .B(n3182), .Z(n3183) );
  XNOR U4328 ( .A(n2916), .B(n3179), .Z(n3182) );
  XNOR U4329 ( .A(n2922), .B(n3178), .Z(n3179) );
  XNOR U4330 ( .A(n3171), .B(n3175), .Z(n3178) );
  XNOR U4331 ( .A(n3170), .B(n3168), .Z(n3175) );
  XNOR U4332 ( .A(n3169), .B(n3167), .Z(n3168) );
  XNOR U4333 ( .A(n2929), .B(n3162), .Z(n3167) );
  XNOR U4334 ( .A(n2928), .B(n3160), .Z(n3162) );
  XNOR U4335 ( .A(n3161), .B(n3156), .Z(n3160) );
  XNOR U4336 ( .A(n3157), .B(n2944), .Z(n3156) );
  XNOR U4337 ( .A(n2939), .B(n3155), .Z(n2944) );
  XNOR U4338 ( .A(n2938), .B(n3150), .Z(n3155) );
  XNOR U4339 ( .A(n2940), .B(n3149), .Z(n3150) );
  XNOR U4340 ( .A(n2943), .B(n3146), .Z(n3149) );
  XNOR U4341 ( .A(n2949), .B(n3145), .Z(n3146) );
  XNOR U4342 ( .A(n3138), .B(n3142), .Z(n3145) );
  XNOR U4343 ( .A(n3137), .B(n3135), .Z(n3142) );
  XNOR U4344 ( .A(n3136), .B(n3134), .Z(n3135) );
  XNOR U4345 ( .A(n2956), .B(n3129), .Z(n3134) );
  XNOR U4346 ( .A(n2955), .B(n3127), .Z(n3129) );
  XNOR U4347 ( .A(n3128), .B(n3123), .Z(n3127) );
  XNOR U4348 ( .A(n3124), .B(n2971), .Z(n3123) );
  XNOR U4349 ( .A(n2966), .B(n3122), .Z(n2971) );
  XNOR U4350 ( .A(n2965), .B(n3117), .Z(n3122) );
  XNOR U4351 ( .A(n2967), .B(n3116), .Z(n3117) );
  XNOR U4352 ( .A(n2970), .B(n3113), .Z(n3116) );
  XNOR U4353 ( .A(n2976), .B(n3112), .Z(n3113) );
  XNOR U4354 ( .A(n3105), .B(n3109), .Z(n3112) );
  XNOR U4355 ( .A(n3104), .B(n3102), .Z(n3109) );
  XNOR U4356 ( .A(n3103), .B(n3101), .Z(n3102) );
  XNOR U4357 ( .A(n2983), .B(n3096), .Z(n3101) );
  XNOR U4358 ( .A(n2982), .B(n3094), .Z(n3096) );
  XNOR U4359 ( .A(n3095), .B(n3090), .Z(n3094) );
  XNOR U4360 ( .A(n3091), .B(n2998), .Z(n3090) );
  XNOR U4361 ( .A(n2993), .B(n3089), .Z(n2998) );
  XNOR U4362 ( .A(n2992), .B(n3084), .Z(n3089) );
  XNOR U4363 ( .A(n2994), .B(n3083), .Z(n3084) );
  XNOR U4364 ( .A(n2997), .B(n3080), .Z(n3083) );
  XNOR U4365 ( .A(n3003), .B(n3079), .Z(n3080) );
  XNOR U4366 ( .A(n3072), .B(n3076), .Z(n3079) );
  XNOR U4367 ( .A(n3071), .B(n3069), .Z(n3076) );
  XNOR U4368 ( .A(n3070), .B(n3068), .Z(n3069) );
  XNOR U4369 ( .A(n3010), .B(n3063), .Z(n3068) );
  XNOR U4370 ( .A(n3009), .B(n3061), .Z(n3063) );
  XNOR U4371 ( .A(n3062), .B(n3057), .Z(n3061) );
  XNOR U4372 ( .A(n3058), .B(n3025), .Z(n3057) );
  XNOR U4373 ( .A(n3020), .B(n3056), .Z(n3025) );
  XNOR U4374 ( .A(n3019), .B(n3051), .Z(n3056) );
  XNOR U4375 ( .A(n3021), .B(n3050), .Z(n3051) );
  XNOR U4376 ( .A(n3024), .B(n3047), .Z(n3050) );
  XNOR U4377 ( .A(n3030), .B(n3046), .Z(n3047) );
  XNOR U4378 ( .A(n3033), .B(n3043), .Z(n3046) );
  XNOR U4379 ( .A(n3032), .B(n3040), .Z(n3043) );
  XOR U4380 ( .A(n3041), .B(n3039), .Z(n3040) );
  XNOR U4381 ( .A(n5572), .B(n5573), .Z(n3039) );
  XOR U4382 ( .A(n5574), .B(n5575), .Z(n5573) );
  XOR U4383 ( .A(n5576), .B(n5577), .Z(n5575) );
  NOR U4384 ( .A(n5578), .B(n5579), .Z(n5576) );
  XOR U4385 ( .A(n5580), .B(n5581), .Z(n5574) );
  NOR U4386 ( .A(n5582), .B(n5583), .Z(n5581) );
  AND U4387 ( .A(n5584), .B(n5585), .Z(n5580) );
  XOR U4388 ( .A(n5586), .B(n5587), .Z(n5572) );
  XOR U4389 ( .A(n5579), .B(n5583), .Z(n5587) );
  XOR U4390 ( .A(n5588), .B(n5585), .Z(n5586) );
  XOR U4391 ( .A(n5589), .B(n5590), .Z(n5588) );
  XOR U4392 ( .A(n5591), .B(n5592), .Z(n5590) );
  XOR U4393 ( .A(n5593), .B(n5594), .Z(n5592) );
  XOR U4394 ( .A(n5595), .B(n5596), .Z(n5591) );
  NOR U4395 ( .A(n5597), .B(n5598), .Z(n5596) );
  AND U4396 ( .A(n5599), .B(n5577), .Z(n5595) );
  XOR U4397 ( .A(n5600), .B(n5601), .Z(n5589) );
  XOR U4398 ( .A(n5602), .B(n5603), .Z(n5601) );
  XOR U4399 ( .A(n5604), .B(n5605), .Z(n5603) );
  XOR U4400 ( .A(n5606), .B(n5607), .Z(n5605) );
  XOR U4401 ( .A(n5608), .B(n5609), .Z(n5607) );
  XOR U4402 ( .A(n5610), .B(n5611), .Z(n5609) );
  XNOR U4403 ( .A(n5612), .B(n5613), .Z(n5608) );
  XOR U4404 ( .A(n5614), .B(n5615), .Z(n5613) );
  NOR U4405 ( .A(n5616), .B(n5611), .Z(n5614) );
  XOR U4406 ( .A(n5617), .B(n5618), .Z(n5606) );
  XOR U4407 ( .A(n5619), .B(n5620), .Z(n5618) );
  XOR U4408 ( .A(n5621), .B(n5622), .Z(n5620) );
  XOR U4409 ( .A(n5623), .B(n5624), .Z(n5622) );
  XOR U4410 ( .A(n5625), .B(n5626), .Z(n5624) );
  XOR U4411 ( .A(n5627), .B(n5628), .Z(n5626) );
  XOR U4412 ( .A(n5629), .B(n5630), .Z(n5628) );
  XOR U4413 ( .A(n5631), .B(n5632), .Z(n5630) );
  NOR U4414 ( .A(n5633), .B(n5634), .Z(n5632) );
  XOR U4415 ( .A(n5635), .B(n5636), .Z(n5629) );
  AND U4416 ( .A(n5631), .B(n5637), .Z(n5635) );
  XOR U4417 ( .A(n5638), .B(n5639), .Z(n5627) );
  XOR U4418 ( .A(n5640), .B(n5641), .Z(n5639) );
  XOR U4419 ( .A(n5642), .B(n5643), .Z(n5641) );
  XOR U4420 ( .A(n5644), .B(n5645), .Z(n5643) );
  XOR U4421 ( .A(n5646), .B(n5647), .Z(n5645) );
  XOR U4422 ( .A(n5648), .B(n5649), .Z(n5647) );
  XOR U4423 ( .A(n5650), .B(n5651), .Z(n5649) );
  XOR U4424 ( .A(n5652), .B(n5653), .Z(n5651) );
  XOR U4425 ( .A(n5654), .B(n5655), .Z(n5653) );
  AND U4426 ( .A(n5656), .B(n5657), .Z(n5655) );
  NOR U4427 ( .A(n5658), .B(n5659), .Z(n5657) );
  NOR U4428 ( .A(n5660), .B(n5661), .Z(n5656) );
  AND U4429 ( .A(n5662), .B(n5663), .Z(n5661) );
  AND U4430 ( .A(n5664), .B(n5665), .Z(n5654) );
  NOR U4431 ( .A(n5666), .B(n5667), .Z(n5665) );
  NOR U4432 ( .A(n5668), .B(n5669), .Z(n5664) );
  AND U4433 ( .A(n5670), .B(n5671), .Z(n5669) );
  XOR U4434 ( .A(n5672), .B(n5673), .Z(n5652) );
  AND U4435 ( .A(n5674), .B(n5675), .Z(n5673) );
  NOR U4436 ( .A(n5676), .B(n5677), .Z(n5675) );
  NOR U4437 ( .A(n5678), .B(n5679), .Z(n5674) );
  AND U4438 ( .A(n5680), .B(n5681), .Z(n5679) );
  AND U4439 ( .A(n5682), .B(n5683), .Z(n5672) );
  NOR U4440 ( .A(n5684), .B(n5685), .Z(n5683) );
  AND U4441 ( .A(n5677), .B(n5686), .Z(n5685) );
  AND U4442 ( .A(n5678), .B(n5687), .Z(n5684) );
  NOR U4443 ( .A(n5688), .B(n5689), .Z(n5682) );
  XOR U4444 ( .A(n5690), .B(n5691), .Z(n5689) );
  AND U4445 ( .A(n5692), .B(n5693), .Z(n5691) );
  NOR U4446 ( .A(n5694), .B(n5695), .Z(n5693) );
  NOR U4447 ( .A(n5696), .B(n5697), .Z(n5692) );
  AND U4448 ( .A(n5698), .B(n5699), .Z(n5697) );
  AND U4449 ( .A(n5700), .B(n5701), .Z(n5690) );
  NOR U4450 ( .A(n5702), .B(n5703), .Z(n5701) );
  AND U4451 ( .A(n5695), .B(n5704), .Z(n5703) );
  AND U4452 ( .A(n5696), .B(n5705), .Z(n5702) );
  NOR U4453 ( .A(n5706), .B(n5707), .Z(n5700) );
  XOR U4454 ( .A(n5708), .B(n5709), .Z(n5707) );
  AND U4455 ( .A(n5710), .B(n5711), .Z(n5709) );
  NOR U4456 ( .A(n5712), .B(n5713), .Z(n5711) );
  NOR U4457 ( .A(n5714), .B(n5715), .Z(n5710) );
  AND U4458 ( .A(n5716), .B(n5717), .Z(n5715) );
  AND U4459 ( .A(n5718), .B(n5719), .Z(n5708) );
  AND U4460 ( .A(n5720), .B(n5721), .Z(n5719) );
  IV U4461 ( .A(n5712), .Z(n5720) );
  NOR U4462 ( .A(n5714), .B(n5722), .Z(n5718) );
  AND U4463 ( .A(n5723), .B(n5724), .Z(n5722) );
  AND U4464 ( .A(n5725), .B(n5726), .Z(n5724) );
  NOR U4465 ( .A(n5727), .B(n5728), .Z(n5725) );
  NOR U4466 ( .A(n5729), .B(n5730), .Z(n5723) );
  AND U4467 ( .A(n5694), .B(n5731), .Z(n5706) );
  AND U4468 ( .A(n5676), .B(n5732), .Z(n5688) );
  XOR U4469 ( .A(n5733), .B(n5734), .Z(n5650) );
  XOR U4470 ( .A(n5735), .B(n5736), .Z(n5734) );
  NOR U4471 ( .A(n5737), .B(n5738), .Z(n5736) );
  AND U4472 ( .A(n5667), .B(n5739), .Z(n5738) );
  AND U4473 ( .A(n5668), .B(n5740), .Z(n5737) );
  NOR U4474 ( .A(n5741), .B(n5742), .Z(n5735) );
  AND U4475 ( .A(n5659), .B(n5743), .Z(n5742) );
  AND U4476 ( .A(n5660), .B(n5744), .Z(n5741) );
  XOR U4477 ( .A(n5745), .B(n5746), .Z(n5733) );
  AND U4478 ( .A(n5666), .B(n5747), .Z(n5746) );
  AND U4479 ( .A(n5658), .B(n5748), .Z(n5745) );
  AND U4480 ( .A(n5749), .B(n5750), .Z(n5648) );
  NOR U4481 ( .A(n5751), .B(n5752), .Z(n5750) );
  NOR U4482 ( .A(n5753), .B(n5754), .Z(n5749) );
  AND U4483 ( .A(n5755), .B(n5756), .Z(n5754) );
  XOR U4484 ( .A(n5757), .B(n5758), .Z(n5646) );
  AND U4485 ( .A(n5759), .B(n5760), .Z(n5758) );
  NOR U4486 ( .A(n5761), .B(n5762), .Z(n5760) );
  NOR U4487 ( .A(n5763), .B(n5764), .Z(n5759) );
  AND U4488 ( .A(n5765), .B(n5766), .Z(n5764) );
  NOR U4489 ( .A(n5767), .B(n5768), .Z(n5757) );
  AND U4490 ( .A(n5762), .B(n5769), .Z(n5768) );
  AND U4491 ( .A(n5763), .B(n5770), .Z(n5767) );
  XOR U4492 ( .A(n5771), .B(n5772), .Z(n5644) );
  XOR U4493 ( .A(n5773), .B(n5774), .Z(n5772) );
  NOR U4494 ( .A(n5775), .B(n5776), .Z(n5774) );
  AND U4495 ( .A(n5752), .B(n5777), .Z(n5776) );
  AND U4496 ( .A(n5753), .B(n5778), .Z(n5775) );
  AND U4497 ( .A(n5761), .B(n5779), .Z(n5773) );
  XOR U4498 ( .A(n5780), .B(n5781), .Z(n5771) );
  AND U4499 ( .A(n5751), .B(n5782), .Z(n5781) );
  AND U4500 ( .A(n5783), .B(n5784), .Z(n5780) );
  AND U4501 ( .A(n5785), .B(n5786), .Z(n5642) );
  NOR U4502 ( .A(n5787), .B(n5788), .Z(n5786) );
  NOR U4503 ( .A(n5789), .B(n5790), .Z(n5785) );
  AND U4504 ( .A(n5791), .B(n5792), .Z(n5790) );
  XOR U4505 ( .A(n5793), .B(n5794), .Z(n5640) );
  AND U4506 ( .A(n5795), .B(n5796), .Z(n5794) );
  NOR U4507 ( .A(n5783), .B(n5797), .Z(n5796) );
  NOR U4508 ( .A(n5798), .B(n5799), .Z(n5795) );
  AND U4509 ( .A(n5800), .B(n5801), .Z(n5799) );
  NOR U4510 ( .A(n5802), .B(n5803), .Z(n5793) );
  AND U4511 ( .A(n5797), .B(n5804), .Z(n5803) );
  AND U4512 ( .A(n5798), .B(n5805), .Z(n5802) );
  XOR U4513 ( .A(n5806), .B(n5807), .Z(n5638) );
  XOR U4514 ( .A(n5808), .B(n5809), .Z(n5807) );
  NOR U4515 ( .A(n5810), .B(n5811), .Z(n5809) );
  AND U4516 ( .A(n5788), .B(n5812), .Z(n5811) );
  AND U4517 ( .A(n5789), .B(n5813), .Z(n5810) );
  NOR U4518 ( .A(n5814), .B(n5815), .Z(n5808) );
  AND U4519 ( .A(n5816), .B(n5817), .Z(n5815) );
  AND U4520 ( .A(n5818), .B(n5819), .Z(n5814) );
  XOR U4521 ( .A(n5820), .B(n5821), .Z(n5806) );
  AND U4522 ( .A(n5787), .B(n5822), .Z(n5821) );
  AND U4523 ( .A(n5823), .B(n5824), .Z(n5820) );
  XOR U4524 ( .A(n5825), .B(n5826), .Z(n5625) );
  NOR U4525 ( .A(n5818), .B(n5827), .Z(n5826) );
  AND U4526 ( .A(n5828), .B(n5829), .Z(n5827) );
  NOR U4527 ( .A(n5823), .B(n5816), .Z(n5825) );
  XOR U4528 ( .A(n5830), .B(n5831), .Z(n5623) );
  XOR U4529 ( .A(n5832), .B(n5833), .Z(n5831) );
  AND U4530 ( .A(n5633), .B(n5834), .Z(n5833) );
  AND U4531 ( .A(n5634), .B(n5835), .Z(n5832) );
  XOR U4532 ( .A(n5836), .B(n5837), .Z(n5830) );
  AND U4533 ( .A(n5636), .B(n5838), .Z(n5837) );
  AND U4534 ( .A(n5839), .B(n5840), .Z(n5836) );
  XNOR U4535 ( .A(n5841), .B(n5842), .Z(n5619) );
  XOR U4536 ( .A(n5843), .B(n5844), .Z(n5617) );
  XOR U4537 ( .A(n5845), .B(n5839), .Z(n5844) );
  AND U4538 ( .A(n5846), .B(n5841), .Z(n5845) );
  XOR U4539 ( .A(n5847), .B(n5848), .Z(n5843) );
  AND U4540 ( .A(n5849), .B(n5850), .Z(n5848) );
  AND U4541 ( .A(n5851), .B(n5621), .Z(n5847) );
  XOR U4542 ( .A(n5852), .B(n5853), .Z(n5604) );
  AND U4543 ( .A(n5854), .B(n5615), .Z(n5853) );
  NOR U4544 ( .A(n5855), .B(n5612), .Z(n5852) );
  XOR U4545 ( .A(n5856), .B(n5857), .Z(n5602) );
  XOR U4546 ( .A(n5858), .B(n5859), .Z(n5857) );
  NOR U4547 ( .A(n5860), .B(n5610), .Z(n5859) );
  NOR U4548 ( .A(n5861), .B(n5593), .Z(n5858) );
  XOR U4549 ( .A(n5862), .B(n5863), .Z(n5856) );
  NOR U4550 ( .A(n5864), .B(n5594), .Z(n5863) );
  NOR U4551 ( .A(n5865), .B(n5866), .Z(n5862) );
  XNOR U4552 ( .A(n5598), .B(n5866), .Z(n5600) );
  XOR U4553 ( .A(n5867), .B(n5868), .Z(n3041) );
  NOR U4554 ( .A(n5869), .B(n5867), .Z(n5868) );
  XOR U4555 ( .A(n5870), .B(n5871), .Z(n3032) );
  NOR U4556 ( .A(n5872), .B(n5870), .Z(n5871) );
  XOR U4557 ( .A(n5873), .B(n5874), .Z(n3033) );
  NOR U4558 ( .A(n5875), .B(n5873), .Z(n5874) );
  XOR U4559 ( .A(n5876), .B(n5877), .Z(n3030) );
  NOR U4560 ( .A(n5878), .B(n5876), .Z(n5877) );
  XOR U4561 ( .A(n5879), .B(n5880), .Z(n3024) );
  NOR U4562 ( .A(n5881), .B(n5879), .Z(n5880) );
  XOR U4563 ( .A(n5882), .B(n5883), .Z(n3021) );
  NOR U4564 ( .A(n5884), .B(n5882), .Z(n5883) );
  XOR U4565 ( .A(n5885), .B(n5886), .Z(n3019) );
  NOR U4566 ( .A(n5887), .B(n5885), .Z(n5886) );
  XOR U4567 ( .A(n5888), .B(n5889), .Z(n3020) );
  NOR U4568 ( .A(n5890), .B(n5888), .Z(n5889) );
  XOR U4569 ( .A(n5891), .B(n5892), .Z(n3058) );
  NOR U4570 ( .A(n5893), .B(n5891), .Z(n5892) );
  XOR U4571 ( .A(n5894), .B(n5895), .Z(n3062) );
  NOR U4572 ( .A(n5896), .B(n5894), .Z(n5895) );
  XOR U4573 ( .A(n5897), .B(n5898), .Z(n3009) );
  NOR U4574 ( .A(n5899), .B(n5897), .Z(n5898) );
  XOR U4575 ( .A(n5900), .B(n5901), .Z(n3010) );
  NOR U4576 ( .A(n5902), .B(n5900), .Z(n5901) );
  XOR U4577 ( .A(n5903), .B(n5904), .Z(n3070) );
  NOR U4578 ( .A(n5905), .B(n5903), .Z(n5904) );
  XOR U4579 ( .A(n5906), .B(n5907), .Z(n3071) );
  NOR U4580 ( .A(n5908), .B(n5906), .Z(n5907) );
  XOR U4581 ( .A(n5909), .B(n5910), .Z(n3072) );
  NOR U4582 ( .A(n5911), .B(n5909), .Z(n5910) );
  XOR U4583 ( .A(n5912), .B(n5913), .Z(n3003) );
  NOR U4584 ( .A(n5914), .B(n5912), .Z(n5913) );
  XOR U4585 ( .A(n5915), .B(n5916), .Z(n2997) );
  NOR U4586 ( .A(n5917), .B(n5915), .Z(n5916) );
  XOR U4587 ( .A(n5918), .B(n5919), .Z(n2994) );
  NOR U4588 ( .A(n5920), .B(n5918), .Z(n5919) );
  XOR U4589 ( .A(n5921), .B(n5922), .Z(n2992) );
  NOR U4590 ( .A(n5923), .B(n5921), .Z(n5922) );
  XOR U4591 ( .A(n5924), .B(n5925), .Z(n2993) );
  NOR U4592 ( .A(n5926), .B(n5924), .Z(n5925) );
  XOR U4593 ( .A(n5927), .B(n5928), .Z(n3091) );
  NOR U4594 ( .A(n5929), .B(n5927), .Z(n5928) );
  XOR U4595 ( .A(n5930), .B(n5931), .Z(n3095) );
  NOR U4596 ( .A(n5932), .B(n5930), .Z(n5931) );
  XOR U4597 ( .A(n5933), .B(n5934), .Z(n2982) );
  NOR U4598 ( .A(n5935), .B(n5933), .Z(n5934) );
  XOR U4599 ( .A(n5936), .B(n5937), .Z(n2983) );
  NOR U4600 ( .A(n5938), .B(n5936), .Z(n5937) );
  XOR U4601 ( .A(n5939), .B(n5940), .Z(n3103) );
  NOR U4602 ( .A(n5941), .B(n5939), .Z(n5940) );
  XOR U4603 ( .A(n5942), .B(n5943), .Z(n3104) );
  NOR U4604 ( .A(n5944), .B(n5942), .Z(n5943) );
  XOR U4605 ( .A(n5945), .B(n5946), .Z(n3105) );
  NOR U4606 ( .A(n5947), .B(n5945), .Z(n5946) );
  XOR U4607 ( .A(n5948), .B(n5949), .Z(n2976) );
  NOR U4608 ( .A(n5950), .B(n5948), .Z(n5949) );
  XOR U4609 ( .A(n5951), .B(n5952), .Z(n2970) );
  NOR U4610 ( .A(n5953), .B(n5951), .Z(n5952) );
  XOR U4611 ( .A(n5954), .B(n5955), .Z(n2967) );
  NOR U4612 ( .A(n5956), .B(n5954), .Z(n5955) );
  XOR U4613 ( .A(n5957), .B(n5958), .Z(n2965) );
  NOR U4614 ( .A(n5959), .B(n5957), .Z(n5958) );
  XOR U4615 ( .A(n5960), .B(n5961), .Z(n2966) );
  NOR U4616 ( .A(n5962), .B(n5960), .Z(n5961) );
  XOR U4617 ( .A(n5963), .B(n5964), .Z(n3124) );
  NOR U4618 ( .A(n5965), .B(n5963), .Z(n5964) );
  XOR U4619 ( .A(n5966), .B(n5967), .Z(n3128) );
  NOR U4620 ( .A(n5968), .B(n5966), .Z(n5967) );
  XOR U4621 ( .A(n5969), .B(n5970), .Z(n2955) );
  NOR U4622 ( .A(n5971), .B(n5969), .Z(n5970) );
  XOR U4623 ( .A(n5972), .B(n5973), .Z(n2956) );
  NOR U4624 ( .A(n5974), .B(n5972), .Z(n5973) );
  XOR U4625 ( .A(n5975), .B(n5976), .Z(n3136) );
  NOR U4626 ( .A(n5977), .B(n5975), .Z(n5976) );
  XOR U4627 ( .A(n5978), .B(n5979), .Z(n3137) );
  NOR U4628 ( .A(n5980), .B(n5978), .Z(n5979) );
  XOR U4629 ( .A(n5981), .B(n5982), .Z(n3138) );
  NOR U4630 ( .A(n5983), .B(n5981), .Z(n5982) );
  XOR U4631 ( .A(n5984), .B(n5985), .Z(n2949) );
  NOR U4632 ( .A(n5986), .B(n5984), .Z(n5985) );
  XOR U4633 ( .A(n5987), .B(n5988), .Z(n2943) );
  NOR U4634 ( .A(n5989), .B(n5987), .Z(n5988) );
  XOR U4635 ( .A(n5990), .B(n5991), .Z(n2940) );
  NOR U4636 ( .A(n5992), .B(n5990), .Z(n5991) );
  XOR U4637 ( .A(n5993), .B(n5994), .Z(n2938) );
  NOR U4638 ( .A(n5995), .B(n5993), .Z(n5994) );
  XOR U4639 ( .A(n5996), .B(n5997), .Z(n2939) );
  NOR U4640 ( .A(n5998), .B(n5996), .Z(n5997) );
  XOR U4641 ( .A(n5999), .B(n6000), .Z(n3157) );
  NOR U4642 ( .A(n6001), .B(n5999), .Z(n6000) );
  XOR U4643 ( .A(n6002), .B(n6003), .Z(n3161) );
  NOR U4644 ( .A(n6004), .B(n6002), .Z(n6003) );
  XOR U4645 ( .A(n6005), .B(n6006), .Z(n2928) );
  NOR U4646 ( .A(n6007), .B(n6005), .Z(n6006) );
  XOR U4647 ( .A(n6008), .B(n6009), .Z(n2929) );
  NOR U4648 ( .A(n6010), .B(n6008), .Z(n6009) );
  XOR U4649 ( .A(n6011), .B(n6012), .Z(n3169) );
  NOR U4650 ( .A(n6013), .B(n6011), .Z(n6012) );
  XOR U4651 ( .A(n6014), .B(n6015), .Z(n3170) );
  NOR U4652 ( .A(n6016), .B(n6014), .Z(n6015) );
  XOR U4653 ( .A(n6017), .B(n6018), .Z(n3171) );
  NOR U4654 ( .A(n6019), .B(n6017), .Z(n6018) );
  XOR U4655 ( .A(n6020), .B(n6021), .Z(n2922) );
  NOR U4656 ( .A(n6022), .B(n6020), .Z(n6021) );
  XOR U4657 ( .A(n6023), .B(n6024), .Z(n2916) );
  NOR U4658 ( .A(n6025), .B(n6023), .Z(n6024) );
  XOR U4659 ( .A(n6026), .B(n6027), .Z(n2913) );
  NOR U4660 ( .A(n6028), .B(n6026), .Z(n6027) );
  XOR U4661 ( .A(n6029), .B(n6030), .Z(n2911) );
  NOR U4662 ( .A(n6031), .B(n6029), .Z(n6030) );
  XOR U4663 ( .A(n6032), .B(n6033), .Z(n2912) );
  NOR U4664 ( .A(n6034), .B(n6032), .Z(n6033) );
  XOR U4665 ( .A(n6035), .B(n6036), .Z(n3190) );
  NOR U4666 ( .A(n6037), .B(n6035), .Z(n6036) );
  XOR U4667 ( .A(n6038), .B(n6039), .Z(n3194) );
  NOR U4668 ( .A(n6040), .B(n6038), .Z(n6039) );
  XOR U4669 ( .A(n6041), .B(n6042), .Z(n2901) );
  NOR U4670 ( .A(n6043), .B(n6041), .Z(n6042) );
  XOR U4671 ( .A(n6044), .B(n6045), .Z(n2902) );
  NOR U4672 ( .A(n6046), .B(n6044), .Z(n6045) );
  XOR U4673 ( .A(n6047), .B(n6048), .Z(n3202) );
  NOR U4674 ( .A(n6049), .B(n6047), .Z(n6048) );
  XOR U4675 ( .A(n6050), .B(n6051), .Z(n3203) );
  NOR U4676 ( .A(n6052), .B(n6050), .Z(n6051) );
  XOR U4677 ( .A(n6053), .B(n6054), .Z(n3204) );
  NOR U4678 ( .A(n6055), .B(n6053), .Z(n6054) );
  XOR U4679 ( .A(n6056), .B(n6057), .Z(n2895) );
  NOR U4680 ( .A(n6058), .B(n6056), .Z(n6057) );
  XOR U4681 ( .A(n6059), .B(n6060), .Z(n2889) );
  NOR U4682 ( .A(n6061), .B(n6059), .Z(n6060) );
  XOR U4683 ( .A(n6062), .B(n6063), .Z(n2886) );
  NOR U4684 ( .A(n6064), .B(n6062), .Z(n6063) );
  XOR U4685 ( .A(n6065), .B(n6066), .Z(n2884) );
  NOR U4686 ( .A(n6067), .B(n6065), .Z(n6066) );
  XOR U4687 ( .A(n6068), .B(n6069), .Z(n2885) );
  NOR U4688 ( .A(n6070), .B(n6068), .Z(n6069) );
  XOR U4689 ( .A(n6071), .B(n6072), .Z(n3223) );
  NOR U4690 ( .A(n6073), .B(n6071), .Z(n6072) );
  XOR U4691 ( .A(n6074), .B(n6075), .Z(n3227) );
  NOR U4692 ( .A(n6076), .B(n6074), .Z(n6075) );
  XOR U4693 ( .A(n6077), .B(n6078), .Z(n2874) );
  NOR U4694 ( .A(n6079), .B(n6077), .Z(n6078) );
  XOR U4695 ( .A(n6080), .B(n6081), .Z(n2875) );
  NOR U4696 ( .A(n6082), .B(n6080), .Z(n6081) );
  XOR U4697 ( .A(n6083), .B(n6084), .Z(n3235) );
  NOR U4698 ( .A(n6085), .B(n6083), .Z(n6084) );
  XOR U4699 ( .A(n6086), .B(n6087), .Z(n3236) );
  NOR U4700 ( .A(n6088), .B(n6086), .Z(n6087) );
  XOR U4701 ( .A(n6089), .B(n6090), .Z(n3237) );
  NOR U4702 ( .A(n6091), .B(n6089), .Z(n6090) );
  XOR U4703 ( .A(n6092), .B(n6093), .Z(n2868) );
  NOR U4704 ( .A(n6094), .B(n6092), .Z(n6093) );
  XOR U4705 ( .A(n6095), .B(n6096), .Z(n2862) );
  NOR U4706 ( .A(n6097), .B(n6095), .Z(n6096) );
  XOR U4707 ( .A(n6098), .B(n6099), .Z(n2859) );
  NOR U4708 ( .A(n6100), .B(n6098), .Z(n6099) );
  XOR U4709 ( .A(n6101), .B(n6102), .Z(n2857) );
  NOR U4710 ( .A(n6103), .B(n6101), .Z(n6102) );
  XOR U4711 ( .A(n6104), .B(n6105), .Z(n2858) );
  NOR U4712 ( .A(n6106), .B(n6104), .Z(n6105) );
  XOR U4713 ( .A(n6107), .B(n6108), .Z(n3256) );
  NOR U4714 ( .A(n6109), .B(n6107), .Z(n6108) );
  XOR U4715 ( .A(n6110), .B(n6111), .Z(n3260) );
  NOR U4716 ( .A(n6112), .B(n6110), .Z(n6111) );
  XOR U4717 ( .A(n6113), .B(n6114), .Z(n2847) );
  NOR U4718 ( .A(n6115), .B(n6113), .Z(n6114) );
  XOR U4719 ( .A(n6116), .B(n6117), .Z(n2848) );
  NOR U4720 ( .A(n6118), .B(n6116), .Z(n6117) );
  XOR U4721 ( .A(n6119), .B(n6120), .Z(n3268) );
  NOR U4722 ( .A(n6121), .B(n6119), .Z(n6120) );
  XOR U4723 ( .A(n6122), .B(n6123), .Z(n3269) );
  NOR U4724 ( .A(n6124), .B(n6122), .Z(n6123) );
  XOR U4725 ( .A(n6125), .B(n6126), .Z(n3270) );
  NOR U4726 ( .A(n6127), .B(n6125), .Z(n6126) );
  XOR U4727 ( .A(n6128), .B(n6129), .Z(n2841) );
  NOR U4728 ( .A(n6130), .B(n6128), .Z(n6129) );
  XOR U4729 ( .A(n6131), .B(n6132), .Z(n2835) );
  NOR U4730 ( .A(n6133), .B(n6131), .Z(n6132) );
  XOR U4731 ( .A(n6134), .B(n6135), .Z(n2832) );
  NOR U4732 ( .A(n6136), .B(n6134), .Z(n6135) );
  XOR U4733 ( .A(n6137), .B(n6138), .Z(n2830) );
  NOR U4734 ( .A(n6139), .B(n6137), .Z(n6138) );
  XOR U4735 ( .A(n6140), .B(n6141), .Z(n2831) );
  NOR U4736 ( .A(n6142), .B(n6140), .Z(n6141) );
  XOR U4737 ( .A(n6143), .B(n6144), .Z(n3289) );
  NOR U4738 ( .A(n6145), .B(n6143), .Z(n6144) );
  XOR U4739 ( .A(n6146), .B(n6147), .Z(n3293) );
  NOR U4740 ( .A(n6148), .B(n6146), .Z(n6147) );
  XOR U4741 ( .A(n6149), .B(n6150), .Z(n2820) );
  NOR U4742 ( .A(n6151), .B(n6149), .Z(n6150) );
  XOR U4743 ( .A(n6152), .B(n6153), .Z(n2821) );
  NOR U4744 ( .A(n6154), .B(n6152), .Z(n6153) );
  XOR U4745 ( .A(n6155), .B(n6156), .Z(n3301) );
  NOR U4746 ( .A(n6157), .B(n6155), .Z(n6156) );
  XOR U4747 ( .A(n6158), .B(n6159), .Z(n3302) );
  NOR U4748 ( .A(n6160), .B(n6158), .Z(n6159) );
  XOR U4749 ( .A(n6161), .B(n6162), .Z(n3303) );
  NOR U4750 ( .A(n6163), .B(n6161), .Z(n6162) );
  XOR U4751 ( .A(n6164), .B(n6165), .Z(n2814) );
  NOR U4752 ( .A(n6166), .B(n6164), .Z(n6165) );
  XOR U4753 ( .A(n6167), .B(n6168), .Z(n2808) );
  NOR U4754 ( .A(n6169), .B(n6167), .Z(n6168) );
  XOR U4755 ( .A(n6170), .B(n6171), .Z(n2805) );
  NOR U4756 ( .A(n6172), .B(n6170), .Z(n6171) );
  XOR U4757 ( .A(n6173), .B(n6174), .Z(n2803) );
  NOR U4758 ( .A(n6175), .B(n6173), .Z(n6174) );
  XOR U4759 ( .A(n6176), .B(n6177), .Z(n2804) );
  NOR U4760 ( .A(n6178), .B(n6176), .Z(n6177) );
  XOR U4761 ( .A(n6179), .B(n6180), .Z(n3322) );
  NOR U4762 ( .A(n6181), .B(n6179), .Z(n6180) );
  XOR U4763 ( .A(n6182), .B(n6183), .Z(n3326) );
  NOR U4764 ( .A(n6184), .B(n6182), .Z(n6183) );
  XOR U4765 ( .A(n6185), .B(n6186), .Z(n2793) );
  NOR U4766 ( .A(n6187), .B(n6185), .Z(n6186) );
  XOR U4767 ( .A(n6188), .B(n6189), .Z(n2794) );
  NOR U4768 ( .A(n6190), .B(n6188), .Z(n6189) );
  XOR U4769 ( .A(n6191), .B(n6192), .Z(n3334) );
  NOR U4770 ( .A(n6193), .B(n6191), .Z(n6192) );
  XOR U4771 ( .A(n6194), .B(n6195), .Z(n3335) );
  NOR U4772 ( .A(n6196), .B(n6194), .Z(n6195) );
  XOR U4773 ( .A(n6197), .B(n6198), .Z(n3336) );
  NOR U4774 ( .A(n6199), .B(n6197), .Z(n6198) );
  XOR U4775 ( .A(n6200), .B(n6201), .Z(n2787) );
  NOR U4776 ( .A(n6202), .B(n6200), .Z(n6201) );
  XOR U4777 ( .A(n6203), .B(n6204), .Z(n2781) );
  NOR U4778 ( .A(n6205), .B(n6203), .Z(n6204) );
  XOR U4779 ( .A(n6206), .B(n6207), .Z(n2778) );
  NOR U4780 ( .A(n6208), .B(n6206), .Z(n6207) );
  XOR U4781 ( .A(n6209), .B(n6210), .Z(n2776) );
  NOR U4782 ( .A(n6211), .B(n6209), .Z(n6210) );
  XOR U4783 ( .A(n6212), .B(n6213), .Z(n2777) );
  NOR U4784 ( .A(n6214), .B(n6212), .Z(n6213) );
  XOR U4785 ( .A(n6215), .B(n6216), .Z(n3355) );
  NOR U4786 ( .A(n6217), .B(n6215), .Z(n6216) );
  XOR U4787 ( .A(n6218), .B(n6219), .Z(n3359) );
  NOR U4788 ( .A(n6220), .B(n6218), .Z(n6219) );
  XOR U4789 ( .A(n6221), .B(n6222), .Z(n2766) );
  NOR U4790 ( .A(n6223), .B(n6221), .Z(n6222) );
  XOR U4791 ( .A(n6224), .B(n6225), .Z(n2767) );
  NOR U4792 ( .A(n6226), .B(n6224), .Z(n6225) );
  XOR U4793 ( .A(n6227), .B(n6228), .Z(n3367) );
  NOR U4794 ( .A(n6229), .B(n6227), .Z(n6228) );
  XOR U4795 ( .A(n6230), .B(n6231), .Z(n3368) );
  NOR U4796 ( .A(n6232), .B(n6230), .Z(n6231) );
  XOR U4797 ( .A(n6233), .B(n6234), .Z(n3369) );
  NOR U4798 ( .A(n6235), .B(n6233), .Z(n6234) );
  XOR U4799 ( .A(n6236), .B(n6237), .Z(n2760) );
  NOR U4800 ( .A(n6238), .B(n6236), .Z(n6237) );
  XOR U4801 ( .A(n6239), .B(n6240), .Z(n2753) );
  NOR U4802 ( .A(n6241), .B(n6239), .Z(n6240) );
  XOR U4803 ( .A(n6242), .B(n6243), .Z(n2749) );
  NOR U4804 ( .A(n6244), .B(n6242), .Z(n6243) );
  XOR U4805 ( .A(n6245), .B(n6246), .Z(n2751) );
  NOR U4806 ( .A(n6247), .B(n6245), .Z(n6246) );
  XOR U4807 ( .A(n6248), .B(n6249), .Z(n3383) );
  NOR U4808 ( .A(n6250), .B(n6248), .Z(n6249) );
  XOR U4809 ( .A(n6251), .B(n6252), .Z(n3384) );
  NOR U4810 ( .A(n6253), .B(n6251), .Z(n6252) );
  XOR U4811 ( .A(n6254), .B(n6255), .Z(n3387) );
  NOR U4812 ( .A(n6256), .B(n6254), .Z(n6255) );
  XOR U4813 ( .A(n6257), .B(n6258), .Z(n3390) );
  NOR U4814 ( .A(n6259), .B(n6257), .Z(n6258) );
  XOR U4815 ( .A(n6260), .B(n6261), .Z(n3393) );
  NOR U4816 ( .A(n6262), .B(n6260), .Z(n6261) );
  XOR U4817 ( .A(n6263), .B(n6264), .Z(n3396) );
  NOR U4818 ( .A(n6265), .B(n6263), .Z(n6264) );
  XOR U4819 ( .A(n6266), .B(n6267), .Z(n3399) );
  NOR U4820 ( .A(n6268), .B(n6266), .Z(n6267) );
  XOR U4821 ( .A(n6269), .B(n6270), .Z(n3402) );
  NOR U4822 ( .A(n6271), .B(n6269), .Z(n6270) );
  XOR U4823 ( .A(n6272), .B(n6273), .Z(n3405) );
  NOR U4824 ( .A(n6274), .B(n6272), .Z(n6273) );
  XOR U4825 ( .A(n6275), .B(n6276), .Z(n3408) );
  NOR U4826 ( .A(n6277), .B(n6275), .Z(n6276) );
  XOR U4827 ( .A(n6278), .B(n6279), .Z(n3411) );
  NOR U4828 ( .A(n6280), .B(n6278), .Z(n6279) );
  XOR U4829 ( .A(n6281), .B(n6282), .Z(n3414) );
  NOR U4830 ( .A(n6283), .B(n6281), .Z(n6282) );
  XOR U4831 ( .A(n6284), .B(n6285), .Z(n3417) );
  NOR U4832 ( .A(n6286), .B(n6284), .Z(n6285) );
  XOR U4833 ( .A(n6287), .B(n6288), .Z(n3420) );
  NOR U4834 ( .A(n6289), .B(n6287), .Z(n6288) );
  XOR U4835 ( .A(n6290), .B(n6291), .Z(n3423) );
  NOR U4836 ( .A(n6292), .B(n6290), .Z(n6291) );
  XOR U4837 ( .A(n6293), .B(n6294), .Z(n3426) );
  NOR U4838 ( .A(n6295), .B(n6293), .Z(n6294) );
  XOR U4839 ( .A(n6296), .B(n6297), .Z(n3429) );
  NOR U4840 ( .A(n6298), .B(n6296), .Z(n6297) );
  XOR U4841 ( .A(n6299), .B(n6300), .Z(n3432) );
  NOR U4842 ( .A(n6301), .B(n6299), .Z(n6300) );
  XOR U4843 ( .A(n6302), .B(n6303), .Z(n3435) );
  NOR U4844 ( .A(n6304), .B(n6302), .Z(n6303) );
  XOR U4845 ( .A(n6305), .B(n6306), .Z(n3438) );
  NOR U4846 ( .A(n6307), .B(n6305), .Z(n6306) );
  XOR U4847 ( .A(n6308), .B(n6309), .Z(n3441) );
  NOR U4848 ( .A(n6310), .B(n6308), .Z(n6309) );
  XOR U4849 ( .A(n6311), .B(n6312), .Z(n3444) );
  NOR U4850 ( .A(n6313), .B(n6311), .Z(n6312) );
  XOR U4851 ( .A(n6314), .B(n6315), .Z(n3447) );
  NOR U4852 ( .A(n6316), .B(n6314), .Z(n6315) );
  XOR U4853 ( .A(n6317), .B(n6318), .Z(n3450) );
  NOR U4854 ( .A(n6319), .B(n6317), .Z(n6318) );
  XOR U4855 ( .A(n6320), .B(n6321), .Z(n3453) );
  NOR U4856 ( .A(n6322), .B(n6320), .Z(n6321) );
  XOR U4857 ( .A(n6323), .B(n6324), .Z(n3456) );
  NOR U4858 ( .A(n6325), .B(n6323), .Z(n6324) );
  XOR U4859 ( .A(n6326), .B(n6327), .Z(n3459) );
  NOR U4860 ( .A(n6328), .B(n6326), .Z(n6327) );
  XOR U4861 ( .A(n6329), .B(n6330), .Z(n3462) );
  NOR U4862 ( .A(n6331), .B(n6329), .Z(n6330) );
  XOR U4863 ( .A(n6332), .B(n6333), .Z(n3465) );
  NOR U4864 ( .A(n6334), .B(n6332), .Z(n6333) );
  XOR U4865 ( .A(n6335), .B(n6336), .Z(n3468) );
  NOR U4866 ( .A(n6337), .B(n6335), .Z(n6336) );
  XOR U4867 ( .A(n6338), .B(n6339), .Z(n3471) );
  NOR U4868 ( .A(n6340), .B(n6338), .Z(n6339) );
  XOR U4869 ( .A(n6341), .B(n6342), .Z(n3474) );
  NOR U4870 ( .A(n6343), .B(n6341), .Z(n6342) );
  XOR U4871 ( .A(n6344), .B(n6345), .Z(n3477) );
  NOR U4872 ( .A(n6346), .B(n6344), .Z(n6345) );
  XOR U4873 ( .A(n6347), .B(n6348), .Z(n3480) );
  NOR U4874 ( .A(n6349), .B(n6347), .Z(n6348) );
  XOR U4875 ( .A(n6350), .B(n6351), .Z(n3483) );
  NOR U4876 ( .A(n6352), .B(n6350), .Z(n6351) );
  XOR U4877 ( .A(n6353), .B(n6354), .Z(n3486) );
  NOR U4878 ( .A(n6355), .B(n6353), .Z(n6354) );
  XOR U4879 ( .A(n6356), .B(n6357), .Z(n3489) );
  NOR U4880 ( .A(n6358), .B(n6356), .Z(n6357) );
  XOR U4881 ( .A(n6359), .B(n6360), .Z(n3492) );
  NOR U4882 ( .A(n6361), .B(n6359), .Z(n6360) );
  XOR U4883 ( .A(n6362), .B(n6363), .Z(n3495) );
  NOR U4884 ( .A(n6364), .B(n6362), .Z(n6363) );
  XOR U4885 ( .A(n6365), .B(n6366), .Z(n3498) );
  NOR U4886 ( .A(n6367), .B(n6365), .Z(n6366) );
  XOR U4887 ( .A(n6368), .B(n6369), .Z(n3501) );
  NOR U4888 ( .A(n6370), .B(n6368), .Z(n6369) );
  XOR U4889 ( .A(n6371), .B(n6372), .Z(n3504) );
  NOR U4890 ( .A(n6373), .B(n6371), .Z(n6372) );
  XOR U4891 ( .A(n6374), .B(n6375), .Z(n3507) );
  NOR U4892 ( .A(n6376), .B(n6374), .Z(n6375) );
  XOR U4893 ( .A(n6377), .B(n6378), .Z(n3510) );
  NOR U4894 ( .A(n6379), .B(n6377), .Z(n6378) );
  XOR U4895 ( .A(n6380), .B(n6381), .Z(n3513) );
  NOR U4896 ( .A(n6382), .B(n6380), .Z(n6381) );
  XOR U4897 ( .A(n6383), .B(n6384), .Z(n3516) );
  NOR U4898 ( .A(n6385), .B(n6383), .Z(n6384) );
  XOR U4899 ( .A(n6386), .B(n6387), .Z(n3519) );
  NOR U4900 ( .A(n6388), .B(n6386), .Z(n6387) );
  XOR U4901 ( .A(n6389), .B(n6390), .Z(n3522) );
  NOR U4902 ( .A(n6391), .B(n6389), .Z(n6390) );
  XOR U4903 ( .A(n6392), .B(n6393), .Z(n3525) );
  NOR U4904 ( .A(n6394), .B(n6392), .Z(n6393) );
  XOR U4905 ( .A(n6395), .B(n6396), .Z(n3528) );
  NOR U4906 ( .A(n6397), .B(n6395), .Z(n6396) );
  XOR U4907 ( .A(n6398), .B(n6399), .Z(n3531) );
  NOR U4908 ( .A(n6400), .B(n6398), .Z(n6399) );
  XOR U4909 ( .A(n6401), .B(n6402), .Z(n3534) );
  NOR U4910 ( .A(n6403), .B(n6401), .Z(n6402) );
  XOR U4911 ( .A(n6404), .B(n6405), .Z(n3537) );
  NOR U4912 ( .A(n6406), .B(n6404), .Z(n6405) );
  XOR U4913 ( .A(n6407), .B(n6408), .Z(n3540) );
  NOR U4914 ( .A(n6409), .B(n6407), .Z(n6408) );
  XOR U4915 ( .A(n6410), .B(n6411), .Z(n3543) );
  NOR U4916 ( .A(n6412), .B(n6410), .Z(n6411) );
  XOR U4917 ( .A(n6413), .B(n6414), .Z(n3546) );
  NOR U4918 ( .A(n6415), .B(n6413), .Z(n6414) );
  XOR U4919 ( .A(n6416), .B(n6417), .Z(n3549) );
  NOR U4920 ( .A(n6418), .B(n6416), .Z(n6417) );
  XOR U4921 ( .A(n6419), .B(n6420), .Z(n3552) );
  NOR U4922 ( .A(n6421), .B(n6419), .Z(n6420) );
  XOR U4923 ( .A(n6422), .B(n6423), .Z(n3555) );
  NOR U4924 ( .A(n6424), .B(n6422), .Z(n6423) );
  XOR U4925 ( .A(n6425), .B(n6426), .Z(n3558) );
  NOR U4926 ( .A(n6427), .B(n6425), .Z(n6426) );
  XOR U4927 ( .A(n6428), .B(n6429), .Z(n3561) );
  NOR U4928 ( .A(n6430), .B(n6428), .Z(n6429) );
  XOR U4929 ( .A(n6431), .B(n6432), .Z(n3564) );
  NOR U4930 ( .A(n6433), .B(n6431), .Z(n6432) );
  XOR U4931 ( .A(n6434), .B(n6435), .Z(n3567) );
  NOR U4932 ( .A(n6436), .B(n6434), .Z(n6435) );
  XOR U4933 ( .A(n6437), .B(n6438), .Z(n3570) );
  NOR U4934 ( .A(n6439), .B(n6437), .Z(n6438) );
  XOR U4935 ( .A(n6440), .B(n6441), .Z(n3573) );
  NOR U4936 ( .A(n6442), .B(n6440), .Z(n6441) );
  XOR U4937 ( .A(n6443), .B(n6444), .Z(n3576) );
  NOR U4938 ( .A(n6445), .B(n6443), .Z(n6444) );
  XOR U4939 ( .A(n6446), .B(n6447), .Z(n3579) );
  NOR U4940 ( .A(n6448), .B(n6446), .Z(n6447) );
  XOR U4941 ( .A(n6449), .B(n6450), .Z(n3582) );
  NOR U4942 ( .A(n6451), .B(n6449), .Z(n6450) );
  XOR U4943 ( .A(n6452), .B(n6453), .Z(n3585) );
  NOR U4944 ( .A(n6454), .B(n6452), .Z(n6453) );
  XOR U4945 ( .A(n6455), .B(n6456), .Z(n3588) );
  NOR U4946 ( .A(n6457), .B(n6455), .Z(n6456) );
  XOR U4947 ( .A(n6458), .B(n6459), .Z(n3591) );
  NOR U4948 ( .A(n6460), .B(n6458), .Z(n6459) );
  XOR U4949 ( .A(n6461), .B(n6462), .Z(n3594) );
  NOR U4950 ( .A(n6463), .B(n6461), .Z(n6462) );
  XOR U4951 ( .A(n6464), .B(n6465), .Z(n3597) );
  NOR U4952 ( .A(n6466), .B(n6464), .Z(n6465) );
  XOR U4953 ( .A(n6467), .B(n6468), .Z(n3600) );
  NOR U4954 ( .A(n6469), .B(n6467), .Z(n6468) );
  XOR U4955 ( .A(n6470), .B(n6471), .Z(n3603) );
  NOR U4956 ( .A(n6472), .B(n6470), .Z(n6471) );
  XOR U4957 ( .A(n6473), .B(n6474), .Z(n3606) );
  NOR U4958 ( .A(n6475), .B(n6473), .Z(n6474) );
  XOR U4959 ( .A(n6476), .B(n6477), .Z(n3609) );
  NOR U4960 ( .A(n6478), .B(n6476), .Z(n6477) );
  XOR U4961 ( .A(n6479), .B(n6480), .Z(n3612) );
  NOR U4962 ( .A(n6481), .B(n6479), .Z(n6480) );
  XOR U4963 ( .A(n6482), .B(n6483), .Z(n3615) );
  NOR U4964 ( .A(n6484), .B(n6482), .Z(n6483) );
  XOR U4965 ( .A(n6485), .B(n6486), .Z(n3618) );
  NOR U4966 ( .A(n6487), .B(n6485), .Z(n6486) );
  XOR U4967 ( .A(n6488), .B(n6489), .Z(n3621) );
  NOR U4968 ( .A(n6490), .B(n6488), .Z(n6489) );
  XOR U4969 ( .A(n6491), .B(n6492), .Z(n3624) );
  NOR U4970 ( .A(n6493), .B(n6491), .Z(n6492) );
  XOR U4971 ( .A(n6494), .B(n6495), .Z(n3627) );
  NOR U4972 ( .A(n6496), .B(n6494), .Z(n6495) );
  XOR U4973 ( .A(n6497), .B(n6498), .Z(n3630) );
  NOR U4974 ( .A(n6499), .B(n6497), .Z(n6498) );
  XOR U4975 ( .A(n6500), .B(n6501), .Z(n3633) );
  NOR U4976 ( .A(n6502), .B(n6500), .Z(n6501) );
  XOR U4977 ( .A(n6503), .B(n6504), .Z(n3636) );
  NOR U4978 ( .A(n6505), .B(n6503), .Z(n6504) );
  XOR U4979 ( .A(n6506), .B(n6507), .Z(n3639) );
  NOR U4980 ( .A(n6508), .B(n6506), .Z(n6507) );
  XOR U4981 ( .A(n6509), .B(n6510), .Z(n3642) );
  NOR U4982 ( .A(n6511), .B(n6509), .Z(n6510) );
  XOR U4983 ( .A(n6512), .B(n6513), .Z(n3645) );
  NOR U4984 ( .A(n6514), .B(n6512), .Z(n6513) );
  XOR U4985 ( .A(n6515), .B(n6516), .Z(n3648) );
  NOR U4986 ( .A(n6517), .B(n6515), .Z(n6516) );
  XOR U4987 ( .A(n6518), .B(n6519), .Z(n3651) );
  NOR U4988 ( .A(n6520), .B(n6518), .Z(n6519) );
  XOR U4989 ( .A(n6521), .B(n6522), .Z(n3654) );
  NOR U4990 ( .A(n6523), .B(n6521), .Z(n6522) );
  XOR U4991 ( .A(n6524), .B(n6525), .Z(n3657) );
  NOR U4992 ( .A(n6526), .B(n6524), .Z(n6525) );
  XOR U4993 ( .A(n6527), .B(n6528), .Z(n3660) );
  NOR U4994 ( .A(n6529), .B(n6527), .Z(n6528) );
  XOR U4995 ( .A(n6530), .B(n6531), .Z(n3663) );
  NOR U4996 ( .A(n6532), .B(n6530), .Z(n6531) );
  XOR U4997 ( .A(n6533), .B(n6534), .Z(n3666) );
  NOR U4998 ( .A(n6535), .B(n6533), .Z(n6534) );
  XOR U4999 ( .A(n6536), .B(n6537), .Z(n3669) );
  NOR U5000 ( .A(n6538), .B(n6536), .Z(n6537) );
  XOR U5001 ( .A(n6539), .B(n6540), .Z(n3672) );
  NOR U5002 ( .A(n6541), .B(n6539), .Z(n6540) );
  XOR U5003 ( .A(n6542), .B(n6543), .Z(n3675) );
  NOR U5004 ( .A(n6544), .B(n6542), .Z(n6543) );
  XOR U5005 ( .A(n6545), .B(n6546), .Z(n3678) );
  NOR U5006 ( .A(n6547), .B(n6545), .Z(n6546) );
  XOR U5007 ( .A(n6548), .B(n6549), .Z(n3681) );
  NOR U5008 ( .A(n6550), .B(n6548), .Z(n6549) );
  XOR U5009 ( .A(n6551), .B(n6552), .Z(n3684) );
  NOR U5010 ( .A(n6553), .B(n6551), .Z(n6552) );
  XOR U5011 ( .A(n6554), .B(n6555), .Z(n3687) );
  NOR U5012 ( .A(n6556), .B(n6554), .Z(n6555) );
  XOR U5013 ( .A(n6557), .B(n6558), .Z(n3690) );
  NOR U5014 ( .A(n6559), .B(n6557), .Z(n6558) );
  XOR U5015 ( .A(n6560), .B(n6561), .Z(n3693) );
  NOR U5016 ( .A(n6562), .B(n6560), .Z(n6561) );
  XOR U5017 ( .A(n6563), .B(n6564), .Z(n3696) );
  NOR U5018 ( .A(n6565), .B(n6563), .Z(n6564) );
  XOR U5019 ( .A(n6566), .B(n6567), .Z(n3699) );
  NOR U5020 ( .A(n6568), .B(n6566), .Z(n6567) );
  XOR U5021 ( .A(n6569), .B(n6570), .Z(n3702) );
  NOR U5022 ( .A(n6571), .B(n6569), .Z(n6570) );
  XOR U5023 ( .A(n6572), .B(n6573), .Z(n3705) );
  NOR U5024 ( .A(n6574), .B(n6572), .Z(n6573) );
  XOR U5025 ( .A(n6575), .B(n6576), .Z(n3708) );
  NOR U5026 ( .A(n6577), .B(n6575), .Z(n6576) );
  XOR U5027 ( .A(n6578), .B(n6579), .Z(n3711) );
  NOR U5028 ( .A(n6580), .B(n6578), .Z(n6579) );
  XOR U5029 ( .A(n6581), .B(n6582), .Z(n3714) );
  NOR U5030 ( .A(n6583), .B(n6581), .Z(n6582) );
  XOR U5031 ( .A(n6584), .B(n6585), .Z(n3717) );
  NOR U5032 ( .A(n6586), .B(n6584), .Z(n6585) );
  XOR U5033 ( .A(n6587), .B(n6588), .Z(n3720) );
  NOR U5034 ( .A(n6589), .B(n6587), .Z(n6588) );
  XOR U5035 ( .A(n6590), .B(n6591), .Z(n3723) );
  NOR U5036 ( .A(n6592), .B(n6590), .Z(n6591) );
  XOR U5037 ( .A(n6593), .B(n6594), .Z(n3726) );
  NOR U5038 ( .A(n6595), .B(n6593), .Z(n6594) );
  XOR U5039 ( .A(n6596), .B(n6597), .Z(n3729) );
  NOR U5040 ( .A(n6598), .B(n6596), .Z(n6597) );
  XOR U5041 ( .A(n6599), .B(n6600), .Z(n3732) );
  NOR U5042 ( .A(n6601), .B(n6599), .Z(n6600) );
  XOR U5043 ( .A(n6602), .B(n6603), .Z(n3735) );
  NOR U5044 ( .A(n6604), .B(n6602), .Z(n6603) );
  XOR U5045 ( .A(n6605), .B(n6606), .Z(n3738) );
  NOR U5046 ( .A(n6607), .B(n6605), .Z(n6606) );
  XOR U5047 ( .A(n6608), .B(n6609), .Z(n3741) );
  NOR U5048 ( .A(n6610), .B(n6608), .Z(n6609) );
  XOR U5049 ( .A(n6611), .B(n6612), .Z(n3744) );
  NOR U5050 ( .A(n6613), .B(n6611), .Z(n6612) );
  XOR U5051 ( .A(n6614), .B(n6615), .Z(n3747) );
  NOR U5052 ( .A(n6616), .B(n6614), .Z(n6615) );
  XOR U5053 ( .A(n6617), .B(n6618), .Z(n3750) );
  NOR U5054 ( .A(n6619), .B(n6617), .Z(n6618) );
  XOR U5055 ( .A(n6620), .B(n6621), .Z(n3753) );
  NOR U5056 ( .A(n6622), .B(n6620), .Z(n6621) );
  XOR U5057 ( .A(n6623), .B(n6624), .Z(n3756) );
  NOR U5058 ( .A(n6625), .B(n6623), .Z(n6624) );
  XOR U5059 ( .A(n6626), .B(n6627), .Z(n3759) );
  NOR U5060 ( .A(n6628), .B(n6626), .Z(n6627) );
  XOR U5061 ( .A(n6629), .B(n6630), .Z(n3762) );
  NOR U5062 ( .A(n6631), .B(n6629), .Z(n6630) );
  XOR U5063 ( .A(n6632), .B(n6633), .Z(n3765) );
  NOR U5064 ( .A(n6634), .B(n6632), .Z(n6633) );
  XOR U5065 ( .A(n6635), .B(n6636), .Z(n3768) );
  NOR U5066 ( .A(n6637), .B(n6635), .Z(n6636) );
  XOR U5067 ( .A(n6638), .B(n6639), .Z(n3771) );
  NOR U5068 ( .A(n6640), .B(n6638), .Z(n6639) );
  XOR U5069 ( .A(n6641), .B(n6642), .Z(n3774) );
  NOR U5070 ( .A(n6643), .B(n6641), .Z(n6642) );
  XOR U5071 ( .A(n6644), .B(n6645), .Z(n3777) );
  NOR U5072 ( .A(n6646), .B(n6644), .Z(n6645) );
  XOR U5073 ( .A(n6647), .B(n6648), .Z(n3780) );
  NOR U5074 ( .A(n6649), .B(n6647), .Z(n6648) );
  XOR U5075 ( .A(n6650), .B(n6651), .Z(n3783) );
  NOR U5076 ( .A(n6652), .B(n6650), .Z(n6651) );
  XOR U5077 ( .A(n6653), .B(n6654), .Z(n3786) );
  NOR U5078 ( .A(n6655), .B(n6653), .Z(n6654) );
  XOR U5079 ( .A(n6656), .B(n6657), .Z(n3789) );
  NOR U5080 ( .A(n6658), .B(n6656), .Z(n6657) );
  XOR U5081 ( .A(n6659), .B(n6660), .Z(n3792) );
  NOR U5082 ( .A(n6661), .B(n6659), .Z(n6660) );
  XOR U5083 ( .A(n6662), .B(n6663), .Z(n3795) );
  NOR U5084 ( .A(n6664), .B(n6662), .Z(n6663) );
  XOR U5085 ( .A(n6665), .B(n6666), .Z(n3798) );
  NOR U5086 ( .A(n6667), .B(n6665), .Z(n6666) );
  XOR U5087 ( .A(n6668), .B(n6669), .Z(n3801) );
  NOR U5088 ( .A(n6670), .B(n6668), .Z(n6669) );
  XOR U5089 ( .A(n6671), .B(n6672), .Z(n3804) );
  NOR U5090 ( .A(n6673), .B(n6671), .Z(n6672) );
  XOR U5091 ( .A(n6674), .B(n6675), .Z(n3807) );
  NOR U5092 ( .A(n6676), .B(n6674), .Z(n6675) );
  XOR U5093 ( .A(n6677), .B(n6678), .Z(n3810) );
  NOR U5094 ( .A(n6679), .B(n6677), .Z(n6678) );
  XOR U5095 ( .A(n6680), .B(n6681), .Z(n3813) );
  NOR U5096 ( .A(n6682), .B(n6680), .Z(n6681) );
  XOR U5097 ( .A(n6683), .B(n6684), .Z(n3816) );
  NOR U5098 ( .A(n6685), .B(n6683), .Z(n6684) );
  XOR U5099 ( .A(n6686), .B(n6687), .Z(n3819) );
  NOR U5100 ( .A(n6688), .B(n6686), .Z(n6687) );
  XOR U5101 ( .A(n6689), .B(n6690), .Z(n3822) );
  NOR U5102 ( .A(n6691), .B(n6689), .Z(n6690) );
  XOR U5103 ( .A(n6692), .B(n6693), .Z(n3825) );
  NOR U5104 ( .A(n6694), .B(n6692), .Z(n6693) );
  XOR U5105 ( .A(n6695), .B(n6696), .Z(n3828) );
  NOR U5106 ( .A(n6697), .B(n6695), .Z(n6696) );
  XOR U5107 ( .A(n6698), .B(n6699), .Z(n3831) );
  NOR U5108 ( .A(n6700), .B(n6698), .Z(n6699) );
  XOR U5109 ( .A(n6701), .B(n6702), .Z(n3834) );
  NOR U5110 ( .A(n6703), .B(n6701), .Z(n6702) );
  XOR U5111 ( .A(n6704), .B(n6705), .Z(n3837) );
  NOR U5112 ( .A(n6706), .B(n6704), .Z(n6705) );
  XOR U5113 ( .A(n6707), .B(n6708), .Z(n3840) );
  NOR U5114 ( .A(n6709), .B(n6707), .Z(n6708) );
  XOR U5115 ( .A(n6710), .B(n6711), .Z(n3843) );
  NOR U5116 ( .A(n6712), .B(n6710), .Z(n6711) );
  XOR U5117 ( .A(n6713), .B(n6714), .Z(n3846) );
  NOR U5118 ( .A(n6715), .B(n6713), .Z(n6714) );
  XOR U5119 ( .A(n6716), .B(n6717), .Z(n3849) );
  NOR U5120 ( .A(n6718), .B(n6716), .Z(n6717) );
  XOR U5121 ( .A(n6719), .B(n6720), .Z(n3852) );
  NOR U5122 ( .A(n6721), .B(n6719), .Z(n6720) );
  XOR U5123 ( .A(n6722), .B(n6723), .Z(n3855) );
  NOR U5124 ( .A(n6724), .B(n6722), .Z(n6723) );
  XOR U5125 ( .A(n6725), .B(n6726), .Z(n3858) );
  NOR U5126 ( .A(n6727), .B(n6725), .Z(n6726) );
  XOR U5127 ( .A(n6728), .B(n6729), .Z(n3861) );
  NOR U5128 ( .A(n6730), .B(n6728), .Z(n6729) );
  XOR U5129 ( .A(n6731), .B(n6732), .Z(n3864) );
  NOR U5130 ( .A(n6733), .B(n6731), .Z(n6732) );
  XOR U5131 ( .A(n6734), .B(n6735), .Z(n3867) );
  NOR U5132 ( .A(n6736), .B(n6734), .Z(n6735) );
  XOR U5133 ( .A(n6737), .B(n6738), .Z(n3870) );
  NOR U5134 ( .A(n6739), .B(n6737), .Z(n6738) );
  XOR U5135 ( .A(n6740), .B(n6741), .Z(n3873) );
  NOR U5136 ( .A(n6742), .B(n6740), .Z(n6741) );
  XOR U5137 ( .A(n6743), .B(n6744), .Z(n3876) );
  NOR U5138 ( .A(n6745), .B(n6743), .Z(n6744) );
  XOR U5139 ( .A(n6746), .B(n6747), .Z(n3879) );
  NOR U5140 ( .A(n6748), .B(n6746), .Z(n6747) );
  XOR U5141 ( .A(n6749), .B(n6750), .Z(n3882) );
  NOR U5142 ( .A(n6751), .B(n6749), .Z(n6750) );
  XOR U5143 ( .A(n6752), .B(n6753), .Z(n3885) );
  NOR U5144 ( .A(n6754), .B(n6752), .Z(n6753) );
  XOR U5145 ( .A(n6755), .B(n6756), .Z(n3888) );
  NOR U5146 ( .A(n6757), .B(n6755), .Z(n6756) );
  XOR U5147 ( .A(n6758), .B(n6759), .Z(n3891) );
  NOR U5148 ( .A(n6760), .B(n6758), .Z(n6759) );
  XOR U5149 ( .A(n6761), .B(n6762), .Z(n3894) );
  NOR U5150 ( .A(n6763), .B(n6761), .Z(n6762) );
  XOR U5151 ( .A(n6764), .B(n6765), .Z(n3897) );
  NOR U5152 ( .A(n6766), .B(n6764), .Z(n6765) );
  XOR U5153 ( .A(n6767), .B(n6768), .Z(n3900) );
  NOR U5154 ( .A(n6769), .B(n6767), .Z(n6768) );
  XOR U5155 ( .A(n6770), .B(n6771), .Z(n3903) );
  NOR U5156 ( .A(n6772), .B(n6770), .Z(n6771) );
  XOR U5157 ( .A(n6773), .B(n6774), .Z(n3906) );
  NOR U5158 ( .A(n6775), .B(n6773), .Z(n6774) );
  XOR U5159 ( .A(n6776), .B(n6777), .Z(n3909) );
  NOR U5160 ( .A(n6778), .B(n6776), .Z(n6777) );
  XOR U5161 ( .A(n6779), .B(n6780), .Z(n3912) );
  NOR U5162 ( .A(n6781), .B(n6779), .Z(n6780) );
  XOR U5163 ( .A(n6782), .B(n6783), .Z(n3915) );
  NOR U5164 ( .A(n6784), .B(n6782), .Z(n6783) );
  XOR U5165 ( .A(n6785), .B(n6786), .Z(n3918) );
  NOR U5166 ( .A(n6787), .B(n6785), .Z(n6786) );
  XOR U5167 ( .A(n6788), .B(n6789), .Z(n3921) );
  NOR U5168 ( .A(n6790), .B(n6788), .Z(n6789) );
  XOR U5169 ( .A(n6791), .B(n6792), .Z(n3924) );
  NOR U5170 ( .A(n6793), .B(n6791), .Z(n6792) );
  XOR U5171 ( .A(n6794), .B(n6795), .Z(n3927) );
  NOR U5172 ( .A(n6796), .B(n6794), .Z(n6795) );
  XOR U5173 ( .A(n6797), .B(n6798), .Z(n3930) );
  NOR U5174 ( .A(n6799), .B(n6797), .Z(n6798) );
  XOR U5175 ( .A(n6800), .B(n6801), .Z(n3933) );
  NOR U5176 ( .A(n6802), .B(n6800), .Z(n6801) );
  XOR U5177 ( .A(n6803), .B(n6804), .Z(n3936) );
  NOR U5178 ( .A(n6805), .B(n6803), .Z(n6804) );
  XOR U5179 ( .A(n6806), .B(n6807), .Z(n3939) );
  NOR U5180 ( .A(n6808), .B(n6806), .Z(n6807) );
  XOR U5181 ( .A(n6809), .B(n6810), .Z(n3942) );
  NOR U5182 ( .A(n6811), .B(n6809), .Z(n6810) );
  XOR U5183 ( .A(n6812), .B(n6813), .Z(n3945) );
  NOR U5184 ( .A(n6814), .B(n6812), .Z(n6813) );
  XOR U5185 ( .A(n6815), .B(n6816), .Z(n3948) );
  NOR U5186 ( .A(n6817), .B(n6815), .Z(n6816) );
  XOR U5187 ( .A(n6818), .B(n6819), .Z(n3951) );
  NOR U5188 ( .A(n6820), .B(n6818), .Z(n6819) );
  XOR U5189 ( .A(n6821), .B(n6822), .Z(n3954) );
  NOR U5190 ( .A(n6823), .B(n6821), .Z(n6822) );
  XOR U5191 ( .A(n6824), .B(n6825), .Z(n3957) );
  NOR U5192 ( .A(n6826), .B(n6824), .Z(n6825) );
  XOR U5193 ( .A(n6827), .B(n6828), .Z(n3960) );
  NOR U5194 ( .A(n6829), .B(n6827), .Z(n6828) );
  XOR U5195 ( .A(n6830), .B(n6831), .Z(n3963) );
  NOR U5196 ( .A(n6832), .B(n6830), .Z(n6831) );
  XOR U5197 ( .A(n6833), .B(n6834), .Z(n3966) );
  NOR U5198 ( .A(n6835), .B(n6833), .Z(n6834) );
  XOR U5199 ( .A(n6836), .B(n6837), .Z(n3969) );
  NOR U5200 ( .A(n6838), .B(n6836), .Z(n6837) );
  XOR U5201 ( .A(n6839), .B(n6840), .Z(n3972) );
  NOR U5202 ( .A(n6841), .B(n6839), .Z(n6840) );
  XOR U5203 ( .A(n6842), .B(n6843), .Z(n3975) );
  NOR U5204 ( .A(n6844), .B(n6842), .Z(n6843) );
  XOR U5205 ( .A(n6845), .B(n6846), .Z(n3978) );
  NOR U5206 ( .A(n6847), .B(n6845), .Z(n6846) );
  XOR U5207 ( .A(n6848), .B(n6849), .Z(n3981) );
  NOR U5208 ( .A(n6850), .B(n6848), .Z(n6849) );
  XOR U5209 ( .A(n6851), .B(n6852), .Z(n3984) );
  NOR U5210 ( .A(n6853), .B(n6851), .Z(n6852) );
  XOR U5211 ( .A(n6854), .B(n6855), .Z(n3987) );
  NOR U5212 ( .A(n6856), .B(n6854), .Z(n6855) );
  XOR U5213 ( .A(n6857), .B(n6858), .Z(n3990) );
  NOR U5214 ( .A(n6859), .B(n6857), .Z(n6858) );
  XOR U5215 ( .A(n6860), .B(n6861), .Z(n3993) );
  NOR U5216 ( .A(n6862), .B(n6860), .Z(n6861) );
  XOR U5217 ( .A(n6863), .B(n6864), .Z(n3996) );
  NOR U5218 ( .A(n6865), .B(n6863), .Z(n6864) );
  XOR U5219 ( .A(n6866), .B(n6867), .Z(n3999) );
  NOR U5220 ( .A(n6868), .B(n6866), .Z(n6867) );
  XOR U5221 ( .A(n6869), .B(n6870), .Z(n4002) );
  NOR U5222 ( .A(n6871), .B(n6869), .Z(n6870) );
  XOR U5223 ( .A(n6872), .B(n6873), .Z(n4005) );
  NOR U5224 ( .A(n6874), .B(n6872), .Z(n6873) );
  XOR U5225 ( .A(n6875), .B(n6876), .Z(n4008) );
  NOR U5226 ( .A(n6877), .B(n6875), .Z(n6876) );
  XOR U5227 ( .A(n6878), .B(n6879), .Z(n4011) );
  NOR U5228 ( .A(n6880), .B(n6878), .Z(n6879) );
  XOR U5229 ( .A(n6881), .B(n6882), .Z(n4014) );
  NOR U5230 ( .A(n6883), .B(n6881), .Z(n6882) );
  XOR U5231 ( .A(n6884), .B(n6885), .Z(n4017) );
  NOR U5232 ( .A(n6886), .B(n6884), .Z(n6885) );
  XOR U5233 ( .A(n6887), .B(n6888), .Z(n4020) );
  NOR U5234 ( .A(n6889), .B(n6887), .Z(n6888) );
  XOR U5235 ( .A(n6890), .B(n6891), .Z(n4023) );
  NOR U5236 ( .A(n6892), .B(n6890), .Z(n6891) );
  XOR U5237 ( .A(n6893), .B(n6894), .Z(n4026) );
  NOR U5238 ( .A(n6895), .B(n6893), .Z(n6894) );
  XOR U5239 ( .A(n6896), .B(n6897), .Z(n4029) );
  NOR U5240 ( .A(n6898), .B(n6896), .Z(n6897) );
  XOR U5241 ( .A(n6899), .B(n6900), .Z(n4032) );
  NOR U5242 ( .A(n6901), .B(n6899), .Z(n6900) );
  XOR U5243 ( .A(n6902), .B(n6903), .Z(n4035) );
  NOR U5244 ( .A(n6904), .B(n6902), .Z(n6903) );
  XOR U5245 ( .A(n6905), .B(n6906), .Z(n4038) );
  NOR U5246 ( .A(n6907), .B(n6905), .Z(n6906) );
  XOR U5247 ( .A(n6908), .B(n6909), .Z(n4041) );
  NOR U5248 ( .A(n6910), .B(n6908), .Z(n6909) );
  XOR U5249 ( .A(n6911), .B(n6912), .Z(n4044) );
  NOR U5250 ( .A(n6913), .B(n6911), .Z(n6912) );
  XOR U5251 ( .A(n6914), .B(n6915), .Z(n4047) );
  NOR U5252 ( .A(n6916), .B(n6914), .Z(n6915) );
  XOR U5253 ( .A(n6917), .B(n6918), .Z(n4050) );
  NOR U5254 ( .A(n6919), .B(n6917), .Z(n6918) );
  XOR U5255 ( .A(n6920), .B(n6921), .Z(n4053) );
  NOR U5256 ( .A(n6922), .B(n6920), .Z(n6921) );
  XOR U5257 ( .A(n6923), .B(n6924), .Z(n4056) );
  NOR U5258 ( .A(n6925), .B(n6923), .Z(n6924) );
  XOR U5259 ( .A(n6926), .B(n6927), .Z(n4059) );
  NOR U5260 ( .A(n6928), .B(n6926), .Z(n6927) );
  XOR U5261 ( .A(n6929), .B(n6930), .Z(n4062) );
  NOR U5262 ( .A(n6931), .B(n6929), .Z(n6930) );
  XOR U5263 ( .A(n6932), .B(n6933), .Z(n4065) );
  NOR U5264 ( .A(n6934), .B(n6932), .Z(n6933) );
  XOR U5265 ( .A(n6935), .B(n6936), .Z(n4068) );
  NOR U5266 ( .A(n6937), .B(n6935), .Z(n6936) );
  XOR U5267 ( .A(n6938), .B(n6939), .Z(n4071) );
  NOR U5268 ( .A(n6940), .B(n6938), .Z(n6939) );
  XOR U5269 ( .A(n6941), .B(n6942), .Z(n4074) );
  NOR U5270 ( .A(n6943), .B(n6941), .Z(n6942) );
  XOR U5271 ( .A(n6944), .B(n6945), .Z(n4077) );
  NOR U5272 ( .A(n6946), .B(n6944), .Z(n6945) );
  XOR U5273 ( .A(n6947), .B(n6948), .Z(n4080) );
  NOR U5274 ( .A(n6949), .B(n6947), .Z(n6948) );
  XOR U5275 ( .A(n6950), .B(n6951), .Z(n4083) );
  NOR U5276 ( .A(n6952), .B(n6950), .Z(n6951) );
  XOR U5277 ( .A(n6953), .B(n6954), .Z(n4086) );
  NOR U5278 ( .A(n6955), .B(n6953), .Z(n6954) );
  XOR U5279 ( .A(n6956), .B(n6957), .Z(n4089) );
  NOR U5280 ( .A(n6958), .B(n6956), .Z(n6957) );
  XOR U5281 ( .A(n6959), .B(n6960), .Z(n4092) );
  NOR U5282 ( .A(n6961), .B(n6959), .Z(n6960) );
  XOR U5283 ( .A(n6962), .B(n6963), .Z(n4095) );
  NOR U5284 ( .A(n6964), .B(n6962), .Z(n6963) );
  XOR U5285 ( .A(n6965), .B(n6966), .Z(n4098) );
  NOR U5286 ( .A(n6967), .B(n6965), .Z(n6966) );
  XOR U5287 ( .A(n6968), .B(n6969), .Z(n4101) );
  NOR U5288 ( .A(n6970), .B(n6968), .Z(n6969) );
  XOR U5289 ( .A(n6971), .B(n6972), .Z(n4104) );
  NOR U5290 ( .A(n6973), .B(n6971), .Z(n6972) );
  XOR U5291 ( .A(n6974), .B(n6975), .Z(n4107) );
  NOR U5292 ( .A(n6976), .B(n6974), .Z(n6975) );
  XOR U5293 ( .A(n6977), .B(n6978), .Z(n4110) );
  NOR U5294 ( .A(n6979), .B(n6977), .Z(n6978) );
  XOR U5295 ( .A(n6980), .B(n6981), .Z(n4113) );
  NOR U5296 ( .A(n6982), .B(n6980), .Z(n6981) );
  XOR U5297 ( .A(n6983), .B(n6984), .Z(n4116) );
  NOR U5298 ( .A(n6985), .B(n6983), .Z(n6984) );
  XOR U5299 ( .A(n6986), .B(n6987), .Z(n4119) );
  NOR U5300 ( .A(n6988), .B(n6986), .Z(n6987) );
  XOR U5301 ( .A(n6989), .B(n6990), .Z(n4122) );
  NOR U5302 ( .A(n6991), .B(n6989), .Z(n6990) );
  XOR U5303 ( .A(n6992), .B(n6993), .Z(n4125) );
  NOR U5304 ( .A(n6994), .B(n6992), .Z(n6993) );
  XOR U5305 ( .A(n6995), .B(n6996), .Z(n4128) );
  NOR U5306 ( .A(n6997), .B(n6995), .Z(n6996) );
  XOR U5307 ( .A(n6998), .B(n6999), .Z(n4131) );
  NOR U5308 ( .A(n7000), .B(n6998), .Z(n6999) );
  XOR U5309 ( .A(n7001), .B(n7002), .Z(n4134) );
  NOR U5310 ( .A(n7003), .B(n7001), .Z(n7002) );
  XOR U5311 ( .A(n7004), .B(n7005), .Z(n4137) );
  NOR U5312 ( .A(n7006), .B(n7004), .Z(n7005) );
  XOR U5313 ( .A(n7007), .B(n7008), .Z(n4140) );
  NOR U5314 ( .A(n7009), .B(n7007), .Z(n7008) );
  XOR U5315 ( .A(n7010), .B(n7011), .Z(n4143) );
  NOR U5316 ( .A(n7012), .B(n7010), .Z(n7011) );
  XOR U5317 ( .A(n7013), .B(n7014), .Z(n4146) );
  NOR U5318 ( .A(n7015), .B(n7013), .Z(n7014) );
  XOR U5319 ( .A(n7016), .B(n7017), .Z(n4149) );
  AND U5320 ( .A(n7018), .B(n7016), .Z(n7017) );
  XOR U5321 ( .A(n7019), .B(n7020), .Z(n4152) );
  AND U5322 ( .A(n74), .B(n7019), .Z(n7020) );
  XNOR U5323 ( .A(n5568), .B(n59), .Z(n5570) );
  IV U5324 ( .A(n56), .Z(n59) );
  XOR U5325 ( .A(n5565), .B(n5564), .Z(n56) );
  XNOR U5326 ( .A(n5562), .B(n5561), .Z(n5564) );
  XNOR U5327 ( .A(n5559), .B(n5558), .Z(n5561) );
  XNOR U5328 ( .A(n5556), .B(n5555), .Z(n5558) );
  XNOR U5329 ( .A(n5553), .B(n5552), .Z(n5555) );
  XNOR U5330 ( .A(n5550), .B(n5549), .Z(n5552) );
  XNOR U5331 ( .A(n5547), .B(n5546), .Z(n5549) );
  XNOR U5332 ( .A(n5544), .B(n5543), .Z(n5546) );
  XNOR U5333 ( .A(n5541), .B(n5540), .Z(n5543) );
  XNOR U5334 ( .A(n5538), .B(n5537), .Z(n5540) );
  XNOR U5335 ( .A(n5535), .B(n5534), .Z(n5537) );
  XNOR U5336 ( .A(n5532), .B(n5531), .Z(n5534) );
  XNOR U5337 ( .A(n5529), .B(n5528), .Z(n5531) );
  XNOR U5338 ( .A(n5526), .B(n5525), .Z(n5528) );
  XNOR U5339 ( .A(n5523), .B(n5522), .Z(n5525) );
  XNOR U5340 ( .A(n5520), .B(n5519), .Z(n5522) );
  XNOR U5341 ( .A(n5517), .B(n5516), .Z(n5519) );
  XNOR U5342 ( .A(n5514), .B(n5513), .Z(n5516) );
  XNOR U5343 ( .A(n5511), .B(n5510), .Z(n5513) );
  XNOR U5344 ( .A(n5508), .B(n5507), .Z(n5510) );
  XNOR U5345 ( .A(n5505), .B(n5504), .Z(n5507) );
  XNOR U5346 ( .A(n5502), .B(n5501), .Z(n5504) );
  XNOR U5347 ( .A(n5499), .B(n5498), .Z(n5501) );
  XNOR U5348 ( .A(n5496), .B(n5495), .Z(n5498) );
  XNOR U5349 ( .A(n5493), .B(n5492), .Z(n5495) );
  XNOR U5350 ( .A(n5490), .B(n5489), .Z(n5492) );
  XNOR U5351 ( .A(n5487), .B(n5486), .Z(n5489) );
  XNOR U5352 ( .A(n5484), .B(n5483), .Z(n5486) );
  XNOR U5353 ( .A(n5481), .B(n5480), .Z(n5483) );
  XNOR U5354 ( .A(n5478), .B(n5477), .Z(n5480) );
  XNOR U5355 ( .A(n5475), .B(n5474), .Z(n5477) );
  XNOR U5356 ( .A(n5472), .B(n5471), .Z(n5474) );
  XNOR U5357 ( .A(n5469), .B(n5468), .Z(n5471) );
  XNOR U5358 ( .A(n5466), .B(n5465), .Z(n5468) );
  XNOR U5359 ( .A(n5463), .B(n5462), .Z(n5465) );
  XNOR U5360 ( .A(n5460), .B(n5459), .Z(n5462) );
  XNOR U5361 ( .A(n5457), .B(n5456), .Z(n5459) );
  XNOR U5362 ( .A(n5454), .B(n5453), .Z(n5456) );
  XNOR U5363 ( .A(n5451), .B(n5450), .Z(n5453) );
  XNOR U5364 ( .A(n5448), .B(n5447), .Z(n5450) );
  XNOR U5365 ( .A(n5445), .B(n5444), .Z(n5447) );
  XNOR U5366 ( .A(n5442), .B(n5441), .Z(n5444) );
  XNOR U5367 ( .A(n5439), .B(n5438), .Z(n5441) );
  XNOR U5368 ( .A(n5436), .B(n5435), .Z(n5438) );
  XNOR U5369 ( .A(n5433), .B(n5432), .Z(n5435) );
  XNOR U5370 ( .A(n5430), .B(n5429), .Z(n5432) );
  XNOR U5371 ( .A(n5427), .B(n5426), .Z(n5429) );
  XNOR U5372 ( .A(n5424), .B(n5423), .Z(n5426) );
  XNOR U5373 ( .A(n5421), .B(n5420), .Z(n5423) );
  XNOR U5374 ( .A(n5418), .B(n5417), .Z(n5420) );
  XNOR U5375 ( .A(n5415), .B(n5414), .Z(n5417) );
  XNOR U5376 ( .A(n5412), .B(n5411), .Z(n5414) );
  XNOR U5377 ( .A(n5409), .B(n5408), .Z(n5411) );
  XNOR U5378 ( .A(n5406), .B(n5405), .Z(n5408) );
  XNOR U5379 ( .A(n5403), .B(n5402), .Z(n5405) );
  XNOR U5380 ( .A(n5400), .B(n5399), .Z(n5402) );
  XNOR U5381 ( .A(n5397), .B(n5396), .Z(n5399) );
  XNOR U5382 ( .A(n5394), .B(n5393), .Z(n5396) );
  XNOR U5383 ( .A(n5391), .B(n5390), .Z(n5393) );
  XNOR U5384 ( .A(n5388), .B(n5387), .Z(n5390) );
  XNOR U5385 ( .A(n5385), .B(n5384), .Z(n5387) );
  XNOR U5386 ( .A(n5382), .B(n5381), .Z(n5384) );
  XNOR U5387 ( .A(n5379), .B(n5378), .Z(n5381) );
  XNOR U5388 ( .A(n5376), .B(n5375), .Z(n5378) );
  XNOR U5389 ( .A(n5373), .B(n5372), .Z(n5375) );
  XNOR U5390 ( .A(n5370), .B(n5369), .Z(n5372) );
  XNOR U5391 ( .A(n5367), .B(n5366), .Z(n5369) );
  XNOR U5392 ( .A(n5364), .B(n5363), .Z(n5366) );
  XNOR U5393 ( .A(n5361), .B(n5360), .Z(n5363) );
  XNOR U5394 ( .A(n5358), .B(n5357), .Z(n5360) );
  XNOR U5395 ( .A(n5355), .B(n5354), .Z(n5357) );
  XNOR U5396 ( .A(n5352), .B(n5351), .Z(n5354) );
  XNOR U5397 ( .A(n5349), .B(n5348), .Z(n5351) );
  XNOR U5398 ( .A(n5346), .B(n5345), .Z(n5348) );
  XNOR U5399 ( .A(n5343), .B(n5342), .Z(n5345) );
  XNOR U5400 ( .A(n5340), .B(n5339), .Z(n5342) );
  XNOR U5401 ( .A(n5337), .B(n5336), .Z(n5339) );
  XNOR U5402 ( .A(n5334), .B(n5333), .Z(n5336) );
  XNOR U5403 ( .A(n5331), .B(n5330), .Z(n5333) );
  XNOR U5404 ( .A(n5328), .B(n5327), .Z(n5330) );
  XNOR U5405 ( .A(n5325), .B(n5324), .Z(n5327) );
  XNOR U5406 ( .A(n5322), .B(n5321), .Z(n5324) );
  XNOR U5407 ( .A(n5319), .B(n5318), .Z(n5321) );
  XNOR U5408 ( .A(n5316), .B(n5315), .Z(n5318) );
  XNOR U5409 ( .A(n5313), .B(n5312), .Z(n5315) );
  XNOR U5410 ( .A(n5310), .B(n5309), .Z(n5312) );
  XNOR U5411 ( .A(n5307), .B(n5306), .Z(n5309) );
  XNOR U5412 ( .A(n5304), .B(n5303), .Z(n5306) );
  XNOR U5413 ( .A(n5301), .B(n5300), .Z(n5303) );
  XNOR U5414 ( .A(n5298), .B(n5297), .Z(n5300) );
  XNOR U5415 ( .A(n5295), .B(n5294), .Z(n5297) );
  XNOR U5416 ( .A(n5292), .B(n5291), .Z(n5294) );
  XNOR U5417 ( .A(n5289), .B(n5288), .Z(n5291) );
  XNOR U5418 ( .A(n5286), .B(n5285), .Z(n5288) );
  XNOR U5419 ( .A(n5283), .B(n5282), .Z(n5285) );
  XNOR U5420 ( .A(n5280), .B(n5279), .Z(n5282) );
  XNOR U5421 ( .A(n5277), .B(n5276), .Z(n5279) );
  XNOR U5422 ( .A(n5274), .B(n5273), .Z(n5276) );
  XNOR U5423 ( .A(n5271), .B(n5270), .Z(n5273) );
  XNOR U5424 ( .A(n5268), .B(n5267), .Z(n5270) );
  XNOR U5425 ( .A(n5265), .B(n5264), .Z(n5267) );
  XNOR U5426 ( .A(n5262), .B(n5261), .Z(n5264) );
  XNOR U5427 ( .A(n5259), .B(n5258), .Z(n5261) );
  XNOR U5428 ( .A(n5256), .B(n5255), .Z(n5258) );
  XNOR U5429 ( .A(n5253), .B(n5252), .Z(n5255) );
  XNOR U5430 ( .A(n5250), .B(n5249), .Z(n5252) );
  XNOR U5431 ( .A(n5247), .B(n5246), .Z(n5249) );
  XNOR U5432 ( .A(n5244), .B(n5243), .Z(n5246) );
  XNOR U5433 ( .A(n5241), .B(n5240), .Z(n5243) );
  XNOR U5434 ( .A(n5238), .B(n5237), .Z(n5240) );
  XNOR U5435 ( .A(n5235), .B(n5234), .Z(n5237) );
  XNOR U5436 ( .A(n5232), .B(n5231), .Z(n5234) );
  XNOR U5437 ( .A(n5229), .B(n5228), .Z(n5231) );
  XNOR U5438 ( .A(n5226), .B(n5225), .Z(n5228) );
  XNOR U5439 ( .A(n5223), .B(n5222), .Z(n5225) );
  XNOR U5440 ( .A(n5220), .B(n5219), .Z(n5222) );
  XNOR U5441 ( .A(n5217), .B(n5216), .Z(n5219) );
  XNOR U5442 ( .A(n5214), .B(n5213), .Z(n5216) );
  XNOR U5443 ( .A(n5211), .B(n5210), .Z(n5213) );
  XNOR U5444 ( .A(n5208), .B(n5207), .Z(n5210) );
  XNOR U5445 ( .A(n5205), .B(n5204), .Z(n5207) );
  XNOR U5446 ( .A(n5202), .B(n5201), .Z(n5204) );
  XNOR U5447 ( .A(n5199), .B(n5198), .Z(n5201) );
  XNOR U5448 ( .A(n5196), .B(n5195), .Z(n5198) );
  XNOR U5449 ( .A(n5193), .B(n5192), .Z(n5195) );
  XNOR U5450 ( .A(n5190), .B(n5189), .Z(n5192) );
  XNOR U5451 ( .A(n5187), .B(n5186), .Z(n5189) );
  XNOR U5452 ( .A(n5184), .B(n5183), .Z(n5186) );
  XNOR U5453 ( .A(n5181), .B(n5180), .Z(n5183) );
  XNOR U5454 ( .A(n5178), .B(n5177), .Z(n5180) );
  XNOR U5455 ( .A(n5175), .B(n5174), .Z(n5177) );
  XNOR U5456 ( .A(n5172), .B(n5171), .Z(n5174) );
  XNOR U5457 ( .A(n5169), .B(n5168), .Z(n5171) );
  XNOR U5458 ( .A(n5166), .B(n5165), .Z(n5168) );
  XNOR U5459 ( .A(n5163), .B(n5162), .Z(n5165) );
  XNOR U5460 ( .A(n5160), .B(n5159), .Z(n5162) );
  XNOR U5461 ( .A(n5157), .B(n5156), .Z(n5159) );
  XNOR U5462 ( .A(n5154), .B(n5153), .Z(n5156) );
  XNOR U5463 ( .A(n5151), .B(n5150), .Z(n5153) );
  XNOR U5464 ( .A(n5148), .B(n5147), .Z(n5150) );
  XNOR U5465 ( .A(n5145), .B(n5144), .Z(n5147) );
  XNOR U5466 ( .A(n5142), .B(n5141), .Z(n5144) );
  XNOR U5467 ( .A(n5139), .B(n5138), .Z(n5141) );
  XNOR U5468 ( .A(n5136), .B(n5135), .Z(n5138) );
  XNOR U5469 ( .A(n5133), .B(n5132), .Z(n5135) );
  XNOR U5470 ( .A(n5130), .B(n5129), .Z(n5132) );
  XNOR U5471 ( .A(n5127), .B(n5126), .Z(n5129) );
  XNOR U5472 ( .A(n5124), .B(n5123), .Z(n5126) );
  XNOR U5473 ( .A(n5121), .B(n5120), .Z(n5123) );
  XNOR U5474 ( .A(n5118), .B(n5117), .Z(n5120) );
  XNOR U5475 ( .A(n5115), .B(n5114), .Z(n5117) );
  XNOR U5476 ( .A(n5112), .B(n5111), .Z(n5114) );
  XNOR U5477 ( .A(n5109), .B(n5108), .Z(n5111) );
  XNOR U5478 ( .A(n5106), .B(n5105), .Z(n5108) );
  XNOR U5479 ( .A(n5103), .B(n5102), .Z(n5105) );
  XNOR U5480 ( .A(n5100), .B(n5099), .Z(n5102) );
  XNOR U5481 ( .A(n5097), .B(n5096), .Z(n5099) );
  XNOR U5482 ( .A(n5094), .B(n5093), .Z(n5096) );
  XNOR U5483 ( .A(n5091), .B(n5090), .Z(n5093) );
  XNOR U5484 ( .A(n5088), .B(n5087), .Z(n5090) );
  XNOR U5485 ( .A(n5085), .B(n5084), .Z(n5087) );
  XNOR U5486 ( .A(n5082), .B(n5081), .Z(n5084) );
  XNOR U5487 ( .A(n5079), .B(n5078), .Z(n5081) );
  XNOR U5488 ( .A(n5076), .B(n5075), .Z(n5078) );
  XNOR U5489 ( .A(n5073), .B(n5072), .Z(n5075) );
  XNOR U5490 ( .A(n5070), .B(n5069), .Z(n5072) );
  XNOR U5491 ( .A(n5067), .B(n5066), .Z(n5069) );
  XNOR U5492 ( .A(n5064), .B(n5063), .Z(n5066) );
  XNOR U5493 ( .A(n5061), .B(n5060), .Z(n5063) );
  XNOR U5494 ( .A(n5058), .B(n5057), .Z(n5060) );
  XNOR U5495 ( .A(n5055), .B(n5054), .Z(n5057) );
  XNOR U5496 ( .A(n5052), .B(n5051), .Z(n5054) );
  XNOR U5497 ( .A(n5049), .B(n5048), .Z(n5051) );
  XNOR U5498 ( .A(n5046), .B(n5045), .Z(n5048) );
  XNOR U5499 ( .A(n5043), .B(n5042), .Z(n5045) );
  XNOR U5500 ( .A(n5040), .B(n5039), .Z(n5042) );
  XNOR U5501 ( .A(n5037), .B(n5036), .Z(n5039) );
  XNOR U5502 ( .A(n5034), .B(n5033), .Z(n5036) );
  XNOR U5503 ( .A(n5031), .B(n5030), .Z(n5033) );
  XNOR U5504 ( .A(n5028), .B(n5027), .Z(n5030) );
  XNOR U5505 ( .A(n5025), .B(n5024), .Z(n5027) );
  XNOR U5506 ( .A(n5022), .B(n5021), .Z(n5024) );
  XNOR U5507 ( .A(n5019), .B(n5018), .Z(n5021) );
  XNOR U5508 ( .A(n5016), .B(n5015), .Z(n5018) );
  XNOR U5509 ( .A(n5013), .B(n5012), .Z(n5015) );
  XNOR U5510 ( .A(n5010), .B(n5009), .Z(n5012) );
  XNOR U5511 ( .A(n5007), .B(n5006), .Z(n5009) );
  XNOR U5512 ( .A(n5004), .B(n5003), .Z(n5006) );
  XNOR U5513 ( .A(n5001), .B(n5000), .Z(n5003) );
  XNOR U5514 ( .A(n4998), .B(n4997), .Z(n5000) );
  XNOR U5515 ( .A(n4995), .B(n4994), .Z(n4997) );
  XNOR U5516 ( .A(n4992), .B(n4991), .Z(n4994) );
  XNOR U5517 ( .A(n4989), .B(n4988), .Z(n4991) );
  XNOR U5518 ( .A(n4986), .B(n4985), .Z(n4988) );
  XNOR U5519 ( .A(n4983), .B(n4982), .Z(n4985) );
  XNOR U5520 ( .A(n4980), .B(n4979), .Z(n4982) );
  XNOR U5521 ( .A(n4977), .B(n4976), .Z(n4979) );
  XNOR U5522 ( .A(n4974), .B(n4973), .Z(n4976) );
  XNOR U5523 ( .A(n4971), .B(n4970), .Z(n4973) );
  XNOR U5524 ( .A(n4968), .B(n4967), .Z(n4970) );
  XNOR U5525 ( .A(n4965), .B(n4964), .Z(n4967) );
  XNOR U5526 ( .A(n4962), .B(n4961), .Z(n4964) );
  XNOR U5527 ( .A(n4959), .B(n4958), .Z(n4961) );
  XNOR U5528 ( .A(n4956), .B(n4955), .Z(n4958) );
  XNOR U5529 ( .A(n4953), .B(n4952), .Z(n4955) );
  XNOR U5530 ( .A(n4950), .B(n4949), .Z(n4952) );
  XNOR U5531 ( .A(n4947), .B(n4946), .Z(n4949) );
  XNOR U5532 ( .A(n4944), .B(n4943), .Z(n4946) );
  XNOR U5533 ( .A(n4941), .B(n4940), .Z(n4943) );
  XNOR U5534 ( .A(n4938), .B(n4937), .Z(n4940) );
  XNOR U5535 ( .A(n4935), .B(n4934), .Z(n4937) );
  XNOR U5536 ( .A(n4932), .B(n4931), .Z(n4934) );
  XNOR U5537 ( .A(n4929), .B(n4928), .Z(n4931) );
  XNOR U5538 ( .A(n4926), .B(n4925), .Z(n4928) );
  XNOR U5539 ( .A(n4923), .B(n4922), .Z(n4925) );
  XNOR U5540 ( .A(n4920), .B(n4919), .Z(n4922) );
  XNOR U5541 ( .A(n4917), .B(n4916), .Z(n4919) );
  XNOR U5542 ( .A(n4914), .B(n4913), .Z(n4916) );
  XNOR U5543 ( .A(n4911), .B(n4910), .Z(n4913) );
  XNOR U5544 ( .A(n4908), .B(n4907), .Z(n4910) );
  XNOR U5545 ( .A(n4905), .B(n4904), .Z(n4907) );
  XNOR U5546 ( .A(n4902), .B(n4901), .Z(n4904) );
  XNOR U5547 ( .A(n4899), .B(n4898), .Z(n4901) );
  XNOR U5548 ( .A(n4896), .B(n4895), .Z(n4898) );
  XNOR U5549 ( .A(n4893), .B(n4892), .Z(n4895) );
  XNOR U5550 ( .A(n4890), .B(n4889), .Z(n4892) );
  XNOR U5551 ( .A(n4887), .B(n4886), .Z(n4889) );
  XNOR U5552 ( .A(n4884), .B(n4883), .Z(n4886) );
  XNOR U5553 ( .A(n4881), .B(n4880), .Z(n4883) );
  XNOR U5554 ( .A(n4878), .B(n4877), .Z(n4880) );
  XNOR U5555 ( .A(n4875), .B(n4874), .Z(n4877) );
  XNOR U5556 ( .A(n4872), .B(n4871), .Z(n4874) );
  XNOR U5557 ( .A(n4869), .B(n4868), .Z(n4871) );
  XNOR U5558 ( .A(n4866), .B(n4865), .Z(n4868) );
  XNOR U5559 ( .A(n4863), .B(n4862), .Z(n4865) );
  XNOR U5560 ( .A(n4860), .B(n4859), .Z(n4862) );
  XNOR U5561 ( .A(n4857), .B(n4856), .Z(n4859) );
  XNOR U5562 ( .A(n4854), .B(n4853), .Z(n4856) );
  XNOR U5563 ( .A(n4851), .B(n4850), .Z(n4853) );
  XNOR U5564 ( .A(n4848), .B(n4847), .Z(n4850) );
  XNOR U5565 ( .A(n4845), .B(n4844), .Z(n4847) );
  XNOR U5566 ( .A(n4842), .B(n4841), .Z(n4844) );
  XNOR U5567 ( .A(n4839), .B(n4838), .Z(n4841) );
  XNOR U5568 ( .A(n4836), .B(n4835), .Z(n4838) );
  XNOR U5569 ( .A(n4833), .B(n4832), .Z(n4835) );
  XNOR U5570 ( .A(n4830), .B(n4829), .Z(n4832) );
  XNOR U5571 ( .A(n4827), .B(n4826), .Z(n4829) );
  XNOR U5572 ( .A(n4824), .B(n4823), .Z(n4826) );
  XNOR U5573 ( .A(n4821), .B(n4820), .Z(n4823) );
  XNOR U5574 ( .A(n4818), .B(n4817), .Z(n4820) );
  XNOR U5575 ( .A(n4815), .B(n4814), .Z(n4817) );
  XNOR U5576 ( .A(n4812), .B(n4811), .Z(n4814) );
  XNOR U5577 ( .A(n4809), .B(n4808), .Z(n4811) );
  XNOR U5578 ( .A(n4806), .B(n4805), .Z(n4808) );
  XNOR U5579 ( .A(n4803), .B(n4802), .Z(n4805) );
  XNOR U5580 ( .A(n4800), .B(n4799), .Z(n4802) );
  XNOR U5581 ( .A(n4797), .B(n4178), .Z(n4799) );
  XOR U5582 ( .A(n4177), .B(n4166), .Z(n4178) );
  XOR U5583 ( .A(n7021), .B(n4164), .Z(n4166) );
  XNOR U5584 ( .A(n4165), .B(n4161), .Z(n4164) );
  XNOR U5585 ( .A(n4160), .B(n4187), .Z(n4161) );
  XNOR U5586 ( .A(n4186), .B(n4796), .Z(n4187) );
  XNOR U5587 ( .A(n4787), .B(n4795), .Z(n4796) );
  XNOR U5588 ( .A(n4786), .B(n4792), .Z(n4795) );
  XNOR U5589 ( .A(n4791), .B(n4196), .Z(n4792) );
  XNOR U5590 ( .A(n4195), .B(n4785), .Z(n4196) );
  XNOR U5591 ( .A(n4776), .B(n4784), .Z(n4785) );
  XNOR U5592 ( .A(n4775), .B(n4781), .Z(n4784) );
  XNOR U5593 ( .A(n4780), .B(n4205), .Z(n4781) );
  XNOR U5594 ( .A(n4204), .B(n4774), .Z(n4205) );
  XNOR U5595 ( .A(n4765), .B(n4773), .Z(n4774) );
  XNOR U5596 ( .A(n4764), .B(n4770), .Z(n4773) );
  XNOR U5597 ( .A(n4769), .B(n4214), .Z(n4770) );
  XNOR U5598 ( .A(n4213), .B(n4763), .Z(n4214) );
  XNOR U5599 ( .A(n4754), .B(n4762), .Z(n4763) );
  XNOR U5600 ( .A(n4753), .B(n4759), .Z(n4762) );
  XNOR U5601 ( .A(n4758), .B(n4223), .Z(n4759) );
  XNOR U5602 ( .A(n4222), .B(n4752), .Z(n4223) );
  XNOR U5603 ( .A(n4743), .B(n4751), .Z(n4752) );
  XNOR U5604 ( .A(n4742), .B(n4748), .Z(n4751) );
  XNOR U5605 ( .A(n4747), .B(n4232), .Z(n4748) );
  XNOR U5606 ( .A(n4231), .B(n4741), .Z(n4232) );
  XNOR U5607 ( .A(n4732), .B(n4740), .Z(n4741) );
  XNOR U5608 ( .A(n4731), .B(n4737), .Z(n4740) );
  XNOR U5609 ( .A(n4736), .B(n4241), .Z(n4737) );
  XNOR U5610 ( .A(n4240), .B(n4730), .Z(n4241) );
  XNOR U5611 ( .A(n4721), .B(n4729), .Z(n4730) );
  XNOR U5612 ( .A(n4720), .B(n4726), .Z(n4729) );
  XNOR U5613 ( .A(n4725), .B(n4250), .Z(n4726) );
  XNOR U5614 ( .A(n4249), .B(n4719), .Z(n4250) );
  XNOR U5615 ( .A(n4710), .B(n4718), .Z(n4719) );
  XNOR U5616 ( .A(n4709), .B(n4715), .Z(n4718) );
  XNOR U5617 ( .A(n4714), .B(n4259), .Z(n4715) );
  XNOR U5618 ( .A(n4258), .B(n4708), .Z(n4259) );
  XNOR U5619 ( .A(n4699), .B(n4707), .Z(n4708) );
  XNOR U5620 ( .A(n4698), .B(n4704), .Z(n4707) );
  XNOR U5621 ( .A(n4703), .B(n4268), .Z(n4704) );
  XNOR U5622 ( .A(n4267), .B(n4697), .Z(n4268) );
  XNOR U5623 ( .A(n4688), .B(n4696), .Z(n4697) );
  XNOR U5624 ( .A(n4687), .B(n4693), .Z(n4696) );
  XNOR U5625 ( .A(n4692), .B(n4277), .Z(n4693) );
  XNOR U5626 ( .A(n4276), .B(n4686), .Z(n4277) );
  XNOR U5627 ( .A(n4677), .B(n4685), .Z(n4686) );
  XNOR U5628 ( .A(n4676), .B(n4682), .Z(n4685) );
  XNOR U5629 ( .A(n4681), .B(n4286), .Z(n4682) );
  XNOR U5630 ( .A(n4285), .B(n4675), .Z(n4286) );
  XNOR U5631 ( .A(n4666), .B(n4674), .Z(n4675) );
  XNOR U5632 ( .A(n4665), .B(n4671), .Z(n4674) );
  XNOR U5633 ( .A(n4670), .B(n4295), .Z(n4671) );
  XNOR U5634 ( .A(n4294), .B(n4664), .Z(n4295) );
  XNOR U5635 ( .A(n4655), .B(n4663), .Z(n4664) );
  XNOR U5636 ( .A(n4654), .B(n4660), .Z(n4663) );
  XNOR U5637 ( .A(n4659), .B(n4304), .Z(n4660) );
  XNOR U5638 ( .A(n4303), .B(n4653), .Z(n4304) );
  XNOR U5639 ( .A(n4644), .B(n4652), .Z(n4653) );
  XNOR U5640 ( .A(n4643), .B(n4649), .Z(n4652) );
  XNOR U5641 ( .A(n4648), .B(n4313), .Z(n4649) );
  XNOR U5642 ( .A(n4312), .B(n4642), .Z(n4313) );
  XNOR U5643 ( .A(n4633), .B(n4641), .Z(n4642) );
  XNOR U5644 ( .A(n4632), .B(n4638), .Z(n4641) );
  XNOR U5645 ( .A(n4637), .B(n4322), .Z(n4638) );
  XNOR U5646 ( .A(n4321), .B(n4631), .Z(n4322) );
  XNOR U5647 ( .A(n4622), .B(n4630), .Z(n4631) );
  XNOR U5648 ( .A(n4621), .B(n4627), .Z(n4630) );
  XNOR U5649 ( .A(n4626), .B(n4331), .Z(n4627) );
  XNOR U5650 ( .A(n4330), .B(n4620), .Z(n4331) );
  XNOR U5651 ( .A(n4611), .B(n4619), .Z(n4620) );
  XNOR U5652 ( .A(n4610), .B(n4616), .Z(n4619) );
  XNOR U5653 ( .A(n4615), .B(n4340), .Z(n4616) );
  XNOR U5654 ( .A(n4339), .B(n4609), .Z(n4340) );
  XNOR U5655 ( .A(n4600), .B(n4608), .Z(n4609) );
  XNOR U5656 ( .A(n4599), .B(n4605), .Z(n4608) );
  XNOR U5657 ( .A(n4604), .B(n4349), .Z(n4605) );
  XNOR U5658 ( .A(n4348), .B(n4598), .Z(n4349) );
  XNOR U5659 ( .A(n4589), .B(n4597), .Z(n4598) );
  XNOR U5660 ( .A(n4588), .B(n4594), .Z(n4597) );
  XNOR U5661 ( .A(n4593), .B(n4358), .Z(n4594) );
  XNOR U5662 ( .A(n4357), .B(n4587), .Z(n4358) );
  XNOR U5663 ( .A(n4578), .B(n4586), .Z(n4587) );
  XNOR U5664 ( .A(n4577), .B(n4583), .Z(n4586) );
  XNOR U5665 ( .A(n4582), .B(n4367), .Z(n4583) );
  XNOR U5666 ( .A(n4366), .B(n4576), .Z(n4367) );
  XNOR U5667 ( .A(n4567), .B(n4575), .Z(n4576) );
  XNOR U5668 ( .A(n4566), .B(n4572), .Z(n4575) );
  XNOR U5669 ( .A(n4571), .B(n4376), .Z(n4572) );
  XNOR U5670 ( .A(n4375), .B(n4565), .Z(n4376) );
  XNOR U5671 ( .A(n4556), .B(n4564), .Z(n4565) );
  XNOR U5672 ( .A(n4555), .B(n4561), .Z(n4564) );
  XNOR U5673 ( .A(n4560), .B(n4385), .Z(n4561) );
  XNOR U5674 ( .A(n4384), .B(n4554), .Z(n4385) );
  XNOR U5675 ( .A(n4545), .B(n4553), .Z(n4554) );
  XNOR U5676 ( .A(n4544), .B(n4550), .Z(n4553) );
  XNOR U5677 ( .A(n4549), .B(n4394), .Z(n4550) );
  XNOR U5678 ( .A(n4393), .B(n4543), .Z(n4394) );
  XNOR U5679 ( .A(n4534), .B(n4542), .Z(n4543) );
  XNOR U5680 ( .A(n4533), .B(n4539), .Z(n4542) );
  XNOR U5681 ( .A(n4538), .B(n4403), .Z(n4539) );
  XNOR U5682 ( .A(n4402), .B(n4532), .Z(n4403) );
  XNOR U5683 ( .A(n4523), .B(n4531), .Z(n4532) );
  XNOR U5684 ( .A(n4522), .B(n4528), .Z(n4531) );
  XNOR U5685 ( .A(n4527), .B(n4412), .Z(n4528) );
  XNOR U5686 ( .A(n4411), .B(n4521), .Z(n4412) );
  XNOR U5687 ( .A(n4512), .B(n4520), .Z(n4521) );
  XNOR U5688 ( .A(n4511), .B(n4517), .Z(n4520) );
  XNOR U5689 ( .A(n4516), .B(n4421), .Z(n4517) );
  XNOR U5690 ( .A(n4420), .B(n4510), .Z(n4421) );
  XNOR U5691 ( .A(n4501), .B(n4509), .Z(n4510) );
  XNOR U5692 ( .A(n4500), .B(n4506), .Z(n4509) );
  XNOR U5693 ( .A(n4505), .B(n4430), .Z(n4506) );
  XNOR U5694 ( .A(n4429), .B(n4499), .Z(n4430) );
  XNOR U5695 ( .A(n4490), .B(n4498), .Z(n4499) );
  XNOR U5696 ( .A(n4489), .B(n4495), .Z(n4498) );
  XNOR U5697 ( .A(n4494), .B(n4477), .Z(n4495) );
  XNOR U5698 ( .A(n4436), .B(n4488), .Z(n4477) );
  XNOR U5699 ( .A(n4479), .B(n4487), .Z(n4488) );
  XNOR U5700 ( .A(n4478), .B(n4484), .Z(n4487) );
  XNOR U5701 ( .A(n4483), .B(n4467), .Z(n4484) );
  XNOR U5702 ( .A(n4439), .B(n4476), .Z(n4467) );
  XNOR U5703 ( .A(n4463), .B(n4473), .Z(n4476) );
  XNOR U5704 ( .A(n4466), .B(n4472), .Z(n4473) );
  XNOR U5705 ( .A(n4435), .B(n4462), .Z(n4472) );
  XNOR U5706 ( .A(n4445), .B(n4461), .Z(n4462) );
  XNOR U5707 ( .A(n4448), .B(n4458), .Z(n4461) );
  XOR U5708 ( .A(n4447), .B(n4455), .Z(n4458) );
  XOR U5709 ( .A(n4456), .B(n4454), .Z(n4455) );
  XOR U5710 ( .A(n7022), .B(n7023), .Z(n4454) );
  XOR U5711 ( .A(n7024), .B(n7025), .Z(n7023) );
  XNOR U5712 ( .A(n7026), .B(n7027), .Z(n7025) );
  NOR U5713 ( .A(n7028), .B(n7027), .Z(n7026) );
  XOR U5714 ( .A(n7029), .B(n7030), .Z(n7024) );
  NOR U5715 ( .A(n7031), .B(n7032), .Z(n7030) );
  NOR U5716 ( .A(n7033), .B(n7034), .Z(n7029) );
  XOR U5717 ( .A(n7035), .B(n7036), .Z(n7022) );
  XOR U5718 ( .A(n7037), .B(n7038), .Z(n7036) );
  XOR U5719 ( .A(n7039), .B(n7040), .Z(n7038) );
  XOR U5720 ( .A(n7041), .B(n7042), .Z(n7040) );
  XOR U5721 ( .A(n7043), .B(n7044), .Z(n7042) );
  AND U5722 ( .A(n7045), .B(n7044), .Z(n7043) );
  XOR U5723 ( .A(n7046), .B(n7047), .Z(n7041) );
  XOR U5724 ( .A(n7048), .B(n7049), .Z(n7047) );
  XOR U5725 ( .A(n7050), .B(n7051), .Z(n7049) );
  XNOR U5726 ( .A(n7052), .B(n7053), .Z(n7051) );
  NOR U5727 ( .A(n7054), .B(n7053), .Z(n7052) );
  XOR U5728 ( .A(n7055), .B(n7056), .Z(n7050) );
  XOR U5729 ( .A(n7057), .B(n7058), .Z(n7056) );
  XNOR U5730 ( .A(n7059), .B(n7060), .Z(n7058) );
  XOR U5731 ( .A(n7061), .B(n7062), .Z(n7057) );
  XOR U5732 ( .A(n7063), .B(n7064), .Z(n7062) );
  XOR U5733 ( .A(n7065), .B(n7066), .Z(n7064) );
  XOR U5734 ( .A(n7067), .B(n7068), .Z(n7066) );
  XOR U5735 ( .A(n7069), .B(n7070), .Z(n7068) );
  XOR U5736 ( .A(n7071), .B(n7072), .Z(n7070) );
  XOR U5737 ( .A(n7073), .B(n7074), .Z(n7072) );
  XOR U5738 ( .A(n7075), .B(n7076), .Z(n7074) );
  XOR U5739 ( .A(n7077), .B(n7078), .Z(n7076) );
  XOR U5740 ( .A(n7079), .B(n7080), .Z(n7078) );
  XOR U5741 ( .A(n7081), .B(n7082), .Z(n7080) );
  XOR U5742 ( .A(n7083), .B(n7084), .Z(n7082) );
  XOR U5743 ( .A(n7085), .B(n7086), .Z(n7084) );
  XOR U5744 ( .A(n7087), .B(n7088), .Z(n7086) );
  XOR U5745 ( .A(n7089), .B(n7090), .Z(n7088) );
  XOR U5746 ( .A(n7091), .B(n7092), .Z(n7090) );
  XOR U5747 ( .A(n7093), .B(n7094), .Z(n7092) );
  AND U5748 ( .A(n7095), .B(n7096), .Z(n7094) );
  AND U5749 ( .A(n7097), .B(n7098), .Z(n7093) );
  XOR U5750 ( .A(n7099), .B(n7100), .Z(n7091) );
  AND U5751 ( .A(n7101), .B(n7102), .Z(n7100) );
  NOR U5752 ( .A(n7103), .B(n7104), .Z(n7102) );
  IV U5753 ( .A(n7105), .Z(n7103) );
  NOR U5754 ( .A(n7106), .B(n7107), .Z(n7105) );
  AND U5755 ( .A(n7108), .B(n7109), .Z(n7101) );
  NOR U5756 ( .A(n7110), .B(n7111), .Z(n7108) );
  NOR U5757 ( .A(n7112), .B(n7113), .Z(n7099) );
  XOR U5758 ( .A(n7114), .B(n7115), .Z(n7089) );
  XOR U5759 ( .A(n7116), .B(n7117), .Z(n7115) );
  NOR U5760 ( .A(n7118), .B(n7119), .Z(n7117) );
  AND U5761 ( .A(n7120), .B(n7121), .Z(n7119) );
  IV U5762 ( .A(n7122), .Z(n7118) );
  NOR U5763 ( .A(n7123), .B(n7124), .Z(n7122) );
  AND U5764 ( .A(n7112), .B(n7125), .Z(n7124) );
  AND U5765 ( .A(n7113), .B(n7126), .Z(n7123) );
  NOR U5766 ( .A(n7127), .B(n7128), .Z(n7116) );
  XOR U5767 ( .A(n7129), .B(n7130), .Z(n7114) );
  NOR U5768 ( .A(n7131), .B(n7132), .Z(n7130) );
  AND U5769 ( .A(n7133), .B(n7134), .Z(n7132) );
  IV U5770 ( .A(n7135), .Z(n7131) );
  NOR U5771 ( .A(n7136), .B(n7137), .Z(n7135) );
  AND U5772 ( .A(n7127), .B(n7138), .Z(n7137) );
  AND U5773 ( .A(n7128), .B(n7139), .Z(n7136) );
  NOR U5774 ( .A(n7140), .B(n7141), .Z(n7129) );
  AND U5775 ( .A(n7142), .B(n7143), .Z(n7087) );
  XOR U5776 ( .A(n7144), .B(n7145), .Z(n7085) );
  AND U5777 ( .A(n7146), .B(n7147), .Z(n7145) );
  NOR U5778 ( .A(n7148), .B(n7149), .Z(n7144) );
  AND U5779 ( .A(n7150), .B(n7151), .Z(n7149) );
  IV U5780 ( .A(n7152), .Z(n7148) );
  NOR U5781 ( .A(n7153), .B(n7154), .Z(n7152) );
  AND U5782 ( .A(n7140), .B(n7155), .Z(n7154) );
  AND U5783 ( .A(n7141), .B(n7156), .Z(n7153) );
  XOR U5784 ( .A(n7157), .B(n7158), .Z(n7083) );
  XOR U5785 ( .A(n7159), .B(n7160), .Z(n7158) );
  NOR U5786 ( .A(n7161), .B(n7162), .Z(n7160) );
  NOR U5787 ( .A(n7163), .B(n7164), .Z(n7159) );
  AND U5788 ( .A(n7165), .B(n7166), .Z(n7164) );
  IV U5789 ( .A(n7167), .Z(n7163) );
  NOR U5790 ( .A(n7168), .B(n7169), .Z(n7167) );
  AND U5791 ( .A(n7161), .B(n7170), .Z(n7169) );
  AND U5792 ( .A(n7162), .B(n7171), .Z(n7168) );
  XOR U5793 ( .A(n7172), .B(n7173), .Z(n7157) );
  NOR U5794 ( .A(n7174), .B(n7175), .Z(n7173) );
  NOR U5795 ( .A(n7176), .B(n7177), .Z(n7172) );
  AND U5796 ( .A(n7178), .B(n7179), .Z(n7177) );
  IV U5797 ( .A(n7180), .Z(n7176) );
  NOR U5798 ( .A(n7181), .B(n7182), .Z(n7180) );
  AND U5799 ( .A(n7174), .B(n7183), .Z(n7182) );
  AND U5800 ( .A(n7175), .B(n7184), .Z(n7181) );
  AND U5801 ( .A(n7185), .B(n7186), .Z(n7081) );
  XOR U5802 ( .A(n7187), .B(n7188), .Z(n7079) );
  AND U5803 ( .A(n7189), .B(n7190), .Z(n7188) );
  AND U5804 ( .A(n7191), .B(n7192), .Z(n7187) );
  XOR U5805 ( .A(n7193), .B(n7194), .Z(n7077) );
  XOR U5806 ( .A(n7195), .B(n7196), .Z(n7194) );
  NOR U5807 ( .A(n7197), .B(n7198), .Z(n7196) );
  NOR U5808 ( .A(n7199), .B(n7200), .Z(n7195) );
  AND U5809 ( .A(n7201), .B(n7202), .Z(n7200) );
  IV U5810 ( .A(n7203), .Z(n7199) );
  NOR U5811 ( .A(n7204), .B(n7205), .Z(n7203) );
  AND U5812 ( .A(n7197), .B(n7206), .Z(n7205) );
  AND U5813 ( .A(n7198), .B(n7207), .Z(n7204) );
  XOR U5814 ( .A(n7208), .B(n7209), .Z(n7193) );
  NOR U5815 ( .A(n7210), .B(n7211), .Z(n7209) );
  NOR U5816 ( .A(n7212), .B(n7213), .Z(n7208) );
  AND U5817 ( .A(n7214), .B(n7215), .Z(n7213) );
  IV U5818 ( .A(n7216), .Z(n7212) );
  NOR U5819 ( .A(n7217), .B(n7218), .Z(n7216) );
  AND U5820 ( .A(n7210), .B(n7219), .Z(n7218) );
  AND U5821 ( .A(n7211), .B(n7220), .Z(n7217) );
  AND U5822 ( .A(n7221), .B(n7222), .Z(n7075) );
  XOR U5823 ( .A(n7223), .B(n7224), .Z(n7073) );
  AND U5824 ( .A(n7225), .B(n7226), .Z(n7224) );
  NOR U5825 ( .A(n7227), .B(n7228), .Z(n7223) );
  XOR U5826 ( .A(n7229), .B(n7230), .Z(n7071) );
  XOR U5827 ( .A(n7231), .B(n7232), .Z(n7230) );
  NOR U5828 ( .A(n7233), .B(n7234), .Z(n7232) );
  AND U5829 ( .A(n7235), .B(n7236), .Z(n7234) );
  IV U5830 ( .A(n7237), .Z(n7233) );
  NOR U5831 ( .A(n7238), .B(n7239), .Z(n7237) );
  AND U5832 ( .A(n7227), .B(n7240), .Z(n7239) );
  AND U5833 ( .A(n7228), .B(n7241), .Z(n7238) );
  NOR U5834 ( .A(n7242), .B(n7243), .Z(n7231) );
  XOR U5835 ( .A(n7244), .B(n7245), .Z(n7229) );
  NOR U5836 ( .A(n7246), .B(n7247), .Z(n7245) );
  AND U5837 ( .A(n7248), .B(n7249), .Z(n7247) );
  IV U5838 ( .A(n7250), .Z(n7246) );
  NOR U5839 ( .A(n7251), .B(n7252), .Z(n7250) );
  AND U5840 ( .A(n7242), .B(n7253), .Z(n7252) );
  AND U5841 ( .A(n7243), .B(n7254), .Z(n7251) );
  NOR U5842 ( .A(n7255), .B(n7256), .Z(n7244) );
  NOR U5843 ( .A(n7257), .B(n7258), .Z(n7069) );
  AND U5844 ( .A(n7259), .B(n7260), .Z(n7258) );
  IV U5845 ( .A(n7261), .Z(n7257) );
  NOR U5846 ( .A(n7262), .B(n7263), .Z(n7261) );
  AND U5847 ( .A(n7255), .B(n7264), .Z(n7263) );
  AND U5848 ( .A(n7256), .B(n7265), .Z(n7262) );
  XOR U5849 ( .A(n7266), .B(n7267), .Z(n7067) );
  NOR U5850 ( .A(n7268), .B(n7269), .Z(n7267) );
  AND U5851 ( .A(n7270), .B(n7271), .Z(n7266) );
  XOR U5852 ( .A(n7272), .B(n7273), .Z(n7065) );
  XOR U5853 ( .A(n7274), .B(n7275), .Z(n7273) );
  AND U5854 ( .A(n7268), .B(n7276), .Z(n7274) );
  XOR U5855 ( .A(n7277), .B(n7278), .Z(n7272) );
  AND U5856 ( .A(n7269), .B(n7279), .Z(n7278) );
  AND U5857 ( .A(n7275), .B(n7280), .Z(n7277) );
  XOR U5858 ( .A(n7281), .B(n7282), .Z(n7061) );
  XOR U5859 ( .A(n7283), .B(n7284), .Z(n7282) );
  AND U5860 ( .A(n7285), .B(n7063), .Z(n7283) );
  XOR U5861 ( .A(n7286), .B(n7287), .Z(n7055) );
  XOR U5862 ( .A(n7288), .B(n7289), .Z(n7287) );
  AND U5863 ( .A(n7059), .B(n7290), .Z(n7289) );
  AND U5864 ( .A(n7291), .B(n7284), .Z(n7288) );
  XOR U5865 ( .A(n7292), .B(n7293), .Z(n7286) );
  AND U5866 ( .A(n7294), .B(n7281), .Z(n7293) );
  NOR U5867 ( .A(n7295), .B(n7060), .Z(n7292) );
  XOR U5868 ( .A(n7296), .B(n7297), .Z(n7048) );
  XOR U5869 ( .A(n7298), .B(n7299), .Z(n7046) );
  XOR U5870 ( .A(n7300), .B(n7301), .Z(n7299) );
  AND U5871 ( .A(n7302), .B(n7301), .Z(n7300) );
  XOR U5872 ( .A(n7303), .B(n7304), .Z(n7298) );
  NOR U5873 ( .A(n7305), .B(n7296), .Z(n7304) );
  NOR U5874 ( .A(n7306), .B(n7297), .Z(n7303) );
  XOR U5875 ( .A(n7307), .B(n7308), .Z(n7039) );
  XOR U5876 ( .A(n7309), .B(n7310), .Z(n7037) );
  XNOR U5877 ( .A(n7311), .B(n7312), .Z(n7310) );
  NOR U5878 ( .A(n7313), .B(n7312), .Z(n7311) );
  XOR U5879 ( .A(n7314), .B(n7315), .Z(n7309) );
  NOR U5880 ( .A(n7316), .B(n7307), .Z(n7315) );
  NOR U5881 ( .A(n7317), .B(n7308), .Z(n7314) );
  XNOR U5882 ( .A(n7034), .B(n7032), .Z(n7035) );
  XNOR U5883 ( .A(n7318), .B(n7319), .Z(n4456) );
  NOR U5884 ( .A(n7320), .B(n7318), .Z(n7319) );
  XOR U5885 ( .A(n7321), .B(n7322), .Z(n4447) );
  NOR U5886 ( .A(n7323), .B(n7321), .Z(n7322) );
  XOR U5887 ( .A(n7324), .B(n7325), .Z(n4448) );
  NOR U5888 ( .A(n7326), .B(n7324), .Z(n7325) );
  XOR U5889 ( .A(n7327), .B(n7328), .Z(n4445) );
  NOR U5890 ( .A(n7329), .B(n7327), .Z(n7328) );
  XOR U5891 ( .A(n7330), .B(n7331), .Z(n4435) );
  NOR U5892 ( .A(n7332), .B(n7330), .Z(n7331) );
  XOR U5893 ( .A(n7333), .B(n7334), .Z(n4466) );
  NOR U5894 ( .A(n7335), .B(n7333), .Z(n7334) );
  XOR U5895 ( .A(n7336), .B(n7337), .Z(n4463) );
  NOR U5896 ( .A(n7338), .B(n7336), .Z(n7337) );
  XOR U5897 ( .A(n7339), .B(n7340), .Z(n4439) );
  NOR U5898 ( .A(n7341), .B(n7339), .Z(n7340) );
  XOR U5899 ( .A(n7342), .B(n7343), .Z(n4483) );
  NOR U5900 ( .A(n7344), .B(n7342), .Z(n7343) );
  XOR U5901 ( .A(n7345), .B(n7346), .Z(n4478) );
  NOR U5902 ( .A(n7347), .B(n7345), .Z(n7346) );
  XOR U5903 ( .A(n7348), .B(n7349), .Z(n4479) );
  NOR U5904 ( .A(n7350), .B(n7348), .Z(n7349) );
  XOR U5905 ( .A(n7351), .B(n7352), .Z(n4436) );
  NOR U5906 ( .A(n7353), .B(n7351), .Z(n7352) );
  XOR U5907 ( .A(n7354), .B(n7355), .Z(n4494) );
  NOR U5908 ( .A(n7356), .B(n7354), .Z(n7355) );
  XOR U5909 ( .A(n7357), .B(n7358), .Z(n4489) );
  NOR U5910 ( .A(n7359), .B(n7357), .Z(n7358) );
  XOR U5911 ( .A(n7360), .B(n7361), .Z(n4490) );
  NOR U5912 ( .A(n7362), .B(n7360), .Z(n7361) );
  XOR U5913 ( .A(n7363), .B(n7364), .Z(n4429) );
  NOR U5914 ( .A(n7365), .B(n7363), .Z(n7364) );
  XOR U5915 ( .A(n7366), .B(n7367), .Z(n4505) );
  NOR U5916 ( .A(n7368), .B(n7366), .Z(n7367) );
  XOR U5917 ( .A(n7369), .B(n7370), .Z(n4500) );
  NOR U5918 ( .A(n7371), .B(n7369), .Z(n7370) );
  XOR U5919 ( .A(n7372), .B(n7373), .Z(n4501) );
  NOR U5920 ( .A(n7374), .B(n7372), .Z(n7373) );
  XOR U5921 ( .A(n7375), .B(n7376), .Z(n4420) );
  NOR U5922 ( .A(n7377), .B(n7375), .Z(n7376) );
  XOR U5923 ( .A(n7378), .B(n7379), .Z(n4516) );
  NOR U5924 ( .A(n7380), .B(n7378), .Z(n7379) );
  XOR U5925 ( .A(n7381), .B(n7382), .Z(n4511) );
  NOR U5926 ( .A(n7383), .B(n7381), .Z(n7382) );
  XOR U5927 ( .A(n7384), .B(n7385), .Z(n4512) );
  NOR U5928 ( .A(n7386), .B(n7384), .Z(n7385) );
  XOR U5929 ( .A(n7387), .B(n7388), .Z(n4411) );
  NOR U5930 ( .A(n7389), .B(n7387), .Z(n7388) );
  XOR U5931 ( .A(n7390), .B(n7391), .Z(n4527) );
  NOR U5932 ( .A(n7392), .B(n7390), .Z(n7391) );
  XOR U5933 ( .A(n7393), .B(n7394), .Z(n4522) );
  NOR U5934 ( .A(n7395), .B(n7393), .Z(n7394) );
  XOR U5935 ( .A(n7396), .B(n7397), .Z(n4523) );
  NOR U5936 ( .A(n7398), .B(n7396), .Z(n7397) );
  XOR U5937 ( .A(n7399), .B(n7400), .Z(n4402) );
  NOR U5938 ( .A(n7401), .B(n7399), .Z(n7400) );
  XOR U5939 ( .A(n7402), .B(n7403), .Z(n4538) );
  NOR U5940 ( .A(n7404), .B(n7402), .Z(n7403) );
  XOR U5941 ( .A(n7405), .B(n7406), .Z(n4533) );
  NOR U5942 ( .A(n7407), .B(n7405), .Z(n7406) );
  XOR U5943 ( .A(n7408), .B(n7409), .Z(n4534) );
  NOR U5944 ( .A(n7410), .B(n7408), .Z(n7409) );
  XOR U5945 ( .A(n7411), .B(n7412), .Z(n4393) );
  NOR U5946 ( .A(n7413), .B(n7411), .Z(n7412) );
  XOR U5947 ( .A(n7414), .B(n7415), .Z(n4549) );
  NOR U5948 ( .A(n7416), .B(n7414), .Z(n7415) );
  XOR U5949 ( .A(n7417), .B(n7418), .Z(n4544) );
  NOR U5950 ( .A(n7419), .B(n7417), .Z(n7418) );
  XOR U5951 ( .A(n7420), .B(n7421), .Z(n4545) );
  NOR U5952 ( .A(n7422), .B(n7420), .Z(n7421) );
  XOR U5953 ( .A(n7423), .B(n7424), .Z(n4384) );
  NOR U5954 ( .A(n7425), .B(n7423), .Z(n7424) );
  XOR U5955 ( .A(n7426), .B(n7427), .Z(n4560) );
  NOR U5956 ( .A(n7428), .B(n7426), .Z(n7427) );
  XOR U5957 ( .A(n7429), .B(n7430), .Z(n4555) );
  NOR U5958 ( .A(n7431), .B(n7429), .Z(n7430) );
  XOR U5959 ( .A(n7432), .B(n7433), .Z(n4556) );
  NOR U5960 ( .A(n7434), .B(n7432), .Z(n7433) );
  XOR U5961 ( .A(n7435), .B(n7436), .Z(n4375) );
  NOR U5962 ( .A(n7437), .B(n7435), .Z(n7436) );
  XOR U5963 ( .A(n7438), .B(n7439), .Z(n4571) );
  NOR U5964 ( .A(n7440), .B(n7438), .Z(n7439) );
  XOR U5965 ( .A(n7441), .B(n7442), .Z(n4566) );
  NOR U5966 ( .A(n7443), .B(n7441), .Z(n7442) );
  XOR U5967 ( .A(n7444), .B(n7445), .Z(n4567) );
  NOR U5968 ( .A(n7446), .B(n7444), .Z(n7445) );
  XOR U5969 ( .A(n7447), .B(n7448), .Z(n4366) );
  NOR U5970 ( .A(n7449), .B(n7447), .Z(n7448) );
  XOR U5971 ( .A(n7450), .B(n7451), .Z(n4582) );
  NOR U5972 ( .A(n7452), .B(n7450), .Z(n7451) );
  XOR U5973 ( .A(n7453), .B(n7454), .Z(n4577) );
  NOR U5974 ( .A(n7455), .B(n7453), .Z(n7454) );
  XOR U5975 ( .A(n7456), .B(n7457), .Z(n4578) );
  NOR U5976 ( .A(n7458), .B(n7456), .Z(n7457) );
  XOR U5977 ( .A(n7459), .B(n7460), .Z(n4357) );
  NOR U5978 ( .A(n7461), .B(n7459), .Z(n7460) );
  XOR U5979 ( .A(n7462), .B(n7463), .Z(n4593) );
  NOR U5980 ( .A(n7464), .B(n7462), .Z(n7463) );
  XOR U5981 ( .A(n7465), .B(n7466), .Z(n4588) );
  NOR U5982 ( .A(n7467), .B(n7465), .Z(n7466) );
  XOR U5983 ( .A(n7468), .B(n7469), .Z(n4589) );
  NOR U5984 ( .A(n7470), .B(n7468), .Z(n7469) );
  XOR U5985 ( .A(n7471), .B(n7472), .Z(n4348) );
  NOR U5986 ( .A(n7473), .B(n7471), .Z(n7472) );
  XOR U5987 ( .A(n7474), .B(n7475), .Z(n4604) );
  NOR U5988 ( .A(n7476), .B(n7474), .Z(n7475) );
  XOR U5989 ( .A(n7477), .B(n7478), .Z(n4599) );
  NOR U5990 ( .A(n7479), .B(n7477), .Z(n7478) );
  XOR U5991 ( .A(n7480), .B(n7481), .Z(n4600) );
  NOR U5992 ( .A(n7482), .B(n7480), .Z(n7481) );
  XOR U5993 ( .A(n7483), .B(n7484), .Z(n4339) );
  NOR U5994 ( .A(n7485), .B(n7483), .Z(n7484) );
  XOR U5995 ( .A(n7486), .B(n7487), .Z(n4615) );
  NOR U5996 ( .A(n7488), .B(n7486), .Z(n7487) );
  XOR U5997 ( .A(n7489), .B(n7490), .Z(n4610) );
  NOR U5998 ( .A(n7491), .B(n7489), .Z(n7490) );
  XOR U5999 ( .A(n7492), .B(n7493), .Z(n4611) );
  NOR U6000 ( .A(n7494), .B(n7492), .Z(n7493) );
  XOR U6001 ( .A(n7495), .B(n7496), .Z(n4330) );
  NOR U6002 ( .A(n7497), .B(n7495), .Z(n7496) );
  XOR U6003 ( .A(n7498), .B(n7499), .Z(n4626) );
  NOR U6004 ( .A(n7500), .B(n7498), .Z(n7499) );
  XOR U6005 ( .A(n7501), .B(n7502), .Z(n4621) );
  NOR U6006 ( .A(n7503), .B(n7501), .Z(n7502) );
  XOR U6007 ( .A(n7504), .B(n7505), .Z(n4622) );
  NOR U6008 ( .A(n7506), .B(n7504), .Z(n7505) );
  XOR U6009 ( .A(n7507), .B(n7508), .Z(n4321) );
  NOR U6010 ( .A(n7509), .B(n7507), .Z(n7508) );
  XOR U6011 ( .A(n7510), .B(n7511), .Z(n4637) );
  NOR U6012 ( .A(n7512), .B(n7510), .Z(n7511) );
  XOR U6013 ( .A(n7513), .B(n7514), .Z(n4632) );
  NOR U6014 ( .A(n7515), .B(n7513), .Z(n7514) );
  XOR U6015 ( .A(n7516), .B(n7517), .Z(n4633) );
  NOR U6016 ( .A(n7518), .B(n7516), .Z(n7517) );
  XOR U6017 ( .A(n7519), .B(n7520), .Z(n4312) );
  NOR U6018 ( .A(n7521), .B(n7519), .Z(n7520) );
  XOR U6019 ( .A(n7522), .B(n7523), .Z(n4648) );
  NOR U6020 ( .A(n7524), .B(n7522), .Z(n7523) );
  XOR U6021 ( .A(n7525), .B(n7526), .Z(n4643) );
  NOR U6022 ( .A(n7527), .B(n7525), .Z(n7526) );
  XOR U6023 ( .A(n7528), .B(n7529), .Z(n4644) );
  NOR U6024 ( .A(n7530), .B(n7528), .Z(n7529) );
  XOR U6025 ( .A(n7531), .B(n7532), .Z(n4303) );
  NOR U6026 ( .A(n7533), .B(n7531), .Z(n7532) );
  XOR U6027 ( .A(n7534), .B(n7535), .Z(n4659) );
  NOR U6028 ( .A(n7536), .B(n7534), .Z(n7535) );
  XOR U6029 ( .A(n7537), .B(n7538), .Z(n4654) );
  NOR U6030 ( .A(n7539), .B(n7537), .Z(n7538) );
  XOR U6031 ( .A(n7540), .B(n7541), .Z(n4655) );
  NOR U6032 ( .A(n7542), .B(n7540), .Z(n7541) );
  XOR U6033 ( .A(n7543), .B(n7544), .Z(n4294) );
  NOR U6034 ( .A(n7545), .B(n7543), .Z(n7544) );
  XOR U6035 ( .A(n7546), .B(n7547), .Z(n4670) );
  NOR U6036 ( .A(n7548), .B(n7546), .Z(n7547) );
  XOR U6037 ( .A(n7549), .B(n7550), .Z(n4665) );
  NOR U6038 ( .A(n7551), .B(n7549), .Z(n7550) );
  XOR U6039 ( .A(n7552), .B(n7553), .Z(n4666) );
  NOR U6040 ( .A(n7554), .B(n7552), .Z(n7553) );
  XOR U6041 ( .A(n7555), .B(n7556), .Z(n4285) );
  NOR U6042 ( .A(n7557), .B(n7555), .Z(n7556) );
  XOR U6043 ( .A(n7558), .B(n7559), .Z(n4681) );
  NOR U6044 ( .A(n7560), .B(n7558), .Z(n7559) );
  XOR U6045 ( .A(n7561), .B(n7562), .Z(n4676) );
  NOR U6046 ( .A(n7563), .B(n7561), .Z(n7562) );
  XOR U6047 ( .A(n7564), .B(n7565), .Z(n4677) );
  NOR U6048 ( .A(n7566), .B(n7564), .Z(n7565) );
  XOR U6049 ( .A(n7567), .B(n7568), .Z(n4276) );
  NOR U6050 ( .A(n7569), .B(n7567), .Z(n7568) );
  XOR U6051 ( .A(n7570), .B(n7571), .Z(n4692) );
  NOR U6052 ( .A(n7572), .B(n7570), .Z(n7571) );
  XOR U6053 ( .A(n7573), .B(n7574), .Z(n4687) );
  NOR U6054 ( .A(n7575), .B(n7573), .Z(n7574) );
  XOR U6055 ( .A(n7576), .B(n7577), .Z(n4688) );
  NOR U6056 ( .A(n7578), .B(n7576), .Z(n7577) );
  XOR U6057 ( .A(n7579), .B(n7580), .Z(n4267) );
  NOR U6058 ( .A(n7581), .B(n7579), .Z(n7580) );
  XOR U6059 ( .A(n7582), .B(n7583), .Z(n4703) );
  NOR U6060 ( .A(n7584), .B(n7582), .Z(n7583) );
  XOR U6061 ( .A(n7585), .B(n7586), .Z(n4698) );
  NOR U6062 ( .A(n7587), .B(n7585), .Z(n7586) );
  XOR U6063 ( .A(n7588), .B(n7589), .Z(n4699) );
  NOR U6064 ( .A(n7590), .B(n7588), .Z(n7589) );
  XOR U6065 ( .A(n7591), .B(n7592), .Z(n4258) );
  NOR U6066 ( .A(n7593), .B(n7591), .Z(n7592) );
  XOR U6067 ( .A(n7594), .B(n7595), .Z(n4714) );
  NOR U6068 ( .A(n7596), .B(n7594), .Z(n7595) );
  XOR U6069 ( .A(n7597), .B(n7598), .Z(n4709) );
  NOR U6070 ( .A(n7599), .B(n7597), .Z(n7598) );
  XOR U6071 ( .A(n7600), .B(n7601), .Z(n4710) );
  NOR U6072 ( .A(n7602), .B(n7600), .Z(n7601) );
  XOR U6073 ( .A(n7603), .B(n7604), .Z(n4249) );
  NOR U6074 ( .A(n7605), .B(n7603), .Z(n7604) );
  XOR U6075 ( .A(n7606), .B(n7607), .Z(n4725) );
  NOR U6076 ( .A(n7608), .B(n7606), .Z(n7607) );
  XOR U6077 ( .A(n7609), .B(n7610), .Z(n4720) );
  NOR U6078 ( .A(n7611), .B(n7609), .Z(n7610) );
  XOR U6079 ( .A(n7612), .B(n7613), .Z(n4721) );
  NOR U6080 ( .A(n7614), .B(n7612), .Z(n7613) );
  XOR U6081 ( .A(n7615), .B(n7616), .Z(n4240) );
  NOR U6082 ( .A(n7617), .B(n7615), .Z(n7616) );
  XOR U6083 ( .A(n7618), .B(n7619), .Z(n4736) );
  NOR U6084 ( .A(n7620), .B(n7618), .Z(n7619) );
  XOR U6085 ( .A(n7621), .B(n7622), .Z(n4731) );
  NOR U6086 ( .A(n7623), .B(n7621), .Z(n7622) );
  XOR U6087 ( .A(n7624), .B(n7625), .Z(n4732) );
  NOR U6088 ( .A(n7626), .B(n7624), .Z(n7625) );
  XOR U6089 ( .A(n7627), .B(n7628), .Z(n4231) );
  NOR U6090 ( .A(n7629), .B(n7627), .Z(n7628) );
  XOR U6091 ( .A(n7630), .B(n7631), .Z(n4747) );
  NOR U6092 ( .A(n7632), .B(n7630), .Z(n7631) );
  XOR U6093 ( .A(n7633), .B(n7634), .Z(n4742) );
  NOR U6094 ( .A(n7635), .B(n7633), .Z(n7634) );
  XOR U6095 ( .A(n7636), .B(n7637), .Z(n4743) );
  NOR U6096 ( .A(n7638), .B(n7636), .Z(n7637) );
  XOR U6097 ( .A(n7639), .B(n7640), .Z(n4222) );
  NOR U6098 ( .A(n7641), .B(n7639), .Z(n7640) );
  XOR U6099 ( .A(n7642), .B(n7643), .Z(n4758) );
  NOR U6100 ( .A(n7644), .B(n7642), .Z(n7643) );
  XOR U6101 ( .A(n7645), .B(n7646), .Z(n4753) );
  NOR U6102 ( .A(n7647), .B(n7645), .Z(n7646) );
  XOR U6103 ( .A(n7648), .B(n7649), .Z(n4754) );
  NOR U6104 ( .A(n7650), .B(n7648), .Z(n7649) );
  XOR U6105 ( .A(n7651), .B(n7652), .Z(n4213) );
  NOR U6106 ( .A(n7653), .B(n7651), .Z(n7652) );
  XOR U6107 ( .A(n7654), .B(n7655), .Z(n4769) );
  NOR U6108 ( .A(n7656), .B(n7654), .Z(n7655) );
  XOR U6109 ( .A(n7657), .B(n7658), .Z(n4764) );
  NOR U6110 ( .A(n7659), .B(n7657), .Z(n7658) );
  XOR U6111 ( .A(n7660), .B(n7661), .Z(n4765) );
  NOR U6112 ( .A(n7662), .B(n7660), .Z(n7661) );
  XOR U6113 ( .A(n7663), .B(n7664), .Z(n4204) );
  NOR U6114 ( .A(n7665), .B(n7663), .Z(n7664) );
  XOR U6115 ( .A(n7666), .B(n7667), .Z(n4780) );
  NOR U6116 ( .A(n7668), .B(n7666), .Z(n7667) );
  XOR U6117 ( .A(n7669), .B(n7670), .Z(n4775) );
  NOR U6118 ( .A(n7671), .B(n7669), .Z(n7670) );
  XOR U6119 ( .A(n7672), .B(n7673), .Z(n4776) );
  NOR U6120 ( .A(n7674), .B(n7672), .Z(n7673) );
  XOR U6121 ( .A(n7675), .B(n7676), .Z(n4195) );
  NOR U6122 ( .A(n7677), .B(n7675), .Z(n7676) );
  XOR U6123 ( .A(n7678), .B(n7679), .Z(n4791) );
  NOR U6124 ( .A(n7680), .B(n7678), .Z(n7679) );
  XOR U6125 ( .A(n7681), .B(n7682), .Z(n4786) );
  NOR U6126 ( .A(n7683), .B(n7681), .Z(n7682) );
  XOR U6127 ( .A(n7684), .B(n7685), .Z(n4787) );
  NOR U6128 ( .A(n7686), .B(n7684), .Z(n7685) );
  XOR U6129 ( .A(n7687), .B(n7688), .Z(n4186) );
  NOR U6130 ( .A(n7689), .B(n7687), .Z(n7688) );
  XOR U6131 ( .A(n7690), .B(n7691), .Z(n4160) );
  NOR U6132 ( .A(n7692), .B(n7690), .Z(n7691) );
  XOR U6133 ( .A(n7693), .B(n7694), .Z(n4165) );
  NOR U6134 ( .A(n7695), .B(n7693), .Z(n7694) );
  IV U6135 ( .A(n4167), .Z(n7021) );
  XNOR U6136 ( .A(n7696), .B(n7697), .Z(n4167) );
  NOR U6137 ( .A(n7698), .B(n7696), .Z(n7697) );
  XOR U6138 ( .A(n7699), .B(n7700), .Z(n4177) );
  NOR U6139 ( .A(n7701), .B(n7699), .Z(n7700) );
  XOR U6140 ( .A(n7702), .B(n7703), .Z(n4797) );
  NOR U6141 ( .A(n7704), .B(n7702), .Z(n7703) );
  XOR U6142 ( .A(n7705), .B(n7706), .Z(n4800) );
  NOR U6143 ( .A(n7707), .B(n7705), .Z(n7706) );
  XOR U6144 ( .A(n7708), .B(n7709), .Z(n4803) );
  NOR U6145 ( .A(n7710), .B(n7708), .Z(n7709) );
  XOR U6146 ( .A(n7711), .B(n7712), .Z(n4806) );
  NOR U6147 ( .A(n7713), .B(n7711), .Z(n7712) );
  XOR U6148 ( .A(n7714), .B(n7715), .Z(n4809) );
  NOR U6149 ( .A(n7716), .B(n7714), .Z(n7715) );
  XOR U6150 ( .A(n7717), .B(n7718), .Z(n4812) );
  NOR U6151 ( .A(n7719), .B(n7717), .Z(n7718) );
  XOR U6152 ( .A(n7720), .B(n7721), .Z(n4815) );
  NOR U6153 ( .A(n7722), .B(n7720), .Z(n7721) );
  XOR U6154 ( .A(n7723), .B(n7724), .Z(n4818) );
  NOR U6155 ( .A(n7725), .B(n7723), .Z(n7724) );
  XOR U6156 ( .A(n7726), .B(n7727), .Z(n4821) );
  NOR U6157 ( .A(n7728), .B(n7726), .Z(n7727) );
  XOR U6158 ( .A(n7729), .B(n7730), .Z(n4824) );
  NOR U6159 ( .A(n7731), .B(n7729), .Z(n7730) );
  XOR U6160 ( .A(n7732), .B(n7733), .Z(n4827) );
  NOR U6161 ( .A(n7734), .B(n7732), .Z(n7733) );
  XOR U6162 ( .A(n7735), .B(n7736), .Z(n4830) );
  NOR U6163 ( .A(n7737), .B(n7735), .Z(n7736) );
  XOR U6164 ( .A(n7738), .B(n7739), .Z(n4833) );
  NOR U6165 ( .A(n7740), .B(n7738), .Z(n7739) );
  XOR U6166 ( .A(n7741), .B(n7742), .Z(n4836) );
  NOR U6167 ( .A(n7743), .B(n7741), .Z(n7742) );
  XOR U6168 ( .A(n7744), .B(n7745), .Z(n4839) );
  NOR U6169 ( .A(n7746), .B(n7744), .Z(n7745) );
  XOR U6170 ( .A(n7747), .B(n7748), .Z(n4842) );
  NOR U6171 ( .A(n7749), .B(n7747), .Z(n7748) );
  XOR U6172 ( .A(n7750), .B(n7751), .Z(n4845) );
  NOR U6173 ( .A(n7752), .B(n7750), .Z(n7751) );
  XOR U6174 ( .A(n7753), .B(n7754), .Z(n4848) );
  NOR U6175 ( .A(n7755), .B(n7753), .Z(n7754) );
  XOR U6176 ( .A(n7756), .B(n7757), .Z(n4851) );
  NOR U6177 ( .A(n7758), .B(n7756), .Z(n7757) );
  XOR U6178 ( .A(n7759), .B(n7760), .Z(n4854) );
  NOR U6179 ( .A(n7761), .B(n7759), .Z(n7760) );
  XOR U6180 ( .A(n7762), .B(n7763), .Z(n4857) );
  NOR U6181 ( .A(n7764), .B(n7762), .Z(n7763) );
  XOR U6182 ( .A(n7765), .B(n7766), .Z(n4860) );
  NOR U6183 ( .A(n7767), .B(n7765), .Z(n7766) );
  XOR U6184 ( .A(n7768), .B(n7769), .Z(n4863) );
  NOR U6185 ( .A(n7770), .B(n7768), .Z(n7769) );
  XOR U6186 ( .A(n7771), .B(n7772), .Z(n4866) );
  NOR U6187 ( .A(n7773), .B(n7771), .Z(n7772) );
  XOR U6188 ( .A(n7774), .B(n7775), .Z(n4869) );
  NOR U6189 ( .A(n7776), .B(n7774), .Z(n7775) );
  XOR U6190 ( .A(n7777), .B(n7778), .Z(n4872) );
  NOR U6191 ( .A(n7779), .B(n7777), .Z(n7778) );
  XOR U6192 ( .A(n7780), .B(n7781), .Z(n4875) );
  NOR U6193 ( .A(n7782), .B(n7780), .Z(n7781) );
  XOR U6194 ( .A(n7783), .B(n7784), .Z(n4878) );
  NOR U6195 ( .A(n7785), .B(n7783), .Z(n7784) );
  XOR U6196 ( .A(n7786), .B(n7787), .Z(n4881) );
  NOR U6197 ( .A(n7788), .B(n7786), .Z(n7787) );
  XOR U6198 ( .A(n7789), .B(n7790), .Z(n4884) );
  NOR U6199 ( .A(n7791), .B(n7789), .Z(n7790) );
  XOR U6200 ( .A(n7792), .B(n7793), .Z(n4887) );
  NOR U6201 ( .A(n7794), .B(n7792), .Z(n7793) );
  XOR U6202 ( .A(n7795), .B(n7796), .Z(n4890) );
  NOR U6203 ( .A(n7797), .B(n7795), .Z(n7796) );
  XOR U6204 ( .A(n7798), .B(n7799), .Z(n4893) );
  NOR U6205 ( .A(n7800), .B(n7798), .Z(n7799) );
  XOR U6206 ( .A(n7801), .B(n7802), .Z(n4896) );
  NOR U6207 ( .A(n7803), .B(n7801), .Z(n7802) );
  XOR U6208 ( .A(n7804), .B(n7805), .Z(n4899) );
  NOR U6209 ( .A(n7806), .B(n7804), .Z(n7805) );
  XOR U6210 ( .A(n7807), .B(n7808), .Z(n4902) );
  NOR U6211 ( .A(n7809), .B(n7807), .Z(n7808) );
  XOR U6212 ( .A(n7810), .B(n7811), .Z(n4905) );
  NOR U6213 ( .A(n7812), .B(n7810), .Z(n7811) );
  XOR U6214 ( .A(n7813), .B(n7814), .Z(n4908) );
  NOR U6215 ( .A(n7815), .B(n7813), .Z(n7814) );
  XOR U6216 ( .A(n7816), .B(n7817), .Z(n4911) );
  NOR U6217 ( .A(n7818), .B(n7816), .Z(n7817) );
  XOR U6218 ( .A(n7819), .B(n7820), .Z(n4914) );
  NOR U6219 ( .A(n7821), .B(n7819), .Z(n7820) );
  XOR U6220 ( .A(n7822), .B(n7823), .Z(n4917) );
  NOR U6221 ( .A(n7824), .B(n7822), .Z(n7823) );
  XOR U6222 ( .A(n7825), .B(n7826), .Z(n4920) );
  NOR U6223 ( .A(n7827), .B(n7825), .Z(n7826) );
  XOR U6224 ( .A(n7828), .B(n7829), .Z(n4923) );
  NOR U6225 ( .A(n7830), .B(n7828), .Z(n7829) );
  XOR U6226 ( .A(n7831), .B(n7832), .Z(n4926) );
  NOR U6227 ( .A(n7833), .B(n7831), .Z(n7832) );
  XOR U6228 ( .A(n7834), .B(n7835), .Z(n4929) );
  NOR U6229 ( .A(n7836), .B(n7834), .Z(n7835) );
  XOR U6230 ( .A(n7837), .B(n7838), .Z(n4932) );
  NOR U6231 ( .A(n7839), .B(n7837), .Z(n7838) );
  XOR U6232 ( .A(n7840), .B(n7841), .Z(n4935) );
  NOR U6233 ( .A(n7842), .B(n7840), .Z(n7841) );
  XOR U6234 ( .A(n7843), .B(n7844), .Z(n4938) );
  NOR U6235 ( .A(n7845), .B(n7843), .Z(n7844) );
  XOR U6236 ( .A(n7846), .B(n7847), .Z(n4941) );
  NOR U6237 ( .A(n7848), .B(n7846), .Z(n7847) );
  XOR U6238 ( .A(n7849), .B(n7850), .Z(n4944) );
  NOR U6239 ( .A(n7851), .B(n7849), .Z(n7850) );
  XOR U6240 ( .A(n7852), .B(n7853), .Z(n4947) );
  NOR U6241 ( .A(n7854), .B(n7852), .Z(n7853) );
  XOR U6242 ( .A(n7855), .B(n7856), .Z(n4950) );
  NOR U6243 ( .A(n7857), .B(n7855), .Z(n7856) );
  XOR U6244 ( .A(n7858), .B(n7859), .Z(n4953) );
  NOR U6245 ( .A(n7860), .B(n7858), .Z(n7859) );
  XOR U6246 ( .A(n7861), .B(n7862), .Z(n4956) );
  NOR U6247 ( .A(n7863), .B(n7861), .Z(n7862) );
  XOR U6248 ( .A(n7864), .B(n7865), .Z(n4959) );
  NOR U6249 ( .A(n7866), .B(n7864), .Z(n7865) );
  XOR U6250 ( .A(n7867), .B(n7868), .Z(n4962) );
  NOR U6251 ( .A(n7869), .B(n7867), .Z(n7868) );
  XOR U6252 ( .A(n7870), .B(n7871), .Z(n4965) );
  NOR U6253 ( .A(n7872), .B(n7870), .Z(n7871) );
  XOR U6254 ( .A(n7873), .B(n7874), .Z(n4968) );
  NOR U6255 ( .A(n7875), .B(n7873), .Z(n7874) );
  XOR U6256 ( .A(n7876), .B(n7877), .Z(n4971) );
  NOR U6257 ( .A(n7878), .B(n7876), .Z(n7877) );
  XOR U6258 ( .A(n7879), .B(n7880), .Z(n4974) );
  NOR U6259 ( .A(n7881), .B(n7879), .Z(n7880) );
  XOR U6260 ( .A(n7882), .B(n7883), .Z(n4977) );
  NOR U6261 ( .A(n7884), .B(n7882), .Z(n7883) );
  XOR U6262 ( .A(n7885), .B(n7886), .Z(n4980) );
  NOR U6263 ( .A(n7887), .B(n7885), .Z(n7886) );
  XOR U6264 ( .A(n7888), .B(n7889), .Z(n4983) );
  NOR U6265 ( .A(n7890), .B(n7888), .Z(n7889) );
  XOR U6266 ( .A(n7891), .B(n7892), .Z(n4986) );
  NOR U6267 ( .A(n7893), .B(n7891), .Z(n7892) );
  XOR U6268 ( .A(n7894), .B(n7895), .Z(n4989) );
  NOR U6269 ( .A(n7896), .B(n7894), .Z(n7895) );
  XOR U6270 ( .A(n7897), .B(n7898), .Z(n4992) );
  NOR U6271 ( .A(n7899), .B(n7897), .Z(n7898) );
  XOR U6272 ( .A(n7900), .B(n7901), .Z(n4995) );
  NOR U6273 ( .A(n7902), .B(n7900), .Z(n7901) );
  XOR U6274 ( .A(n7903), .B(n7904), .Z(n4998) );
  NOR U6275 ( .A(n7905), .B(n7903), .Z(n7904) );
  XOR U6276 ( .A(n7906), .B(n7907), .Z(n5001) );
  NOR U6277 ( .A(n7908), .B(n7906), .Z(n7907) );
  XOR U6278 ( .A(n7909), .B(n7910), .Z(n5004) );
  NOR U6279 ( .A(n7911), .B(n7909), .Z(n7910) );
  XOR U6280 ( .A(n7912), .B(n7913), .Z(n5007) );
  NOR U6281 ( .A(n7914), .B(n7912), .Z(n7913) );
  XOR U6282 ( .A(n7915), .B(n7916), .Z(n5010) );
  NOR U6283 ( .A(n7917), .B(n7915), .Z(n7916) );
  XOR U6284 ( .A(n7918), .B(n7919), .Z(n5013) );
  NOR U6285 ( .A(n7920), .B(n7918), .Z(n7919) );
  XOR U6286 ( .A(n7921), .B(n7922), .Z(n5016) );
  NOR U6287 ( .A(n7923), .B(n7921), .Z(n7922) );
  XOR U6288 ( .A(n7924), .B(n7925), .Z(n5019) );
  NOR U6289 ( .A(n7926), .B(n7924), .Z(n7925) );
  XOR U6290 ( .A(n7927), .B(n7928), .Z(n5022) );
  NOR U6291 ( .A(n7929), .B(n7927), .Z(n7928) );
  XOR U6292 ( .A(n7930), .B(n7931), .Z(n5025) );
  NOR U6293 ( .A(n7932), .B(n7930), .Z(n7931) );
  XOR U6294 ( .A(n7933), .B(n7934), .Z(n5028) );
  NOR U6295 ( .A(n7935), .B(n7933), .Z(n7934) );
  XOR U6296 ( .A(n7936), .B(n7937), .Z(n5031) );
  NOR U6297 ( .A(n7938), .B(n7936), .Z(n7937) );
  XOR U6298 ( .A(n7939), .B(n7940), .Z(n5034) );
  NOR U6299 ( .A(n7941), .B(n7939), .Z(n7940) );
  XOR U6300 ( .A(n7942), .B(n7943), .Z(n5037) );
  NOR U6301 ( .A(n7944), .B(n7942), .Z(n7943) );
  XOR U6302 ( .A(n7945), .B(n7946), .Z(n5040) );
  NOR U6303 ( .A(n7947), .B(n7945), .Z(n7946) );
  XOR U6304 ( .A(n7948), .B(n7949), .Z(n5043) );
  NOR U6305 ( .A(n7950), .B(n7948), .Z(n7949) );
  XOR U6306 ( .A(n7951), .B(n7952), .Z(n5046) );
  NOR U6307 ( .A(n7953), .B(n7951), .Z(n7952) );
  XOR U6308 ( .A(n7954), .B(n7955), .Z(n5049) );
  NOR U6309 ( .A(n7956), .B(n7954), .Z(n7955) );
  XOR U6310 ( .A(n7957), .B(n7958), .Z(n5052) );
  NOR U6311 ( .A(n7959), .B(n7957), .Z(n7958) );
  XOR U6312 ( .A(n7960), .B(n7961), .Z(n5055) );
  NOR U6313 ( .A(n7962), .B(n7960), .Z(n7961) );
  XOR U6314 ( .A(n7963), .B(n7964), .Z(n5058) );
  NOR U6315 ( .A(n7965), .B(n7963), .Z(n7964) );
  XOR U6316 ( .A(n7966), .B(n7967), .Z(n5061) );
  NOR U6317 ( .A(n7968), .B(n7966), .Z(n7967) );
  XOR U6318 ( .A(n7969), .B(n7970), .Z(n5064) );
  NOR U6319 ( .A(n7971), .B(n7969), .Z(n7970) );
  XOR U6320 ( .A(n7972), .B(n7973), .Z(n5067) );
  NOR U6321 ( .A(n7974), .B(n7972), .Z(n7973) );
  XOR U6322 ( .A(n7975), .B(n7976), .Z(n5070) );
  NOR U6323 ( .A(n7977), .B(n7975), .Z(n7976) );
  XOR U6324 ( .A(n7978), .B(n7979), .Z(n5073) );
  NOR U6325 ( .A(n7980), .B(n7978), .Z(n7979) );
  XOR U6326 ( .A(n7981), .B(n7982), .Z(n5076) );
  NOR U6327 ( .A(n7983), .B(n7981), .Z(n7982) );
  XOR U6328 ( .A(n7984), .B(n7985), .Z(n5079) );
  NOR U6329 ( .A(n7986), .B(n7984), .Z(n7985) );
  XOR U6330 ( .A(n7987), .B(n7988), .Z(n5082) );
  NOR U6331 ( .A(n7989), .B(n7987), .Z(n7988) );
  XOR U6332 ( .A(n7990), .B(n7991), .Z(n5085) );
  NOR U6333 ( .A(n7992), .B(n7990), .Z(n7991) );
  XOR U6334 ( .A(n7993), .B(n7994), .Z(n5088) );
  NOR U6335 ( .A(n7995), .B(n7993), .Z(n7994) );
  XOR U6336 ( .A(n7996), .B(n7997), .Z(n5091) );
  NOR U6337 ( .A(n7998), .B(n7996), .Z(n7997) );
  XOR U6338 ( .A(n7999), .B(n8000), .Z(n5094) );
  NOR U6339 ( .A(n8001), .B(n7999), .Z(n8000) );
  XOR U6340 ( .A(n8002), .B(n8003), .Z(n5097) );
  NOR U6341 ( .A(n8004), .B(n8002), .Z(n8003) );
  XOR U6342 ( .A(n8005), .B(n8006), .Z(n5100) );
  NOR U6343 ( .A(n8007), .B(n8005), .Z(n8006) );
  XOR U6344 ( .A(n8008), .B(n8009), .Z(n5103) );
  NOR U6345 ( .A(n8010), .B(n8008), .Z(n8009) );
  XOR U6346 ( .A(n8011), .B(n8012), .Z(n5106) );
  NOR U6347 ( .A(n8013), .B(n8011), .Z(n8012) );
  XOR U6348 ( .A(n8014), .B(n8015), .Z(n5109) );
  NOR U6349 ( .A(n8016), .B(n8014), .Z(n8015) );
  XOR U6350 ( .A(n8017), .B(n8018), .Z(n5112) );
  NOR U6351 ( .A(n8019), .B(n8017), .Z(n8018) );
  XOR U6352 ( .A(n8020), .B(n8021), .Z(n5115) );
  NOR U6353 ( .A(n8022), .B(n8020), .Z(n8021) );
  XOR U6354 ( .A(n8023), .B(n8024), .Z(n5118) );
  NOR U6355 ( .A(n8025), .B(n8023), .Z(n8024) );
  XOR U6356 ( .A(n8026), .B(n8027), .Z(n5121) );
  NOR U6357 ( .A(n8028), .B(n8026), .Z(n8027) );
  XOR U6358 ( .A(n8029), .B(n8030), .Z(n5124) );
  NOR U6359 ( .A(n8031), .B(n8029), .Z(n8030) );
  XOR U6360 ( .A(n8032), .B(n8033), .Z(n5127) );
  NOR U6361 ( .A(n8034), .B(n8032), .Z(n8033) );
  XOR U6362 ( .A(n8035), .B(n8036), .Z(n5130) );
  NOR U6363 ( .A(n8037), .B(n8035), .Z(n8036) );
  XOR U6364 ( .A(n8038), .B(n8039), .Z(n5133) );
  NOR U6365 ( .A(n8040), .B(n8038), .Z(n8039) );
  XOR U6366 ( .A(n8041), .B(n8042), .Z(n5136) );
  NOR U6367 ( .A(n8043), .B(n8041), .Z(n8042) );
  XOR U6368 ( .A(n8044), .B(n8045), .Z(n5139) );
  NOR U6369 ( .A(n8046), .B(n8044), .Z(n8045) );
  XOR U6370 ( .A(n8047), .B(n8048), .Z(n5142) );
  NOR U6371 ( .A(n8049), .B(n8047), .Z(n8048) );
  XOR U6372 ( .A(n8050), .B(n8051), .Z(n5145) );
  NOR U6373 ( .A(n8052), .B(n8050), .Z(n8051) );
  XOR U6374 ( .A(n8053), .B(n8054), .Z(n5148) );
  NOR U6375 ( .A(n8055), .B(n8053), .Z(n8054) );
  XOR U6376 ( .A(n8056), .B(n8057), .Z(n5151) );
  NOR U6377 ( .A(n8058), .B(n8056), .Z(n8057) );
  XOR U6378 ( .A(n8059), .B(n8060), .Z(n5154) );
  NOR U6379 ( .A(n8061), .B(n8059), .Z(n8060) );
  XOR U6380 ( .A(n8062), .B(n8063), .Z(n5157) );
  NOR U6381 ( .A(n8064), .B(n8062), .Z(n8063) );
  XOR U6382 ( .A(n8065), .B(n8066), .Z(n5160) );
  NOR U6383 ( .A(n8067), .B(n8065), .Z(n8066) );
  XOR U6384 ( .A(n8068), .B(n8069), .Z(n5163) );
  NOR U6385 ( .A(n8070), .B(n8068), .Z(n8069) );
  XOR U6386 ( .A(n8071), .B(n8072), .Z(n5166) );
  NOR U6387 ( .A(n8073), .B(n8071), .Z(n8072) );
  XOR U6388 ( .A(n8074), .B(n8075), .Z(n5169) );
  NOR U6389 ( .A(n8076), .B(n8074), .Z(n8075) );
  XOR U6390 ( .A(n8077), .B(n8078), .Z(n5172) );
  NOR U6391 ( .A(n8079), .B(n8077), .Z(n8078) );
  XOR U6392 ( .A(n8080), .B(n8081), .Z(n5175) );
  NOR U6393 ( .A(n8082), .B(n8080), .Z(n8081) );
  XOR U6394 ( .A(n8083), .B(n8084), .Z(n5178) );
  NOR U6395 ( .A(n8085), .B(n8083), .Z(n8084) );
  XOR U6396 ( .A(n8086), .B(n8087), .Z(n5181) );
  NOR U6397 ( .A(n8088), .B(n8086), .Z(n8087) );
  XOR U6398 ( .A(n8089), .B(n8090), .Z(n5184) );
  NOR U6399 ( .A(n8091), .B(n8089), .Z(n8090) );
  XOR U6400 ( .A(n8092), .B(n8093), .Z(n5187) );
  NOR U6401 ( .A(n8094), .B(n8092), .Z(n8093) );
  XOR U6402 ( .A(n8095), .B(n8096), .Z(n5190) );
  NOR U6403 ( .A(n8097), .B(n8095), .Z(n8096) );
  XOR U6404 ( .A(n8098), .B(n8099), .Z(n5193) );
  NOR U6405 ( .A(n8100), .B(n8098), .Z(n8099) );
  XOR U6406 ( .A(n8101), .B(n8102), .Z(n5196) );
  NOR U6407 ( .A(n8103), .B(n8101), .Z(n8102) );
  XOR U6408 ( .A(n8104), .B(n8105), .Z(n5199) );
  NOR U6409 ( .A(n8106), .B(n8104), .Z(n8105) );
  XOR U6410 ( .A(n8107), .B(n8108), .Z(n5202) );
  NOR U6411 ( .A(n8109), .B(n8107), .Z(n8108) );
  XOR U6412 ( .A(n8110), .B(n8111), .Z(n5205) );
  NOR U6413 ( .A(n8112), .B(n8110), .Z(n8111) );
  XOR U6414 ( .A(n8113), .B(n8114), .Z(n5208) );
  NOR U6415 ( .A(n8115), .B(n8113), .Z(n8114) );
  XOR U6416 ( .A(n8116), .B(n8117), .Z(n5211) );
  NOR U6417 ( .A(n8118), .B(n8116), .Z(n8117) );
  XOR U6418 ( .A(n8119), .B(n8120), .Z(n5214) );
  NOR U6419 ( .A(n8121), .B(n8119), .Z(n8120) );
  XOR U6420 ( .A(n8122), .B(n8123), .Z(n5217) );
  NOR U6421 ( .A(n8124), .B(n8122), .Z(n8123) );
  XOR U6422 ( .A(n8125), .B(n8126), .Z(n5220) );
  NOR U6423 ( .A(n8127), .B(n8125), .Z(n8126) );
  XOR U6424 ( .A(n8128), .B(n8129), .Z(n5223) );
  NOR U6425 ( .A(n8130), .B(n8128), .Z(n8129) );
  XOR U6426 ( .A(n8131), .B(n8132), .Z(n5226) );
  NOR U6427 ( .A(n8133), .B(n8131), .Z(n8132) );
  XOR U6428 ( .A(n8134), .B(n8135), .Z(n5229) );
  NOR U6429 ( .A(n8136), .B(n8134), .Z(n8135) );
  XOR U6430 ( .A(n8137), .B(n8138), .Z(n5232) );
  NOR U6431 ( .A(n8139), .B(n8137), .Z(n8138) );
  XOR U6432 ( .A(n8140), .B(n8141), .Z(n5235) );
  NOR U6433 ( .A(n8142), .B(n8140), .Z(n8141) );
  XOR U6434 ( .A(n8143), .B(n8144), .Z(n5238) );
  NOR U6435 ( .A(n8145), .B(n8143), .Z(n8144) );
  XOR U6436 ( .A(n8146), .B(n8147), .Z(n5241) );
  NOR U6437 ( .A(n8148), .B(n8146), .Z(n8147) );
  XOR U6438 ( .A(n8149), .B(n8150), .Z(n5244) );
  NOR U6439 ( .A(n8151), .B(n8149), .Z(n8150) );
  XOR U6440 ( .A(n8152), .B(n8153), .Z(n5247) );
  NOR U6441 ( .A(n8154), .B(n8152), .Z(n8153) );
  XOR U6442 ( .A(n8155), .B(n8156), .Z(n5250) );
  NOR U6443 ( .A(n8157), .B(n8155), .Z(n8156) );
  XOR U6444 ( .A(n8158), .B(n8159), .Z(n5253) );
  NOR U6445 ( .A(n8160), .B(n8158), .Z(n8159) );
  XOR U6446 ( .A(n8161), .B(n8162), .Z(n5256) );
  NOR U6447 ( .A(n8163), .B(n8161), .Z(n8162) );
  XOR U6448 ( .A(n8164), .B(n8165), .Z(n5259) );
  NOR U6449 ( .A(n8166), .B(n8164), .Z(n8165) );
  XOR U6450 ( .A(n8167), .B(n8168), .Z(n5262) );
  NOR U6451 ( .A(n8169), .B(n8167), .Z(n8168) );
  XOR U6452 ( .A(n8170), .B(n8171), .Z(n5265) );
  NOR U6453 ( .A(n8172), .B(n8170), .Z(n8171) );
  XOR U6454 ( .A(n8173), .B(n8174), .Z(n5268) );
  NOR U6455 ( .A(n8175), .B(n8173), .Z(n8174) );
  XOR U6456 ( .A(n8176), .B(n8177), .Z(n5271) );
  NOR U6457 ( .A(n8178), .B(n8176), .Z(n8177) );
  XOR U6458 ( .A(n8179), .B(n8180), .Z(n5274) );
  NOR U6459 ( .A(n8181), .B(n8179), .Z(n8180) );
  XOR U6460 ( .A(n8182), .B(n8183), .Z(n5277) );
  NOR U6461 ( .A(n8184), .B(n8182), .Z(n8183) );
  XOR U6462 ( .A(n8185), .B(n8186), .Z(n5280) );
  NOR U6463 ( .A(n8187), .B(n8185), .Z(n8186) );
  XOR U6464 ( .A(n8188), .B(n8189), .Z(n5283) );
  NOR U6465 ( .A(n8190), .B(n8188), .Z(n8189) );
  XOR U6466 ( .A(n8191), .B(n8192), .Z(n5286) );
  NOR U6467 ( .A(n8193), .B(n8191), .Z(n8192) );
  XOR U6468 ( .A(n8194), .B(n8195), .Z(n5289) );
  NOR U6469 ( .A(n8196), .B(n8194), .Z(n8195) );
  XOR U6470 ( .A(n8197), .B(n8198), .Z(n5292) );
  NOR U6471 ( .A(n8199), .B(n8197), .Z(n8198) );
  XOR U6472 ( .A(n8200), .B(n8201), .Z(n5295) );
  NOR U6473 ( .A(n8202), .B(n8200), .Z(n8201) );
  XOR U6474 ( .A(n8203), .B(n8204), .Z(n5298) );
  NOR U6475 ( .A(n8205), .B(n8203), .Z(n8204) );
  XOR U6476 ( .A(n8206), .B(n8207), .Z(n5301) );
  NOR U6477 ( .A(n8208), .B(n8206), .Z(n8207) );
  XOR U6478 ( .A(n8209), .B(n8210), .Z(n5304) );
  NOR U6479 ( .A(n8211), .B(n8209), .Z(n8210) );
  XOR U6480 ( .A(n8212), .B(n8213), .Z(n5307) );
  NOR U6481 ( .A(n8214), .B(n8212), .Z(n8213) );
  XOR U6482 ( .A(n8215), .B(n8216), .Z(n5310) );
  NOR U6483 ( .A(n8217), .B(n8215), .Z(n8216) );
  XOR U6484 ( .A(n8218), .B(n8219), .Z(n5313) );
  NOR U6485 ( .A(n8220), .B(n8218), .Z(n8219) );
  XOR U6486 ( .A(n8221), .B(n8222), .Z(n5316) );
  NOR U6487 ( .A(n8223), .B(n8221), .Z(n8222) );
  XOR U6488 ( .A(n8224), .B(n8225), .Z(n5319) );
  NOR U6489 ( .A(n8226), .B(n8224), .Z(n8225) );
  XOR U6490 ( .A(n8227), .B(n8228), .Z(n5322) );
  NOR U6491 ( .A(n8229), .B(n8227), .Z(n8228) );
  XOR U6492 ( .A(n8230), .B(n8231), .Z(n5325) );
  NOR U6493 ( .A(n8232), .B(n8230), .Z(n8231) );
  XOR U6494 ( .A(n8233), .B(n8234), .Z(n5328) );
  NOR U6495 ( .A(n8235), .B(n8233), .Z(n8234) );
  XOR U6496 ( .A(n8236), .B(n8237), .Z(n5331) );
  NOR U6497 ( .A(n8238), .B(n8236), .Z(n8237) );
  XOR U6498 ( .A(n8239), .B(n8240), .Z(n5334) );
  NOR U6499 ( .A(n8241), .B(n8239), .Z(n8240) );
  XOR U6500 ( .A(n8242), .B(n8243), .Z(n5337) );
  NOR U6501 ( .A(n8244), .B(n8242), .Z(n8243) );
  XOR U6502 ( .A(n8245), .B(n8246), .Z(n5340) );
  NOR U6503 ( .A(n8247), .B(n8245), .Z(n8246) );
  XOR U6504 ( .A(n8248), .B(n8249), .Z(n5343) );
  NOR U6505 ( .A(n8250), .B(n8248), .Z(n8249) );
  XOR U6506 ( .A(n8251), .B(n8252), .Z(n5346) );
  NOR U6507 ( .A(n8253), .B(n8251), .Z(n8252) );
  XOR U6508 ( .A(n8254), .B(n8255), .Z(n5349) );
  NOR U6509 ( .A(n8256), .B(n8254), .Z(n8255) );
  XOR U6510 ( .A(n8257), .B(n8258), .Z(n5352) );
  NOR U6511 ( .A(n8259), .B(n8257), .Z(n8258) );
  XOR U6512 ( .A(n8260), .B(n8261), .Z(n5355) );
  NOR U6513 ( .A(n8262), .B(n8260), .Z(n8261) );
  XOR U6514 ( .A(n8263), .B(n8264), .Z(n5358) );
  NOR U6515 ( .A(n8265), .B(n8263), .Z(n8264) );
  XOR U6516 ( .A(n8266), .B(n8267), .Z(n5361) );
  NOR U6517 ( .A(n8268), .B(n8266), .Z(n8267) );
  XOR U6518 ( .A(n8269), .B(n8270), .Z(n5364) );
  NOR U6519 ( .A(n8271), .B(n8269), .Z(n8270) );
  XOR U6520 ( .A(n8272), .B(n8273), .Z(n5367) );
  NOR U6521 ( .A(n8274), .B(n8272), .Z(n8273) );
  XOR U6522 ( .A(n8275), .B(n8276), .Z(n5370) );
  NOR U6523 ( .A(n8277), .B(n8275), .Z(n8276) );
  XOR U6524 ( .A(n8278), .B(n8279), .Z(n5373) );
  NOR U6525 ( .A(n8280), .B(n8278), .Z(n8279) );
  XOR U6526 ( .A(n8281), .B(n8282), .Z(n5376) );
  NOR U6527 ( .A(n8283), .B(n8281), .Z(n8282) );
  XOR U6528 ( .A(n8284), .B(n8285), .Z(n5379) );
  NOR U6529 ( .A(n8286), .B(n8284), .Z(n8285) );
  XOR U6530 ( .A(n8287), .B(n8288), .Z(n5382) );
  NOR U6531 ( .A(n8289), .B(n8287), .Z(n8288) );
  XOR U6532 ( .A(n8290), .B(n8291), .Z(n5385) );
  NOR U6533 ( .A(n8292), .B(n8290), .Z(n8291) );
  XOR U6534 ( .A(n8293), .B(n8294), .Z(n5388) );
  NOR U6535 ( .A(n8295), .B(n8293), .Z(n8294) );
  XOR U6536 ( .A(n8296), .B(n8297), .Z(n5391) );
  NOR U6537 ( .A(n8298), .B(n8296), .Z(n8297) );
  XOR U6538 ( .A(n8299), .B(n8300), .Z(n5394) );
  NOR U6539 ( .A(n8301), .B(n8299), .Z(n8300) );
  XOR U6540 ( .A(n8302), .B(n8303), .Z(n5397) );
  NOR U6541 ( .A(n8304), .B(n8302), .Z(n8303) );
  XOR U6542 ( .A(n8305), .B(n8306), .Z(n5400) );
  NOR U6543 ( .A(n8307), .B(n8305), .Z(n8306) );
  XOR U6544 ( .A(n8308), .B(n8309), .Z(n5403) );
  NOR U6545 ( .A(n8310), .B(n8308), .Z(n8309) );
  XOR U6546 ( .A(n8311), .B(n8312), .Z(n5406) );
  NOR U6547 ( .A(n8313), .B(n8311), .Z(n8312) );
  XOR U6548 ( .A(n8314), .B(n8315), .Z(n5409) );
  NOR U6549 ( .A(n8316), .B(n8314), .Z(n8315) );
  XOR U6550 ( .A(n8317), .B(n8318), .Z(n5412) );
  NOR U6551 ( .A(n8319), .B(n8317), .Z(n8318) );
  XOR U6552 ( .A(n8320), .B(n8321), .Z(n5415) );
  NOR U6553 ( .A(n8322), .B(n8320), .Z(n8321) );
  XOR U6554 ( .A(n8323), .B(n8324), .Z(n5418) );
  NOR U6555 ( .A(n8325), .B(n8323), .Z(n8324) );
  XOR U6556 ( .A(n8326), .B(n8327), .Z(n5421) );
  NOR U6557 ( .A(n8328), .B(n8326), .Z(n8327) );
  XOR U6558 ( .A(n8329), .B(n8330), .Z(n5424) );
  NOR U6559 ( .A(n8331), .B(n8329), .Z(n8330) );
  XOR U6560 ( .A(n8332), .B(n8333), .Z(n5427) );
  NOR U6561 ( .A(n8334), .B(n8332), .Z(n8333) );
  XOR U6562 ( .A(n8335), .B(n8336), .Z(n5430) );
  NOR U6563 ( .A(n8337), .B(n8335), .Z(n8336) );
  XOR U6564 ( .A(n8338), .B(n8339), .Z(n5433) );
  NOR U6565 ( .A(n8340), .B(n8338), .Z(n8339) );
  XOR U6566 ( .A(n8341), .B(n8342), .Z(n5436) );
  NOR U6567 ( .A(n8343), .B(n8341), .Z(n8342) );
  XOR U6568 ( .A(n8344), .B(n8345), .Z(n5439) );
  NOR U6569 ( .A(n8346), .B(n8344), .Z(n8345) );
  XOR U6570 ( .A(n8347), .B(n8348), .Z(n5442) );
  NOR U6571 ( .A(n8349), .B(n8347), .Z(n8348) );
  XOR U6572 ( .A(n8350), .B(n8351), .Z(n5445) );
  NOR U6573 ( .A(n8352), .B(n8350), .Z(n8351) );
  XOR U6574 ( .A(n8353), .B(n8354), .Z(n5448) );
  NOR U6575 ( .A(n8355), .B(n8353), .Z(n8354) );
  XOR U6576 ( .A(n8356), .B(n8357), .Z(n5451) );
  NOR U6577 ( .A(n8358), .B(n8356), .Z(n8357) );
  XOR U6578 ( .A(n8359), .B(n8360), .Z(n5454) );
  NOR U6579 ( .A(n8361), .B(n8359), .Z(n8360) );
  XOR U6580 ( .A(n8362), .B(n8363), .Z(n5457) );
  NOR U6581 ( .A(n8364), .B(n8362), .Z(n8363) );
  XOR U6582 ( .A(n8365), .B(n8366), .Z(n5460) );
  NOR U6583 ( .A(n8367), .B(n8365), .Z(n8366) );
  XOR U6584 ( .A(n8368), .B(n8369), .Z(n5463) );
  NOR U6585 ( .A(n8370), .B(n8368), .Z(n8369) );
  XOR U6586 ( .A(n8371), .B(n8372), .Z(n5466) );
  NOR U6587 ( .A(n8373), .B(n8371), .Z(n8372) );
  XOR U6588 ( .A(n8374), .B(n8375), .Z(n5469) );
  NOR U6589 ( .A(n8376), .B(n8374), .Z(n8375) );
  XOR U6590 ( .A(n8377), .B(n8378), .Z(n5472) );
  NOR U6591 ( .A(n8379), .B(n8377), .Z(n8378) );
  XOR U6592 ( .A(n8380), .B(n8381), .Z(n5475) );
  NOR U6593 ( .A(n8382), .B(n8380), .Z(n8381) );
  XOR U6594 ( .A(n8383), .B(n8384), .Z(n5478) );
  NOR U6595 ( .A(n8385), .B(n8383), .Z(n8384) );
  XOR U6596 ( .A(n8386), .B(n8387), .Z(n5481) );
  NOR U6597 ( .A(n8388), .B(n8386), .Z(n8387) );
  XOR U6598 ( .A(n8389), .B(n8390), .Z(n5484) );
  NOR U6599 ( .A(n8391), .B(n8389), .Z(n8390) );
  XOR U6600 ( .A(n8392), .B(n8393), .Z(n5487) );
  NOR U6601 ( .A(n8394), .B(n8392), .Z(n8393) );
  XOR U6602 ( .A(n8395), .B(n8396), .Z(n5490) );
  NOR U6603 ( .A(n8397), .B(n8395), .Z(n8396) );
  XOR U6604 ( .A(n8398), .B(n8399), .Z(n5493) );
  NOR U6605 ( .A(n8400), .B(n8398), .Z(n8399) );
  XOR U6606 ( .A(n8401), .B(n8402), .Z(n5496) );
  NOR U6607 ( .A(n8403), .B(n8401), .Z(n8402) );
  XOR U6608 ( .A(n8404), .B(n8405), .Z(n5499) );
  NOR U6609 ( .A(n8406), .B(n8404), .Z(n8405) );
  XOR U6610 ( .A(n8407), .B(n8408), .Z(n5502) );
  NOR U6611 ( .A(n8409), .B(n8407), .Z(n8408) );
  XOR U6612 ( .A(n8410), .B(n8411), .Z(n5505) );
  NOR U6613 ( .A(n8412), .B(n8410), .Z(n8411) );
  XOR U6614 ( .A(n8413), .B(n8414), .Z(n5508) );
  NOR U6615 ( .A(n8415), .B(n8413), .Z(n8414) );
  XOR U6616 ( .A(n8416), .B(n8417), .Z(n5511) );
  NOR U6617 ( .A(n8418), .B(n8416), .Z(n8417) );
  XOR U6618 ( .A(n8419), .B(n8420), .Z(n5514) );
  NOR U6619 ( .A(n8421), .B(n8419), .Z(n8420) );
  XOR U6620 ( .A(n8422), .B(n8423), .Z(n5517) );
  NOR U6621 ( .A(n8424), .B(n8422), .Z(n8423) );
  XOR U6622 ( .A(n8425), .B(n8426), .Z(n5520) );
  NOR U6623 ( .A(n8427), .B(n8425), .Z(n8426) );
  XOR U6624 ( .A(n8428), .B(n8429), .Z(n5523) );
  NOR U6625 ( .A(n8430), .B(n8428), .Z(n8429) );
  XOR U6626 ( .A(n8431), .B(n8432), .Z(n5526) );
  NOR U6627 ( .A(n8433), .B(n8431), .Z(n8432) );
  XOR U6628 ( .A(n8434), .B(n8435), .Z(n5529) );
  NOR U6629 ( .A(n8436), .B(n8434), .Z(n8435) );
  XOR U6630 ( .A(n8437), .B(n8438), .Z(n5532) );
  NOR U6631 ( .A(n8439), .B(n8437), .Z(n8438) );
  XOR U6632 ( .A(n8440), .B(n8441), .Z(n5535) );
  NOR U6633 ( .A(n8442), .B(n8440), .Z(n8441) );
  XOR U6634 ( .A(n8443), .B(n8444), .Z(n5538) );
  NOR U6635 ( .A(n8445), .B(n8443), .Z(n8444) );
  XOR U6636 ( .A(n8446), .B(n8447), .Z(n5541) );
  NOR U6637 ( .A(n8448), .B(n8446), .Z(n8447) );
  XOR U6638 ( .A(n8449), .B(n8450), .Z(n5544) );
  NOR U6639 ( .A(n8451), .B(n8449), .Z(n8450) );
  XOR U6640 ( .A(n8452), .B(n8453), .Z(n5547) );
  NOR U6641 ( .A(n8454), .B(n8452), .Z(n8453) );
  XOR U6642 ( .A(n8455), .B(n8456), .Z(n5550) );
  NOR U6643 ( .A(n8457), .B(n8455), .Z(n8456) );
  XOR U6644 ( .A(n8458), .B(n8459), .Z(n5553) );
  NOR U6645 ( .A(n8460), .B(n8458), .Z(n8459) );
  XOR U6646 ( .A(n8461), .B(n8462), .Z(n5556) );
  NOR U6647 ( .A(n8463), .B(n8461), .Z(n8462) );
  XOR U6648 ( .A(n8464), .B(n8465), .Z(n5559) );
  NOR U6649 ( .A(n8466), .B(n8464), .Z(n8465) );
  XOR U6650 ( .A(n8467), .B(n8468), .Z(n5562) );
  NOR U6651 ( .A(n8469), .B(n8467), .Z(n8468) );
  XOR U6652 ( .A(n8470), .B(n8471), .Z(n5565) );
  NOR U6653 ( .A(n72), .B(n8472), .Z(n8471) );
  IV U6654 ( .A(n8470), .Z(n8472) );
  XOR U6655 ( .A(n8473), .B(n8474), .Z(n5568) );
  AND U6656 ( .A(n8475), .B(n8476), .Z(n8474) );
  XOR U6657 ( .A(n8473), .B(n74), .Z(n8476) );
  XOR U6658 ( .A(n7019), .B(n7018), .Z(n74) );
  XNOR U6659 ( .A(n7016), .B(n7015), .Z(n7018) );
  XNOR U6660 ( .A(n7013), .B(n7012), .Z(n7015) );
  XNOR U6661 ( .A(n7010), .B(n7009), .Z(n7012) );
  XNOR U6662 ( .A(n7007), .B(n7006), .Z(n7009) );
  XNOR U6663 ( .A(n7004), .B(n7003), .Z(n7006) );
  XNOR U6664 ( .A(n7001), .B(n7000), .Z(n7003) );
  XNOR U6665 ( .A(n6998), .B(n6997), .Z(n7000) );
  XNOR U6666 ( .A(n6995), .B(n6994), .Z(n6997) );
  XNOR U6667 ( .A(n6992), .B(n6991), .Z(n6994) );
  XNOR U6668 ( .A(n6989), .B(n6988), .Z(n6991) );
  XNOR U6669 ( .A(n6986), .B(n6985), .Z(n6988) );
  XNOR U6670 ( .A(n6983), .B(n6982), .Z(n6985) );
  XNOR U6671 ( .A(n6980), .B(n6979), .Z(n6982) );
  XNOR U6672 ( .A(n6977), .B(n6976), .Z(n6979) );
  XNOR U6673 ( .A(n6974), .B(n6973), .Z(n6976) );
  XNOR U6674 ( .A(n6971), .B(n6970), .Z(n6973) );
  XNOR U6675 ( .A(n6968), .B(n6967), .Z(n6970) );
  XNOR U6676 ( .A(n6965), .B(n6964), .Z(n6967) );
  XNOR U6677 ( .A(n6962), .B(n6961), .Z(n6964) );
  XNOR U6678 ( .A(n6959), .B(n6958), .Z(n6961) );
  XNOR U6679 ( .A(n6956), .B(n6955), .Z(n6958) );
  XNOR U6680 ( .A(n6953), .B(n6952), .Z(n6955) );
  XNOR U6681 ( .A(n6950), .B(n6949), .Z(n6952) );
  XNOR U6682 ( .A(n6947), .B(n6946), .Z(n6949) );
  XNOR U6683 ( .A(n6944), .B(n6943), .Z(n6946) );
  XNOR U6684 ( .A(n6941), .B(n6940), .Z(n6943) );
  XNOR U6685 ( .A(n6938), .B(n6937), .Z(n6940) );
  XNOR U6686 ( .A(n6935), .B(n6934), .Z(n6937) );
  XNOR U6687 ( .A(n6932), .B(n6931), .Z(n6934) );
  XNOR U6688 ( .A(n6929), .B(n6928), .Z(n6931) );
  XNOR U6689 ( .A(n6926), .B(n6925), .Z(n6928) );
  XNOR U6690 ( .A(n6923), .B(n6922), .Z(n6925) );
  XNOR U6691 ( .A(n6920), .B(n6919), .Z(n6922) );
  XNOR U6692 ( .A(n6917), .B(n6916), .Z(n6919) );
  XNOR U6693 ( .A(n6914), .B(n6913), .Z(n6916) );
  XNOR U6694 ( .A(n6911), .B(n6910), .Z(n6913) );
  XNOR U6695 ( .A(n6908), .B(n6907), .Z(n6910) );
  XNOR U6696 ( .A(n6905), .B(n6904), .Z(n6907) );
  XNOR U6697 ( .A(n6902), .B(n6901), .Z(n6904) );
  XNOR U6698 ( .A(n6899), .B(n6898), .Z(n6901) );
  XNOR U6699 ( .A(n6896), .B(n6895), .Z(n6898) );
  XNOR U6700 ( .A(n6893), .B(n6892), .Z(n6895) );
  XNOR U6701 ( .A(n6890), .B(n6889), .Z(n6892) );
  XNOR U6702 ( .A(n6887), .B(n6886), .Z(n6889) );
  XNOR U6703 ( .A(n6884), .B(n6883), .Z(n6886) );
  XNOR U6704 ( .A(n6881), .B(n6880), .Z(n6883) );
  XNOR U6705 ( .A(n6878), .B(n6877), .Z(n6880) );
  XNOR U6706 ( .A(n6875), .B(n6874), .Z(n6877) );
  XNOR U6707 ( .A(n6872), .B(n6871), .Z(n6874) );
  XNOR U6708 ( .A(n6869), .B(n6868), .Z(n6871) );
  XNOR U6709 ( .A(n6866), .B(n6865), .Z(n6868) );
  XNOR U6710 ( .A(n6863), .B(n6862), .Z(n6865) );
  XNOR U6711 ( .A(n6860), .B(n6859), .Z(n6862) );
  XNOR U6712 ( .A(n6857), .B(n6856), .Z(n6859) );
  XNOR U6713 ( .A(n6854), .B(n6853), .Z(n6856) );
  XNOR U6714 ( .A(n6851), .B(n6850), .Z(n6853) );
  XNOR U6715 ( .A(n6848), .B(n6847), .Z(n6850) );
  XNOR U6716 ( .A(n6845), .B(n6844), .Z(n6847) );
  XNOR U6717 ( .A(n6842), .B(n6841), .Z(n6844) );
  XNOR U6718 ( .A(n6839), .B(n6838), .Z(n6841) );
  XNOR U6719 ( .A(n6836), .B(n6835), .Z(n6838) );
  XNOR U6720 ( .A(n6833), .B(n6832), .Z(n6835) );
  XNOR U6721 ( .A(n6830), .B(n6829), .Z(n6832) );
  XNOR U6722 ( .A(n6827), .B(n6826), .Z(n6829) );
  XNOR U6723 ( .A(n6824), .B(n6823), .Z(n6826) );
  XNOR U6724 ( .A(n6821), .B(n6820), .Z(n6823) );
  XNOR U6725 ( .A(n6818), .B(n6817), .Z(n6820) );
  XNOR U6726 ( .A(n6815), .B(n6814), .Z(n6817) );
  XNOR U6727 ( .A(n6812), .B(n6811), .Z(n6814) );
  XNOR U6728 ( .A(n6809), .B(n6808), .Z(n6811) );
  XNOR U6729 ( .A(n6806), .B(n6805), .Z(n6808) );
  XNOR U6730 ( .A(n6803), .B(n6802), .Z(n6805) );
  XNOR U6731 ( .A(n6800), .B(n6799), .Z(n6802) );
  XNOR U6732 ( .A(n6797), .B(n6796), .Z(n6799) );
  XNOR U6733 ( .A(n6794), .B(n6793), .Z(n6796) );
  XNOR U6734 ( .A(n6791), .B(n6790), .Z(n6793) );
  XNOR U6735 ( .A(n6788), .B(n6787), .Z(n6790) );
  XNOR U6736 ( .A(n6785), .B(n6784), .Z(n6787) );
  XNOR U6737 ( .A(n6782), .B(n6781), .Z(n6784) );
  XNOR U6738 ( .A(n6779), .B(n6778), .Z(n6781) );
  XNOR U6739 ( .A(n6776), .B(n6775), .Z(n6778) );
  XNOR U6740 ( .A(n6773), .B(n6772), .Z(n6775) );
  XNOR U6741 ( .A(n6770), .B(n6769), .Z(n6772) );
  XNOR U6742 ( .A(n6767), .B(n6766), .Z(n6769) );
  XNOR U6743 ( .A(n6764), .B(n6763), .Z(n6766) );
  XNOR U6744 ( .A(n6761), .B(n6760), .Z(n6763) );
  XNOR U6745 ( .A(n6758), .B(n6757), .Z(n6760) );
  XNOR U6746 ( .A(n6755), .B(n6754), .Z(n6757) );
  XNOR U6747 ( .A(n6752), .B(n6751), .Z(n6754) );
  XNOR U6748 ( .A(n6749), .B(n6748), .Z(n6751) );
  XNOR U6749 ( .A(n6746), .B(n6745), .Z(n6748) );
  XNOR U6750 ( .A(n6743), .B(n6742), .Z(n6745) );
  XNOR U6751 ( .A(n6740), .B(n6739), .Z(n6742) );
  XNOR U6752 ( .A(n6737), .B(n6736), .Z(n6739) );
  XNOR U6753 ( .A(n6734), .B(n6733), .Z(n6736) );
  XNOR U6754 ( .A(n6731), .B(n6730), .Z(n6733) );
  XNOR U6755 ( .A(n6728), .B(n6727), .Z(n6730) );
  XNOR U6756 ( .A(n6725), .B(n6724), .Z(n6727) );
  XNOR U6757 ( .A(n6722), .B(n6721), .Z(n6724) );
  XNOR U6758 ( .A(n6719), .B(n6718), .Z(n6721) );
  XNOR U6759 ( .A(n6716), .B(n6715), .Z(n6718) );
  XNOR U6760 ( .A(n6713), .B(n6712), .Z(n6715) );
  XNOR U6761 ( .A(n6710), .B(n6709), .Z(n6712) );
  XNOR U6762 ( .A(n6707), .B(n6706), .Z(n6709) );
  XNOR U6763 ( .A(n6704), .B(n6703), .Z(n6706) );
  XNOR U6764 ( .A(n6701), .B(n6700), .Z(n6703) );
  XNOR U6765 ( .A(n6698), .B(n6697), .Z(n6700) );
  XNOR U6766 ( .A(n6695), .B(n6694), .Z(n6697) );
  XNOR U6767 ( .A(n6692), .B(n6691), .Z(n6694) );
  XNOR U6768 ( .A(n6689), .B(n6688), .Z(n6691) );
  XNOR U6769 ( .A(n6686), .B(n6685), .Z(n6688) );
  XNOR U6770 ( .A(n6683), .B(n6682), .Z(n6685) );
  XNOR U6771 ( .A(n6680), .B(n6679), .Z(n6682) );
  XNOR U6772 ( .A(n6677), .B(n6676), .Z(n6679) );
  XNOR U6773 ( .A(n6674), .B(n6673), .Z(n6676) );
  XNOR U6774 ( .A(n6671), .B(n6670), .Z(n6673) );
  XNOR U6775 ( .A(n6668), .B(n6667), .Z(n6670) );
  XNOR U6776 ( .A(n6665), .B(n6664), .Z(n6667) );
  XNOR U6777 ( .A(n6662), .B(n6661), .Z(n6664) );
  XNOR U6778 ( .A(n6659), .B(n6658), .Z(n6661) );
  XNOR U6779 ( .A(n6656), .B(n6655), .Z(n6658) );
  XNOR U6780 ( .A(n6653), .B(n6652), .Z(n6655) );
  XNOR U6781 ( .A(n6650), .B(n6649), .Z(n6652) );
  XNOR U6782 ( .A(n6647), .B(n6646), .Z(n6649) );
  XNOR U6783 ( .A(n6644), .B(n6643), .Z(n6646) );
  XNOR U6784 ( .A(n6641), .B(n6640), .Z(n6643) );
  XNOR U6785 ( .A(n6638), .B(n6637), .Z(n6640) );
  XNOR U6786 ( .A(n6635), .B(n6634), .Z(n6637) );
  XNOR U6787 ( .A(n6632), .B(n6631), .Z(n6634) );
  XNOR U6788 ( .A(n6629), .B(n6628), .Z(n6631) );
  XNOR U6789 ( .A(n6626), .B(n6625), .Z(n6628) );
  XNOR U6790 ( .A(n6623), .B(n6622), .Z(n6625) );
  XNOR U6791 ( .A(n6620), .B(n6619), .Z(n6622) );
  XNOR U6792 ( .A(n6617), .B(n6616), .Z(n6619) );
  XNOR U6793 ( .A(n6614), .B(n6613), .Z(n6616) );
  XNOR U6794 ( .A(n6611), .B(n6610), .Z(n6613) );
  XNOR U6795 ( .A(n6608), .B(n6607), .Z(n6610) );
  XNOR U6796 ( .A(n6605), .B(n6604), .Z(n6607) );
  XNOR U6797 ( .A(n6602), .B(n6601), .Z(n6604) );
  XNOR U6798 ( .A(n6599), .B(n6598), .Z(n6601) );
  XNOR U6799 ( .A(n6596), .B(n6595), .Z(n6598) );
  XNOR U6800 ( .A(n6593), .B(n6592), .Z(n6595) );
  XNOR U6801 ( .A(n6590), .B(n6589), .Z(n6592) );
  XNOR U6802 ( .A(n6587), .B(n6586), .Z(n6589) );
  XNOR U6803 ( .A(n6584), .B(n6583), .Z(n6586) );
  XNOR U6804 ( .A(n6581), .B(n6580), .Z(n6583) );
  XNOR U6805 ( .A(n6578), .B(n6577), .Z(n6580) );
  XNOR U6806 ( .A(n6575), .B(n6574), .Z(n6577) );
  XNOR U6807 ( .A(n6572), .B(n6571), .Z(n6574) );
  XNOR U6808 ( .A(n6569), .B(n6568), .Z(n6571) );
  XNOR U6809 ( .A(n6566), .B(n6565), .Z(n6568) );
  XNOR U6810 ( .A(n6563), .B(n6562), .Z(n6565) );
  XNOR U6811 ( .A(n6560), .B(n6559), .Z(n6562) );
  XNOR U6812 ( .A(n6557), .B(n6556), .Z(n6559) );
  XNOR U6813 ( .A(n6554), .B(n6553), .Z(n6556) );
  XNOR U6814 ( .A(n6551), .B(n6550), .Z(n6553) );
  XNOR U6815 ( .A(n6548), .B(n6547), .Z(n6550) );
  XNOR U6816 ( .A(n6545), .B(n6544), .Z(n6547) );
  XNOR U6817 ( .A(n6542), .B(n6541), .Z(n6544) );
  XNOR U6818 ( .A(n6539), .B(n6538), .Z(n6541) );
  XNOR U6819 ( .A(n6536), .B(n6535), .Z(n6538) );
  XNOR U6820 ( .A(n6533), .B(n6532), .Z(n6535) );
  XNOR U6821 ( .A(n6530), .B(n6529), .Z(n6532) );
  XNOR U6822 ( .A(n6527), .B(n6526), .Z(n6529) );
  XNOR U6823 ( .A(n6524), .B(n6523), .Z(n6526) );
  XNOR U6824 ( .A(n6521), .B(n6520), .Z(n6523) );
  XNOR U6825 ( .A(n6518), .B(n6517), .Z(n6520) );
  XNOR U6826 ( .A(n6515), .B(n6514), .Z(n6517) );
  XNOR U6827 ( .A(n6512), .B(n6511), .Z(n6514) );
  XNOR U6828 ( .A(n6509), .B(n6508), .Z(n6511) );
  XNOR U6829 ( .A(n6506), .B(n6505), .Z(n6508) );
  XNOR U6830 ( .A(n6503), .B(n6502), .Z(n6505) );
  XNOR U6831 ( .A(n6500), .B(n6499), .Z(n6502) );
  XNOR U6832 ( .A(n6497), .B(n6496), .Z(n6499) );
  XNOR U6833 ( .A(n6494), .B(n6493), .Z(n6496) );
  XNOR U6834 ( .A(n6491), .B(n6490), .Z(n6493) );
  XNOR U6835 ( .A(n6488), .B(n6487), .Z(n6490) );
  XNOR U6836 ( .A(n6485), .B(n6484), .Z(n6487) );
  XNOR U6837 ( .A(n6482), .B(n6481), .Z(n6484) );
  XNOR U6838 ( .A(n6479), .B(n6478), .Z(n6481) );
  XNOR U6839 ( .A(n6476), .B(n6475), .Z(n6478) );
  XNOR U6840 ( .A(n6473), .B(n6472), .Z(n6475) );
  XNOR U6841 ( .A(n6470), .B(n6469), .Z(n6472) );
  XNOR U6842 ( .A(n6467), .B(n6466), .Z(n6469) );
  XNOR U6843 ( .A(n6464), .B(n6463), .Z(n6466) );
  XNOR U6844 ( .A(n6461), .B(n6460), .Z(n6463) );
  XNOR U6845 ( .A(n6458), .B(n6457), .Z(n6460) );
  XNOR U6846 ( .A(n6455), .B(n6454), .Z(n6457) );
  XNOR U6847 ( .A(n6452), .B(n6451), .Z(n6454) );
  XNOR U6848 ( .A(n6449), .B(n6448), .Z(n6451) );
  XNOR U6849 ( .A(n6446), .B(n6445), .Z(n6448) );
  XNOR U6850 ( .A(n6443), .B(n6442), .Z(n6445) );
  XNOR U6851 ( .A(n6440), .B(n6439), .Z(n6442) );
  XNOR U6852 ( .A(n6437), .B(n6436), .Z(n6439) );
  XNOR U6853 ( .A(n6434), .B(n6433), .Z(n6436) );
  XNOR U6854 ( .A(n6431), .B(n6430), .Z(n6433) );
  XNOR U6855 ( .A(n6428), .B(n6427), .Z(n6430) );
  XNOR U6856 ( .A(n6425), .B(n6424), .Z(n6427) );
  XNOR U6857 ( .A(n6422), .B(n6421), .Z(n6424) );
  XNOR U6858 ( .A(n6419), .B(n6418), .Z(n6421) );
  XNOR U6859 ( .A(n6416), .B(n6415), .Z(n6418) );
  XNOR U6860 ( .A(n6413), .B(n6412), .Z(n6415) );
  XNOR U6861 ( .A(n6410), .B(n6409), .Z(n6412) );
  XNOR U6862 ( .A(n6407), .B(n6406), .Z(n6409) );
  XNOR U6863 ( .A(n6404), .B(n6403), .Z(n6406) );
  XNOR U6864 ( .A(n6401), .B(n6400), .Z(n6403) );
  XNOR U6865 ( .A(n6398), .B(n6397), .Z(n6400) );
  XNOR U6866 ( .A(n6395), .B(n6394), .Z(n6397) );
  XNOR U6867 ( .A(n6392), .B(n6391), .Z(n6394) );
  XNOR U6868 ( .A(n6389), .B(n6388), .Z(n6391) );
  XNOR U6869 ( .A(n6386), .B(n6385), .Z(n6388) );
  XNOR U6870 ( .A(n6383), .B(n6382), .Z(n6385) );
  XNOR U6871 ( .A(n6380), .B(n6379), .Z(n6382) );
  XNOR U6872 ( .A(n6377), .B(n6376), .Z(n6379) );
  XNOR U6873 ( .A(n6374), .B(n6373), .Z(n6376) );
  XNOR U6874 ( .A(n6371), .B(n6370), .Z(n6373) );
  XNOR U6875 ( .A(n6368), .B(n6367), .Z(n6370) );
  XNOR U6876 ( .A(n6365), .B(n6364), .Z(n6367) );
  XNOR U6877 ( .A(n6362), .B(n6361), .Z(n6364) );
  XNOR U6878 ( .A(n6359), .B(n6358), .Z(n6361) );
  XNOR U6879 ( .A(n6356), .B(n6355), .Z(n6358) );
  XNOR U6880 ( .A(n6353), .B(n6352), .Z(n6355) );
  XNOR U6881 ( .A(n6350), .B(n6349), .Z(n6352) );
  XNOR U6882 ( .A(n6347), .B(n6346), .Z(n6349) );
  XNOR U6883 ( .A(n6344), .B(n6343), .Z(n6346) );
  XNOR U6884 ( .A(n6341), .B(n6340), .Z(n6343) );
  XNOR U6885 ( .A(n6338), .B(n6337), .Z(n6340) );
  XNOR U6886 ( .A(n6335), .B(n6334), .Z(n6337) );
  XNOR U6887 ( .A(n6332), .B(n6331), .Z(n6334) );
  XNOR U6888 ( .A(n6329), .B(n6328), .Z(n6331) );
  XNOR U6889 ( .A(n6326), .B(n6325), .Z(n6328) );
  XNOR U6890 ( .A(n6323), .B(n6322), .Z(n6325) );
  XNOR U6891 ( .A(n6320), .B(n6319), .Z(n6322) );
  XNOR U6892 ( .A(n6317), .B(n6316), .Z(n6319) );
  XNOR U6893 ( .A(n6314), .B(n6313), .Z(n6316) );
  XNOR U6894 ( .A(n6311), .B(n6310), .Z(n6313) );
  XNOR U6895 ( .A(n6308), .B(n6307), .Z(n6310) );
  XNOR U6896 ( .A(n6305), .B(n6304), .Z(n6307) );
  XNOR U6897 ( .A(n6302), .B(n6301), .Z(n6304) );
  XNOR U6898 ( .A(n6299), .B(n6298), .Z(n6301) );
  XNOR U6899 ( .A(n6296), .B(n6295), .Z(n6298) );
  XNOR U6900 ( .A(n6293), .B(n6292), .Z(n6295) );
  XNOR U6901 ( .A(n6290), .B(n6289), .Z(n6292) );
  XNOR U6902 ( .A(n6287), .B(n6286), .Z(n6289) );
  XNOR U6903 ( .A(n6284), .B(n6283), .Z(n6286) );
  XNOR U6904 ( .A(n6281), .B(n6280), .Z(n6283) );
  XNOR U6905 ( .A(n6278), .B(n6277), .Z(n6280) );
  XNOR U6906 ( .A(n6275), .B(n6274), .Z(n6277) );
  XNOR U6907 ( .A(n6272), .B(n6271), .Z(n6274) );
  XNOR U6908 ( .A(n6269), .B(n6268), .Z(n6271) );
  XNOR U6909 ( .A(n6266), .B(n6265), .Z(n6268) );
  XNOR U6910 ( .A(n6263), .B(n6262), .Z(n6265) );
  XNOR U6911 ( .A(n6260), .B(n6259), .Z(n6262) );
  XNOR U6912 ( .A(n6257), .B(n6256), .Z(n6259) );
  XNOR U6913 ( .A(n6254), .B(n6253), .Z(n6256) );
  XNOR U6914 ( .A(n6251), .B(n6250), .Z(n6253) );
  XNOR U6915 ( .A(n6248), .B(n6247), .Z(n6250) );
  XNOR U6916 ( .A(n6245), .B(n6244), .Z(n6247) );
  XNOR U6917 ( .A(n6242), .B(n6241), .Z(n6244) );
  XNOR U6918 ( .A(n6239), .B(n6238), .Z(n6241) );
  XNOR U6919 ( .A(n6236), .B(n6235), .Z(n6238) );
  XNOR U6920 ( .A(n6233), .B(n6232), .Z(n6235) );
  XNOR U6921 ( .A(n6230), .B(n6229), .Z(n6232) );
  XNOR U6922 ( .A(n6227), .B(n6226), .Z(n6229) );
  XNOR U6923 ( .A(n6224), .B(n6223), .Z(n6226) );
  XNOR U6924 ( .A(n6221), .B(n6220), .Z(n6223) );
  XNOR U6925 ( .A(n6218), .B(n6217), .Z(n6220) );
  XNOR U6926 ( .A(n6215), .B(n6214), .Z(n6217) );
  XNOR U6927 ( .A(n6212), .B(n6211), .Z(n6214) );
  XNOR U6928 ( .A(n6209), .B(n6208), .Z(n6211) );
  XNOR U6929 ( .A(n6206), .B(n6205), .Z(n6208) );
  XNOR U6930 ( .A(n6203), .B(n6202), .Z(n6205) );
  XNOR U6931 ( .A(n6200), .B(n6199), .Z(n6202) );
  XNOR U6932 ( .A(n6197), .B(n6196), .Z(n6199) );
  XNOR U6933 ( .A(n6194), .B(n6193), .Z(n6196) );
  XNOR U6934 ( .A(n6191), .B(n6190), .Z(n6193) );
  XNOR U6935 ( .A(n6188), .B(n6187), .Z(n6190) );
  XNOR U6936 ( .A(n6185), .B(n6184), .Z(n6187) );
  XNOR U6937 ( .A(n6182), .B(n6181), .Z(n6184) );
  XNOR U6938 ( .A(n6179), .B(n6178), .Z(n6181) );
  XNOR U6939 ( .A(n6176), .B(n6175), .Z(n6178) );
  XNOR U6940 ( .A(n6173), .B(n6172), .Z(n6175) );
  XNOR U6941 ( .A(n6170), .B(n6169), .Z(n6172) );
  XNOR U6942 ( .A(n6167), .B(n6166), .Z(n6169) );
  XNOR U6943 ( .A(n6164), .B(n6163), .Z(n6166) );
  XNOR U6944 ( .A(n6161), .B(n6160), .Z(n6163) );
  XNOR U6945 ( .A(n6158), .B(n6157), .Z(n6160) );
  XNOR U6946 ( .A(n6155), .B(n6154), .Z(n6157) );
  XNOR U6947 ( .A(n6152), .B(n6151), .Z(n6154) );
  XNOR U6948 ( .A(n6149), .B(n6148), .Z(n6151) );
  XNOR U6949 ( .A(n6146), .B(n6145), .Z(n6148) );
  XNOR U6950 ( .A(n6143), .B(n6142), .Z(n6145) );
  XNOR U6951 ( .A(n6140), .B(n6139), .Z(n6142) );
  XNOR U6952 ( .A(n6137), .B(n6136), .Z(n6139) );
  XNOR U6953 ( .A(n6134), .B(n6133), .Z(n6136) );
  XNOR U6954 ( .A(n6131), .B(n6130), .Z(n6133) );
  XNOR U6955 ( .A(n6128), .B(n6127), .Z(n6130) );
  XNOR U6956 ( .A(n6125), .B(n6124), .Z(n6127) );
  XNOR U6957 ( .A(n6122), .B(n6121), .Z(n6124) );
  XNOR U6958 ( .A(n6119), .B(n6118), .Z(n6121) );
  XNOR U6959 ( .A(n6116), .B(n6115), .Z(n6118) );
  XNOR U6960 ( .A(n6113), .B(n6112), .Z(n6115) );
  XNOR U6961 ( .A(n6110), .B(n6109), .Z(n6112) );
  XNOR U6962 ( .A(n6107), .B(n6106), .Z(n6109) );
  XNOR U6963 ( .A(n6104), .B(n6103), .Z(n6106) );
  XNOR U6964 ( .A(n6101), .B(n6100), .Z(n6103) );
  XNOR U6965 ( .A(n6098), .B(n6097), .Z(n6100) );
  XNOR U6966 ( .A(n6095), .B(n6094), .Z(n6097) );
  XNOR U6967 ( .A(n6092), .B(n6091), .Z(n6094) );
  XNOR U6968 ( .A(n6089), .B(n6088), .Z(n6091) );
  XNOR U6969 ( .A(n6086), .B(n6085), .Z(n6088) );
  XNOR U6970 ( .A(n6083), .B(n6082), .Z(n6085) );
  XNOR U6971 ( .A(n6080), .B(n6079), .Z(n6082) );
  XNOR U6972 ( .A(n6077), .B(n6076), .Z(n6079) );
  XNOR U6973 ( .A(n6074), .B(n6073), .Z(n6076) );
  XNOR U6974 ( .A(n6071), .B(n6070), .Z(n6073) );
  XNOR U6975 ( .A(n6068), .B(n6067), .Z(n6070) );
  XNOR U6976 ( .A(n6065), .B(n6064), .Z(n6067) );
  XNOR U6977 ( .A(n6062), .B(n6061), .Z(n6064) );
  XNOR U6978 ( .A(n6059), .B(n6058), .Z(n6061) );
  XNOR U6979 ( .A(n6056), .B(n6055), .Z(n6058) );
  XNOR U6980 ( .A(n6053), .B(n6052), .Z(n6055) );
  XNOR U6981 ( .A(n6050), .B(n6049), .Z(n6052) );
  XNOR U6982 ( .A(n6047), .B(n6046), .Z(n6049) );
  XNOR U6983 ( .A(n6044), .B(n6043), .Z(n6046) );
  XNOR U6984 ( .A(n6041), .B(n6040), .Z(n6043) );
  XNOR U6985 ( .A(n6038), .B(n6037), .Z(n6040) );
  XNOR U6986 ( .A(n6035), .B(n6034), .Z(n6037) );
  XNOR U6987 ( .A(n6032), .B(n6031), .Z(n6034) );
  XNOR U6988 ( .A(n6029), .B(n6028), .Z(n6031) );
  XNOR U6989 ( .A(n6026), .B(n6025), .Z(n6028) );
  XNOR U6990 ( .A(n6023), .B(n6022), .Z(n6025) );
  XNOR U6991 ( .A(n6020), .B(n6019), .Z(n6022) );
  XNOR U6992 ( .A(n6017), .B(n6016), .Z(n6019) );
  XNOR U6993 ( .A(n6014), .B(n6013), .Z(n6016) );
  XNOR U6994 ( .A(n6011), .B(n6010), .Z(n6013) );
  XNOR U6995 ( .A(n6008), .B(n6007), .Z(n6010) );
  XNOR U6996 ( .A(n6005), .B(n6004), .Z(n6007) );
  XNOR U6997 ( .A(n6002), .B(n6001), .Z(n6004) );
  XNOR U6998 ( .A(n5999), .B(n5998), .Z(n6001) );
  XNOR U6999 ( .A(n5996), .B(n5995), .Z(n5998) );
  XNOR U7000 ( .A(n5993), .B(n5992), .Z(n5995) );
  XNOR U7001 ( .A(n5990), .B(n5989), .Z(n5992) );
  XNOR U7002 ( .A(n5987), .B(n5986), .Z(n5989) );
  XNOR U7003 ( .A(n5984), .B(n5983), .Z(n5986) );
  XNOR U7004 ( .A(n5981), .B(n5980), .Z(n5983) );
  XNOR U7005 ( .A(n5978), .B(n5977), .Z(n5980) );
  XNOR U7006 ( .A(n5975), .B(n5974), .Z(n5977) );
  XNOR U7007 ( .A(n5972), .B(n5971), .Z(n5974) );
  XNOR U7008 ( .A(n5969), .B(n5968), .Z(n5971) );
  XNOR U7009 ( .A(n5966), .B(n5965), .Z(n5968) );
  XNOR U7010 ( .A(n5963), .B(n5962), .Z(n5965) );
  XNOR U7011 ( .A(n5960), .B(n5959), .Z(n5962) );
  XNOR U7012 ( .A(n5957), .B(n5956), .Z(n5959) );
  XNOR U7013 ( .A(n5954), .B(n5953), .Z(n5956) );
  XNOR U7014 ( .A(n5951), .B(n5950), .Z(n5953) );
  XNOR U7015 ( .A(n5948), .B(n5947), .Z(n5950) );
  XNOR U7016 ( .A(n5945), .B(n5944), .Z(n5947) );
  XNOR U7017 ( .A(n5942), .B(n5941), .Z(n5944) );
  XNOR U7018 ( .A(n5939), .B(n5938), .Z(n5941) );
  XNOR U7019 ( .A(n5936), .B(n5935), .Z(n5938) );
  XNOR U7020 ( .A(n5933), .B(n5932), .Z(n5935) );
  XNOR U7021 ( .A(n5930), .B(n5929), .Z(n5932) );
  XNOR U7022 ( .A(n5927), .B(n5926), .Z(n5929) );
  XNOR U7023 ( .A(n5924), .B(n5923), .Z(n5926) );
  XNOR U7024 ( .A(n5921), .B(n5920), .Z(n5923) );
  XNOR U7025 ( .A(n5918), .B(n5917), .Z(n5920) );
  XNOR U7026 ( .A(n5915), .B(n5914), .Z(n5917) );
  XNOR U7027 ( .A(n5912), .B(n5911), .Z(n5914) );
  XNOR U7028 ( .A(n5909), .B(n5908), .Z(n5911) );
  XNOR U7029 ( .A(n5906), .B(n5905), .Z(n5908) );
  XNOR U7030 ( .A(n5903), .B(n5902), .Z(n5905) );
  XNOR U7031 ( .A(n5900), .B(n5899), .Z(n5902) );
  XNOR U7032 ( .A(n5897), .B(n5896), .Z(n5899) );
  XNOR U7033 ( .A(n5894), .B(n5893), .Z(n5896) );
  XNOR U7034 ( .A(n5891), .B(n5890), .Z(n5893) );
  XNOR U7035 ( .A(n5888), .B(n5887), .Z(n5890) );
  XNOR U7036 ( .A(n5885), .B(n5884), .Z(n5887) );
  XNOR U7037 ( .A(n5882), .B(n5881), .Z(n5884) );
  XNOR U7038 ( .A(n5879), .B(n5878), .Z(n5881) );
  XNOR U7039 ( .A(n5876), .B(n5875), .Z(n5878) );
  XNOR U7040 ( .A(n5873), .B(n5872), .Z(n5875) );
  XNOR U7041 ( .A(n5870), .B(n5869), .Z(n5872) );
  XOR U7042 ( .A(n5867), .B(n5584), .Z(n5869) );
  XNOR U7043 ( .A(n5585), .B(n5582), .Z(n5584) );
  XNOR U7044 ( .A(n5583), .B(n5578), .Z(n5582) );
  XOR U7045 ( .A(n5579), .B(n5599), .Z(n5578) );
  XOR U7046 ( .A(n8477), .B(n5597), .Z(n5599) );
  XNOR U7047 ( .A(n5598), .B(n5865), .Z(n5597) );
  XNOR U7048 ( .A(n5866), .B(n5864), .Z(n5865) );
  XNOR U7049 ( .A(n5594), .B(n5861), .Z(n5864) );
  XNOR U7050 ( .A(n5593), .B(n5616), .Z(n5861) );
  XNOR U7051 ( .A(n5611), .B(n5860), .Z(n5616) );
  XNOR U7052 ( .A(n5610), .B(n5855), .Z(n5860) );
  XOR U7053 ( .A(n5612), .B(n5854), .Z(n5855) );
  XOR U7054 ( .A(n5615), .B(n5851), .Z(n5854) );
  XOR U7055 ( .A(n5621), .B(n5849), .Z(n5851) );
  XOR U7056 ( .A(n5850), .B(n5846), .Z(n5849) );
  XOR U7057 ( .A(n5841), .B(n5840), .Z(n5846) );
  XOR U7058 ( .A(n5637), .B(n5839), .Z(n5840) );
  AND U7059 ( .A(n8478), .B(n8479), .Z(n5839) );
  XOR U7060 ( .A(n5838), .B(n5631), .Z(n5637) );
  AND U7061 ( .A(n8480), .B(n8481), .Z(n5631) );
  XOR U7062 ( .A(n5835), .B(n5636), .Z(n5838) );
  AND U7063 ( .A(n8482), .B(n8483), .Z(n5636) );
  XOR U7064 ( .A(n5834), .B(n5634), .Z(n5835) );
  AND U7065 ( .A(n8484), .B(n8485), .Z(n5634) );
  XNOR U7066 ( .A(n5828), .B(n5633), .Z(n5834) );
  AND U7067 ( .A(n8486), .B(n8487), .Z(n5633) );
  XNOR U7068 ( .A(n5819), .B(n5829), .Z(n5828) );
  AND U7069 ( .A(n8488), .B(n8489), .Z(n5829) );
  XOR U7070 ( .A(n5817), .B(n5818), .Z(n5819) );
  AND U7071 ( .A(n8490), .B(n8491), .Z(n5818) );
  XOR U7072 ( .A(n5824), .B(n5816), .Z(n5817) );
  AND U7073 ( .A(n8492), .B(n8493), .Z(n5816) );
  XNOR U7074 ( .A(n5791), .B(n5823), .Z(n5824) );
  AND U7075 ( .A(n8494), .B(n8495), .Z(n5823) );
  XNOR U7076 ( .A(n5813), .B(n5792), .Z(n5791) );
  AND U7077 ( .A(n8496), .B(n8497), .Z(n5792) );
  XOR U7078 ( .A(n5812), .B(n5789), .Z(n5813) );
  AND U7079 ( .A(n8498), .B(n8499), .Z(n5789) );
  XOR U7080 ( .A(n5822), .B(n5788), .Z(n5812) );
  AND U7081 ( .A(n8500), .B(n8501), .Z(n5788) );
  XNOR U7082 ( .A(n5800), .B(n5787), .Z(n5822) );
  AND U7083 ( .A(n8502), .B(n8503), .Z(n5787) );
  XNOR U7084 ( .A(n5805), .B(n5801), .Z(n5800) );
  AND U7085 ( .A(n8504), .B(n8505), .Z(n5801) );
  XOR U7086 ( .A(n5804), .B(n5798), .Z(n5805) );
  AND U7087 ( .A(n8506), .B(n8507), .Z(n5798) );
  XOR U7088 ( .A(n5784), .B(n5797), .Z(n5804) );
  AND U7089 ( .A(n8508), .B(n8509), .Z(n5797) );
  XNOR U7090 ( .A(n5755), .B(n5783), .Z(n5784) );
  AND U7091 ( .A(n8510), .B(n8511), .Z(n5783) );
  XNOR U7092 ( .A(n5778), .B(n5756), .Z(n5755) );
  AND U7093 ( .A(n8512), .B(n8513), .Z(n5756) );
  XOR U7094 ( .A(n5777), .B(n5753), .Z(n5778) );
  AND U7095 ( .A(n8514), .B(n8515), .Z(n5753) );
  XOR U7096 ( .A(n5782), .B(n5752), .Z(n5777) );
  AND U7097 ( .A(n8516), .B(n8517), .Z(n5752) );
  XNOR U7098 ( .A(n5765), .B(n5751), .Z(n5782) );
  AND U7099 ( .A(n8518), .B(n8519), .Z(n5751) );
  XNOR U7100 ( .A(n5770), .B(n5766), .Z(n5765) );
  AND U7101 ( .A(n8520), .B(n8521), .Z(n5766) );
  XOR U7102 ( .A(n5769), .B(n5763), .Z(n5770) );
  AND U7103 ( .A(n8522), .B(n8523), .Z(n5763) );
  XOR U7104 ( .A(n5779), .B(n5762), .Z(n5769) );
  AND U7105 ( .A(n8524), .B(n8525), .Z(n5762) );
  XNOR U7106 ( .A(n5662), .B(n5761), .Z(n5779) );
  AND U7107 ( .A(n8526), .B(n8527), .Z(n5761) );
  XNOR U7108 ( .A(n5744), .B(n5663), .Z(n5662) );
  AND U7109 ( .A(n8528), .B(n8529), .Z(n5663) );
  XOR U7110 ( .A(n5743), .B(n5660), .Z(n5744) );
  AND U7111 ( .A(n8530), .B(n8531), .Z(n5660) );
  XOR U7112 ( .A(n5748), .B(n5659), .Z(n5743) );
  AND U7113 ( .A(n8532), .B(n8533), .Z(n5659) );
  XNOR U7114 ( .A(n5670), .B(n5658), .Z(n5748) );
  AND U7115 ( .A(n8534), .B(n8535), .Z(n5658) );
  XNOR U7116 ( .A(n5740), .B(n5671), .Z(n5670) );
  AND U7117 ( .A(n8536), .B(n8537), .Z(n5671) );
  XOR U7118 ( .A(n5739), .B(n5668), .Z(n5740) );
  AND U7119 ( .A(n8538), .B(n8539), .Z(n5668) );
  XOR U7120 ( .A(n5747), .B(n5667), .Z(n5739) );
  AND U7121 ( .A(n8540), .B(n8541), .Z(n5667) );
  XNOR U7122 ( .A(n5680), .B(n5666), .Z(n5747) );
  AND U7123 ( .A(n8542), .B(n8543), .Z(n5666) );
  XNOR U7124 ( .A(n5687), .B(n5681), .Z(n5680) );
  AND U7125 ( .A(n8544), .B(n8545), .Z(n5681) );
  XOR U7126 ( .A(n5686), .B(n5678), .Z(n5687) );
  AND U7127 ( .A(n8546), .B(n8547), .Z(n5678) );
  XOR U7128 ( .A(n5732), .B(n5677), .Z(n5686) );
  AND U7129 ( .A(n8548), .B(n8549), .Z(n5677) );
  XNOR U7130 ( .A(n5698), .B(n5676), .Z(n5732) );
  AND U7131 ( .A(n8550), .B(n8551), .Z(n5676) );
  XNOR U7132 ( .A(n5705), .B(n5699), .Z(n5698) );
  AND U7133 ( .A(n8552), .B(n8553), .Z(n5699) );
  XOR U7134 ( .A(n5704), .B(n5696), .Z(n5705) );
  AND U7135 ( .A(n8554), .B(n8555), .Z(n5696) );
  XOR U7136 ( .A(n5731), .B(n5695), .Z(n5704) );
  AND U7137 ( .A(n8556), .B(n8557), .Z(n5695) );
  XNOR U7138 ( .A(n5716), .B(n5694), .Z(n5731) );
  AND U7139 ( .A(n8558), .B(n8559), .Z(n5694) );
  XOR U7140 ( .A(n8560), .B(n5717), .Z(n5716) );
  AND U7141 ( .A(n8561), .B(n8562), .Z(n5717) );
  XOR U7142 ( .A(n8563), .B(n8564), .Z(n8560) );
  XOR U7143 ( .A(n8565), .B(n8566), .Z(n8564) );
  XOR U7144 ( .A(n5729), .B(n5730), .Z(n8566) );
  AND U7145 ( .A(n8567), .B(n8568), .Z(n5730) );
  AND U7146 ( .A(n8569), .B(n8570), .Z(n5729) );
  XNOR U7147 ( .A(n5727), .B(n5726), .Z(n8565) );
  IV U7148 ( .A(n8571), .Z(n5726) );
  AND U7149 ( .A(n8572), .B(n8573), .Z(n8571) );
  AND U7150 ( .A(n8574), .B(n8575), .Z(n5727) );
  XOR U7151 ( .A(n8576), .B(n8577), .Z(n8563) );
  XNOR U7152 ( .A(n5712), .B(n5721), .Z(n8577) );
  IV U7153 ( .A(n5713), .Z(n5721) );
  AND U7154 ( .A(n8578), .B(n8579), .Z(n5713) );
  AND U7155 ( .A(n8580), .B(n8581), .Z(n5712) );
  XOR U7156 ( .A(n5728), .B(n5714), .Z(n8576) );
  AND U7157 ( .A(n8582), .B(n8583), .Z(n5714) );
  XNOR U7158 ( .A(n8584), .B(n8585), .Z(n5728) );
  AND U7159 ( .A(n8586), .B(n8587), .Z(n8585) );
  NOR U7160 ( .A(n8588), .B(n8589), .Z(n8587) );
  NOR U7161 ( .A(n8590), .B(n8591), .Z(n8586) );
  AND U7162 ( .A(n8592), .B(n8593), .Z(n8591) );
  AND U7163 ( .A(n8594), .B(n8595), .Z(n8584) );
  NOR U7164 ( .A(n8596), .B(n8597), .Z(n8595) );
  AND U7165 ( .A(n8589), .B(n8598), .Z(n8597) );
  AND U7166 ( .A(n8590), .B(n8599), .Z(n8596) );
  NOR U7167 ( .A(n8600), .B(n8601), .Z(n8594) );
  XOR U7168 ( .A(n8602), .B(n8603), .Z(n8601) );
  AND U7169 ( .A(n8604), .B(n8605), .Z(n8603) );
  NOR U7170 ( .A(n8606), .B(n8607), .Z(n8605) );
  NOR U7171 ( .A(n8608), .B(n8609), .Z(n8604) );
  AND U7172 ( .A(n8610), .B(n8611), .Z(n8609) );
  AND U7173 ( .A(n8612), .B(n8613), .Z(n8602) );
  NOR U7174 ( .A(n8614), .B(n8615), .Z(n8613) );
  AND U7175 ( .A(n8607), .B(n8616), .Z(n8615) );
  AND U7176 ( .A(n8608), .B(n8617), .Z(n8614) );
  NOR U7177 ( .A(n8618), .B(n8619), .Z(n8612) );
  XOR U7178 ( .A(n8620), .B(n8621), .Z(n8619) );
  AND U7179 ( .A(n8622), .B(n8623), .Z(n8621) );
  NOR U7180 ( .A(n8624), .B(n8625), .Z(n8623) );
  NOR U7181 ( .A(n8626), .B(n8627), .Z(n8622) );
  AND U7182 ( .A(n8628), .B(n8629), .Z(n8627) );
  AND U7183 ( .A(n8630), .B(n8631), .Z(n8620) );
  NOR U7184 ( .A(n8632), .B(n8633), .Z(n8631) );
  AND U7185 ( .A(n8625), .B(n8634), .Z(n8633) );
  AND U7186 ( .A(n8626), .B(n8635), .Z(n8632) );
  NOR U7187 ( .A(n8636), .B(n8637), .Z(n8630) );
  XOR U7188 ( .A(n8638), .B(n8639), .Z(n8637) );
  AND U7189 ( .A(n8640), .B(n8641), .Z(n8639) );
  NOR U7190 ( .A(n8642), .B(n8643), .Z(n8641) );
  NOR U7191 ( .A(n8644), .B(n8645), .Z(n8640) );
  AND U7192 ( .A(n8646), .B(n8647), .Z(n8645) );
  AND U7193 ( .A(n8648), .B(n8649), .Z(n8638) );
  NOR U7194 ( .A(n8650), .B(n8651), .Z(n8649) );
  AND U7195 ( .A(n8643), .B(n8652), .Z(n8651) );
  AND U7196 ( .A(n8644), .B(n8653), .Z(n8650) );
  NOR U7197 ( .A(n8654), .B(n8655), .Z(n8648) );
  AND U7198 ( .A(n8656), .B(n8657), .Z(n8655) );
  AND U7199 ( .A(n8658), .B(n8659), .Z(n8657) );
  AND U7200 ( .A(n8660), .B(n8661), .Z(n8659) );
  AND U7201 ( .A(n8662), .B(n8663), .Z(n8661) );
  NOR U7202 ( .A(n8664), .B(n8665), .Z(n8662) );
  NOR U7203 ( .A(n8666), .B(n8667), .Z(n8660) );
  AND U7204 ( .A(n8668), .B(n8669), .Z(n8658) );
  NOR U7205 ( .A(n8670), .B(n8671), .Z(n8669) );
  NOR U7206 ( .A(n8672), .B(n8673), .Z(n8668) );
  AND U7207 ( .A(n8674), .B(n8675), .Z(n8656) );
  AND U7208 ( .A(n8676), .B(n8677), .Z(n8675) );
  NOR U7209 ( .A(n8678), .B(n8679), .Z(n8677) );
  NOR U7210 ( .A(n8680), .B(n8681), .Z(n8676) );
  AND U7211 ( .A(n8682), .B(n8683), .Z(n8674) );
  NOR U7212 ( .A(n8684), .B(n8685), .Z(n8683) );
  NOR U7213 ( .A(n8686), .B(n8687), .Z(n8682) );
  AND U7214 ( .A(n8642), .B(n8688), .Z(n8654) );
  AND U7215 ( .A(n8624), .B(n8689), .Z(n8636) );
  AND U7216 ( .A(n8606), .B(n8690), .Z(n8618) );
  AND U7217 ( .A(n8588), .B(n8691), .Z(n8600) );
  XOR U7218 ( .A(n8692), .B(n8693), .Z(n5841) );
  AND U7219 ( .A(n8692), .B(n8694), .Z(n8693) );
  IV U7220 ( .A(n5842), .Z(n5850) );
  XNOR U7221 ( .A(n8695), .B(n8696), .Z(n5842) );
  AND U7222 ( .A(n8695), .B(n8697), .Z(n8696) );
  XOR U7223 ( .A(n8698), .B(n8699), .Z(n5621) );
  AND U7224 ( .A(n8698), .B(n8700), .Z(n8699) );
  XOR U7225 ( .A(n8701), .B(n8702), .Z(n5615) );
  AND U7226 ( .A(n8701), .B(n8703), .Z(n8702) );
  XNOR U7227 ( .A(n8704), .B(n8705), .Z(n5612) );
  AND U7228 ( .A(n8704), .B(n8706), .Z(n8705) );
  XNOR U7229 ( .A(n8707), .B(n8708), .Z(n5610) );
  AND U7230 ( .A(n8709), .B(n8707), .Z(n8708) );
  XOR U7231 ( .A(n8710), .B(n8711), .Z(n5611) );
  NOR U7232 ( .A(n8712), .B(n8710), .Z(n8711) );
  XOR U7233 ( .A(n8713), .B(n8714), .Z(n5593) );
  NOR U7234 ( .A(n8715), .B(n8713), .Z(n8714) );
  XOR U7235 ( .A(n8716), .B(n8717), .Z(n5594) );
  NOR U7236 ( .A(n8718), .B(n8716), .Z(n8717) );
  XOR U7237 ( .A(n8719), .B(n8720), .Z(n5866) );
  NOR U7238 ( .A(n8721), .B(n8719), .Z(n8720) );
  XOR U7239 ( .A(n8722), .B(n8723), .Z(n5598) );
  NOR U7240 ( .A(n8724), .B(n8722), .Z(n8723) );
  IV U7241 ( .A(n5577), .Z(n8477) );
  XNOR U7242 ( .A(n8725), .B(n8726), .Z(n5577) );
  NOR U7243 ( .A(n8727), .B(n8725), .Z(n8726) );
  XOR U7244 ( .A(n8728), .B(n8729), .Z(n5579) );
  NOR U7245 ( .A(n8730), .B(n8728), .Z(n8729) );
  XOR U7246 ( .A(n8731), .B(n8732), .Z(n5583) );
  NOR U7247 ( .A(n8733), .B(n8731), .Z(n8732) );
  XNOR U7248 ( .A(n8734), .B(n8735), .Z(n5585) );
  NOR U7249 ( .A(n8736), .B(n8734), .Z(n8735) );
  XOR U7250 ( .A(n8737), .B(n8738), .Z(n5867) );
  NOR U7251 ( .A(n8739), .B(n8737), .Z(n8738) );
  XOR U7252 ( .A(n8740), .B(n8741), .Z(n5870) );
  NOR U7253 ( .A(n8742), .B(n8740), .Z(n8741) );
  XOR U7254 ( .A(n8743), .B(n8744), .Z(n5873) );
  NOR U7255 ( .A(n8745), .B(n8743), .Z(n8744) );
  XOR U7256 ( .A(n8746), .B(n8747), .Z(n5876) );
  NOR U7257 ( .A(n8748), .B(n8746), .Z(n8747) );
  XOR U7258 ( .A(n8749), .B(n8750), .Z(n5879) );
  NOR U7259 ( .A(n8751), .B(n8749), .Z(n8750) );
  XOR U7260 ( .A(n8752), .B(n8753), .Z(n5882) );
  NOR U7261 ( .A(n8754), .B(n8752), .Z(n8753) );
  XOR U7262 ( .A(n8755), .B(n8756), .Z(n5885) );
  NOR U7263 ( .A(n8757), .B(n8755), .Z(n8756) );
  XOR U7264 ( .A(n8758), .B(n8759), .Z(n5888) );
  NOR U7265 ( .A(n8760), .B(n8758), .Z(n8759) );
  XOR U7266 ( .A(n8761), .B(n8762), .Z(n5891) );
  NOR U7267 ( .A(n8763), .B(n8761), .Z(n8762) );
  XOR U7268 ( .A(n8764), .B(n8765), .Z(n5894) );
  NOR U7269 ( .A(n8766), .B(n8764), .Z(n8765) );
  XOR U7270 ( .A(n8767), .B(n8768), .Z(n5897) );
  NOR U7271 ( .A(n8769), .B(n8767), .Z(n8768) );
  XOR U7272 ( .A(n8770), .B(n8771), .Z(n5900) );
  NOR U7273 ( .A(n8772), .B(n8770), .Z(n8771) );
  XOR U7274 ( .A(n8773), .B(n8774), .Z(n5903) );
  NOR U7275 ( .A(n8775), .B(n8773), .Z(n8774) );
  XOR U7276 ( .A(n8776), .B(n8777), .Z(n5906) );
  NOR U7277 ( .A(n8778), .B(n8776), .Z(n8777) );
  XOR U7278 ( .A(n8779), .B(n8780), .Z(n5909) );
  NOR U7279 ( .A(n8781), .B(n8779), .Z(n8780) );
  XOR U7280 ( .A(n8782), .B(n8783), .Z(n5912) );
  NOR U7281 ( .A(n8784), .B(n8782), .Z(n8783) );
  XOR U7282 ( .A(n8785), .B(n8786), .Z(n5915) );
  NOR U7283 ( .A(n8787), .B(n8785), .Z(n8786) );
  XOR U7284 ( .A(n8788), .B(n8789), .Z(n5918) );
  NOR U7285 ( .A(n8790), .B(n8788), .Z(n8789) );
  XOR U7286 ( .A(n8791), .B(n8792), .Z(n5921) );
  NOR U7287 ( .A(n8793), .B(n8791), .Z(n8792) );
  XOR U7288 ( .A(n8794), .B(n8795), .Z(n5924) );
  NOR U7289 ( .A(n8796), .B(n8794), .Z(n8795) );
  XOR U7290 ( .A(n8797), .B(n8798), .Z(n5927) );
  NOR U7291 ( .A(n8799), .B(n8797), .Z(n8798) );
  XOR U7292 ( .A(n8800), .B(n8801), .Z(n5930) );
  NOR U7293 ( .A(n8802), .B(n8800), .Z(n8801) );
  XOR U7294 ( .A(n8803), .B(n8804), .Z(n5933) );
  NOR U7295 ( .A(n8805), .B(n8803), .Z(n8804) );
  XOR U7296 ( .A(n8806), .B(n8807), .Z(n5936) );
  NOR U7297 ( .A(n8808), .B(n8806), .Z(n8807) );
  XOR U7298 ( .A(n8809), .B(n8810), .Z(n5939) );
  NOR U7299 ( .A(n8811), .B(n8809), .Z(n8810) );
  XOR U7300 ( .A(n8812), .B(n8813), .Z(n5942) );
  NOR U7301 ( .A(n8814), .B(n8812), .Z(n8813) );
  XOR U7302 ( .A(n8815), .B(n8816), .Z(n5945) );
  NOR U7303 ( .A(n8817), .B(n8815), .Z(n8816) );
  XOR U7304 ( .A(n8818), .B(n8819), .Z(n5948) );
  NOR U7305 ( .A(n8820), .B(n8818), .Z(n8819) );
  XOR U7306 ( .A(n8821), .B(n8822), .Z(n5951) );
  NOR U7307 ( .A(n8823), .B(n8821), .Z(n8822) );
  XOR U7308 ( .A(n8824), .B(n8825), .Z(n5954) );
  NOR U7309 ( .A(n8826), .B(n8824), .Z(n8825) );
  XOR U7310 ( .A(n8827), .B(n8828), .Z(n5957) );
  NOR U7311 ( .A(n8829), .B(n8827), .Z(n8828) );
  XOR U7312 ( .A(n8830), .B(n8831), .Z(n5960) );
  NOR U7313 ( .A(n8832), .B(n8830), .Z(n8831) );
  XOR U7314 ( .A(n8833), .B(n8834), .Z(n5963) );
  NOR U7315 ( .A(n8835), .B(n8833), .Z(n8834) );
  XOR U7316 ( .A(n8836), .B(n8837), .Z(n5966) );
  NOR U7317 ( .A(n8838), .B(n8836), .Z(n8837) );
  XOR U7318 ( .A(n8839), .B(n8840), .Z(n5969) );
  NOR U7319 ( .A(n8841), .B(n8839), .Z(n8840) );
  XOR U7320 ( .A(n8842), .B(n8843), .Z(n5972) );
  NOR U7321 ( .A(n8844), .B(n8842), .Z(n8843) );
  XOR U7322 ( .A(n8845), .B(n8846), .Z(n5975) );
  NOR U7323 ( .A(n8847), .B(n8845), .Z(n8846) );
  XOR U7324 ( .A(n8848), .B(n8849), .Z(n5978) );
  NOR U7325 ( .A(n8850), .B(n8848), .Z(n8849) );
  XOR U7326 ( .A(n8851), .B(n8852), .Z(n5981) );
  NOR U7327 ( .A(n8853), .B(n8851), .Z(n8852) );
  XOR U7328 ( .A(n8854), .B(n8855), .Z(n5984) );
  NOR U7329 ( .A(n8856), .B(n8854), .Z(n8855) );
  XOR U7330 ( .A(n8857), .B(n8858), .Z(n5987) );
  NOR U7331 ( .A(n8859), .B(n8857), .Z(n8858) );
  XOR U7332 ( .A(n8860), .B(n8861), .Z(n5990) );
  NOR U7333 ( .A(n8862), .B(n8860), .Z(n8861) );
  XOR U7334 ( .A(n8863), .B(n8864), .Z(n5993) );
  NOR U7335 ( .A(n8865), .B(n8863), .Z(n8864) );
  XOR U7336 ( .A(n8866), .B(n8867), .Z(n5996) );
  NOR U7337 ( .A(n8868), .B(n8866), .Z(n8867) );
  XOR U7338 ( .A(n8869), .B(n8870), .Z(n5999) );
  NOR U7339 ( .A(n8871), .B(n8869), .Z(n8870) );
  XOR U7340 ( .A(n8872), .B(n8873), .Z(n6002) );
  NOR U7341 ( .A(n8874), .B(n8872), .Z(n8873) );
  XOR U7342 ( .A(n8875), .B(n8876), .Z(n6005) );
  NOR U7343 ( .A(n8877), .B(n8875), .Z(n8876) );
  XOR U7344 ( .A(n8878), .B(n8879), .Z(n6008) );
  NOR U7345 ( .A(n8880), .B(n8878), .Z(n8879) );
  XOR U7346 ( .A(n8881), .B(n8882), .Z(n6011) );
  NOR U7347 ( .A(n8883), .B(n8881), .Z(n8882) );
  XOR U7348 ( .A(n8884), .B(n8885), .Z(n6014) );
  NOR U7349 ( .A(n8886), .B(n8884), .Z(n8885) );
  XOR U7350 ( .A(n8887), .B(n8888), .Z(n6017) );
  NOR U7351 ( .A(n8889), .B(n8887), .Z(n8888) );
  XOR U7352 ( .A(n8890), .B(n8891), .Z(n6020) );
  NOR U7353 ( .A(n8892), .B(n8890), .Z(n8891) );
  XOR U7354 ( .A(n8893), .B(n8894), .Z(n6023) );
  NOR U7355 ( .A(n8895), .B(n8893), .Z(n8894) );
  XOR U7356 ( .A(n8896), .B(n8897), .Z(n6026) );
  NOR U7357 ( .A(n8898), .B(n8896), .Z(n8897) );
  XOR U7358 ( .A(n8899), .B(n8900), .Z(n6029) );
  NOR U7359 ( .A(n8901), .B(n8899), .Z(n8900) );
  XOR U7360 ( .A(n8902), .B(n8903), .Z(n6032) );
  NOR U7361 ( .A(n8904), .B(n8902), .Z(n8903) );
  XOR U7362 ( .A(n8905), .B(n8906), .Z(n6035) );
  NOR U7363 ( .A(n8907), .B(n8905), .Z(n8906) );
  XOR U7364 ( .A(n8908), .B(n8909), .Z(n6038) );
  NOR U7365 ( .A(n8910), .B(n8908), .Z(n8909) );
  XOR U7366 ( .A(n8911), .B(n8912), .Z(n6041) );
  NOR U7367 ( .A(n8913), .B(n8911), .Z(n8912) );
  XOR U7368 ( .A(n8914), .B(n8915), .Z(n6044) );
  NOR U7369 ( .A(n8916), .B(n8914), .Z(n8915) );
  XOR U7370 ( .A(n8917), .B(n8918), .Z(n6047) );
  NOR U7371 ( .A(n8919), .B(n8917), .Z(n8918) );
  XOR U7372 ( .A(n8920), .B(n8921), .Z(n6050) );
  NOR U7373 ( .A(n8922), .B(n8920), .Z(n8921) );
  XOR U7374 ( .A(n8923), .B(n8924), .Z(n6053) );
  NOR U7375 ( .A(n8925), .B(n8923), .Z(n8924) );
  XOR U7376 ( .A(n8926), .B(n8927), .Z(n6056) );
  NOR U7377 ( .A(n8928), .B(n8926), .Z(n8927) );
  XOR U7378 ( .A(n8929), .B(n8930), .Z(n6059) );
  NOR U7379 ( .A(n8931), .B(n8929), .Z(n8930) );
  XOR U7380 ( .A(n8932), .B(n8933), .Z(n6062) );
  NOR U7381 ( .A(n8934), .B(n8932), .Z(n8933) );
  XOR U7382 ( .A(n8935), .B(n8936), .Z(n6065) );
  NOR U7383 ( .A(n8937), .B(n8935), .Z(n8936) );
  XOR U7384 ( .A(n8938), .B(n8939), .Z(n6068) );
  NOR U7385 ( .A(n8940), .B(n8938), .Z(n8939) );
  XOR U7386 ( .A(n8941), .B(n8942), .Z(n6071) );
  NOR U7387 ( .A(n8943), .B(n8941), .Z(n8942) );
  XOR U7388 ( .A(n8944), .B(n8945), .Z(n6074) );
  NOR U7389 ( .A(n8946), .B(n8944), .Z(n8945) );
  XOR U7390 ( .A(n8947), .B(n8948), .Z(n6077) );
  NOR U7391 ( .A(n8949), .B(n8947), .Z(n8948) );
  XOR U7392 ( .A(n8950), .B(n8951), .Z(n6080) );
  NOR U7393 ( .A(n8952), .B(n8950), .Z(n8951) );
  XOR U7394 ( .A(n8953), .B(n8954), .Z(n6083) );
  NOR U7395 ( .A(n8955), .B(n8953), .Z(n8954) );
  XOR U7396 ( .A(n8956), .B(n8957), .Z(n6086) );
  NOR U7397 ( .A(n8958), .B(n8956), .Z(n8957) );
  XOR U7398 ( .A(n8959), .B(n8960), .Z(n6089) );
  NOR U7399 ( .A(n8961), .B(n8959), .Z(n8960) );
  XOR U7400 ( .A(n8962), .B(n8963), .Z(n6092) );
  NOR U7401 ( .A(n8964), .B(n8962), .Z(n8963) );
  XOR U7402 ( .A(n8965), .B(n8966), .Z(n6095) );
  NOR U7403 ( .A(n8967), .B(n8965), .Z(n8966) );
  XOR U7404 ( .A(n8968), .B(n8969), .Z(n6098) );
  NOR U7405 ( .A(n8970), .B(n8968), .Z(n8969) );
  XOR U7406 ( .A(n8971), .B(n8972), .Z(n6101) );
  NOR U7407 ( .A(n8973), .B(n8971), .Z(n8972) );
  XOR U7408 ( .A(n8974), .B(n8975), .Z(n6104) );
  NOR U7409 ( .A(n8976), .B(n8974), .Z(n8975) );
  XOR U7410 ( .A(n8977), .B(n8978), .Z(n6107) );
  NOR U7411 ( .A(n8979), .B(n8977), .Z(n8978) );
  XOR U7412 ( .A(n8980), .B(n8981), .Z(n6110) );
  NOR U7413 ( .A(n8982), .B(n8980), .Z(n8981) );
  XOR U7414 ( .A(n8983), .B(n8984), .Z(n6113) );
  NOR U7415 ( .A(n8985), .B(n8983), .Z(n8984) );
  XOR U7416 ( .A(n8986), .B(n8987), .Z(n6116) );
  NOR U7417 ( .A(n8988), .B(n8986), .Z(n8987) );
  XOR U7418 ( .A(n8989), .B(n8990), .Z(n6119) );
  NOR U7419 ( .A(n8991), .B(n8989), .Z(n8990) );
  XOR U7420 ( .A(n8992), .B(n8993), .Z(n6122) );
  NOR U7421 ( .A(n8994), .B(n8992), .Z(n8993) );
  XOR U7422 ( .A(n8995), .B(n8996), .Z(n6125) );
  NOR U7423 ( .A(n8997), .B(n8995), .Z(n8996) );
  XOR U7424 ( .A(n8998), .B(n8999), .Z(n6128) );
  NOR U7425 ( .A(n9000), .B(n8998), .Z(n8999) );
  XOR U7426 ( .A(n9001), .B(n9002), .Z(n6131) );
  NOR U7427 ( .A(n9003), .B(n9001), .Z(n9002) );
  XOR U7428 ( .A(n9004), .B(n9005), .Z(n6134) );
  NOR U7429 ( .A(n9006), .B(n9004), .Z(n9005) );
  XOR U7430 ( .A(n9007), .B(n9008), .Z(n6137) );
  NOR U7431 ( .A(n9009), .B(n9007), .Z(n9008) );
  XOR U7432 ( .A(n9010), .B(n9011), .Z(n6140) );
  NOR U7433 ( .A(n9012), .B(n9010), .Z(n9011) );
  XOR U7434 ( .A(n9013), .B(n9014), .Z(n6143) );
  NOR U7435 ( .A(n9015), .B(n9013), .Z(n9014) );
  XOR U7436 ( .A(n9016), .B(n9017), .Z(n6146) );
  NOR U7437 ( .A(n9018), .B(n9016), .Z(n9017) );
  XOR U7438 ( .A(n9019), .B(n9020), .Z(n6149) );
  NOR U7439 ( .A(n9021), .B(n9019), .Z(n9020) );
  XOR U7440 ( .A(n9022), .B(n9023), .Z(n6152) );
  NOR U7441 ( .A(n9024), .B(n9022), .Z(n9023) );
  XOR U7442 ( .A(n9025), .B(n9026), .Z(n6155) );
  NOR U7443 ( .A(n9027), .B(n9025), .Z(n9026) );
  XOR U7444 ( .A(n9028), .B(n9029), .Z(n6158) );
  NOR U7445 ( .A(n9030), .B(n9028), .Z(n9029) );
  XOR U7446 ( .A(n9031), .B(n9032), .Z(n6161) );
  NOR U7447 ( .A(n9033), .B(n9031), .Z(n9032) );
  XOR U7448 ( .A(n9034), .B(n9035), .Z(n6164) );
  NOR U7449 ( .A(n9036), .B(n9034), .Z(n9035) );
  XOR U7450 ( .A(n9037), .B(n9038), .Z(n6167) );
  NOR U7451 ( .A(n9039), .B(n9037), .Z(n9038) );
  XOR U7452 ( .A(n9040), .B(n9041), .Z(n6170) );
  NOR U7453 ( .A(n9042), .B(n9040), .Z(n9041) );
  XOR U7454 ( .A(n9043), .B(n9044), .Z(n6173) );
  NOR U7455 ( .A(n9045), .B(n9043), .Z(n9044) );
  XOR U7456 ( .A(n9046), .B(n9047), .Z(n6176) );
  NOR U7457 ( .A(n9048), .B(n9046), .Z(n9047) );
  XOR U7458 ( .A(n9049), .B(n9050), .Z(n6179) );
  NOR U7459 ( .A(n9051), .B(n9049), .Z(n9050) );
  XOR U7460 ( .A(n9052), .B(n9053), .Z(n6182) );
  NOR U7461 ( .A(n9054), .B(n9052), .Z(n9053) );
  XOR U7462 ( .A(n9055), .B(n9056), .Z(n6185) );
  NOR U7463 ( .A(n9057), .B(n9055), .Z(n9056) );
  XOR U7464 ( .A(n9058), .B(n9059), .Z(n6188) );
  NOR U7465 ( .A(n9060), .B(n9058), .Z(n9059) );
  XOR U7466 ( .A(n9061), .B(n9062), .Z(n6191) );
  NOR U7467 ( .A(n9063), .B(n9061), .Z(n9062) );
  XOR U7468 ( .A(n9064), .B(n9065), .Z(n6194) );
  NOR U7469 ( .A(n9066), .B(n9064), .Z(n9065) );
  XOR U7470 ( .A(n9067), .B(n9068), .Z(n6197) );
  NOR U7471 ( .A(n9069), .B(n9067), .Z(n9068) );
  XOR U7472 ( .A(n9070), .B(n9071), .Z(n6200) );
  NOR U7473 ( .A(n9072), .B(n9070), .Z(n9071) );
  XOR U7474 ( .A(n9073), .B(n9074), .Z(n6203) );
  NOR U7475 ( .A(n9075), .B(n9073), .Z(n9074) );
  XOR U7476 ( .A(n9076), .B(n9077), .Z(n6206) );
  NOR U7477 ( .A(n9078), .B(n9076), .Z(n9077) );
  XOR U7478 ( .A(n9079), .B(n9080), .Z(n6209) );
  NOR U7479 ( .A(n9081), .B(n9079), .Z(n9080) );
  XOR U7480 ( .A(n9082), .B(n9083), .Z(n6212) );
  NOR U7481 ( .A(n9084), .B(n9082), .Z(n9083) );
  XOR U7482 ( .A(n9085), .B(n9086), .Z(n6215) );
  NOR U7483 ( .A(n9087), .B(n9085), .Z(n9086) );
  XOR U7484 ( .A(n9088), .B(n9089), .Z(n6218) );
  NOR U7485 ( .A(n9090), .B(n9088), .Z(n9089) );
  XOR U7486 ( .A(n9091), .B(n9092), .Z(n6221) );
  NOR U7487 ( .A(n9093), .B(n9091), .Z(n9092) );
  XOR U7488 ( .A(n9094), .B(n9095), .Z(n6224) );
  NOR U7489 ( .A(n9096), .B(n9094), .Z(n9095) );
  XOR U7490 ( .A(n9097), .B(n9098), .Z(n6227) );
  NOR U7491 ( .A(n9099), .B(n9097), .Z(n9098) );
  XOR U7492 ( .A(n9100), .B(n9101), .Z(n6230) );
  NOR U7493 ( .A(n9102), .B(n9100), .Z(n9101) );
  XOR U7494 ( .A(n9103), .B(n9104), .Z(n6233) );
  NOR U7495 ( .A(n9105), .B(n9103), .Z(n9104) );
  XOR U7496 ( .A(n9106), .B(n9107), .Z(n6236) );
  NOR U7497 ( .A(n9108), .B(n9106), .Z(n9107) );
  XOR U7498 ( .A(n9109), .B(n9110), .Z(n6239) );
  NOR U7499 ( .A(n9111), .B(n9109), .Z(n9110) );
  XOR U7500 ( .A(n9112), .B(n9113), .Z(n6242) );
  NOR U7501 ( .A(n9114), .B(n9112), .Z(n9113) );
  XOR U7502 ( .A(n9115), .B(n9116), .Z(n6245) );
  NOR U7503 ( .A(n9117), .B(n9115), .Z(n9116) );
  XOR U7504 ( .A(n9118), .B(n9119), .Z(n6248) );
  NOR U7505 ( .A(n9120), .B(n9118), .Z(n9119) );
  XOR U7506 ( .A(n9121), .B(n9122), .Z(n6251) );
  NOR U7507 ( .A(n9123), .B(n9121), .Z(n9122) );
  XOR U7508 ( .A(n9124), .B(n9125), .Z(n6254) );
  NOR U7509 ( .A(n9126), .B(n9124), .Z(n9125) );
  XOR U7510 ( .A(n9127), .B(n9128), .Z(n6257) );
  NOR U7511 ( .A(n9129), .B(n9127), .Z(n9128) );
  XOR U7512 ( .A(n9130), .B(n9131), .Z(n6260) );
  NOR U7513 ( .A(n9132), .B(n9130), .Z(n9131) );
  XOR U7514 ( .A(n9133), .B(n9134), .Z(n6263) );
  NOR U7515 ( .A(n9135), .B(n9133), .Z(n9134) );
  XOR U7516 ( .A(n9136), .B(n9137), .Z(n6266) );
  NOR U7517 ( .A(n9138), .B(n9136), .Z(n9137) );
  XOR U7518 ( .A(n9139), .B(n9140), .Z(n6269) );
  NOR U7519 ( .A(n9141), .B(n9139), .Z(n9140) );
  XOR U7520 ( .A(n9142), .B(n9143), .Z(n6272) );
  NOR U7521 ( .A(n9144), .B(n9142), .Z(n9143) );
  XOR U7522 ( .A(n9145), .B(n9146), .Z(n6275) );
  NOR U7523 ( .A(n9147), .B(n9145), .Z(n9146) );
  XOR U7524 ( .A(n9148), .B(n9149), .Z(n6278) );
  NOR U7525 ( .A(n9150), .B(n9148), .Z(n9149) );
  XOR U7526 ( .A(n9151), .B(n9152), .Z(n6281) );
  NOR U7527 ( .A(n9153), .B(n9151), .Z(n9152) );
  XOR U7528 ( .A(n9154), .B(n9155), .Z(n6284) );
  NOR U7529 ( .A(n9156), .B(n9154), .Z(n9155) );
  XOR U7530 ( .A(n9157), .B(n9158), .Z(n6287) );
  NOR U7531 ( .A(n9159), .B(n9157), .Z(n9158) );
  XOR U7532 ( .A(n9160), .B(n9161), .Z(n6290) );
  NOR U7533 ( .A(n9162), .B(n9160), .Z(n9161) );
  XOR U7534 ( .A(n9163), .B(n9164), .Z(n6293) );
  NOR U7535 ( .A(n9165), .B(n9163), .Z(n9164) );
  XOR U7536 ( .A(n9166), .B(n9167), .Z(n6296) );
  NOR U7537 ( .A(n9168), .B(n9166), .Z(n9167) );
  XOR U7538 ( .A(n9169), .B(n9170), .Z(n6299) );
  NOR U7539 ( .A(n9171), .B(n9169), .Z(n9170) );
  XOR U7540 ( .A(n9172), .B(n9173), .Z(n6302) );
  NOR U7541 ( .A(n9174), .B(n9172), .Z(n9173) );
  XOR U7542 ( .A(n9175), .B(n9176), .Z(n6305) );
  NOR U7543 ( .A(n9177), .B(n9175), .Z(n9176) );
  XOR U7544 ( .A(n9178), .B(n9179), .Z(n6308) );
  NOR U7545 ( .A(n9180), .B(n9178), .Z(n9179) );
  XOR U7546 ( .A(n9181), .B(n9182), .Z(n6311) );
  NOR U7547 ( .A(n9183), .B(n9181), .Z(n9182) );
  XOR U7548 ( .A(n9184), .B(n9185), .Z(n6314) );
  NOR U7549 ( .A(n9186), .B(n9184), .Z(n9185) );
  XOR U7550 ( .A(n9187), .B(n9188), .Z(n6317) );
  NOR U7551 ( .A(n9189), .B(n9187), .Z(n9188) );
  XOR U7552 ( .A(n9190), .B(n9191), .Z(n6320) );
  NOR U7553 ( .A(n9192), .B(n9190), .Z(n9191) );
  XOR U7554 ( .A(n9193), .B(n9194), .Z(n6323) );
  NOR U7555 ( .A(n9195), .B(n9193), .Z(n9194) );
  XOR U7556 ( .A(n9196), .B(n9197), .Z(n6326) );
  NOR U7557 ( .A(n9198), .B(n9196), .Z(n9197) );
  XOR U7558 ( .A(n9199), .B(n9200), .Z(n6329) );
  NOR U7559 ( .A(n9201), .B(n9199), .Z(n9200) );
  XOR U7560 ( .A(n9202), .B(n9203), .Z(n6332) );
  NOR U7561 ( .A(n9204), .B(n9202), .Z(n9203) );
  XOR U7562 ( .A(n9205), .B(n9206), .Z(n6335) );
  NOR U7563 ( .A(n9207), .B(n9205), .Z(n9206) );
  XOR U7564 ( .A(n9208), .B(n9209), .Z(n6338) );
  NOR U7565 ( .A(n9210), .B(n9208), .Z(n9209) );
  XOR U7566 ( .A(n9211), .B(n9212), .Z(n6341) );
  NOR U7567 ( .A(n9213), .B(n9211), .Z(n9212) );
  XOR U7568 ( .A(n9214), .B(n9215), .Z(n6344) );
  NOR U7569 ( .A(n9216), .B(n9214), .Z(n9215) );
  XOR U7570 ( .A(n9217), .B(n9218), .Z(n6347) );
  NOR U7571 ( .A(n9219), .B(n9217), .Z(n9218) );
  XOR U7572 ( .A(n9220), .B(n9221), .Z(n6350) );
  NOR U7573 ( .A(n9222), .B(n9220), .Z(n9221) );
  XOR U7574 ( .A(n9223), .B(n9224), .Z(n6353) );
  NOR U7575 ( .A(n9225), .B(n9223), .Z(n9224) );
  XOR U7576 ( .A(n9226), .B(n9227), .Z(n6356) );
  NOR U7577 ( .A(n9228), .B(n9226), .Z(n9227) );
  XOR U7578 ( .A(n9229), .B(n9230), .Z(n6359) );
  NOR U7579 ( .A(n9231), .B(n9229), .Z(n9230) );
  XOR U7580 ( .A(n9232), .B(n9233), .Z(n6362) );
  NOR U7581 ( .A(n9234), .B(n9232), .Z(n9233) );
  XOR U7582 ( .A(n9235), .B(n9236), .Z(n6365) );
  NOR U7583 ( .A(n9237), .B(n9235), .Z(n9236) );
  XOR U7584 ( .A(n9238), .B(n9239), .Z(n6368) );
  NOR U7585 ( .A(n9240), .B(n9238), .Z(n9239) );
  XOR U7586 ( .A(n9241), .B(n9242), .Z(n6371) );
  NOR U7587 ( .A(n9243), .B(n9241), .Z(n9242) );
  XOR U7588 ( .A(n9244), .B(n9245), .Z(n6374) );
  NOR U7589 ( .A(n9246), .B(n9244), .Z(n9245) );
  XOR U7590 ( .A(n9247), .B(n9248), .Z(n6377) );
  NOR U7591 ( .A(n9249), .B(n9247), .Z(n9248) );
  XOR U7592 ( .A(n9250), .B(n9251), .Z(n6380) );
  NOR U7593 ( .A(n9252), .B(n9250), .Z(n9251) );
  XOR U7594 ( .A(n9253), .B(n9254), .Z(n6383) );
  NOR U7595 ( .A(n9255), .B(n9253), .Z(n9254) );
  XOR U7596 ( .A(n9256), .B(n9257), .Z(n6386) );
  NOR U7597 ( .A(n9258), .B(n9256), .Z(n9257) );
  XOR U7598 ( .A(n9259), .B(n9260), .Z(n6389) );
  NOR U7599 ( .A(n9261), .B(n9259), .Z(n9260) );
  XOR U7600 ( .A(n9262), .B(n9263), .Z(n6392) );
  NOR U7601 ( .A(n9264), .B(n9262), .Z(n9263) );
  XOR U7602 ( .A(n9265), .B(n9266), .Z(n6395) );
  NOR U7603 ( .A(n9267), .B(n9265), .Z(n9266) );
  XOR U7604 ( .A(n9268), .B(n9269), .Z(n6398) );
  NOR U7605 ( .A(n9270), .B(n9268), .Z(n9269) );
  XOR U7606 ( .A(n9271), .B(n9272), .Z(n6401) );
  NOR U7607 ( .A(n9273), .B(n9271), .Z(n9272) );
  XOR U7608 ( .A(n9274), .B(n9275), .Z(n6404) );
  NOR U7609 ( .A(n9276), .B(n9274), .Z(n9275) );
  XOR U7610 ( .A(n9277), .B(n9278), .Z(n6407) );
  NOR U7611 ( .A(n9279), .B(n9277), .Z(n9278) );
  XOR U7612 ( .A(n9280), .B(n9281), .Z(n6410) );
  NOR U7613 ( .A(n9282), .B(n9280), .Z(n9281) );
  XOR U7614 ( .A(n9283), .B(n9284), .Z(n6413) );
  NOR U7615 ( .A(n9285), .B(n9283), .Z(n9284) );
  XOR U7616 ( .A(n9286), .B(n9287), .Z(n6416) );
  NOR U7617 ( .A(n9288), .B(n9286), .Z(n9287) );
  XOR U7618 ( .A(n9289), .B(n9290), .Z(n6419) );
  NOR U7619 ( .A(n9291), .B(n9289), .Z(n9290) );
  XOR U7620 ( .A(n9292), .B(n9293), .Z(n6422) );
  NOR U7621 ( .A(n9294), .B(n9292), .Z(n9293) );
  XOR U7622 ( .A(n9295), .B(n9296), .Z(n6425) );
  NOR U7623 ( .A(n9297), .B(n9295), .Z(n9296) );
  XOR U7624 ( .A(n9298), .B(n9299), .Z(n6428) );
  NOR U7625 ( .A(n9300), .B(n9298), .Z(n9299) );
  XOR U7626 ( .A(n9301), .B(n9302), .Z(n6431) );
  NOR U7627 ( .A(n9303), .B(n9301), .Z(n9302) );
  XOR U7628 ( .A(n9304), .B(n9305), .Z(n6434) );
  NOR U7629 ( .A(n9306), .B(n9304), .Z(n9305) );
  XOR U7630 ( .A(n9307), .B(n9308), .Z(n6437) );
  NOR U7631 ( .A(n9309), .B(n9307), .Z(n9308) );
  XOR U7632 ( .A(n9310), .B(n9311), .Z(n6440) );
  NOR U7633 ( .A(n9312), .B(n9310), .Z(n9311) );
  XOR U7634 ( .A(n9313), .B(n9314), .Z(n6443) );
  NOR U7635 ( .A(n9315), .B(n9313), .Z(n9314) );
  XOR U7636 ( .A(n9316), .B(n9317), .Z(n6446) );
  NOR U7637 ( .A(n9318), .B(n9316), .Z(n9317) );
  XOR U7638 ( .A(n9319), .B(n9320), .Z(n6449) );
  NOR U7639 ( .A(n9321), .B(n9319), .Z(n9320) );
  XOR U7640 ( .A(n9322), .B(n9323), .Z(n6452) );
  NOR U7641 ( .A(n9324), .B(n9322), .Z(n9323) );
  XOR U7642 ( .A(n9325), .B(n9326), .Z(n6455) );
  NOR U7643 ( .A(n9327), .B(n9325), .Z(n9326) );
  XOR U7644 ( .A(n9328), .B(n9329), .Z(n6458) );
  NOR U7645 ( .A(n9330), .B(n9328), .Z(n9329) );
  XOR U7646 ( .A(n9331), .B(n9332), .Z(n6461) );
  NOR U7647 ( .A(n9333), .B(n9331), .Z(n9332) );
  XOR U7648 ( .A(n9334), .B(n9335), .Z(n6464) );
  NOR U7649 ( .A(n9336), .B(n9334), .Z(n9335) );
  XOR U7650 ( .A(n9337), .B(n9338), .Z(n6467) );
  NOR U7651 ( .A(n9339), .B(n9337), .Z(n9338) );
  XOR U7652 ( .A(n9340), .B(n9341), .Z(n6470) );
  NOR U7653 ( .A(n9342), .B(n9340), .Z(n9341) );
  XOR U7654 ( .A(n9343), .B(n9344), .Z(n6473) );
  NOR U7655 ( .A(n9345), .B(n9343), .Z(n9344) );
  XOR U7656 ( .A(n9346), .B(n9347), .Z(n6476) );
  NOR U7657 ( .A(n9348), .B(n9346), .Z(n9347) );
  XOR U7658 ( .A(n9349), .B(n9350), .Z(n6479) );
  NOR U7659 ( .A(n9351), .B(n9349), .Z(n9350) );
  XOR U7660 ( .A(n9352), .B(n9353), .Z(n6482) );
  NOR U7661 ( .A(n9354), .B(n9352), .Z(n9353) );
  XOR U7662 ( .A(n9355), .B(n9356), .Z(n6485) );
  NOR U7663 ( .A(n9357), .B(n9355), .Z(n9356) );
  XOR U7664 ( .A(n9358), .B(n9359), .Z(n6488) );
  NOR U7665 ( .A(n9360), .B(n9358), .Z(n9359) );
  XOR U7666 ( .A(n9361), .B(n9362), .Z(n6491) );
  NOR U7667 ( .A(n9363), .B(n9361), .Z(n9362) );
  XOR U7668 ( .A(n9364), .B(n9365), .Z(n6494) );
  NOR U7669 ( .A(n9366), .B(n9364), .Z(n9365) );
  XOR U7670 ( .A(n9367), .B(n9368), .Z(n6497) );
  NOR U7671 ( .A(n9369), .B(n9367), .Z(n9368) );
  XOR U7672 ( .A(n9370), .B(n9371), .Z(n6500) );
  NOR U7673 ( .A(n9372), .B(n9370), .Z(n9371) );
  XOR U7674 ( .A(n9373), .B(n9374), .Z(n6503) );
  NOR U7675 ( .A(n9375), .B(n9373), .Z(n9374) );
  XOR U7676 ( .A(n9376), .B(n9377), .Z(n6506) );
  NOR U7677 ( .A(n9378), .B(n9376), .Z(n9377) );
  XOR U7678 ( .A(n9379), .B(n9380), .Z(n6509) );
  NOR U7679 ( .A(n9381), .B(n9379), .Z(n9380) );
  XOR U7680 ( .A(n9382), .B(n9383), .Z(n6512) );
  NOR U7681 ( .A(n9384), .B(n9382), .Z(n9383) );
  XOR U7682 ( .A(n9385), .B(n9386), .Z(n6515) );
  NOR U7683 ( .A(n9387), .B(n9385), .Z(n9386) );
  XOR U7684 ( .A(n9388), .B(n9389), .Z(n6518) );
  NOR U7685 ( .A(n9390), .B(n9388), .Z(n9389) );
  XOR U7686 ( .A(n9391), .B(n9392), .Z(n6521) );
  NOR U7687 ( .A(n9393), .B(n9391), .Z(n9392) );
  XOR U7688 ( .A(n9394), .B(n9395), .Z(n6524) );
  NOR U7689 ( .A(n9396), .B(n9394), .Z(n9395) );
  XOR U7690 ( .A(n9397), .B(n9398), .Z(n6527) );
  NOR U7691 ( .A(n9399), .B(n9397), .Z(n9398) );
  XOR U7692 ( .A(n9400), .B(n9401), .Z(n6530) );
  NOR U7693 ( .A(n9402), .B(n9400), .Z(n9401) );
  XOR U7694 ( .A(n9403), .B(n9404), .Z(n6533) );
  NOR U7695 ( .A(n9405), .B(n9403), .Z(n9404) );
  XOR U7696 ( .A(n9406), .B(n9407), .Z(n6536) );
  NOR U7697 ( .A(n9408), .B(n9406), .Z(n9407) );
  XOR U7698 ( .A(n9409), .B(n9410), .Z(n6539) );
  NOR U7699 ( .A(n9411), .B(n9409), .Z(n9410) );
  XOR U7700 ( .A(n9412), .B(n9413), .Z(n6542) );
  NOR U7701 ( .A(n9414), .B(n9412), .Z(n9413) );
  XOR U7702 ( .A(n9415), .B(n9416), .Z(n6545) );
  NOR U7703 ( .A(n9417), .B(n9415), .Z(n9416) );
  XOR U7704 ( .A(n9418), .B(n9419), .Z(n6548) );
  NOR U7705 ( .A(n9420), .B(n9418), .Z(n9419) );
  XOR U7706 ( .A(n9421), .B(n9422), .Z(n6551) );
  NOR U7707 ( .A(n9423), .B(n9421), .Z(n9422) );
  XOR U7708 ( .A(n9424), .B(n9425), .Z(n6554) );
  NOR U7709 ( .A(n9426), .B(n9424), .Z(n9425) );
  XOR U7710 ( .A(n9427), .B(n9428), .Z(n6557) );
  NOR U7711 ( .A(n9429), .B(n9427), .Z(n9428) );
  XOR U7712 ( .A(n9430), .B(n9431), .Z(n6560) );
  NOR U7713 ( .A(n9432), .B(n9430), .Z(n9431) );
  XOR U7714 ( .A(n9433), .B(n9434), .Z(n6563) );
  NOR U7715 ( .A(n9435), .B(n9433), .Z(n9434) );
  XOR U7716 ( .A(n9436), .B(n9437), .Z(n6566) );
  NOR U7717 ( .A(n9438), .B(n9436), .Z(n9437) );
  XOR U7718 ( .A(n9439), .B(n9440), .Z(n6569) );
  NOR U7719 ( .A(n9441), .B(n9439), .Z(n9440) );
  XOR U7720 ( .A(n9442), .B(n9443), .Z(n6572) );
  NOR U7721 ( .A(n9444), .B(n9442), .Z(n9443) );
  XOR U7722 ( .A(n9445), .B(n9446), .Z(n6575) );
  NOR U7723 ( .A(n9447), .B(n9445), .Z(n9446) );
  XOR U7724 ( .A(n9448), .B(n9449), .Z(n6578) );
  NOR U7725 ( .A(n9450), .B(n9448), .Z(n9449) );
  XOR U7726 ( .A(n9451), .B(n9452), .Z(n6581) );
  NOR U7727 ( .A(n9453), .B(n9451), .Z(n9452) );
  XOR U7728 ( .A(n9454), .B(n9455), .Z(n6584) );
  NOR U7729 ( .A(n9456), .B(n9454), .Z(n9455) );
  XOR U7730 ( .A(n9457), .B(n9458), .Z(n6587) );
  NOR U7731 ( .A(n9459), .B(n9457), .Z(n9458) );
  XOR U7732 ( .A(n9460), .B(n9461), .Z(n6590) );
  NOR U7733 ( .A(n9462), .B(n9460), .Z(n9461) );
  XOR U7734 ( .A(n9463), .B(n9464), .Z(n6593) );
  NOR U7735 ( .A(n9465), .B(n9463), .Z(n9464) );
  XOR U7736 ( .A(n9466), .B(n9467), .Z(n6596) );
  NOR U7737 ( .A(n9468), .B(n9466), .Z(n9467) );
  XOR U7738 ( .A(n9469), .B(n9470), .Z(n6599) );
  NOR U7739 ( .A(n9471), .B(n9469), .Z(n9470) );
  XOR U7740 ( .A(n9472), .B(n9473), .Z(n6602) );
  NOR U7741 ( .A(n9474), .B(n9472), .Z(n9473) );
  XOR U7742 ( .A(n9475), .B(n9476), .Z(n6605) );
  NOR U7743 ( .A(n9477), .B(n9475), .Z(n9476) );
  XOR U7744 ( .A(n9478), .B(n9479), .Z(n6608) );
  NOR U7745 ( .A(n9480), .B(n9478), .Z(n9479) );
  XOR U7746 ( .A(n9481), .B(n9482), .Z(n6611) );
  NOR U7747 ( .A(n9483), .B(n9481), .Z(n9482) );
  XOR U7748 ( .A(n9484), .B(n9485), .Z(n6614) );
  NOR U7749 ( .A(n9486), .B(n9484), .Z(n9485) );
  XOR U7750 ( .A(n9487), .B(n9488), .Z(n6617) );
  NOR U7751 ( .A(n9489), .B(n9487), .Z(n9488) );
  XOR U7752 ( .A(n9490), .B(n9491), .Z(n6620) );
  NOR U7753 ( .A(n9492), .B(n9490), .Z(n9491) );
  XOR U7754 ( .A(n9493), .B(n9494), .Z(n6623) );
  NOR U7755 ( .A(n9495), .B(n9493), .Z(n9494) );
  XOR U7756 ( .A(n9496), .B(n9497), .Z(n6626) );
  NOR U7757 ( .A(n9498), .B(n9496), .Z(n9497) );
  XOR U7758 ( .A(n9499), .B(n9500), .Z(n6629) );
  NOR U7759 ( .A(n9501), .B(n9499), .Z(n9500) );
  XOR U7760 ( .A(n9502), .B(n9503), .Z(n6632) );
  NOR U7761 ( .A(n9504), .B(n9502), .Z(n9503) );
  XOR U7762 ( .A(n9505), .B(n9506), .Z(n6635) );
  NOR U7763 ( .A(n9507), .B(n9505), .Z(n9506) );
  XOR U7764 ( .A(n9508), .B(n9509), .Z(n6638) );
  NOR U7765 ( .A(n9510), .B(n9508), .Z(n9509) );
  XOR U7766 ( .A(n9511), .B(n9512), .Z(n6641) );
  NOR U7767 ( .A(n9513), .B(n9511), .Z(n9512) );
  XOR U7768 ( .A(n9514), .B(n9515), .Z(n6644) );
  NOR U7769 ( .A(n9516), .B(n9514), .Z(n9515) );
  XOR U7770 ( .A(n9517), .B(n9518), .Z(n6647) );
  NOR U7771 ( .A(n9519), .B(n9517), .Z(n9518) );
  XOR U7772 ( .A(n9520), .B(n9521), .Z(n6650) );
  NOR U7773 ( .A(n9522), .B(n9520), .Z(n9521) );
  XOR U7774 ( .A(n9523), .B(n9524), .Z(n6653) );
  NOR U7775 ( .A(n9525), .B(n9523), .Z(n9524) );
  XOR U7776 ( .A(n9526), .B(n9527), .Z(n6656) );
  NOR U7777 ( .A(n9528), .B(n9526), .Z(n9527) );
  XOR U7778 ( .A(n9529), .B(n9530), .Z(n6659) );
  NOR U7779 ( .A(n9531), .B(n9529), .Z(n9530) );
  XOR U7780 ( .A(n9532), .B(n9533), .Z(n6662) );
  NOR U7781 ( .A(n9534), .B(n9532), .Z(n9533) );
  XOR U7782 ( .A(n9535), .B(n9536), .Z(n6665) );
  NOR U7783 ( .A(n9537), .B(n9535), .Z(n9536) );
  XOR U7784 ( .A(n9538), .B(n9539), .Z(n6668) );
  NOR U7785 ( .A(n9540), .B(n9538), .Z(n9539) );
  XOR U7786 ( .A(n9541), .B(n9542), .Z(n6671) );
  NOR U7787 ( .A(n9543), .B(n9541), .Z(n9542) );
  XOR U7788 ( .A(n9544), .B(n9545), .Z(n6674) );
  NOR U7789 ( .A(n9546), .B(n9544), .Z(n9545) );
  XOR U7790 ( .A(n9547), .B(n9548), .Z(n6677) );
  NOR U7791 ( .A(n9549), .B(n9547), .Z(n9548) );
  XOR U7792 ( .A(n9550), .B(n9551), .Z(n6680) );
  NOR U7793 ( .A(n9552), .B(n9550), .Z(n9551) );
  XOR U7794 ( .A(n9553), .B(n9554), .Z(n6683) );
  NOR U7795 ( .A(n9555), .B(n9553), .Z(n9554) );
  XOR U7796 ( .A(n9556), .B(n9557), .Z(n6686) );
  NOR U7797 ( .A(n9558), .B(n9556), .Z(n9557) );
  XOR U7798 ( .A(n9559), .B(n9560), .Z(n6689) );
  NOR U7799 ( .A(n9561), .B(n9559), .Z(n9560) );
  XOR U7800 ( .A(n9562), .B(n9563), .Z(n6692) );
  NOR U7801 ( .A(n9564), .B(n9562), .Z(n9563) );
  XOR U7802 ( .A(n9565), .B(n9566), .Z(n6695) );
  NOR U7803 ( .A(n9567), .B(n9565), .Z(n9566) );
  XOR U7804 ( .A(n9568), .B(n9569), .Z(n6698) );
  NOR U7805 ( .A(n9570), .B(n9568), .Z(n9569) );
  XOR U7806 ( .A(n9571), .B(n9572), .Z(n6701) );
  NOR U7807 ( .A(n9573), .B(n9571), .Z(n9572) );
  XOR U7808 ( .A(n9574), .B(n9575), .Z(n6704) );
  NOR U7809 ( .A(n9576), .B(n9574), .Z(n9575) );
  XOR U7810 ( .A(n9577), .B(n9578), .Z(n6707) );
  NOR U7811 ( .A(n9579), .B(n9577), .Z(n9578) );
  XOR U7812 ( .A(n9580), .B(n9581), .Z(n6710) );
  NOR U7813 ( .A(n9582), .B(n9580), .Z(n9581) );
  XOR U7814 ( .A(n9583), .B(n9584), .Z(n6713) );
  NOR U7815 ( .A(n9585), .B(n9583), .Z(n9584) );
  XOR U7816 ( .A(n9586), .B(n9587), .Z(n6716) );
  NOR U7817 ( .A(n9588), .B(n9586), .Z(n9587) );
  XOR U7818 ( .A(n9589), .B(n9590), .Z(n6719) );
  NOR U7819 ( .A(n9591), .B(n9589), .Z(n9590) );
  XOR U7820 ( .A(n9592), .B(n9593), .Z(n6722) );
  NOR U7821 ( .A(n9594), .B(n9592), .Z(n9593) );
  XOR U7822 ( .A(n9595), .B(n9596), .Z(n6725) );
  NOR U7823 ( .A(n9597), .B(n9595), .Z(n9596) );
  XOR U7824 ( .A(n9598), .B(n9599), .Z(n6728) );
  NOR U7825 ( .A(n9600), .B(n9598), .Z(n9599) );
  XOR U7826 ( .A(n9601), .B(n9602), .Z(n6731) );
  NOR U7827 ( .A(n9603), .B(n9601), .Z(n9602) );
  XOR U7828 ( .A(n9604), .B(n9605), .Z(n6734) );
  NOR U7829 ( .A(n9606), .B(n9604), .Z(n9605) );
  XOR U7830 ( .A(n9607), .B(n9608), .Z(n6737) );
  NOR U7831 ( .A(n9609), .B(n9607), .Z(n9608) );
  XOR U7832 ( .A(n9610), .B(n9611), .Z(n6740) );
  NOR U7833 ( .A(n9612), .B(n9610), .Z(n9611) );
  XOR U7834 ( .A(n9613), .B(n9614), .Z(n6743) );
  NOR U7835 ( .A(n9615), .B(n9613), .Z(n9614) );
  XOR U7836 ( .A(n9616), .B(n9617), .Z(n6746) );
  NOR U7837 ( .A(n9618), .B(n9616), .Z(n9617) );
  XOR U7838 ( .A(n9619), .B(n9620), .Z(n6749) );
  NOR U7839 ( .A(n9621), .B(n9619), .Z(n9620) );
  XOR U7840 ( .A(n9622), .B(n9623), .Z(n6752) );
  NOR U7841 ( .A(n9624), .B(n9622), .Z(n9623) );
  XOR U7842 ( .A(n9625), .B(n9626), .Z(n6755) );
  NOR U7843 ( .A(n9627), .B(n9625), .Z(n9626) );
  XOR U7844 ( .A(n9628), .B(n9629), .Z(n6758) );
  NOR U7845 ( .A(n9630), .B(n9628), .Z(n9629) );
  XOR U7846 ( .A(n9631), .B(n9632), .Z(n6761) );
  NOR U7847 ( .A(n9633), .B(n9631), .Z(n9632) );
  XOR U7848 ( .A(n9634), .B(n9635), .Z(n6764) );
  NOR U7849 ( .A(n9636), .B(n9634), .Z(n9635) );
  XOR U7850 ( .A(n9637), .B(n9638), .Z(n6767) );
  NOR U7851 ( .A(n9639), .B(n9637), .Z(n9638) );
  XOR U7852 ( .A(n9640), .B(n9641), .Z(n6770) );
  NOR U7853 ( .A(n9642), .B(n9640), .Z(n9641) );
  XOR U7854 ( .A(n9643), .B(n9644), .Z(n6773) );
  NOR U7855 ( .A(n9645), .B(n9643), .Z(n9644) );
  XOR U7856 ( .A(n9646), .B(n9647), .Z(n6776) );
  NOR U7857 ( .A(n9648), .B(n9646), .Z(n9647) );
  XOR U7858 ( .A(n9649), .B(n9650), .Z(n6779) );
  NOR U7859 ( .A(n9651), .B(n9649), .Z(n9650) );
  XOR U7860 ( .A(n9652), .B(n9653), .Z(n6782) );
  NOR U7861 ( .A(n9654), .B(n9652), .Z(n9653) );
  XOR U7862 ( .A(n9655), .B(n9656), .Z(n6785) );
  NOR U7863 ( .A(n9657), .B(n9655), .Z(n9656) );
  XOR U7864 ( .A(n9658), .B(n9659), .Z(n6788) );
  NOR U7865 ( .A(n9660), .B(n9658), .Z(n9659) );
  XOR U7866 ( .A(n9661), .B(n9662), .Z(n6791) );
  NOR U7867 ( .A(n9663), .B(n9661), .Z(n9662) );
  XOR U7868 ( .A(n9664), .B(n9665), .Z(n6794) );
  NOR U7869 ( .A(n9666), .B(n9664), .Z(n9665) );
  XOR U7870 ( .A(n9667), .B(n9668), .Z(n6797) );
  NOR U7871 ( .A(n9669), .B(n9667), .Z(n9668) );
  XOR U7872 ( .A(n9670), .B(n9671), .Z(n6800) );
  NOR U7873 ( .A(n9672), .B(n9670), .Z(n9671) );
  XOR U7874 ( .A(n9673), .B(n9674), .Z(n6803) );
  NOR U7875 ( .A(n9675), .B(n9673), .Z(n9674) );
  XOR U7876 ( .A(n9676), .B(n9677), .Z(n6806) );
  NOR U7877 ( .A(n9678), .B(n9676), .Z(n9677) );
  XOR U7878 ( .A(n9679), .B(n9680), .Z(n6809) );
  NOR U7879 ( .A(n9681), .B(n9679), .Z(n9680) );
  XOR U7880 ( .A(n9682), .B(n9683), .Z(n6812) );
  NOR U7881 ( .A(n9684), .B(n9682), .Z(n9683) );
  XOR U7882 ( .A(n9685), .B(n9686), .Z(n6815) );
  NOR U7883 ( .A(n9687), .B(n9685), .Z(n9686) );
  XOR U7884 ( .A(n9688), .B(n9689), .Z(n6818) );
  NOR U7885 ( .A(n9690), .B(n9688), .Z(n9689) );
  XOR U7886 ( .A(n9691), .B(n9692), .Z(n6821) );
  NOR U7887 ( .A(n9693), .B(n9691), .Z(n9692) );
  XOR U7888 ( .A(n9694), .B(n9695), .Z(n6824) );
  NOR U7889 ( .A(n9696), .B(n9694), .Z(n9695) );
  XOR U7890 ( .A(n9697), .B(n9698), .Z(n6827) );
  NOR U7891 ( .A(n9699), .B(n9697), .Z(n9698) );
  XOR U7892 ( .A(n9700), .B(n9701), .Z(n6830) );
  NOR U7893 ( .A(n9702), .B(n9700), .Z(n9701) );
  XOR U7894 ( .A(n9703), .B(n9704), .Z(n6833) );
  NOR U7895 ( .A(n9705), .B(n9703), .Z(n9704) );
  XOR U7896 ( .A(n9706), .B(n9707), .Z(n6836) );
  NOR U7897 ( .A(n9708), .B(n9706), .Z(n9707) );
  XOR U7898 ( .A(n9709), .B(n9710), .Z(n6839) );
  NOR U7899 ( .A(n9711), .B(n9709), .Z(n9710) );
  XOR U7900 ( .A(n9712), .B(n9713), .Z(n6842) );
  NOR U7901 ( .A(n9714), .B(n9712), .Z(n9713) );
  XOR U7902 ( .A(n9715), .B(n9716), .Z(n6845) );
  NOR U7903 ( .A(n9717), .B(n9715), .Z(n9716) );
  XOR U7904 ( .A(n9718), .B(n9719), .Z(n6848) );
  NOR U7905 ( .A(n9720), .B(n9718), .Z(n9719) );
  XOR U7906 ( .A(n9721), .B(n9722), .Z(n6851) );
  NOR U7907 ( .A(n9723), .B(n9721), .Z(n9722) );
  XOR U7908 ( .A(n9724), .B(n9725), .Z(n6854) );
  NOR U7909 ( .A(n9726), .B(n9724), .Z(n9725) );
  XOR U7910 ( .A(n9727), .B(n9728), .Z(n6857) );
  NOR U7911 ( .A(n9729), .B(n9727), .Z(n9728) );
  XOR U7912 ( .A(n9730), .B(n9731), .Z(n6860) );
  NOR U7913 ( .A(n9732), .B(n9730), .Z(n9731) );
  XOR U7914 ( .A(n9733), .B(n9734), .Z(n6863) );
  NOR U7915 ( .A(n9735), .B(n9733), .Z(n9734) );
  XOR U7916 ( .A(n9736), .B(n9737), .Z(n6866) );
  NOR U7917 ( .A(n9738), .B(n9736), .Z(n9737) );
  XOR U7918 ( .A(n9739), .B(n9740), .Z(n6869) );
  NOR U7919 ( .A(n9741), .B(n9739), .Z(n9740) );
  XOR U7920 ( .A(n9742), .B(n9743), .Z(n6872) );
  NOR U7921 ( .A(n9744), .B(n9742), .Z(n9743) );
  XOR U7922 ( .A(n9745), .B(n9746), .Z(n6875) );
  NOR U7923 ( .A(n9747), .B(n9745), .Z(n9746) );
  XOR U7924 ( .A(n9748), .B(n9749), .Z(n6878) );
  NOR U7925 ( .A(n9750), .B(n9748), .Z(n9749) );
  XOR U7926 ( .A(n9751), .B(n9752), .Z(n6881) );
  NOR U7927 ( .A(n9753), .B(n9751), .Z(n9752) );
  XOR U7928 ( .A(n9754), .B(n9755), .Z(n6884) );
  NOR U7929 ( .A(n9756), .B(n9754), .Z(n9755) );
  XOR U7930 ( .A(n9757), .B(n9758), .Z(n6887) );
  NOR U7931 ( .A(n9759), .B(n9757), .Z(n9758) );
  XOR U7932 ( .A(n9760), .B(n9761), .Z(n6890) );
  NOR U7933 ( .A(n9762), .B(n9760), .Z(n9761) );
  XOR U7934 ( .A(n9763), .B(n9764), .Z(n6893) );
  NOR U7935 ( .A(n9765), .B(n9763), .Z(n9764) );
  XOR U7936 ( .A(n9766), .B(n9767), .Z(n6896) );
  NOR U7937 ( .A(n9768), .B(n9766), .Z(n9767) );
  XOR U7938 ( .A(n9769), .B(n9770), .Z(n6899) );
  NOR U7939 ( .A(n9771), .B(n9769), .Z(n9770) );
  XOR U7940 ( .A(n9772), .B(n9773), .Z(n6902) );
  NOR U7941 ( .A(n9774), .B(n9772), .Z(n9773) );
  XOR U7942 ( .A(n9775), .B(n9776), .Z(n6905) );
  NOR U7943 ( .A(n9777), .B(n9775), .Z(n9776) );
  XOR U7944 ( .A(n9778), .B(n9779), .Z(n6908) );
  NOR U7945 ( .A(n9780), .B(n9778), .Z(n9779) );
  XOR U7946 ( .A(n9781), .B(n9782), .Z(n6911) );
  NOR U7947 ( .A(n9783), .B(n9781), .Z(n9782) );
  XOR U7948 ( .A(n9784), .B(n9785), .Z(n6914) );
  NOR U7949 ( .A(n9786), .B(n9784), .Z(n9785) );
  XOR U7950 ( .A(n9787), .B(n9788), .Z(n6917) );
  NOR U7951 ( .A(n9789), .B(n9787), .Z(n9788) );
  XOR U7952 ( .A(n9790), .B(n9791), .Z(n6920) );
  NOR U7953 ( .A(n9792), .B(n9790), .Z(n9791) );
  XOR U7954 ( .A(n9793), .B(n9794), .Z(n6923) );
  NOR U7955 ( .A(n9795), .B(n9793), .Z(n9794) );
  XOR U7956 ( .A(n9796), .B(n9797), .Z(n6926) );
  NOR U7957 ( .A(n9798), .B(n9796), .Z(n9797) );
  XOR U7958 ( .A(n9799), .B(n9800), .Z(n6929) );
  NOR U7959 ( .A(n9801), .B(n9799), .Z(n9800) );
  XOR U7960 ( .A(n9802), .B(n9803), .Z(n6932) );
  NOR U7961 ( .A(n9804), .B(n9802), .Z(n9803) );
  XOR U7962 ( .A(n9805), .B(n9806), .Z(n6935) );
  NOR U7963 ( .A(n9807), .B(n9805), .Z(n9806) );
  XOR U7964 ( .A(n9808), .B(n9809), .Z(n6938) );
  NOR U7965 ( .A(n9810), .B(n9808), .Z(n9809) );
  XOR U7966 ( .A(n9811), .B(n9812), .Z(n6941) );
  NOR U7967 ( .A(n9813), .B(n9811), .Z(n9812) );
  XOR U7968 ( .A(n9814), .B(n9815), .Z(n6944) );
  NOR U7969 ( .A(n9816), .B(n9814), .Z(n9815) );
  XOR U7970 ( .A(n9817), .B(n9818), .Z(n6947) );
  NOR U7971 ( .A(n9819), .B(n9817), .Z(n9818) );
  XOR U7972 ( .A(n9820), .B(n9821), .Z(n6950) );
  NOR U7973 ( .A(n9822), .B(n9820), .Z(n9821) );
  XOR U7974 ( .A(n9823), .B(n9824), .Z(n6953) );
  NOR U7975 ( .A(n9825), .B(n9823), .Z(n9824) );
  XOR U7976 ( .A(n9826), .B(n9827), .Z(n6956) );
  NOR U7977 ( .A(n9828), .B(n9826), .Z(n9827) );
  XOR U7978 ( .A(n9829), .B(n9830), .Z(n6959) );
  NOR U7979 ( .A(n9831), .B(n9829), .Z(n9830) );
  XOR U7980 ( .A(n9832), .B(n9833), .Z(n6962) );
  NOR U7981 ( .A(n9834), .B(n9832), .Z(n9833) );
  XOR U7982 ( .A(n9835), .B(n9836), .Z(n6965) );
  NOR U7983 ( .A(n9837), .B(n9835), .Z(n9836) );
  XOR U7984 ( .A(n9838), .B(n9839), .Z(n6968) );
  NOR U7985 ( .A(n9840), .B(n9838), .Z(n9839) );
  XOR U7986 ( .A(n9841), .B(n9842), .Z(n6971) );
  NOR U7987 ( .A(n9843), .B(n9841), .Z(n9842) );
  XOR U7988 ( .A(n9844), .B(n9845), .Z(n6974) );
  NOR U7989 ( .A(n9846), .B(n9844), .Z(n9845) );
  XOR U7990 ( .A(n9847), .B(n9848), .Z(n6977) );
  NOR U7991 ( .A(n9849), .B(n9847), .Z(n9848) );
  XOR U7992 ( .A(n9850), .B(n9851), .Z(n6980) );
  NOR U7993 ( .A(n9852), .B(n9850), .Z(n9851) );
  XOR U7994 ( .A(n9853), .B(n9854), .Z(n6983) );
  NOR U7995 ( .A(n9855), .B(n9853), .Z(n9854) );
  XOR U7996 ( .A(n9856), .B(n9857), .Z(n6986) );
  NOR U7997 ( .A(n9858), .B(n9856), .Z(n9857) );
  XOR U7998 ( .A(n9859), .B(n9860), .Z(n6989) );
  NOR U7999 ( .A(n9861), .B(n9859), .Z(n9860) );
  XOR U8000 ( .A(n9862), .B(n9863), .Z(n6992) );
  NOR U8001 ( .A(n9864), .B(n9862), .Z(n9863) );
  XOR U8002 ( .A(n9865), .B(n9866), .Z(n6995) );
  NOR U8003 ( .A(n9867), .B(n9865), .Z(n9866) );
  XOR U8004 ( .A(n9868), .B(n9869), .Z(n6998) );
  NOR U8005 ( .A(n9870), .B(n9868), .Z(n9869) );
  XOR U8006 ( .A(n9871), .B(n9872), .Z(n7001) );
  NOR U8007 ( .A(n9873), .B(n9871), .Z(n9872) );
  XOR U8008 ( .A(n9874), .B(n9875), .Z(n7004) );
  NOR U8009 ( .A(n9876), .B(n9874), .Z(n9875) );
  XOR U8010 ( .A(n9877), .B(n9878), .Z(n7007) );
  NOR U8011 ( .A(n9879), .B(n9877), .Z(n9878) );
  XOR U8012 ( .A(n9880), .B(n9881), .Z(n7010) );
  NOR U8013 ( .A(n9882), .B(n9880), .Z(n9881) );
  XOR U8014 ( .A(n9883), .B(n9884), .Z(n7013) );
  NOR U8015 ( .A(n9885), .B(n9883), .Z(n9884) );
  XOR U8016 ( .A(n9886), .B(n9887), .Z(n7016) );
  AND U8017 ( .A(n9888), .B(n9886), .Z(n9887) );
  XOR U8018 ( .A(n9889), .B(n9890), .Z(n7019) );
  AND U8019 ( .A(n89), .B(n9889), .Z(n9890) );
  XNOR U8020 ( .A(n9891), .B(n8473), .Z(n8475) );
  IV U8021 ( .A(n72), .Z(n9891) );
  XOR U8022 ( .A(n8470), .B(n8469), .Z(n72) );
  XNOR U8023 ( .A(n8467), .B(n8466), .Z(n8469) );
  XNOR U8024 ( .A(n8464), .B(n8463), .Z(n8466) );
  XNOR U8025 ( .A(n8461), .B(n8460), .Z(n8463) );
  XNOR U8026 ( .A(n8458), .B(n8457), .Z(n8460) );
  XNOR U8027 ( .A(n8455), .B(n8454), .Z(n8457) );
  XNOR U8028 ( .A(n8452), .B(n8451), .Z(n8454) );
  XNOR U8029 ( .A(n8449), .B(n8448), .Z(n8451) );
  XNOR U8030 ( .A(n8446), .B(n8445), .Z(n8448) );
  XNOR U8031 ( .A(n8443), .B(n8442), .Z(n8445) );
  XNOR U8032 ( .A(n8440), .B(n8439), .Z(n8442) );
  XNOR U8033 ( .A(n8437), .B(n8436), .Z(n8439) );
  XNOR U8034 ( .A(n8434), .B(n8433), .Z(n8436) );
  XNOR U8035 ( .A(n8431), .B(n8430), .Z(n8433) );
  XNOR U8036 ( .A(n8428), .B(n8427), .Z(n8430) );
  XNOR U8037 ( .A(n8425), .B(n8424), .Z(n8427) );
  XNOR U8038 ( .A(n8422), .B(n8421), .Z(n8424) );
  XNOR U8039 ( .A(n8419), .B(n8418), .Z(n8421) );
  XNOR U8040 ( .A(n8416), .B(n8415), .Z(n8418) );
  XNOR U8041 ( .A(n8413), .B(n8412), .Z(n8415) );
  XNOR U8042 ( .A(n8410), .B(n8409), .Z(n8412) );
  XNOR U8043 ( .A(n8407), .B(n8406), .Z(n8409) );
  XNOR U8044 ( .A(n8404), .B(n8403), .Z(n8406) );
  XNOR U8045 ( .A(n8401), .B(n8400), .Z(n8403) );
  XNOR U8046 ( .A(n8398), .B(n8397), .Z(n8400) );
  XNOR U8047 ( .A(n8395), .B(n8394), .Z(n8397) );
  XNOR U8048 ( .A(n8392), .B(n8391), .Z(n8394) );
  XNOR U8049 ( .A(n8389), .B(n8388), .Z(n8391) );
  XNOR U8050 ( .A(n8386), .B(n8385), .Z(n8388) );
  XNOR U8051 ( .A(n8383), .B(n8382), .Z(n8385) );
  XNOR U8052 ( .A(n8380), .B(n8379), .Z(n8382) );
  XNOR U8053 ( .A(n8377), .B(n8376), .Z(n8379) );
  XNOR U8054 ( .A(n8374), .B(n8373), .Z(n8376) );
  XNOR U8055 ( .A(n8371), .B(n8370), .Z(n8373) );
  XNOR U8056 ( .A(n8368), .B(n8367), .Z(n8370) );
  XNOR U8057 ( .A(n8365), .B(n8364), .Z(n8367) );
  XNOR U8058 ( .A(n8362), .B(n8361), .Z(n8364) );
  XNOR U8059 ( .A(n8359), .B(n8358), .Z(n8361) );
  XNOR U8060 ( .A(n8356), .B(n8355), .Z(n8358) );
  XNOR U8061 ( .A(n8353), .B(n8352), .Z(n8355) );
  XNOR U8062 ( .A(n8350), .B(n8349), .Z(n8352) );
  XNOR U8063 ( .A(n8347), .B(n8346), .Z(n8349) );
  XNOR U8064 ( .A(n8344), .B(n8343), .Z(n8346) );
  XNOR U8065 ( .A(n8341), .B(n8340), .Z(n8343) );
  XNOR U8066 ( .A(n8338), .B(n8337), .Z(n8340) );
  XNOR U8067 ( .A(n8335), .B(n8334), .Z(n8337) );
  XNOR U8068 ( .A(n8332), .B(n8331), .Z(n8334) );
  XNOR U8069 ( .A(n8329), .B(n8328), .Z(n8331) );
  XNOR U8070 ( .A(n8326), .B(n8325), .Z(n8328) );
  XNOR U8071 ( .A(n8323), .B(n8322), .Z(n8325) );
  XNOR U8072 ( .A(n8320), .B(n8319), .Z(n8322) );
  XNOR U8073 ( .A(n8317), .B(n8316), .Z(n8319) );
  XNOR U8074 ( .A(n8314), .B(n8313), .Z(n8316) );
  XNOR U8075 ( .A(n8311), .B(n8310), .Z(n8313) );
  XNOR U8076 ( .A(n8308), .B(n8307), .Z(n8310) );
  XNOR U8077 ( .A(n8305), .B(n8304), .Z(n8307) );
  XNOR U8078 ( .A(n8302), .B(n8301), .Z(n8304) );
  XNOR U8079 ( .A(n8299), .B(n8298), .Z(n8301) );
  XNOR U8080 ( .A(n8296), .B(n8295), .Z(n8298) );
  XNOR U8081 ( .A(n8293), .B(n8292), .Z(n8295) );
  XNOR U8082 ( .A(n8290), .B(n8289), .Z(n8292) );
  XNOR U8083 ( .A(n8287), .B(n8286), .Z(n8289) );
  XNOR U8084 ( .A(n8284), .B(n8283), .Z(n8286) );
  XNOR U8085 ( .A(n8281), .B(n8280), .Z(n8283) );
  XNOR U8086 ( .A(n8278), .B(n8277), .Z(n8280) );
  XNOR U8087 ( .A(n8275), .B(n8274), .Z(n8277) );
  XNOR U8088 ( .A(n8272), .B(n8271), .Z(n8274) );
  XNOR U8089 ( .A(n8269), .B(n8268), .Z(n8271) );
  XNOR U8090 ( .A(n8266), .B(n8265), .Z(n8268) );
  XNOR U8091 ( .A(n8263), .B(n8262), .Z(n8265) );
  XNOR U8092 ( .A(n8260), .B(n8259), .Z(n8262) );
  XNOR U8093 ( .A(n8257), .B(n8256), .Z(n8259) );
  XNOR U8094 ( .A(n8254), .B(n8253), .Z(n8256) );
  XNOR U8095 ( .A(n8251), .B(n8250), .Z(n8253) );
  XNOR U8096 ( .A(n8248), .B(n8247), .Z(n8250) );
  XNOR U8097 ( .A(n8245), .B(n8244), .Z(n8247) );
  XNOR U8098 ( .A(n8242), .B(n8241), .Z(n8244) );
  XNOR U8099 ( .A(n8239), .B(n8238), .Z(n8241) );
  XNOR U8100 ( .A(n8236), .B(n8235), .Z(n8238) );
  XNOR U8101 ( .A(n8233), .B(n8232), .Z(n8235) );
  XNOR U8102 ( .A(n8230), .B(n8229), .Z(n8232) );
  XNOR U8103 ( .A(n8227), .B(n8226), .Z(n8229) );
  XNOR U8104 ( .A(n8224), .B(n8223), .Z(n8226) );
  XNOR U8105 ( .A(n8221), .B(n8220), .Z(n8223) );
  XNOR U8106 ( .A(n8218), .B(n8217), .Z(n8220) );
  XNOR U8107 ( .A(n8215), .B(n8214), .Z(n8217) );
  XNOR U8108 ( .A(n8212), .B(n8211), .Z(n8214) );
  XNOR U8109 ( .A(n8209), .B(n8208), .Z(n8211) );
  XNOR U8110 ( .A(n8206), .B(n8205), .Z(n8208) );
  XNOR U8111 ( .A(n8203), .B(n8202), .Z(n8205) );
  XNOR U8112 ( .A(n8200), .B(n8199), .Z(n8202) );
  XNOR U8113 ( .A(n8197), .B(n8196), .Z(n8199) );
  XNOR U8114 ( .A(n8194), .B(n8193), .Z(n8196) );
  XNOR U8115 ( .A(n8191), .B(n8190), .Z(n8193) );
  XNOR U8116 ( .A(n8188), .B(n8187), .Z(n8190) );
  XNOR U8117 ( .A(n8185), .B(n8184), .Z(n8187) );
  XNOR U8118 ( .A(n8182), .B(n8181), .Z(n8184) );
  XNOR U8119 ( .A(n8179), .B(n8178), .Z(n8181) );
  XNOR U8120 ( .A(n8176), .B(n8175), .Z(n8178) );
  XNOR U8121 ( .A(n8173), .B(n8172), .Z(n8175) );
  XNOR U8122 ( .A(n8170), .B(n8169), .Z(n8172) );
  XNOR U8123 ( .A(n8167), .B(n8166), .Z(n8169) );
  XNOR U8124 ( .A(n8164), .B(n8163), .Z(n8166) );
  XNOR U8125 ( .A(n8161), .B(n8160), .Z(n8163) );
  XNOR U8126 ( .A(n8158), .B(n8157), .Z(n8160) );
  XNOR U8127 ( .A(n8155), .B(n8154), .Z(n8157) );
  XNOR U8128 ( .A(n8152), .B(n8151), .Z(n8154) );
  XNOR U8129 ( .A(n8149), .B(n8148), .Z(n8151) );
  XNOR U8130 ( .A(n8146), .B(n8145), .Z(n8148) );
  XNOR U8131 ( .A(n8143), .B(n8142), .Z(n8145) );
  XNOR U8132 ( .A(n8140), .B(n8139), .Z(n8142) );
  XNOR U8133 ( .A(n8137), .B(n8136), .Z(n8139) );
  XNOR U8134 ( .A(n8134), .B(n8133), .Z(n8136) );
  XNOR U8135 ( .A(n8131), .B(n8130), .Z(n8133) );
  XNOR U8136 ( .A(n8128), .B(n8127), .Z(n8130) );
  XNOR U8137 ( .A(n8125), .B(n8124), .Z(n8127) );
  XNOR U8138 ( .A(n8122), .B(n8121), .Z(n8124) );
  XNOR U8139 ( .A(n8119), .B(n8118), .Z(n8121) );
  XNOR U8140 ( .A(n8116), .B(n8115), .Z(n8118) );
  XNOR U8141 ( .A(n8113), .B(n8112), .Z(n8115) );
  XNOR U8142 ( .A(n8110), .B(n8109), .Z(n8112) );
  XNOR U8143 ( .A(n8107), .B(n8106), .Z(n8109) );
  XNOR U8144 ( .A(n8104), .B(n8103), .Z(n8106) );
  XNOR U8145 ( .A(n8101), .B(n8100), .Z(n8103) );
  XNOR U8146 ( .A(n8098), .B(n8097), .Z(n8100) );
  XNOR U8147 ( .A(n8095), .B(n8094), .Z(n8097) );
  XNOR U8148 ( .A(n8092), .B(n8091), .Z(n8094) );
  XNOR U8149 ( .A(n8089), .B(n8088), .Z(n8091) );
  XNOR U8150 ( .A(n8086), .B(n8085), .Z(n8088) );
  XNOR U8151 ( .A(n8083), .B(n8082), .Z(n8085) );
  XNOR U8152 ( .A(n8080), .B(n8079), .Z(n8082) );
  XNOR U8153 ( .A(n8077), .B(n8076), .Z(n8079) );
  XNOR U8154 ( .A(n8074), .B(n8073), .Z(n8076) );
  XNOR U8155 ( .A(n8071), .B(n8070), .Z(n8073) );
  XNOR U8156 ( .A(n8068), .B(n8067), .Z(n8070) );
  XNOR U8157 ( .A(n8065), .B(n8064), .Z(n8067) );
  XNOR U8158 ( .A(n8062), .B(n8061), .Z(n8064) );
  XNOR U8159 ( .A(n8059), .B(n8058), .Z(n8061) );
  XNOR U8160 ( .A(n8056), .B(n8055), .Z(n8058) );
  XNOR U8161 ( .A(n8053), .B(n8052), .Z(n8055) );
  XNOR U8162 ( .A(n8050), .B(n8049), .Z(n8052) );
  XNOR U8163 ( .A(n8047), .B(n8046), .Z(n8049) );
  XNOR U8164 ( .A(n8044), .B(n8043), .Z(n8046) );
  XNOR U8165 ( .A(n8041), .B(n8040), .Z(n8043) );
  XNOR U8166 ( .A(n8038), .B(n8037), .Z(n8040) );
  XNOR U8167 ( .A(n8035), .B(n8034), .Z(n8037) );
  XNOR U8168 ( .A(n8032), .B(n8031), .Z(n8034) );
  XNOR U8169 ( .A(n8029), .B(n8028), .Z(n8031) );
  XNOR U8170 ( .A(n8026), .B(n8025), .Z(n8028) );
  XNOR U8171 ( .A(n8023), .B(n8022), .Z(n8025) );
  XNOR U8172 ( .A(n8020), .B(n8019), .Z(n8022) );
  XNOR U8173 ( .A(n8017), .B(n8016), .Z(n8019) );
  XNOR U8174 ( .A(n8014), .B(n8013), .Z(n8016) );
  XNOR U8175 ( .A(n8011), .B(n8010), .Z(n8013) );
  XNOR U8176 ( .A(n8008), .B(n8007), .Z(n8010) );
  XNOR U8177 ( .A(n8005), .B(n8004), .Z(n8007) );
  XNOR U8178 ( .A(n8002), .B(n8001), .Z(n8004) );
  XNOR U8179 ( .A(n7999), .B(n7998), .Z(n8001) );
  XNOR U8180 ( .A(n7996), .B(n7995), .Z(n7998) );
  XNOR U8181 ( .A(n7993), .B(n7992), .Z(n7995) );
  XNOR U8182 ( .A(n7990), .B(n7989), .Z(n7992) );
  XNOR U8183 ( .A(n7987), .B(n7986), .Z(n7989) );
  XNOR U8184 ( .A(n7984), .B(n7983), .Z(n7986) );
  XNOR U8185 ( .A(n7981), .B(n7980), .Z(n7983) );
  XNOR U8186 ( .A(n7978), .B(n7977), .Z(n7980) );
  XNOR U8187 ( .A(n7975), .B(n7974), .Z(n7977) );
  XNOR U8188 ( .A(n7972), .B(n7971), .Z(n7974) );
  XNOR U8189 ( .A(n7969), .B(n7968), .Z(n7971) );
  XNOR U8190 ( .A(n7966), .B(n7965), .Z(n7968) );
  XNOR U8191 ( .A(n7963), .B(n7962), .Z(n7965) );
  XNOR U8192 ( .A(n7960), .B(n7959), .Z(n7962) );
  XNOR U8193 ( .A(n7957), .B(n7956), .Z(n7959) );
  XNOR U8194 ( .A(n7954), .B(n7953), .Z(n7956) );
  XNOR U8195 ( .A(n7951), .B(n7950), .Z(n7953) );
  XNOR U8196 ( .A(n7948), .B(n7947), .Z(n7950) );
  XNOR U8197 ( .A(n7945), .B(n7944), .Z(n7947) );
  XNOR U8198 ( .A(n7942), .B(n7941), .Z(n7944) );
  XNOR U8199 ( .A(n7939), .B(n7938), .Z(n7941) );
  XNOR U8200 ( .A(n7936), .B(n7935), .Z(n7938) );
  XNOR U8201 ( .A(n7933), .B(n7932), .Z(n7935) );
  XNOR U8202 ( .A(n7930), .B(n7929), .Z(n7932) );
  XNOR U8203 ( .A(n7927), .B(n7926), .Z(n7929) );
  XNOR U8204 ( .A(n7924), .B(n7923), .Z(n7926) );
  XNOR U8205 ( .A(n7921), .B(n7920), .Z(n7923) );
  XNOR U8206 ( .A(n7918), .B(n7917), .Z(n7920) );
  XNOR U8207 ( .A(n7915), .B(n7914), .Z(n7917) );
  XNOR U8208 ( .A(n7912), .B(n7911), .Z(n7914) );
  XNOR U8209 ( .A(n7909), .B(n7908), .Z(n7911) );
  XNOR U8210 ( .A(n7906), .B(n7905), .Z(n7908) );
  XNOR U8211 ( .A(n7903), .B(n7902), .Z(n7905) );
  XNOR U8212 ( .A(n7900), .B(n7899), .Z(n7902) );
  XNOR U8213 ( .A(n7897), .B(n7896), .Z(n7899) );
  XNOR U8214 ( .A(n7894), .B(n7893), .Z(n7896) );
  XNOR U8215 ( .A(n7891), .B(n7890), .Z(n7893) );
  XNOR U8216 ( .A(n7888), .B(n7887), .Z(n7890) );
  XNOR U8217 ( .A(n7885), .B(n7884), .Z(n7887) );
  XNOR U8218 ( .A(n7882), .B(n7881), .Z(n7884) );
  XNOR U8219 ( .A(n7879), .B(n7878), .Z(n7881) );
  XNOR U8220 ( .A(n7876), .B(n7875), .Z(n7878) );
  XNOR U8221 ( .A(n7873), .B(n7872), .Z(n7875) );
  XNOR U8222 ( .A(n7870), .B(n7869), .Z(n7872) );
  XNOR U8223 ( .A(n7867), .B(n7866), .Z(n7869) );
  XNOR U8224 ( .A(n7864), .B(n7863), .Z(n7866) );
  XNOR U8225 ( .A(n7861), .B(n7860), .Z(n7863) );
  XNOR U8226 ( .A(n7858), .B(n7857), .Z(n7860) );
  XNOR U8227 ( .A(n7855), .B(n7854), .Z(n7857) );
  XNOR U8228 ( .A(n7852), .B(n7851), .Z(n7854) );
  XNOR U8229 ( .A(n7849), .B(n7848), .Z(n7851) );
  XNOR U8230 ( .A(n7846), .B(n7845), .Z(n7848) );
  XNOR U8231 ( .A(n7843), .B(n7842), .Z(n7845) );
  XNOR U8232 ( .A(n7840), .B(n7839), .Z(n7842) );
  XNOR U8233 ( .A(n7837), .B(n7836), .Z(n7839) );
  XNOR U8234 ( .A(n7834), .B(n7833), .Z(n7836) );
  XNOR U8235 ( .A(n7831), .B(n7830), .Z(n7833) );
  XNOR U8236 ( .A(n7828), .B(n7827), .Z(n7830) );
  XNOR U8237 ( .A(n7825), .B(n7824), .Z(n7827) );
  XNOR U8238 ( .A(n7822), .B(n7821), .Z(n7824) );
  XNOR U8239 ( .A(n7819), .B(n7818), .Z(n7821) );
  XNOR U8240 ( .A(n7816), .B(n7815), .Z(n7818) );
  XNOR U8241 ( .A(n7813), .B(n7812), .Z(n7815) );
  XNOR U8242 ( .A(n7810), .B(n7809), .Z(n7812) );
  XNOR U8243 ( .A(n7807), .B(n7806), .Z(n7809) );
  XNOR U8244 ( .A(n7804), .B(n7803), .Z(n7806) );
  XNOR U8245 ( .A(n7801), .B(n7800), .Z(n7803) );
  XNOR U8246 ( .A(n7798), .B(n7797), .Z(n7800) );
  XNOR U8247 ( .A(n7795), .B(n7794), .Z(n7797) );
  XNOR U8248 ( .A(n7792), .B(n7791), .Z(n7794) );
  XNOR U8249 ( .A(n7789), .B(n7788), .Z(n7791) );
  XNOR U8250 ( .A(n7786), .B(n7785), .Z(n7788) );
  XNOR U8251 ( .A(n7783), .B(n7782), .Z(n7785) );
  XNOR U8252 ( .A(n7780), .B(n7779), .Z(n7782) );
  XNOR U8253 ( .A(n7777), .B(n7776), .Z(n7779) );
  XNOR U8254 ( .A(n7774), .B(n7773), .Z(n7776) );
  XNOR U8255 ( .A(n7771), .B(n7770), .Z(n7773) );
  XNOR U8256 ( .A(n7768), .B(n7767), .Z(n7770) );
  XNOR U8257 ( .A(n7765), .B(n7764), .Z(n7767) );
  XNOR U8258 ( .A(n7762), .B(n7761), .Z(n7764) );
  XNOR U8259 ( .A(n7759), .B(n7758), .Z(n7761) );
  XNOR U8260 ( .A(n7756), .B(n7755), .Z(n7758) );
  XNOR U8261 ( .A(n7753), .B(n7752), .Z(n7755) );
  XNOR U8262 ( .A(n7750), .B(n7749), .Z(n7752) );
  XNOR U8263 ( .A(n7747), .B(n7746), .Z(n7749) );
  XNOR U8264 ( .A(n7744), .B(n7743), .Z(n7746) );
  XNOR U8265 ( .A(n7741), .B(n7740), .Z(n7743) );
  XNOR U8266 ( .A(n7738), .B(n7737), .Z(n7740) );
  XNOR U8267 ( .A(n7735), .B(n7734), .Z(n7737) );
  XNOR U8268 ( .A(n7732), .B(n7731), .Z(n7734) );
  XNOR U8269 ( .A(n7729), .B(n7728), .Z(n7731) );
  XNOR U8270 ( .A(n7726), .B(n7725), .Z(n7728) );
  XNOR U8271 ( .A(n7723), .B(n7722), .Z(n7725) );
  XNOR U8272 ( .A(n7720), .B(n7719), .Z(n7722) );
  XNOR U8273 ( .A(n7717), .B(n7716), .Z(n7719) );
  XNOR U8274 ( .A(n7714), .B(n7713), .Z(n7716) );
  XNOR U8275 ( .A(n7711), .B(n7710), .Z(n7713) );
  XNOR U8276 ( .A(n7708), .B(n7707), .Z(n7710) );
  XNOR U8277 ( .A(n7705), .B(n7704), .Z(n7707) );
  XNOR U8278 ( .A(n7702), .B(n7701), .Z(n7704) );
  XNOR U8279 ( .A(n7699), .B(n7698), .Z(n7701) );
  XNOR U8280 ( .A(n7696), .B(n7695), .Z(n7698) );
  XNOR U8281 ( .A(n7693), .B(n7692), .Z(n7695) );
  XNOR U8282 ( .A(n7690), .B(n7689), .Z(n7692) );
  XNOR U8283 ( .A(n7687), .B(n7686), .Z(n7689) );
  XNOR U8284 ( .A(n7684), .B(n7683), .Z(n7686) );
  XNOR U8285 ( .A(n7681), .B(n7680), .Z(n7683) );
  XNOR U8286 ( .A(n7678), .B(n7677), .Z(n7680) );
  XNOR U8287 ( .A(n7675), .B(n7674), .Z(n7677) );
  XNOR U8288 ( .A(n7672), .B(n7671), .Z(n7674) );
  XNOR U8289 ( .A(n7669), .B(n7668), .Z(n7671) );
  XNOR U8290 ( .A(n7666), .B(n7665), .Z(n7668) );
  XNOR U8291 ( .A(n7663), .B(n7662), .Z(n7665) );
  XNOR U8292 ( .A(n7660), .B(n7659), .Z(n7662) );
  XNOR U8293 ( .A(n7657), .B(n7656), .Z(n7659) );
  XNOR U8294 ( .A(n7654), .B(n7653), .Z(n7656) );
  XNOR U8295 ( .A(n7651), .B(n7650), .Z(n7653) );
  XNOR U8296 ( .A(n7648), .B(n7647), .Z(n7650) );
  XNOR U8297 ( .A(n7645), .B(n7644), .Z(n7647) );
  XNOR U8298 ( .A(n7642), .B(n7641), .Z(n7644) );
  XNOR U8299 ( .A(n7639), .B(n7638), .Z(n7641) );
  XNOR U8300 ( .A(n7636), .B(n7635), .Z(n7638) );
  XNOR U8301 ( .A(n7633), .B(n7632), .Z(n7635) );
  XNOR U8302 ( .A(n7630), .B(n7629), .Z(n7632) );
  XNOR U8303 ( .A(n7627), .B(n7626), .Z(n7629) );
  XNOR U8304 ( .A(n7624), .B(n7623), .Z(n7626) );
  XNOR U8305 ( .A(n7621), .B(n7620), .Z(n7623) );
  XNOR U8306 ( .A(n7618), .B(n7617), .Z(n7620) );
  XNOR U8307 ( .A(n7615), .B(n7614), .Z(n7617) );
  XNOR U8308 ( .A(n7612), .B(n7611), .Z(n7614) );
  XNOR U8309 ( .A(n7609), .B(n7608), .Z(n7611) );
  XNOR U8310 ( .A(n7606), .B(n7605), .Z(n7608) );
  XNOR U8311 ( .A(n7603), .B(n7602), .Z(n7605) );
  XNOR U8312 ( .A(n7600), .B(n7599), .Z(n7602) );
  XNOR U8313 ( .A(n7597), .B(n7596), .Z(n7599) );
  XNOR U8314 ( .A(n7594), .B(n7593), .Z(n7596) );
  XNOR U8315 ( .A(n7591), .B(n7590), .Z(n7593) );
  XNOR U8316 ( .A(n7588), .B(n7587), .Z(n7590) );
  XNOR U8317 ( .A(n7585), .B(n7584), .Z(n7587) );
  XNOR U8318 ( .A(n7582), .B(n7581), .Z(n7584) );
  XNOR U8319 ( .A(n7579), .B(n7578), .Z(n7581) );
  XNOR U8320 ( .A(n7576), .B(n7575), .Z(n7578) );
  XNOR U8321 ( .A(n7573), .B(n7572), .Z(n7575) );
  XNOR U8322 ( .A(n7570), .B(n7569), .Z(n7572) );
  XNOR U8323 ( .A(n7567), .B(n7566), .Z(n7569) );
  XNOR U8324 ( .A(n7564), .B(n7563), .Z(n7566) );
  XNOR U8325 ( .A(n7561), .B(n7560), .Z(n7563) );
  XNOR U8326 ( .A(n7558), .B(n7557), .Z(n7560) );
  XNOR U8327 ( .A(n7555), .B(n7554), .Z(n7557) );
  XNOR U8328 ( .A(n7552), .B(n7551), .Z(n7554) );
  XNOR U8329 ( .A(n7549), .B(n7548), .Z(n7551) );
  XNOR U8330 ( .A(n7546), .B(n7545), .Z(n7548) );
  XNOR U8331 ( .A(n7543), .B(n7542), .Z(n7545) );
  XNOR U8332 ( .A(n7540), .B(n7539), .Z(n7542) );
  XNOR U8333 ( .A(n7537), .B(n7536), .Z(n7539) );
  XNOR U8334 ( .A(n7534), .B(n7533), .Z(n7536) );
  XNOR U8335 ( .A(n7531), .B(n7530), .Z(n7533) );
  XNOR U8336 ( .A(n7528), .B(n7527), .Z(n7530) );
  XNOR U8337 ( .A(n7525), .B(n7524), .Z(n7527) );
  XNOR U8338 ( .A(n7522), .B(n7521), .Z(n7524) );
  XNOR U8339 ( .A(n7519), .B(n7518), .Z(n7521) );
  XNOR U8340 ( .A(n7516), .B(n7515), .Z(n7518) );
  XNOR U8341 ( .A(n7513), .B(n7512), .Z(n7515) );
  XNOR U8342 ( .A(n7510), .B(n7509), .Z(n7512) );
  XNOR U8343 ( .A(n7507), .B(n7506), .Z(n7509) );
  XNOR U8344 ( .A(n7504), .B(n7503), .Z(n7506) );
  XNOR U8345 ( .A(n7501), .B(n7500), .Z(n7503) );
  XNOR U8346 ( .A(n7498), .B(n7497), .Z(n7500) );
  XNOR U8347 ( .A(n7495), .B(n7494), .Z(n7497) );
  XNOR U8348 ( .A(n7492), .B(n7491), .Z(n7494) );
  XNOR U8349 ( .A(n7489), .B(n7488), .Z(n7491) );
  XNOR U8350 ( .A(n7486), .B(n7485), .Z(n7488) );
  XNOR U8351 ( .A(n7483), .B(n7482), .Z(n7485) );
  XNOR U8352 ( .A(n7480), .B(n7479), .Z(n7482) );
  XNOR U8353 ( .A(n7477), .B(n7476), .Z(n7479) );
  XNOR U8354 ( .A(n7474), .B(n7473), .Z(n7476) );
  XNOR U8355 ( .A(n7471), .B(n7470), .Z(n7473) );
  XNOR U8356 ( .A(n7468), .B(n7467), .Z(n7470) );
  XNOR U8357 ( .A(n7465), .B(n7464), .Z(n7467) );
  XNOR U8358 ( .A(n7462), .B(n7461), .Z(n7464) );
  XNOR U8359 ( .A(n7459), .B(n7458), .Z(n7461) );
  XNOR U8360 ( .A(n7456), .B(n7455), .Z(n7458) );
  XNOR U8361 ( .A(n7453), .B(n7452), .Z(n7455) );
  XNOR U8362 ( .A(n7450), .B(n7449), .Z(n7452) );
  XNOR U8363 ( .A(n7447), .B(n7446), .Z(n7449) );
  XNOR U8364 ( .A(n7444), .B(n7443), .Z(n7446) );
  XNOR U8365 ( .A(n7441), .B(n7440), .Z(n7443) );
  XNOR U8366 ( .A(n7438), .B(n7437), .Z(n7440) );
  XNOR U8367 ( .A(n7435), .B(n7434), .Z(n7437) );
  XNOR U8368 ( .A(n7432), .B(n7431), .Z(n7434) );
  XNOR U8369 ( .A(n7429), .B(n7428), .Z(n7431) );
  XNOR U8370 ( .A(n7426), .B(n7425), .Z(n7428) );
  XNOR U8371 ( .A(n7423), .B(n7422), .Z(n7425) );
  XNOR U8372 ( .A(n7420), .B(n7419), .Z(n7422) );
  XNOR U8373 ( .A(n7417), .B(n7416), .Z(n7419) );
  XNOR U8374 ( .A(n7414), .B(n7413), .Z(n7416) );
  XNOR U8375 ( .A(n7411), .B(n7410), .Z(n7413) );
  XNOR U8376 ( .A(n7408), .B(n7407), .Z(n7410) );
  XNOR U8377 ( .A(n7405), .B(n7404), .Z(n7407) );
  XNOR U8378 ( .A(n7402), .B(n7401), .Z(n7404) );
  XNOR U8379 ( .A(n7399), .B(n7398), .Z(n7401) );
  XNOR U8380 ( .A(n7396), .B(n7395), .Z(n7398) );
  XNOR U8381 ( .A(n7393), .B(n7392), .Z(n7395) );
  XNOR U8382 ( .A(n7390), .B(n7389), .Z(n7392) );
  XNOR U8383 ( .A(n7387), .B(n7386), .Z(n7389) );
  XNOR U8384 ( .A(n7384), .B(n7383), .Z(n7386) );
  XNOR U8385 ( .A(n7381), .B(n7380), .Z(n7383) );
  XNOR U8386 ( .A(n7378), .B(n7377), .Z(n7380) );
  XNOR U8387 ( .A(n7375), .B(n7374), .Z(n7377) );
  XNOR U8388 ( .A(n7372), .B(n7371), .Z(n7374) );
  XNOR U8389 ( .A(n7369), .B(n7368), .Z(n7371) );
  XNOR U8390 ( .A(n7366), .B(n7365), .Z(n7368) );
  XNOR U8391 ( .A(n7363), .B(n7362), .Z(n7365) );
  XNOR U8392 ( .A(n7360), .B(n7359), .Z(n7362) );
  XNOR U8393 ( .A(n7357), .B(n7356), .Z(n7359) );
  XNOR U8394 ( .A(n7354), .B(n7353), .Z(n7356) );
  XNOR U8395 ( .A(n7351), .B(n7350), .Z(n7353) );
  XNOR U8396 ( .A(n7348), .B(n7347), .Z(n7350) );
  XNOR U8397 ( .A(n7345), .B(n7344), .Z(n7347) );
  XNOR U8398 ( .A(n7342), .B(n7341), .Z(n7344) );
  XNOR U8399 ( .A(n7339), .B(n7338), .Z(n7341) );
  XNOR U8400 ( .A(n7336), .B(n7335), .Z(n7338) );
  XNOR U8401 ( .A(n7333), .B(n7332), .Z(n7335) );
  XNOR U8402 ( .A(n7330), .B(n7329), .Z(n7332) );
  XNOR U8403 ( .A(n7327), .B(n7326), .Z(n7329) );
  XNOR U8404 ( .A(n7324), .B(n7323), .Z(n7326) );
  XNOR U8405 ( .A(n7321), .B(n7320), .Z(n7323) );
  XOR U8406 ( .A(n7318), .B(n7045), .Z(n7320) );
  XOR U8407 ( .A(n9892), .B(n7033), .Z(n7045) );
  XNOR U8408 ( .A(n7034), .B(n7031), .Z(n7033) );
  XNOR U8409 ( .A(n7032), .B(n7028), .Z(n7031) );
  XNOR U8410 ( .A(n7027), .B(n7054), .Z(n7028) );
  XNOR U8411 ( .A(n7053), .B(n7317), .Z(n7054) );
  XNOR U8412 ( .A(n7308), .B(n7316), .Z(n7317) );
  XNOR U8413 ( .A(n7307), .B(n7313), .Z(n7316) );
  XNOR U8414 ( .A(n7312), .B(n7295), .Z(n7313) );
  XNOR U8415 ( .A(n7060), .B(n7306), .Z(n7295) );
  XNOR U8416 ( .A(n7297), .B(n7305), .Z(n7306) );
  XOR U8417 ( .A(n7296), .B(n7302), .Z(n7305) );
  XOR U8418 ( .A(n7301), .B(n7285), .Z(n7302) );
  XOR U8419 ( .A(n7063), .B(n7294), .Z(n7285) );
  XOR U8420 ( .A(n7281), .B(n7291), .Z(n7294) );
  XOR U8421 ( .A(n7284), .B(n7290), .Z(n7291) );
  XOR U8422 ( .A(n7280), .B(n7059), .Z(n7290) );
  AND U8423 ( .A(n9893), .B(n9894), .Z(n7059) );
  XOR U8424 ( .A(n7279), .B(n7275), .Z(n7280) );
  AND U8425 ( .A(n9895), .B(n9896), .Z(n7275) );
  XOR U8426 ( .A(n7276), .B(n7269), .Z(n7279) );
  AND U8427 ( .A(n9897), .B(n9898), .Z(n7269) );
  XNOR U8428 ( .A(n7270), .B(n7268), .Z(n7276) );
  AND U8429 ( .A(n9899), .B(n9900), .Z(n7268) );
  XOR U8430 ( .A(n7221), .B(n7271), .Z(n7270) );
  AND U8431 ( .A(n9901), .B(n9902), .Z(n7271) );
  XNOR U8432 ( .A(n7265), .B(n7222), .Z(n7221) );
  AND U8433 ( .A(n9903), .B(n9904), .Z(n7222) );
  XOR U8434 ( .A(n7264), .B(n7256), .Z(n7265) );
  AND U8435 ( .A(n9905), .B(n9906), .Z(n7256) );
  XNOR U8436 ( .A(n7259), .B(n7255), .Z(n7264) );
  AND U8437 ( .A(n9907), .B(n9908), .Z(n7255) );
  XOR U8438 ( .A(n7225), .B(n7260), .Z(n7259) );
  AND U8439 ( .A(n9909), .B(n9910), .Z(n7260) );
  XNOR U8440 ( .A(n7254), .B(n7226), .Z(n7225) );
  AND U8441 ( .A(n9911), .B(n9912), .Z(n7226) );
  XOR U8442 ( .A(n7253), .B(n7243), .Z(n7254) );
  AND U8443 ( .A(n9913), .B(n9914), .Z(n7243) );
  XNOR U8444 ( .A(n7248), .B(n7242), .Z(n7253) );
  AND U8445 ( .A(n9915), .B(n9916), .Z(n7242) );
  XOR U8446 ( .A(n7185), .B(n7249), .Z(n7248) );
  AND U8447 ( .A(n9917), .B(n9918), .Z(n7249) );
  XNOR U8448 ( .A(n7241), .B(n7186), .Z(n7185) );
  AND U8449 ( .A(n9919), .B(n9920), .Z(n7186) );
  XOR U8450 ( .A(n7240), .B(n7228), .Z(n7241) );
  AND U8451 ( .A(n9921), .B(n9922), .Z(n7228) );
  XNOR U8452 ( .A(n7235), .B(n7227), .Z(n7240) );
  AND U8453 ( .A(n9923), .B(n9924), .Z(n7227) );
  XOR U8454 ( .A(n7189), .B(n7236), .Z(n7235) );
  AND U8455 ( .A(n9925), .B(n9926), .Z(n7236) );
  XNOR U8456 ( .A(n7220), .B(n7190), .Z(n7189) );
  AND U8457 ( .A(n9927), .B(n9928), .Z(n7190) );
  XOR U8458 ( .A(n7219), .B(n7211), .Z(n7220) );
  AND U8459 ( .A(n9929), .B(n9930), .Z(n7211) );
  XNOR U8460 ( .A(n7214), .B(n7210), .Z(n7219) );
  AND U8461 ( .A(n9931), .B(n9932), .Z(n7210) );
  XOR U8462 ( .A(n7191), .B(n7215), .Z(n7214) );
  AND U8463 ( .A(n9933), .B(n9934), .Z(n7215) );
  XNOR U8464 ( .A(n7207), .B(n7192), .Z(n7191) );
  AND U8465 ( .A(n9935), .B(n9936), .Z(n7192) );
  XOR U8466 ( .A(n7206), .B(n7198), .Z(n7207) );
  AND U8467 ( .A(n9937), .B(n9938), .Z(n7198) );
  XNOR U8468 ( .A(n7201), .B(n7197), .Z(n7206) );
  AND U8469 ( .A(n9939), .B(n9940), .Z(n7197) );
  XOR U8470 ( .A(n7142), .B(n7202), .Z(n7201) );
  AND U8471 ( .A(n9941), .B(n9942), .Z(n7202) );
  XNOR U8472 ( .A(n7184), .B(n7143), .Z(n7142) );
  AND U8473 ( .A(n9943), .B(n9944), .Z(n7143) );
  XOR U8474 ( .A(n7183), .B(n7175), .Z(n7184) );
  AND U8475 ( .A(n9945), .B(n9946), .Z(n7175) );
  XNOR U8476 ( .A(n7178), .B(n7174), .Z(n7183) );
  AND U8477 ( .A(n9947), .B(n9948), .Z(n7174) );
  XOR U8478 ( .A(n7146), .B(n7179), .Z(n7178) );
  AND U8479 ( .A(n9949), .B(n9950), .Z(n7179) );
  XNOR U8480 ( .A(n7171), .B(n7147), .Z(n7146) );
  AND U8481 ( .A(n9951), .B(n9952), .Z(n7147) );
  XOR U8482 ( .A(n7170), .B(n7162), .Z(n7171) );
  AND U8483 ( .A(n9953), .B(n9954), .Z(n7162) );
  XNOR U8484 ( .A(n7165), .B(n7161), .Z(n7170) );
  AND U8485 ( .A(n9955), .B(n9956), .Z(n7161) );
  XOR U8486 ( .A(n7095), .B(n7166), .Z(n7165) );
  AND U8487 ( .A(n9957), .B(n9958), .Z(n7166) );
  XNOR U8488 ( .A(n7156), .B(n7096), .Z(n7095) );
  AND U8489 ( .A(n9959), .B(n9960), .Z(n7096) );
  XOR U8490 ( .A(n7155), .B(n7141), .Z(n7156) );
  AND U8491 ( .A(n9961), .B(n9962), .Z(n7141) );
  XNOR U8492 ( .A(n7150), .B(n7140), .Z(n7155) );
  AND U8493 ( .A(n9963), .B(n9964), .Z(n7140) );
  XOR U8494 ( .A(n7097), .B(n7151), .Z(n7150) );
  AND U8495 ( .A(n9965), .B(n9966), .Z(n7151) );
  XNOR U8496 ( .A(n7139), .B(n7098), .Z(n7097) );
  AND U8497 ( .A(n9967), .B(n9968), .Z(n7098) );
  XOR U8498 ( .A(n7138), .B(n7128), .Z(n7139) );
  AND U8499 ( .A(n9969), .B(n9970), .Z(n7128) );
  XNOR U8500 ( .A(n7133), .B(n7127), .Z(n7138) );
  AND U8501 ( .A(n9971), .B(n9972), .Z(n7127) );
  XOR U8502 ( .A(n9973), .B(n7126), .Z(n7133) );
  XOR U8503 ( .A(n7125), .B(n7113), .Z(n7126) );
  AND U8504 ( .A(n9974), .B(n9975), .Z(n7113) );
  XNOR U8505 ( .A(n7120), .B(n7112), .Z(n7125) );
  AND U8506 ( .A(n9976), .B(n9977), .Z(n7112) );
  XOR U8507 ( .A(n9978), .B(n9979), .Z(n7120) );
  XOR U8508 ( .A(n7110), .B(n9980), .Z(n9979) );
  XOR U8509 ( .A(n7106), .B(n7104), .Z(n9980) );
  AND U8510 ( .A(n9981), .B(n9982), .Z(n7104) );
  AND U8511 ( .A(n9983), .B(n9984), .Z(n7106) );
  AND U8512 ( .A(n9985), .B(n9986), .Z(n7110) );
  XNOR U8513 ( .A(n9987), .B(n7107), .Z(n9978) );
  XOR U8514 ( .A(n9988), .B(n9989), .Z(n7107) );
  XOR U8515 ( .A(n9990), .B(n9991), .Z(n9989) );
  XOR U8516 ( .A(n9992), .B(n9993), .Z(n9991) );
  NOR U8517 ( .A(n9994), .B(n9995), .Z(n9993) );
  NOR U8518 ( .A(n9996), .B(n9997), .Z(n9992) );
  AND U8519 ( .A(n9998), .B(n9999), .Z(n9997) );
  IV U8520 ( .A(n10000), .Z(n9996) );
  NOR U8521 ( .A(n10001), .B(n10002), .Z(n10000) );
  AND U8522 ( .A(n9994), .B(n10003), .Z(n10002) );
  AND U8523 ( .A(n9995), .B(n10004), .Z(n10001) );
  NOR U8524 ( .A(n10005), .B(n10006), .Z(n9990) );
  AND U8525 ( .A(n10007), .B(n10008), .Z(n10006) );
  IV U8526 ( .A(n10009), .Z(n10005) );
  NOR U8527 ( .A(n10010), .B(n10011), .Z(n10009) );
  AND U8528 ( .A(n10012), .B(n10013), .Z(n10011) );
  AND U8529 ( .A(n10014), .B(n10015), .Z(n10010) );
  XOR U8530 ( .A(n10016), .B(n10017), .Z(n9988) );
  XOR U8531 ( .A(n10018), .B(n10019), .Z(n10017) );
  XOR U8532 ( .A(n10020), .B(n10021), .Z(n10019) );
  XOR U8533 ( .A(n10022), .B(n10023), .Z(n10021) );
  AND U8534 ( .A(n10024), .B(n10025), .Z(n10023) );
  AND U8535 ( .A(n10026), .B(n10027), .Z(n10022) );
  XOR U8536 ( .A(n10028), .B(n10029), .Z(n10020) );
  AND U8537 ( .A(n10030), .B(n10031), .Z(n10029) );
  AND U8538 ( .A(n10032), .B(n10033), .Z(n10028) );
  AND U8539 ( .A(n10034), .B(n10035), .Z(n10033) );
  AND U8540 ( .A(n10036), .B(n10037), .Z(n10035) );
  NOR U8541 ( .A(n10038), .B(n10039), .Z(n10037) );
  IV U8542 ( .A(n10040), .Z(n10038) );
  NOR U8543 ( .A(n10041), .B(n10042), .Z(n10040) );
  NOR U8544 ( .A(n10043), .B(n10044), .Z(n10036) );
  AND U8545 ( .A(n10045), .B(n10046), .Z(n10034) );
  NOR U8546 ( .A(n10047), .B(n10048), .Z(n10046) );
  NOR U8547 ( .A(n10049), .B(n10050), .Z(n10045) );
  AND U8548 ( .A(n10051), .B(n10052), .Z(n10032) );
  AND U8549 ( .A(n10053), .B(n10054), .Z(n10052) );
  NOR U8550 ( .A(n10055), .B(n10056), .Z(n10054) );
  NOR U8551 ( .A(n10057), .B(n10058), .Z(n10053) );
  AND U8552 ( .A(n10059), .B(n10060), .Z(n10051) );
  NOR U8553 ( .A(n10061), .B(n10062), .Z(n10060) );
  NOR U8554 ( .A(n10063), .B(n10064), .Z(n10059) );
  XOR U8555 ( .A(n10065), .B(n10066), .Z(n10018) );
  XOR U8556 ( .A(n10067), .B(n10068), .Z(n10066) );
  NOR U8557 ( .A(n10069), .B(n10070), .Z(n10068) );
  NOR U8558 ( .A(n10071), .B(n10072), .Z(n10067) );
  AND U8559 ( .A(n10073), .B(n10074), .Z(n10072) );
  IV U8560 ( .A(n10075), .Z(n10071) );
  NOR U8561 ( .A(n10076), .B(n10077), .Z(n10075) );
  AND U8562 ( .A(n10069), .B(n10078), .Z(n10077) );
  AND U8563 ( .A(n10070), .B(n10079), .Z(n10076) );
  XOR U8564 ( .A(n10080), .B(n10081), .Z(n10065) );
  NOR U8565 ( .A(n10082), .B(n10083), .Z(n10081) );
  NOR U8566 ( .A(n10084), .B(n10085), .Z(n10080) );
  AND U8567 ( .A(n10086), .B(n10087), .Z(n10085) );
  IV U8568 ( .A(n10088), .Z(n10084) );
  NOR U8569 ( .A(n10089), .B(n10090), .Z(n10088) );
  AND U8570 ( .A(n10082), .B(n10091), .Z(n10090) );
  AND U8571 ( .A(n10083), .B(n10092), .Z(n10089) );
  XNOR U8572 ( .A(n10093), .B(n10094), .Z(n10016) );
  AND U8573 ( .A(n10095), .B(n10096), .Z(n10094) );
  NOR U8574 ( .A(n10012), .B(n10014), .Z(n10093) );
  XNOR U8575 ( .A(n7111), .B(n7121), .Z(n9987) );
  AND U8576 ( .A(n10097), .B(n10098), .Z(n7121) );
  AND U8577 ( .A(n10099), .B(n10100), .Z(n7111) );
  XOR U8578 ( .A(n7109), .B(n7134), .Z(n9973) );
  AND U8579 ( .A(n10101), .B(n10102), .Z(n7134) );
  IV U8580 ( .A(n10103), .Z(n7109) );
  AND U8581 ( .A(n10104), .B(n10105), .Z(n10103) );
  XOR U8582 ( .A(n10106), .B(n10107), .Z(n7284) );
  AND U8583 ( .A(n10106), .B(n10108), .Z(n10107) );
  XOR U8584 ( .A(n10109), .B(n10110), .Z(n7281) );
  AND U8585 ( .A(n10109), .B(n10111), .Z(n10110) );
  XOR U8586 ( .A(n10112), .B(n10113), .Z(n7063) );
  AND U8587 ( .A(n10112), .B(n10114), .Z(n10113) );
  XOR U8588 ( .A(n10115), .B(n10116), .Z(n7301) );
  AND U8589 ( .A(n10115), .B(n10117), .Z(n10116) );
  XNOR U8590 ( .A(n10118), .B(n10119), .Z(n7296) );
  AND U8591 ( .A(n10118), .B(n10120), .Z(n10119) );
  XNOR U8592 ( .A(n10121), .B(n10122), .Z(n7297) );
  AND U8593 ( .A(n10123), .B(n10121), .Z(n10122) );
  XOR U8594 ( .A(n10124), .B(n10125), .Z(n7060) );
  NOR U8595 ( .A(n10126), .B(n10124), .Z(n10125) );
  XOR U8596 ( .A(n10127), .B(n10128), .Z(n7312) );
  NOR U8597 ( .A(n10129), .B(n10127), .Z(n10128) );
  XOR U8598 ( .A(n10130), .B(n10131), .Z(n7307) );
  NOR U8599 ( .A(n10132), .B(n10130), .Z(n10131) );
  XOR U8600 ( .A(n10133), .B(n10134), .Z(n7308) );
  NOR U8601 ( .A(n10135), .B(n10133), .Z(n10134) );
  XOR U8602 ( .A(n10136), .B(n10137), .Z(n7053) );
  NOR U8603 ( .A(n10138), .B(n10136), .Z(n10137) );
  XOR U8604 ( .A(n10139), .B(n10140), .Z(n7027) );
  NOR U8605 ( .A(n10141), .B(n10139), .Z(n10140) );
  XOR U8606 ( .A(n10142), .B(n10143), .Z(n7032) );
  NOR U8607 ( .A(n10144), .B(n10142), .Z(n10143) );
  XOR U8608 ( .A(n10145), .B(n10146), .Z(n7034) );
  NOR U8609 ( .A(n10147), .B(n10145), .Z(n10146) );
  IV U8610 ( .A(n7044), .Z(n9892) );
  XNOR U8611 ( .A(n10148), .B(n10149), .Z(n7044) );
  NOR U8612 ( .A(n10150), .B(n10148), .Z(n10149) );
  XOR U8613 ( .A(n10151), .B(n10152), .Z(n7318) );
  NOR U8614 ( .A(n10153), .B(n10151), .Z(n10152) );
  XOR U8615 ( .A(n10154), .B(n10155), .Z(n7321) );
  NOR U8616 ( .A(n10156), .B(n10154), .Z(n10155) );
  XOR U8617 ( .A(n10157), .B(n10158), .Z(n7324) );
  NOR U8618 ( .A(n10159), .B(n10157), .Z(n10158) );
  XOR U8619 ( .A(n10160), .B(n10161), .Z(n7327) );
  NOR U8620 ( .A(n10162), .B(n10160), .Z(n10161) );
  XOR U8621 ( .A(n10163), .B(n10164), .Z(n7330) );
  NOR U8622 ( .A(n10165), .B(n10163), .Z(n10164) );
  XOR U8623 ( .A(n10166), .B(n10167), .Z(n7333) );
  NOR U8624 ( .A(n10168), .B(n10166), .Z(n10167) );
  XOR U8625 ( .A(n10169), .B(n10170), .Z(n7336) );
  NOR U8626 ( .A(n10171), .B(n10169), .Z(n10170) );
  XOR U8627 ( .A(n10172), .B(n10173), .Z(n7339) );
  NOR U8628 ( .A(n10174), .B(n10172), .Z(n10173) );
  XOR U8629 ( .A(n10175), .B(n10176), .Z(n7342) );
  NOR U8630 ( .A(n10177), .B(n10175), .Z(n10176) );
  XOR U8631 ( .A(n10178), .B(n10179), .Z(n7345) );
  NOR U8632 ( .A(n10180), .B(n10178), .Z(n10179) );
  XOR U8633 ( .A(n10181), .B(n10182), .Z(n7348) );
  NOR U8634 ( .A(n10183), .B(n10181), .Z(n10182) );
  XOR U8635 ( .A(n10184), .B(n10185), .Z(n7351) );
  NOR U8636 ( .A(n10186), .B(n10184), .Z(n10185) );
  XOR U8637 ( .A(n10187), .B(n10188), .Z(n7354) );
  NOR U8638 ( .A(n10189), .B(n10187), .Z(n10188) );
  XOR U8639 ( .A(n10190), .B(n10191), .Z(n7357) );
  NOR U8640 ( .A(n10192), .B(n10190), .Z(n10191) );
  XOR U8641 ( .A(n10193), .B(n10194), .Z(n7360) );
  NOR U8642 ( .A(n10195), .B(n10193), .Z(n10194) );
  XOR U8643 ( .A(n10196), .B(n10197), .Z(n7363) );
  NOR U8644 ( .A(n10198), .B(n10196), .Z(n10197) );
  XOR U8645 ( .A(n10199), .B(n10200), .Z(n7366) );
  NOR U8646 ( .A(n10201), .B(n10199), .Z(n10200) );
  XOR U8647 ( .A(n10202), .B(n10203), .Z(n7369) );
  NOR U8648 ( .A(n10204), .B(n10202), .Z(n10203) );
  XOR U8649 ( .A(n10205), .B(n10206), .Z(n7372) );
  NOR U8650 ( .A(n10207), .B(n10205), .Z(n10206) );
  XOR U8651 ( .A(n10208), .B(n10209), .Z(n7375) );
  NOR U8652 ( .A(n10210), .B(n10208), .Z(n10209) );
  XOR U8653 ( .A(n10211), .B(n10212), .Z(n7378) );
  NOR U8654 ( .A(n10213), .B(n10211), .Z(n10212) );
  XOR U8655 ( .A(n10214), .B(n10215), .Z(n7381) );
  NOR U8656 ( .A(n10216), .B(n10214), .Z(n10215) );
  XOR U8657 ( .A(n10217), .B(n10218), .Z(n7384) );
  NOR U8658 ( .A(n10219), .B(n10217), .Z(n10218) );
  XOR U8659 ( .A(n10220), .B(n10221), .Z(n7387) );
  NOR U8660 ( .A(n10222), .B(n10220), .Z(n10221) );
  XOR U8661 ( .A(n10223), .B(n10224), .Z(n7390) );
  NOR U8662 ( .A(n10225), .B(n10223), .Z(n10224) );
  XOR U8663 ( .A(n10226), .B(n10227), .Z(n7393) );
  NOR U8664 ( .A(n10228), .B(n10226), .Z(n10227) );
  XOR U8665 ( .A(n10229), .B(n10230), .Z(n7396) );
  NOR U8666 ( .A(n10231), .B(n10229), .Z(n10230) );
  XOR U8667 ( .A(n10232), .B(n10233), .Z(n7399) );
  NOR U8668 ( .A(n10234), .B(n10232), .Z(n10233) );
  XOR U8669 ( .A(n10235), .B(n10236), .Z(n7402) );
  NOR U8670 ( .A(n10237), .B(n10235), .Z(n10236) );
  XOR U8671 ( .A(n10238), .B(n10239), .Z(n7405) );
  NOR U8672 ( .A(n10240), .B(n10238), .Z(n10239) );
  XOR U8673 ( .A(n10241), .B(n10242), .Z(n7408) );
  NOR U8674 ( .A(n10243), .B(n10241), .Z(n10242) );
  XOR U8675 ( .A(n10244), .B(n10245), .Z(n7411) );
  NOR U8676 ( .A(n10246), .B(n10244), .Z(n10245) );
  XOR U8677 ( .A(n10247), .B(n10248), .Z(n7414) );
  NOR U8678 ( .A(n10249), .B(n10247), .Z(n10248) );
  XOR U8679 ( .A(n10250), .B(n10251), .Z(n7417) );
  NOR U8680 ( .A(n10252), .B(n10250), .Z(n10251) );
  XOR U8681 ( .A(n10253), .B(n10254), .Z(n7420) );
  NOR U8682 ( .A(n10255), .B(n10253), .Z(n10254) );
  XOR U8683 ( .A(n10256), .B(n10257), .Z(n7423) );
  NOR U8684 ( .A(n10258), .B(n10256), .Z(n10257) );
  XOR U8685 ( .A(n10259), .B(n10260), .Z(n7426) );
  NOR U8686 ( .A(n10261), .B(n10259), .Z(n10260) );
  XOR U8687 ( .A(n10262), .B(n10263), .Z(n7429) );
  NOR U8688 ( .A(n10264), .B(n10262), .Z(n10263) );
  XOR U8689 ( .A(n10265), .B(n10266), .Z(n7432) );
  NOR U8690 ( .A(n10267), .B(n10265), .Z(n10266) );
  XOR U8691 ( .A(n10268), .B(n10269), .Z(n7435) );
  NOR U8692 ( .A(n10270), .B(n10268), .Z(n10269) );
  XOR U8693 ( .A(n10271), .B(n10272), .Z(n7438) );
  NOR U8694 ( .A(n10273), .B(n10271), .Z(n10272) );
  XOR U8695 ( .A(n10274), .B(n10275), .Z(n7441) );
  NOR U8696 ( .A(n10276), .B(n10274), .Z(n10275) );
  XOR U8697 ( .A(n10277), .B(n10278), .Z(n7444) );
  NOR U8698 ( .A(n10279), .B(n10277), .Z(n10278) );
  XOR U8699 ( .A(n10280), .B(n10281), .Z(n7447) );
  NOR U8700 ( .A(n10282), .B(n10280), .Z(n10281) );
  XOR U8701 ( .A(n10283), .B(n10284), .Z(n7450) );
  NOR U8702 ( .A(n10285), .B(n10283), .Z(n10284) );
  XOR U8703 ( .A(n10286), .B(n10287), .Z(n7453) );
  NOR U8704 ( .A(n10288), .B(n10286), .Z(n10287) );
  XOR U8705 ( .A(n10289), .B(n10290), .Z(n7456) );
  NOR U8706 ( .A(n10291), .B(n10289), .Z(n10290) );
  XOR U8707 ( .A(n10292), .B(n10293), .Z(n7459) );
  NOR U8708 ( .A(n10294), .B(n10292), .Z(n10293) );
  XOR U8709 ( .A(n10295), .B(n10296), .Z(n7462) );
  NOR U8710 ( .A(n10297), .B(n10295), .Z(n10296) );
  XOR U8711 ( .A(n10298), .B(n10299), .Z(n7465) );
  NOR U8712 ( .A(n10300), .B(n10298), .Z(n10299) );
  XOR U8713 ( .A(n10301), .B(n10302), .Z(n7468) );
  NOR U8714 ( .A(n10303), .B(n10301), .Z(n10302) );
  XOR U8715 ( .A(n10304), .B(n10305), .Z(n7471) );
  NOR U8716 ( .A(n10306), .B(n10304), .Z(n10305) );
  XOR U8717 ( .A(n10307), .B(n10308), .Z(n7474) );
  NOR U8718 ( .A(n10309), .B(n10307), .Z(n10308) );
  XOR U8719 ( .A(n10310), .B(n10311), .Z(n7477) );
  NOR U8720 ( .A(n10312), .B(n10310), .Z(n10311) );
  XOR U8721 ( .A(n10313), .B(n10314), .Z(n7480) );
  NOR U8722 ( .A(n10315), .B(n10313), .Z(n10314) );
  XOR U8723 ( .A(n10316), .B(n10317), .Z(n7483) );
  NOR U8724 ( .A(n10318), .B(n10316), .Z(n10317) );
  XOR U8725 ( .A(n10319), .B(n10320), .Z(n7486) );
  NOR U8726 ( .A(n10321), .B(n10319), .Z(n10320) );
  XOR U8727 ( .A(n10322), .B(n10323), .Z(n7489) );
  NOR U8728 ( .A(n10324), .B(n10322), .Z(n10323) );
  XOR U8729 ( .A(n10325), .B(n10326), .Z(n7492) );
  NOR U8730 ( .A(n10327), .B(n10325), .Z(n10326) );
  XOR U8731 ( .A(n10328), .B(n10329), .Z(n7495) );
  NOR U8732 ( .A(n10330), .B(n10328), .Z(n10329) );
  XOR U8733 ( .A(n10331), .B(n10332), .Z(n7498) );
  NOR U8734 ( .A(n10333), .B(n10331), .Z(n10332) );
  XOR U8735 ( .A(n10334), .B(n10335), .Z(n7501) );
  NOR U8736 ( .A(n10336), .B(n10334), .Z(n10335) );
  XOR U8737 ( .A(n10337), .B(n10338), .Z(n7504) );
  NOR U8738 ( .A(n10339), .B(n10337), .Z(n10338) );
  XOR U8739 ( .A(n10340), .B(n10341), .Z(n7507) );
  NOR U8740 ( .A(n10342), .B(n10340), .Z(n10341) );
  XOR U8741 ( .A(n10343), .B(n10344), .Z(n7510) );
  NOR U8742 ( .A(n10345), .B(n10343), .Z(n10344) );
  XOR U8743 ( .A(n10346), .B(n10347), .Z(n7513) );
  NOR U8744 ( .A(n10348), .B(n10346), .Z(n10347) );
  XOR U8745 ( .A(n10349), .B(n10350), .Z(n7516) );
  NOR U8746 ( .A(n10351), .B(n10349), .Z(n10350) );
  XOR U8747 ( .A(n10352), .B(n10353), .Z(n7519) );
  NOR U8748 ( .A(n10354), .B(n10352), .Z(n10353) );
  XOR U8749 ( .A(n10355), .B(n10356), .Z(n7522) );
  NOR U8750 ( .A(n10357), .B(n10355), .Z(n10356) );
  XOR U8751 ( .A(n10358), .B(n10359), .Z(n7525) );
  NOR U8752 ( .A(n10360), .B(n10358), .Z(n10359) );
  XOR U8753 ( .A(n10361), .B(n10362), .Z(n7528) );
  NOR U8754 ( .A(n10363), .B(n10361), .Z(n10362) );
  XOR U8755 ( .A(n10364), .B(n10365), .Z(n7531) );
  NOR U8756 ( .A(n10366), .B(n10364), .Z(n10365) );
  XOR U8757 ( .A(n10367), .B(n10368), .Z(n7534) );
  NOR U8758 ( .A(n10369), .B(n10367), .Z(n10368) );
  XOR U8759 ( .A(n10370), .B(n10371), .Z(n7537) );
  NOR U8760 ( .A(n10372), .B(n10370), .Z(n10371) );
  XOR U8761 ( .A(n10373), .B(n10374), .Z(n7540) );
  NOR U8762 ( .A(n10375), .B(n10373), .Z(n10374) );
  XOR U8763 ( .A(n10376), .B(n10377), .Z(n7543) );
  NOR U8764 ( .A(n10378), .B(n10376), .Z(n10377) );
  XOR U8765 ( .A(n10379), .B(n10380), .Z(n7546) );
  NOR U8766 ( .A(n10381), .B(n10379), .Z(n10380) );
  XOR U8767 ( .A(n10382), .B(n10383), .Z(n7549) );
  NOR U8768 ( .A(n10384), .B(n10382), .Z(n10383) );
  XOR U8769 ( .A(n10385), .B(n10386), .Z(n7552) );
  NOR U8770 ( .A(n10387), .B(n10385), .Z(n10386) );
  XOR U8771 ( .A(n10388), .B(n10389), .Z(n7555) );
  NOR U8772 ( .A(n10390), .B(n10388), .Z(n10389) );
  XOR U8773 ( .A(n10391), .B(n10392), .Z(n7558) );
  NOR U8774 ( .A(n10393), .B(n10391), .Z(n10392) );
  XOR U8775 ( .A(n10394), .B(n10395), .Z(n7561) );
  NOR U8776 ( .A(n10396), .B(n10394), .Z(n10395) );
  XOR U8777 ( .A(n10397), .B(n10398), .Z(n7564) );
  NOR U8778 ( .A(n10399), .B(n10397), .Z(n10398) );
  XOR U8779 ( .A(n10400), .B(n10401), .Z(n7567) );
  NOR U8780 ( .A(n10402), .B(n10400), .Z(n10401) );
  XOR U8781 ( .A(n10403), .B(n10404), .Z(n7570) );
  NOR U8782 ( .A(n10405), .B(n10403), .Z(n10404) );
  XOR U8783 ( .A(n10406), .B(n10407), .Z(n7573) );
  NOR U8784 ( .A(n10408), .B(n10406), .Z(n10407) );
  XOR U8785 ( .A(n10409), .B(n10410), .Z(n7576) );
  NOR U8786 ( .A(n10411), .B(n10409), .Z(n10410) );
  XOR U8787 ( .A(n10412), .B(n10413), .Z(n7579) );
  NOR U8788 ( .A(n10414), .B(n10412), .Z(n10413) );
  XOR U8789 ( .A(n10415), .B(n10416), .Z(n7582) );
  NOR U8790 ( .A(n10417), .B(n10415), .Z(n10416) );
  XOR U8791 ( .A(n10418), .B(n10419), .Z(n7585) );
  NOR U8792 ( .A(n10420), .B(n10418), .Z(n10419) );
  XOR U8793 ( .A(n10421), .B(n10422), .Z(n7588) );
  NOR U8794 ( .A(n10423), .B(n10421), .Z(n10422) );
  XOR U8795 ( .A(n10424), .B(n10425), .Z(n7591) );
  NOR U8796 ( .A(n10426), .B(n10424), .Z(n10425) );
  XOR U8797 ( .A(n10427), .B(n10428), .Z(n7594) );
  NOR U8798 ( .A(n10429), .B(n10427), .Z(n10428) );
  XOR U8799 ( .A(n10430), .B(n10431), .Z(n7597) );
  NOR U8800 ( .A(n10432), .B(n10430), .Z(n10431) );
  XOR U8801 ( .A(n10433), .B(n10434), .Z(n7600) );
  NOR U8802 ( .A(n10435), .B(n10433), .Z(n10434) );
  XOR U8803 ( .A(n10436), .B(n10437), .Z(n7603) );
  NOR U8804 ( .A(n10438), .B(n10436), .Z(n10437) );
  XOR U8805 ( .A(n10439), .B(n10440), .Z(n7606) );
  NOR U8806 ( .A(n10441), .B(n10439), .Z(n10440) );
  XOR U8807 ( .A(n10442), .B(n10443), .Z(n7609) );
  NOR U8808 ( .A(n10444), .B(n10442), .Z(n10443) );
  XOR U8809 ( .A(n10445), .B(n10446), .Z(n7612) );
  NOR U8810 ( .A(n10447), .B(n10445), .Z(n10446) );
  XOR U8811 ( .A(n10448), .B(n10449), .Z(n7615) );
  NOR U8812 ( .A(n10450), .B(n10448), .Z(n10449) );
  XOR U8813 ( .A(n10451), .B(n10452), .Z(n7618) );
  NOR U8814 ( .A(n10453), .B(n10451), .Z(n10452) );
  XOR U8815 ( .A(n10454), .B(n10455), .Z(n7621) );
  NOR U8816 ( .A(n10456), .B(n10454), .Z(n10455) );
  XOR U8817 ( .A(n10457), .B(n10458), .Z(n7624) );
  NOR U8818 ( .A(n10459), .B(n10457), .Z(n10458) );
  XOR U8819 ( .A(n10460), .B(n10461), .Z(n7627) );
  NOR U8820 ( .A(n10462), .B(n10460), .Z(n10461) );
  XOR U8821 ( .A(n10463), .B(n10464), .Z(n7630) );
  NOR U8822 ( .A(n10465), .B(n10463), .Z(n10464) );
  XOR U8823 ( .A(n10466), .B(n10467), .Z(n7633) );
  NOR U8824 ( .A(n10468), .B(n10466), .Z(n10467) );
  XOR U8825 ( .A(n10469), .B(n10470), .Z(n7636) );
  NOR U8826 ( .A(n10471), .B(n10469), .Z(n10470) );
  XOR U8827 ( .A(n10472), .B(n10473), .Z(n7639) );
  NOR U8828 ( .A(n10474), .B(n10472), .Z(n10473) );
  XOR U8829 ( .A(n10475), .B(n10476), .Z(n7642) );
  NOR U8830 ( .A(n10477), .B(n10475), .Z(n10476) );
  XOR U8831 ( .A(n10478), .B(n10479), .Z(n7645) );
  NOR U8832 ( .A(n10480), .B(n10478), .Z(n10479) );
  XOR U8833 ( .A(n10481), .B(n10482), .Z(n7648) );
  NOR U8834 ( .A(n10483), .B(n10481), .Z(n10482) );
  XOR U8835 ( .A(n10484), .B(n10485), .Z(n7651) );
  NOR U8836 ( .A(n10486), .B(n10484), .Z(n10485) );
  XOR U8837 ( .A(n10487), .B(n10488), .Z(n7654) );
  NOR U8838 ( .A(n10489), .B(n10487), .Z(n10488) );
  XOR U8839 ( .A(n10490), .B(n10491), .Z(n7657) );
  NOR U8840 ( .A(n10492), .B(n10490), .Z(n10491) );
  XOR U8841 ( .A(n10493), .B(n10494), .Z(n7660) );
  NOR U8842 ( .A(n10495), .B(n10493), .Z(n10494) );
  XOR U8843 ( .A(n10496), .B(n10497), .Z(n7663) );
  NOR U8844 ( .A(n10498), .B(n10496), .Z(n10497) );
  XOR U8845 ( .A(n10499), .B(n10500), .Z(n7666) );
  NOR U8846 ( .A(n10501), .B(n10499), .Z(n10500) );
  XOR U8847 ( .A(n10502), .B(n10503), .Z(n7669) );
  NOR U8848 ( .A(n10504), .B(n10502), .Z(n10503) );
  XOR U8849 ( .A(n10505), .B(n10506), .Z(n7672) );
  NOR U8850 ( .A(n10507), .B(n10505), .Z(n10506) );
  XOR U8851 ( .A(n10508), .B(n10509), .Z(n7675) );
  NOR U8852 ( .A(n10510), .B(n10508), .Z(n10509) );
  XOR U8853 ( .A(n10511), .B(n10512), .Z(n7678) );
  NOR U8854 ( .A(n10513), .B(n10511), .Z(n10512) );
  XOR U8855 ( .A(n10514), .B(n10515), .Z(n7681) );
  NOR U8856 ( .A(n10516), .B(n10514), .Z(n10515) );
  XOR U8857 ( .A(n10517), .B(n10518), .Z(n7684) );
  NOR U8858 ( .A(n10519), .B(n10517), .Z(n10518) );
  XOR U8859 ( .A(n10520), .B(n10521), .Z(n7687) );
  NOR U8860 ( .A(n10522), .B(n10520), .Z(n10521) );
  XOR U8861 ( .A(n10523), .B(n10524), .Z(n7690) );
  NOR U8862 ( .A(n10525), .B(n10523), .Z(n10524) );
  XOR U8863 ( .A(n10526), .B(n10527), .Z(n7693) );
  NOR U8864 ( .A(n10528), .B(n10526), .Z(n10527) );
  XOR U8865 ( .A(n10529), .B(n10530), .Z(n7696) );
  NOR U8866 ( .A(n10531), .B(n10529), .Z(n10530) );
  XOR U8867 ( .A(n10532), .B(n10533), .Z(n7699) );
  NOR U8868 ( .A(n10534), .B(n10532), .Z(n10533) );
  XOR U8869 ( .A(n10535), .B(n10536), .Z(n7702) );
  NOR U8870 ( .A(n10537), .B(n10535), .Z(n10536) );
  XOR U8871 ( .A(n10538), .B(n10539), .Z(n7705) );
  NOR U8872 ( .A(n10540), .B(n10538), .Z(n10539) );
  XOR U8873 ( .A(n10541), .B(n10542), .Z(n7708) );
  NOR U8874 ( .A(n10543), .B(n10541), .Z(n10542) );
  XOR U8875 ( .A(n10544), .B(n10545), .Z(n7711) );
  NOR U8876 ( .A(n10546), .B(n10544), .Z(n10545) );
  XOR U8877 ( .A(n10547), .B(n10548), .Z(n7714) );
  NOR U8878 ( .A(n10549), .B(n10547), .Z(n10548) );
  XOR U8879 ( .A(n10550), .B(n10551), .Z(n7717) );
  NOR U8880 ( .A(n10552), .B(n10550), .Z(n10551) );
  XOR U8881 ( .A(n10553), .B(n10554), .Z(n7720) );
  NOR U8882 ( .A(n10555), .B(n10553), .Z(n10554) );
  XOR U8883 ( .A(n10556), .B(n10557), .Z(n7723) );
  NOR U8884 ( .A(n10558), .B(n10556), .Z(n10557) );
  XOR U8885 ( .A(n10559), .B(n10560), .Z(n7726) );
  NOR U8886 ( .A(n10561), .B(n10559), .Z(n10560) );
  XOR U8887 ( .A(n10562), .B(n10563), .Z(n7729) );
  NOR U8888 ( .A(n10564), .B(n10562), .Z(n10563) );
  XOR U8889 ( .A(n10565), .B(n10566), .Z(n7732) );
  NOR U8890 ( .A(n10567), .B(n10565), .Z(n10566) );
  XOR U8891 ( .A(n10568), .B(n10569), .Z(n7735) );
  NOR U8892 ( .A(n10570), .B(n10568), .Z(n10569) );
  XOR U8893 ( .A(n10571), .B(n10572), .Z(n7738) );
  NOR U8894 ( .A(n10573), .B(n10571), .Z(n10572) );
  XOR U8895 ( .A(n10574), .B(n10575), .Z(n7741) );
  NOR U8896 ( .A(n10576), .B(n10574), .Z(n10575) );
  XOR U8897 ( .A(n10577), .B(n10578), .Z(n7744) );
  NOR U8898 ( .A(n10579), .B(n10577), .Z(n10578) );
  XOR U8899 ( .A(n10580), .B(n10581), .Z(n7747) );
  NOR U8900 ( .A(n10582), .B(n10580), .Z(n10581) );
  XOR U8901 ( .A(n10583), .B(n10584), .Z(n7750) );
  NOR U8902 ( .A(n10585), .B(n10583), .Z(n10584) );
  XOR U8903 ( .A(n10586), .B(n10587), .Z(n7753) );
  NOR U8904 ( .A(n10588), .B(n10586), .Z(n10587) );
  XOR U8905 ( .A(n10589), .B(n10590), .Z(n7756) );
  NOR U8906 ( .A(n10591), .B(n10589), .Z(n10590) );
  XOR U8907 ( .A(n10592), .B(n10593), .Z(n7759) );
  NOR U8908 ( .A(n10594), .B(n10592), .Z(n10593) );
  XOR U8909 ( .A(n10595), .B(n10596), .Z(n7762) );
  NOR U8910 ( .A(n10597), .B(n10595), .Z(n10596) );
  XOR U8911 ( .A(n10598), .B(n10599), .Z(n7765) );
  NOR U8912 ( .A(n10600), .B(n10598), .Z(n10599) );
  XOR U8913 ( .A(n10601), .B(n10602), .Z(n7768) );
  NOR U8914 ( .A(n10603), .B(n10601), .Z(n10602) );
  XOR U8915 ( .A(n10604), .B(n10605), .Z(n7771) );
  NOR U8916 ( .A(n10606), .B(n10604), .Z(n10605) );
  XOR U8917 ( .A(n10607), .B(n10608), .Z(n7774) );
  NOR U8918 ( .A(n10609), .B(n10607), .Z(n10608) );
  XOR U8919 ( .A(n10610), .B(n10611), .Z(n7777) );
  NOR U8920 ( .A(n10612), .B(n10610), .Z(n10611) );
  XOR U8921 ( .A(n10613), .B(n10614), .Z(n7780) );
  NOR U8922 ( .A(n10615), .B(n10613), .Z(n10614) );
  XOR U8923 ( .A(n10616), .B(n10617), .Z(n7783) );
  NOR U8924 ( .A(n10618), .B(n10616), .Z(n10617) );
  XOR U8925 ( .A(n10619), .B(n10620), .Z(n7786) );
  NOR U8926 ( .A(n10621), .B(n10619), .Z(n10620) );
  XOR U8927 ( .A(n10622), .B(n10623), .Z(n7789) );
  NOR U8928 ( .A(n10624), .B(n10622), .Z(n10623) );
  XOR U8929 ( .A(n10625), .B(n10626), .Z(n7792) );
  NOR U8930 ( .A(n10627), .B(n10625), .Z(n10626) );
  XOR U8931 ( .A(n10628), .B(n10629), .Z(n7795) );
  NOR U8932 ( .A(n10630), .B(n10628), .Z(n10629) );
  XOR U8933 ( .A(n10631), .B(n10632), .Z(n7798) );
  NOR U8934 ( .A(n10633), .B(n10631), .Z(n10632) );
  XOR U8935 ( .A(n10634), .B(n10635), .Z(n7801) );
  NOR U8936 ( .A(n10636), .B(n10634), .Z(n10635) );
  XOR U8937 ( .A(n10637), .B(n10638), .Z(n7804) );
  NOR U8938 ( .A(n10639), .B(n10637), .Z(n10638) );
  XOR U8939 ( .A(n10640), .B(n10641), .Z(n7807) );
  NOR U8940 ( .A(n10642), .B(n10640), .Z(n10641) );
  XOR U8941 ( .A(n10643), .B(n10644), .Z(n7810) );
  NOR U8942 ( .A(n10645), .B(n10643), .Z(n10644) );
  XOR U8943 ( .A(n10646), .B(n10647), .Z(n7813) );
  NOR U8944 ( .A(n10648), .B(n10646), .Z(n10647) );
  XOR U8945 ( .A(n10649), .B(n10650), .Z(n7816) );
  NOR U8946 ( .A(n10651), .B(n10649), .Z(n10650) );
  XOR U8947 ( .A(n10652), .B(n10653), .Z(n7819) );
  NOR U8948 ( .A(n10654), .B(n10652), .Z(n10653) );
  XOR U8949 ( .A(n10655), .B(n10656), .Z(n7822) );
  NOR U8950 ( .A(n10657), .B(n10655), .Z(n10656) );
  XOR U8951 ( .A(n10658), .B(n10659), .Z(n7825) );
  NOR U8952 ( .A(n10660), .B(n10658), .Z(n10659) );
  XOR U8953 ( .A(n10661), .B(n10662), .Z(n7828) );
  NOR U8954 ( .A(n10663), .B(n10661), .Z(n10662) );
  XOR U8955 ( .A(n10664), .B(n10665), .Z(n7831) );
  NOR U8956 ( .A(n10666), .B(n10664), .Z(n10665) );
  XOR U8957 ( .A(n10667), .B(n10668), .Z(n7834) );
  NOR U8958 ( .A(n10669), .B(n10667), .Z(n10668) );
  XOR U8959 ( .A(n10670), .B(n10671), .Z(n7837) );
  NOR U8960 ( .A(n10672), .B(n10670), .Z(n10671) );
  XOR U8961 ( .A(n10673), .B(n10674), .Z(n7840) );
  NOR U8962 ( .A(n10675), .B(n10673), .Z(n10674) );
  XOR U8963 ( .A(n10676), .B(n10677), .Z(n7843) );
  NOR U8964 ( .A(n10678), .B(n10676), .Z(n10677) );
  XOR U8965 ( .A(n10679), .B(n10680), .Z(n7846) );
  NOR U8966 ( .A(n10681), .B(n10679), .Z(n10680) );
  XOR U8967 ( .A(n10682), .B(n10683), .Z(n7849) );
  NOR U8968 ( .A(n10684), .B(n10682), .Z(n10683) );
  XOR U8969 ( .A(n10685), .B(n10686), .Z(n7852) );
  NOR U8970 ( .A(n10687), .B(n10685), .Z(n10686) );
  XOR U8971 ( .A(n10688), .B(n10689), .Z(n7855) );
  NOR U8972 ( .A(n10690), .B(n10688), .Z(n10689) );
  XOR U8973 ( .A(n10691), .B(n10692), .Z(n7858) );
  NOR U8974 ( .A(n10693), .B(n10691), .Z(n10692) );
  XOR U8975 ( .A(n10694), .B(n10695), .Z(n7861) );
  NOR U8976 ( .A(n10696), .B(n10694), .Z(n10695) );
  XOR U8977 ( .A(n10697), .B(n10698), .Z(n7864) );
  NOR U8978 ( .A(n10699), .B(n10697), .Z(n10698) );
  XOR U8979 ( .A(n10700), .B(n10701), .Z(n7867) );
  NOR U8980 ( .A(n10702), .B(n10700), .Z(n10701) );
  XOR U8981 ( .A(n10703), .B(n10704), .Z(n7870) );
  NOR U8982 ( .A(n10705), .B(n10703), .Z(n10704) );
  XOR U8983 ( .A(n10706), .B(n10707), .Z(n7873) );
  NOR U8984 ( .A(n10708), .B(n10706), .Z(n10707) );
  XOR U8985 ( .A(n10709), .B(n10710), .Z(n7876) );
  NOR U8986 ( .A(n10711), .B(n10709), .Z(n10710) );
  XOR U8987 ( .A(n10712), .B(n10713), .Z(n7879) );
  NOR U8988 ( .A(n10714), .B(n10712), .Z(n10713) );
  XOR U8989 ( .A(n10715), .B(n10716), .Z(n7882) );
  NOR U8990 ( .A(n10717), .B(n10715), .Z(n10716) );
  XOR U8991 ( .A(n10718), .B(n10719), .Z(n7885) );
  NOR U8992 ( .A(n10720), .B(n10718), .Z(n10719) );
  XOR U8993 ( .A(n10721), .B(n10722), .Z(n7888) );
  NOR U8994 ( .A(n10723), .B(n10721), .Z(n10722) );
  XOR U8995 ( .A(n10724), .B(n10725), .Z(n7891) );
  NOR U8996 ( .A(n10726), .B(n10724), .Z(n10725) );
  XOR U8997 ( .A(n10727), .B(n10728), .Z(n7894) );
  NOR U8998 ( .A(n10729), .B(n10727), .Z(n10728) );
  XOR U8999 ( .A(n10730), .B(n10731), .Z(n7897) );
  NOR U9000 ( .A(n10732), .B(n10730), .Z(n10731) );
  XOR U9001 ( .A(n10733), .B(n10734), .Z(n7900) );
  NOR U9002 ( .A(n10735), .B(n10733), .Z(n10734) );
  XOR U9003 ( .A(n10736), .B(n10737), .Z(n7903) );
  NOR U9004 ( .A(n10738), .B(n10736), .Z(n10737) );
  XOR U9005 ( .A(n10739), .B(n10740), .Z(n7906) );
  NOR U9006 ( .A(n10741), .B(n10739), .Z(n10740) );
  XOR U9007 ( .A(n10742), .B(n10743), .Z(n7909) );
  NOR U9008 ( .A(n10744), .B(n10742), .Z(n10743) );
  XOR U9009 ( .A(n10745), .B(n10746), .Z(n7912) );
  NOR U9010 ( .A(n10747), .B(n10745), .Z(n10746) );
  XOR U9011 ( .A(n10748), .B(n10749), .Z(n7915) );
  NOR U9012 ( .A(n10750), .B(n10748), .Z(n10749) );
  XOR U9013 ( .A(n10751), .B(n10752), .Z(n7918) );
  NOR U9014 ( .A(n10753), .B(n10751), .Z(n10752) );
  XOR U9015 ( .A(n10754), .B(n10755), .Z(n7921) );
  NOR U9016 ( .A(n10756), .B(n10754), .Z(n10755) );
  XOR U9017 ( .A(n10757), .B(n10758), .Z(n7924) );
  NOR U9018 ( .A(n10759), .B(n10757), .Z(n10758) );
  XOR U9019 ( .A(n10760), .B(n10761), .Z(n7927) );
  NOR U9020 ( .A(n10762), .B(n10760), .Z(n10761) );
  XOR U9021 ( .A(n10763), .B(n10764), .Z(n7930) );
  NOR U9022 ( .A(n10765), .B(n10763), .Z(n10764) );
  XOR U9023 ( .A(n10766), .B(n10767), .Z(n7933) );
  NOR U9024 ( .A(n10768), .B(n10766), .Z(n10767) );
  XOR U9025 ( .A(n10769), .B(n10770), .Z(n7936) );
  NOR U9026 ( .A(n10771), .B(n10769), .Z(n10770) );
  XOR U9027 ( .A(n10772), .B(n10773), .Z(n7939) );
  NOR U9028 ( .A(n10774), .B(n10772), .Z(n10773) );
  XOR U9029 ( .A(n10775), .B(n10776), .Z(n7942) );
  NOR U9030 ( .A(n10777), .B(n10775), .Z(n10776) );
  XOR U9031 ( .A(n10778), .B(n10779), .Z(n7945) );
  NOR U9032 ( .A(n10780), .B(n10778), .Z(n10779) );
  XOR U9033 ( .A(n10781), .B(n10782), .Z(n7948) );
  NOR U9034 ( .A(n10783), .B(n10781), .Z(n10782) );
  XOR U9035 ( .A(n10784), .B(n10785), .Z(n7951) );
  NOR U9036 ( .A(n10786), .B(n10784), .Z(n10785) );
  XOR U9037 ( .A(n10787), .B(n10788), .Z(n7954) );
  NOR U9038 ( .A(n10789), .B(n10787), .Z(n10788) );
  XOR U9039 ( .A(n10790), .B(n10791), .Z(n7957) );
  NOR U9040 ( .A(n10792), .B(n10790), .Z(n10791) );
  XOR U9041 ( .A(n10793), .B(n10794), .Z(n7960) );
  NOR U9042 ( .A(n10795), .B(n10793), .Z(n10794) );
  XOR U9043 ( .A(n10796), .B(n10797), .Z(n7963) );
  NOR U9044 ( .A(n10798), .B(n10796), .Z(n10797) );
  XOR U9045 ( .A(n10799), .B(n10800), .Z(n7966) );
  NOR U9046 ( .A(n10801), .B(n10799), .Z(n10800) );
  XOR U9047 ( .A(n10802), .B(n10803), .Z(n7969) );
  NOR U9048 ( .A(n10804), .B(n10802), .Z(n10803) );
  XOR U9049 ( .A(n10805), .B(n10806), .Z(n7972) );
  NOR U9050 ( .A(n10807), .B(n10805), .Z(n10806) );
  XOR U9051 ( .A(n10808), .B(n10809), .Z(n7975) );
  NOR U9052 ( .A(n10810), .B(n10808), .Z(n10809) );
  XOR U9053 ( .A(n10811), .B(n10812), .Z(n7978) );
  NOR U9054 ( .A(n10813), .B(n10811), .Z(n10812) );
  XOR U9055 ( .A(n10814), .B(n10815), .Z(n7981) );
  NOR U9056 ( .A(n10816), .B(n10814), .Z(n10815) );
  XOR U9057 ( .A(n10817), .B(n10818), .Z(n7984) );
  NOR U9058 ( .A(n10819), .B(n10817), .Z(n10818) );
  XOR U9059 ( .A(n10820), .B(n10821), .Z(n7987) );
  NOR U9060 ( .A(n10822), .B(n10820), .Z(n10821) );
  XOR U9061 ( .A(n10823), .B(n10824), .Z(n7990) );
  NOR U9062 ( .A(n10825), .B(n10823), .Z(n10824) );
  XOR U9063 ( .A(n10826), .B(n10827), .Z(n7993) );
  NOR U9064 ( .A(n10828), .B(n10826), .Z(n10827) );
  XOR U9065 ( .A(n10829), .B(n10830), .Z(n7996) );
  NOR U9066 ( .A(n10831), .B(n10829), .Z(n10830) );
  XOR U9067 ( .A(n10832), .B(n10833), .Z(n7999) );
  NOR U9068 ( .A(n10834), .B(n10832), .Z(n10833) );
  XOR U9069 ( .A(n10835), .B(n10836), .Z(n8002) );
  NOR U9070 ( .A(n10837), .B(n10835), .Z(n10836) );
  XOR U9071 ( .A(n10838), .B(n10839), .Z(n8005) );
  NOR U9072 ( .A(n10840), .B(n10838), .Z(n10839) );
  XOR U9073 ( .A(n10841), .B(n10842), .Z(n8008) );
  NOR U9074 ( .A(n10843), .B(n10841), .Z(n10842) );
  XOR U9075 ( .A(n10844), .B(n10845), .Z(n8011) );
  NOR U9076 ( .A(n10846), .B(n10844), .Z(n10845) );
  XOR U9077 ( .A(n10847), .B(n10848), .Z(n8014) );
  NOR U9078 ( .A(n10849), .B(n10847), .Z(n10848) );
  XOR U9079 ( .A(n10850), .B(n10851), .Z(n8017) );
  NOR U9080 ( .A(n10852), .B(n10850), .Z(n10851) );
  XOR U9081 ( .A(n10853), .B(n10854), .Z(n8020) );
  NOR U9082 ( .A(n10855), .B(n10853), .Z(n10854) );
  XOR U9083 ( .A(n10856), .B(n10857), .Z(n8023) );
  NOR U9084 ( .A(n10858), .B(n10856), .Z(n10857) );
  XOR U9085 ( .A(n10859), .B(n10860), .Z(n8026) );
  NOR U9086 ( .A(n10861), .B(n10859), .Z(n10860) );
  XOR U9087 ( .A(n10862), .B(n10863), .Z(n8029) );
  NOR U9088 ( .A(n10864), .B(n10862), .Z(n10863) );
  XOR U9089 ( .A(n10865), .B(n10866), .Z(n8032) );
  NOR U9090 ( .A(n10867), .B(n10865), .Z(n10866) );
  XOR U9091 ( .A(n10868), .B(n10869), .Z(n8035) );
  NOR U9092 ( .A(n10870), .B(n10868), .Z(n10869) );
  XOR U9093 ( .A(n10871), .B(n10872), .Z(n8038) );
  NOR U9094 ( .A(n10873), .B(n10871), .Z(n10872) );
  XOR U9095 ( .A(n10874), .B(n10875), .Z(n8041) );
  NOR U9096 ( .A(n10876), .B(n10874), .Z(n10875) );
  XOR U9097 ( .A(n10877), .B(n10878), .Z(n8044) );
  NOR U9098 ( .A(n10879), .B(n10877), .Z(n10878) );
  XOR U9099 ( .A(n10880), .B(n10881), .Z(n8047) );
  NOR U9100 ( .A(n10882), .B(n10880), .Z(n10881) );
  XOR U9101 ( .A(n10883), .B(n10884), .Z(n8050) );
  NOR U9102 ( .A(n10885), .B(n10883), .Z(n10884) );
  XOR U9103 ( .A(n10886), .B(n10887), .Z(n8053) );
  NOR U9104 ( .A(n10888), .B(n10886), .Z(n10887) );
  XOR U9105 ( .A(n10889), .B(n10890), .Z(n8056) );
  NOR U9106 ( .A(n10891), .B(n10889), .Z(n10890) );
  XOR U9107 ( .A(n10892), .B(n10893), .Z(n8059) );
  NOR U9108 ( .A(n10894), .B(n10892), .Z(n10893) );
  XOR U9109 ( .A(n10895), .B(n10896), .Z(n8062) );
  NOR U9110 ( .A(n10897), .B(n10895), .Z(n10896) );
  XOR U9111 ( .A(n10898), .B(n10899), .Z(n8065) );
  NOR U9112 ( .A(n10900), .B(n10898), .Z(n10899) );
  XOR U9113 ( .A(n10901), .B(n10902), .Z(n8068) );
  NOR U9114 ( .A(n10903), .B(n10901), .Z(n10902) );
  XOR U9115 ( .A(n10904), .B(n10905), .Z(n8071) );
  NOR U9116 ( .A(n10906), .B(n10904), .Z(n10905) );
  XOR U9117 ( .A(n10907), .B(n10908), .Z(n8074) );
  NOR U9118 ( .A(n10909), .B(n10907), .Z(n10908) );
  XOR U9119 ( .A(n10910), .B(n10911), .Z(n8077) );
  NOR U9120 ( .A(n10912), .B(n10910), .Z(n10911) );
  XOR U9121 ( .A(n10913), .B(n10914), .Z(n8080) );
  NOR U9122 ( .A(n10915), .B(n10913), .Z(n10914) );
  XOR U9123 ( .A(n10916), .B(n10917), .Z(n8083) );
  NOR U9124 ( .A(n10918), .B(n10916), .Z(n10917) );
  XOR U9125 ( .A(n10919), .B(n10920), .Z(n8086) );
  NOR U9126 ( .A(n10921), .B(n10919), .Z(n10920) );
  XOR U9127 ( .A(n10922), .B(n10923), .Z(n8089) );
  NOR U9128 ( .A(n10924), .B(n10922), .Z(n10923) );
  XOR U9129 ( .A(n10925), .B(n10926), .Z(n8092) );
  NOR U9130 ( .A(n10927), .B(n10925), .Z(n10926) );
  XOR U9131 ( .A(n10928), .B(n10929), .Z(n8095) );
  NOR U9132 ( .A(n10930), .B(n10928), .Z(n10929) );
  XOR U9133 ( .A(n10931), .B(n10932), .Z(n8098) );
  NOR U9134 ( .A(n10933), .B(n10931), .Z(n10932) );
  XOR U9135 ( .A(n10934), .B(n10935), .Z(n8101) );
  NOR U9136 ( .A(n10936), .B(n10934), .Z(n10935) );
  XOR U9137 ( .A(n10937), .B(n10938), .Z(n8104) );
  NOR U9138 ( .A(n10939), .B(n10937), .Z(n10938) );
  XOR U9139 ( .A(n10940), .B(n10941), .Z(n8107) );
  NOR U9140 ( .A(n10942), .B(n10940), .Z(n10941) );
  XOR U9141 ( .A(n10943), .B(n10944), .Z(n8110) );
  NOR U9142 ( .A(n10945), .B(n10943), .Z(n10944) );
  XOR U9143 ( .A(n10946), .B(n10947), .Z(n8113) );
  NOR U9144 ( .A(n10948), .B(n10946), .Z(n10947) );
  XOR U9145 ( .A(n10949), .B(n10950), .Z(n8116) );
  NOR U9146 ( .A(n10951), .B(n10949), .Z(n10950) );
  XOR U9147 ( .A(n10952), .B(n10953), .Z(n8119) );
  NOR U9148 ( .A(n10954), .B(n10952), .Z(n10953) );
  XOR U9149 ( .A(n10955), .B(n10956), .Z(n8122) );
  NOR U9150 ( .A(n10957), .B(n10955), .Z(n10956) );
  XOR U9151 ( .A(n10958), .B(n10959), .Z(n8125) );
  NOR U9152 ( .A(n10960), .B(n10958), .Z(n10959) );
  XOR U9153 ( .A(n10961), .B(n10962), .Z(n8128) );
  NOR U9154 ( .A(n10963), .B(n10961), .Z(n10962) );
  XOR U9155 ( .A(n10964), .B(n10965), .Z(n8131) );
  NOR U9156 ( .A(n10966), .B(n10964), .Z(n10965) );
  XOR U9157 ( .A(n10967), .B(n10968), .Z(n8134) );
  NOR U9158 ( .A(n10969), .B(n10967), .Z(n10968) );
  XOR U9159 ( .A(n10970), .B(n10971), .Z(n8137) );
  NOR U9160 ( .A(n10972), .B(n10970), .Z(n10971) );
  XOR U9161 ( .A(n10973), .B(n10974), .Z(n8140) );
  NOR U9162 ( .A(n10975), .B(n10973), .Z(n10974) );
  XOR U9163 ( .A(n10976), .B(n10977), .Z(n8143) );
  NOR U9164 ( .A(n10978), .B(n10976), .Z(n10977) );
  XOR U9165 ( .A(n10979), .B(n10980), .Z(n8146) );
  NOR U9166 ( .A(n10981), .B(n10979), .Z(n10980) );
  XOR U9167 ( .A(n10982), .B(n10983), .Z(n8149) );
  NOR U9168 ( .A(n10984), .B(n10982), .Z(n10983) );
  XOR U9169 ( .A(n10985), .B(n10986), .Z(n8152) );
  NOR U9170 ( .A(n10987), .B(n10985), .Z(n10986) );
  XOR U9171 ( .A(n10988), .B(n10989), .Z(n8155) );
  NOR U9172 ( .A(n10990), .B(n10988), .Z(n10989) );
  XOR U9173 ( .A(n10991), .B(n10992), .Z(n8158) );
  NOR U9174 ( .A(n10993), .B(n10991), .Z(n10992) );
  XOR U9175 ( .A(n10994), .B(n10995), .Z(n8161) );
  NOR U9176 ( .A(n10996), .B(n10994), .Z(n10995) );
  XOR U9177 ( .A(n10997), .B(n10998), .Z(n8164) );
  NOR U9178 ( .A(n10999), .B(n10997), .Z(n10998) );
  XOR U9179 ( .A(n11000), .B(n11001), .Z(n8167) );
  NOR U9180 ( .A(n11002), .B(n11000), .Z(n11001) );
  XOR U9181 ( .A(n11003), .B(n11004), .Z(n8170) );
  NOR U9182 ( .A(n11005), .B(n11003), .Z(n11004) );
  XOR U9183 ( .A(n11006), .B(n11007), .Z(n8173) );
  NOR U9184 ( .A(n11008), .B(n11006), .Z(n11007) );
  XOR U9185 ( .A(n11009), .B(n11010), .Z(n8176) );
  NOR U9186 ( .A(n11011), .B(n11009), .Z(n11010) );
  XOR U9187 ( .A(n11012), .B(n11013), .Z(n8179) );
  NOR U9188 ( .A(n11014), .B(n11012), .Z(n11013) );
  XOR U9189 ( .A(n11015), .B(n11016), .Z(n8182) );
  NOR U9190 ( .A(n11017), .B(n11015), .Z(n11016) );
  XOR U9191 ( .A(n11018), .B(n11019), .Z(n8185) );
  NOR U9192 ( .A(n11020), .B(n11018), .Z(n11019) );
  XOR U9193 ( .A(n11021), .B(n11022), .Z(n8188) );
  NOR U9194 ( .A(n11023), .B(n11021), .Z(n11022) );
  XOR U9195 ( .A(n11024), .B(n11025), .Z(n8191) );
  NOR U9196 ( .A(n11026), .B(n11024), .Z(n11025) );
  XOR U9197 ( .A(n11027), .B(n11028), .Z(n8194) );
  NOR U9198 ( .A(n11029), .B(n11027), .Z(n11028) );
  XOR U9199 ( .A(n11030), .B(n11031), .Z(n8197) );
  NOR U9200 ( .A(n11032), .B(n11030), .Z(n11031) );
  XOR U9201 ( .A(n11033), .B(n11034), .Z(n8200) );
  NOR U9202 ( .A(n11035), .B(n11033), .Z(n11034) );
  XOR U9203 ( .A(n11036), .B(n11037), .Z(n8203) );
  NOR U9204 ( .A(n11038), .B(n11036), .Z(n11037) );
  XOR U9205 ( .A(n11039), .B(n11040), .Z(n8206) );
  NOR U9206 ( .A(n11041), .B(n11039), .Z(n11040) );
  XOR U9207 ( .A(n11042), .B(n11043), .Z(n8209) );
  NOR U9208 ( .A(n11044), .B(n11042), .Z(n11043) );
  XOR U9209 ( .A(n11045), .B(n11046), .Z(n8212) );
  NOR U9210 ( .A(n11047), .B(n11045), .Z(n11046) );
  XOR U9211 ( .A(n11048), .B(n11049), .Z(n8215) );
  NOR U9212 ( .A(n11050), .B(n11048), .Z(n11049) );
  XOR U9213 ( .A(n11051), .B(n11052), .Z(n8218) );
  NOR U9214 ( .A(n11053), .B(n11051), .Z(n11052) );
  XOR U9215 ( .A(n11054), .B(n11055), .Z(n8221) );
  NOR U9216 ( .A(n11056), .B(n11054), .Z(n11055) );
  XOR U9217 ( .A(n11057), .B(n11058), .Z(n8224) );
  NOR U9218 ( .A(n11059), .B(n11057), .Z(n11058) );
  XOR U9219 ( .A(n11060), .B(n11061), .Z(n8227) );
  NOR U9220 ( .A(n11062), .B(n11060), .Z(n11061) );
  XOR U9221 ( .A(n11063), .B(n11064), .Z(n8230) );
  NOR U9222 ( .A(n11065), .B(n11063), .Z(n11064) );
  XOR U9223 ( .A(n11066), .B(n11067), .Z(n8233) );
  NOR U9224 ( .A(n11068), .B(n11066), .Z(n11067) );
  XOR U9225 ( .A(n11069), .B(n11070), .Z(n8236) );
  NOR U9226 ( .A(n11071), .B(n11069), .Z(n11070) );
  XOR U9227 ( .A(n11072), .B(n11073), .Z(n8239) );
  NOR U9228 ( .A(n11074), .B(n11072), .Z(n11073) );
  XOR U9229 ( .A(n11075), .B(n11076), .Z(n8242) );
  NOR U9230 ( .A(n11077), .B(n11075), .Z(n11076) );
  XOR U9231 ( .A(n11078), .B(n11079), .Z(n8245) );
  NOR U9232 ( .A(n11080), .B(n11078), .Z(n11079) );
  XOR U9233 ( .A(n11081), .B(n11082), .Z(n8248) );
  NOR U9234 ( .A(n11083), .B(n11081), .Z(n11082) );
  XOR U9235 ( .A(n11084), .B(n11085), .Z(n8251) );
  NOR U9236 ( .A(n11086), .B(n11084), .Z(n11085) );
  XOR U9237 ( .A(n11087), .B(n11088), .Z(n8254) );
  NOR U9238 ( .A(n11089), .B(n11087), .Z(n11088) );
  XOR U9239 ( .A(n11090), .B(n11091), .Z(n8257) );
  NOR U9240 ( .A(n11092), .B(n11090), .Z(n11091) );
  XOR U9241 ( .A(n11093), .B(n11094), .Z(n8260) );
  NOR U9242 ( .A(n11095), .B(n11093), .Z(n11094) );
  XOR U9243 ( .A(n11096), .B(n11097), .Z(n8263) );
  NOR U9244 ( .A(n11098), .B(n11096), .Z(n11097) );
  XOR U9245 ( .A(n11099), .B(n11100), .Z(n8266) );
  NOR U9246 ( .A(n11101), .B(n11099), .Z(n11100) );
  XOR U9247 ( .A(n11102), .B(n11103), .Z(n8269) );
  NOR U9248 ( .A(n11104), .B(n11102), .Z(n11103) );
  XOR U9249 ( .A(n11105), .B(n11106), .Z(n8272) );
  NOR U9250 ( .A(n11107), .B(n11105), .Z(n11106) );
  XOR U9251 ( .A(n11108), .B(n11109), .Z(n8275) );
  NOR U9252 ( .A(n11110), .B(n11108), .Z(n11109) );
  XOR U9253 ( .A(n11111), .B(n11112), .Z(n8278) );
  NOR U9254 ( .A(n11113), .B(n11111), .Z(n11112) );
  XOR U9255 ( .A(n11114), .B(n11115), .Z(n8281) );
  NOR U9256 ( .A(n11116), .B(n11114), .Z(n11115) );
  XOR U9257 ( .A(n11117), .B(n11118), .Z(n8284) );
  NOR U9258 ( .A(n11119), .B(n11117), .Z(n11118) );
  XOR U9259 ( .A(n11120), .B(n11121), .Z(n8287) );
  NOR U9260 ( .A(n11122), .B(n11120), .Z(n11121) );
  XOR U9261 ( .A(n11123), .B(n11124), .Z(n8290) );
  NOR U9262 ( .A(n11125), .B(n11123), .Z(n11124) );
  XOR U9263 ( .A(n11126), .B(n11127), .Z(n8293) );
  NOR U9264 ( .A(n11128), .B(n11126), .Z(n11127) );
  XOR U9265 ( .A(n11129), .B(n11130), .Z(n8296) );
  NOR U9266 ( .A(n11131), .B(n11129), .Z(n11130) );
  XOR U9267 ( .A(n11132), .B(n11133), .Z(n8299) );
  NOR U9268 ( .A(n11134), .B(n11132), .Z(n11133) );
  XOR U9269 ( .A(n11135), .B(n11136), .Z(n8302) );
  NOR U9270 ( .A(n11137), .B(n11135), .Z(n11136) );
  XOR U9271 ( .A(n11138), .B(n11139), .Z(n8305) );
  NOR U9272 ( .A(n11140), .B(n11138), .Z(n11139) );
  XOR U9273 ( .A(n11141), .B(n11142), .Z(n8308) );
  NOR U9274 ( .A(n11143), .B(n11141), .Z(n11142) );
  XOR U9275 ( .A(n11144), .B(n11145), .Z(n8311) );
  NOR U9276 ( .A(n11146), .B(n11144), .Z(n11145) );
  XOR U9277 ( .A(n11147), .B(n11148), .Z(n8314) );
  NOR U9278 ( .A(n11149), .B(n11147), .Z(n11148) );
  XOR U9279 ( .A(n11150), .B(n11151), .Z(n8317) );
  NOR U9280 ( .A(n11152), .B(n11150), .Z(n11151) );
  XOR U9281 ( .A(n11153), .B(n11154), .Z(n8320) );
  NOR U9282 ( .A(n11155), .B(n11153), .Z(n11154) );
  XOR U9283 ( .A(n11156), .B(n11157), .Z(n8323) );
  NOR U9284 ( .A(n11158), .B(n11156), .Z(n11157) );
  XOR U9285 ( .A(n11159), .B(n11160), .Z(n8326) );
  NOR U9286 ( .A(n11161), .B(n11159), .Z(n11160) );
  XOR U9287 ( .A(n11162), .B(n11163), .Z(n8329) );
  NOR U9288 ( .A(n11164), .B(n11162), .Z(n11163) );
  XOR U9289 ( .A(n11165), .B(n11166), .Z(n8332) );
  NOR U9290 ( .A(n11167), .B(n11165), .Z(n11166) );
  XOR U9291 ( .A(n11168), .B(n11169), .Z(n8335) );
  NOR U9292 ( .A(n11170), .B(n11168), .Z(n11169) );
  XOR U9293 ( .A(n11171), .B(n11172), .Z(n8338) );
  NOR U9294 ( .A(n11173), .B(n11171), .Z(n11172) );
  XOR U9295 ( .A(n11174), .B(n11175), .Z(n8341) );
  NOR U9296 ( .A(n11176), .B(n11174), .Z(n11175) );
  XOR U9297 ( .A(n11177), .B(n11178), .Z(n8344) );
  NOR U9298 ( .A(n11179), .B(n11177), .Z(n11178) );
  XOR U9299 ( .A(n11180), .B(n11181), .Z(n8347) );
  NOR U9300 ( .A(n11182), .B(n11180), .Z(n11181) );
  XOR U9301 ( .A(n11183), .B(n11184), .Z(n8350) );
  NOR U9302 ( .A(n11185), .B(n11183), .Z(n11184) );
  XOR U9303 ( .A(n11186), .B(n11187), .Z(n8353) );
  NOR U9304 ( .A(n11188), .B(n11186), .Z(n11187) );
  XOR U9305 ( .A(n11189), .B(n11190), .Z(n8356) );
  NOR U9306 ( .A(n11191), .B(n11189), .Z(n11190) );
  XOR U9307 ( .A(n11192), .B(n11193), .Z(n8359) );
  NOR U9308 ( .A(n11194), .B(n11192), .Z(n11193) );
  XOR U9309 ( .A(n11195), .B(n11196), .Z(n8362) );
  NOR U9310 ( .A(n11197), .B(n11195), .Z(n11196) );
  XOR U9311 ( .A(n11198), .B(n11199), .Z(n8365) );
  NOR U9312 ( .A(n11200), .B(n11198), .Z(n11199) );
  XOR U9313 ( .A(n11201), .B(n11202), .Z(n8368) );
  NOR U9314 ( .A(n11203), .B(n11201), .Z(n11202) );
  XOR U9315 ( .A(n11204), .B(n11205), .Z(n8371) );
  NOR U9316 ( .A(n11206), .B(n11204), .Z(n11205) );
  XOR U9317 ( .A(n11207), .B(n11208), .Z(n8374) );
  NOR U9318 ( .A(n11209), .B(n11207), .Z(n11208) );
  XOR U9319 ( .A(n11210), .B(n11211), .Z(n8377) );
  NOR U9320 ( .A(n11212), .B(n11210), .Z(n11211) );
  XOR U9321 ( .A(n11213), .B(n11214), .Z(n8380) );
  NOR U9322 ( .A(n11215), .B(n11213), .Z(n11214) );
  XOR U9323 ( .A(n11216), .B(n11217), .Z(n8383) );
  NOR U9324 ( .A(n11218), .B(n11216), .Z(n11217) );
  XOR U9325 ( .A(n11219), .B(n11220), .Z(n8386) );
  NOR U9326 ( .A(n11221), .B(n11219), .Z(n11220) );
  XOR U9327 ( .A(n11222), .B(n11223), .Z(n8389) );
  NOR U9328 ( .A(n11224), .B(n11222), .Z(n11223) );
  XOR U9329 ( .A(n11225), .B(n11226), .Z(n8392) );
  NOR U9330 ( .A(n11227), .B(n11225), .Z(n11226) );
  XOR U9331 ( .A(n11228), .B(n11229), .Z(n8395) );
  NOR U9332 ( .A(n11230), .B(n11228), .Z(n11229) );
  XOR U9333 ( .A(n11231), .B(n11232), .Z(n8398) );
  NOR U9334 ( .A(n11233), .B(n11231), .Z(n11232) );
  XOR U9335 ( .A(n11234), .B(n11235), .Z(n8401) );
  NOR U9336 ( .A(n11236), .B(n11234), .Z(n11235) );
  XOR U9337 ( .A(n11237), .B(n11238), .Z(n8404) );
  NOR U9338 ( .A(n11239), .B(n11237), .Z(n11238) );
  XOR U9339 ( .A(n11240), .B(n11241), .Z(n8407) );
  NOR U9340 ( .A(n11242), .B(n11240), .Z(n11241) );
  XOR U9341 ( .A(n11243), .B(n11244), .Z(n8410) );
  NOR U9342 ( .A(n11245), .B(n11243), .Z(n11244) );
  XOR U9343 ( .A(n11246), .B(n11247), .Z(n8413) );
  NOR U9344 ( .A(n11248), .B(n11246), .Z(n11247) );
  XOR U9345 ( .A(n11249), .B(n11250), .Z(n8416) );
  NOR U9346 ( .A(n11251), .B(n11249), .Z(n11250) );
  XOR U9347 ( .A(n11252), .B(n11253), .Z(n8419) );
  NOR U9348 ( .A(n11254), .B(n11252), .Z(n11253) );
  XOR U9349 ( .A(n11255), .B(n11256), .Z(n8422) );
  NOR U9350 ( .A(n11257), .B(n11255), .Z(n11256) );
  XOR U9351 ( .A(n11258), .B(n11259), .Z(n8425) );
  NOR U9352 ( .A(n11260), .B(n11258), .Z(n11259) );
  XOR U9353 ( .A(n11261), .B(n11262), .Z(n8428) );
  NOR U9354 ( .A(n11263), .B(n11261), .Z(n11262) );
  XOR U9355 ( .A(n11264), .B(n11265), .Z(n8431) );
  NOR U9356 ( .A(n11266), .B(n11264), .Z(n11265) );
  XOR U9357 ( .A(n11267), .B(n11268), .Z(n8434) );
  NOR U9358 ( .A(n11269), .B(n11267), .Z(n11268) );
  XOR U9359 ( .A(n11270), .B(n11271), .Z(n8437) );
  NOR U9360 ( .A(n11272), .B(n11270), .Z(n11271) );
  XOR U9361 ( .A(n11273), .B(n11274), .Z(n8440) );
  NOR U9362 ( .A(n11275), .B(n11273), .Z(n11274) );
  XOR U9363 ( .A(n11276), .B(n11277), .Z(n8443) );
  NOR U9364 ( .A(n11278), .B(n11276), .Z(n11277) );
  XOR U9365 ( .A(n11279), .B(n11280), .Z(n8446) );
  NOR U9366 ( .A(n11281), .B(n11279), .Z(n11280) );
  XOR U9367 ( .A(n11282), .B(n11283), .Z(n8449) );
  NOR U9368 ( .A(n11284), .B(n11282), .Z(n11283) );
  XOR U9369 ( .A(n11285), .B(n11286), .Z(n8452) );
  NOR U9370 ( .A(n11287), .B(n11285), .Z(n11286) );
  XOR U9371 ( .A(n11288), .B(n11289), .Z(n8455) );
  NOR U9372 ( .A(n11290), .B(n11288), .Z(n11289) );
  XOR U9373 ( .A(n11291), .B(n11292), .Z(n8458) );
  NOR U9374 ( .A(n11293), .B(n11291), .Z(n11292) );
  XOR U9375 ( .A(n11294), .B(n11295), .Z(n8461) );
  NOR U9376 ( .A(n11296), .B(n11294), .Z(n11295) );
  XOR U9377 ( .A(n11297), .B(n11298), .Z(n8464) );
  NOR U9378 ( .A(n11299), .B(n11297), .Z(n11298) );
  XOR U9379 ( .A(n11300), .B(n11301), .Z(n8467) );
  NOR U9380 ( .A(n11302), .B(n11300), .Z(n11301) );
  XOR U9381 ( .A(n11303), .B(n11304), .Z(n8470) );
  NOR U9382 ( .A(n87), .B(n11305), .Z(n11304) );
  IV U9383 ( .A(n11303), .Z(n11305) );
  XOR U9384 ( .A(n11306), .B(n11307), .Z(n8473) );
  AND U9385 ( .A(n11308), .B(n11309), .Z(n11307) );
  XOR U9386 ( .A(n11306), .B(n89), .Z(n11309) );
  XOR U9387 ( .A(n9889), .B(n9888), .Z(n89) );
  XNOR U9388 ( .A(n9886), .B(n9885), .Z(n9888) );
  XNOR U9389 ( .A(n9883), .B(n9882), .Z(n9885) );
  XNOR U9390 ( .A(n9880), .B(n9879), .Z(n9882) );
  XNOR U9391 ( .A(n9877), .B(n9876), .Z(n9879) );
  XNOR U9392 ( .A(n9874), .B(n9873), .Z(n9876) );
  XNOR U9393 ( .A(n9871), .B(n9870), .Z(n9873) );
  XNOR U9394 ( .A(n9868), .B(n9867), .Z(n9870) );
  XNOR U9395 ( .A(n9865), .B(n9864), .Z(n9867) );
  XNOR U9396 ( .A(n9862), .B(n9861), .Z(n9864) );
  XNOR U9397 ( .A(n9859), .B(n9858), .Z(n9861) );
  XNOR U9398 ( .A(n9856), .B(n9855), .Z(n9858) );
  XNOR U9399 ( .A(n9853), .B(n9852), .Z(n9855) );
  XNOR U9400 ( .A(n9850), .B(n9849), .Z(n9852) );
  XNOR U9401 ( .A(n9847), .B(n9846), .Z(n9849) );
  XNOR U9402 ( .A(n9844), .B(n9843), .Z(n9846) );
  XNOR U9403 ( .A(n9841), .B(n9840), .Z(n9843) );
  XNOR U9404 ( .A(n9838), .B(n9837), .Z(n9840) );
  XNOR U9405 ( .A(n9835), .B(n9834), .Z(n9837) );
  XNOR U9406 ( .A(n9832), .B(n9831), .Z(n9834) );
  XNOR U9407 ( .A(n9829), .B(n9828), .Z(n9831) );
  XNOR U9408 ( .A(n9826), .B(n9825), .Z(n9828) );
  XNOR U9409 ( .A(n9823), .B(n9822), .Z(n9825) );
  XNOR U9410 ( .A(n9820), .B(n9819), .Z(n9822) );
  XNOR U9411 ( .A(n9817), .B(n9816), .Z(n9819) );
  XNOR U9412 ( .A(n9814), .B(n9813), .Z(n9816) );
  XNOR U9413 ( .A(n9811), .B(n9810), .Z(n9813) );
  XNOR U9414 ( .A(n9808), .B(n9807), .Z(n9810) );
  XNOR U9415 ( .A(n9805), .B(n9804), .Z(n9807) );
  XNOR U9416 ( .A(n9802), .B(n9801), .Z(n9804) );
  XNOR U9417 ( .A(n9799), .B(n9798), .Z(n9801) );
  XNOR U9418 ( .A(n9796), .B(n9795), .Z(n9798) );
  XNOR U9419 ( .A(n9793), .B(n9792), .Z(n9795) );
  XNOR U9420 ( .A(n9790), .B(n9789), .Z(n9792) );
  XNOR U9421 ( .A(n9787), .B(n9786), .Z(n9789) );
  XNOR U9422 ( .A(n9784), .B(n9783), .Z(n9786) );
  XNOR U9423 ( .A(n9781), .B(n9780), .Z(n9783) );
  XNOR U9424 ( .A(n9778), .B(n9777), .Z(n9780) );
  XNOR U9425 ( .A(n9775), .B(n9774), .Z(n9777) );
  XNOR U9426 ( .A(n9772), .B(n9771), .Z(n9774) );
  XNOR U9427 ( .A(n9769), .B(n9768), .Z(n9771) );
  XNOR U9428 ( .A(n9766), .B(n9765), .Z(n9768) );
  XNOR U9429 ( .A(n9763), .B(n9762), .Z(n9765) );
  XNOR U9430 ( .A(n9760), .B(n9759), .Z(n9762) );
  XNOR U9431 ( .A(n9757), .B(n9756), .Z(n9759) );
  XNOR U9432 ( .A(n9754), .B(n9753), .Z(n9756) );
  XNOR U9433 ( .A(n9751), .B(n9750), .Z(n9753) );
  XNOR U9434 ( .A(n9748), .B(n9747), .Z(n9750) );
  XNOR U9435 ( .A(n9745), .B(n9744), .Z(n9747) );
  XNOR U9436 ( .A(n9742), .B(n9741), .Z(n9744) );
  XNOR U9437 ( .A(n9739), .B(n9738), .Z(n9741) );
  XNOR U9438 ( .A(n9736), .B(n9735), .Z(n9738) );
  XNOR U9439 ( .A(n9733), .B(n9732), .Z(n9735) );
  XNOR U9440 ( .A(n9730), .B(n9729), .Z(n9732) );
  XNOR U9441 ( .A(n9727), .B(n9726), .Z(n9729) );
  XNOR U9442 ( .A(n9724), .B(n9723), .Z(n9726) );
  XNOR U9443 ( .A(n9721), .B(n9720), .Z(n9723) );
  XNOR U9444 ( .A(n9718), .B(n9717), .Z(n9720) );
  XNOR U9445 ( .A(n9715), .B(n9714), .Z(n9717) );
  XNOR U9446 ( .A(n9712), .B(n9711), .Z(n9714) );
  XNOR U9447 ( .A(n9709), .B(n9708), .Z(n9711) );
  XNOR U9448 ( .A(n9706), .B(n9705), .Z(n9708) );
  XNOR U9449 ( .A(n9703), .B(n9702), .Z(n9705) );
  XNOR U9450 ( .A(n9700), .B(n9699), .Z(n9702) );
  XNOR U9451 ( .A(n9697), .B(n9696), .Z(n9699) );
  XNOR U9452 ( .A(n9694), .B(n9693), .Z(n9696) );
  XNOR U9453 ( .A(n9691), .B(n9690), .Z(n9693) );
  XNOR U9454 ( .A(n9688), .B(n9687), .Z(n9690) );
  XNOR U9455 ( .A(n9685), .B(n9684), .Z(n9687) );
  XNOR U9456 ( .A(n9682), .B(n9681), .Z(n9684) );
  XNOR U9457 ( .A(n9679), .B(n9678), .Z(n9681) );
  XNOR U9458 ( .A(n9676), .B(n9675), .Z(n9678) );
  XNOR U9459 ( .A(n9673), .B(n9672), .Z(n9675) );
  XNOR U9460 ( .A(n9670), .B(n9669), .Z(n9672) );
  XNOR U9461 ( .A(n9667), .B(n9666), .Z(n9669) );
  XNOR U9462 ( .A(n9664), .B(n9663), .Z(n9666) );
  XNOR U9463 ( .A(n9661), .B(n9660), .Z(n9663) );
  XNOR U9464 ( .A(n9658), .B(n9657), .Z(n9660) );
  XNOR U9465 ( .A(n9655), .B(n9654), .Z(n9657) );
  XNOR U9466 ( .A(n9652), .B(n9651), .Z(n9654) );
  XNOR U9467 ( .A(n9649), .B(n9648), .Z(n9651) );
  XNOR U9468 ( .A(n9646), .B(n9645), .Z(n9648) );
  XNOR U9469 ( .A(n9643), .B(n9642), .Z(n9645) );
  XNOR U9470 ( .A(n9640), .B(n9639), .Z(n9642) );
  XNOR U9471 ( .A(n9637), .B(n9636), .Z(n9639) );
  XNOR U9472 ( .A(n9634), .B(n9633), .Z(n9636) );
  XNOR U9473 ( .A(n9631), .B(n9630), .Z(n9633) );
  XNOR U9474 ( .A(n9628), .B(n9627), .Z(n9630) );
  XNOR U9475 ( .A(n9625), .B(n9624), .Z(n9627) );
  XNOR U9476 ( .A(n9622), .B(n9621), .Z(n9624) );
  XNOR U9477 ( .A(n9619), .B(n9618), .Z(n9621) );
  XNOR U9478 ( .A(n9616), .B(n9615), .Z(n9618) );
  XNOR U9479 ( .A(n9613), .B(n9612), .Z(n9615) );
  XNOR U9480 ( .A(n9610), .B(n9609), .Z(n9612) );
  XNOR U9481 ( .A(n9607), .B(n9606), .Z(n9609) );
  XNOR U9482 ( .A(n9604), .B(n9603), .Z(n9606) );
  XNOR U9483 ( .A(n9601), .B(n9600), .Z(n9603) );
  XNOR U9484 ( .A(n9598), .B(n9597), .Z(n9600) );
  XNOR U9485 ( .A(n9595), .B(n9594), .Z(n9597) );
  XNOR U9486 ( .A(n9592), .B(n9591), .Z(n9594) );
  XNOR U9487 ( .A(n9589), .B(n9588), .Z(n9591) );
  XNOR U9488 ( .A(n9586), .B(n9585), .Z(n9588) );
  XNOR U9489 ( .A(n9583), .B(n9582), .Z(n9585) );
  XNOR U9490 ( .A(n9580), .B(n9579), .Z(n9582) );
  XNOR U9491 ( .A(n9577), .B(n9576), .Z(n9579) );
  XNOR U9492 ( .A(n9574), .B(n9573), .Z(n9576) );
  XNOR U9493 ( .A(n9571), .B(n9570), .Z(n9573) );
  XNOR U9494 ( .A(n9568), .B(n9567), .Z(n9570) );
  XNOR U9495 ( .A(n9565), .B(n9564), .Z(n9567) );
  XNOR U9496 ( .A(n9562), .B(n9561), .Z(n9564) );
  XNOR U9497 ( .A(n9559), .B(n9558), .Z(n9561) );
  XNOR U9498 ( .A(n9556), .B(n9555), .Z(n9558) );
  XNOR U9499 ( .A(n9553), .B(n9552), .Z(n9555) );
  XNOR U9500 ( .A(n9550), .B(n9549), .Z(n9552) );
  XNOR U9501 ( .A(n9547), .B(n9546), .Z(n9549) );
  XNOR U9502 ( .A(n9544), .B(n9543), .Z(n9546) );
  XNOR U9503 ( .A(n9541), .B(n9540), .Z(n9543) );
  XNOR U9504 ( .A(n9538), .B(n9537), .Z(n9540) );
  XNOR U9505 ( .A(n9535), .B(n9534), .Z(n9537) );
  XNOR U9506 ( .A(n9532), .B(n9531), .Z(n9534) );
  XNOR U9507 ( .A(n9529), .B(n9528), .Z(n9531) );
  XNOR U9508 ( .A(n9526), .B(n9525), .Z(n9528) );
  XNOR U9509 ( .A(n9523), .B(n9522), .Z(n9525) );
  XNOR U9510 ( .A(n9520), .B(n9519), .Z(n9522) );
  XNOR U9511 ( .A(n9517), .B(n9516), .Z(n9519) );
  XNOR U9512 ( .A(n9514), .B(n9513), .Z(n9516) );
  XNOR U9513 ( .A(n9511), .B(n9510), .Z(n9513) );
  XNOR U9514 ( .A(n9508), .B(n9507), .Z(n9510) );
  XNOR U9515 ( .A(n9505), .B(n9504), .Z(n9507) );
  XNOR U9516 ( .A(n9502), .B(n9501), .Z(n9504) );
  XNOR U9517 ( .A(n9499), .B(n9498), .Z(n9501) );
  XNOR U9518 ( .A(n9496), .B(n9495), .Z(n9498) );
  XNOR U9519 ( .A(n9493), .B(n9492), .Z(n9495) );
  XNOR U9520 ( .A(n9490), .B(n9489), .Z(n9492) );
  XNOR U9521 ( .A(n9487), .B(n9486), .Z(n9489) );
  XNOR U9522 ( .A(n9484), .B(n9483), .Z(n9486) );
  XNOR U9523 ( .A(n9481), .B(n9480), .Z(n9483) );
  XNOR U9524 ( .A(n9478), .B(n9477), .Z(n9480) );
  XNOR U9525 ( .A(n9475), .B(n9474), .Z(n9477) );
  XNOR U9526 ( .A(n9472), .B(n9471), .Z(n9474) );
  XNOR U9527 ( .A(n9469), .B(n9468), .Z(n9471) );
  XNOR U9528 ( .A(n9466), .B(n9465), .Z(n9468) );
  XNOR U9529 ( .A(n9463), .B(n9462), .Z(n9465) );
  XNOR U9530 ( .A(n9460), .B(n9459), .Z(n9462) );
  XNOR U9531 ( .A(n9457), .B(n9456), .Z(n9459) );
  XNOR U9532 ( .A(n9454), .B(n9453), .Z(n9456) );
  XNOR U9533 ( .A(n9451), .B(n9450), .Z(n9453) );
  XNOR U9534 ( .A(n9448), .B(n9447), .Z(n9450) );
  XNOR U9535 ( .A(n9445), .B(n9444), .Z(n9447) );
  XNOR U9536 ( .A(n9442), .B(n9441), .Z(n9444) );
  XNOR U9537 ( .A(n9439), .B(n9438), .Z(n9441) );
  XNOR U9538 ( .A(n9436), .B(n9435), .Z(n9438) );
  XNOR U9539 ( .A(n9433), .B(n9432), .Z(n9435) );
  XNOR U9540 ( .A(n9430), .B(n9429), .Z(n9432) );
  XNOR U9541 ( .A(n9427), .B(n9426), .Z(n9429) );
  XNOR U9542 ( .A(n9424), .B(n9423), .Z(n9426) );
  XNOR U9543 ( .A(n9421), .B(n9420), .Z(n9423) );
  XNOR U9544 ( .A(n9418), .B(n9417), .Z(n9420) );
  XNOR U9545 ( .A(n9415), .B(n9414), .Z(n9417) );
  XNOR U9546 ( .A(n9412), .B(n9411), .Z(n9414) );
  XNOR U9547 ( .A(n9409), .B(n9408), .Z(n9411) );
  XNOR U9548 ( .A(n9406), .B(n9405), .Z(n9408) );
  XNOR U9549 ( .A(n9403), .B(n9402), .Z(n9405) );
  XNOR U9550 ( .A(n9400), .B(n9399), .Z(n9402) );
  XNOR U9551 ( .A(n9397), .B(n9396), .Z(n9399) );
  XNOR U9552 ( .A(n9394), .B(n9393), .Z(n9396) );
  XNOR U9553 ( .A(n9391), .B(n9390), .Z(n9393) );
  XNOR U9554 ( .A(n9388), .B(n9387), .Z(n9390) );
  XNOR U9555 ( .A(n9385), .B(n9384), .Z(n9387) );
  XNOR U9556 ( .A(n9382), .B(n9381), .Z(n9384) );
  XNOR U9557 ( .A(n9379), .B(n9378), .Z(n9381) );
  XNOR U9558 ( .A(n9376), .B(n9375), .Z(n9378) );
  XNOR U9559 ( .A(n9373), .B(n9372), .Z(n9375) );
  XNOR U9560 ( .A(n9370), .B(n9369), .Z(n9372) );
  XNOR U9561 ( .A(n9367), .B(n9366), .Z(n9369) );
  XNOR U9562 ( .A(n9364), .B(n9363), .Z(n9366) );
  XNOR U9563 ( .A(n9361), .B(n9360), .Z(n9363) );
  XNOR U9564 ( .A(n9358), .B(n9357), .Z(n9360) );
  XNOR U9565 ( .A(n9355), .B(n9354), .Z(n9357) );
  XNOR U9566 ( .A(n9352), .B(n9351), .Z(n9354) );
  XNOR U9567 ( .A(n9349), .B(n9348), .Z(n9351) );
  XNOR U9568 ( .A(n9346), .B(n9345), .Z(n9348) );
  XNOR U9569 ( .A(n9343), .B(n9342), .Z(n9345) );
  XNOR U9570 ( .A(n9340), .B(n9339), .Z(n9342) );
  XNOR U9571 ( .A(n9337), .B(n9336), .Z(n9339) );
  XNOR U9572 ( .A(n9334), .B(n9333), .Z(n9336) );
  XNOR U9573 ( .A(n9331), .B(n9330), .Z(n9333) );
  XNOR U9574 ( .A(n9328), .B(n9327), .Z(n9330) );
  XNOR U9575 ( .A(n9325), .B(n9324), .Z(n9327) );
  XNOR U9576 ( .A(n9322), .B(n9321), .Z(n9324) );
  XNOR U9577 ( .A(n9319), .B(n9318), .Z(n9321) );
  XNOR U9578 ( .A(n9316), .B(n9315), .Z(n9318) );
  XNOR U9579 ( .A(n9313), .B(n9312), .Z(n9315) );
  XNOR U9580 ( .A(n9310), .B(n9309), .Z(n9312) );
  XNOR U9581 ( .A(n9307), .B(n9306), .Z(n9309) );
  XNOR U9582 ( .A(n9304), .B(n9303), .Z(n9306) );
  XNOR U9583 ( .A(n9301), .B(n9300), .Z(n9303) );
  XNOR U9584 ( .A(n9298), .B(n9297), .Z(n9300) );
  XNOR U9585 ( .A(n9295), .B(n9294), .Z(n9297) );
  XNOR U9586 ( .A(n9292), .B(n9291), .Z(n9294) );
  XNOR U9587 ( .A(n9289), .B(n9288), .Z(n9291) );
  XNOR U9588 ( .A(n9286), .B(n9285), .Z(n9288) );
  XNOR U9589 ( .A(n9283), .B(n9282), .Z(n9285) );
  XNOR U9590 ( .A(n9280), .B(n9279), .Z(n9282) );
  XNOR U9591 ( .A(n9277), .B(n9276), .Z(n9279) );
  XNOR U9592 ( .A(n9274), .B(n9273), .Z(n9276) );
  XNOR U9593 ( .A(n9271), .B(n9270), .Z(n9273) );
  XNOR U9594 ( .A(n9268), .B(n9267), .Z(n9270) );
  XNOR U9595 ( .A(n9265), .B(n9264), .Z(n9267) );
  XNOR U9596 ( .A(n9262), .B(n9261), .Z(n9264) );
  XNOR U9597 ( .A(n9259), .B(n9258), .Z(n9261) );
  XNOR U9598 ( .A(n9256), .B(n9255), .Z(n9258) );
  XNOR U9599 ( .A(n9253), .B(n9252), .Z(n9255) );
  XNOR U9600 ( .A(n9250), .B(n9249), .Z(n9252) );
  XNOR U9601 ( .A(n9247), .B(n9246), .Z(n9249) );
  XNOR U9602 ( .A(n9244), .B(n9243), .Z(n9246) );
  XNOR U9603 ( .A(n9241), .B(n9240), .Z(n9243) );
  XNOR U9604 ( .A(n9238), .B(n9237), .Z(n9240) );
  XNOR U9605 ( .A(n9235), .B(n9234), .Z(n9237) );
  XNOR U9606 ( .A(n9232), .B(n9231), .Z(n9234) );
  XNOR U9607 ( .A(n9229), .B(n9228), .Z(n9231) );
  XNOR U9608 ( .A(n9226), .B(n9225), .Z(n9228) );
  XNOR U9609 ( .A(n9223), .B(n9222), .Z(n9225) );
  XNOR U9610 ( .A(n9220), .B(n9219), .Z(n9222) );
  XNOR U9611 ( .A(n9217), .B(n9216), .Z(n9219) );
  XNOR U9612 ( .A(n9214), .B(n9213), .Z(n9216) );
  XNOR U9613 ( .A(n9211), .B(n9210), .Z(n9213) );
  XNOR U9614 ( .A(n9208), .B(n9207), .Z(n9210) );
  XNOR U9615 ( .A(n9205), .B(n9204), .Z(n9207) );
  XNOR U9616 ( .A(n9202), .B(n9201), .Z(n9204) );
  XNOR U9617 ( .A(n9199), .B(n9198), .Z(n9201) );
  XNOR U9618 ( .A(n9196), .B(n9195), .Z(n9198) );
  XNOR U9619 ( .A(n9193), .B(n9192), .Z(n9195) );
  XNOR U9620 ( .A(n9190), .B(n9189), .Z(n9192) );
  XNOR U9621 ( .A(n9187), .B(n9186), .Z(n9189) );
  XNOR U9622 ( .A(n9184), .B(n9183), .Z(n9186) );
  XNOR U9623 ( .A(n9181), .B(n9180), .Z(n9183) );
  XNOR U9624 ( .A(n9178), .B(n9177), .Z(n9180) );
  XNOR U9625 ( .A(n9175), .B(n9174), .Z(n9177) );
  XNOR U9626 ( .A(n9172), .B(n9171), .Z(n9174) );
  XNOR U9627 ( .A(n9169), .B(n9168), .Z(n9171) );
  XNOR U9628 ( .A(n9166), .B(n9165), .Z(n9168) );
  XNOR U9629 ( .A(n9163), .B(n9162), .Z(n9165) );
  XNOR U9630 ( .A(n9160), .B(n9159), .Z(n9162) );
  XNOR U9631 ( .A(n9157), .B(n9156), .Z(n9159) );
  XNOR U9632 ( .A(n9154), .B(n9153), .Z(n9156) );
  XNOR U9633 ( .A(n9151), .B(n9150), .Z(n9153) );
  XNOR U9634 ( .A(n9148), .B(n9147), .Z(n9150) );
  XNOR U9635 ( .A(n9145), .B(n9144), .Z(n9147) );
  XNOR U9636 ( .A(n9142), .B(n9141), .Z(n9144) );
  XNOR U9637 ( .A(n9139), .B(n9138), .Z(n9141) );
  XNOR U9638 ( .A(n9136), .B(n9135), .Z(n9138) );
  XNOR U9639 ( .A(n9133), .B(n9132), .Z(n9135) );
  XNOR U9640 ( .A(n9130), .B(n9129), .Z(n9132) );
  XNOR U9641 ( .A(n9127), .B(n9126), .Z(n9129) );
  XNOR U9642 ( .A(n9124), .B(n9123), .Z(n9126) );
  XNOR U9643 ( .A(n9121), .B(n9120), .Z(n9123) );
  XNOR U9644 ( .A(n9118), .B(n9117), .Z(n9120) );
  XNOR U9645 ( .A(n9115), .B(n9114), .Z(n9117) );
  XNOR U9646 ( .A(n9112), .B(n9111), .Z(n9114) );
  XNOR U9647 ( .A(n9109), .B(n9108), .Z(n9111) );
  XNOR U9648 ( .A(n9106), .B(n9105), .Z(n9108) );
  XNOR U9649 ( .A(n9103), .B(n9102), .Z(n9105) );
  XNOR U9650 ( .A(n9100), .B(n9099), .Z(n9102) );
  XNOR U9651 ( .A(n9097), .B(n9096), .Z(n9099) );
  XNOR U9652 ( .A(n9094), .B(n9093), .Z(n9096) );
  XNOR U9653 ( .A(n9091), .B(n9090), .Z(n9093) );
  XNOR U9654 ( .A(n9088), .B(n9087), .Z(n9090) );
  XNOR U9655 ( .A(n9085), .B(n9084), .Z(n9087) );
  XNOR U9656 ( .A(n9082), .B(n9081), .Z(n9084) );
  XNOR U9657 ( .A(n9079), .B(n9078), .Z(n9081) );
  XNOR U9658 ( .A(n9076), .B(n9075), .Z(n9078) );
  XNOR U9659 ( .A(n9073), .B(n9072), .Z(n9075) );
  XNOR U9660 ( .A(n9070), .B(n9069), .Z(n9072) );
  XNOR U9661 ( .A(n9067), .B(n9066), .Z(n9069) );
  XNOR U9662 ( .A(n9064), .B(n9063), .Z(n9066) );
  XNOR U9663 ( .A(n9061), .B(n9060), .Z(n9063) );
  XNOR U9664 ( .A(n9058), .B(n9057), .Z(n9060) );
  XNOR U9665 ( .A(n9055), .B(n9054), .Z(n9057) );
  XNOR U9666 ( .A(n9052), .B(n9051), .Z(n9054) );
  XNOR U9667 ( .A(n9049), .B(n9048), .Z(n9051) );
  XNOR U9668 ( .A(n9046), .B(n9045), .Z(n9048) );
  XNOR U9669 ( .A(n9043), .B(n9042), .Z(n9045) );
  XNOR U9670 ( .A(n9040), .B(n9039), .Z(n9042) );
  XNOR U9671 ( .A(n9037), .B(n9036), .Z(n9039) );
  XNOR U9672 ( .A(n9034), .B(n9033), .Z(n9036) );
  XNOR U9673 ( .A(n9031), .B(n9030), .Z(n9033) );
  XNOR U9674 ( .A(n9028), .B(n9027), .Z(n9030) );
  XNOR U9675 ( .A(n9025), .B(n9024), .Z(n9027) );
  XNOR U9676 ( .A(n9022), .B(n9021), .Z(n9024) );
  XNOR U9677 ( .A(n9019), .B(n9018), .Z(n9021) );
  XNOR U9678 ( .A(n9016), .B(n9015), .Z(n9018) );
  XNOR U9679 ( .A(n9013), .B(n9012), .Z(n9015) );
  XNOR U9680 ( .A(n9010), .B(n9009), .Z(n9012) );
  XNOR U9681 ( .A(n9007), .B(n9006), .Z(n9009) );
  XNOR U9682 ( .A(n9004), .B(n9003), .Z(n9006) );
  XNOR U9683 ( .A(n9001), .B(n9000), .Z(n9003) );
  XNOR U9684 ( .A(n8998), .B(n8997), .Z(n9000) );
  XNOR U9685 ( .A(n8995), .B(n8994), .Z(n8997) );
  XNOR U9686 ( .A(n8992), .B(n8991), .Z(n8994) );
  XNOR U9687 ( .A(n8989), .B(n8988), .Z(n8991) );
  XNOR U9688 ( .A(n8986), .B(n8985), .Z(n8988) );
  XNOR U9689 ( .A(n8983), .B(n8982), .Z(n8985) );
  XNOR U9690 ( .A(n8980), .B(n8979), .Z(n8982) );
  XNOR U9691 ( .A(n8977), .B(n8976), .Z(n8979) );
  XNOR U9692 ( .A(n8974), .B(n8973), .Z(n8976) );
  XNOR U9693 ( .A(n8971), .B(n8970), .Z(n8973) );
  XNOR U9694 ( .A(n8968), .B(n8967), .Z(n8970) );
  XNOR U9695 ( .A(n8965), .B(n8964), .Z(n8967) );
  XNOR U9696 ( .A(n8962), .B(n8961), .Z(n8964) );
  XNOR U9697 ( .A(n8959), .B(n8958), .Z(n8961) );
  XNOR U9698 ( .A(n8956), .B(n8955), .Z(n8958) );
  XNOR U9699 ( .A(n8953), .B(n8952), .Z(n8955) );
  XNOR U9700 ( .A(n8950), .B(n8949), .Z(n8952) );
  XNOR U9701 ( .A(n8947), .B(n8946), .Z(n8949) );
  XNOR U9702 ( .A(n8944), .B(n8943), .Z(n8946) );
  XNOR U9703 ( .A(n8941), .B(n8940), .Z(n8943) );
  XNOR U9704 ( .A(n8938), .B(n8937), .Z(n8940) );
  XNOR U9705 ( .A(n8935), .B(n8934), .Z(n8937) );
  XNOR U9706 ( .A(n8932), .B(n8931), .Z(n8934) );
  XNOR U9707 ( .A(n8929), .B(n8928), .Z(n8931) );
  XNOR U9708 ( .A(n8926), .B(n8925), .Z(n8928) );
  XNOR U9709 ( .A(n8923), .B(n8922), .Z(n8925) );
  XNOR U9710 ( .A(n8920), .B(n8919), .Z(n8922) );
  XNOR U9711 ( .A(n8917), .B(n8916), .Z(n8919) );
  XNOR U9712 ( .A(n8914), .B(n8913), .Z(n8916) );
  XNOR U9713 ( .A(n8911), .B(n8910), .Z(n8913) );
  XNOR U9714 ( .A(n8908), .B(n8907), .Z(n8910) );
  XNOR U9715 ( .A(n8905), .B(n8904), .Z(n8907) );
  XNOR U9716 ( .A(n8902), .B(n8901), .Z(n8904) );
  XNOR U9717 ( .A(n8899), .B(n8898), .Z(n8901) );
  XNOR U9718 ( .A(n8896), .B(n8895), .Z(n8898) );
  XNOR U9719 ( .A(n8893), .B(n8892), .Z(n8895) );
  XNOR U9720 ( .A(n8890), .B(n8889), .Z(n8892) );
  XNOR U9721 ( .A(n8887), .B(n8886), .Z(n8889) );
  XNOR U9722 ( .A(n8884), .B(n8883), .Z(n8886) );
  XNOR U9723 ( .A(n8881), .B(n8880), .Z(n8883) );
  XNOR U9724 ( .A(n8878), .B(n8877), .Z(n8880) );
  XNOR U9725 ( .A(n8875), .B(n8874), .Z(n8877) );
  XNOR U9726 ( .A(n8872), .B(n8871), .Z(n8874) );
  XNOR U9727 ( .A(n8869), .B(n8868), .Z(n8871) );
  XNOR U9728 ( .A(n8866), .B(n8865), .Z(n8868) );
  XNOR U9729 ( .A(n8863), .B(n8862), .Z(n8865) );
  XNOR U9730 ( .A(n8860), .B(n8859), .Z(n8862) );
  XNOR U9731 ( .A(n8857), .B(n8856), .Z(n8859) );
  XNOR U9732 ( .A(n8854), .B(n8853), .Z(n8856) );
  XNOR U9733 ( .A(n8851), .B(n8850), .Z(n8853) );
  XNOR U9734 ( .A(n8848), .B(n8847), .Z(n8850) );
  XNOR U9735 ( .A(n8845), .B(n8844), .Z(n8847) );
  XNOR U9736 ( .A(n8842), .B(n8841), .Z(n8844) );
  XNOR U9737 ( .A(n8839), .B(n8838), .Z(n8841) );
  XNOR U9738 ( .A(n8836), .B(n8835), .Z(n8838) );
  XNOR U9739 ( .A(n8833), .B(n8832), .Z(n8835) );
  XNOR U9740 ( .A(n8830), .B(n8829), .Z(n8832) );
  XNOR U9741 ( .A(n8827), .B(n8826), .Z(n8829) );
  XNOR U9742 ( .A(n8824), .B(n8823), .Z(n8826) );
  XNOR U9743 ( .A(n8821), .B(n8820), .Z(n8823) );
  XNOR U9744 ( .A(n8818), .B(n8817), .Z(n8820) );
  XNOR U9745 ( .A(n8815), .B(n8814), .Z(n8817) );
  XNOR U9746 ( .A(n8812), .B(n8811), .Z(n8814) );
  XNOR U9747 ( .A(n8809), .B(n8808), .Z(n8811) );
  XNOR U9748 ( .A(n8806), .B(n8805), .Z(n8808) );
  XNOR U9749 ( .A(n8803), .B(n8802), .Z(n8805) );
  XNOR U9750 ( .A(n8800), .B(n8799), .Z(n8802) );
  XNOR U9751 ( .A(n8797), .B(n8796), .Z(n8799) );
  XNOR U9752 ( .A(n8794), .B(n8793), .Z(n8796) );
  XNOR U9753 ( .A(n8791), .B(n8790), .Z(n8793) );
  XNOR U9754 ( .A(n8788), .B(n8787), .Z(n8790) );
  XNOR U9755 ( .A(n8785), .B(n8784), .Z(n8787) );
  XNOR U9756 ( .A(n8782), .B(n8781), .Z(n8784) );
  XNOR U9757 ( .A(n8779), .B(n8778), .Z(n8781) );
  XNOR U9758 ( .A(n8776), .B(n8775), .Z(n8778) );
  XNOR U9759 ( .A(n8773), .B(n8772), .Z(n8775) );
  XNOR U9760 ( .A(n8770), .B(n8769), .Z(n8772) );
  XNOR U9761 ( .A(n8767), .B(n8766), .Z(n8769) );
  XNOR U9762 ( .A(n8764), .B(n8763), .Z(n8766) );
  XNOR U9763 ( .A(n8761), .B(n8760), .Z(n8763) );
  XNOR U9764 ( .A(n8758), .B(n8757), .Z(n8760) );
  XNOR U9765 ( .A(n8755), .B(n8754), .Z(n8757) );
  XNOR U9766 ( .A(n8752), .B(n8751), .Z(n8754) );
  XNOR U9767 ( .A(n8749), .B(n8748), .Z(n8751) );
  XNOR U9768 ( .A(n8746), .B(n8745), .Z(n8748) );
  XNOR U9769 ( .A(n8743), .B(n8742), .Z(n8745) );
  XNOR U9770 ( .A(n8740), .B(n8739), .Z(n8742) );
  XNOR U9771 ( .A(n8737), .B(n8736), .Z(n8739) );
  XNOR U9772 ( .A(n8734), .B(n8733), .Z(n8736) );
  XNOR U9773 ( .A(n8731), .B(n8730), .Z(n8733) );
  XNOR U9774 ( .A(n8728), .B(n8727), .Z(n8730) );
  XNOR U9775 ( .A(n8725), .B(n8724), .Z(n8727) );
  XNOR U9776 ( .A(n8722), .B(n8721), .Z(n8724) );
  XNOR U9777 ( .A(n8719), .B(n8718), .Z(n8721) );
  XNOR U9778 ( .A(n8716), .B(n8715), .Z(n8718) );
  XOR U9779 ( .A(n11310), .B(n8712), .Z(n8715) );
  XOR U9780 ( .A(n8710), .B(n8709), .Z(n8712) );
  XOR U9781 ( .A(n8707), .B(n8706), .Z(n8709) );
  XOR U9782 ( .A(n8703), .B(n8704), .Z(n8706) );
  AND U9783 ( .A(n11311), .B(n11312), .Z(n8704) );
  XOR U9784 ( .A(n8700), .B(n8701), .Z(n8703) );
  AND U9785 ( .A(n11313), .B(n11314), .Z(n8701) );
  XOR U9786 ( .A(n8697), .B(n8698), .Z(n8700) );
  AND U9787 ( .A(n11315), .B(n11316), .Z(n8698) );
  XOR U9788 ( .A(n8694), .B(n8695), .Z(n8697) );
  AND U9789 ( .A(n11317), .B(n11318), .Z(n8695) );
  XNOR U9790 ( .A(n8478), .B(n8692), .Z(n8694) );
  AND U9791 ( .A(n11319), .B(n11320), .Z(n8692) );
  XOR U9792 ( .A(n8480), .B(n8479), .Z(n8478) );
  AND U9793 ( .A(n11321), .B(n11322), .Z(n8479) );
  XOR U9794 ( .A(n8482), .B(n8481), .Z(n8480) );
  AND U9795 ( .A(n11323), .B(n11324), .Z(n8481) );
  XOR U9796 ( .A(n8484), .B(n8483), .Z(n8482) );
  AND U9797 ( .A(n11325), .B(n11326), .Z(n8483) );
  XOR U9798 ( .A(n8486), .B(n8485), .Z(n8484) );
  AND U9799 ( .A(n11327), .B(n11328), .Z(n8485) );
  XOR U9800 ( .A(n8488), .B(n8487), .Z(n8486) );
  AND U9801 ( .A(n11329), .B(n11330), .Z(n8487) );
  XOR U9802 ( .A(n8490), .B(n8489), .Z(n8488) );
  AND U9803 ( .A(n11331), .B(n11332), .Z(n8489) );
  XOR U9804 ( .A(n8492), .B(n8491), .Z(n8490) );
  AND U9805 ( .A(n11333), .B(n11334), .Z(n8491) );
  XOR U9806 ( .A(n8494), .B(n8493), .Z(n8492) );
  AND U9807 ( .A(n11335), .B(n11336), .Z(n8493) );
  XOR U9808 ( .A(n8496), .B(n8495), .Z(n8494) );
  AND U9809 ( .A(n11337), .B(n11338), .Z(n8495) );
  XOR U9810 ( .A(n8498), .B(n8497), .Z(n8496) );
  AND U9811 ( .A(n11339), .B(n11340), .Z(n8497) );
  XOR U9812 ( .A(n8500), .B(n8499), .Z(n8498) );
  AND U9813 ( .A(n11341), .B(n11342), .Z(n8499) );
  XOR U9814 ( .A(n8502), .B(n8501), .Z(n8500) );
  AND U9815 ( .A(n11343), .B(n11344), .Z(n8501) );
  XOR U9816 ( .A(n8504), .B(n8503), .Z(n8502) );
  AND U9817 ( .A(n11345), .B(n11346), .Z(n8503) );
  XOR U9818 ( .A(n8506), .B(n8505), .Z(n8504) );
  AND U9819 ( .A(n11347), .B(n11348), .Z(n8505) );
  XOR U9820 ( .A(n8508), .B(n8507), .Z(n8506) );
  AND U9821 ( .A(n11349), .B(n11350), .Z(n8507) );
  XOR U9822 ( .A(n8510), .B(n8509), .Z(n8508) );
  AND U9823 ( .A(n11351), .B(n11352), .Z(n8509) );
  XOR U9824 ( .A(n8512), .B(n8511), .Z(n8510) );
  AND U9825 ( .A(n11353), .B(n11354), .Z(n8511) );
  XOR U9826 ( .A(n8514), .B(n8513), .Z(n8512) );
  AND U9827 ( .A(n11355), .B(n11356), .Z(n8513) );
  XOR U9828 ( .A(n8516), .B(n8515), .Z(n8514) );
  AND U9829 ( .A(n11357), .B(n11358), .Z(n8515) );
  XOR U9830 ( .A(n8518), .B(n8517), .Z(n8516) );
  AND U9831 ( .A(n11359), .B(n11360), .Z(n8517) );
  XOR U9832 ( .A(n8520), .B(n8519), .Z(n8518) );
  AND U9833 ( .A(n11361), .B(n11362), .Z(n8519) );
  XOR U9834 ( .A(n8522), .B(n8521), .Z(n8520) );
  AND U9835 ( .A(n11363), .B(n11364), .Z(n8521) );
  XOR U9836 ( .A(n8524), .B(n8523), .Z(n8522) );
  AND U9837 ( .A(n11365), .B(n11366), .Z(n8523) );
  XOR U9838 ( .A(n8526), .B(n8525), .Z(n8524) );
  AND U9839 ( .A(n11367), .B(n11368), .Z(n8525) );
  XOR U9840 ( .A(n8528), .B(n8527), .Z(n8526) );
  AND U9841 ( .A(n11369), .B(n11370), .Z(n8527) );
  XOR U9842 ( .A(n8530), .B(n8529), .Z(n8528) );
  AND U9843 ( .A(n11371), .B(n11372), .Z(n8529) );
  XOR U9844 ( .A(n8532), .B(n8531), .Z(n8530) );
  AND U9845 ( .A(n11373), .B(n11374), .Z(n8531) );
  XOR U9846 ( .A(n8534), .B(n8533), .Z(n8532) );
  AND U9847 ( .A(n11375), .B(n11376), .Z(n8533) );
  XOR U9848 ( .A(n8536), .B(n8535), .Z(n8534) );
  AND U9849 ( .A(n11377), .B(n11378), .Z(n8535) );
  XOR U9850 ( .A(n8538), .B(n8537), .Z(n8536) );
  AND U9851 ( .A(n11379), .B(n11380), .Z(n8537) );
  XOR U9852 ( .A(n8540), .B(n8539), .Z(n8538) );
  AND U9853 ( .A(n11381), .B(n11382), .Z(n8539) );
  XOR U9854 ( .A(n8542), .B(n8541), .Z(n8540) );
  AND U9855 ( .A(n11383), .B(n11384), .Z(n8541) );
  XOR U9856 ( .A(n8544), .B(n8543), .Z(n8542) );
  AND U9857 ( .A(n11385), .B(n11386), .Z(n8543) );
  XOR U9858 ( .A(n8546), .B(n8545), .Z(n8544) );
  AND U9859 ( .A(n11387), .B(n11388), .Z(n8545) );
  XOR U9860 ( .A(n8548), .B(n8547), .Z(n8546) );
  AND U9861 ( .A(n11389), .B(n11390), .Z(n8547) );
  XOR U9862 ( .A(n8550), .B(n8549), .Z(n8548) );
  AND U9863 ( .A(n11391), .B(n11392), .Z(n8549) );
  XOR U9864 ( .A(n8552), .B(n8551), .Z(n8550) );
  AND U9865 ( .A(n11393), .B(n11394), .Z(n8551) );
  XOR U9866 ( .A(n8554), .B(n8553), .Z(n8552) );
  AND U9867 ( .A(n11395), .B(n11396), .Z(n8553) );
  XOR U9868 ( .A(n8556), .B(n8555), .Z(n8554) );
  AND U9869 ( .A(n11397), .B(n11398), .Z(n8555) );
  XOR U9870 ( .A(n8558), .B(n8557), .Z(n8556) );
  AND U9871 ( .A(n11399), .B(n11400), .Z(n8557) );
  XOR U9872 ( .A(n8561), .B(n8559), .Z(n8558) );
  AND U9873 ( .A(n11401), .B(n11402), .Z(n8559) );
  XOR U9874 ( .A(n8582), .B(n8562), .Z(n8561) );
  AND U9875 ( .A(n11403), .B(n11404), .Z(n8562) );
  XOR U9876 ( .A(n8578), .B(n8583), .Z(n8582) );
  AND U9877 ( .A(n11405), .B(n11406), .Z(n8583) );
  XOR U9878 ( .A(n8580), .B(n8579), .Z(n8578) );
  AND U9879 ( .A(n11407), .B(n11408), .Z(n8579) );
  XOR U9880 ( .A(n8567), .B(n8581), .Z(n8580) );
  AND U9881 ( .A(n11409), .B(n11410), .Z(n8581) );
  XOR U9882 ( .A(n8569), .B(n8568), .Z(n8567) );
  AND U9883 ( .A(n11411), .B(n11412), .Z(n8568) );
  XOR U9884 ( .A(n8572), .B(n8570), .Z(n8569) );
  AND U9885 ( .A(n11413), .B(n11414), .Z(n8570) );
  XOR U9886 ( .A(n8574), .B(n8573), .Z(n8572) );
  AND U9887 ( .A(n11415), .B(n11416), .Z(n8573) );
  XOR U9888 ( .A(n8592), .B(n8575), .Z(n8574) );
  AND U9889 ( .A(n11417), .B(n11418), .Z(n8575) );
  XNOR U9890 ( .A(n8599), .B(n8593), .Z(n8592) );
  AND U9891 ( .A(n11419), .B(n11420), .Z(n8593) );
  XOR U9892 ( .A(n8598), .B(n8590), .Z(n8599) );
  AND U9893 ( .A(n11421), .B(n11422), .Z(n8590) );
  XOR U9894 ( .A(n8691), .B(n8589), .Z(n8598) );
  AND U9895 ( .A(n11423), .B(n11424), .Z(n8589) );
  XNOR U9896 ( .A(n8610), .B(n8588), .Z(n8691) );
  AND U9897 ( .A(n11425), .B(n11426), .Z(n8588) );
  XNOR U9898 ( .A(n8617), .B(n8611), .Z(n8610) );
  AND U9899 ( .A(n11427), .B(n11428), .Z(n8611) );
  XOR U9900 ( .A(n8616), .B(n8608), .Z(n8617) );
  AND U9901 ( .A(n11429), .B(n11430), .Z(n8608) );
  XOR U9902 ( .A(n8690), .B(n8607), .Z(n8616) );
  AND U9903 ( .A(n11431), .B(n11432), .Z(n8607) );
  XNOR U9904 ( .A(n8628), .B(n8606), .Z(n8690) );
  AND U9905 ( .A(n11433), .B(n11434), .Z(n8606) );
  XNOR U9906 ( .A(n8635), .B(n8629), .Z(n8628) );
  AND U9907 ( .A(n11435), .B(n11436), .Z(n8629) );
  XOR U9908 ( .A(n8634), .B(n8626), .Z(n8635) );
  AND U9909 ( .A(n11437), .B(n11438), .Z(n8626) );
  XOR U9910 ( .A(n8689), .B(n8625), .Z(n8634) );
  AND U9911 ( .A(n11439), .B(n11440), .Z(n8625) );
  XNOR U9912 ( .A(n8646), .B(n8624), .Z(n8689) );
  AND U9913 ( .A(n11441), .B(n11442), .Z(n8624) );
  XNOR U9914 ( .A(n8653), .B(n8647), .Z(n8646) );
  AND U9915 ( .A(n11443), .B(n11444), .Z(n8647) );
  XOR U9916 ( .A(n8652), .B(n8644), .Z(n8653) );
  AND U9917 ( .A(n11445), .B(n11446), .Z(n8644) );
  XOR U9918 ( .A(n8688), .B(n8643), .Z(n8652) );
  AND U9919 ( .A(n11447), .B(n11448), .Z(n8643) );
  XNOR U9920 ( .A(n11449), .B(n11450), .Z(n8688) );
  XOR U9921 ( .A(n8686), .B(n8687), .Z(n11450) );
  AND U9922 ( .A(n11451), .B(n11452), .Z(n8687) );
  AND U9923 ( .A(n11453), .B(n11454), .Z(n8686) );
  XOR U9924 ( .A(n11455), .B(n8642), .Z(n11449) );
  AND U9925 ( .A(n11456), .B(n11457), .Z(n8642) );
  XOR U9926 ( .A(n11458), .B(n11459), .Z(n11455) );
  XOR U9927 ( .A(n11460), .B(n11461), .Z(n11459) );
  XOR U9928 ( .A(n8679), .B(n8680), .Z(n11461) );
  AND U9929 ( .A(n11462), .B(n11463), .Z(n8680) );
  AND U9930 ( .A(n11464), .B(n11465), .Z(n8679) );
  XOR U9931 ( .A(n8673), .B(n8678), .Z(n11460) );
  AND U9932 ( .A(n11466), .B(n11467), .Z(n8678) );
  AND U9933 ( .A(n11468), .B(n11469), .Z(n8673) );
  XOR U9934 ( .A(n11470), .B(n11471), .Z(n11458) );
  XOR U9935 ( .A(n8681), .B(n8684), .Z(n11471) );
  AND U9936 ( .A(n11472), .B(n11473), .Z(n8684) );
  AND U9937 ( .A(n11474), .B(n11475), .Z(n8681) );
  XOR U9938 ( .A(n11476), .B(n8685), .Z(n11470) );
  AND U9939 ( .A(n11477), .B(n11478), .Z(n8685) );
  XOR U9940 ( .A(n11479), .B(n11480), .Z(n11476) );
  XOR U9941 ( .A(n11481), .B(n11482), .Z(n11480) );
  XOR U9942 ( .A(n8666), .B(n8667), .Z(n11482) );
  AND U9943 ( .A(n11483), .B(n11484), .Z(n8667) );
  AND U9944 ( .A(n11485), .B(n11486), .Z(n8666) );
  XNOR U9945 ( .A(n8664), .B(n8663), .Z(n11481) );
  IV U9946 ( .A(n11487), .Z(n8663) );
  AND U9947 ( .A(n11488), .B(n11489), .Z(n11487) );
  AND U9948 ( .A(n11490), .B(n11491), .Z(n8664) );
  XOR U9949 ( .A(n11492), .B(n11493), .Z(n11479) );
  XOR U9950 ( .A(n8670), .B(n8671), .Z(n11493) );
  AND U9951 ( .A(n11494), .B(n11495), .Z(n8671) );
  AND U9952 ( .A(n11496), .B(n11497), .Z(n8670) );
  XOR U9953 ( .A(n8665), .B(n8672), .Z(n11492) );
  AND U9954 ( .A(n11498), .B(n11499), .Z(n8672) );
  XNOR U9955 ( .A(n11500), .B(n11501), .Z(n8665) );
  AND U9956 ( .A(n11502), .B(n11503), .Z(n11501) );
  NOR U9957 ( .A(n11504), .B(n11505), .Z(n11503) );
  NOR U9958 ( .A(n11506), .B(n11507), .Z(n11502) );
  AND U9959 ( .A(n11508), .B(n11509), .Z(n11507) );
  AND U9960 ( .A(n11510), .B(n11511), .Z(n11500) );
  NOR U9961 ( .A(n11512), .B(n11513), .Z(n11511) );
  AND U9962 ( .A(n11505), .B(n11514), .Z(n11513) );
  AND U9963 ( .A(n11506), .B(n11515), .Z(n11512) );
  NOR U9964 ( .A(n11516), .B(n11517), .Z(n11510) );
  XOR U9965 ( .A(n11518), .B(n11519), .Z(n11517) );
  AND U9966 ( .A(n11520), .B(n11521), .Z(n11519) );
  NOR U9967 ( .A(n11522), .B(n11523), .Z(n11521) );
  NOR U9968 ( .A(n11524), .B(n11525), .Z(n11520) );
  AND U9969 ( .A(n11526), .B(n11527), .Z(n11525) );
  AND U9970 ( .A(n11528), .B(n11529), .Z(n11518) );
  NOR U9971 ( .A(n11530), .B(n11531), .Z(n11529) );
  AND U9972 ( .A(n11523), .B(n11532), .Z(n11531) );
  AND U9973 ( .A(n11524), .B(n11533), .Z(n11530) );
  NOR U9974 ( .A(n11534), .B(n11535), .Z(n11528) );
  AND U9975 ( .A(n11536), .B(n11537), .Z(n11535) );
  AND U9976 ( .A(n11538), .B(n11539), .Z(n11537) );
  AND U9977 ( .A(n11540), .B(n11541), .Z(n11539) );
  NOR U9978 ( .A(n11542), .B(n11543), .Z(n11540) );
  NOR U9979 ( .A(n11544), .B(n11545), .Z(n11538) );
  AND U9980 ( .A(n11546), .B(n11547), .Z(n11536) );
  NOR U9981 ( .A(n11548), .B(n11549), .Z(n11547) );
  NOR U9982 ( .A(n11550), .B(n11551), .Z(n11546) );
  AND U9983 ( .A(n11522), .B(n11552), .Z(n11534) );
  AND U9984 ( .A(n11504), .B(n11553), .Z(n11516) );
  XOR U9985 ( .A(n11554), .B(n11555), .Z(n8707) );
  AND U9986 ( .A(n11554), .B(n11556), .Z(n11555) );
  XNOR U9987 ( .A(n11557), .B(n11558), .Z(n8710) );
  AND U9988 ( .A(n11557), .B(n11559), .Z(n11558) );
  IV U9989 ( .A(n8713), .Z(n11310) );
  XNOR U9990 ( .A(n11560), .B(n11561), .Z(n8713) );
  AND U9991 ( .A(n11560), .B(n11562), .Z(n11561) );
  XNOR U9992 ( .A(n11563), .B(n11564), .Z(n8716) );
  AND U9993 ( .A(n11563), .B(n11565), .Z(n11564) );
  XNOR U9994 ( .A(n11566), .B(n11567), .Z(n8719) );
  AND U9995 ( .A(n11568), .B(n11566), .Z(n11567) );
  XOR U9996 ( .A(n11569), .B(n11570), .Z(n8722) );
  NOR U9997 ( .A(n11571), .B(n11569), .Z(n11570) );
  XOR U9998 ( .A(n11572), .B(n11573), .Z(n8725) );
  NOR U9999 ( .A(n11574), .B(n11572), .Z(n11573) );
  XOR U10000 ( .A(n11575), .B(n11576), .Z(n8728) );
  NOR U10001 ( .A(n11577), .B(n11575), .Z(n11576) );
  XOR U10002 ( .A(n11578), .B(n11579), .Z(n8731) );
  NOR U10003 ( .A(n11580), .B(n11578), .Z(n11579) );
  XOR U10004 ( .A(n11581), .B(n11582), .Z(n8734) );
  NOR U10005 ( .A(n11583), .B(n11581), .Z(n11582) );
  XOR U10006 ( .A(n11584), .B(n11585), .Z(n8737) );
  NOR U10007 ( .A(n11586), .B(n11584), .Z(n11585) );
  XOR U10008 ( .A(n11587), .B(n11588), .Z(n8740) );
  NOR U10009 ( .A(n11589), .B(n11587), .Z(n11588) );
  XOR U10010 ( .A(n11590), .B(n11591), .Z(n8743) );
  NOR U10011 ( .A(n11592), .B(n11590), .Z(n11591) );
  XOR U10012 ( .A(n11593), .B(n11594), .Z(n8746) );
  NOR U10013 ( .A(n11595), .B(n11593), .Z(n11594) );
  XOR U10014 ( .A(n11596), .B(n11597), .Z(n8749) );
  NOR U10015 ( .A(n11598), .B(n11596), .Z(n11597) );
  XOR U10016 ( .A(n11599), .B(n11600), .Z(n8752) );
  NOR U10017 ( .A(n11601), .B(n11599), .Z(n11600) );
  XOR U10018 ( .A(n11602), .B(n11603), .Z(n8755) );
  NOR U10019 ( .A(n11604), .B(n11602), .Z(n11603) );
  XOR U10020 ( .A(n11605), .B(n11606), .Z(n8758) );
  NOR U10021 ( .A(n11607), .B(n11605), .Z(n11606) );
  XOR U10022 ( .A(n11608), .B(n11609), .Z(n8761) );
  NOR U10023 ( .A(n11610), .B(n11608), .Z(n11609) );
  XOR U10024 ( .A(n11611), .B(n11612), .Z(n8764) );
  NOR U10025 ( .A(n11613), .B(n11611), .Z(n11612) );
  XOR U10026 ( .A(n11614), .B(n11615), .Z(n8767) );
  NOR U10027 ( .A(n11616), .B(n11614), .Z(n11615) );
  XOR U10028 ( .A(n11617), .B(n11618), .Z(n8770) );
  NOR U10029 ( .A(n11619), .B(n11617), .Z(n11618) );
  XOR U10030 ( .A(n11620), .B(n11621), .Z(n8773) );
  NOR U10031 ( .A(n11622), .B(n11620), .Z(n11621) );
  XOR U10032 ( .A(n11623), .B(n11624), .Z(n8776) );
  NOR U10033 ( .A(n11625), .B(n11623), .Z(n11624) );
  XOR U10034 ( .A(n11626), .B(n11627), .Z(n8779) );
  NOR U10035 ( .A(n11628), .B(n11626), .Z(n11627) );
  XOR U10036 ( .A(n11629), .B(n11630), .Z(n8782) );
  NOR U10037 ( .A(n11631), .B(n11629), .Z(n11630) );
  XOR U10038 ( .A(n11632), .B(n11633), .Z(n8785) );
  NOR U10039 ( .A(n11634), .B(n11632), .Z(n11633) );
  XOR U10040 ( .A(n11635), .B(n11636), .Z(n8788) );
  NOR U10041 ( .A(n11637), .B(n11635), .Z(n11636) );
  XOR U10042 ( .A(n11638), .B(n11639), .Z(n8791) );
  NOR U10043 ( .A(n11640), .B(n11638), .Z(n11639) );
  XOR U10044 ( .A(n11641), .B(n11642), .Z(n8794) );
  NOR U10045 ( .A(n11643), .B(n11641), .Z(n11642) );
  XOR U10046 ( .A(n11644), .B(n11645), .Z(n8797) );
  NOR U10047 ( .A(n11646), .B(n11644), .Z(n11645) );
  XOR U10048 ( .A(n11647), .B(n11648), .Z(n8800) );
  NOR U10049 ( .A(n11649), .B(n11647), .Z(n11648) );
  XOR U10050 ( .A(n11650), .B(n11651), .Z(n8803) );
  NOR U10051 ( .A(n11652), .B(n11650), .Z(n11651) );
  XOR U10052 ( .A(n11653), .B(n11654), .Z(n8806) );
  NOR U10053 ( .A(n11655), .B(n11653), .Z(n11654) );
  XOR U10054 ( .A(n11656), .B(n11657), .Z(n8809) );
  NOR U10055 ( .A(n11658), .B(n11656), .Z(n11657) );
  XOR U10056 ( .A(n11659), .B(n11660), .Z(n8812) );
  NOR U10057 ( .A(n11661), .B(n11659), .Z(n11660) );
  XOR U10058 ( .A(n11662), .B(n11663), .Z(n8815) );
  NOR U10059 ( .A(n11664), .B(n11662), .Z(n11663) );
  XOR U10060 ( .A(n11665), .B(n11666), .Z(n8818) );
  NOR U10061 ( .A(n11667), .B(n11665), .Z(n11666) );
  XOR U10062 ( .A(n11668), .B(n11669), .Z(n8821) );
  NOR U10063 ( .A(n11670), .B(n11668), .Z(n11669) );
  XOR U10064 ( .A(n11671), .B(n11672), .Z(n8824) );
  NOR U10065 ( .A(n11673), .B(n11671), .Z(n11672) );
  XOR U10066 ( .A(n11674), .B(n11675), .Z(n8827) );
  NOR U10067 ( .A(n11676), .B(n11674), .Z(n11675) );
  XOR U10068 ( .A(n11677), .B(n11678), .Z(n8830) );
  NOR U10069 ( .A(n11679), .B(n11677), .Z(n11678) );
  XOR U10070 ( .A(n11680), .B(n11681), .Z(n8833) );
  NOR U10071 ( .A(n11682), .B(n11680), .Z(n11681) );
  XOR U10072 ( .A(n11683), .B(n11684), .Z(n8836) );
  NOR U10073 ( .A(n11685), .B(n11683), .Z(n11684) );
  XOR U10074 ( .A(n11686), .B(n11687), .Z(n8839) );
  NOR U10075 ( .A(n11688), .B(n11686), .Z(n11687) );
  XOR U10076 ( .A(n11689), .B(n11690), .Z(n8842) );
  NOR U10077 ( .A(n11691), .B(n11689), .Z(n11690) );
  XOR U10078 ( .A(n11692), .B(n11693), .Z(n8845) );
  NOR U10079 ( .A(n11694), .B(n11692), .Z(n11693) );
  XOR U10080 ( .A(n11695), .B(n11696), .Z(n8848) );
  NOR U10081 ( .A(n11697), .B(n11695), .Z(n11696) );
  XOR U10082 ( .A(n11698), .B(n11699), .Z(n8851) );
  NOR U10083 ( .A(n11700), .B(n11698), .Z(n11699) );
  XOR U10084 ( .A(n11701), .B(n11702), .Z(n8854) );
  NOR U10085 ( .A(n11703), .B(n11701), .Z(n11702) );
  XOR U10086 ( .A(n11704), .B(n11705), .Z(n8857) );
  NOR U10087 ( .A(n11706), .B(n11704), .Z(n11705) );
  XOR U10088 ( .A(n11707), .B(n11708), .Z(n8860) );
  NOR U10089 ( .A(n11709), .B(n11707), .Z(n11708) );
  XOR U10090 ( .A(n11710), .B(n11711), .Z(n8863) );
  NOR U10091 ( .A(n11712), .B(n11710), .Z(n11711) );
  XOR U10092 ( .A(n11713), .B(n11714), .Z(n8866) );
  NOR U10093 ( .A(n11715), .B(n11713), .Z(n11714) );
  XOR U10094 ( .A(n11716), .B(n11717), .Z(n8869) );
  NOR U10095 ( .A(n11718), .B(n11716), .Z(n11717) );
  XOR U10096 ( .A(n11719), .B(n11720), .Z(n8872) );
  NOR U10097 ( .A(n11721), .B(n11719), .Z(n11720) );
  XOR U10098 ( .A(n11722), .B(n11723), .Z(n8875) );
  NOR U10099 ( .A(n11724), .B(n11722), .Z(n11723) );
  XOR U10100 ( .A(n11725), .B(n11726), .Z(n8878) );
  NOR U10101 ( .A(n11727), .B(n11725), .Z(n11726) );
  XOR U10102 ( .A(n11728), .B(n11729), .Z(n8881) );
  NOR U10103 ( .A(n11730), .B(n11728), .Z(n11729) );
  XOR U10104 ( .A(n11731), .B(n11732), .Z(n8884) );
  NOR U10105 ( .A(n11733), .B(n11731), .Z(n11732) );
  XOR U10106 ( .A(n11734), .B(n11735), .Z(n8887) );
  NOR U10107 ( .A(n11736), .B(n11734), .Z(n11735) );
  XOR U10108 ( .A(n11737), .B(n11738), .Z(n8890) );
  NOR U10109 ( .A(n11739), .B(n11737), .Z(n11738) );
  XOR U10110 ( .A(n11740), .B(n11741), .Z(n8893) );
  NOR U10111 ( .A(n11742), .B(n11740), .Z(n11741) );
  XOR U10112 ( .A(n11743), .B(n11744), .Z(n8896) );
  NOR U10113 ( .A(n11745), .B(n11743), .Z(n11744) );
  XOR U10114 ( .A(n11746), .B(n11747), .Z(n8899) );
  NOR U10115 ( .A(n11748), .B(n11746), .Z(n11747) );
  XOR U10116 ( .A(n11749), .B(n11750), .Z(n8902) );
  NOR U10117 ( .A(n11751), .B(n11749), .Z(n11750) );
  XOR U10118 ( .A(n11752), .B(n11753), .Z(n8905) );
  NOR U10119 ( .A(n11754), .B(n11752), .Z(n11753) );
  XOR U10120 ( .A(n11755), .B(n11756), .Z(n8908) );
  NOR U10121 ( .A(n11757), .B(n11755), .Z(n11756) );
  XOR U10122 ( .A(n11758), .B(n11759), .Z(n8911) );
  NOR U10123 ( .A(n11760), .B(n11758), .Z(n11759) );
  XOR U10124 ( .A(n11761), .B(n11762), .Z(n8914) );
  NOR U10125 ( .A(n11763), .B(n11761), .Z(n11762) );
  XOR U10126 ( .A(n11764), .B(n11765), .Z(n8917) );
  NOR U10127 ( .A(n11766), .B(n11764), .Z(n11765) );
  XOR U10128 ( .A(n11767), .B(n11768), .Z(n8920) );
  NOR U10129 ( .A(n11769), .B(n11767), .Z(n11768) );
  XOR U10130 ( .A(n11770), .B(n11771), .Z(n8923) );
  NOR U10131 ( .A(n11772), .B(n11770), .Z(n11771) );
  XOR U10132 ( .A(n11773), .B(n11774), .Z(n8926) );
  NOR U10133 ( .A(n11775), .B(n11773), .Z(n11774) );
  XOR U10134 ( .A(n11776), .B(n11777), .Z(n8929) );
  NOR U10135 ( .A(n11778), .B(n11776), .Z(n11777) );
  XOR U10136 ( .A(n11779), .B(n11780), .Z(n8932) );
  NOR U10137 ( .A(n11781), .B(n11779), .Z(n11780) );
  XOR U10138 ( .A(n11782), .B(n11783), .Z(n8935) );
  NOR U10139 ( .A(n11784), .B(n11782), .Z(n11783) );
  XOR U10140 ( .A(n11785), .B(n11786), .Z(n8938) );
  NOR U10141 ( .A(n11787), .B(n11785), .Z(n11786) );
  XOR U10142 ( .A(n11788), .B(n11789), .Z(n8941) );
  NOR U10143 ( .A(n11790), .B(n11788), .Z(n11789) );
  XOR U10144 ( .A(n11791), .B(n11792), .Z(n8944) );
  NOR U10145 ( .A(n11793), .B(n11791), .Z(n11792) );
  XOR U10146 ( .A(n11794), .B(n11795), .Z(n8947) );
  NOR U10147 ( .A(n11796), .B(n11794), .Z(n11795) );
  XOR U10148 ( .A(n11797), .B(n11798), .Z(n8950) );
  NOR U10149 ( .A(n11799), .B(n11797), .Z(n11798) );
  XOR U10150 ( .A(n11800), .B(n11801), .Z(n8953) );
  NOR U10151 ( .A(n11802), .B(n11800), .Z(n11801) );
  XOR U10152 ( .A(n11803), .B(n11804), .Z(n8956) );
  NOR U10153 ( .A(n11805), .B(n11803), .Z(n11804) );
  XOR U10154 ( .A(n11806), .B(n11807), .Z(n8959) );
  NOR U10155 ( .A(n11808), .B(n11806), .Z(n11807) );
  XOR U10156 ( .A(n11809), .B(n11810), .Z(n8962) );
  NOR U10157 ( .A(n11811), .B(n11809), .Z(n11810) );
  XOR U10158 ( .A(n11812), .B(n11813), .Z(n8965) );
  NOR U10159 ( .A(n11814), .B(n11812), .Z(n11813) );
  XOR U10160 ( .A(n11815), .B(n11816), .Z(n8968) );
  NOR U10161 ( .A(n11817), .B(n11815), .Z(n11816) );
  XOR U10162 ( .A(n11818), .B(n11819), .Z(n8971) );
  NOR U10163 ( .A(n11820), .B(n11818), .Z(n11819) );
  XOR U10164 ( .A(n11821), .B(n11822), .Z(n8974) );
  NOR U10165 ( .A(n11823), .B(n11821), .Z(n11822) );
  XOR U10166 ( .A(n11824), .B(n11825), .Z(n8977) );
  NOR U10167 ( .A(n11826), .B(n11824), .Z(n11825) );
  XOR U10168 ( .A(n11827), .B(n11828), .Z(n8980) );
  NOR U10169 ( .A(n11829), .B(n11827), .Z(n11828) );
  XOR U10170 ( .A(n11830), .B(n11831), .Z(n8983) );
  NOR U10171 ( .A(n11832), .B(n11830), .Z(n11831) );
  XOR U10172 ( .A(n11833), .B(n11834), .Z(n8986) );
  NOR U10173 ( .A(n11835), .B(n11833), .Z(n11834) );
  XOR U10174 ( .A(n11836), .B(n11837), .Z(n8989) );
  NOR U10175 ( .A(n11838), .B(n11836), .Z(n11837) );
  XOR U10176 ( .A(n11839), .B(n11840), .Z(n8992) );
  NOR U10177 ( .A(n11841), .B(n11839), .Z(n11840) );
  XOR U10178 ( .A(n11842), .B(n11843), .Z(n8995) );
  NOR U10179 ( .A(n11844), .B(n11842), .Z(n11843) );
  XOR U10180 ( .A(n11845), .B(n11846), .Z(n8998) );
  NOR U10181 ( .A(n11847), .B(n11845), .Z(n11846) );
  XOR U10182 ( .A(n11848), .B(n11849), .Z(n9001) );
  NOR U10183 ( .A(n11850), .B(n11848), .Z(n11849) );
  XOR U10184 ( .A(n11851), .B(n11852), .Z(n9004) );
  NOR U10185 ( .A(n11853), .B(n11851), .Z(n11852) );
  XOR U10186 ( .A(n11854), .B(n11855), .Z(n9007) );
  NOR U10187 ( .A(n11856), .B(n11854), .Z(n11855) );
  XOR U10188 ( .A(n11857), .B(n11858), .Z(n9010) );
  NOR U10189 ( .A(n11859), .B(n11857), .Z(n11858) );
  XOR U10190 ( .A(n11860), .B(n11861), .Z(n9013) );
  NOR U10191 ( .A(n11862), .B(n11860), .Z(n11861) );
  XOR U10192 ( .A(n11863), .B(n11864), .Z(n9016) );
  NOR U10193 ( .A(n11865), .B(n11863), .Z(n11864) );
  XOR U10194 ( .A(n11866), .B(n11867), .Z(n9019) );
  NOR U10195 ( .A(n11868), .B(n11866), .Z(n11867) );
  XOR U10196 ( .A(n11869), .B(n11870), .Z(n9022) );
  NOR U10197 ( .A(n11871), .B(n11869), .Z(n11870) );
  XOR U10198 ( .A(n11872), .B(n11873), .Z(n9025) );
  NOR U10199 ( .A(n11874), .B(n11872), .Z(n11873) );
  XOR U10200 ( .A(n11875), .B(n11876), .Z(n9028) );
  NOR U10201 ( .A(n11877), .B(n11875), .Z(n11876) );
  XOR U10202 ( .A(n11878), .B(n11879), .Z(n9031) );
  NOR U10203 ( .A(n11880), .B(n11878), .Z(n11879) );
  XOR U10204 ( .A(n11881), .B(n11882), .Z(n9034) );
  NOR U10205 ( .A(n11883), .B(n11881), .Z(n11882) );
  XOR U10206 ( .A(n11884), .B(n11885), .Z(n9037) );
  NOR U10207 ( .A(n11886), .B(n11884), .Z(n11885) );
  XOR U10208 ( .A(n11887), .B(n11888), .Z(n9040) );
  NOR U10209 ( .A(n11889), .B(n11887), .Z(n11888) );
  XOR U10210 ( .A(n11890), .B(n11891), .Z(n9043) );
  NOR U10211 ( .A(n11892), .B(n11890), .Z(n11891) );
  XOR U10212 ( .A(n11893), .B(n11894), .Z(n9046) );
  NOR U10213 ( .A(n11895), .B(n11893), .Z(n11894) );
  XOR U10214 ( .A(n11896), .B(n11897), .Z(n9049) );
  NOR U10215 ( .A(n11898), .B(n11896), .Z(n11897) );
  XOR U10216 ( .A(n11899), .B(n11900), .Z(n9052) );
  NOR U10217 ( .A(n11901), .B(n11899), .Z(n11900) );
  XOR U10218 ( .A(n11902), .B(n11903), .Z(n9055) );
  NOR U10219 ( .A(n11904), .B(n11902), .Z(n11903) );
  XOR U10220 ( .A(n11905), .B(n11906), .Z(n9058) );
  NOR U10221 ( .A(n11907), .B(n11905), .Z(n11906) );
  XOR U10222 ( .A(n11908), .B(n11909), .Z(n9061) );
  NOR U10223 ( .A(n11910), .B(n11908), .Z(n11909) );
  XOR U10224 ( .A(n11911), .B(n11912), .Z(n9064) );
  NOR U10225 ( .A(n11913), .B(n11911), .Z(n11912) );
  XOR U10226 ( .A(n11914), .B(n11915), .Z(n9067) );
  NOR U10227 ( .A(n11916), .B(n11914), .Z(n11915) );
  XOR U10228 ( .A(n11917), .B(n11918), .Z(n9070) );
  NOR U10229 ( .A(n11919), .B(n11917), .Z(n11918) );
  XOR U10230 ( .A(n11920), .B(n11921), .Z(n9073) );
  NOR U10231 ( .A(n11922), .B(n11920), .Z(n11921) );
  XOR U10232 ( .A(n11923), .B(n11924), .Z(n9076) );
  NOR U10233 ( .A(n11925), .B(n11923), .Z(n11924) );
  XOR U10234 ( .A(n11926), .B(n11927), .Z(n9079) );
  NOR U10235 ( .A(n11928), .B(n11926), .Z(n11927) );
  XOR U10236 ( .A(n11929), .B(n11930), .Z(n9082) );
  NOR U10237 ( .A(n11931), .B(n11929), .Z(n11930) );
  XOR U10238 ( .A(n11932), .B(n11933), .Z(n9085) );
  NOR U10239 ( .A(n11934), .B(n11932), .Z(n11933) );
  XOR U10240 ( .A(n11935), .B(n11936), .Z(n9088) );
  NOR U10241 ( .A(n11937), .B(n11935), .Z(n11936) );
  XOR U10242 ( .A(n11938), .B(n11939), .Z(n9091) );
  NOR U10243 ( .A(n11940), .B(n11938), .Z(n11939) );
  XOR U10244 ( .A(n11941), .B(n11942), .Z(n9094) );
  NOR U10245 ( .A(n11943), .B(n11941), .Z(n11942) );
  XOR U10246 ( .A(n11944), .B(n11945), .Z(n9097) );
  NOR U10247 ( .A(n11946), .B(n11944), .Z(n11945) );
  XOR U10248 ( .A(n11947), .B(n11948), .Z(n9100) );
  NOR U10249 ( .A(n11949), .B(n11947), .Z(n11948) );
  XOR U10250 ( .A(n11950), .B(n11951), .Z(n9103) );
  NOR U10251 ( .A(n11952), .B(n11950), .Z(n11951) );
  XOR U10252 ( .A(n11953), .B(n11954), .Z(n9106) );
  NOR U10253 ( .A(n11955), .B(n11953), .Z(n11954) );
  XOR U10254 ( .A(n11956), .B(n11957), .Z(n9109) );
  NOR U10255 ( .A(n11958), .B(n11956), .Z(n11957) );
  XOR U10256 ( .A(n11959), .B(n11960), .Z(n9112) );
  NOR U10257 ( .A(n11961), .B(n11959), .Z(n11960) );
  XOR U10258 ( .A(n11962), .B(n11963), .Z(n9115) );
  NOR U10259 ( .A(n11964), .B(n11962), .Z(n11963) );
  XOR U10260 ( .A(n11965), .B(n11966), .Z(n9118) );
  NOR U10261 ( .A(n11967), .B(n11965), .Z(n11966) );
  XOR U10262 ( .A(n11968), .B(n11969), .Z(n9121) );
  NOR U10263 ( .A(n11970), .B(n11968), .Z(n11969) );
  XOR U10264 ( .A(n11971), .B(n11972), .Z(n9124) );
  NOR U10265 ( .A(n11973), .B(n11971), .Z(n11972) );
  XOR U10266 ( .A(n11974), .B(n11975), .Z(n9127) );
  NOR U10267 ( .A(n11976), .B(n11974), .Z(n11975) );
  XOR U10268 ( .A(n11977), .B(n11978), .Z(n9130) );
  NOR U10269 ( .A(n11979), .B(n11977), .Z(n11978) );
  XOR U10270 ( .A(n11980), .B(n11981), .Z(n9133) );
  NOR U10271 ( .A(n11982), .B(n11980), .Z(n11981) );
  XOR U10272 ( .A(n11983), .B(n11984), .Z(n9136) );
  NOR U10273 ( .A(n11985), .B(n11983), .Z(n11984) );
  XOR U10274 ( .A(n11986), .B(n11987), .Z(n9139) );
  NOR U10275 ( .A(n11988), .B(n11986), .Z(n11987) );
  XOR U10276 ( .A(n11989), .B(n11990), .Z(n9142) );
  NOR U10277 ( .A(n11991), .B(n11989), .Z(n11990) );
  XOR U10278 ( .A(n11992), .B(n11993), .Z(n9145) );
  NOR U10279 ( .A(n11994), .B(n11992), .Z(n11993) );
  XOR U10280 ( .A(n11995), .B(n11996), .Z(n9148) );
  NOR U10281 ( .A(n11997), .B(n11995), .Z(n11996) );
  XOR U10282 ( .A(n11998), .B(n11999), .Z(n9151) );
  NOR U10283 ( .A(n12000), .B(n11998), .Z(n11999) );
  XOR U10284 ( .A(n12001), .B(n12002), .Z(n9154) );
  NOR U10285 ( .A(n12003), .B(n12001), .Z(n12002) );
  XOR U10286 ( .A(n12004), .B(n12005), .Z(n9157) );
  NOR U10287 ( .A(n12006), .B(n12004), .Z(n12005) );
  XOR U10288 ( .A(n12007), .B(n12008), .Z(n9160) );
  NOR U10289 ( .A(n12009), .B(n12007), .Z(n12008) );
  XOR U10290 ( .A(n12010), .B(n12011), .Z(n9163) );
  NOR U10291 ( .A(n12012), .B(n12010), .Z(n12011) );
  XOR U10292 ( .A(n12013), .B(n12014), .Z(n9166) );
  NOR U10293 ( .A(n12015), .B(n12013), .Z(n12014) );
  XOR U10294 ( .A(n12016), .B(n12017), .Z(n9169) );
  NOR U10295 ( .A(n12018), .B(n12016), .Z(n12017) );
  XOR U10296 ( .A(n12019), .B(n12020), .Z(n9172) );
  NOR U10297 ( .A(n12021), .B(n12019), .Z(n12020) );
  XOR U10298 ( .A(n12022), .B(n12023), .Z(n9175) );
  NOR U10299 ( .A(n12024), .B(n12022), .Z(n12023) );
  XOR U10300 ( .A(n12025), .B(n12026), .Z(n9178) );
  NOR U10301 ( .A(n12027), .B(n12025), .Z(n12026) );
  XOR U10302 ( .A(n12028), .B(n12029), .Z(n9181) );
  NOR U10303 ( .A(n12030), .B(n12028), .Z(n12029) );
  XOR U10304 ( .A(n12031), .B(n12032), .Z(n9184) );
  NOR U10305 ( .A(n12033), .B(n12031), .Z(n12032) );
  XOR U10306 ( .A(n12034), .B(n12035), .Z(n9187) );
  NOR U10307 ( .A(n12036), .B(n12034), .Z(n12035) );
  XOR U10308 ( .A(n12037), .B(n12038), .Z(n9190) );
  NOR U10309 ( .A(n12039), .B(n12037), .Z(n12038) );
  XOR U10310 ( .A(n12040), .B(n12041), .Z(n9193) );
  NOR U10311 ( .A(n12042), .B(n12040), .Z(n12041) );
  XOR U10312 ( .A(n12043), .B(n12044), .Z(n9196) );
  NOR U10313 ( .A(n12045), .B(n12043), .Z(n12044) );
  XOR U10314 ( .A(n12046), .B(n12047), .Z(n9199) );
  NOR U10315 ( .A(n12048), .B(n12046), .Z(n12047) );
  XOR U10316 ( .A(n12049), .B(n12050), .Z(n9202) );
  NOR U10317 ( .A(n12051), .B(n12049), .Z(n12050) );
  XOR U10318 ( .A(n12052), .B(n12053), .Z(n9205) );
  NOR U10319 ( .A(n12054), .B(n12052), .Z(n12053) );
  XOR U10320 ( .A(n12055), .B(n12056), .Z(n9208) );
  NOR U10321 ( .A(n12057), .B(n12055), .Z(n12056) );
  XOR U10322 ( .A(n12058), .B(n12059), .Z(n9211) );
  NOR U10323 ( .A(n12060), .B(n12058), .Z(n12059) );
  XOR U10324 ( .A(n12061), .B(n12062), .Z(n9214) );
  NOR U10325 ( .A(n12063), .B(n12061), .Z(n12062) );
  XOR U10326 ( .A(n12064), .B(n12065), .Z(n9217) );
  NOR U10327 ( .A(n12066), .B(n12064), .Z(n12065) );
  XOR U10328 ( .A(n12067), .B(n12068), .Z(n9220) );
  NOR U10329 ( .A(n12069), .B(n12067), .Z(n12068) );
  XOR U10330 ( .A(n12070), .B(n12071), .Z(n9223) );
  NOR U10331 ( .A(n12072), .B(n12070), .Z(n12071) );
  XOR U10332 ( .A(n12073), .B(n12074), .Z(n9226) );
  NOR U10333 ( .A(n12075), .B(n12073), .Z(n12074) );
  XOR U10334 ( .A(n12076), .B(n12077), .Z(n9229) );
  NOR U10335 ( .A(n12078), .B(n12076), .Z(n12077) );
  XOR U10336 ( .A(n12079), .B(n12080), .Z(n9232) );
  NOR U10337 ( .A(n12081), .B(n12079), .Z(n12080) );
  XOR U10338 ( .A(n12082), .B(n12083), .Z(n9235) );
  NOR U10339 ( .A(n12084), .B(n12082), .Z(n12083) );
  XOR U10340 ( .A(n12085), .B(n12086), .Z(n9238) );
  NOR U10341 ( .A(n12087), .B(n12085), .Z(n12086) );
  XOR U10342 ( .A(n12088), .B(n12089), .Z(n9241) );
  NOR U10343 ( .A(n12090), .B(n12088), .Z(n12089) );
  XOR U10344 ( .A(n12091), .B(n12092), .Z(n9244) );
  NOR U10345 ( .A(n12093), .B(n12091), .Z(n12092) );
  XOR U10346 ( .A(n12094), .B(n12095), .Z(n9247) );
  NOR U10347 ( .A(n12096), .B(n12094), .Z(n12095) );
  XOR U10348 ( .A(n12097), .B(n12098), .Z(n9250) );
  NOR U10349 ( .A(n12099), .B(n12097), .Z(n12098) );
  XOR U10350 ( .A(n12100), .B(n12101), .Z(n9253) );
  NOR U10351 ( .A(n12102), .B(n12100), .Z(n12101) );
  XOR U10352 ( .A(n12103), .B(n12104), .Z(n9256) );
  NOR U10353 ( .A(n12105), .B(n12103), .Z(n12104) );
  XOR U10354 ( .A(n12106), .B(n12107), .Z(n9259) );
  NOR U10355 ( .A(n12108), .B(n12106), .Z(n12107) );
  XOR U10356 ( .A(n12109), .B(n12110), .Z(n9262) );
  NOR U10357 ( .A(n12111), .B(n12109), .Z(n12110) );
  XOR U10358 ( .A(n12112), .B(n12113), .Z(n9265) );
  NOR U10359 ( .A(n12114), .B(n12112), .Z(n12113) );
  XOR U10360 ( .A(n12115), .B(n12116), .Z(n9268) );
  NOR U10361 ( .A(n12117), .B(n12115), .Z(n12116) );
  XOR U10362 ( .A(n12118), .B(n12119), .Z(n9271) );
  NOR U10363 ( .A(n12120), .B(n12118), .Z(n12119) );
  XOR U10364 ( .A(n12121), .B(n12122), .Z(n9274) );
  NOR U10365 ( .A(n12123), .B(n12121), .Z(n12122) );
  XOR U10366 ( .A(n12124), .B(n12125), .Z(n9277) );
  NOR U10367 ( .A(n12126), .B(n12124), .Z(n12125) );
  XOR U10368 ( .A(n12127), .B(n12128), .Z(n9280) );
  NOR U10369 ( .A(n12129), .B(n12127), .Z(n12128) );
  XOR U10370 ( .A(n12130), .B(n12131), .Z(n9283) );
  NOR U10371 ( .A(n12132), .B(n12130), .Z(n12131) );
  XOR U10372 ( .A(n12133), .B(n12134), .Z(n9286) );
  NOR U10373 ( .A(n12135), .B(n12133), .Z(n12134) );
  XOR U10374 ( .A(n12136), .B(n12137), .Z(n9289) );
  NOR U10375 ( .A(n12138), .B(n12136), .Z(n12137) );
  XOR U10376 ( .A(n12139), .B(n12140), .Z(n9292) );
  NOR U10377 ( .A(n12141), .B(n12139), .Z(n12140) );
  XOR U10378 ( .A(n12142), .B(n12143), .Z(n9295) );
  NOR U10379 ( .A(n12144), .B(n12142), .Z(n12143) );
  XOR U10380 ( .A(n12145), .B(n12146), .Z(n9298) );
  NOR U10381 ( .A(n12147), .B(n12145), .Z(n12146) );
  XOR U10382 ( .A(n12148), .B(n12149), .Z(n9301) );
  NOR U10383 ( .A(n12150), .B(n12148), .Z(n12149) );
  XOR U10384 ( .A(n12151), .B(n12152), .Z(n9304) );
  NOR U10385 ( .A(n12153), .B(n12151), .Z(n12152) );
  XOR U10386 ( .A(n12154), .B(n12155), .Z(n9307) );
  NOR U10387 ( .A(n12156), .B(n12154), .Z(n12155) );
  XOR U10388 ( .A(n12157), .B(n12158), .Z(n9310) );
  NOR U10389 ( .A(n12159), .B(n12157), .Z(n12158) );
  XOR U10390 ( .A(n12160), .B(n12161), .Z(n9313) );
  NOR U10391 ( .A(n12162), .B(n12160), .Z(n12161) );
  XOR U10392 ( .A(n12163), .B(n12164), .Z(n9316) );
  NOR U10393 ( .A(n12165), .B(n12163), .Z(n12164) );
  XOR U10394 ( .A(n12166), .B(n12167), .Z(n9319) );
  NOR U10395 ( .A(n12168), .B(n12166), .Z(n12167) );
  XOR U10396 ( .A(n12169), .B(n12170), .Z(n9322) );
  NOR U10397 ( .A(n12171), .B(n12169), .Z(n12170) );
  XOR U10398 ( .A(n12172), .B(n12173), .Z(n9325) );
  NOR U10399 ( .A(n12174), .B(n12172), .Z(n12173) );
  XOR U10400 ( .A(n12175), .B(n12176), .Z(n9328) );
  NOR U10401 ( .A(n12177), .B(n12175), .Z(n12176) );
  XOR U10402 ( .A(n12178), .B(n12179), .Z(n9331) );
  NOR U10403 ( .A(n12180), .B(n12178), .Z(n12179) );
  XOR U10404 ( .A(n12181), .B(n12182), .Z(n9334) );
  NOR U10405 ( .A(n12183), .B(n12181), .Z(n12182) );
  XOR U10406 ( .A(n12184), .B(n12185), .Z(n9337) );
  NOR U10407 ( .A(n12186), .B(n12184), .Z(n12185) );
  XOR U10408 ( .A(n12187), .B(n12188), .Z(n9340) );
  NOR U10409 ( .A(n12189), .B(n12187), .Z(n12188) );
  XOR U10410 ( .A(n12190), .B(n12191), .Z(n9343) );
  NOR U10411 ( .A(n12192), .B(n12190), .Z(n12191) );
  XOR U10412 ( .A(n12193), .B(n12194), .Z(n9346) );
  NOR U10413 ( .A(n12195), .B(n12193), .Z(n12194) );
  XOR U10414 ( .A(n12196), .B(n12197), .Z(n9349) );
  NOR U10415 ( .A(n12198), .B(n12196), .Z(n12197) );
  XOR U10416 ( .A(n12199), .B(n12200), .Z(n9352) );
  NOR U10417 ( .A(n12201), .B(n12199), .Z(n12200) );
  XOR U10418 ( .A(n12202), .B(n12203), .Z(n9355) );
  NOR U10419 ( .A(n12204), .B(n12202), .Z(n12203) );
  XOR U10420 ( .A(n12205), .B(n12206), .Z(n9358) );
  NOR U10421 ( .A(n12207), .B(n12205), .Z(n12206) );
  XOR U10422 ( .A(n12208), .B(n12209), .Z(n9361) );
  NOR U10423 ( .A(n12210), .B(n12208), .Z(n12209) );
  XOR U10424 ( .A(n12211), .B(n12212), .Z(n9364) );
  NOR U10425 ( .A(n12213), .B(n12211), .Z(n12212) );
  XOR U10426 ( .A(n12214), .B(n12215), .Z(n9367) );
  NOR U10427 ( .A(n12216), .B(n12214), .Z(n12215) );
  XOR U10428 ( .A(n12217), .B(n12218), .Z(n9370) );
  NOR U10429 ( .A(n12219), .B(n12217), .Z(n12218) );
  XOR U10430 ( .A(n12220), .B(n12221), .Z(n9373) );
  NOR U10431 ( .A(n12222), .B(n12220), .Z(n12221) );
  XOR U10432 ( .A(n12223), .B(n12224), .Z(n9376) );
  NOR U10433 ( .A(n12225), .B(n12223), .Z(n12224) );
  XOR U10434 ( .A(n12226), .B(n12227), .Z(n9379) );
  NOR U10435 ( .A(n12228), .B(n12226), .Z(n12227) );
  XOR U10436 ( .A(n12229), .B(n12230), .Z(n9382) );
  NOR U10437 ( .A(n12231), .B(n12229), .Z(n12230) );
  XOR U10438 ( .A(n12232), .B(n12233), .Z(n9385) );
  NOR U10439 ( .A(n12234), .B(n12232), .Z(n12233) );
  XOR U10440 ( .A(n12235), .B(n12236), .Z(n9388) );
  NOR U10441 ( .A(n12237), .B(n12235), .Z(n12236) );
  XOR U10442 ( .A(n12238), .B(n12239), .Z(n9391) );
  NOR U10443 ( .A(n12240), .B(n12238), .Z(n12239) );
  XOR U10444 ( .A(n12241), .B(n12242), .Z(n9394) );
  NOR U10445 ( .A(n12243), .B(n12241), .Z(n12242) );
  XOR U10446 ( .A(n12244), .B(n12245), .Z(n9397) );
  NOR U10447 ( .A(n12246), .B(n12244), .Z(n12245) );
  XOR U10448 ( .A(n12247), .B(n12248), .Z(n9400) );
  NOR U10449 ( .A(n12249), .B(n12247), .Z(n12248) );
  XOR U10450 ( .A(n12250), .B(n12251), .Z(n9403) );
  NOR U10451 ( .A(n12252), .B(n12250), .Z(n12251) );
  XOR U10452 ( .A(n12253), .B(n12254), .Z(n9406) );
  NOR U10453 ( .A(n12255), .B(n12253), .Z(n12254) );
  XOR U10454 ( .A(n12256), .B(n12257), .Z(n9409) );
  NOR U10455 ( .A(n12258), .B(n12256), .Z(n12257) );
  XOR U10456 ( .A(n12259), .B(n12260), .Z(n9412) );
  NOR U10457 ( .A(n12261), .B(n12259), .Z(n12260) );
  XOR U10458 ( .A(n12262), .B(n12263), .Z(n9415) );
  NOR U10459 ( .A(n12264), .B(n12262), .Z(n12263) );
  XOR U10460 ( .A(n12265), .B(n12266), .Z(n9418) );
  NOR U10461 ( .A(n12267), .B(n12265), .Z(n12266) );
  XOR U10462 ( .A(n12268), .B(n12269), .Z(n9421) );
  NOR U10463 ( .A(n12270), .B(n12268), .Z(n12269) );
  XOR U10464 ( .A(n12271), .B(n12272), .Z(n9424) );
  NOR U10465 ( .A(n12273), .B(n12271), .Z(n12272) );
  XOR U10466 ( .A(n12274), .B(n12275), .Z(n9427) );
  NOR U10467 ( .A(n12276), .B(n12274), .Z(n12275) );
  XOR U10468 ( .A(n12277), .B(n12278), .Z(n9430) );
  NOR U10469 ( .A(n12279), .B(n12277), .Z(n12278) );
  XOR U10470 ( .A(n12280), .B(n12281), .Z(n9433) );
  NOR U10471 ( .A(n12282), .B(n12280), .Z(n12281) );
  XOR U10472 ( .A(n12283), .B(n12284), .Z(n9436) );
  NOR U10473 ( .A(n12285), .B(n12283), .Z(n12284) );
  XOR U10474 ( .A(n12286), .B(n12287), .Z(n9439) );
  NOR U10475 ( .A(n12288), .B(n12286), .Z(n12287) );
  XOR U10476 ( .A(n12289), .B(n12290), .Z(n9442) );
  NOR U10477 ( .A(n12291), .B(n12289), .Z(n12290) );
  XOR U10478 ( .A(n12292), .B(n12293), .Z(n9445) );
  NOR U10479 ( .A(n12294), .B(n12292), .Z(n12293) );
  XOR U10480 ( .A(n12295), .B(n12296), .Z(n9448) );
  NOR U10481 ( .A(n12297), .B(n12295), .Z(n12296) );
  XOR U10482 ( .A(n12298), .B(n12299), .Z(n9451) );
  NOR U10483 ( .A(n12300), .B(n12298), .Z(n12299) );
  XOR U10484 ( .A(n12301), .B(n12302), .Z(n9454) );
  NOR U10485 ( .A(n12303), .B(n12301), .Z(n12302) );
  XOR U10486 ( .A(n12304), .B(n12305), .Z(n9457) );
  NOR U10487 ( .A(n12306), .B(n12304), .Z(n12305) );
  XOR U10488 ( .A(n12307), .B(n12308), .Z(n9460) );
  NOR U10489 ( .A(n12309), .B(n12307), .Z(n12308) );
  XOR U10490 ( .A(n12310), .B(n12311), .Z(n9463) );
  NOR U10491 ( .A(n12312), .B(n12310), .Z(n12311) );
  XOR U10492 ( .A(n12313), .B(n12314), .Z(n9466) );
  NOR U10493 ( .A(n12315), .B(n12313), .Z(n12314) );
  XOR U10494 ( .A(n12316), .B(n12317), .Z(n9469) );
  NOR U10495 ( .A(n12318), .B(n12316), .Z(n12317) );
  XOR U10496 ( .A(n12319), .B(n12320), .Z(n9472) );
  NOR U10497 ( .A(n12321), .B(n12319), .Z(n12320) );
  XOR U10498 ( .A(n12322), .B(n12323), .Z(n9475) );
  NOR U10499 ( .A(n12324), .B(n12322), .Z(n12323) );
  XOR U10500 ( .A(n12325), .B(n12326), .Z(n9478) );
  NOR U10501 ( .A(n12327), .B(n12325), .Z(n12326) );
  XOR U10502 ( .A(n12328), .B(n12329), .Z(n9481) );
  NOR U10503 ( .A(n12330), .B(n12328), .Z(n12329) );
  XOR U10504 ( .A(n12331), .B(n12332), .Z(n9484) );
  NOR U10505 ( .A(n12333), .B(n12331), .Z(n12332) );
  XOR U10506 ( .A(n12334), .B(n12335), .Z(n9487) );
  NOR U10507 ( .A(n12336), .B(n12334), .Z(n12335) );
  XOR U10508 ( .A(n12337), .B(n12338), .Z(n9490) );
  NOR U10509 ( .A(n12339), .B(n12337), .Z(n12338) );
  XOR U10510 ( .A(n12340), .B(n12341), .Z(n9493) );
  NOR U10511 ( .A(n12342), .B(n12340), .Z(n12341) );
  XOR U10512 ( .A(n12343), .B(n12344), .Z(n9496) );
  NOR U10513 ( .A(n12345), .B(n12343), .Z(n12344) );
  XOR U10514 ( .A(n12346), .B(n12347), .Z(n9499) );
  NOR U10515 ( .A(n12348), .B(n12346), .Z(n12347) );
  XOR U10516 ( .A(n12349), .B(n12350), .Z(n9502) );
  NOR U10517 ( .A(n12351), .B(n12349), .Z(n12350) );
  XOR U10518 ( .A(n12352), .B(n12353), .Z(n9505) );
  NOR U10519 ( .A(n12354), .B(n12352), .Z(n12353) );
  XOR U10520 ( .A(n12355), .B(n12356), .Z(n9508) );
  NOR U10521 ( .A(n12357), .B(n12355), .Z(n12356) );
  XOR U10522 ( .A(n12358), .B(n12359), .Z(n9511) );
  NOR U10523 ( .A(n12360), .B(n12358), .Z(n12359) );
  XOR U10524 ( .A(n12361), .B(n12362), .Z(n9514) );
  NOR U10525 ( .A(n12363), .B(n12361), .Z(n12362) );
  XOR U10526 ( .A(n12364), .B(n12365), .Z(n9517) );
  NOR U10527 ( .A(n12366), .B(n12364), .Z(n12365) );
  XOR U10528 ( .A(n12367), .B(n12368), .Z(n9520) );
  NOR U10529 ( .A(n12369), .B(n12367), .Z(n12368) );
  XOR U10530 ( .A(n12370), .B(n12371), .Z(n9523) );
  NOR U10531 ( .A(n12372), .B(n12370), .Z(n12371) );
  XOR U10532 ( .A(n12373), .B(n12374), .Z(n9526) );
  NOR U10533 ( .A(n12375), .B(n12373), .Z(n12374) );
  XOR U10534 ( .A(n12376), .B(n12377), .Z(n9529) );
  NOR U10535 ( .A(n12378), .B(n12376), .Z(n12377) );
  XOR U10536 ( .A(n12379), .B(n12380), .Z(n9532) );
  NOR U10537 ( .A(n12381), .B(n12379), .Z(n12380) );
  XOR U10538 ( .A(n12382), .B(n12383), .Z(n9535) );
  NOR U10539 ( .A(n12384), .B(n12382), .Z(n12383) );
  XOR U10540 ( .A(n12385), .B(n12386), .Z(n9538) );
  NOR U10541 ( .A(n12387), .B(n12385), .Z(n12386) );
  XOR U10542 ( .A(n12388), .B(n12389), .Z(n9541) );
  NOR U10543 ( .A(n12390), .B(n12388), .Z(n12389) );
  XOR U10544 ( .A(n12391), .B(n12392), .Z(n9544) );
  NOR U10545 ( .A(n12393), .B(n12391), .Z(n12392) );
  XOR U10546 ( .A(n12394), .B(n12395), .Z(n9547) );
  NOR U10547 ( .A(n12396), .B(n12394), .Z(n12395) );
  XOR U10548 ( .A(n12397), .B(n12398), .Z(n9550) );
  NOR U10549 ( .A(n12399), .B(n12397), .Z(n12398) );
  XOR U10550 ( .A(n12400), .B(n12401), .Z(n9553) );
  NOR U10551 ( .A(n12402), .B(n12400), .Z(n12401) );
  XOR U10552 ( .A(n12403), .B(n12404), .Z(n9556) );
  NOR U10553 ( .A(n12405), .B(n12403), .Z(n12404) );
  XOR U10554 ( .A(n12406), .B(n12407), .Z(n9559) );
  NOR U10555 ( .A(n12408), .B(n12406), .Z(n12407) );
  XOR U10556 ( .A(n12409), .B(n12410), .Z(n9562) );
  NOR U10557 ( .A(n12411), .B(n12409), .Z(n12410) );
  XOR U10558 ( .A(n12412), .B(n12413), .Z(n9565) );
  NOR U10559 ( .A(n12414), .B(n12412), .Z(n12413) );
  XOR U10560 ( .A(n12415), .B(n12416), .Z(n9568) );
  NOR U10561 ( .A(n12417), .B(n12415), .Z(n12416) );
  XOR U10562 ( .A(n12418), .B(n12419), .Z(n9571) );
  NOR U10563 ( .A(n12420), .B(n12418), .Z(n12419) );
  XOR U10564 ( .A(n12421), .B(n12422), .Z(n9574) );
  NOR U10565 ( .A(n12423), .B(n12421), .Z(n12422) );
  XOR U10566 ( .A(n12424), .B(n12425), .Z(n9577) );
  NOR U10567 ( .A(n12426), .B(n12424), .Z(n12425) );
  XOR U10568 ( .A(n12427), .B(n12428), .Z(n9580) );
  NOR U10569 ( .A(n12429), .B(n12427), .Z(n12428) );
  XOR U10570 ( .A(n12430), .B(n12431), .Z(n9583) );
  NOR U10571 ( .A(n12432), .B(n12430), .Z(n12431) );
  XOR U10572 ( .A(n12433), .B(n12434), .Z(n9586) );
  NOR U10573 ( .A(n12435), .B(n12433), .Z(n12434) );
  XOR U10574 ( .A(n12436), .B(n12437), .Z(n9589) );
  NOR U10575 ( .A(n12438), .B(n12436), .Z(n12437) );
  XOR U10576 ( .A(n12439), .B(n12440), .Z(n9592) );
  NOR U10577 ( .A(n12441), .B(n12439), .Z(n12440) );
  XOR U10578 ( .A(n12442), .B(n12443), .Z(n9595) );
  NOR U10579 ( .A(n12444), .B(n12442), .Z(n12443) );
  XOR U10580 ( .A(n12445), .B(n12446), .Z(n9598) );
  NOR U10581 ( .A(n12447), .B(n12445), .Z(n12446) );
  XOR U10582 ( .A(n12448), .B(n12449), .Z(n9601) );
  NOR U10583 ( .A(n12450), .B(n12448), .Z(n12449) );
  XOR U10584 ( .A(n12451), .B(n12452), .Z(n9604) );
  NOR U10585 ( .A(n12453), .B(n12451), .Z(n12452) );
  XOR U10586 ( .A(n12454), .B(n12455), .Z(n9607) );
  NOR U10587 ( .A(n12456), .B(n12454), .Z(n12455) );
  XOR U10588 ( .A(n12457), .B(n12458), .Z(n9610) );
  NOR U10589 ( .A(n12459), .B(n12457), .Z(n12458) );
  XOR U10590 ( .A(n12460), .B(n12461), .Z(n9613) );
  NOR U10591 ( .A(n12462), .B(n12460), .Z(n12461) );
  XOR U10592 ( .A(n12463), .B(n12464), .Z(n9616) );
  NOR U10593 ( .A(n12465), .B(n12463), .Z(n12464) );
  XOR U10594 ( .A(n12466), .B(n12467), .Z(n9619) );
  NOR U10595 ( .A(n12468), .B(n12466), .Z(n12467) );
  XOR U10596 ( .A(n12469), .B(n12470), .Z(n9622) );
  NOR U10597 ( .A(n12471), .B(n12469), .Z(n12470) );
  XOR U10598 ( .A(n12472), .B(n12473), .Z(n9625) );
  NOR U10599 ( .A(n12474), .B(n12472), .Z(n12473) );
  XOR U10600 ( .A(n12475), .B(n12476), .Z(n9628) );
  NOR U10601 ( .A(n12477), .B(n12475), .Z(n12476) );
  XOR U10602 ( .A(n12478), .B(n12479), .Z(n9631) );
  NOR U10603 ( .A(n12480), .B(n12478), .Z(n12479) );
  XOR U10604 ( .A(n12481), .B(n12482), .Z(n9634) );
  NOR U10605 ( .A(n12483), .B(n12481), .Z(n12482) );
  XOR U10606 ( .A(n12484), .B(n12485), .Z(n9637) );
  NOR U10607 ( .A(n12486), .B(n12484), .Z(n12485) );
  XOR U10608 ( .A(n12487), .B(n12488), .Z(n9640) );
  NOR U10609 ( .A(n12489), .B(n12487), .Z(n12488) );
  XOR U10610 ( .A(n12490), .B(n12491), .Z(n9643) );
  NOR U10611 ( .A(n12492), .B(n12490), .Z(n12491) );
  XOR U10612 ( .A(n12493), .B(n12494), .Z(n9646) );
  NOR U10613 ( .A(n12495), .B(n12493), .Z(n12494) );
  XOR U10614 ( .A(n12496), .B(n12497), .Z(n9649) );
  NOR U10615 ( .A(n12498), .B(n12496), .Z(n12497) );
  XOR U10616 ( .A(n12499), .B(n12500), .Z(n9652) );
  NOR U10617 ( .A(n12501), .B(n12499), .Z(n12500) );
  XOR U10618 ( .A(n12502), .B(n12503), .Z(n9655) );
  NOR U10619 ( .A(n12504), .B(n12502), .Z(n12503) );
  XOR U10620 ( .A(n12505), .B(n12506), .Z(n9658) );
  NOR U10621 ( .A(n12507), .B(n12505), .Z(n12506) );
  XOR U10622 ( .A(n12508), .B(n12509), .Z(n9661) );
  NOR U10623 ( .A(n12510), .B(n12508), .Z(n12509) );
  XOR U10624 ( .A(n12511), .B(n12512), .Z(n9664) );
  NOR U10625 ( .A(n12513), .B(n12511), .Z(n12512) );
  XOR U10626 ( .A(n12514), .B(n12515), .Z(n9667) );
  NOR U10627 ( .A(n12516), .B(n12514), .Z(n12515) );
  XOR U10628 ( .A(n12517), .B(n12518), .Z(n9670) );
  NOR U10629 ( .A(n12519), .B(n12517), .Z(n12518) );
  XOR U10630 ( .A(n12520), .B(n12521), .Z(n9673) );
  NOR U10631 ( .A(n12522), .B(n12520), .Z(n12521) );
  XOR U10632 ( .A(n12523), .B(n12524), .Z(n9676) );
  NOR U10633 ( .A(n12525), .B(n12523), .Z(n12524) );
  XOR U10634 ( .A(n12526), .B(n12527), .Z(n9679) );
  NOR U10635 ( .A(n12528), .B(n12526), .Z(n12527) );
  XOR U10636 ( .A(n12529), .B(n12530), .Z(n9682) );
  NOR U10637 ( .A(n12531), .B(n12529), .Z(n12530) );
  XOR U10638 ( .A(n12532), .B(n12533), .Z(n9685) );
  NOR U10639 ( .A(n12534), .B(n12532), .Z(n12533) );
  XOR U10640 ( .A(n12535), .B(n12536), .Z(n9688) );
  NOR U10641 ( .A(n12537), .B(n12535), .Z(n12536) );
  XOR U10642 ( .A(n12538), .B(n12539), .Z(n9691) );
  NOR U10643 ( .A(n12540), .B(n12538), .Z(n12539) );
  XOR U10644 ( .A(n12541), .B(n12542), .Z(n9694) );
  NOR U10645 ( .A(n12543), .B(n12541), .Z(n12542) );
  XOR U10646 ( .A(n12544), .B(n12545), .Z(n9697) );
  NOR U10647 ( .A(n12546), .B(n12544), .Z(n12545) );
  XOR U10648 ( .A(n12547), .B(n12548), .Z(n9700) );
  NOR U10649 ( .A(n12549), .B(n12547), .Z(n12548) );
  XOR U10650 ( .A(n12550), .B(n12551), .Z(n9703) );
  NOR U10651 ( .A(n12552), .B(n12550), .Z(n12551) );
  XOR U10652 ( .A(n12553), .B(n12554), .Z(n9706) );
  NOR U10653 ( .A(n12555), .B(n12553), .Z(n12554) );
  XOR U10654 ( .A(n12556), .B(n12557), .Z(n9709) );
  NOR U10655 ( .A(n12558), .B(n12556), .Z(n12557) );
  XOR U10656 ( .A(n12559), .B(n12560), .Z(n9712) );
  NOR U10657 ( .A(n12561), .B(n12559), .Z(n12560) );
  XOR U10658 ( .A(n12562), .B(n12563), .Z(n9715) );
  NOR U10659 ( .A(n12564), .B(n12562), .Z(n12563) );
  XOR U10660 ( .A(n12565), .B(n12566), .Z(n9718) );
  NOR U10661 ( .A(n12567), .B(n12565), .Z(n12566) );
  XOR U10662 ( .A(n12568), .B(n12569), .Z(n9721) );
  NOR U10663 ( .A(n12570), .B(n12568), .Z(n12569) );
  XOR U10664 ( .A(n12571), .B(n12572), .Z(n9724) );
  NOR U10665 ( .A(n12573), .B(n12571), .Z(n12572) );
  XOR U10666 ( .A(n12574), .B(n12575), .Z(n9727) );
  NOR U10667 ( .A(n12576), .B(n12574), .Z(n12575) );
  XOR U10668 ( .A(n12577), .B(n12578), .Z(n9730) );
  NOR U10669 ( .A(n12579), .B(n12577), .Z(n12578) );
  XOR U10670 ( .A(n12580), .B(n12581), .Z(n9733) );
  NOR U10671 ( .A(n12582), .B(n12580), .Z(n12581) );
  XOR U10672 ( .A(n12583), .B(n12584), .Z(n9736) );
  NOR U10673 ( .A(n12585), .B(n12583), .Z(n12584) );
  XOR U10674 ( .A(n12586), .B(n12587), .Z(n9739) );
  NOR U10675 ( .A(n12588), .B(n12586), .Z(n12587) );
  XOR U10676 ( .A(n12589), .B(n12590), .Z(n9742) );
  NOR U10677 ( .A(n12591), .B(n12589), .Z(n12590) );
  XOR U10678 ( .A(n12592), .B(n12593), .Z(n9745) );
  NOR U10679 ( .A(n12594), .B(n12592), .Z(n12593) );
  XOR U10680 ( .A(n12595), .B(n12596), .Z(n9748) );
  NOR U10681 ( .A(n12597), .B(n12595), .Z(n12596) );
  XOR U10682 ( .A(n12598), .B(n12599), .Z(n9751) );
  NOR U10683 ( .A(n12600), .B(n12598), .Z(n12599) );
  XOR U10684 ( .A(n12601), .B(n12602), .Z(n9754) );
  NOR U10685 ( .A(n12603), .B(n12601), .Z(n12602) );
  XOR U10686 ( .A(n12604), .B(n12605), .Z(n9757) );
  NOR U10687 ( .A(n12606), .B(n12604), .Z(n12605) );
  XOR U10688 ( .A(n12607), .B(n12608), .Z(n9760) );
  NOR U10689 ( .A(n12609), .B(n12607), .Z(n12608) );
  XOR U10690 ( .A(n12610), .B(n12611), .Z(n9763) );
  NOR U10691 ( .A(n12612), .B(n12610), .Z(n12611) );
  XOR U10692 ( .A(n12613), .B(n12614), .Z(n9766) );
  NOR U10693 ( .A(n12615), .B(n12613), .Z(n12614) );
  XOR U10694 ( .A(n12616), .B(n12617), .Z(n9769) );
  NOR U10695 ( .A(n12618), .B(n12616), .Z(n12617) );
  XOR U10696 ( .A(n12619), .B(n12620), .Z(n9772) );
  NOR U10697 ( .A(n12621), .B(n12619), .Z(n12620) );
  XOR U10698 ( .A(n12622), .B(n12623), .Z(n9775) );
  NOR U10699 ( .A(n12624), .B(n12622), .Z(n12623) );
  XOR U10700 ( .A(n12625), .B(n12626), .Z(n9778) );
  NOR U10701 ( .A(n12627), .B(n12625), .Z(n12626) );
  XOR U10702 ( .A(n12628), .B(n12629), .Z(n9781) );
  NOR U10703 ( .A(n12630), .B(n12628), .Z(n12629) );
  XOR U10704 ( .A(n12631), .B(n12632), .Z(n9784) );
  NOR U10705 ( .A(n12633), .B(n12631), .Z(n12632) );
  XOR U10706 ( .A(n12634), .B(n12635), .Z(n9787) );
  NOR U10707 ( .A(n12636), .B(n12634), .Z(n12635) );
  XOR U10708 ( .A(n12637), .B(n12638), .Z(n9790) );
  NOR U10709 ( .A(n12639), .B(n12637), .Z(n12638) );
  XOR U10710 ( .A(n12640), .B(n12641), .Z(n9793) );
  NOR U10711 ( .A(n12642), .B(n12640), .Z(n12641) );
  XOR U10712 ( .A(n12643), .B(n12644), .Z(n9796) );
  NOR U10713 ( .A(n12645), .B(n12643), .Z(n12644) );
  XOR U10714 ( .A(n12646), .B(n12647), .Z(n9799) );
  NOR U10715 ( .A(n12648), .B(n12646), .Z(n12647) );
  XOR U10716 ( .A(n12649), .B(n12650), .Z(n9802) );
  NOR U10717 ( .A(n12651), .B(n12649), .Z(n12650) );
  XOR U10718 ( .A(n12652), .B(n12653), .Z(n9805) );
  NOR U10719 ( .A(n12654), .B(n12652), .Z(n12653) );
  XOR U10720 ( .A(n12655), .B(n12656), .Z(n9808) );
  NOR U10721 ( .A(n12657), .B(n12655), .Z(n12656) );
  XOR U10722 ( .A(n12658), .B(n12659), .Z(n9811) );
  NOR U10723 ( .A(n12660), .B(n12658), .Z(n12659) );
  XOR U10724 ( .A(n12661), .B(n12662), .Z(n9814) );
  NOR U10725 ( .A(n12663), .B(n12661), .Z(n12662) );
  XOR U10726 ( .A(n12664), .B(n12665), .Z(n9817) );
  NOR U10727 ( .A(n12666), .B(n12664), .Z(n12665) );
  XOR U10728 ( .A(n12667), .B(n12668), .Z(n9820) );
  NOR U10729 ( .A(n12669), .B(n12667), .Z(n12668) );
  XOR U10730 ( .A(n12670), .B(n12671), .Z(n9823) );
  NOR U10731 ( .A(n12672), .B(n12670), .Z(n12671) );
  XOR U10732 ( .A(n12673), .B(n12674), .Z(n9826) );
  NOR U10733 ( .A(n12675), .B(n12673), .Z(n12674) );
  XOR U10734 ( .A(n12676), .B(n12677), .Z(n9829) );
  NOR U10735 ( .A(n12678), .B(n12676), .Z(n12677) );
  XOR U10736 ( .A(n12679), .B(n12680), .Z(n9832) );
  NOR U10737 ( .A(n12681), .B(n12679), .Z(n12680) );
  XOR U10738 ( .A(n12682), .B(n12683), .Z(n9835) );
  NOR U10739 ( .A(n12684), .B(n12682), .Z(n12683) );
  XOR U10740 ( .A(n12685), .B(n12686), .Z(n9838) );
  NOR U10741 ( .A(n12687), .B(n12685), .Z(n12686) );
  XOR U10742 ( .A(n12688), .B(n12689), .Z(n9841) );
  NOR U10743 ( .A(n12690), .B(n12688), .Z(n12689) );
  XOR U10744 ( .A(n12691), .B(n12692), .Z(n9844) );
  NOR U10745 ( .A(n12693), .B(n12691), .Z(n12692) );
  XOR U10746 ( .A(n12694), .B(n12695), .Z(n9847) );
  NOR U10747 ( .A(n12696), .B(n12694), .Z(n12695) );
  XOR U10748 ( .A(n12697), .B(n12698), .Z(n9850) );
  NOR U10749 ( .A(n12699), .B(n12697), .Z(n12698) );
  XOR U10750 ( .A(n12700), .B(n12701), .Z(n9853) );
  NOR U10751 ( .A(n12702), .B(n12700), .Z(n12701) );
  XOR U10752 ( .A(n12703), .B(n12704), .Z(n9856) );
  NOR U10753 ( .A(n12705), .B(n12703), .Z(n12704) );
  XOR U10754 ( .A(n12706), .B(n12707), .Z(n9859) );
  NOR U10755 ( .A(n12708), .B(n12706), .Z(n12707) );
  XOR U10756 ( .A(n12709), .B(n12710), .Z(n9862) );
  NOR U10757 ( .A(n12711), .B(n12709), .Z(n12710) );
  XOR U10758 ( .A(n12712), .B(n12713), .Z(n9865) );
  NOR U10759 ( .A(n12714), .B(n12712), .Z(n12713) );
  XOR U10760 ( .A(n12715), .B(n12716), .Z(n9868) );
  NOR U10761 ( .A(n12717), .B(n12715), .Z(n12716) );
  XOR U10762 ( .A(n12718), .B(n12719), .Z(n9871) );
  NOR U10763 ( .A(n12720), .B(n12718), .Z(n12719) );
  XOR U10764 ( .A(n12721), .B(n12722), .Z(n9874) );
  NOR U10765 ( .A(n12723), .B(n12721), .Z(n12722) );
  XOR U10766 ( .A(n12724), .B(n12725), .Z(n9877) );
  NOR U10767 ( .A(n12726), .B(n12724), .Z(n12725) );
  XOR U10768 ( .A(n12727), .B(n12728), .Z(n9880) );
  NOR U10769 ( .A(n12729), .B(n12727), .Z(n12728) );
  XOR U10770 ( .A(n12730), .B(n12731), .Z(n9883) );
  NOR U10771 ( .A(n12732), .B(n12730), .Z(n12731) );
  XOR U10772 ( .A(n12733), .B(n12734), .Z(n9886) );
  AND U10773 ( .A(n12735), .B(n12733), .Z(n12734) );
  XOR U10774 ( .A(n12736), .B(n12737), .Z(n9889) );
  AND U10775 ( .A(n104), .B(n12736), .Z(n12737) );
  XNOR U10776 ( .A(n12738), .B(n11306), .Z(n11308) );
  IV U10777 ( .A(n87), .Z(n12738) );
  XOR U10778 ( .A(n11303), .B(n11302), .Z(n87) );
  XNOR U10779 ( .A(n11300), .B(n11299), .Z(n11302) );
  XNOR U10780 ( .A(n11297), .B(n11296), .Z(n11299) );
  XNOR U10781 ( .A(n11294), .B(n11293), .Z(n11296) );
  XNOR U10782 ( .A(n11291), .B(n11290), .Z(n11293) );
  XNOR U10783 ( .A(n11288), .B(n11287), .Z(n11290) );
  XNOR U10784 ( .A(n11285), .B(n11284), .Z(n11287) );
  XNOR U10785 ( .A(n11282), .B(n11281), .Z(n11284) );
  XNOR U10786 ( .A(n11279), .B(n11278), .Z(n11281) );
  XNOR U10787 ( .A(n11276), .B(n11275), .Z(n11278) );
  XNOR U10788 ( .A(n11273), .B(n11272), .Z(n11275) );
  XNOR U10789 ( .A(n11270), .B(n11269), .Z(n11272) );
  XNOR U10790 ( .A(n11267), .B(n11266), .Z(n11269) );
  XNOR U10791 ( .A(n11264), .B(n11263), .Z(n11266) );
  XNOR U10792 ( .A(n11261), .B(n11260), .Z(n11263) );
  XNOR U10793 ( .A(n11258), .B(n11257), .Z(n11260) );
  XNOR U10794 ( .A(n11255), .B(n11254), .Z(n11257) );
  XNOR U10795 ( .A(n11252), .B(n11251), .Z(n11254) );
  XNOR U10796 ( .A(n11249), .B(n11248), .Z(n11251) );
  XNOR U10797 ( .A(n11246), .B(n11245), .Z(n11248) );
  XNOR U10798 ( .A(n11243), .B(n11242), .Z(n11245) );
  XNOR U10799 ( .A(n11240), .B(n11239), .Z(n11242) );
  XNOR U10800 ( .A(n11237), .B(n11236), .Z(n11239) );
  XNOR U10801 ( .A(n11234), .B(n11233), .Z(n11236) );
  XNOR U10802 ( .A(n11231), .B(n11230), .Z(n11233) );
  XNOR U10803 ( .A(n11228), .B(n11227), .Z(n11230) );
  XNOR U10804 ( .A(n11225), .B(n11224), .Z(n11227) );
  XNOR U10805 ( .A(n11222), .B(n11221), .Z(n11224) );
  XNOR U10806 ( .A(n11219), .B(n11218), .Z(n11221) );
  XNOR U10807 ( .A(n11216), .B(n11215), .Z(n11218) );
  XNOR U10808 ( .A(n11213), .B(n11212), .Z(n11215) );
  XNOR U10809 ( .A(n11210), .B(n11209), .Z(n11212) );
  XNOR U10810 ( .A(n11207), .B(n11206), .Z(n11209) );
  XNOR U10811 ( .A(n11204), .B(n11203), .Z(n11206) );
  XNOR U10812 ( .A(n11201), .B(n11200), .Z(n11203) );
  XNOR U10813 ( .A(n11198), .B(n11197), .Z(n11200) );
  XNOR U10814 ( .A(n11195), .B(n11194), .Z(n11197) );
  XNOR U10815 ( .A(n11192), .B(n11191), .Z(n11194) );
  XNOR U10816 ( .A(n11189), .B(n11188), .Z(n11191) );
  XNOR U10817 ( .A(n11186), .B(n11185), .Z(n11188) );
  XNOR U10818 ( .A(n11183), .B(n11182), .Z(n11185) );
  XNOR U10819 ( .A(n11180), .B(n11179), .Z(n11182) );
  XNOR U10820 ( .A(n11177), .B(n11176), .Z(n11179) );
  XNOR U10821 ( .A(n11174), .B(n11173), .Z(n11176) );
  XNOR U10822 ( .A(n11171), .B(n11170), .Z(n11173) );
  XNOR U10823 ( .A(n11168), .B(n11167), .Z(n11170) );
  XNOR U10824 ( .A(n11165), .B(n11164), .Z(n11167) );
  XNOR U10825 ( .A(n11162), .B(n11161), .Z(n11164) );
  XNOR U10826 ( .A(n11159), .B(n11158), .Z(n11161) );
  XNOR U10827 ( .A(n11156), .B(n11155), .Z(n11158) );
  XNOR U10828 ( .A(n11153), .B(n11152), .Z(n11155) );
  XNOR U10829 ( .A(n11150), .B(n11149), .Z(n11152) );
  XNOR U10830 ( .A(n11147), .B(n11146), .Z(n11149) );
  XNOR U10831 ( .A(n11144), .B(n11143), .Z(n11146) );
  XNOR U10832 ( .A(n11141), .B(n11140), .Z(n11143) );
  XNOR U10833 ( .A(n11138), .B(n11137), .Z(n11140) );
  XNOR U10834 ( .A(n11135), .B(n11134), .Z(n11137) );
  XNOR U10835 ( .A(n11132), .B(n11131), .Z(n11134) );
  XNOR U10836 ( .A(n11129), .B(n11128), .Z(n11131) );
  XNOR U10837 ( .A(n11126), .B(n11125), .Z(n11128) );
  XNOR U10838 ( .A(n11123), .B(n11122), .Z(n11125) );
  XNOR U10839 ( .A(n11120), .B(n11119), .Z(n11122) );
  XNOR U10840 ( .A(n11117), .B(n11116), .Z(n11119) );
  XNOR U10841 ( .A(n11114), .B(n11113), .Z(n11116) );
  XNOR U10842 ( .A(n11111), .B(n11110), .Z(n11113) );
  XNOR U10843 ( .A(n11108), .B(n11107), .Z(n11110) );
  XNOR U10844 ( .A(n11105), .B(n11104), .Z(n11107) );
  XNOR U10845 ( .A(n11102), .B(n11101), .Z(n11104) );
  XNOR U10846 ( .A(n11099), .B(n11098), .Z(n11101) );
  XNOR U10847 ( .A(n11096), .B(n11095), .Z(n11098) );
  XNOR U10848 ( .A(n11093), .B(n11092), .Z(n11095) );
  XNOR U10849 ( .A(n11090), .B(n11089), .Z(n11092) );
  XNOR U10850 ( .A(n11087), .B(n11086), .Z(n11089) );
  XNOR U10851 ( .A(n11084), .B(n11083), .Z(n11086) );
  XNOR U10852 ( .A(n11081), .B(n11080), .Z(n11083) );
  XNOR U10853 ( .A(n11078), .B(n11077), .Z(n11080) );
  XNOR U10854 ( .A(n11075), .B(n11074), .Z(n11077) );
  XNOR U10855 ( .A(n11072), .B(n11071), .Z(n11074) );
  XNOR U10856 ( .A(n11069), .B(n11068), .Z(n11071) );
  XNOR U10857 ( .A(n11066), .B(n11065), .Z(n11068) );
  XNOR U10858 ( .A(n11063), .B(n11062), .Z(n11065) );
  XNOR U10859 ( .A(n11060), .B(n11059), .Z(n11062) );
  XNOR U10860 ( .A(n11057), .B(n11056), .Z(n11059) );
  XNOR U10861 ( .A(n11054), .B(n11053), .Z(n11056) );
  XNOR U10862 ( .A(n11051), .B(n11050), .Z(n11053) );
  XNOR U10863 ( .A(n11048), .B(n11047), .Z(n11050) );
  XNOR U10864 ( .A(n11045), .B(n11044), .Z(n11047) );
  XNOR U10865 ( .A(n11042), .B(n11041), .Z(n11044) );
  XNOR U10866 ( .A(n11039), .B(n11038), .Z(n11041) );
  XNOR U10867 ( .A(n11036), .B(n11035), .Z(n11038) );
  XNOR U10868 ( .A(n11033), .B(n11032), .Z(n11035) );
  XNOR U10869 ( .A(n11030), .B(n11029), .Z(n11032) );
  XNOR U10870 ( .A(n11027), .B(n11026), .Z(n11029) );
  XNOR U10871 ( .A(n11024), .B(n11023), .Z(n11026) );
  XNOR U10872 ( .A(n11021), .B(n11020), .Z(n11023) );
  XNOR U10873 ( .A(n11018), .B(n11017), .Z(n11020) );
  XNOR U10874 ( .A(n11015), .B(n11014), .Z(n11017) );
  XNOR U10875 ( .A(n11012), .B(n11011), .Z(n11014) );
  XNOR U10876 ( .A(n11009), .B(n11008), .Z(n11011) );
  XNOR U10877 ( .A(n11006), .B(n11005), .Z(n11008) );
  XNOR U10878 ( .A(n11003), .B(n11002), .Z(n11005) );
  XNOR U10879 ( .A(n11000), .B(n10999), .Z(n11002) );
  XNOR U10880 ( .A(n10997), .B(n10996), .Z(n10999) );
  XNOR U10881 ( .A(n10994), .B(n10993), .Z(n10996) );
  XNOR U10882 ( .A(n10991), .B(n10990), .Z(n10993) );
  XNOR U10883 ( .A(n10988), .B(n10987), .Z(n10990) );
  XNOR U10884 ( .A(n10985), .B(n10984), .Z(n10987) );
  XNOR U10885 ( .A(n10982), .B(n10981), .Z(n10984) );
  XNOR U10886 ( .A(n10979), .B(n10978), .Z(n10981) );
  XNOR U10887 ( .A(n10976), .B(n10975), .Z(n10978) );
  XNOR U10888 ( .A(n10973), .B(n10972), .Z(n10975) );
  XNOR U10889 ( .A(n10970), .B(n10969), .Z(n10972) );
  XNOR U10890 ( .A(n10967), .B(n10966), .Z(n10969) );
  XNOR U10891 ( .A(n10964), .B(n10963), .Z(n10966) );
  XNOR U10892 ( .A(n10961), .B(n10960), .Z(n10963) );
  XNOR U10893 ( .A(n10958), .B(n10957), .Z(n10960) );
  XNOR U10894 ( .A(n10955), .B(n10954), .Z(n10957) );
  XNOR U10895 ( .A(n10952), .B(n10951), .Z(n10954) );
  XNOR U10896 ( .A(n10949), .B(n10948), .Z(n10951) );
  XNOR U10897 ( .A(n10946), .B(n10945), .Z(n10948) );
  XNOR U10898 ( .A(n10943), .B(n10942), .Z(n10945) );
  XNOR U10899 ( .A(n10940), .B(n10939), .Z(n10942) );
  XNOR U10900 ( .A(n10937), .B(n10936), .Z(n10939) );
  XNOR U10901 ( .A(n10934), .B(n10933), .Z(n10936) );
  XNOR U10902 ( .A(n10931), .B(n10930), .Z(n10933) );
  XNOR U10903 ( .A(n10928), .B(n10927), .Z(n10930) );
  XNOR U10904 ( .A(n10925), .B(n10924), .Z(n10927) );
  XNOR U10905 ( .A(n10922), .B(n10921), .Z(n10924) );
  XNOR U10906 ( .A(n10919), .B(n10918), .Z(n10921) );
  XNOR U10907 ( .A(n10916), .B(n10915), .Z(n10918) );
  XNOR U10908 ( .A(n10913), .B(n10912), .Z(n10915) );
  XNOR U10909 ( .A(n10910), .B(n10909), .Z(n10912) );
  XNOR U10910 ( .A(n10907), .B(n10906), .Z(n10909) );
  XNOR U10911 ( .A(n10904), .B(n10903), .Z(n10906) );
  XNOR U10912 ( .A(n10901), .B(n10900), .Z(n10903) );
  XNOR U10913 ( .A(n10898), .B(n10897), .Z(n10900) );
  XNOR U10914 ( .A(n10895), .B(n10894), .Z(n10897) );
  XNOR U10915 ( .A(n10892), .B(n10891), .Z(n10894) );
  XNOR U10916 ( .A(n10889), .B(n10888), .Z(n10891) );
  XNOR U10917 ( .A(n10886), .B(n10885), .Z(n10888) );
  XNOR U10918 ( .A(n10883), .B(n10882), .Z(n10885) );
  XNOR U10919 ( .A(n10880), .B(n10879), .Z(n10882) );
  XNOR U10920 ( .A(n10877), .B(n10876), .Z(n10879) );
  XNOR U10921 ( .A(n10874), .B(n10873), .Z(n10876) );
  XNOR U10922 ( .A(n10871), .B(n10870), .Z(n10873) );
  XNOR U10923 ( .A(n10868), .B(n10867), .Z(n10870) );
  XNOR U10924 ( .A(n10865), .B(n10864), .Z(n10867) );
  XNOR U10925 ( .A(n10862), .B(n10861), .Z(n10864) );
  XNOR U10926 ( .A(n10859), .B(n10858), .Z(n10861) );
  XNOR U10927 ( .A(n10856), .B(n10855), .Z(n10858) );
  XNOR U10928 ( .A(n10853), .B(n10852), .Z(n10855) );
  XNOR U10929 ( .A(n10850), .B(n10849), .Z(n10852) );
  XNOR U10930 ( .A(n10847), .B(n10846), .Z(n10849) );
  XNOR U10931 ( .A(n10844), .B(n10843), .Z(n10846) );
  XNOR U10932 ( .A(n10841), .B(n10840), .Z(n10843) );
  XNOR U10933 ( .A(n10838), .B(n10837), .Z(n10840) );
  XNOR U10934 ( .A(n10835), .B(n10834), .Z(n10837) );
  XNOR U10935 ( .A(n10832), .B(n10831), .Z(n10834) );
  XNOR U10936 ( .A(n10829), .B(n10828), .Z(n10831) );
  XNOR U10937 ( .A(n10826), .B(n10825), .Z(n10828) );
  XNOR U10938 ( .A(n10823), .B(n10822), .Z(n10825) );
  XNOR U10939 ( .A(n10820), .B(n10819), .Z(n10822) );
  XNOR U10940 ( .A(n10817), .B(n10816), .Z(n10819) );
  XNOR U10941 ( .A(n10814), .B(n10813), .Z(n10816) );
  XNOR U10942 ( .A(n10811), .B(n10810), .Z(n10813) );
  XNOR U10943 ( .A(n10808), .B(n10807), .Z(n10810) );
  XNOR U10944 ( .A(n10805), .B(n10804), .Z(n10807) );
  XNOR U10945 ( .A(n10802), .B(n10801), .Z(n10804) );
  XNOR U10946 ( .A(n10799), .B(n10798), .Z(n10801) );
  XNOR U10947 ( .A(n10796), .B(n10795), .Z(n10798) );
  XNOR U10948 ( .A(n10793), .B(n10792), .Z(n10795) );
  XNOR U10949 ( .A(n10790), .B(n10789), .Z(n10792) );
  XNOR U10950 ( .A(n10787), .B(n10786), .Z(n10789) );
  XNOR U10951 ( .A(n10784), .B(n10783), .Z(n10786) );
  XNOR U10952 ( .A(n10781), .B(n10780), .Z(n10783) );
  XNOR U10953 ( .A(n10778), .B(n10777), .Z(n10780) );
  XNOR U10954 ( .A(n10775), .B(n10774), .Z(n10777) );
  XNOR U10955 ( .A(n10772), .B(n10771), .Z(n10774) );
  XNOR U10956 ( .A(n10769), .B(n10768), .Z(n10771) );
  XNOR U10957 ( .A(n10766), .B(n10765), .Z(n10768) );
  XNOR U10958 ( .A(n10763), .B(n10762), .Z(n10765) );
  XNOR U10959 ( .A(n10760), .B(n10759), .Z(n10762) );
  XNOR U10960 ( .A(n10757), .B(n10756), .Z(n10759) );
  XNOR U10961 ( .A(n10754), .B(n10753), .Z(n10756) );
  XNOR U10962 ( .A(n10751), .B(n10750), .Z(n10753) );
  XNOR U10963 ( .A(n10748), .B(n10747), .Z(n10750) );
  XNOR U10964 ( .A(n10745), .B(n10744), .Z(n10747) );
  XNOR U10965 ( .A(n10742), .B(n10741), .Z(n10744) );
  XNOR U10966 ( .A(n10739), .B(n10738), .Z(n10741) );
  XNOR U10967 ( .A(n10736), .B(n10735), .Z(n10738) );
  XNOR U10968 ( .A(n10733), .B(n10732), .Z(n10735) );
  XNOR U10969 ( .A(n10730), .B(n10729), .Z(n10732) );
  XNOR U10970 ( .A(n10727), .B(n10726), .Z(n10729) );
  XNOR U10971 ( .A(n10724), .B(n10723), .Z(n10726) );
  XNOR U10972 ( .A(n10721), .B(n10720), .Z(n10723) );
  XNOR U10973 ( .A(n10718), .B(n10717), .Z(n10720) );
  XNOR U10974 ( .A(n10715), .B(n10714), .Z(n10717) );
  XNOR U10975 ( .A(n10712), .B(n10711), .Z(n10714) );
  XNOR U10976 ( .A(n10709), .B(n10708), .Z(n10711) );
  XNOR U10977 ( .A(n10706), .B(n10705), .Z(n10708) );
  XNOR U10978 ( .A(n10703), .B(n10702), .Z(n10705) );
  XNOR U10979 ( .A(n10700), .B(n10699), .Z(n10702) );
  XNOR U10980 ( .A(n10697), .B(n10696), .Z(n10699) );
  XNOR U10981 ( .A(n10694), .B(n10693), .Z(n10696) );
  XNOR U10982 ( .A(n10691), .B(n10690), .Z(n10693) );
  XNOR U10983 ( .A(n10688), .B(n10687), .Z(n10690) );
  XNOR U10984 ( .A(n10685), .B(n10684), .Z(n10687) );
  XNOR U10985 ( .A(n10682), .B(n10681), .Z(n10684) );
  XNOR U10986 ( .A(n10679), .B(n10678), .Z(n10681) );
  XNOR U10987 ( .A(n10676), .B(n10675), .Z(n10678) );
  XNOR U10988 ( .A(n10673), .B(n10672), .Z(n10675) );
  XNOR U10989 ( .A(n10670), .B(n10669), .Z(n10672) );
  XNOR U10990 ( .A(n10667), .B(n10666), .Z(n10669) );
  XNOR U10991 ( .A(n10664), .B(n10663), .Z(n10666) );
  XNOR U10992 ( .A(n10661), .B(n10660), .Z(n10663) );
  XNOR U10993 ( .A(n10658), .B(n10657), .Z(n10660) );
  XNOR U10994 ( .A(n10655), .B(n10654), .Z(n10657) );
  XNOR U10995 ( .A(n10652), .B(n10651), .Z(n10654) );
  XNOR U10996 ( .A(n10649), .B(n10648), .Z(n10651) );
  XNOR U10997 ( .A(n10646), .B(n10645), .Z(n10648) );
  XNOR U10998 ( .A(n10643), .B(n10642), .Z(n10645) );
  XNOR U10999 ( .A(n10640), .B(n10639), .Z(n10642) );
  XNOR U11000 ( .A(n10637), .B(n10636), .Z(n10639) );
  XNOR U11001 ( .A(n10634), .B(n10633), .Z(n10636) );
  XNOR U11002 ( .A(n10631), .B(n10630), .Z(n10633) );
  XNOR U11003 ( .A(n10628), .B(n10627), .Z(n10630) );
  XNOR U11004 ( .A(n10625), .B(n10624), .Z(n10627) );
  XNOR U11005 ( .A(n10622), .B(n10621), .Z(n10624) );
  XNOR U11006 ( .A(n10619), .B(n10618), .Z(n10621) );
  XNOR U11007 ( .A(n10616), .B(n10615), .Z(n10618) );
  XNOR U11008 ( .A(n10613), .B(n10612), .Z(n10615) );
  XNOR U11009 ( .A(n10610), .B(n10609), .Z(n10612) );
  XNOR U11010 ( .A(n10607), .B(n10606), .Z(n10609) );
  XNOR U11011 ( .A(n10604), .B(n10603), .Z(n10606) );
  XNOR U11012 ( .A(n10601), .B(n10600), .Z(n10603) );
  XNOR U11013 ( .A(n10598), .B(n10597), .Z(n10600) );
  XNOR U11014 ( .A(n10595), .B(n10594), .Z(n10597) );
  XNOR U11015 ( .A(n10592), .B(n10591), .Z(n10594) );
  XNOR U11016 ( .A(n10589), .B(n10588), .Z(n10591) );
  XNOR U11017 ( .A(n10586), .B(n10585), .Z(n10588) );
  XNOR U11018 ( .A(n10583), .B(n10582), .Z(n10585) );
  XNOR U11019 ( .A(n10580), .B(n10579), .Z(n10582) );
  XNOR U11020 ( .A(n10577), .B(n10576), .Z(n10579) );
  XNOR U11021 ( .A(n10574), .B(n10573), .Z(n10576) );
  XNOR U11022 ( .A(n10571), .B(n10570), .Z(n10573) );
  XNOR U11023 ( .A(n10568), .B(n10567), .Z(n10570) );
  XNOR U11024 ( .A(n10565), .B(n10564), .Z(n10567) );
  XNOR U11025 ( .A(n10562), .B(n10561), .Z(n10564) );
  XNOR U11026 ( .A(n10559), .B(n10558), .Z(n10561) );
  XNOR U11027 ( .A(n10556), .B(n10555), .Z(n10558) );
  XNOR U11028 ( .A(n10553), .B(n10552), .Z(n10555) );
  XNOR U11029 ( .A(n10550), .B(n10549), .Z(n10552) );
  XNOR U11030 ( .A(n10547), .B(n10546), .Z(n10549) );
  XNOR U11031 ( .A(n10544), .B(n10543), .Z(n10546) );
  XNOR U11032 ( .A(n10541), .B(n10540), .Z(n10543) );
  XNOR U11033 ( .A(n10538), .B(n10537), .Z(n10540) );
  XNOR U11034 ( .A(n10535), .B(n10534), .Z(n10537) );
  XNOR U11035 ( .A(n10532), .B(n10531), .Z(n10534) );
  XNOR U11036 ( .A(n10529), .B(n10528), .Z(n10531) );
  XNOR U11037 ( .A(n10526), .B(n10525), .Z(n10528) );
  XNOR U11038 ( .A(n10523), .B(n10522), .Z(n10525) );
  XNOR U11039 ( .A(n10520), .B(n10519), .Z(n10522) );
  XNOR U11040 ( .A(n10517), .B(n10516), .Z(n10519) );
  XNOR U11041 ( .A(n10514), .B(n10513), .Z(n10516) );
  XNOR U11042 ( .A(n10511), .B(n10510), .Z(n10513) );
  XNOR U11043 ( .A(n10508), .B(n10507), .Z(n10510) );
  XNOR U11044 ( .A(n10505), .B(n10504), .Z(n10507) );
  XNOR U11045 ( .A(n10502), .B(n10501), .Z(n10504) );
  XNOR U11046 ( .A(n10499), .B(n10498), .Z(n10501) );
  XNOR U11047 ( .A(n10496), .B(n10495), .Z(n10498) );
  XNOR U11048 ( .A(n10493), .B(n10492), .Z(n10495) );
  XNOR U11049 ( .A(n10490), .B(n10489), .Z(n10492) );
  XNOR U11050 ( .A(n10487), .B(n10486), .Z(n10489) );
  XNOR U11051 ( .A(n10484), .B(n10483), .Z(n10486) );
  XNOR U11052 ( .A(n10481), .B(n10480), .Z(n10483) );
  XNOR U11053 ( .A(n10478), .B(n10477), .Z(n10480) );
  XNOR U11054 ( .A(n10475), .B(n10474), .Z(n10477) );
  XNOR U11055 ( .A(n10472), .B(n10471), .Z(n10474) );
  XNOR U11056 ( .A(n10469), .B(n10468), .Z(n10471) );
  XNOR U11057 ( .A(n10466), .B(n10465), .Z(n10468) );
  XNOR U11058 ( .A(n10463), .B(n10462), .Z(n10465) );
  XNOR U11059 ( .A(n10460), .B(n10459), .Z(n10462) );
  XNOR U11060 ( .A(n10457), .B(n10456), .Z(n10459) );
  XNOR U11061 ( .A(n10454), .B(n10453), .Z(n10456) );
  XNOR U11062 ( .A(n10451), .B(n10450), .Z(n10453) );
  XNOR U11063 ( .A(n10448), .B(n10447), .Z(n10450) );
  XNOR U11064 ( .A(n10445), .B(n10444), .Z(n10447) );
  XNOR U11065 ( .A(n10442), .B(n10441), .Z(n10444) );
  XNOR U11066 ( .A(n10439), .B(n10438), .Z(n10441) );
  XNOR U11067 ( .A(n10436), .B(n10435), .Z(n10438) );
  XNOR U11068 ( .A(n10433), .B(n10432), .Z(n10435) );
  XNOR U11069 ( .A(n10430), .B(n10429), .Z(n10432) );
  XNOR U11070 ( .A(n10427), .B(n10426), .Z(n10429) );
  XNOR U11071 ( .A(n10424), .B(n10423), .Z(n10426) );
  XNOR U11072 ( .A(n10421), .B(n10420), .Z(n10423) );
  XNOR U11073 ( .A(n10418), .B(n10417), .Z(n10420) );
  XNOR U11074 ( .A(n10415), .B(n10414), .Z(n10417) );
  XNOR U11075 ( .A(n10412), .B(n10411), .Z(n10414) );
  XNOR U11076 ( .A(n10409), .B(n10408), .Z(n10411) );
  XNOR U11077 ( .A(n10406), .B(n10405), .Z(n10408) );
  XNOR U11078 ( .A(n10403), .B(n10402), .Z(n10405) );
  XNOR U11079 ( .A(n10400), .B(n10399), .Z(n10402) );
  XNOR U11080 ( .A(n10397), .B(n10396), .Z(n10399) );
  XNOR U11081 ( .A(n10394), .B(n10393), .Z(n10396) );
  XNOR U11082 ( .A(n10391), .B(n10390), .Z(n10393) );
  XNOR U11083 ( .A(n10388), .B(n10387), .Z(n10390) );
  XNOR U11084 ( .A(n10385), .B(n10384), .Z(n10387) );
  XNOR U11085 ( .A(n10382), .B(n10381), .Z(n10384) );
  XNOR U11086 ( .A(n10379), .B(n10378), .Z(n10381) );
  XNOR U11087 ( .A(n10376), .B(n10375), .Z(n10378) );
  XNOR U11088 ( .A(n10373), .B(n10372), .Z(n10375) );
  XNOR U11089 ( .A(n10370), .B(n10369), .Z(n10372) );
  XNOR U11090 ( .A(n10367), .B(n10366), .Z(n10369) );
  XNOR U11091 ( .A(n10364), .B(n10363), .Z(n10366) );
  XNOR U11092 ( .A(n10361), .B(n10360), .Z(n10363) );
  XNOR U11093 ( .A(n10358), .B(n10357), .Z(n10360) );
  XNOR U11094 ( .A(n10355), .B(n10354), .Z(n10357) );
  XNOR U11095 ( .A(n10352), .B(n10351), .Z(n10354) );
  XNOR U11096 ( .A(n10349), .B(n10348), .Z(n10351) );
  XNOR U11097 ( .A(n10346), .B(n10345), .Z(n10348) );
  XNOR U11098 ( .A(n10343), .B(n10342), .Z(n10345) );
  XNOR U11099 ( .A(n10340), .B(n10339), .Z(n10342) );
  XNOR U11100 ( .A(n10337), .B(n10336), .Z(n10339) );
  XNOR U11101 ( .A(n10334), .B(n10333), .Z(n10336) );
  XNOR U11102 ( .A(n10331), .B(n10330), .Z(n10333) );
  XNOR U11103 ( .A(n10328), .B(n10327), .Z(n10330) );
  XNOR U11104 ( .A(n10325), .B(n10324), .Z(n10327) );
  XNOR U11105 ( .A(n10322), .B(n10321), .Z(n10324) );
  XNOR U11106 ( .A(n10319), .B(n10318), .Z(n10321) );
  XNOR U11107 ( .A(n10316), .B(n10315), .Z(n10318) );
  XNOR U11108 ( .A(n10313), .B(n10312), .Z(n10315) );
  XNOR U11109 ( .A(n10310), .B(n10309), .Z(n10312) );
  XNOR U11110 ( .A(n10307), .B(n10306), .Z(n10309) );
  XNOR U11111 ( .A(n10304), .B(n10303), .Z(n10306) );
  XNOR U11112 ( .A(n10301), .B(n10300), .Z(n10303) );
  XNOR U11113 ( .A(n10298), .B(n10297), .Z(n10300) );
  XNOR U11114 ( .A(n10295), .B(n10294), .Z(n10297) );
  XNOR U11115 ( .A(n10292), .B(n10291), .Z(n10294) );
  XNOR U11116 ( .A(n10289), .B(n10288), .Z(n10291) );
  XNOR U11117 ( .A(n10286), .B(n10285), .Z(n10288) );
  XNOR U11118 ( .A(n10283), .B(n10282), .Z(n10285) );
  XNOR U11119 ( .A(n10280), .B(n10279), .Z(n10282) );
  XNOR U11120 ( .A(n10277), .B(n10276), .Z(n10279) );
  XNOR U11121 ( .A(n10274), .B(n10273), .Z(n10276) );
  XNOR U11122 ( .A(n10271), .B(n10270), .Z(n10273) );
  XNOR U11123 ( .A(n10268), .B(n10267), .Z(n10270) );
  XNOR U11124 ( .A(n10265), .B(n10264), .Z(n10267) );
  XNOR U11125 ( .A(n10262), .B(n10261), .Z(n10264) );
  XNOR U11126 ( .A(n10259), .B(n10258), .Z(n10261) );
  XNOR U11127 ( .A(n10256), .B(n10255), .Z(n10258) );
  XNOR U11128 ( .A(n10253), .B(n10252), .Z(n10255) );
  XNOR U11129 ( .A(n10250), .B(n10249), .Z(n10252) );
  XNOR U11130 ( .A(n10247), .B(n10246), .Z(n10249) );
  XNOR U11131 ( .A(n10244), .B(n10243), .Z(n10246) );
  XNOR U11132 ( .A(n10241), .B(n10240), .Z(n10243) );
  XNOR U11133 ( .A(n10238), .B(n10237), .Z(n10240) );
  XNOR U11134 ( .A(n10235), .B(n10234), .Z(n10237) );
  XNOR U11135 ( .A(n10232), .B(n10231), .Z(n10234) );
  XNOR U11136 ( .A(n10229), .B(n10228), .Z(n10231) );
  XNOR U11137 ( .A(n10226), .B(n10225), .Z(n10228) );
  XNOR U11138 ( .A(n10223), .B(n10222), .Z(n10225) );
  XNOR U11139 ( .A(n10220), .B(n10219), .Z(n10222) );
  XNOR U11140 ( .A(n10217), .B(n10216), .Z(n10219) );
  XNOR U11141 ( .A(n10214), .B(n10213), .Z(n10216) );
  XNOR U11142 ( .A(n10211), .B(n10210), .Z(n10213) );
  XNOR U11143 ( .A(n10208), .B(n10207), .Z(n10210) );
  XNOR U11144 ( .A(n10205), .B(n10204), .Z(n10207) );
  XNOR U11145 ( .A(n10202), .B(n10201), .Z(n10204) );
  XNOR U11146 ( .A(n10199), .B(n10198), .Z(n10201) );
  XNOR U11147 ( .A(n10196), .B(n10195), .Z(n10198) );
  XNOR U11148 ( .A(n10193), .B(n10192), .Z(n10195) );
  XNOR U11149 ( .A(n10190), .B(n10189), .Z(n10192) );
  XNOR U11150 ( .A(n10187), .B(n10186), .Z(n10189) );
  XNOR U11151 ( .A(n10184), .B(n10183), .Z(n10186) );
  XNOR U11152 ( .A(n10181), .B(n10180), .Z(n10183) );
  XNOR U11153 ( .A(n10178), .B(n10177), .Z(n10180) );
  XNOR U11154 ( .A(n10175), .B(n10174), .Z(n10177) );
  XNOR U11155 ( .A(n10172), .B(n10171), .Z(n10174) );
  XNOR U11156 ( .A(n10169), .B(n10168), .Z(n10171) );
  XNOR U11157 ( .A(n10166), .B(n10165), .Z(n10168) );
  XNOR U11158 ( .A(n10163), .B(n10162), .Z(n10165) );
  XNOR U11159 ( .A(n10160), .B(n10159), .Z(n10162) );
  XNOR U11160 ( .A(n10157), .B(n10156), .Z(n10159) );
  XNOR U11161 ( .A(n10154), .B(n10153), .Z(n10156) );
  XNOR U11162 ( .A(n10151), .B(n10150), .Z(n10153) );
  XNOR U11163 ( .A(n10148), .B(n10147), .Z(n10150) );
  XNOR U11164 ( .A(n10145), .B(n10144), .Z(n10147) );
  XNOR U11165 ( .A(n10142), .B(n10141), .Z(n10144) );
  XNOR U11166 ( .A(n10139), .B(n10138), .Z(n10141) );
  XNOR U11167 ( .A(n10136), .B(n10135), .Z(n10138) );
  XNOR U11168 ( .A(n10133), .B(n10132), .Z(n10135) );
  XNOR U11169 ( .A(n10130), .B(n10129), .Z(n10132) );
  XOR U11170 ( .A(n12739), .B(n10126), .Z(n10129) );
  XOR U11171 ( .A(n10124), .B(n10123), .Z(n10126) );
  XOR U11172 ( .A(n10121), .B(n10120), .Z(n10123) );
  XOR U11173 ( .A(n10117), .B(n10118), .Z(n10120) );
  AND U11174 ( .A(n12740), .B(n12741), .Z(n10118) );
  XOR U11175 ( .A(n10114), .B(n10115), .Z(n10117) );
  AND U11176 ( .A(n12742), .B(n12743), .Z(n10115) );
  XOR U11177 ( .A(n10111), .B(n10112), .Z(n10114) );
  AND U11178 ( .A(n12744), .B(n12745), .Z(n10112) );
  XOR U11179 ( .A(n10108), .B(n10109), .Z(n10111) );
  AND U11180 ( .A(n12746), .B(n12747), .Z(n10109) );
  XNOR U11181 ( .A(n9893), .B(n10106), .Z(n10108) );
  AND U11182 ( .A(n12748), .B(n12749), .Z(n10106) );
  XOR U11183 ( .A(n9895), .B(n9894), .Z(n9893) );
  AND U11184 ( .A(n12750), .B(n12751), .Z(n9894) );
  XOR U11185 ( .A(n9897), .B(n9896), .Z(n9895) );
  AND U11186 ( .A(n12752), .B(n12753), .Z(n9896) );
  XOR U11187 ( .A(n9899), .B(n9898), .Z(n9897) );
  AND U11188 ( .A(n12754), .B(n12755), .Z(n9898) );
  XOR U11189 ( .A(n9901), .B(n9900), .Z(n9899) );
  AND U11190 ( .A(n12756), .B(n12757), .Z(n9900) );
  XOR U11191 ( .A(n9903), .B(n9902), .Z(n9901) );
  AND U11192 ( .A(n12758), .B(n12759), .Z(n9902) );
  XOR U11193 ( .A(n9905), .B(n9904), .Z(n9903) );
  AND U11194 ( .A(n12760), .B(n12761), .Z(n9904) );
  XOR U11195 ( .A(n9907), .B(n9906), .Z(n9905) );
  AND U11196 ( .A(n12762), .B(n12763), .Z(n9906) );
  XOR U11197 ( .A(n9909), .B(n9908), .Z(n9907) );
  AND U11198 ( .A(n12764), .B(n12765), .Z(n9908) );
  XOR U11199 ( .A(n9911), .B(n9910), .Z(n9909) );
  AND U11200 ( .A(n12766), .B(n12767), .Z(n9910) );
  XOR U11201 ( .A(n9913), .B(n9912), .Z(n9911) );
  AND U11202 ( .A(n12768), .B(n12769), .Z(n9912) );
  XOR U11203 ( .A(n9915), .B(n9914), .Z(n9913) );
  AND U11204 ( .A(n12770), .B(n12771), .Z(n9914) );
  XOR U11205 ( .A(n9917), .B(n9916), .Z(n9915) );
  AND U11206 ( .A(n12772), .B(n12773), .Z(n9916) );
  XOR U11207 ( .A(n9919), .B(n9918), .Z(n9917) );
  AND U11208 ( .A(n12774), .B(n12775), .Z(n9918) );
  XOR U11209 ( .A(n9921), .B(n9920), .Z(n9919) );
  AND U11210 ( .A(n12776), .B(n12777), .Z(n9920) );
  XOR U11211 ( .A(n9923), .B(n9922), .Z(n9921) );
  AND U11212 ( .A(n12778), .B(n12779), .Z(n9922) );
  XOR U11213 ( .A(n9925), .B(n9924), .Z(n9923) );
  AND U11214 ( .A(n12780), .B(n12781), .Z(n9924) );
  XOR U11215 ( .A(n9927), .B(n9926), .Z(n9925) );
  AND U11216 ( .A(n12782), .B(n12783), .Z(n9926) );
  XOR U11217 ( .A(n9929), .B(n9928), .Z(n9927) );
  AND U11218 ( .A(n12784), .B(n12785), .Z(n9928) );
  XOR U11219 ( .A(n9931), .B(n9930), .Z(n9929) );
  AND U11220 ( .A(n12786), .B(n12787), .Z(n9930) );
  XOR U11221 ( .A(n9933), .B(n9932), .Z(n9931) );
  AND U11222 ( .A(n12788), .B(n12789), .Z(n9932) );
  XOR U11223 ( .A(n9935), .B(n9934), .Z(n9933) );
  AND U11224 ( .A(n12790), .B(n12791), .Z(n9934) );
  XOR U11225 ( .A(n9937), .B(n9936), .Z(n9935) );
  AND U11226 ( .A(n12792), .B(n12793), .Z(n9936) );
  XOR U11227 ( .A(n9939), .B(n9938), .Z(n9937) );
  AND U11228 ( .A(n12794), .B(n12795), .Z(n9938) );
  XOR U11229 ( .A(n9941), .B(n9940), .Z(n9939) );
  AND U11230 ( .A(n12796), .B(n12797), .Z(n9940) );
  XOR U11231 ( .A(n9943), .B(n9942), .Z(n9941) );
  AND U11232 ( .A(n12798), .B(n12799), .Z(n9942) );
  XOR U11233 ( .A(n9945), .B(n9944), .Z(n9943) );
  AND U11234 ( .A(n12800), .B(n12801), .Z(n9944) );
  XOR U11235 ( .A(n9947), .B(n9946), .Z(n9945) );
  AND U11236 ( .A(n12802), .B(n12803), .Z(n9946) );
  XOR U11237 ( .A(n9949), .B(n9948), .Z(n9947) );
  AND U11238 ( .A(n12804), .B(n12805), .Z(n9948) );
  XOR U11239 ( .A(n9951), .B(n9950), .Z(n9949) );
  AND U11240 ( .A(n12806), .B(n12807), .Z(n9950) );
  XOR U11241 ( .A(n9953), .B(n9952), .Z(n9951) );
  AND U11242 ( .A(n12808), .B(n12809), .Z(n9952) );
  XOR U11243 ( .A(n9955), .B(n9954), .Z(n9953) );
  AND U11244 ( .A(n12810), .B(n12811), .Z(n9954) );
  XOR U11245 ( .A(n9957), .B(n9956), .Z(n9955) );
  AND U11246 ( .A(n12812), .B(n12813), .Z(n9956) );
  XOR U11247 ( .A(n9959), .B(n9958), .Z(n9957) );
  AND U11248 ( .A(n12814), .B(n12815), .Z(n9958) );
  XOR U11249 ( .A(n9961), .B(n9960), .Z(n9959) );
  AND U11250 ( .A(n12816), .B(n12817), .Z(n9960) );
  XOR U11251 ( .A(n9963), .B(n9962), .Z(n9961) );
  AND U11252 ( .A(n12818), .B(n12819), .Z(n9962) );
  XOR U11253 ( .A(n9965), .B(n9964), .Z(n9963) );
  AND U11254 ( .A(n12820), .B(n12821), .Z(n9964) );
  XOR U11255 ( .A(n9967), .B(n9966), .Z(n9965) );
  AND U11256 ( .A(n12822), .B(n12823), .Z(n9966) );
  XOR U11257 ( .A(n9969), .B(n9968), .Z(n9967) );
  AND U11258 ( .A(n12824), .B(n12825), .Z(n9968) );
  XOR U11259 ( .A(n9971), .B(n9970), .Z(n9969) );
  AND U11260 ( .A(n12826), .B(n12827), .Z(n9970) );
  XOR U11261 ( .A(n10101), .B(n9972), .Z(n9971) );
  AND U11262 ( .A(n12828), .B(n12829), .Z(n9972) );
  XOR U11263 ( .A(n10104), .B(n10102), .Z(n10101) );
  AND U11264 ( .A(n12830), .B(n12831), .Z(n10102) );
  XOR U11265 ( .A(n9974), .B(n10105), .Z(n10104) );
  AND U11266 ( .A(n12832), .B(n12833), .Z(n10105) );
  XOR U11267 ( .A(n9976), .B(n9975), .Z(n9974) );
  AND U11268 ( .A(n12834), .B(n12835), .Z(n9975) );
  XOR U11269 ( .A(n10097), .B(n9977), .Z(n9976) );
  AND U11270 ( .A(n12836), .B(n12837), .Z(n9977) );
  XOR U11271 ( .A(n10099), .B(n10098), .Z(n10097) );
  AND U11272 ( .A(n12838), .B(n12839), .Z(n10098) );
  XOR U11273 ( .A(n9985), .B(n10100), .Z(n10099) );
  AND U11274 ( .A(n12840), .B(n12841), .Z(n10100) );
  XOR U11275 ( .A(n9981), .B(n9986), .Z(n9985) );
  AND U11276 ( .A(n12842), .B(n12843), .Z(n9986) );
  XOR U11277 ( .A(n9983), .B(n9982), .Z(n9981) );
  AND U11278 ( .A(n12844), .B(n12845), .Z(n9982) );
  XOR U11279 ( .A(n10095), .B(n9984), .Z(n9983) );
  AND U11280 ( .A(n12846), .B(n12847), .Z(n9984) );
  XNOR U11281 ( .A(n10004), .B(n10096), .Z(n10095) );
  AND U11282 ( .A(n12848), .B(n12849), .Z(n10096) );
  XOR U11283 ( .A(n10003), .B(n9995), .Z(n10004) );
  AND U11284 ( .A(n12850), .B(n12851), .Z(n9995) );
  XNOR U11285 ( .A(n9998), .B(n9994), .Z(n10003) );
  AND U11286 ( .A(n12852), .B(n12853), .Z(n9994) );
  XOR U11287 ( .A(n10024), .B(n9999), .Z(n9998) );
  AND U11288 ( .A(n12854), .B(n12855), .Z(n9999) );
  XNOR U11289 ( .A(n10015), .B(n10025), .Z(n10024) );
  AND U11290 ( .A(n12856), .B(n12857), .Z(n10025) );
  XOR U11291 ( .A(n10013), .B(n10014), .Z(n10015) );
  AND U11292 ( .A(n12858), .B(n12859), .Z(n10014) );
  XNOR U11293 ( .A(n10007), .B(n10012), .Z(n10013) );
  AND U11294 ( .A(n12860), .B(n12861), .Z(n10012) );
  XOR U11295 ( .A(n10026), .B(n10008), .Z(n10007) );
  AND U11296 ( .A(n12862), .B(n12863), .Z(n10008) );
  XNOR U11297 ( .A(n10092), .B(n10027), .Z(n10026) );
  AND U11298 ( .A(n12864), .B(n12865), .Z(n10027) );
  XOR U11299 ( .A(n10091), .B(n10083), .Z(n10092) );
  AND U11300 ( .A(n12866), .B(n12867), .Z(n10083) );
  XNOR U11301 ( .A(n10086), .B(n10082), .Z(n10091) );
  AND U11302 ( .A(n12868), .B(n12869), .Z(n10082) );
  XOR U11303 ( .A(n10030), .B(n10087), .Z(n10086) );
  AND U11304 ( .A(n12870), .B(n12871), .Z(n10087) );
  XNOR U11305 ( .A(n10079), .B(n10031), .Z(n10030) );
  AND U11306 ( .A(n12872), .B(n12873), .Z(n10031) );
  XOR U11307 ( .A(n10078), .B(n10070), .Z(n10079) );
  AND U11308 ( .A(n12874), .B(n12875), .Z(n10070) );
  XNOR U11309 ( .A(n10073), .B(n10069), .Z(n10078) );
  AND U11310 ( .A(n12876), .B(n12877), .Z(n10069) );
  XOR U11311 ( .A(n12878), .B(n12879), .Z(n10073) );
  XOR U11312 ( .A(n10063), .B(n10064), .Z(n12879) );
  AND U11313 ( .A(n12880), .B(n12881), .Z(n10064) );
  AND U11314 ( .A(n12882), .B(n12883), .Z(n10063) );
  XOR U11315 ( .A(n12884), .B(n10074), .Z(n12878) );
  AND U11316 ( .A(n12885), .B(n12886), .Z(n10074) );
  XOR U11317 ( .A(n12887), .B(n12888), .Z(n12884) );
  XOR U11318 ( .A(n12889), .B(n12890), .Z(n12888) );
  XOR U11319 ( .A(n10056), .B(n10057), .Z(n12890) );
  AND U11320 ( .A(n12891), .B(n12892), .Z(n10057) );
  AND U11321 ( .A(n12893), .B(n12894), .Z(n10056) );
  XOR U11322 ( .A(n10050), .B(n10055), .Z(n12889) );
  AND U11323 ( .A(n12895), .B(n12896), .Z(n10055) );
  AND U11324 ( .A(n12897), .B(n12898), .Z(n10050) );
  XOR U11325 ( .A(n12899), .B(n12900), .Z(n12887) );
  XOR U11326 ( .A(n10058), .B(n10061), .Z(n12900) );
  AND U11327 ( .A(n12901), .B(n12902), .Z(n10061) );
  AND U11328 ( .A(n12903), .B(n12904), .Z(n10058) );
  XOR U11329 ( .A(n12905), .B(n10062), .Z(n12899) );
  AND U11330 ( .A(n12906), .B(n12907), .Z(n10062) );
  XOR U11331 ( .A(n12908), .B(n12909), .Z(n12905) );
  XOR U11332 ( .A(n12910), .B(n12911), .Z(n12909) );
  XOR U11333 ( .A(n10043), .B(n10044), .Z(n12911) );
  AND U11334 ( .A(n12912), .B(n12913), .Z(n10044) );
  AND U11335 ( .A(n12914), .B(n12915), .Z(n10043) );
  XOR U11336 ( .A(n10041), .B(n10039), .Z(n12910) );
  AND U11337 ( .A(n12916), .B(n12917), .Z(n10039) );
  AND U11338 ( .A(n12918), .B(n12919), .Z(n10041) );
  XOR U11339 ( .A(n12920), .B(n12921), .Z(n12908) );
  XOR U11340 ( .A(n10047), .B(n10048), .Z(n12921) );
  AND U11341 ( .A(n12922), .B(n12923), .Z(n10048) );
  AND U11342 ( .A(n12924), .B(n12925), .Z(n10047) );
  XOR U11343 ( .A(n10042), .B(n10049), .Z(n12920) );
  AND U11344 ( .A(n12926), .B(n12927), .Z(n10049) );
  XOR U11345 ( .A(n12928), .B(n12929), .Z(n10042) );
  XOR U11346 ( .A(n12930), .B(n12931), .Z(n12929) );
  XOR U11347 ( .A(n12932), .B(n12933), .Z(n12931) );
  NOR U11348 ( .A(n12934), .B(n12935), .Z(n12933) );
  NOR U11349 ( .A(n12936), .B(n12937), .Z(n12932) );
  AND U11350 ( .A(n12938), .B(n12939), .Z(n12937) );
  IV U11351 ( .A(n12940), .Z(n12936) );
  NOR U11352 ( .A(n12941), .B(n12942), .Z(n12940) );
  AND U11353 ( .A(n12934), .B(n12943), .Z(n12942) );
  AND U11354 ( .A(n12935), .B(n12944), .Z(n12941) );
  XOR U11355 ( .A(n12945), .B(n12946), .Z(n12930) );
  NOR U11356 ( .A(n12947), .B(n12948), .Z(n12946) );
  NOR U11357 ( .A(n12949), .B(n12950), .Z(n12945) );
  AND U11358 ( .A(n12951), .B(n12952), .Z(n12950) );
  IV U11359 ( .A(n12953), .Z(n12949) );
  NOR U11360 ( .A(n12954), .B(n12955), .Z(n12953) );
  AND U11361 ( .A(n12947), .B(n12956), .Z(n12955) );
  AND U11362 ( .A(n12948), .B(n12957), .Z(n12954) );
  XOR U11363 ( .A(n12958), .B(n12959), .Z(n12928) );
  AND U11364 ( .A(n12960), .B(n12961), .Z(n12959) );
  XNOR U11365 ( .A(n12962), .B(n12963), .Z(n12958) );
  AND U11366 ( .A(n12964), .B(n12965), .Z(n12963) );
  AND U11367 ( .A(n12966), .B(n12967), .Z(n12962) );
  AND U11368 ( .A(n12968), .B(n12969), .Z(n12967) );
  NOR U11369 ( .A(n12970), .B(n12971), .Z(n12969) );
  IV U11370 ( .A(n12972), .Z(n12970) );
  NOR U11371 ( .A(n12973), .B(n12974), .Z(n12972) );
  NOR U11372 ( .A(n12975), .B(n12976), .Z(n12968) );
  AND U11373 ( .A(n12977), .B(n12978), .Z(n12966) );
  NOR U11374 ( .A(n12979), .B(n12980), .Z(n12978) );
  NOR U11375 ( .A(n12981), .B(n12982), .Z(n12977) );
  XOR U11376 ( .A(n12983), .B(n12984), .Z(n10121) );
  AND U11377 ( .A(n12983), .B(n12985), .Z(n12984) );
  XNOR U11378 ( .A(n12986), .B(n12987), .Z(n10124) );
  AND U11379 ( .A(n12986), .B(n12988), .Z(n12987) );
  IV U11380 ( .A(n10127), .Z(n12739) );
  XNOR U11381 ( .A(n12989), .B(n12990), .Z(n10127) );
  AND U11382 ( .A(n12989), .B(n12991), .Z(n12990) );
  XNOR U11383 ( .A(n12992), .B(n12993), .Z(n10130) );
  AND U11384 ( .A(n12992), .B(n12994), .Z(n12993) );
  XNOR U11385 ( .A(n12995), .B(n12996), .Z(n10133) );
  AND U11386 ( .A(n12997), .B(n12995), .Z(n12996) );
  XOR U11387 ( .A(n12998), .B(n12999), .Z(n10136) );
  NOR U11388 ( .A(n13000), .B(n12998), .Z(n12999) );
  XOR U11389 ( .A(n13001), .B(n13002), .Z(n10139) );
  NOR U11390 ( .A(n13003), .B(n13001), .Z(n13002) );
  XOR U11391 ( .A(n13004), .B(n13005), .Z(n10142) );
  NOR U11392 ( .A(n13006), .B(n13004), .Z(n13005) );
  XOR U11393 ( .A(n13007), .B(n13008), .Z(n10145) );
  NOR U11394 ( .A(n13009), .B(n13007), .Z(n13008) );
  XOR U11395 ( .A(n13010), .B(n13011), .Z(n10148) );
  NOR U11396 ( .A(n13012), .B(n13010), .Z(n13011) );
  XOR U11397 ( .A(n13013), .B(n13014), .Z(n10151) );
  NOR U11398 ( .A(n13015), .B(n13013), .Z(n13014) );
  XOR U11399 ( .A(n13016), .B(n13017), .Z(n10154) );
  NOR U11400 ( .A(n13018), .B(n13016), .Z(n13017) );
  XOR U11401 ( .A(n13019), .B(n13020), .Z(n10157) );
  NOR U11402 ( .A(n13021), .B(n13019), .Z(n13020) );
  XOR U11403 ( .A(n13022), .B(n13023), .Z(n10160) );
  NOR U11404 ( .A(n13024), .B(n13022), .Z(n13023) );
  XOR U11405 ( .A(n13025), .B(n13026), .Z(n10163) );
  NOR U11406 ( .A(n13027), .B(n13025), .Z(n13026) );
  XOR U11407 ( .A(n13028), .B(n13029), .Z(n10166) );
  NOR U11408 ( .A(n13030), .B(n13028), .Z(n13029) );
  XOR U11409 ( .A(n13031), .B(n13032), .Z(n10169) );
  NOR U11410 ( .A(n13033), .B(n13031), .Z(n13032) );
  XOR U11411 ( .A(n13034), .B(n13035), .Z(n10172) );
  NOR U11412 ( .A(n13036), .B(n13034), .Z(n13035) );
  XOR U11413 ( .A(n13037), .B(n13038), .Z(n10175) );
  NOR U11414 ( .A(n13039), .B(n13037), .Z(n13038) );
  XOR U11415 ( .A(n13040), .B(n13041), .Z(n10178) );
  NOR U11416 ( .A(n13042), .B(n13040), .Z(n13041) );
  XOR U11417 ( .A(n13043), .B(n13044), .Z(n10181) );
  NOR U11418 ( .A(n13045), .B(n13043), .Z(n13044) );
  XOR U11419 ( .A(n13046), .B(n13047), .Z(n10184) );
  NOR U11420 ( .A(n13048), .B(n13046), .Z(n13047) );
  XOR U11421 ( .A(n13049), .B(n13050), .Z(n10187) );
  NOR U11422 ( .A(n13051), .B(n13049), .Z(n13050) );
  XOR U11423 ( .A(n13052), .B(n13053), .Z(n10190) );
  NOR U11424 ( .A(n13054), .B(n13052), .Z(n13053) );
  XOR U11425 ( .A(n13055), .B(n13056), .Z(n10193) );
  NOR U11426 ( .A(n13057), .B(n13055), .Z(n13056) );
  XOR U11427 ( .A(n13058), .B(n13059), .Z(n10196) );
  NOR U11428 ( .A(n13060), .B(n13058), .Z(n13059) );
  XOR U11429 ( .A(n13061), .B(n13062), .Z(n10199) );
  NOR U11430 ( .A(n13063), .B(n13061), .Z(n13062) );
  XOR U11431 ( .A(n13064), .B(n13065), .Z(n10202) );
  NOR U11432 ( .A(n13066), .B(n13064), .Z(n13065) );
  XOR U11433 ( .A(n13067), .B(n13068), .Z(n10205) );
  NOR U11434 ( .A(n13069), .B(n13067), .Z(n13068) );
  XOR U11435 ( .A(n13070), .B(n13071), .Z(n10208) );
  NOR U11436 ( .A(n13072), .B(n13070), .Z(n13071) );
  XOR U11437 ( .A(n13073), .B(n13074), .Z(n10211) );
  NOR U11438 ( .A(n13075), .B(n13073), .Z(n13074) );
  XOR U11439 ( .A(n13076), .B(n13077), .Z(n10214) );
  NOR U11440 ( .A(n13078), .B(n13076), .Z(n13077) );
  XOR U11441 ( .A(n13079), .B(n13080), .Z(n10217) );
  NOR U11442 ( .A(n13081), .B(n13079), .Z(n13080) );
  XOR U11443 ( .A(n13082), .B(n13083), .Z(n10220) );
  NOR U11444 ( .A(n13084), .B(n13082), .Z(n13083) );
  XOR U11445 ( .A(n13085), .B(n13086), .Z(n10223) );
  NOR U11446 ( .A(n13087), .B(n13085), .Z(n13086) );
  XOR U11447 ( .A(n13088), .B(n13089), .Z(n10226) );
  NOR U11448 ( .A(n13090), .B(n13088), .Z(n13089) );
  XOR U11449 ( .A(n13091), .B(n13092), .Z(n10229) );
  NOR U11450 ( .A(n13093), .B(n13091), .Z(n13092) );
  XOR U11451 ( .A(n13094), .B(n13095), .Z(n10232) );
  NOR U11452 ( .A(n13096), .B(n13094), .Z(n13095) );
  XOR U11453 ( .A(n13097), .B(n13098), .Z(n10235) );
  NOR U11454 ( .A(n13099), .B(n13097), .Z(n13098) );
  XOR U11455 ( .A(n13100), .B(n13101), .Z(n10238) );
  NOR U11456 ( .A(n13102), .B(n13100), .Z(n13101) );
  XOR U11457 ( .A(n13103), .B(n13104), .Z(n10241) );
  NOR U11458 ( .A(n13105), .B(n13103), .Z(n13104) );
  XOR U11459 ( .A(n13106), .B(n13107), .Z(n10244) );
  NOR U11460 ( .A(n13108), .B(n13106), .Z(n13107) );
  XOR U11461 ( .A(n13109), .B(n13110), .Z(n10247) );
  NOR U11462 ( .A(n13111), .B(n13109), .Z(n13110) );
  XOR U11463 ( .A(n13112), .B(n13113), .Z(n10250) );
  NOR U11464 ( .A(n13114), .B(n13112), .Z(n13113) );
  XOR U11465 ( .A(n13115), .B(n13116), .Z(n10253) );
  NOR U11466 ( .A(n13117), .B(n13115), .Z(n13116) );
  XOR U11467 ( .A(n13118), .B(n13119), .Z(n10256) );
  NOR U11468 ( .A(n13120), .B(n13118), .Z(n13119) );
  XOR U11469 ( .A(n13121), .B(n13122), .Z(n10259) );
  NOR U11470 ( .A(n13123), .B(n13121), .Z(n13122) );
  XOR U11471 ( .A(n13124), .B(n13125), .Z(n10262) );
  NOR U11472 ( .A(n13126), .B(n13124), .Z(n13125) );
  XOR U11473 ( .A(n13127), .B(n13128), .Z(n10265) );
  NOR U11474 ( .A(n13129), .B(n13127), .Z(n13128) );
  XOR U11475 ( .A(n13130), .B(n13131), .Z(n10268) );
  NOR U11476 ( .A(n13132), .B(n13130), .Z(n13131) );
  XOR U11477 ( .A(n13133), .B(n13134), .Z(n10271) );
  NOR U11478 ( .A(n13135), .B(n13133), .Z(n13134) );
  XOR U11479 ( .A(n13136), .B(n13137), .Z(n10274) );
  NOR U11480 ( .A(n13138), .B(n13136), .Z(n13137) );
  XOR U11481 ( .A(n13139), .B(n13140), .Z(n10277) );
  NOR U11482 ( .A(n13141), .B(n13139), .Z(n13140) );
  XOR U11483 ( .A(n13142), .B(n13143), .Z(n10280) );
  NOR U11484 ( .A(n13144), .B(n13142), .Z(n13143) );
  XOR U11485 ( .A(n13145), .B(n13146), .Z(n10283) );
  NOR U11486 ( .A(n13147), .B(n13145), .Z(n13146) );
  XOR U11487 ( .A(n13148), .B(n13149), .Z(n10286) );
  NOR U11488 ( .A(n13150), .B(n13148), .Z(n13149) );
  XOR U11489 ( .A(n13151), .B(n13152), .Z(n10289) );
  NOR U11490 ( .A(n13153), .B(n13151), .Z(n13152) );
  XOR U11491 ( .A(n13154), .B(n13155), .Z(n10292) );
  NOR U11492 ( .A(n13156), .B(n13154), .Z(n13155) );
  XOR U11493 ( .A(n13157), .B(n13158), .Z(n10295) );
  NOR U11494 ( .A(n13159), .B(n13157), .Z(n13158) );
  XOR U11495 ( .A(n13160), .B(n13161), .Z(n10298) );
  NOR U11496 ( .A(n13162), .B(n13160), .Z(n13161) );
  XOR U11497 ( .A(n13163), .B(n13164), .Z(n10301) );
  NOR U11498 ( .A(n13165), .B(n13163), .Z(n13164) );
  XOR U11499 ( .A(n13166), .B(n13167), .Z(n10304) );
  NOR U11500 ( .A(n13168), .B(n13166), .Z(n13167) );
  XOR U11501 ( .A(n13169), .B(n13170), .Z(n10307) );
  NOR U11502 ( .A(n13171), .B(n13169), .Z(n13170) );
  XOR U11503 ( .A(n13172), .B(n13173), .Z(n10310) );
  NOR U11504 ( .A(n13174), .B(n13172), .Z(n13173) );
  XOR U11505 ( .A(n13175), .B(n13176), .Z(n10313) );
  NOR U11506 ( .A(n13177), .B(n13175), .Z(n13176) );
  XOR U11507 ( .A(n13178), .B(n13179), .Z(n10316) );
  NOR U11508 ( .A(n13180), .B(n13178), .Z(n13179) );
  XOR U11509 ( .A(n13181), .B(n13182), .Z(n10319) );
  NOR U11510 ( .A(n13183), .B(n13181), .Z(n13182) );
  XOR U11511 ( .A(n13184), .B(n13185), .Z(n10322) );
  NOR U11512 ( .A(n13186), .B(n13184), .Z(n13185) );
  XOR U11513 ( .A(n13187), .B(n13188), .Z(n10325) );
  NOR U11514 ( .A(n13189), .B(n13187), .Z(n13188) );
  XOR U11515 ( .A(n13190), .B(n13191), .Z(n10328) );
  NOR U11516 ( .A(n13192), .B(n13190), .Z(n13191) );
  XOR U11517 ( .A(n13193), .B(n13194), .Z(n10331) );
  NOR U11518 ( .A(n13195), .B(n13193), .Z(n13194) );
  XOR U11519 ( .A(n13196), .B(n13197), .Z(n10334) );
  NOR U11520 ( .A(n13198), .B(n13196), .Z(n13197) );
  XOR U11521 ( .A(n13199), .B(n13200), .Z(n10337) );
  NOR U11522 ( .A(n13201), .B(n13199), .Z(n13200) );
  XOR U11523 ( .A(n13202), .B(n13203), .Z(n10340) );
  NOR U11524 ( .A(n13204), .B(n13202), .Z(n13203) );
  XOR U11525 ( .A(n13205), .B(n13206), .Z(n10343) );
  NOR U11526 ( .A(n13207), .B(n13205), .Z(n13206) );
  XOR U11527 ( .A(n13208), .B(n13209), .Z(n10346) );
  NOR U11528 ( .A(n13210), .B(n13208), .Z(n13209) );
  XOR U11529 ( .A(n13211), .B(n13212), .Z(n10349) );
  NOR U11530 ( .A(n13213), .B(n13211), .Z(n13212) );
  XOR U11531 ( .A(n13214), .B(n13215), .Z(n10352) );
  NOR U11532 ( .A(n13216), .B(n13214), .Z(n13215) );
  XOR U11533 ( .A(n13217), .B(n13218), .Z(n10355) );
  NOR U11534 ( .A(n13219), .B(n13217), .Z(n13218) );
  XOR U11535 ( .A(n13220), .B(n13221), .Z(n10358) );
  NOR U11536 ( .A(n13222), .B(n13220), .Z(n13221) );
  XOR U11537 ( .A(n13223), .B(n13224), .Z(n10361) );
  NOR U11538 ( .A(n13225), .B(n13223), .Z(n13224) );
  XOR U11539 ( .A(n13226), .B(n13227), .Z(n10364) );
  NOR U11540 ( .A(n13228), .B(n13226), .Z(n13227) );
  XOR U11541 ( .A(n13229), .B(n13230), .Z(n10367) );
  NOR U11542 ( .A(n13231), .B(n13229), .Z(n13230) );
  XOR U11543 ( .A(n13232), .B(n13233), .Z(n10370) );
  NOR U11544 ( .A(n13234), .B(n13232), .Z(n13233) );
  XOR U11545 ( .A(n13235), .B(n13236), .Z(n10373) );
  NOR U11546 ( .A(n13237), .B(n13235), .Z(n13236) );
  XOR U11547 ( .A(n13238), .B(n13239), .Z(n10376) );
  NOR U11548 ( .A(n13240), .B(n13238), .Z(n13239) );
  XOR U11549 ( .A(n13241), .B(n13242), .Z(n10379) );
  NOR U11550 ( .A(n13243), .B(n13241), .Z(n13242) );
  XOR U11551 ( .A(n13244), .B(n13245), .Z(n10382) );
  NOR U11552 ( .A(n13246), .B(n13244), .Z(n13245) );
  XOR U11553 ( .A(n13247), .B(n13248), .Z(n10385) );
  NOR U11554 ( .A(n13249), .B(n13247), .Z(n13248) );
  XOR U11555 ( .A(n13250), .B(n13251), .Z(n10388) );
  NOR U11556 ( .A(n13252), .B(n13250), .Z(n13251) );
  XOR U11557 ( .A(n13253), .B(n13254), .Z(n10391) );
  NOR U11558 ( .A(n13255), .B(n13253), .Z(n13254) );
  XOR U11559 ( .A(n13256), .B(n13257), .Z(n10394) );
  NOR U11560 ( .A(n13258), .B(n13256), .Z(n13257) );
  XOR U11561 ( .A(n13259), .B(n13260), .Z(n10397) );
  NOR U11562 ( .A(n13261), .B(n13259), .Z(n13260) );
  XOR U11563 ( .A(n13262), .B(n13263), .Z(n10400) );
  NOR U11564 ( .A(n13264), .B(n13262), .Z(n13263) );
  XOR U11565 ( .A(n13265), .B(n13266), .Z(n10403) );
  NOR U11566 ( .A(n13267), .B(n13265), .Z(n13266) );
  XOR U11567 ( .A(n13268), .B(n13269), .Z(n10406) );
  NOR U11568 ( .A(n13270), .B(n13268), .Z(n13269) );
  XOR U11569 ( .A(n13271), .B(n13272), .Z(n10409) );
  NOR U11570 ( .A(n13273), .B(n13271), .Z(n13272) );
  XOR U11571 ( .A(n13274), .B(n13275), .Z(n10412) );
  NOR U11572 ( .A(n13276), .B(n13274), .Z(n13275) );
  XOR U11573 ( .A(n13277), .B(n13278), .Z(n10415) );
  NOR U11574 ( .A(n13279), .B(n13277), .Z(n13278) );
  XOR U11575 ( .A(n13280), .B(n13281), .Z(n10418) );
  NOR U11576 ( .A(n13282), .B(n13280), .Z(n13281) );
  XOR U11577 ( .A(n13283), .B(n13284), .Z(n10421) );
  NOR U11578 ( .A(n13285), .B(n13283), .Z(n13284) );
  XOR U11579 ( .A(n13286), .B(n13287), .Z(n10424) );
  NOR U11580 ( .A(n13288), .B(n13286), .Z(n13287) );
  XOR U11581 ( .A(n13289), .B(n13290), .Z(n10427) );
  NOR U11582 ( .A(n13291), .B(n13289), .Z(n13290) );
  XOR U11583 ( .A(n13292), .B(n13293), .Z(n10430) );
  NOR U11584 ( .A(n13294), .B(n13292), .Z(n13293) );
  XOR U11585 ( .A(n13295), .B(n13296), .Z(n10433) );
  NOR U11586 ( .A(n13297), .B(n13295), .Z(n13296) );
  XOR U11587 ( .A(n13298), .B(n13299), .Z(n10436) );
  NOR U11588 ( .A(n13300), .B(n13298), .Z(n13299) );
  XOR U11589 ( .A(n13301), .B(n13302), .Z(n10439) );
  NOR U11590 ( .A(n13303), .B(n13301), .Z(n13302) );
  XOR U11591 ( .A(n13304), .B(n13305), .Z(n10442) );
  NOR U11592 ( .A(n13306), .B(n13304), .Z(n13305) );
  XOR U11593 ( .A(n13307), .B(n13308), .Z(n10445) );
  NOR U11594 ( .A(n13309), .B(n13307), .Z(n13308) );
  XOR U11595 ( .A(n13310), .B(n13311), .Z(n10448) );
  NOR U11596 ( .A(n13312), .B(n13310), .Z(n13311) );
  XOR U11597 ( .A(n13313), .B(n13314), .Z(n10451) );
  NOR U11598 ( .A(n13315), .B(n13313), .Z(n13314) );
  XOR U11599 ( .A(n13316), .B(n13317), .Z(n10454) );
  NOR U11600 ( .A(n13318), .B(n13316), .Z(n13317) );
  XOR U11601 ( .A(n13319), .B(n13320), .Z(n10457) );
  NOR U11602 ( .A(n13321), .B(n13319), .Z(n13320) );
  XOR U11603 ( .A(n13322), .B(n13323), .Z(n10460) );
  NOR U11604 ( .A(n13324), .B(n13322), .Z(n13323) );
  XOR U11605 ( .A(n13325), .B(n13326), .Z(n10463) );
  NOR U11606 ( .A(n13327), .B(n13325), .Z(n13326) );
  XOR U11607 ( .A(n13328), .B(n13329), .Z(n10466) );
  NOR U11608 ( .A(n13330), .B(n13328), .Z(n13329) );
  XOR U11609 ( .A(n13331), .B(n13332), .Z(n10469) );
  NOR U11610 ( .A(n13333), .B(n13331), .Z(n13332) );
  XOR U11611 ( .A(n13334), .B(n13335), .Z(n10472) );
  NOR U11612 ( .A(n13336), .B(n13334), .Z(n13335) );
  XOR U11613 ( .A(n13337), .B(n13338), .Z(n10475) );
  NOR U11614 ( .A(n13339), .B(n13337), .Z(n13338) );
  XOR U11615 ( .A(n13340), .B(n13341), .Z(n10478) );
  NOR U11616 ( .A(n13342), .B(n13340), .Z(n13341) );
  XOR U11617 ( .A(n13343), .B(n13344), .Z(n10481) );
  NOR U11618 ( .A(n13345), .B(n13343), .Z(n13344) );
  XOR U11619 ( .A(n13346), .B(n13347), .Z(n10484) );
  NOR U11620 ( .A(n13348), .B(n13346), .Z(n13347) );
  XOR U11621 ( .A(n13349), .B(n13350), .Z(n10487) );
  NOR U11622 ( .A(n13351), .B(n13349), .Z(n13350) );
  XOR U11623 ( .A(n13352), .B(n13353), .Z(n10490) );
  NOR U11624 ( .A(n13354), .B(n13352), .Z(n13353) );
  XOR U11625 ( .A(n13355), .B(n13356), .Z(n10493) );
  NOR U11626 ( .A(n13357), .B(n13355), .Z(n13356) );
  XOR U11627 ( .A(n13358), .B(n13359), .Z(n10496) );
  NOR U11628 ( .A(n13360), .B(n13358), .Z(n13359) );
  XOR U11629 ( .A(n13361), .B(n13362), .Z(n10499) );
  NOR U11630 ( .A(n13363), .B(n13361), .Z(n13362) );
  XOR U11631 ( .A(n13364), .B(n13365), .Z(n10502) );
  NOR U11632 ( .A(n13366), .B(n13364), .Z(n13365) );
  XOR U11633 ( .A(n13367), .B(n13368), .Z(n10505) );
  NOR U11634 ( .A(n13369), .B(n13367), .Z(n13368) );
  XOR U11635 ( .A(n13370), .B(n13371), .Z(n10508) );
  NOR U11636 ( .A(n13372), .B(n13370), .Z(n13371) );
  XOR U11637 ( .A(n13373), .B(n13374), .Z(n10511) );
  NOR U11638 ( .A(n13375), .B(n13373), .Z(n13374) );
  XOR U11639 ( .A(n13376), .B(n13377), .Z(n10514) );
  NOR U11640 ( .A(n13378), .B(n13376), .Z(n13377) );
  XOR U11641 ( .A(n13379), .B(n13380), .Z(n10517) );
  NOR U11642 ( .A(n13381), .B(n13379), .Z(n13380) );
  XOR U11643 ( .A(n13382), .B(n13383), .Z(n10520) );
  NOR U11644 ( .A(n13384), .B(n13382), .Z(n13383) );
  XOR U11645 ( .A(n13385), .B(n13386), .Z(n10523) );
  NOR U11646 ( .A(n13387), .B(n13385), .Z(n13386) );
  XOR U11647 ( .A(n13388), .B(n13389), .Z(n10526) );
  NOR U11648 ( .A(n13390), .B(n13388), .Z(n13389) );
  XOR U11649 ( .A(n13391), .B(n13392), .Z(n10529) );
  NOR U11650 ( .A(n13393), .B(n13391), .Z(n13392) );
  XOR U11651 ( .A(n13394), .B(n13395), .Z(n10532) );
  NOR U11652 ( .A(n13396), .B(n13394), .Z(n13395) );
  XOR U11653 ( .A(n13397), .B(n13398), .Z(n10535) );
  NOR U11654 ( .A(n13399), .B(n13397), .Z(n13398) );
  XOR U11655 ( .A(n13400), .B(n13401), .Z(n10538) );
  NOR U11656 ( .A(n13402), .B(n13400), .Z(n13401) );
  XOR U11657 ( .A(n13403), .B(n13404), .Z(n10541) );
  NOR U11658 ( .A(n13405), .B(n13403), .Z(n13404) );
  XOR U11659 ( .A(n13406), .B(n13407), .Z(n10544) );
  NOR U11660 ( .A(n13408), .B(n13406), .Z(n13407) );
  XOR U11661 ( .A(n13409), .B(n13410), .Z(n10547) );
  NOR U11662 ( .A(n13411), .B(n13409), .Z(n13410) );
  XOR U11663 ( .A(n13412), .B(n13413), .Z(n10550) );
  NOR U11664 ( .A(n13414), .B(n13412), .Z(n13413) );
  XOR U11665 ( .A(n13415), .B(n13416), .Z(n10553) );
  NOR U11666 ( .A(n13417), .B(n13415), .Z(n13416) );
  XOR U11667 ( .A(n13418), .B(n13419), .Z(n10556) );
  NOR U11668 ( .A(n13420), .B(n13418), .Z(n13419) );
  XOR U11669 ( .A(n13421), .B(n13422), .Z(n10559) );
  NOR U11670 ( .A(n13423), .B(n13421), .Z(n13422) );
  XOR U11671 ( .A(n13424), .B(n13425), .Z(n10562) );
  NOR U11672 ( .A(n13426), .B(n13424), .Z(n13425) );
  XOR U11673 ( .A(n13427), .B(n13428), .Z(n10565) );
  NOR U11674 ( .A(n13429), .B(n13427), .Z(n13428) );
  XOR U11675 ( .A(n13430), .B(n13431), .Z(n10568) );
  NOR U11676 ( .A(n13432), .B(n13430), .Z(n13431) );
  XOR U11677 ( .A(n13433), .B(n13434), .Z(n10571) );
  NOR U11678 ( .A(n13435), .B(n13433), .Z(n13434) );
  XOR U11679 ( .A(n13436), .B(n13437), .Z(n10574) );
  NOR U11680 ( .A(n13438), .B(n13436), .Z(n13437) );
  XOR U11681 ( .A(n13439), .B(n13440), .Z(n10577) );
  NOR U11682 ( .A(n13441), .B(n13439), .Z(n13440) );
  XOR U11683 ( .A(n13442), .B(n13443), .Z(n10580) );
  NOR U11684 ( .A(n13444), .B(n13442), .Z(n13443) );
  XOR U11685 ( .A(n13445), .B(n13446), .Z(n10583) );
  NOR U11686 ( .A(n13447), .B(n13445), .Z(n13446) );
  XOR U11687 ( .A(n13448), .B(n13449), .Z(n10586) );
  NOR U11688 ( .A(n13450), .B(n13448), .Z(n13449) );
  XOR U11689 ( .A(n13451), .B(n13452), .Z(n10589) );
  NOR U11690 ( .A(n13453), .B(n13451), .Z(n13452) );
  XOR U11691 ( .A(n13454), .B(n13455), .Z(n10592) );
  NOR U11692 ( .A(n13456), .B(n13454), .Z(n13455) );
  XOR U11693 ( .A(n13457), .B(n13458), .Z(n10595) );
  NOR U11694 ( .A(n13459), .B(n13457), .Z(n13458) );
  XOR U11695 ( .A(n13460), .B(n13461), .Z(n10598) );
  NOR U11696 ( .A(n13462), .B(n13460), .Z(n13461) );
  XOR U11697 ( .A(n13463), .B(n13464), .Z(n10601) );
  NOR U11698 ( .A(n13465), .B(n13463), .Z(n13464) );
  XOR U11699 ( .A(n13466), .B(n13467), .Z(n10604) );
  NOR U11700 ( .A(n13468), .B(n13466), .Z(n13467) );
  XOR U11701 ( .A(n13469), .B(n13470), .Z(n10607) );
  NOR U11702 ( .A(n13471), .B(n13469), .Z(n13470) );
  XOR U11703 ( .A(n13472), .B(n13473), .Z(n10610) );
  NOR U11704 ( .A(n13474), .B(n13472), .Z(n13473) );
  XOR U11705 ( .A(n13475), .B(n13476), .Z(n10613) );
  NOR U11706 ( .A(n13477), .B(n13475), .Z(n13476) );
  XOR U11707 ( .A(n13478), .B(n13479), .Z(n10616) );
  NOR U11708 ( .A(n13480), .B(n13478), .Z(n13479) );
  XOR U11709 ( .A(n13481), .B(n13482), .Z(n10619) );
  NOR U11710 ( .A(n13483), .B(n13481), .Z(n13482) );
  XOR U11711 ( .A(n13484), .B(n13485), .Z(n10622) );
  NOR U11712 ( .A(n13486), .B(n13484), .Z(n13485) );
  XOR U11713 ( .A(n13487), .B(n13488), .Z(n10625) );
  NOR U11714 ( .A(n13489), .B(n13487), .Z(n13488) );
  XOR U11715 ( .A(n13490), .B(n13491), .Z(n10628) );
  NOR U11716 ( .A(n13492), .B(n13490), .Z(n13491) );
  XOR U11717 ( .A(n13493), .B(n13494), .Z(n10631) );
  NOR U11718 ( .A(n13495), .B(n13493), .Z(n13494) );
  XOR U11719 ( .A(n13496), .B(n13497), .Z(n10634) );
  NOR U11720 ( .A(n13498), .B(n13496), .Z(n13497) );
  XOR U11721 ( .A(n13499), .B(n13500), .Z(n10637) );
  NOR U11722 ( .A(n13501), .B(n13499), .Z(n13500) );
  XOR U11723 ( .A(n13502), .B(n13503), .Z(n10640) );
  NOR U11724 ( .A(n13504), .B(n13502), .Z(n13503) );
  XOR U11725 ( .A(n13505), .B(n13506), .Z(n10643) );
  NOR U11726 ( .A(n13507), .B(n13505), .Z(n13506) );
  XOR U11727 ( .A(n13508), .B(n13509), .Z(n10646) );
  NOR U11728 ( .A(n13510), .B(n13508), .Z(n13509) );
  XOR U11729 ( .A(n13511), .B(n13512), .Z(n10649) );
  NOR U11730 ( .A(n13513), .B(n13511), .Z(n13512) );
  XOR U11731 ( .A(n13514), .B(n13515), .Z(n10652) );
  NOR U11732 ( .A(n13516), .B(n13514), .Z(n13515) );
  XOR U11733 ( .A(n13517), .B(n13518), .Z(n10655) );
  NOR U11734 ( .A(n13519), .B(n13517), .Z(n13518) );
  XOR U11735 ( .A(n13520), .B(n13521), .Z(n10658) );
  NOR U11736 ( .A(n13522), .B(n13520), .Z(n13521) );
  XOR U11737 ( .A(n13523), .B(n13524), .Z(n10661) );
  NOR U11738 ( .A(n13525), .B(n13523), .Z(n13524) );
  XOR U11739 ( .A(n13526), .B(n13527), .Z(n10664) );
  NOR U11740 ( .A(n13528), .B(n13526), .Z(n13527) );
  XOR U11741 ( .A(n13529), .B(n13530), .Z(n10667) );
  NOR U11742 ( .A(n13531), .B(n13529), .Z(n13530) );
  XOR U11743 ( .A(n13532), .B(n13533), .Z(n10670) );
  NOR U11744 ( .A(n13534), .B(n13532), .Z(n13533) );
  XOR U11745 ( .A(n13535), .B(n13536), .Z(n10673) );
  NOR U11746 ( .A(n13537), .B(n13535), .Z(n13536) );
  XOR U11747 ( .A(n13538), .B(n13539), .Z(n10676) );
  NOR U11748 ( .A(n13540), .B(n13538), .Z(n13539) );
  XOR U11749 ( .A(n13541), .B(n13542), .Z(n10679) );
  NOR U11750 ( .A(n13543), .B(n13541), .Z(n13542) );
  XOR U11751 ( .A(n13544), .B(n13545), .Z(n10682) );
  NOR U11752 ( .A(n13546), .B(n13544), .Z(n13545) );
  XOR U11753 ( .A(n13547), .B(n13548), .Z(n10685) );
  NOR U11754 ( .A(n13549), .B(n13547), .Z(n13548) );
  XOR U11755 ( .A(n13550), .B(n13551), .Z(n10688) );
  NOR U11756 ( .A(n13552), .B(n13550), .Z(n13551) );
  XOR U11757 ( .A(n13553), .B(n13554), .Z(n10691) );
  NOR U11758 ( .A(n13555), .B(n13553), .Z(n13554) );
  XOR U11759 ( .A(n13556), .B(n13557), .Z(n10694) );
  NOR U11760 ( .A(n13558), .B(n13556), .Z(n13557) );
  XOR U11761 ( .A(n13559), .B(n13560), .Z(n10697) );
  NOR U11762 ( .A(n13561), .B(n13559), .Z(n13560) );
  XOR U11763 ( .A(n13562), .B(n13563), .Z(n10700) );
  NOR U11764 ( .A(n13564), .B(n13562), .Z(n13563) );
  XOR U11765 ( .A(n13565), .B(n13566), .Z(n10703) );
  NOR U11766 ( .A(n13567), .B(n13565), .Z(n13566) );
  XOR U11767 ( .A(n13568), .B(n13569), .Z(n10706) );
  NOR U11768 ( .A(n13570), .B(n13568), .Z(n13569) );
  XOR U11769 ( .A(n13571), .B(n13572), .Z(n10709) );
  NOR U11770 ( .A(n13573), .B(n13571), .Z(n13572) );
  XOR U11771 ( .A(n13574), .B(n13575), .Z(n10712) );
  NOR U11772 ( .A(n13576), .B(n13574), .Z(n13575) );
  XOR U11773 ( .A(n13577), .B(n13578), .Z(n10715) );
  NOR U11774 ( .A(n13579), .B(n13577), .Z(n13578) );
  XOR U11775 ( .A(n13580), .B(n13581), .Z(n10718) );
  NOR U11776 ( .A(n13582), .B(n13580), .Z(n13581) );
  XOR U11777 ( .A(n13583), .B(n13584), .Z(n10721) );
  NOR U11778 ( .A(n13585), .B(n13583), .Z(n13584) );
  XOR U11779 ( .A(n13586), .B(n13587), .Z(n10724) );
  NOR U11780 ( .A(n13588), .B(n13586), .Z(n13587) );
  XOR U11781 ( .A(n13589), .B(n13590), .Z(n10727) );
  NOR U11782 ( .A(n13591), .B(n13589), .Z(n13590) );
  XOR U11783 ( .A(n13592), .B(n13593), .Z(n10730) );
  NOR U11784 ( .A(n13594), .B(n13592), .Z(n13593) );
  XOR U11785 ( .A(n13595), .B(n13596), .Z(n10733) );
  NOR U11786 ( .A(n13597), .B(n13595), .Z(n13596) );
  XOR U11787 ( .A(n13598), .B(n13599), .Z(n10736) );
  NOR U11788 ( .A(n13600), .B(n13598), .Z(n13599) );
  XOR U11789 ( .A(n13601), .B(n13602), .Z(n10739) );
  NOR U11790 ( .A(n13603), .B(n13601), .Z(n13602) );
  XOR U11791 ( .A(n13604), .B(n13605), .Z(n10742) );
  NOR U11792 ( .A(n13606), .B(n13604), .Z(n13605) );
  XOR U11793 ( .A(n13607), .B(n13608), .Z(n10745) );
  NOR U11794 ( .A(n13609), .B(n13607), .Z(n13608) );
  XOR U11795 ( .A(n13610), .B(n13611), .Z(n10748) );
  NOR U11796 ( .A(n13612), .B(n13610), .Z(n13611) );
  XOR U11797 ( .A(n13613), .B(n13614), .Z(n10751) );
  NOR U11798 ( .A(n13615), .B(n13613), .Z(n13614) );
  XOR U11799 ( .A(n13616), .B(n13617), .Z(n10754) );
  NOR U11800 ( .A(n13618), .B(n13616), .Z(n13617) );
  XOR U11801 ( .A(n13619), .B(n13620), .Z(n10757) );
  NOR U11802 ( .A(n13621), .B(n13619), .Z(n13620) );
  XOR U11803 ( .A(n13622), .B(n13623), .Z(n10760) );
  NOR U11804 ( .A(n13624), .B(n13622), .Z(n13623) );
  XOR U11805 ( .A(n13625), .B(n13626), .Z(n10763) );
  NOR U11806 ( .A(n13627), .B(n13625), .Z(n13626) );
  XOR U11807 ( .A(n13628), .B(n13629), .Z(n10766) );
  NOR U11808 ( .A(n13630), .B(n13628), .Z(n13629) );
  XOR U11809 ( .A(n13631), .B(n13632), .Z(n10769) );
  NOR U11810 ( .A(n13633), .B(n13631), .Z(n13632) );
  XOR U11811 ( .A(n13634), .B(n13635), .Z(n10772) );
  NOR U11812 ( .A(n13636), .B(n13634), .Z(n13635) );
  XOR U11813 ( .A(n13637), .B(n13638), .Z(n10775) );
  NOR U11814 ( .A(n13639), .B(n13637), .Z(n13638) );
  XOR U11815 ( .A(n13640), .B(n13641), .Z(n10778) );
  NOR U11816 ( .A(n13642), .B(n13640), .Z(n13641) );
  XOR U11817 ( .A(n13643), .B(n13644), .Z(n10781) );
  NOR U11818 ( .A(n13645), .B(n13643), .Z(n13644) );
  XOR U11819 ( .A(n13646), .B(n13647), .Z(n10784) );
  NOR U11820 ( .A(n13648), .B(n13646), .Z(n13647) );
  XOR U11821 ( .A(n13649), .B(n13650), .Z(n10787) );
  NOR U11822 ( .A(n13651), .B(n13649), .Z(n13650) );
  XOR U11823 ( .A(n13652), .B(n13653), .Z(n10790) );
  NOR U11824 ( .A(n13654), .B(n13652), .Z(n13653) );
  XOR U11825 ( .A(n13655), .B(n13656), .Z(n10793) );
  NOR U11826 ( .A(n13657), .B(n13655), .Z(n13656) );
  XOR U11827 ( .A(n13658), .B(n13659), .Z(n10796) );
  NOR U11828 ( .A(n13660), .B(n13658), .Z(n13659) );
  XOR U11829 ( .A(n13661), .B(n13662), .Z(n10799) );
  NOR U11830 ( .A(n13663), .B(n13661), .Z(n13662) );
  XOR U11831 ( .A(n13664), .B(n13665), .Z(n10802) );
  NOR U11832 ( .A(n13666), .B(n13664), .Z(n13665) );
  XOR U11833 ( .A(n13667), .B(n13668), .Z(n10805) );
  NOR U11834 ( .A(n13669), .B(n13667), .Z(n13668) );
  XOR U11835 ( .A(n13670), .B(n13671), .Z(n10808) );
  NOR U11836 ( .A(n13672), .B(n13670), .Z(n13671) );
  XOR U11837 ( .A(n13673), .B(n13674), .Z(n10811) );
  NOR U11838 ( .A(n13675), .B(n13673), .Z(n13674) );
  XOR U11839 ( .A(n13676), .B(n13677), .Z(n10814) );
  NOR U11840 ( .A(n13678), .B(n13676), .Z(n13677) );
  XOR U11841 ( .A(n13679), .B(n13680), .Z(n10817) );
  NOR U11842 ( .A(n13681), .B(n13679), .Z(n13680) );
  XOR U11843 ( .A(n13682), .B(n13683), .Z(n10820) );
  NOR U11844 ( .A(n13684), .B(n13682), .Z(n13683) );
  XOR U11845 ( .A(n13685), .B(n13686), .Z(n10823) );
  NOR U11846 ( .A(n13687), .B(n13685), .Z(n13686) );
  XOR U11847 ( .A(n13688), .B(n13689), .Z(n10826) );
  NOR U11848 ( .A(n13690), .B(n13688), .Z(n13689) );
  XOR U11849 ( .A(n13691), .B(n13692), .Z(n10829) );
  NOR U11850 ( .A(n13693), .B(n13691), .Z(n13692) );
  XOR U11851 ( .A(n13694), .B(n13695), .Z(n10832) );
  NOR U11852 ( .A(n13696), .B(n13694), .Z(n13695) );
  XOR U11853 ( .A(n13697), .B(n13698), .Z(n10835) );
  NOR U11854 ( .A(n13699), .B(n13697), .Z(n13698) );
  XOR U11855 ( .A(n13700), .B(n13701), .Z(n10838) );
  NOR U11856 ( .A(n13702), .B(n13700), .Z(n13701) );
  XOR U11857 ( .A(n13703), .B(n13704), .Z(n10841) );
  NOR U11858 ( .A(n13705), .B(n13703), .Z(n13704) );
  XOR U11859 ( .A(n13706), .B(n13707), .Z(n10844) );
  NOR U11860 ( .A(n13708), .B(n13706), .Z(n13707) );
  XOR U11861 ( .A(n13709), .B(n13710), .Z(n10847) );
  NOR U11862 ( .A(n13711), .B(n13709), .Z(n13710) );
  XOR U11863 ( .A(n13712), .B(n13713), .Z(n10850) );
  NOR U11864 ( .A(n13714), .B(n13712), .Z(n13713) );
  XOR U11865 ( .A(n13715), .B(n13716), .Z(n10853) );
  NOR U11866 ( .A(n13717), .B(n13715), .Z(n13716) );
  XOR U11867 ( .A(n13718), .B(n13719), .Z(n10856) );
  NOR U11868 ( .A(n13720), .B(n13718), .Z(n13719) );
  XOR U11869 ( .A(n13721), .B(n13722), .Z(n10859) );
  NOR U11870 ( .A(n13723), .B(n13721), .Z(n13722) );
  XOR U11871 ( .A(n13724), .B(n13725), .Z(n10862) );
  NOR U11872 ( .A(n13726), .B(n13724), .Z(n13725) );
  XOR U11873 ( .A(n13727), .B(n13728), .Z(n10865) );
  NOR U11874 ( .A(n13729), .B(n13727), .Z(n13728) );
  XOR U11875 ( .A(n13730), .B(n13731), .Z(n10868) );
  NOR U11876 ( .A(n13732), .B(n13730), .Z(n13731) );
  XOR U11877 ( .A(n13733), .B(n13734), .Z(n10871) );
  NOR U11878 ( .A(n13735), .B(n13733), .Z(n13734) );
  XOR U11879 ( .A(n13736), .B(n13737), .Z(n10874) );
  NOR U11880 ( .A(n13738), .B(n13736), .Z(n13737) );
  XOR U11881 ( .A(n13739), .B(n13740), .Z(n10877) );
  NOR U11882 ( .A(n13741), .B(n13739), .Z(n13740) );
  XOR U11883 ( .A(n13742), .B(n13743), .Z(n10880) );
  NOR U11884 ( .A(n13744), .B(n13742), .Z(n13743) );
  XOR U11885 ( .A(n13745), .B(n13746), .Z(n10883) );
  NOR U11886 ( .A(n13747), .B(n13745), .Z(n13746) );
  XOR U11887 ( .A(n13748), .B(n13749), .Z(n10886) );
  NOR U11888 ( .A(n13750), .B(n13748), .Z(n13749) );
  XOR U11889 ( .A(n13751), .B(n13752), .Z(n10889) );
  NOR U11890 ( .A(n13753), .B(n13751), .Z(n13752) );
  XOR U11891 ( .A(n13754), .B(n13755), .Z(n10892) );
  NOR U11892 ( .A(n13756), .B(n13754), .Z(n13755) );
  XOR U11893 ( .A(n13757), .B(n13758), .Z(n10895) );
  NOR U11894 ( .A(n13759), .B(n13757), .Z(n13758) );
  XOR U11895 ( .A(n13760), .B(n13761), .Z(n10898) );
  NOR U11896 ( .A(n13762), .B(n13760), .Z(n13761) );
  XOR U11897 ( .A(n13763), .B(n13764), .Z(n10901) );
  NOR U11898 ( .A(n13765), .B(n13763), .Z(n13764) );
  XOR U11899 ( .A(n13766), .B(n13767), .Z(n10904) );
  NOR U11900 ( .A(n13768), .B(n13766), .Z(n13767) );
  XOR U11901 ( .A(n13769), .B(n13770), .Z(n10907) );
  NOR U11902 ( .A(n13771), .B(n13769), .Z(n13770) );
  XOR U11903 ( .A(n13772), .B(n13773), .Z(n10910) );
  NOR U11904 ( .A(n13774), .B(n13772), .Z(n13773) );
  XOR U11905 ( .A(n13775), .B(n13776), .Z(n10913) );
  NOR U11906 ( .A(n13777), .B(n13775), .Z(n13776) );
  XOR U11907 ( .A(n13778), .B(n13779), .Z(n10916) );
  NOR U11908 ( .A(n13780), .B(n13778), .Z(n13779) );
  XOR U11909 ( .A(n13781), .B(n13782), .Z(n10919) );
  NOR U11910 ( .A(n13783), .B(n13781), .Z(n13782) );
  XOR U11911 ( .A(n13784), .B(n13785), .Z(n10922) );
  NOR U11912 ( .A(n13786), .B(n13784), .Z(n13785) );
  XOR U11913 ( .A(n13787), .B(n13788), .Z(n10925) );
  NOR U11914 ( .A(n13789), .B(n13787), .Z(n13788) );
  XOR U11915 ( .A(n13790), .B(n13791), .Z(n10928) );
  NOR U11916 ( .A(n13792), .B(n13790), .Z(n13791) );
  XOR U11917 ( .A(n13793), .B(n13794), .Z(n10931) );
  NOR U11918 ( .A(n13795), .B(n13793), .Z(n13794) );
  XOR U11919 ( .A(n13796), .B(n13797), .Z(n10934) );
  NOR U11920 ( .A(n13798), .B(n13796), .Z(n13797) );
  XOR U11921 ( .A(n13799), .B(n13800), .Z(n10937) );
  NOR U11922 ( .A(n13801), .B(n13799), .Z(n13800) );
  XOR U11923 ( .A(n13802), .B(n13803), .Z(n10940) );
  NOR U11924 ( .A(n13804), .B(n13802), .Z(n13803) );
  XOR U11925 ( .A(n13805), .B(n13806), .Z(n10943) );
  NOR U11926 ( .A(n13807), .B(n13805), .Z(n13806) );
  XOR U11927 ( .A(n13808), .B(n13809), .Z(n10946) );
  NOR U11928 ( .A(n13810), .B(n13808), .Z(n13809) );
  XOR U11929 ( .A(n13811), .B(n13812), .Z(n10949) );
  NOR U11930 ( .A(n13813), .B(n13811), .Z(n13812) );
  XOR U11931 ( .A(n13814), .B(n13815), .Z(n10952) );
  NOR U11932 ( .A(n13816), .B(n13814), .Z(n13815) );
  XOR U11933 ( .A(n13817), .B(n13818), .Z(n10955) );
  NOR U11934 ( .A(n13819), .B(n13817), .Z(n13818) );
  XOR U11935 ( .A(n13820), .B(n13821), .Z(n10958) );
  NOR U11936 ( .A(n13822), .B(n13820), .Z(n13821) );
  XOR U11937 ( .A(n13823), .B(n13824), .Z(n10961) );
  NOR U11938 ( .A(n13825), .B(n13823), .Z(n13824) );
  XOR U11939 ( .A(n13826), .B(n13827), .Z(n10964) );
  NOR U11940 ( .A(n13828), .B(n13826), .Z(n13827) );
  XOR U11941 ( .A(n13829), .B(n13830), .Z(n10967) );
  NOR U11942 ( .A(n13831), .B(n13829), .Z(n13830) );
  XOR U11943 ( .A(n13832), .B(n13833), .Z(n10970) );
  NOR U11944 ( .A(n13834), .B(n13832), .Z(n13833) );
  XOR U11945 ( .A(n13835), .B(n13836), .Z(n10973) );
  NOR U11946 ( .A(n13837), .B(n13835), .Z(n13836) );
  XOR U11947 ( .A(n13838), .B(n13839), .Z(n10976) );
  NOR U11948 ( .A(n13840), .B(n13838), .Z(n13839) );
  XOR U11949 ( .A(n13841), .B(n13842), .Z(n10979) );
  NOR U11950 ( .A(n13843), .B(n13841), .Z(n13842) );
  XOR U11951 ( .A(n13844), .B(n13845), .Z(n10982) );
  NOR U11952 ( .A(n13846), .B(n13844), .Z(n13845) );
  XOR U11953 ( .A(n13847), .B(n13848), .Z(n10985) );
  NOR U11954 ( .A(n13849), .B(n13847), .Z(n13848) );
  XOR U11955 ( .A(n13850), .B(n13851), .Z(n10988) );
  NOR U11956 ( .A(n13852), .B(n13850), .Z(n13851) );
  XOR U11957 ( .A(n13853), .B(n13854), .Z(n10991) );
  NOR U11958 ( .A(n13855), .B(n13853), .Z(n13854) );
  XOR U11959 ( .A(n13856), .B(n13857), .Z(n10994) );
  NOR U11960 ( .A(n13858), .B(n13856), .Z(n13857) );
  XOR U11961 ( .A(n13859), .B(n13860), .Z(n10997) );
  NOR U11962 ( .A(n13861), .B(n13859), .Z(n13860) );
  XOR U11963 ( .A(n13862), .B(n13863), .Z(n11000) );
  NOR U11964 ( .A(n13864), .B(n13862), .Z(n13863) );
  XOR U11965 ( .A(n13865), .B(n13866), .Z(n11003) );
  NOR U11966 ( .A(n13867), .B(n13865), .Z(n13866) );
  XOR U11967 ( .A(n13868), .B(n13869), .Z(n11006) );
  NOR U11968 ( .A(n13870), .B(n13868), .Z(n13869) );
  XOR U11969 ( .A(n13871), .B(n13872), .Z(n11009) );
  NOR U11970 ( .A(n13873), .B(n13871), .Z(n13872) );
  XOR U11971 ( .A(n13874), .B(n13875), .Z(n11012) );
  NOR U11972 ( .A(n13876), .B(n13874), .Z(n13875) );
  XOR U11973 ( .A(n13877), .B(n13878), .Z(n11015) );
  NOR U11974 ( .A(n13879), .B(n13877), .Z(n13878) );
  XOR U11975 ( .A(n13880), .B(n13881), .Z(n11018) );
  NOR U11976 ( .A(n13882), .B(n13880), .Z(n13881) );
  XOR U11977 ( .A(n13883), .B(n13884), .Z(n11021) );
  NOR U11978 ( .A(n13885), .B(n13883), .Z(n13884) );
  XOR U11979 ( .A(n13886), .B(n13887), .Z(n11024) );
  NOR U11980 ( .A(n13888), .B(n13886), .Z(n13887) );
  XOR U11981 ( .A(n13889), .B(n13890), .Z(n11027) );
  NOR U11982 ( .A(n13891), .B(n13889), .Z(n13890) );
  XOR U11983 ( .A(n13892), .B(n13893), .Z(n11030) );
  NOR U11984 ( .A(n13894), .B(n13892), .Z(n13893) );
  XOR U11985 ( .A(n13895), .B(n13896), .Z(n11033) );
  NOR U11986 ( .A(n13897), .B(n13895), .Z(n13896) );
  XOR U11987 ( .A(n13898), .B(n13899), .Z(n11036) );
  NOR U11988 ( .A(n13900), .B(n13898), .Z(n13899) );
  XOR U11989 ( .A(n13901), .B(n13902), .Z(n11039) );
  NOR U11990 ( .A(n13903), .B(n13901), .Z(n13902) );
  XOR U11991 ( .A(n13904), .B(n13905), .Z(n11042) );
  NOR U11992 ( .A(n13906), .B(n13904), .Z(n13905) );
  XOR U11993 ( .A(n13907), .B(n13908), .Z(n11045) );
  NOR U11994 ( .A(n13909), .B(n13907), .Z(n13908) );
  XOR U11995 ( .A(n13910), .B(n13911), .Z(n11048) );
  NOR U11996 ( .A(n13912), .B(n13910), .Z(n13911) );
  XOR U11997 ( .A(n13913), .B(n13914), .Z(n11051) );
  NOR U11998 ( .A(n13915), .B(n13913), .Z(n13914) );
  XOR U11999 ( .A(n13916), .B(n13917), .Z(n11054) );
  NOR U12000 ( .A(n13918), .B(n13916), .Z(n13917) );
  XOR U12001 ( .A(n13919), .B(n13920), .Z(n11057) );
  NOR U12002 ( .A(n13921), .B(n13919), .Z(n13920) );
  XOR U12003 ( .A(n13922), .B(n13923), .Z(n11060) );
  NOR U12004 ( .A(n13924), .B(n13922), .Z(n13923) );
  XOR U12005 ( .A(n13925), .B(n13926), .Z(n11063) );
  NOR U12006 ( .A(n13927), .B(n13925), .Z(n13926) );
  XOR U12007 ( .A(n13928), .B(n13929), .Z(n11066) );
  NOR U12008 ( .A(n13930), .B(n13928), .Z(n13929) );
  XOR U12009 ( .A(n13931), .B(n13932), .Z(n11069) );
  NOR U12010 ( .A(n13933), .B(n13931), .Z(n13932) );
  XOR U12011 ( .A(n13934), .B(n13935), .Z(n11072) );
  NOR U12012 ( .A(n13936), .B(n13934), .Z(n13935) );
  XOR U12013 ( .A(n13937), .B(n13938), .Z(n11075) );
  NOR U12014 ( .A(n13939), .B(n13937), .Z(n13938) );
  XOR U12015 ( .A(n13940), .B(n13941), .Z(n11078) );
  NOR U12016 ( .A(n13942), .B(n13940), .Z(n13941) );
  XOR U12017 ( .A(n13943), .B(n13944), .Z(n11081) );
  NOR U12018 ( .A(n13945), .B(n13943), .Z(n13944) );
  XOR U12019 ( .A(n13946), .B(n13947), .Z(n11084) );
  NOR U12020 ( .A(n13948), .B(n13946), .Z(n13947) );
  XOR U12021 ( .A(n13949), .B(n13950), .Z(n11087) );
  NOR U12022 ( .A(n13951), .B(n13949), .Z(n13950) );
  XOR U12023 ( .A(n13952), .B(n13953), .Z(n11090) );
  NOR U12024 ( .A(n13954), .B(n13952), .Z(n13953) );
  XOR U12025 ( .A(n13955), .B(n13956), .Z(n11093) );
  NOR U12026 ( .A(n13957), .B(n13955), .Z(n13956) );
  XOR U12027 ( .A(n13958), .B(n13959), .Z(n11096) );
  NOR U12028 ( .A(n13960), .B(n13958), .Z(n13959) );
  XOR U12029 ( .A(n13961), .B(n13962), .Z(n11099) );
  NOR U12030 ( .A(n13963), .B(n13961), .Z(n13962) );
  XOR U12031 ( .A(n13964), .B(n13965), .Z(n11102) );
  NOR U12032 ( .A(n13966), .B(n13964), .Z(n13965) );
  XOR U12033 ( .A(n13967), .B(n13968), .Z(n11105) );
  NOR U12034 ( .A(n13969), .B(n13967), .Z(n13968) );
  XOR U12035 ( .A(n13970), .B(n13971), .Z(n11108) );
  NOR U12036 ( .A(n13972), .B(n13970), .Z(n13971) );
  XOR U12037 ( .A(n13973), .B(n13974), .Z(n11111) );
  NOR U12038 ( .A(n13975), .B(n13973), .Z(n13974) );
  XOR U12039 ( .A(n13976), .B(n13977), .Z(n11114) );
  NOR U12040 ( .A(n13978), .B(n13976), .Z(n13977) );
  XOR U12041 ( .A(n13979), .B(n13980), .Z(n11117) );
  NOR U12042 ( .A(n13981), .B(n13979), .Z(n13980) );
  XOR U12043 ( .A(n13982), .B(n13983), .Z(n11120) );
  NOR U12044 ( .A(n13984), .B(n13982), .Z(n13983) );
  XOR U12045 ( .A(n13985), .B(n13986), .Z(n11123) );
  NOR U12046 ( .A(n13987), .B(n13985), .Z(n13986) );
  XOR U12047 ( .A(n13988), .B(n13989), .Z(n11126) );
  NOR U12048 ( .A(n13990), .B(n13988), .Z(n13989) );
  XOR U12049 ( .A(n13991), .B(n13992), .Z(n11129) );
  NOR U12050 ( .A(n13993), .B(n13991), .Z(n13992) );
  XOR U12051 ( .A(n13994), .B(n13995), .Z(n11132) );
  NOR U12052 ( .A(n13996), .B(n13994), .Z(n13995) );
  XOR U12053 ( .A(n13997), .B(n13998), .Z(n11135) );
  NOR U12054 ( .A(n13999), .B(n13997), .Z(n13998) );
  XOR U12055 ( .A(n14000), .B(n14001), .Z(n11138) );
  NOR U12056 ( .A(n14002), .B(n14000), .Z(n14001) );
  XOR U12057 ( .A(n14003), .B(n14004), .Z(n11141) );
  NOR U12058 ( .A(n14005), .B(n14003), .Z(n14004) );
  XOR U12059 ( .A(n14006), .B(n14007), .Z(n11144) );
  NOR U12060 ( .A(n14008), .B(n14006), .Z(n14007) );
  XOR U12061 ( .A(n14009), .B(n14010), .Z(n11147) );
  NOR U12062 ( .A(n14011), .B(n14009), .Z(n14010) );
  XOR U12063 ( .A(n14012), .B(n14013), .Z(n11150) );
  NOR U12064 ( .A(n14014), .B(n14012), .Z(n14013) );
  XOR U12065 ( .A(n14015), .B(n14016), .Z(n11153) );
  NOR U12066 ( .A(n14017), .B(n14015), .Z(n14016) );
  XOR U12067 ( .A(n14018), .B(n14019), .Z(n11156) );
  NOR U12068 ( .A(n14020), .B(n14018), .Z(n14019) );
  XOR U12069 ( .A(n14021), .B(n14022), .Z(n11159) );
  NOR U12070 ( .A(n14023), .B(n14021), .Z(n14022) );
  XOR U12071 ( .A(n14024), .B(n14025), .Z(n11162) );
  NOR U12072 ( .A(n14026), .B(n14024), .Z(n14025) );
  XOR U12073 ( .A(n14027), .B(n14028), .Z(n11165) );
  NOR U12074 ( .A(n14029), .B(n14027), .Z(n14028) );
  XOR U12075 ( .A(n14030), .B(n14031), .Z(n11168) );
  NOR U12076 ( .A(n14032), .B(n14030), .Z(n14031) );
  XOR U12077 ( .A(n14033), .B(n14034), .Z(n11171) );
  NOR U12078 ( .A(n14035), .B(n14033), .Z(n14034) );
  XOR U12079 ( .A(n14036), .B(n14037), .Z(n11174) );
  NOR U12080 ( .A(n14038), .B(n14036), .Z(n14037) );
  XOR U12081 ( .A(n14039), .B(n14040), .Z(n11177) );
  NOR U12082 ( .A(n14041), .B(n14039), .Z(n14040) );
  XOR U12083 ( .A(n14042), .B(n14043), .Z(n11180) );
  NOR U12084 ( .A(n14044), .B(n14042), .Z(n14043) );
  XOR U12085 ( .A(n14045), .B(n14046), .Z(n11183) );
  NOR U12086 ( .A(n14047), .B(n14045), .Z(n14046) );
  XOR U12087 ( .A(n14048), .B(n14049), .Z(n11186) );
  NOR U12088 ( .A(n14050), .B(n14048), .Z(n14049) );
  XOR U12089 ( .A(n14051), .B(n14052), .Z(n11189) );
  NOR U12090 ( .A(n14053), .B(n14051), .Z(n14052) );
  XOR U12091 ( .A(n14054), .B(n14055), .Z(n11192) );
  NOR U12092 ( .A(n14056), .B(n14054), .Z(n14055) );
  XOR U12093 ( .A(n14057), .B(n14058), .Z(n11195) );
  NOR U12094 ( .A(n14059), .B(n14057), .Z(n14058) );
  XOR U12095 ( .A(n14060), .B(n14061), .Z(n11198) );
  NOR U12096 ( .A(n14062), .B(n14060), .Z(n14061) );
  XOR U12097 ( .A(n14063), .B(n14064), .Z(n11201) );
  NOR U12098 ( .A(n14065), .B(n14063), .Z(n14064) );
  XOR U12099 ( .A(n14066), .B(n14067), .Z(n11204) );
  NOR U12100 ( .A(n14068), .B(n14066), .Z(n14067) );
  XOR U12101 ( .A(n14069), .B(n14070), .Z(n11207) );
  NOR U12102 ( .A(n14071), .B(n14069), .Z(n14070) );
  XOR U12103 ( .A(n14072), .B(n14073), .Z(n11210) );
  NOR U12104 ( .A(n14074), .B(n14072), .Z(n14073) );
  XOR U12105 ( .A(n14075), .B(n14076), .Z(n11213) );
  NOR U12106 ( .A(n14077), .B(n14075), .Z(n14076) );
  XOR U12107 ( .A(n14078), .B(n14079), .Z(n11216) );
  NOR U12108 ( .A(n14080), .B(n14078), .Z(n14079) );
  XOR U12109 ( .A(n14081), .B(n14082), .Z(n11219) );
  NOR U12110 ( .A(n14083), .B(n14081), .Z(n14082) );
  XOR U12111 ( .A(n14084), .B(n14085), .Z(n11222) );
  NOR U12112 ( .A(n14086), .B(n14084), .Z(n14085) );
  XOR U12113 ( .A(n14087), .B(n14088), .Z(n11225) );
  NOR U12114 ( .A(n14089), .B(n14087), .Z(n14088) );
  XOR U12115 ( .A(n14090), .B(n14091), .Z(n11228) );
  NOR U12116 ( .A(n14092), .B(n14090), .Z(n14091) );
  XOR U12117 ( .A(n14093), .B(n14094), .Z(n11231) );
  NOR U12118 ( .A(n14095), .B(n14093), .Z(n14094) );
  XOR U12119 ( .A(n14096), .B(n14097), .Z(n11234) );
  NOR U12120 ( .A(n14098), .B(n14096), .Z(n14097) );
  XOR U12121 ( .A(n14099), .B(n14100), .Z(n11237) );
  NOR U12122 ( .A(n14101), .B(n14099), .Z(n14100) );
  XOR U12123 ( .A(n14102), .B(n14103), .Z(n11240) );
  NOR U12124 ( .A(n14104), .B(n14102), .Z(n14103) );
  XOR U12125 ( .A(n14105), .B(n14106), .Z(n11243) );
  NOR U12126 ( .A(n14107), .B(n14105), .Z(n14106) );
  XOR U12127 ( .A(n14108), .B(n14109), .Z(n11246) );
  NOR U12128 ( .A(n14110), .B(n14108), .Z(n14109) );
  XOR U12129 ( .A(n14111), .B(n14112), .Z(n11249) );
  NOR U12130 ( .A(n14113), .B(n14111), .Z(n14112) );
  XOR U12131 ( .A(n14114), .B(n14115), .Z(n11252) );
  NOR U12132 ( .A(n14116), .B(n14114), .Z(n14115) );
  XOR U12133 ( .A(n14117), .B(n14118), .Z(n11255) );
  NOR U12134 ( .A(n14119), .B(n14117), .Z(n14118) );
  XOR U12135 ( .A(n14120), .B(n14121), .Z(n11258) );
  NOR U12136 ( .A(n14122), .B(n14120), .Z(n14121) );
  XOR U12137 ( .A(n14123), .B(n14124), .Z(n11261) );
  NOR U12138 ( .A(n14125), .B(n14123), .Z(n14124) );
  XOR U12139 ( .A(n14126), .B(n14127), .Z(n11264) );
  NOR U12140 ( .A(n14128), .B(n14126), .Z(n14127) );
  XOR U12141 ( .A(n14129), .B(n14130), .Z(n11267) );
  NOR U12142 ( .A(n14131), .B(n14129), .Z(n14130) );
  XOR U12143 ( .A(n14132), .B(n14133), .Z(n11270) );
  NOR U12144 ( .A(n14134), .B(n14132), .Z(n14133) );
  XOR U12145 ( .A(n14135), .B(n14136), .Z(n11273) );
  NOR U12146 ( .A(n14137), .B(n14135), .Z(n14136) );
  XOR U12147 ( .A(n14138), .B(n14139), .Z(n11276) );
  NOR U12148 ( .A(n14140), .B(n14138), .Z(n14139) );
  XOR U12149 ( .A(n14141), .B(n14142), .Z(n11279) );
  NOR U12150 ( .A(n14143), .B(n14141), .Z(n14142) );
  XOR U12151 ( .A(n14144), .B(n14145), .Z(n11282) );
  NOR U12152 ( .A(n14146), .B(n14144), .Z(n14145) );
  XOR U12153 ( .A(n14147), .B(n14148), .Z(n11285) );
  NOR U12154 ( .A(n14149), .B(n14147), .Z(n14148) );
  XOR U12155 ( .A(n14150), .B(n14151), .Z(n11288) );
  NOR U12156 ( .A(n14152), .B(n14150), .Z(n14151) );
  XOR U12157 ( .A(n14153), .B(n14154), .Z(n11291) );
  NOR U12158 ( .A(n14155), .B(n14153), .Z(n14154) );
  XOR U12159 ( .A(n14156), .B(n14157), .Z(n11294) );
  NOR U12160 ( .A(n14158), .B(n14156), .Z(n14157) );
  XOR U12161 ( .A(n14159), .B(n14160), .Z(n11297) );
  NOR U12162 ( .A(n14161), .B(n14159), .Z(n14160) );
  XOR U12163 ( .A(n14162), .B(n14163), .Z(n11300) );
  NOR U12164 ( .A(n14164), .B(n14162), .Z(n14163) );
  XOR U12165 ( .A(n14165), .B(n14166), .Z(n11303) );
  NOR U12166 ( .A(n102), .B(n14167), .Z(n14166) );
  IV U12167 ( .A(n14165), .Z(n14167) );
  XOR U12168 ( .A(n14168), .B(n14169), .Z(n11306) );
  AND U12169 ( .A(n14170), .B(n14171), .Z(n14169) );
  XOR U12170 ( .A(n14168), .B(n104), .Z(n14171) );
  XOR U12171 ( .A(n12736), .B(n12735), .Z(n104) );
  XNOR U12172 ( .A(n12733), .B(n12732), .Z(n12735) );
  XNOR U12173 ( .A(n12730), .B(n12729), .Z(n12732) );
  XNOR U12174 ( .A(n12727), .B(n12726), .Z(n12729) );
  XNOR U12175 ( .A(n12724), .B(n12723), .Z(n12726) );
  XNOR U12176 ( .A(n12721), .B(n12720), .Z(n12723) );
  XNOR U12177 ( .A(n12718), .B(n12717), .Z(n12720) );
  XNOR U12178 ( .A(n12715), .B(n12714), .Z(n12717) );
  XNOR U12179 ( .A(n12712), .B(n12711), .Z(n12714) );
  XNOR U12180 ( .A(n12709), .B(n12708), .Z(n12711) );
  XNOR U12181 ( .A(n12706), .B(n12705), .Z(n12708) );
  XNOR U12182 ( .A(n12703), .B(n12702), .Z(n12705) );
  XNOR U12183 ( .A(n12700), .B(n12699), .Z(n12702) );
  XNOR U12184 ( .A(n12697), .B(n12696), .Z(n12699) );
  XNOR U12185 ( .A(n12694), .B(n12693), .Z(n12696) );
  XNOR U12186 ( .A(n12691), .B(n12690), .Z(n12693) );
  XNOR U12187 ( .A(n12688), .B(n12687), .Z(n12690) );
  XNOR U12188 ( .A(n12685), .B(n12684), .Z(n12687) );
  XNOR U12189 ( .A(n12682), .B(n12681), .Z(n12684) );
  XNOR U12190 ( .A(n12679), .B(n12678), .Z(n12681) );
  XNOR U12191 ( .A(n12676), .B(n12675), .Z(n12678) );
  XNOR U12192 ( .A(n12673), .B(n12672), .Z(n12675) );
  XNOR U12193 ( .A(n12670), .B(n12669), .Z(n12672) );
  XNOR U12194 ( .A(n12667), .B(n12666), .Z(n12669) );
  XNOR U12195 ( .A(n12664), .B(n12663), .Z(n12666) );
  XNOR U12196 ( .A(n12661), .B(n12660), .Z(n12663) );
  XNOR U12197 ( .A(n12658), .B(n12657), .Z(n12660) );
  XNOR U12198 ( .A(n12655), .B(n12654), .Z(n12657) );
  XNOR U12199 ( .A(n12652), .B(n12651), .Z(n12654) );
  XNOR U12200 ( .A(n12649), .B(n12648), .Z(n12651) );
  XNOR U12201 ( .A(n12646), .B(n12645), .Z(n12648) );
  XNOR U12202 ( .A(n12643), .B(n12642), .Z(n12645) );
  XNOR U12203 ( .A(n12640), .B(n12639), .Z(n12642) );
  XNOR U12204 ( .A(n12637), .B(n12636), .Z(n12639) );
  XNOR U12205 ( .A(n12634), .B(n12633), .Z(n12636) );
  XNOR U12206 ( .A(n12631), .B(n12630), .Z(n12633) );
  XNOR U12207 ( .A(n12628), .B(n12627), .Z(n12630) );
  XNOR U12208 ( .A(n12625), .B(n12624), .Z(n12627) );
  XNOR U12209 ( .A(n12622), .B(n12621), .Z(n12624) );
  XNOR U12210 ( .A(n12619), .B(n12618), .Z(n12621) );
  XNOR U12211 ( .A(n12616), .B(n12615), .Z(n12618) );
  XNOR U12212 ( .A(n12613), .B(n12612), .Z(n12615) );
  XNOR U12213 ( .A(n12610), .B(n12609), .Z(n12612) );
  XNOR U12214 ( .A(n12607), .B(n12606), .Z(n12609) );
  XNOR U12215 ( .A(n12604), .B(n12603), .Z(n12606) );
  XNOR U12216 ( .A(n12601), .B(n12600), .Z(n12603) );
  XNOR U12217 ( .A(n12598), .B(n12597), .Z(n12600) );
  XNOR U12218 ( .A(n12595), .B(n12594), .Z(n12597) );
  XNOR U12219 ( .A(n12592), .B(n12591), .Z(n12594) );
  XNOR U12220 ( .A(n12589), .B(n12588), .Z(n12591) );
  XNOR U12221 ( .A(n12586), .B(n12585), .Z(n12588) );
  XNOR U12222 ( .A(n12583), .B(n12582), .Z(n12585) );
  XNOR U12223 ( .A(n12580), .B(n12579), .Z(n12582) );
  XNOR U12224 ( .A(n12577), .B(n12576), .Z(n12579) );
  XNOR U12225 ( .A(n12574), .B(n12573), .Z(n12576) );
  XNOR U12226 ( .A(n12571), .B(n12570), .Z(n12573) );
  XNOR U12227 ( .A(n12568), .B(n12567), .Z(n12570) );
  XNOR U12228 ( .A(n12565), .B(n12564), .Z(n12567) );
  XNOR U12229 ( .A(n12562), .B(n12561), .Z(n12564) );
  XNOR U12230 ( .A(n12559), .B(n12558), .Z(n12561) );
  XNOR U12231 ( .A(n12556), .B(n12555), .Z(n12558) );
  XNOR U12232 ( .A(n12553), .B(n12552), .Z(n12555) );
  XNOR U12233 ( .A(n12550), .B(n12549), .Z(n12552) );
  XNOR U12234 ( .A(n12547), .B(n12546), .Z(n12549) );
  XNOR U12235 ( .A(n12544), .B(n12543), .Z(n12546) );
  XNOR U12236 ( .A(n12541), .B(n12540), .Z(n12543) );
  XNOR U12237 ( .A(n12538), .B(n12537), .Z(n12540) );
  XNOR U12238 ( .A(n12535), .B(n12534), .Z(n12537) );
  XNOR U12239 ( .A(n12532), .B(n12531), .Z(n12534) );
  XNOR U12240 ( .A(n12529), .B(n12528), .Z(n12531) );
  XNOR U12241 ( .A(n12526), .B(n12525), .Z(n12528) );
  XNOR U12242 ( .A(n12523), .B(n12522), .Z(n12525) );
  XNOR U12243 ( .A(n12520), .B(n12519), .Z(n12522) );
  XNOR U12244 ( .A(n12517), .B(n12516), .Z(n12519) );
  XNOR U12245 ( .A(n12514), .B(n12513), .Z(n12516) );
  XNOR U12246 ( .A(n12511), .B(n12510), .Z(n12513) );
  XNOR U12247 ( .A(n12508), .B(n12507), .Z(n12510) );
  XNOR U12248 ( .A(n12505), .B(n12504), .Z(n12507) );
  XNOR U12249 ( .A(n12502), .B(n12501), .Z(n12504) );
  XNOR U12250 ( .A(n12499), .B(n12498), .Z(n12501) );
  XNOR U12251 ( .A(n12496), .B(n12495), .Z(n12498) );
  XNOR U12252 ( .A(n12493), .B(n12492), .Z(n12495) );
  XNOR U12253 ( .A(n12490), .B(n12489), .Z(n12492) );
  XNOR U12254 ( .A(n12487), .B(n12486), .Z(n12489) );
  XNOR U12255 ( .A(n12484), .B(n12483), .Z(n12486) );
  XNOR U12256 ( .A(n12481), .B(n12480), .Z(n12483) );
  XNOR U12257 ( .A(n12478), .B(n12477), .Z(n12480) );
  XNOR U12258 ( .A(n12475), .B(n12474), .Z(n12477) );
  XNOR U12259 ( .A(n12472), .B(n12471), .Z(n12474) );
  XNOR U12260 ( .A(n12469), .B(n12468), .Z(n12471) );
  XNOR U12261 ( .A(n12466), .B(n12465), .Z(n12468) );
  XNOR U12262 ( .A(n12463), .B(n12462), .Z(n12465) );
  XNOR U12263 ( .A(n12460), .B(n12459), .Z(n12462) );
  XNOR U12264 ( .A(n12457), .B(n12456), .Z(n12459) );
  XNOR U12265 ( .A(n12454), .B(n12453), .Z(n12456) );
  XNOR U12266 ( .A(n12451), .B(n12450), .Z(n12453) );
  XNOR U12267 ( .A(n12448), .B(n12447), .Z(n12450) );
  XNOR U12268 ( .A(n12445), .B(n12444), .Z(n12447) );
  XNOR U12269 ( .A(n12442), .B(n12441), .Z(n12444) );
  XNOR U12270 ( .A(n12439), .B(n12438), .Z(n12441) );
  XNOR U12271 ( .A(n12436), .B(n12435), .Z(n12438) );
  XNOR U12272 ( .A(n12433), .B(n12432), .Z(n12435) );
  XNOR U12273 ( .A(n12430), .B(n12429), .Z(n12432) );
  XNOR U12274 ( .A(n12427), .B(n12426), .Z(n12429) );
  XNOR U12275 ( .A(n12424), .B(n12423), .Z(n12426) );
  XNOR U12276 ( .A(n12421), .B(n12420), .Z(n12423) );
  XNOR U12277 ( .A(n12418), .B(n12417), .Z(n12420) );
  XNOR U12278 ( .A(n12415), .B(n12414), .Z(n12417) );
  XNOR U12279 ( .A(n12412), .B(n12411), .Z(n12414) );
  XNOR U12280 ( .A(n12409), .B(n12408), .Z(n12411) );
  XNOR U12281 ( .A(n12406), .B(n12405), .Z(n12408) );
  XNOR U12282 ( .A(n12403), .B(n12402), .Z(n12405) );
  XNOR U12283 ( .A(n12400), .B(n12399), .Z(n12402) );
  XNOR U12284 ( .A(n12397), .B(n12396), .Z(n12399) );
  XNOR U12285 ( .A(n12394), .B(n12393), .Z(n12396) );
  XNOR U12286 ( .A(n12391), .B(n12390), .Z(n12393) );
  XNOR U12287 ( .A(n12388), .B(n12387), .Z(n12390) );
  XNOR U12288 ( .A(n12385), .B(n12384), .Z(n12387) );
  XNOR U12289 ( .A(n12382), .B(n12381), .Z(n12384) );
  XNOR U12290 ( .A(n12379), .B(n12378), .Z(n12381) );
  XNOR U12291 ( .A(n12376), .B(n12375), .Z(n12378) );
  XNOR U12292 ( .A(n12373), .B(n12372), .Z(n12375) );
  XNOR U12293 ( .A(n12370), .B(n12369), .Z(n12372) );
  XNOR U12294 ( .A(n12367), .B(n12366), .Z(n12369) );
  XNOR U12295 ( .A(n12364), .B(n12363), .Z(n12366) );
  XNOR U12296 ( .A(n12361), .B(n12360), .Z(n12363) );
  XNOR U12297 ( .A(n12358), .B(n12357), .Z(n12360) );
  XNOR U12298 ( .A(n12355), .B(n12354), .Z(n12357) );
  XNOR U12299 ( .A(n12352), .B(n12351), .Z(n12354) );
  XNOR U12300 ( .A(n12349), .B(n12348), .Z(n12351) );
  XNOR U12301 ( .A(n12346), .B(n12345), .Z(n12348) );
  XNOR U12302 ( .A(n12343), .B(n12342), .Z(n12345) );
  XNOR U12303 ( .A(n12340), .B(n12339), .Z(n12342) );
  XNOR U12304 ( .A(n12337), .B(n12336), .Z(n12339) );
  XNOR U12305 ( .A(n12334), .B(n12333), .Z(n12336) );
  XNOR U12306 ( .A(n12331), .B(n12330), .Z(n12333) );
  XNOR U12307 ( .A(n12328), .B(n12327), .Z(n12330) );
  XNOR U12308 ( .A(n12325), .B(n12324), .Z(n12327) );
  XNOR U12309 ( .A(n12322), .B(n12321), .Z(n12324) );
  XNOR U12310 ( .A(n12319), .B(n12318), .Z(n12321) );
  XNOR U12311 ( .A(n12316), .B(n12315), .Z(n12318) );
  XNOR U12312 ( .A(n12313), .B(n12312), .Z(n12315) );
  XNOR U12313 ( .A(n12310), .B(n12309), .Z(n12312) );
  XNOR U12314 ( .A(n12307), .B(n12306), .Z(n12309) );
  XNOR U12315 ( .A(n12304), .B(n12303), .Z(n12306) );
  XNOR U12316 ( .A(n12301), .B(n12300), .Z(n12303) );
  XNOR U12317 ( .A(n12298), .B(n12297), .Z(n12300) );
  XNOR U12318 ( .A(n12295), .B(n12294), .Z(n12297) );
  XNOR U12319 ( .A(n12292), .B(n12291), .Z(n12294) );
  XNOR U12320 ( .A(n12289), .B(n12288), .Z(n12291) );
  XNOR U12321 ( .A(n12286), .B(n12285), .Z(n12288) );
  XNOR U12322 ( .A(n12283), .B(n12282), .Z(n12285) );
  XNOR U12323 ( .A(n12280), .B(n12279), .Z(n12282) );
  XNOR U12324 ( .A(n12277), .B(n12276), .Z(n12279) );
  XNOR U12325 ( .A(n12274), .B(n12273), .Z(n12276) );
  XNOR U12326 ( .A(n12271), .B(n12270), .Z(n12273) );
  XNOR U12327 ( .A(n12268), .B(n12267), .Z(n12270) );
  XNOR U12328 ( .A(n12265), .B(n12264), .Z(n12267) );
  XNOR U12329 ( .A(n12262), .B(n12261), .Z(n12264) );
  XNOR U12330 ( .A(n12259), .B(n12258), .Z(n12261) );
  XNOR U12331 ( .A(n12256), .B(n12255), .Z(n12258) );
  XNOR U12332 ( .A(n12253), .B(n12252), .Z(n12255) );
  XNOR U12333 ( .A(n12250), .B(n12249), .Z(n12252) );
  XNOR U12334 ( .A(n12247), .B(n12246), .Z(n12249) );
  XNOR U12335 ( .A(n12244), .B(n12243), .Z(n12246) );
  XNOR U12336 ( .A(n12241), .B(n12240), .Z(n12243) );
  XNOR U12337 ( .A(n12238), .B(n12237), .Z(n12240) );
  XNOR U12338 ( .A(n12235), .B(n12234), .Z(n12237) );
  XNOR U12339 ( .A(n12232), .B(n12231), .Z(n12234) );
  XNOR U12340 ( .A(n12229), .B(n12228), .Z(n12231) );
  XNOR U12341 ( .A(n12226), .B(n12225), .Z(n12228) );
  XNOR U12342 ( .A(n12223), .B(n12222), .Z(n12225) );
  XNOR U12343 ( .A(n12220), .B(n12219), .Z(n12222) );
  XNOR U12344 ( .A(n12217), .B(n12216), .Z(n12219) );
  XNOR U12345 ( .A(n12214), .B(n12213), .Z(n12216) );
  XNOR U12346 ( .A(n12211), .B(n12210), .Z(n12213) );
  XNOR U12347 ( .A(n12208), .B(n12207), .Z(n12210) );
  XNOR U12348 ( .A(n12205), .B(n12204), .Z(n12207) );
  XNOR U12349 ( .A(n12202), .B(n12201), .Z(n12204) );
  XNOR U12350 ( .A(n12199), .B(n12198), .Z(n12201) );
  XNOR U12351 ( .A(n12196), .B(n12195), .Z(n12198) );
  XNOR U12352 ( .A(n12193), .B(n12192), .Z(n12195) );
  XNOR U12353 ( .A(n12190), .B(n12189), .Z(n12192) );
  XNOR U12354 ( .A(n12187), .B(n12186), .Z(n12189) );
  XNOR U12355 ( .A(n12184), .B(n12183), .Z(n12186) );
  XNOR U12356 ( .A(n12181), .B(n12180), .Z(n12183) );
  XNOR U12357 ( .A(n12178), .B(n12177), .Z(n12180) );
  XNOR U12358 ( .A(n12175), .B(n12174), .Z(n12177) );
  XNOR U12359 ( .A(n12172), .B(n12171), .Z(n12174) );
  XNOR U12360 ( .A(n12169), .B(n12168), .Z(n12171) );
  XNOR U12361 ( .A(n12166), .B(n12165), .Z(n12168) );
  XNOR U12362 ( .A(n12163), .B(n12162), .Z(n12165) );
  XNOR U12363 ( .A(n12160), .B(n12159), .Z(n12162) );
  XNOR U12364 ( .A(n12157), .B(n12156), .Z(n12159) );
  XNOR U12365 ( .A(n12154), .B(n12153), .Z(n12156) );
  XNOR U12366 ( .A(n12151), .B(n12150), .Z(n12153) );
  XNOR U12367 ( .A(n12148), .B(n12147), .Z(n12150) );
  XNOR U12368 ( .A(n12145), .B(n12144), .Z(n12147) );
  XNOR U12369 ( .A(n12142), .B(n12141), .Z(n12144) );
  XNOR U12370 ( .A(n12139), .B(n12138), .Z(n12141) );
  XNOR U12371 ( .A(n12136), .B(n12135), .Z(n12138) );
  XNOR U12372 ( .A(n12133), .B(n12132), .Z(n12135) );
  XNOR U12373 ( .A(n12130), .B(n12129), .Z(n12132) );
  XNOR U12374 ( .A(n12127), .B(n12126), .Z(n12129) );
  XNOR U12375 ( .A(n12124), .B(n12123), .Z(n12126) );
  XNOR U12376 ( .A(n12121), .B(n12120), .Z(n12123) );
  XNOR U12377 ( .A(n12118), .B(n12117), .Z(n12120) );
  XNOR U12378 ( .A(n12115), .B(n12114), .Z(n12117) );
  XNOR U12379 ( .A(n12112), .B(n12111), .Z(n12114) );
  XNOR U12380 ( .A(n12109), .B(n12108), .Z(n12111) );
  XNOR U12381 ( .A(n12106), .B(n12105), .Z(n12108) );
  XNOR U12382 ( .A(n12103), .B(n12102), .Z(n12105) );
  XNOR U12383 ( .A(n12100), .B(n12099), .Z(n12102) );
  XNOR U12384 ( .A(n12097), .B(n12096), .Z(n12099) );
  XNOR U12385 ( .A(n12094), .B(n12093), .Z(n12096) );
  XNOR U12386 ( .A(n12091), .B(n12090), .Z(n12093) );
  XNOR U12387 ( .A(n12088), .B(n12087), .Z(n12090) );
  XNOR U12388 ( .A(n12085), .B(n12084), .Z(n12087) );
  XNOR U12389 ( .A(n12082), .B(n12081), .Z(n12084) );
  XNOR U12390 ( .A(n12079), .B(n12078), .Z(n12081) );
  XNOR U12391 ( .A(n12076), .B(n12075), .Z(n12078) );
  XNOR U12392 ( .A(n12073), .B(n12072), .Z(n12075) );
  XNOR U12393 ( .A(n12070), .B(n12069), .Z(n12072) );
  XNOR U12394 ( .A(n12067), .B(n12066), .Z(n12069) );
  XNOR U12395 ( .A(n12064), .B(n12063), .Z(n12066) );
  XNOR U12396 ( .A(n12061), .B(n12060), .Z(n12063) );
  XNOR U12397 ( .A(n12058), .B(n12057), .Z(n12060) );
  XNOR U12398 ( .A(n12055), .B(n12054), .Z(n12057) );
  XNOR U12399 ( .A(n12052), .B(n12051), .Z(n12054) );
  XNOR U12400 ( .A(n12049), .B(n12048), .Z(n12051) );
  XNOR U12401 ( .A(n12046), .B(n12045), .Z(n12048) );
  XNOR U12402 ( .A(n12043), .B(n12042), .Z(n12045) );
  XNOR U12403 ( .A(n12040), .B(n12039), .Z(n12042) );
  XNOR U12404 ( .A(n12037), .B(n12036), .Z(n12039) );
  XNOR U12405 ( .A(n12034), .B(n12033), .Z(n12036) );
  XNOR U12406 ( .A(n12031), .B(n12030), .Z(n12033) );
  XNOR U12407 ( .A(n12028), .B(n12027), .Z(n12030) );
  XNOR U12408 ( .A(n12025), .B(n12024), .Z(n12027) );
  XNOR U12409 ( .A(n12022), .B(n12021), .Z(n12024) );
  XNOR U12410 ( .A(n12019), .B(n12018), .Z(n12021) );
  XNOR U12411 ( .A(n12016), .B(n12015), .Z(n12018) );
  XNOR U12412 ( .A(n12013), .B(n12012), .Z(n12015) );
  XNOR U12413 ( .A(n12010), .B(n12009), .Z(n12012) );
  XNOR U12414 ( .A(n12007), .B(n12006), .Z(n12009) );
  XNOR U12415 ( .A(n12004), .B(n12003), .Z(n12006) );
  XNOR U12416 ( .A(n12001), .B(n12000), .Z(n12003) );
  XNOR U12417 ( .A(n11998), .B(n11997), .Z(n12000) );
  XNOR U12418 ( .A(n11995), .B(n11994), .Z(n11997) );
  XNOR U12419 ( .A(n11992), .B(n11991), .Z(n11994) );
  XNOR U12420 ( .A(n11989), .B(n11988), .Z(n11991) );
  XNOR U12421 ( .A(n11986), .B(n11985), .Z(n11988) );
  XNOR U12422 ( .A(n11983), .B(n11982), .Z(n11985) );
  XNOR U12423 ( .A(n11980), .B(n11979), .Z(n11982) );
  XNOR U12424 ( .A(n11977), .B(n11976), .Z(n11979) );
  XNOR U12425 ( .A(n11974), .B(n11973), .Z(n11976) );
  XNOR U12426 ( .A(n11971), .B(n11970), .Z(n11973) );
  XNOR U12427 ( .A(n11968), .B(n11967), .Z(n11970) );
  XNOR U12428 ( .A(n11965), .B(n11964), .Z(n11967) );
  XNOR U12429 ( .A(n11962), .B(n11961), .Z(n11964) );
  XNOR U12430 ( .A(n11959), .B(n11958), .Z(n11961) );
  XNOR U12431 ( .A(n11956), .B(n11955), .Z(n11958) );
  XNOR U12432 ( .A(n11953), .B(n11952), .Z(n11955) );
  XNOR U12433 ( .A(n11950), .B(n11949), .Z(n11952) );
  XNOR U12434 ( .A(n11947), .B(n11946), .Z(n11949) );
  XNOR U12435 ( .A(n11944), .B(n11943), .Z(n11946) );
  XNOR U12436 ( .A(n11941), .B(n11940), .Z(n11943) );
  XNOR U12437 ( .A(n11938), .B(n11937), .Z(n11940) );
  XNOR U12438 ( .A(n11935), .B(n11934), .Z(n11937) );
  XNOR U12439 ( .A(n11932), .B(n11931), .Z(n11934) );
  XNOR U12440 ( .A(n11929), .B(n11928), .Z(n11931) );
  XNOR U12441 ( .A(n11926), .B(n11925), .Z(n11928) );
  XNOR U12442 ( .A(n11923), .B(n11922), .Z(n11925) );
  XNOR U12443 ( .A(n11920), .B(n11919), .Z(n11922) );
  XNOR U12444 ( .A(n11917), .B(n11916), .Z(n11919) );
  XNOR U12445 ( .A(n11914), .B(n11913), .Z(n11916) );
  XNOR U12446 ( .A(n11911), .B(n11910), .Z(n11913) );
  XNOR U12447 ( .A(n11908), .B(n11907), .Z(n11910) );
  XNOR U12448 ( .A(n11905), .B(n11904), .Z(n11907) );
  XNOR U12449 ( .A(n11902), .B(n11901), .Z(n11904) );
  XNOR U12450 ( .A(n11899), .B(n11898), .Z(n11901) );
  XNOR U12451 ( .A(n11896), .B(n11895), .Z(n11898) );
  XNOR U12452 ( .A(n11893), .B(n11892), .Z(n11895) );
  XNOR U12453 ( .A(n11890), .B(n11889), .Z(n11892) );
  XNOR U12454 ( .A(n11887), .B(n11886), .Z(n11889) );
  XNOR U12455 ( .A(n11884), .B(n11883), .Z(n11886) );
  XNOR U12456 ( .A(n11881), .B(n11880), .Z(n11883) );
  XNOR U12457 ( .A(n11878), .B(n11877), .Z(n11880) );
  XNOR U12458 ( .A(n11875), .B(n11874), .Z(n11877) );
  XNOR U12459 ( .A(n11872), .B(n11871), .Z(n11874) );
  XNOR U12460 ( .A(n11869), .B(n11868), .Z(n11871) );
  XNOR U12461 ( .A(n11866), .B(n11865), .Z(n11868) );
  XNOR U12462 ( .A(n11863), .B(n11862), .Z(n11865) );
  XNOR U12463 ( .A(n11860), .B(n11859), .Z(n11862) );
  XNOR U12464 ( .A(n11857), .B(n11856), .Z(n11859) );
  XNOR U12465 ( .A(n11854), .B(n11853), .Z(n11856) );
  XNOR U12466 ( .A(n11851), .B(n11850), .Z(n11853) );
  XNOR U12467 ( .A(n11848), .B(n11847), .Z(n11850) );
  XNOR U12468 ( .A(n11845), .B(n11844), .Z(n11847) );
  XNOR U12469 ( .A(n11842), .B(n11841), .Z(n11844) );
  XNOR U12470 ( .A(n11839), .B(n11838), .Z(n11841) );
  XNOR U12471 ( .A(n11836), .B(n11835), .Z(n11838) );
  XNOR U12472 ( .A(n11833), .B(n11832), .Z(n11835) );
  XNOR U12473 ( .A(n11830), .B(n11829), .Z(n11832) );
  XNOR U12474 ( .A(n11827), .B(n11826), .Z(n11829) );
  XNOR U12475 ( .A(n11824), .B(n11823), .Z(n11826) );
  XNOR U12476 ( .A(n11821), .B(n11820), .Z(n11823) );
  XNOR U12477 ( .A(n11818), .B(n11817), .Z(n11820) );
  XNOR U12478 ( .A(n11815), .B(n11814), .Z(n11817) );
  XNOR U12479 ( .A(n11812), .B(n11811), .Z(n11814) );
  XNOR U12480 ( .A(n11809), .B(n11808), .Z(n11811) );
  XNOR U12481 ( .A(n11806), .B(n11805), .Z(n11808) );
  XNOR U12482 ( .A(n11803), .B(n11802), .Z(n11805) );
  XNOR U12483 ( .A(n11800), .B(n11799), .Z(n11802) );
  XNOR U12484 ( .A(n11797), .B(n11796), .Z(n11799) );
  XNOR U12485 ( .A(n11794), .B(n11793), .Z(n11796) );
  XNOR U12486 ( .A(n11791), .B(n11790), .Z(n11793) );
  XNOR U12487 ( .A(n11788), .B(n11787), .Z(n11790) );
  XNOR U12488 ( .A(n11785), .B(n11784), .Z(n11787) );
  XNOR U12489 ( .A(n11782), .B(n11781), .Z(n11784) );
  XNOR U12490 ( .A(n11779), .B(n11778), .Z(n11781) );
  XNOR U12491 ( .A(n11776), .B(n11775), .Z(n11778) );
  XNOR U12492 ( .A(n11773), .B(n11772), .Z(n11775) );
  XNOR U12493 ( .A(n11770), .B(n11769), .Z(n11772) );
  XNOR U12494 ( .A(n11767), .B(n11766), .Z(n11769) );
  XNOR U12495 ( .A(n11764), .B(n11763), .Z(n11766) );
  XNOR U12496 ( .A(n11761), .B(n11760), .Z(n11763) );
  XNOR U12497 ( .A(n11758), .B(n11757), .Z(n11760) );
  XNOR U12498 ( .A(n11755), .B(n11754), .Z(n11757) );
  XNOR U12499 ( .A(n11752), .B(n11751), .Z(n11754) );
  XNOR U12500 ( .A(n11749), .B(n11748), .Z(n11751) );
  XNOR U12501 ( .A(n11746), .B(n11745), .Z(n11748) );
  XNOR U12502 ( .A(n11743), .B(n11742), .Z(n11745) );
  XNOR U12503 ( .A(n11740), .B(n11739), .Z(n11742) );
  XNOR U12504 ( .A(n11737), .B(n11736), .Z(n11739) );
  XNOR U12505 ( .A(n11734), .B(n11733), .Z(n11736) );
  XNOR U12506 ( .A(n11731), .B(n11730), .Z(n11733) );
  XNOR U12507 ( .A(n11728), .B(n11727), .Z(n11730) );
  XNOR U12508 ( .A(n11725), .B(n11724), .Z(n11727) );
  XNOR U12509 ( .A(n11722), .B(n11721), .Z(n11724) );
  XNOR U12510 ( .A(n11719), .B(n11718), .Z(n11721) );
  XNOR U12511 ( .A(n11716), .B(n11715), .Z(n11718) );
  XNOR U12512 ( .A(n11713), .B(n11712), .Z(n11715) );
  XNOR U12513 ( .A(n11710), .B(n11709), .Z(n11712) );
  XNOR U12514 ( .A(n11707), .B(n11706), .Z(n11709) );
  XNOR U12515 ( .A(n11704), .B(n11703), .Z(n11706) );
  XNOR U12516 ( .A(n11701), .B(n11700), .Z(n11703) );
  XNOR U12517 ( .A(n11698), .B(n11697), .Z(n11700) );
  XNOR U12518 ( .A(n11695), .B(n11694), .Z(n11697) );
  XNOR U12519 ( .A(n11692), .B(n11691), .Z(n11694) );
  XNOR U12520 ( .A(n11689), .B(n11688), .Z(n11691) );
  XNOR U12521 ( .A(n11686), .B(n11685), .Z(n11688) );
  XNOR U12522 ( .A(n11683), .B(n11682), .Z(n11685) );
  XNOR U12523 ( .A(n11680), .B(n11679), .Z(n11682) );
  XNOR U12524 ( .A(n11677), .B(n11676), .Z(n11679) );
  XNOR U12525 ( .A(n11674), .B(n11673), .Z(n11676) );
  XNOR U12526 ( .A(n11671), .B(n11670), .Z(n11673) );
  XNOR U12527 ( .A(n11668), .B(n11667), .Z(n11670) );
  XNOR U12528 ( .A(n11665), .B(n11664), .Z(n11667) );
  XNOR U12529 ( .A(n11662), .B(n11661), .Z(n11664) );
  XNOR U12530 ( .A(n11659), .B(n11658), .Z(n11661) );
  XNOR U12531 ( .A(n11656), .B(n11655), .Z(n11658) );
  XNOR U12532 ( .A(n11653), .B(n11652), .Z(n11655) );
  XNOR U12533 ( .A(n11650), .B(n11649), .Z(n11652) );
  XNOR U12534 ( .A(n11647), .B(n11646), .Z(n11649) );
  XNOR U12535 ( .A(n11644), .B(n11643), .Z(n11646) );
  XNOR U12536 ( .A(n11641), .B(n11640), .Z(n11643) );
  XNOR U12537 ( .A(n11638), .B(n11637), .Z(n11640) );
  XNOR U12538 ( .A(n11635), .B(n11634), .Z(n11637) );
  XNOR U12539 ( .A(n11632), .B(n11631), .Z(n11634) );
  XNOR U12540 ( .A(n11629), .B(n11628), .Z(n11631) );
  XNOR U12541 ( .A(n11626), .B(n11625), .Z(n11628) );
  XNOR U12542 ( .A(n11623), .B(n11622), .Z(n11625) );
  XNOR U12543 ( .A(n11620), .B(n11619), .Z(n11622) );
  XNOR U12544 ( .A(n11617), .B(n11616), .Z(n11619) );
  XNOR U12545 ( .A(n11614), .B(n11613), .Z(n11616) );
  XNOR U12546 ( .A(n11611), .B(n11610), .Z(n11613) );
  XNOR U12547 ( .A(n11608), .B(n11607), .Z(n11610) );
  XNOR U12548 ( .A(n11605), .B(n11604), .Z(n11607) );
  XNOR U12549 ( .A(n11602), .B(n11601), .Z(n11604) );
  XNOR U12550 ( .A(n11599), .B(n11598), .Z(n11601) );
  XNOR U12551 ( .A(n11596), .B(n11595), .Z(n11598) );
  XNOR U12552 ( .A(n11593), .B(n11592), .Z(n11595) );
  XNOR U12553 ( .A(n11590), .B(n11589), .Z(n11592) );
  XNOR U12554 ( .A(n11587), .B(n11586), .Z(n11589) );
  XNOR U12555 ( .A(n11584), .B(n11583), .Z(n11586) );
  XNOR U12556 ( .A(n11581), .B(n11580), .Z(n11583) );
  XNOR U12557 ( .A(n11578), .B(n11577), .Z(n11580) );
  XNOR U12558 ( .A(n11575), .B(n11574), .Z(n11577) );
  XNOR U12559 ( .A(n11572), .B(n11571), .Z(n11574) );
  XOR U12560 ( .A(n11569), .B(n11568), .Z(n11571) );
  XOR U12561 ( .A(n11566), .B(n11565), .Z(n11568) );
  XOR U12562 ( .A(n11562), .B(n11563), .Z(n11565) );
  AND U12563 ( .A(n14172), .B(n14173), .Z(n11563) );
  XOR U12564 ( .A(n11559), .B(n11560), .Z(n11562) );
  AND U12565 ( .A(n14174), .B(n14175), .Z(n11560) );
  XOR U12566 ( .A(n11556), .B(n11557), .Z(n11559) );
  AND U12567 ( .A(n14176), .B(n14177), .Z(n11557) );
  XNOR U12568 ( .A(n11311), .B(n11554), .Z(n11556) );
  AND U12569 ( .A(n14178), .B(n14179), .Z(n11554) );
  XOR U12570 ( .A(n11313), .B(n11312), .Z(n11311) );
  AND U12571 ( .A(n14180), .B(n14181), .Z(n11312) );
  XOR U12572 ( .A(n11315), .B(n11314), .Z(n11313) );
  AND U12573 ( .A(n14182), .B(n14183), .Z(n11314) );
  XOR U12574 ( .A(n11317), .B(n11316), .Z(n11315) );
  AND U12575 ( .A(n14184), .B(n14185), .Z(n11316) );
  XOR U12576 ( .A(n11319), .B(n11318), .Z(n11317) );
  AND U12577 ( .A(n14186), .B(n14187), .Z(n11318) );
  XOR U12578 ( .A(n11321), .B(n11320), .Z(n11319) );
  AND U12579 ( .A(n14188), .B(n14189), .Z(n11320) );
  XOR U12580 ( .A(n11323), .B(n11322), .Z(n11321) );
  AND U12581 ( .A(n14190), .B(n14191), .Z(n11322) );
  XOR U12582 ( .A(n11325), .B(n11324), .Z(n11323) );
  AND U12583 ( .A(n14192), .B(n14193), .Z(n11324) );
  XOR U12584 ( .A(n11327), .B(n11326), .Z(n11325) );
  AND U12585 ( .A(n14194), .B(n14195), .Z(n11326) );
  XOR U12586 ( .A(n11329), .B(n11328), .Z(n11327) );
  AND U12587 ( .A(n14196), .B(n14197), .Z(n11328) );
  XOR U12588 ( .A(n11331), .B(n11330), .Z(n11329) );
  AND U12589 ( .A(n14198), .B(n14199), .Z(n11330) );
  XOR U12590 ( .A(n11333), .B(n11332), .Z(n11331) );
  AND U12591 ( .A(n14200), .B(n14201), .Z(n11332) );
  XOR U12592 ( .A(n11335), .B(n11334), .Z(n11333) );
  AND U12593 ( .A(n14202), .B(n14203), .Z(n11334) );
  XOR U12594 ( .A(n11337), .B(n11336), .Z(n11335) );
  AND U12595 ( .A(n14204), .B(n14205), .Z(n11336) );
  XOR U12596 ( .A(n11339), .B(n11338), .Z(n11337) );
  AND U12597 ( .A(n14206), .B(n14207), .Z(n11338) );
  XOR U12598 ( .A(n11341), .B(n11340), .Z(n11339) );
  AND U12599 ( .A(n14208), .B(n14209), .Z(n11340) );
  XOR U12600 ( .A(n11343), .B(n11342), .Z(n11341) );
  AND U12601 ( .A(n14210), .B(n14211), .Z(n11342) );
  XOR U12602 ( .A(n11345), .B(n11344), .Z(n11343) );
  AND U12603 ( .A(n14212), .B(n14213), .Z(n11344) );
  XOR U12604 ( .A(n11347), .B(n11346), .Z(n11345) );
  AND U12605 ( .A(n14214), .B(n14215), .Z(n11346) );
  XOR U12606 ( .A(n11349), .B(n11348), .Z(n11347) );
  AND U12607 ( .A(n14216), .B(n14217), .Z(n11348) );
  XOR U12608 ( .A(n11351), .B(n11350), .Z(n11349) );
  AND U12609 ( .A(n14218), .B(n14219), .Z(n11350) );
  XOR U12610 ( .A(n11353), .B(n11352), .Z(n11351) );
  AND U12611 ( .A(n14220), .B(n14221), .Z(n11352) );
  XOR U12612 ( .A(n11355), .B(n11354), .Z(n11353) );
  AND U12613 ( .A(n14222), .B(n14223), .Z(n11354) );
  XOR U12614 ( .A(n11357), .B(n11356), .Z(n11355) );
  AND U12615 ( .A(n14224), .B(n14225), .Z(n11356) );
  XOR U12616 ( .A(n11359), .B(n11358), .Z(n11357) );
  AND U12617 ( .A(n14226), .B(n14227), .Z(n11358) );
  XOR U12618 ( .A(n11361), .B(n11360), .Z(n11359) );
  AND U12619 ( .A(n14228), .B(n14229), .Z(n11360) );
  XOR U12620 ( .A(n11363), .B(n11362), .Z(n11361) );
  AND U12621 ( .A(n14230), .B(n14231), .Z(n11362) );
  XOR U12622 ( .A(n11365), .B(n11364), .Z(n11363) );
  AND U12623 ( .A(n14232), .B(n14233), .Z(n11364) );
  XOR U12624 ( .A(n11367), .B(n11366), .Z(n11365) );
  AND U12625 ( .A(n14234), .B(n14235), .Z(n11366) );
  XOR U12626 ( .A(n11369), .B(n11368), .Z(n11367) );
  AND U12627 ( .A(n14236), .B(n14237), .Z(n11368) );
  XOR U12628 ( .A(n11371), .B(n11370), .Z(n11369) );
  AND U12629 ( .A(n14238), .B(n14239), .Z(n11370) );
  XOR U12630 ( .A(n11373), .B(n11372), .Z(n11371) );
  AND U12631 ( .A(n14240), .B(n14241), .Z(n11372) );
  XOR U12632 ( .A(n11375), .B(n11374), .Z(n11373) );
  AND U12633 ( .A(n14242), .B(n14243), .Z(n11374) );
  XOR U12634 ( .A(n11377), .B(n11376), .Z(n11375) );
  AND U12635 ( .A(n14244), .B(n14245), .Z(n11376) );
  XOR U12636 ( .A(n11379), .B(n11378), .Z(n11377) );
  AND U12637 ( .A(n14246), .B(n14247), .Z(n11378) );
  XOR U12638 ( .A(n11381), .B(n11380), .Z(n11379) );
  AND U12639 ( .A(n14248), .B(n14249), .Z(n11380) );
  XOR U12640 ( .A(n11383), .B(n11382), .Z(n11381) );
  AND U12641 ( .A(n14250), .B(n14251), .Z(n11382) );
  XOR U12642 ( .A(n11385), .B(n11384), .Z(n11383) );
  AND U12643 ( .A(n14252), .B(n14253), .Z(n11384) );
  XOR U12644 ( .A(n11387), .B(n11386), .Z(n11385) );
  AND U12645 ( .A(n14254), .B(n14255), .Z(n11386) );
  XOR U12646 ( .A(n11389), .B(n11388), .Z(n11387) );
  AND U12647 ( .A(n14256), .B(n14257), .Z(n11388) );
  XOR U12648 ( .A(n11391), .B(n11390), .Z(n11389) );
  AND U12649 ( .A(n14258), .B(n14259), .Z(n11390) );
  XOR U12650 ( .A(n11393), .B(n11392), .Z(n11391) );
  AND U12651 ( .A(n14260), .B(n14261), .Z(n11392) );
  XOR U12652 ( .A(n11395), .B(n11394), .Z(n11393) );
  AND U12653 ( .A(n14262), .B(n14263), .Z(n11394) );
  XOR U12654 ( .A(n11397), .B(n11396), .Z(n11395) );
  AND U12655 ( .A(n14264), .B(n14265), .Z(n11396) );
  XOR U12656 ( .A(n11399), .B(n11398), .Z(n11397) );
  AND U12657 ( .A(n14266), .B(n14267), .Z(n11398) );
  XOR U12658 ( .A(n11401), .B(n11400), .Z(n11399) );
  AND U12659 ( .A(n14268), .B(n14269), .Z(n11400) );
  XOR U12660 ( .A(n11403), .B(n11402), .Z(n11401) );
  AND U12661 ( .A(n14270), .B(n14271), .Z(n11402) );
  XOR U12662 ( .A(n11405), .B(n11404), .Z(n11403) );
  AND U12663 ( .A(n14272), .B(n14273), .Z(n11404) );
  XOR U12664 ( .A(n11407), .B(n11406), .Z(n11405) );
  AND U12665 ( .A(n14274), .B(n14275), .Z(n11406) );
  XOR U12666 ( .A(n11409), .B(n11408), .Z(n11407) );
  AND U12667 ( .A(n14276), .B(n14277), .Z(n11408) );
  XOR U12668 ( .A(n11411), .B(n11410), .Z(n11409) );
  AND U12669 ( .A(n14278), .B(n14279), .Z(n11410) );
  XOR U12670 ( .A(n11413), .B(n11412), .Z(n11411) );
  AND U12671 ( .A(n14280), .B(n14281), .Z(n11412) );
  XOR U12672 ( .A(n11415), .B(n11414), .Z(n11413) );
  AND U12673 ( .A(n14282), .B(n14283), .Z(n11414) );
  XOR U12674 ( .A(n11417), .B(n11416), .Z(n11415) );
  AND U12675 ( .A(n14284), .B(n14285), .Z(n11416) );
  XOR U12676 ( .A(n11419), .B(n11418), .Z(n11417) );
  AND U12677 ( .A(n14286), .B(n14287), .Z(n11418) );
  XOR U12678 ( .A(n11421), .B(n11420), .Z(n11419) );
  AND U12679 ( .A(n14288), .B(n14289), .Z(n11420) );
  XOR U12680 ( .A(n11423), .B(n11422), .Z(n11421) );
  AND U12681 ( .A(n14290), .B(n14291), .Z(n11422) );
  XOR U12682 ( .A(n11425), .B(n11424), .Z(n11423) );
  AND U12683 ( .A(n14292), .B(n14293), .Z(n11424) );
  XOR U12684 ( .A(n11427), .B(n11426), .Z(n11425) );
  AND U12685 ( .A(n14294), .B(n14295), .Z(n11426) );
  XOR U12686 ( .A(n11429), .B(n11428), .Z(n11427) );
  AND U12687 ( .A(n14296), .B(n14297), .Z(n11428) );
  XOR U12688 ( .A(n11431), .B(n11430), .Z(n11429) );
  AND U12689 ( .A(n14298), .B(n14299), .Z(n11430) );
  XOR U12690 ( .A(n11433), .B(n11432), .Z(n11431) );
  AND U12691 ( .A(n14300), .B(n14301), .Z(n11432) );
  XOR U12692 ( .A(n11435), .B(n11434), .Z(n11433) );
  AND U12693 ( .A(n14302), .B(n14303), .Z(n11434) );
  XOR U12694 ( .A(n11437), .B(n11436), .Z(n11435) );
  AND U12695 ( .A(n14304), .B(n14305), .Z(n11436) );
  XOR U12696 ( .A(n11439), .B(n11438), .Z(n11437) );
  AND U12697 ( .A(n14306), .B(n14307), .Z(n11438) );
  XOR U12698 ( .A(n11441), .B(n11440), .Z(n11439) );
  AND U12699 ( .A(n14308), .B(n14309), .Z(n11440) );
  XOR U12700 ( .A(n11443), .B(n11442), .Z(n11441) );
  AND U12701 ( .A(n14310), .B(n14311), .Z(n11442) );
  XOR U12702 ( .A(n11445), .B(n11444), .Z(n11443) );
  AND U12703 ( .A(n14312), .B(n14313), .Z(n11444) );
  XOR U12704 ( .A(n11447), .B(n11446), .Z(n11445) );
  AND U12705 ( .A(n14314), .B(n14315), .Z(n11446) );
  XOR U12706 ( .A(n11456), .B(n11448), .Z(n11447) );
  AND U12707 ( .A(n14316), .B(n14317), .Z(n11448) );
  XOR U12708 ( .A(n11451), .B(n11457), .Z(n11456) );
  AND U12709 ( .A(n14318), .B(n14319), .Z(n11457) );
  XOR U12710 ( .A(n11453), .B(n11452), .Z(n11451) );
  AND U12711 ( .A(n14320), .B(n14321), .Z(n11452) );
  XOR U12712 ( .A(n11477), .B(n11454), .Z(n11453) );
  AND U12713 ( .A(n14322), .B(n14323), .Z(n11454) );
  XOR U12714 ( .A(n11472), .B(n11478), .Z(n11477) );
  AND U12715 ( .A(n14324), .B(n14325), .Z(n11478) );
  XOR U12716 ( .A(n11474), .B(n11473), .Z(n11472) );
  AND U12717 ( .A(n14326), .B(n14327), .Z(n11473) );
  XOR U12718 ( .A(n11462), .B(n11475), .Z(n11474) );
  AND U12719 ( .A(n14328), .B(n14329), .Z(n11475) );
  XOR U12720 ( .A(n11464), .B(n11463), .Z(n11462) );
  AND U12721 ( .A(n14330), .B(n14331), .Z(n11463) );
  XOR U12722 ( .A(n11466), .B(n11465), .Z(n11464) );
  AND U12723 ( .A(n14332), .B(n14333), .Z(n11465) );
  XOR U12724 ( .A(n11468), .B(n11467), .Z(n11466) );
  AND U12725 ( .A(n14334), .B(n14335), .Z(n11467) );
  XOR U12726 ( .A(n11498), .B(n11469), .Z(n11468) );
  AND U12727 ( .A(n14336), .B(n14337), .Z(n11469) );
  XOR U12728 ( .A(n11494), .B(n11499), .Z(n11498) );
  AND U12729 ( .A(n14338), .B(n14339), .Z(n11499) );
  XOR U12730 ( .A(n11496), .B(n11495), .Z(n11494) );
  AND U12731 ( .A(n14340), .B(n14341), .Z(n11495) );
  XOR U12732 ( .A(n11483), .B(n11497), .Z(n11496) );
  AND U12733 ( .A(n14342), .B(n14343), .Z(n11497) );
  XOR U12734 ( .A(n11485), .B(n11484), .Z(n11483) );
  AND U12735 ( .A(n14344), .B(n14345), .Z(n11484) );
  XOR U12736 ( .A(n11488), .B(n11486), .Z(n11485) );
  AND U12737 ( .A(n14346), .B(n14347), .Z(n11486) );
  XOR U12738 ( .A(n11490), .B(n11489), .Z(n11488) );
  AND U12739 ( .A(n14348), .B(n14349), .Z(n11489) );
  XOR U12740 ( .A(n11508), .B(n11491), .Z(n11490) );
  AND U12741 ( .A(n14350), .B(n14351), .Z(n11491) );
  XNOR U12742 ( .A(n11515), .B(n11509), .Z(n11508) );
  AND U12743 ( .A(n14352), .B(n14353), .Z(n11509) );
  XOR U12744 ( .A(n11514), .B(n11506), .Z(n11515) );
  AND U12745 ( .A(n14354), .B(n14355), .Z(n11506) );
  XOR U12746 ( .A(n11553), .B(n11505), .Z(n11514) );
  AND U12747 ( .A(n14356), .B(n14357), .Z(n11505) );
  XNOR U12748 ( .A(n11526), .B(n11504), .Z(n11553) );
  AND U12749 ( .A(n14358), .B(n14359), .Z(n11504) );
  XNOR U12750 ( .A(n11533), .B(n11527), .Z(n11526) );
  AND U12751 ( .A(n14360), .B(n14361), .Z(n11527) );
  XOR U12752 ( .A(n11532), .B(n11524), .Z(n11533) );
  AND U12753 ( .A(n14362), .B(n14363), .Z(n11524) );
  XOR U12754 ( .A(n11552), .B(n11523), .Z(n11532) );
  AND U12755 ( .A(n14364), .B(n14365), .Z(n11523) );
  XNOR U12756 ( .A(n14366), .B(n14367), .Z(n11552) );
  XOR U12757 ( .A(n14368), .B(n14369), .Z(n14367) );
  XOR U12758 ( .A(n14370), .B(n14371), .Z(n14369) );
  XNOR U12759 ( .A(n11550), .B(n11543), .Z(n14371) );
  XNOR U12760 ( .A(n14372), .B(n14373), .Z(n11543) );
  AND U12761 ( .A(n14374), .B(n14375), .Z(n14373) );
  NOR U12762 ( .A(n14376), .B(n14377), .Z(n14375) );
  NOR U12763 ( .A(n14378), .B(n14379), .Z(n14374) );
  AND U12764 ( .A(n14380), .B(n14381), .Z(n14379) );
  AND U12765 ( .A(n14382), .B(n14383), .Z(n14372) );
  NOR U12766 ( .A(n14384), .B(n14385), .Z(n14383) );
  AND U12767 ( .A(n14377), .B(n14386), .Z(n14385) );
  AND U12768 ( .A(n14378), .B(n14387), .Z(n14384) );
  NOR U12769 ( .A(n14388), .B(n14389), .Z(n14382) );
  AND U12770 ( .A(n14390), .B(n14391), .Z(n14389) );
  NOR U12771 ( .A(n14392), .B(n14393), .Z(n14391) );
  IV U12772 ( .A(n14394), .Z(n14392) );
  NOR U12773 ( .A(n14395), .B(n14396), .Z(n14394) );
  NOR U12774 ( .A(n14397), .B(n14398), .Z(n14390) );
  AND U12775 ( .A(n14376), .B(n14399), .Z(n14388) );
  AND U12776 ( .A(n14400), .B(n14401), .Z(n11550) );
  XOR U12777 ( .A(n11548), .B(n11549), .Z(n14370) );
  AND U12778 ( .A(n14402), .B(n14403), .Z(n11549) );
  AND U12779 ( .A(n14404), .B(n14405), .Z(n11548) );
  XOR U12780 ( .A(n14406), .B(n14407), .Z(n14368) );
  XOR U12781 ( .A(n11544), .B(n11545), .Z(n14407) );
  AND U12782 ( .A(n14408), .B(n14409), .Z(n11545) );
  AND U12783 ( .A(n14410), .B(n14411), .Z(n11544) );
  XNOR U12784 ( .A(n11542), .B(n11541), .Z(n14406) );
  IV U12785 ( .A(n14412), .Z(n11541) );
  AND U12786 ( .A(n14413), .B(n14414), .Z(n14412) );
  AND U12787 ( .A(n14415), .B(n14416), .Z(n11542) );
  XNOR U12788 ( .A(n11551), .B(n11522), .Z(n14366) );
  AND U12789 ( .A(n14417), .B(n14418), .Z(n11522) );
  AND U12790 ( .A(n14419), .B(n14420), .Z(n11551) );
  XOR U12791 ( .A(n14421), .B(n14422), .Z(n11566) );
  AND U12792 ( .A(n14421), .B(n14423), .Z(n14422) );
  XNOR U12793 ( .A(n14424), .B(n14425), .Z(n11569) );
  AND U12794 ( .A(n14424), .B(n14426), .Z(n14425) );
  XNOR U12795 ( .A(n14427), .B(n14428), .Z(n11572) );
  AND U12796 ( .A(n14427), .B(n14429), .Z(n14428) );
  XNOR U12797 ( .A(n14430), .B(n14431), .Z(n11575) );
  AND U12798 ( .A(n14430), .B(n14432), .Z(n14431) );
  XNOR U12799 ( .A(n14433), .B(n14434), .Z(n11578) );
  AND U12800 ( .A(n14435), .B(n14433), .Z(n14434) );
  XOR U12801 ( .A(n14436), .B(n14437), .Z(n11581) );
  NOR U12802 ( .A(n14438), .B(n14436), .Z(n14437) );
  XOR U12803 ( .A(n14439), .B(n14440), .Z(n11584) );
  NOR U12804 ( .A(n14441), .B(n14439), .Z(n14440) );
  XOR U12805 ( .A(n14442), .B(n14443), .Z(n11587) );
  NOR U12806 ( .A(n14444), .B(n14442), .Z(n14443) );
  XOR U12807 ( .A(n14445), .B(n14446), .Z(n11590) );
  NOR U12808 ( .A(n14447), .B(n14445), .Z(n14446) );
  XOR U12809 ( .A(n14448), .B(n14449), .Z(n11593) );
  NOR U12810 ( .A(n14450), .B(n14448), .Z(n14449) );
  XOR U12811 ( .A(n14451), .B(n14452), .Z(n11596) );
  NOR U12812 ( .A(n14453), .B(n14451), .Z(n14452) );
  XOR U12813 ( .A(n14454), .B(n14455), .Z(n11599) );
  NOR U12814 ( .A(n14456), .B(n14454), .Z(n14455) );
  XOR U12815 ( .A(n14457), .B(n14458), .Z(n11602) );
  NOR U12816 ( .A(n14459), .B(n14457), .Z(n14458) );
  XOR U12817 ( .A(n14460), .B(n14461), .Z(n11605) );
  NOR U12818 ( .A(n14462), .B(n14460), .Z(n14461) );
  XOR U12819 ( .A(n14463), .B(n14464), .Z(n11608) );
  NOR U12820 ( .A(n14465), .B(n14463), .Z(n14464) );
  XOR U12821 ( .A(n14466), .B(n14467), .Z(n11611) );
  NOR U12822 ( .A(n14468), .B(n14466), .Z(n14467) );
  XOR U12823 ( .A(n14469), .B(n14470), .Z(n11614) );
  NOR U12824 ( .A(n14471), .B(n14469), .Z(n14470) );
  XOR U12825 ( .A(n14472), .B(n14473), .Z(n11617) );
  NOR U12826 ( .A(n14474), .B(n14472), .Z(n14473) );
  XOR U12827 ( .A(n14475), .B(n14476), .Z(n11620) );
  NOR U12828 ( .A(n14477), .B(n14475), .Z(n14476) );
  XOR U12829 ( .A(n14478), .B(n14479), .Z(n11623) );
  NOR U12830 ( .A(n14480), .B(n14478), .Z(n14479) );
  XOR U12831 ( .A(n14481), .B(n14482), .Z(n11626) );
  NOR U12832 ( .A(n14483), .B(n14481), .Z(n14482) );
  XOR U12833 ( .A(n14484), .B(n14485), .Z(n11629) );
  NOR U12834 ( .A(n14486), .B(n14484), .Z(n14485) );
  XOR U12835 ( .A(n14487), .B(n14488), .Z(n11632) );
  NOR U12836 ( .A(n14489), .B(n14487), .Z(n14488) );
  XOR U12837 ( .A(n14490), .B(n14491), .Z(n11635) );
  NOR U12838 ( .A(n14492), .B(n14490), .Z(n14491) );
  XOR U12839 ( .A(n14493), .B(n14494), .Z(n11638) );
  NOR U12840 ( .A(n14495), .B(n14493), .Z(n14494) );
  XOR U12841 ( .A(n14496), .B(n14497), .Z(n11641) );
  NOR U12842 ( .A(n14498), .B(n14496), .Z(n14497) );
  XOR U12843 ( .A(n14499), .B(n14500), .Z(n11644) );
  NOR U12844 ( .A(n14501), .B(n14499), .Z(n14500) );
  XOR U12845 ( .A(n14502), .B(n14503), .Z(n11647) );
  NOR U12846 ( .A(n14504), .B(n14502), .Z(n14503) );
  XOR U12847 ( .A(n14505), .B(n14506), .Z(n11650) );
  NOR U12848 ( .A(n14507), .B(n14505), .Z(n14506) );
  XOR U12849 ( .A(n14508), .B(n14509), .Z(n11653) );
  NOR U12850 ( .A(n14510), .B(n14508), .Z(n14509) );
  XOR U12851 ( .A(n14511), .B(n14512), .Z(n11656) );
  NOR U12852 ( .A(n14513), .B(n14511), .Z(n14512) );
  XOR U12853 ( .A(n14514), .B(n14515), .Z(n11659) );
  NOR U12854 ( .A(n14516), .B(n14514), .Z(n14515) );
  XOR U12855 ( .A(n14517), .B(n14518), .Z(n11662) );
  NOR U12856 ( .A(n14519), .B(n14517), .Z(n14518) );
  XOR U12857 ( .A(n14520), .B(n14521), .Z(n11665) );
  NOR U12858 ( .A(n14522), .B(n14520), .Z(n14521) );
  XOR U12859 ( .A(n14523), .B(n14524), .Z(n11668) );
  NOR U12860 ( .A(n14525), .B(n14523), .Z(n14524) );
  XOR U12861 ( .A(n14526), .B(n14527), .Z(n11671) );
  NOR U12862 ( .A(n14528), .B(n14526), .Z(n14527) );
  XOR U12863 ( .A(n14529), .B(n14530), .Z(n11674) );
  NOR U12864 ( .A(n14531), .B(n14529), .Z(n14530) );
  XOR U12865 ( .A(n14532), .B(n14533), .Z(n11677) );
  NOR U12866 ( .A(n14534), .B(n14532), .Z(n14533) );
  XOR U12867 ( .A(n14535), .B(n14536), .Z(n11680) );
  NOR U12868 ( .A(n14537), .B(n14535), .Z(n14536) );
  XOR U12869 ( .A(n14538), .B(n14539), .Z(n11683) );
  NOR U12870 ( .A(n14540), .B(n14538), .Z(n14539) );
  XOR U12871 ( .A(n14541), .B(n14542), .Z(n11686) );
  NOR U12872 ( .A(n14543), .B(n14541), .Z(n14542) );
  XOR U12873 ( .A(n14544), .B(n14545), .Z(n11689) );
  NOR U12874 ( .A(n14546), .B(n14544), .Z(n14545) );
  XOR U12875 ( .A(n14547), .B(n14548), .Z(n11692) );
  NOR U12876 ( .A(n14549), .B(n14547), .Z(n14548) );
  XOR U12877 ( .A(n14550), .B(n14551), .Z(n11695) );
  NOR U12878 ( .A(n14552), .B(n14550), .Z(n14551) );
  XOR U12879 ( .A(n14553), .B(n14554), .Z(n11698) );
  NOR U12880 ( .A(n14555), .B(n14553), .Z(n14554) );
  XOR U12881 ( .A(n14556), .B(n14557), .Z(n11701) );
  NOR U12882 ( .A(n14558), .B(n14556), .Z(n14557) );
  XOR U12883 ( .A(n14559), .B(n14560), .Z(n11704) );
  NOR U12884 ( .A(n14561), .B(n14559), .Z(n14560) );
  XOR U12885 ( .A(n14562), .B(n14563), .Z(n11707) );
  NOR U12886 ( .A(n14564), .B(n14562), .Z(n14563) );
  XOR U12887 ( .A(n14565), .B(n14566), .Z(n11710) );
  NOR U12888 ( .A(n14567), .B(n14565), .Z(n14566) );
  XOR U12889 ( .A(n14568), .B(n14569), .Z(n11713) );
  NOR U12890 ( .A(n14570), .B(n14568), .Z(n14569) );
  XOR U12891 ( .A(n14571), .B(n14572), .Z(n11716) );
  NOR U12892 ( .A(n14573), .B(n14571), .Z(n14572) );
  XOR U12893 ( .A(n14574), .B(n14575), .Z(n11719) );
  NOR U12894 ( .A(n14576), .B(n14574), .Z(n14575) );
  XOR U12895 ( .A(n14577), .B(n14578), .Z(n11722) );
  NOR U12896 ( .A(n14579), .B(n14577), .Z(n14578) );
  XOR U12897 ( .A(n14580), .B(n14581), .Z(n11725) );
  NOR U12898 ( .A(n14582), .B(n14580), .Z(n14581) );
  XOR U12899 ( .A(n14583), .B(n14584), .Z(n11728) );
  NOR U12900 ( .A(n14585), .B(n14583), .Z(n14584) );
  XOR U12901 ( .A(n14586), .B(n14587), .Z(n11731) );
  NOR U12902 ( .A(n14588), .B(n14586), .Z(n14587) );
  XOR U12903 ( .A(n14589), .B(n14590), .Z(n11734) );
  NOR U12904 ( .A(n14591), .B(n14589), .Z(n14590) );
  XOR U12905 ( .A(n14592), .B(n14593), .Z(n11737) );
  NOR U12906 ( .A(n14594), .B(n14592), .Z(n14593) );
  XOR U12907 ( .A(n14595), .B(n14596), .Z(n11740) );
  NOR U12908 ( .A(n14597), .B(n14595), .Z(n14596) );
  XOR U12909 ( .A(n14598), .B(n14599), .Z(n11743) );
  NOR U12910 ( .A(n14600), .B(n14598), .Z(n14599) );
  XOR U12911 ( .A(n14601), .B(n14602), .Z(n11746) );
  NOR U12912 ( .A(n14603), .B(n14601), .Z(n14602) );
  XOR U12913 ( .A(n14604), .B(n14605), .Z(n11749) );
  NOR U12914 ( .A(n14606), .B(n14604), .Z(n14605) );
  XOR U12915 ( .A(n14607), .B(n14608), .Z(n11752) );
  NOR U12916 ( .A(n14609), .B(n14607), .Z(n14608) );
  XOR U12917 ( .A(n14610), .B(n14611), .Z(n11755) );
  NOR U12918 ( .A(n14612), .B(n14610), .Z(n14611) );
  XOR U12919 ( .A(n14613), .B(n14614), .Z(n11758) );
  NOR U12920 ( .A(n14615), .B(n14613), .Z(n14614) );
  XOR U12921 ( .A(n14616), .B(n14617), .Z(n11761) );
  NOR U12922 ( .A(n14618), .B(n14616), .Z(n14617) );
  XOR U12923 ( .A(n14619), .B(n14620), .Z(n11764) );
  NOR U12924 ( .A(n14621), .B(n14619), .Z(n14620) );
  XOR U12925 ( .A(n14622), .B(n14623), .Z(n11767) );
  NOR U12926 ( .A(n14624), .B(n14622), .Z(n14623) );
  XOR U12927 ( .A(n14625), .B(n14626), .Z(n11770) );
  NOR U12928 ( .A(n14627), .B(n14625), .Z(n14626) );
  XOR U12929 ( .A(n14628), .B(n14629), .Z(n11773) );
  NOR U12930 ( .A(n14630), .B(n14628), .Z(n14629) );
  XOR U12931 ( .A(n14631), .B(n14632), .Z(n11776) );
  NOR U12932 ( .A(n14633), .B(n14631), .Z(n14632) );
  XOR U12933 ( .A(n14634), .B(n14635), .Z(n11779) );
  NOR U12934 ( .A(n14636), .B(n14634), .Z(n14635) );
  XOR U12935 ( .A(n14637), .B(n14638), .Z(n11782) );
  NOR U12936 ( .A(n14639), .B(n14637), .Z(n14638) );
  XOR U12937 ( .A(n14640), .B(n14641), .Z(n11785) );
  NOR U12938 ( .A(n14642), .B(n14640), .Z(n14641) );
  XOR U12939 ( .A(n14643), .B(n14644), .Z(n11788) );
  NOR U12940 ( .A(n14645), .B(n14643), .Z(n14644) );
  XOR U12941 ( .A(n14646), .B(n14647), .Z(n11791) );
  NOR U12942 ( .A(n14648), .B(n14646), .Z(n14647) );
  XOR U12943 ( .A(n14649), .B(n14650), .Z(n11794) );
  NOR U12944 ( .A(n14651), .B(n14649), .Z(n14650) );
  XOR U12945 ( .A(n14652), .B(n14653), .Z(n11797) );
  NOR U12946 ( .A(n14654), .B(n14652), .Z(n14653) );
  XOR U12947 ( .A(n14655), .B(n14656), .Z(n11800) );
  NOR U12948 ( .A(n14657), .B(n14655), .Z(n14656) );
  XOR U12949 ( .A(n14658), .B(n14659), .Z(n11803) );
  NOR U12950 ( .A(n14660), .B(n14658), .Z(n14659) );
  XOR U12951 ( .A(n14661), .B(n14662), .Z(n11806) );
  NOR U12952 ( .A(n14663), .B(n14661), .Z(n14662) );
  XOR U12953 ( .A(n14664), .B(n14665), .Z(n11809) );
  NOR U12954 ( .A(n14666), .B(n14664), .Z(n14665) );
  XOR U12955 ( .A(n14667), .B(n14668), .Z(n11812) );
  NOR U12956 ( .A(n14669), .B(n14667), .Z(n14668) );
  XOR U12957 ( .A(n14670), .B(n14671), .Z(n11815) );
  NOR U12958 ( .A(n14672), .B(n14670), .Z(n14671) );
  XOR U12959 ( .A(n14673), .B(n14674), .Z(n11818) );
  NOR U12960 ( .A(n14675), .B(n14673), .Z(n14674) );
  XOR U12961 ( .A(n14676), .B(n14677), .Z(n11821) );
  NOR U12962 ( .A(n14678), .B(n14676), .Z(n14677) );
  XOR U12963 ( .A(n14679), .B(n14680), .Z(n11824) );
  NOR U12964 ( .A(n14681), .B(n14679), .Z(n14680) );
  XOR U12965 ( .A(n14682), .B(n14683), .Z(n11827) );
  NOR U12966 ( .A(n14684), .B(n14682), .Z(n14683) );
  XOR U12967 ( .A(n14685), .B(n14686), .Z(n11830) );
  NOR U12968 ( .A(n14687), .B(n14685), .Z(n14686) );
  XOR U12969 ( .A(n14688), .B(n14689), .Z(n11833) );
  NOR U12970 ( .A(n14690), .B(n14688), .Z(n14689) );
  XOR U12971 ( .A(n14691), .B(n14692), .Z(n11836) );
  NOR U12972 ( .A(n14693), .B(n14691), .Z(n14692) );
  XOR U12973 ( .A(n14694), .B(n14695), .Z(n11839) );
  NOR U12974 ( .A(n14696), .B(n14694), .Z(n14695) );
  XOR U12975 ( .A(n14697), .B(n14698), .Z(n11842) );
  NOR U12976 ( .A(n14699), .B(n14697), .Z(n14698) );
  XOR U12977 ( .A(n14700), .B(n14701), .Z(n11845) );
  NOR U12978 ( .A(n14702), .B(n14700), .Z(n14701) );
  XOR U12979 ( .A(n14703), .B(n14704), .Z(n11848) );
  NOR U12980 ( .A(n14705), .B(n14703), .Z(n14704) );
  XOR U12981 ( .A(n14706), .B(n14707), .Z(n11851) );
  NOR U12982 ( .A(n14708), .B(n14706), .Z(n14707) );
  XOR U12983 ( .A(n14709), .B(n14710), .Z(n11854) );
  NOR U12984 ( .A(n14711), .B(n14709), .Z(n14710) );
  XOR U12985 ( .A(n14712), .B(n14713), .Z(n11857) );
  NOR U12986 ( .A(n14714), .B(n14712), .Z(n14713) );
  XOR U12987 ( .A(n14715), .B(n14716), .Z(n11860) );
  NOR U12988 ( .A(n14717), .B(n14715), .Z(n14716) );
  XOR U12989 ( .A(n14718), .B(n14719), .Z(n11863) );
  NOR U12990 ( .A(n14720), .B(n14718), .Z(n14719) );
  XOR U12991 ( .A(n14721), .B(n14722), .Z(n11866) );
  NOR U12992 ( .A(n14723), .B(n14721), .Z(n14722) );
  XOR U12993 ( .A(n14724), .B(n14725), .Z(n11869) );
  NOR U12994 ( .A(n14726), .B(n14724), .Z(n14725) );
  XOR U12995 ( .A(n14727), .B(n14728), .Z(n11872) );
  NOR U12996 ( .A(n14729), .B(n14727), .Z(n14728) );
  XOR U12997 ( .A(n14730), .B(n14731), .Z(n11875) );
  NOR U12998 ( .A(n14732), .B(n14730), .Z(n14731) );
  XOR U12999 ( .A(n14733), .B(n14734), .Z(n11878) );
  NOR U13000 ( .A(n14735), .B(n14733), .Z(n14734) );
  XOR U13001 ( .A(n14736), .B(n14737), .Z(n11881) );
  NOR U13002 ( .A(n14738), .B(n14736), .Z(n14737) );
  XOR U13003 ( .A(n14739), .B(n14740), .Z(n11884) );
  NOR U13004 ( .A(n14741), .B(n14739), .Z(n14740) );
  XOR U13005 ( .A(n14742), .B(n14743), .Z(n11887) );
  NOR U13006 ( .A(n14744), .B(n14742), .Z(n14743) );
  XOR U13007 ( .A(n14745), .B(n14746), .Z(n11890) );
  NOR U13008 ( .A(n14747), .B(n14745), .Z(n14746) );
  XOR U13009 ( .A(n14748), .B(n14749), .Z(n11893) );
  NOR U13010 ( .A(n14750), .B(n14748), .Z(n14749) );
  XOR U13011 ( .A(n14751), .B(n14752), .Z(n11896) );
  NOR U13012 ( .A(n14753), .B(n14751), .Z(n14752) );
  XOR U13013 ( .A(n14754), .B(n14755), .Z(n11899) );
  NOR U13014 ( .A(n14756), .B(n14754), .Z(n14755) );
  XOR U13015 ( .A(n14757), .B(n14758), .Z(n11902) );
  NOR U13016 ( .A(n14759), .B(n14757), .Z(n14758) );
  XOR U13017 ( .A(n14760), .B(n14761), .Z(n11905) );
  NOR U13018 ( .A(n14762), .B(n14760), .Z(n14761) );
  XOR U13019 ( .A(n14763), .B(n14764), .Z(n11908) );
  NOR U13020 ( .A(n14765), .B(n14763), .Z(n14764) );
  XOR U13021 ( .A(n14766), .B(n14767), .Z(n11911) );
  NOR U13022 ( .A(n14768), .B(n14766), .Z(n14767) );
  XOR U13023 ( .A(n14769), .B(n14770), .Z(n11914) );
  NOR U13024 ( .A(n14771), .B(n14769), .Z(n14770) );
  XOR U13025 ( .A(n14772), .B(n14773), .Z(n11917) );
  NOR U13026 ( .A(n14774), .B(n14772), .Z(n14773) );
  XOR U13027 ( .A(n14775), .B(n14776), .Z(n11920) );
  NOR U13028 ( .A(n14777), .B(n14775), .Z(n14776) );
  XOR U13029 ( .A(n14778), .B(n14779), .Z(n11923) );
  NOR U13030 ( .A(n14780), .B(n14778), .Z(n14779) );
  XOR U13031 ( .A(n14781), .B(n14782), .Z(n11926) );
  NOR U13032 ( .A(n14783), .B(n14781), .Z(n14782) );
  XOR U13033 ( .A(n14784), .B(n14785), .Z(n11929) );
  NOR U13034 ( .A(n14786), .B(n14784), .Z(n14785) );
  XOR U13035 ( .A(n14787), .B(n14788), .Z(n11932) );
  NOR U13036 ( .A(n14789), .B(n14787), .Z(n14788) );
  XOR U13037 ( .A(n14790), .B(n14791), .Z(n11935) );
  NOR U13038 ( .A(n14792), .B(n14790), .Z(n14791) );
  XOR U13039 ( .A(n14793), .B(n14794), .Z(n11938) );
  NOR U13040 ( .A(n14795), .B(n14793), .Z(n14794) );
  XOR U13041 ( .A(n14796), .B(n14797), .Z(n11941) );
  NOR U13042 ( .A(n14798), .B(n14796), .Z(n14797) );
  XOR U13043 ( .A(n14799), .B(n14800), .Z(n11944) );
  NOR U13044 ( .A(n14801), .B(n14799), .Z(n14800) );
  XOR U13045 ( .A(n14802), .B(n14803), .Z(n11947) );
  NOR U13046 ( .A(n14804), .B(n14802), .Z(n14803) );
  XOR U13047 ( .A(n14805), .B(n14806), .Z(n11950) );
  NOR U13048 ( .A(n14807), .B(n14805), .Z(n14806) );
  XOR U13049 ( .A(n14808), .B(n14809), .Z(n11953) );
  NOR U13050 ( .A(n14810), .B(n14808), .Z(n14809) );
  XOR U13051 ( .A(n14811), .B(n14812), .Z(n11956) );
  NOR U13052 ( .A(n14813), .B(n14811), .Z(n14812) );
  XOR U13053 ( .A(n14814), .B(n14815), .Z(n11959) );
  NOR U13054 ( .A(n14816), .B(n14814), .Z(n14815) );
  XOR U13055 ( .A(n14817), .B(n14818), .Z(n11962) );
  NOR U13056 ( .A(n14819), .B(n14817), .Z(n14818) );
  XOR U13057 ( .A(n14820), .B(n14821), .Z(n11965) );
  NOR U13058 ( .A(n14822), .B(n14820), .Z(n14821) );
  XOR U13059 ( .A(n14823), .B(n14824), .Z(n11968) );
  NOR U13060 ( .A(n14825), .B(n14823), .Z(n14824) );
  XOR U13061 ( .A(n14826), .B(n14827), .Z(n11971) );
  NOR U13062 ( .A(n14828), .B(n14826), .Z(n14827) );
  XOR U13063 ( .A(n14829), .B(n14830), .Z(n11974) );
  NOR U13064 ( .A(n14831), .B(n14829), .Z(n14830) );
  XOR U13065 ( .A(n14832), .B(n14833), .Z(n11977) );
  NOR U13066 ( .A(n14834), .B(n14832), .Z(n14833) );
  XOR U13067 ( .A(n14835), .B(n14836), .Z(n11980) );
  NOR U13068 ( .A(n14837), .B(n14835), .Z(n14836) );
  XOR U13069 ( .A(n14838), .B(n14839), .Z(n11983) );
  NOR U13070 ( .A(n14840), .B(n14838), .Z(n14839) );
  XOR U13071 ( .A(n14841), .B(n14842), .Z(n11986) );
  NOR U13072 ( .A(n14843), .B(n14841), .Z(n14842) );
  XOR U13073 ( .A(n14844), .B(n14845), .Z(n11989) );
  NOR U13074 ( .A(n14846), .B(n14844), .Z(n14845) );
  XOR U13075 ( .A(n14847), .B(n14848), .Z(n11992) );
  NOR U13076 ( .A(n14849), .B(n14847), .Z(n14848) );
  XOR U13077 ( .A(n14850), .B(n14851), .Z(n11995) );
  NOR U13078 ( .A(n14852), .B(n14850), .Z(n14851) );
  XOR U13079 ( .A(n14853), .B(n14854), .Z(n11998) );
  NOR U13080 ( .A(n14855), .B(n14853), .Z(n14854) );
  XOR U13081 ( .A(n14856), .B(n14857), .Z(n12001) );
  NOR U13082 ( .A(n14858), .B(n14856), .Z(n14857) );
  XOR U13083 ( .A(n14859), .B(n14860), .Z(n12004) );
  NOR U13084 ( .A(n14861), .B(n14859), .Z(n14860) );
  XOR U13085 ( .A(n14862), .B(n14863), .Z(n12007) );
  NOR U13086 ( .A(n14864), .B(n14862), .Z(n14863) );
  XOR U13087 ( .A(n14865), .B(n14866), .Z(n12010) );
  NOR U13088 ( .A(n14867), .B(n14865), .Z(n14866) );
  XOR U13089 ( .A(n14868), .B(n14869), .Z(n12013) );
  NOR U13090 ( .A(n14870), .B(n14868), .Z(n14869) );
  XOR U13091 ( .A(n14871), .B(n14872), .Z(n12016) );
  NOR U13092 ( .A(n14873), .B(n14871), .Z(n14872) );
  XOR U13093 ( .A(n14874), .B(n14875), .Z(n12019) );
  NOR U13094 ( .A(n14876), .B(n14874), .Z(n14875) );
  XOR U13095 ( .A(n14877), .B(n14878), .Z(n12022) );
  NOR U13096 ( .A(n14879), .B(n14877), .Z(n14878) );
  XOR U13097 ( .A(n14880), .B(n14881), .Z(n12025) );
  NOR U13098 ( .A(n14882), .B(n14880), .Z(n14881) );
  XOR U13099 ( .A(n14883), .B(n14884), .Z(n12028) );
  NOR U13100 ( .A(n14885), .B(n14883), .Z(n14884) );
  XOR U13101 ( .A(n14886), .B(n14887), .Z(n12031) );
  NOR U13102 ( .A(n14888), .B(n14886), .Z(n14887) );
  XOR U13103 ( .A(n14889), .B(n14890), .Z(n12034) );
  NOR U13104 ( .A(n14891), .B(n14889), .Z(n14890) );
  XOR U13105 ( .A(n14892), .B(n14893), .Z(n12037) );
  NOR U13106 ( .A(n14894), .B(n14892), .Z(n14893) );
  XOR U13107 ( .A(n14895), .B(n14896), .Z(n12040) );
  NOR U13108 ( .A(n14897), .B(n14895), .Z(n14896) );
  XOR U13109 ( .A(n14898), .B(n14899), .Z(n12043) );
  NOR U13110 ( .A(n14900), .B(n14898), .Z(n14899) );
  XOR U13111 ( .A(n14901), .B(n14902), .Z(n12046) );
  NOR U13112 ( .A(n14903), .B(n14901), .Z(n14902) );
  XOR U13113 ( .A(n14904), .B(n14905), .Z(n12049) );
  NOR U13114 ( .A(n14906), .B(n14904), .Z(n14905) );
  XOR U13115 ( .A(n14907), .B(n14908), .Z(n12052) );
  NOR U13116 ( .A(n14909), .B(n14907), .Z(n14908) );
  XOR U13117 ( .A(n14910), .B(n14911), .Z(n12055) );
  NOR U13118 ( .A(n14912), .B(n14910), .Z(n14911) );
  XOR U13119 ( .A(n14913), .B(n14914), .Z(n12058) );
  NOR U13120 ( .A(n14915), .B(n14913), .Z(n14914) );
  XOR U13121 ( .A(n14916), .B(n14917), .Z(n12061) );
  NOR U13122 ( .A(n14918), .B(n14916), .Z(n14917) );
  XOR U13123 ( .A(n14919), .B(n14920), .Z(n12064) );
  NOR U13124 ( .A(n14921), .B(n14919), .Z(n14920) );
  XOR U13125 ( .A(n14922), .B(n14923), .Z(n12067) );
  NOR U13126 ( .A(n14924), .B(n14922), .Z(n14923) );
  XOR U13127 ( .A(n14925), .B(n14926), .Z(n12070) );
  NOR U13128 ( .A(n14927), .B(n14925), .Z(n14926) );
  XOR U13129 ( .A(n14928), .B(n14929), .Z(n12073) );
  NOR U13130 ( .A(n14930), .B(n14928), .Z(n14929) );
  XOR U13131 ( .A(n14931), .B(n14932), .Z(n12076) );
  NOR U13132 ( .A(n14933), .B(n14931), .Z(n14932) );
  XOR U13133 ( .A(n14934), .B(n14935), .Z(n12079) );
  NOR U13134 ( .A(n14936), .B(n14934), .Z(n14935) );
  XOR U13135 ( .A(n14937), .B(n14938), .Z(n12082) );
  NOR U13136 ( .A(n14939), .B(n14937), .Z(n14938) );
  XOR U13137 ( .A(n14940), .B(n14941), .Z(n12085) );
  NOR U13138 ( .A(n14942), .B(n14940), .Z(n14941) );
  XOR U13139 ( .A(n14943), .B(n14944), .Z(n12088) );
  NOR U13140 ( .A(n14945), .B(n14943), .Z(n14944) );
  XOR U13141 ( .A(n14946), .B(n14947), .Z(n12091) );
  NOR U13142 ( .A(n14948), .B(n14946), .Z(n14947) );
  XOR U13143 ( .A(n14949), .B(n14950), .Z(n12094) );
  NOR U13144 ( .A(n14951), .B(n14949), .Z(n14950) );
  XOR U13145 ( .A(n14952), .B(n14953), .Z(n12097) );
  NOR U13146 ( .A(n14954), .B(n14952), .Z(n14953) );
  XOR U13147 ( .A(n14955), .B(n14956), .Z(n12100) );
  NOR U13148 ( .A(n14957), .B(n14955), .Z(n14956) );
  XOR U13149 ( .A(n14958), .B(n14959), .Z(n12103) );
  NOR U13150 ( .A(n14960), .B(n14958), .Z(n14959) );
  XOR U13151 ( .A(n14961), .B(n14962), .Z(n12106) );
  NOR U13152 ( .A(n14963), .B(n14961), .Z(n14962) );
  XOR U13153 ( .A(n14964), .B(n14965), .Z(n12109) );
  NOR U13154 ( .A(n14966), .B(n14964), .Z(n14965) );
  XOR U13155 ( .A(n14967), .B(n14968), .Z(n12112) );
  NOR U13156 ( .A(n14969), .B(n14967), .Z(n14968) );
  XOR U13157 ( .A(n14970), .B(n14971), .Z(n12115) );
  NOR U13158 ( .A(n14972), .B(n14970), .Z(n14971) );
  XOR U13159 ( .A(n14973), .B(n14974), .Z(n12118) );
  NOR U13160 ( .A(n14975), .B(n14973), .Z(n14974) );
  XOR U13161 ( .A(n14976), .B(n14977), .Z(n12121) );
  NOR U13162 ( .A(n14978), .B(n14976), .Z(n14977) );
  XOR U13163 ( .A(n14979), .B(n14980), .Z(n12124) );
  NOR U13164 ( .A(n14981), .B(n14979), .Z(n14980) );
  XOR U13165 ( .A(n14982), .B(n14983), .Z(n12127) );
  NOR U13166 ( .A(n14984), .B(n14982), .Z(n14983) );
  XOR U13167 ( .A(n14985), .B(n14986), .Z(n12130) );
  NOR U13168 ( .A(n14987), .B(n14985), .Z(n14986) );
  XOR U13169 ( .A(n14988), .B(n14989), .Z(n12133) );
  NOR U13170 ( .A(n14990), .B(n14988), .Z(n14989) );
  XOR U13171 ( .A(n14991), .B(n14992), .Z(n12136) );
  NOR U13172 ( .A(n14993), .B(n14991), .Z(n14992) );
  XOR U13173 ( .A(n14994), .B(n14995), .Z(n12139) );
  NOR U13174 ( .A(n14996), .B(n14994), .Z(n14995) );
  XOR U13175 ( .A(n14997), .B(n14998), .Z(n12142) );
  NOR U13176 ( .A(n14999), .B(n14997), .Z(n14998) );
  XOR U13177 ( .A(n15000), .B(n15001), .Z(n12145) );
  NOR U13178 ( .A(n15002), .B(n15000), .Z(n15001) );
  XOR U13179 ( .A(n15003), .B(n15004), .Z(n12148) );
  NOR U13180 ( .A(n15005), .B(n15003), .Z(n15004) );
  XOR U13181 ( .A(n15006), .B(n15007), .Z(n12151) );
  NOR U13182 ( .A(n15008), .B(n15006), .Z(n15007) );
  XOR U13183 ( .A(n15009), .B(n15010), .Z(n12154) );
  NOR U13184 ( .A(n15011), .B(n15009), .Z(n15010) );
  XOR U13185 ( .A(n15012), .B(n15013), .Z(n12157) );
  NOR U13186 ( .A(n15014), .B(n15012), .Z(n15013) );
  XOR U13187 ( .A(n15015), .B(n15016), .Z(n12160) );
  NOR U13188 ( .A(n15017), .B(n15015), .Z(n15016) );
  XOR U13189 ( .A(n15018), .B(n15019), .Z(n12163) );
  NOR U13190 ( .A(n15020), .B(n15018), .Z(n15019) );
  XOR U13191 ( .A(n15021), .B(n15022), .Z(n12166) );
  NOR U13192 ( .A(n15023), .B(n15021), .Z(n15022) );
  XOR U13193 ( .A(n15024), .B(n15025), .Z(n12169) );
  NOR U13194 ( .A(n15026), .B(n15024), .Z(n15025) );
  XOR U13195 ( .A(n15027), .B(n15028), .Z(n12172) );
  NOR U13196 ( .A(n15029), .B(n15027), .Z(n15028) );
  XOR U13197 ( .A(n15030), .B(n15031), .Z(n12175) );
  NOR U13198 ( .A(n15032), .B(n15030), .Z(n15031) );
  XOR U13199 ( .A(n15033), .B(n15034), .Z(n12178) );
  NOR U13200 ( .A(n15035), .B(n15033), .Z(n15034) );
  XOR U13201 ( .A(n15036), .B(n15037), .Z(n12181) );
  NOR U13202 ( .A(n15038), .B(n15036), .Z(n15037) );
  XOR U13203 ( .A(n15039), .B(n15040), .Z(n12184) );
  NOR U13204 ( .A(n15041), .B(n15039), .Z(n15040) );
  XOR U13205 ( .A(n15042), .B(n15043), .Z(n12187) );
  NOR U13206 ( .A(n15044), .B(n15042), .Z(n15043) );
  XOR U13207 ( .A(n15045), .B(n15046), .Z(n12190) );
  NOR U13208 ( .A(n15047), .B(n15045), .Z(n15046) );
  XOR U13209 ( .A(n15048), .B(n15049), .Z(n12193) );
  NOR U13210 ( .A(n15050), .B(n15048), .Z(n15049) );
  XOR U13211 ( .A(n15051), .B(n15052), .Z(n12196) );
  NOR U13212 ( .A(n15053), .B(n15051), .Z(n15052) );
  XOR U13213 ( .A(n15054), .B(n15055), .Z(n12199) );
  NOR U13214 ( .A(n15056), .B(n15054), .Z(n15055) );
  XOR U13215 ( .A(n15057), .B(n15058), .Z(n12202) );
  NOR U13216 ( .A(n15059), .B(n15057), .Z(n15058) );
  XOR U13217 ( .A(n15060), .B(n15061), .Z(n12205) );
  NOR U13218 ( .A(n15062), .B(n15060), .Z(n15061) );
  XOR U13219 ( .A(n15063), .B(n15064), .Z(n12208) );
  NOR U13220 ( .A(n15065), .B(n15063), .Z(n15064) );
  XOR U13221 ( .A(n15066), .B(n15067), .Z(n12211) );
  NOR U13222 ( .A(n15068), .B(n15066), .Z(n15067) );
  XOR U13223 ( .A(n15069), .B(n15070), .Z(n12214) );
  NOR U13224 ( .A(n15071), .B(n15069), .Z(n15070) );
  XOR U13225 ( .A(n15072), .B(n15073), .Z(n12217) );
  NOR U13226 ( .A(n15074), .B(n15072), .Z(n15073) );
  XOR U13227 ( .A(n15075), .B(n15076), .Z(n12220) );
  NOR U13228 ( .A(n15077), .B(n15075), .Z(n15076) );
  XOR U13229 ( .A(n15078), .B(n15079), .Z(n12223) );
  NOR U13230 ( .A(n15080), .B(n15078), .Z(n15079) );
  XOR U13231 ( .A(n15081), .B(n15082), .Z(n12226) );
  NOR U13232 ( .A(n15083), .B(n15081), .Z(n15082) );
  XOR U13233 ( .A(n15084), .B(n15085), .Z(n12229) );
  NOR U13234 ( .A(n15086), .B(n15084), .Z(n15085) );
  XOR U13235 ( .A(n15087), .B(n15088), .Z(n12232) );
  NOR U13236 ( .A(n15089), .B(n15087), .Z(n15088) );
  XOR U13237 ( .A(n15090), .B(n15091), .Z(n12235) );
  NOR U13238 ( .A(n15092), .B(n15090), .Z(n15091) );
  XOR U13239 ( .A(n15093), .B(n15094), .Z(n12238) );
  NOR U13240 ( .A(n15095), .B(n15093), .Z(n15094) );
  XOR U13241 ( .A(n15096), .B(n15097), .Z(n12241) );
  NOR U13242 ( .A(n15098), .B(n15096), .Z(n15097) );
  XOR U13243 ( .A(n15099), .B(n15100), .Z(n12244) );
  NOR U13244 ( .A(n15101), .B(n15099), .Z(n15100) );
  XOR U13245 ( .A(n15102), .B(n15103), .Z(n12247) );
  NOR U13246 ( .A(n15104), .B(n15102), .Z(n15103) );
  XOR U13247 ( .A(n15105), .B(n15106), .Z(n12250) );
  NOR U13248 ( .A(n15107), .B(n15105), .Z(n15106) );
  XOR U13249 ( .A(n15108), .B(n15109), .Z(n12253) );
  NOR U13250 ( .A(n15110), .B(n15108), .Z(n15109) );
  XOR U13251 ( .A(n15111), .B(n15112), .Z(n12256) );
  NOR U13252 ( .A(n15113), .B(n15111), .Z(n15112) );
  XOR U13253 ( .A(n15114), .B(n15115), .Z(n12259) );
  NOR U13254 ( .A(n15116), .B(n15114), .Z(n15115) );
  XOR U13255 ( .A(n15117), .B(n15118), .Z(n12262) );
  NOR U13256 ( .A(n15119), .B(n15117), .Z(n15118) );
  XOR U13257 ( .A(n15120), .B(n15121), .Z(n12265) );
  NOR U13258 ( .A(n15122), .B(n15120), .Z(n15121) );
  XOR U13259 ( .A(n15123), .B(n15124), .Z(n12268) );
  NOR U13260 ( .A(n15125), .B(n15123), .Z(n15124) );
  XOR U13261 ( .A(n15126), .B(n15127), .Z(n12271) );
  NOR U13262 ( .A(n15128), .B(n15126), .Z(n15127) );
  XOR U13263 ( .A(n15129), .B(n15130), .Z(n12274) );
  NOR U13264 ( .A(n15131), .B(n15129), .Z(n15130) );
  XOR U13265 ( .A(n15132), .B(n15133), .Z(n12277) );
  NOR U13266 ( .A(n15134), .B(n15132), .Z(n15133) );
  XOR U13267 ( .A(n15135), .B(n15136), .Z(n12280) );
  NOR U13268 ( .A(n15137), .B(n15135), .Z(n15136) );
  XOR U13269 ( .A(n15138), .B(n15139), .Z(n12283) );
  NOR U13270 ( .A(n15140), .B(n15138), .Z(n15139) );
  XOR U13271 ( .A(n15141), .B(n15142), .Z(n12286) );
  NOR U13272 ( .A(n15143), .B(n15141), .Z(n15142) );
  XOR U13273 ( .A(n15144), .B(n15145), .Z(n12289) );
  NOR U13274 ( .A(n15146), .B(n15144), .Z(n15145) );
  XOR U13275 ( .A(n15147), .B(n15148), .Z(n12292) );
  NOR U13276 ( .A(n15149), .B(n15147), .Z(n15148) );
  XOR U13277 ( .A(n15150), .B(n15151), .Z(n12295) );
  NOR U13278 ( .A(n15152), .B(n15150), .Z(n15151) );
  XOR U13279 ( .A(n15153), .B(n15154), .Z(n12298) );
  NOR U13280 ( .A(n15155), .B(n15153), .Z(n15154) );
  XOR U13281 ( .A(n15156), .B(n15157), .Z(n12301) );
  NOR U13282 ( .A(n15158), .B(n15156), .Z(n15157) );
  XOR U13283 ( .A(n15159), .B(n15160), .Z(n12304) );
  NOR U13284 ( .A(n15161), .B(n15159), .Z(n15160) );
  XOR U13285 ( .A(n15162), .B(n15163), .Z(n12307) );
  NOR U13286 ( .A(n15164), .B(n15162), .Z(n15163) );
  XOR U13287 ( .A(n15165), .B(n15166), .Z(n12310) );
  NOR U13288 ( .A(n15167), .B(n15165), .Z(n15166) );
  XOR U13289 ( .A(n15168), .B(n15169), .Z(n12313) );
  NOR U13290 ( .A(n15170), .B(n15168), .Z(n15169) );
  XOR U13291 ( .A(n15171), .B(n15172), .Z(n12316) );
  NOR U13292 ( .A(n15173), .B(n15171), .Z(n15172) );
  XOR U13293 ( .A(n15174), .B(n15175), .Z(n12319) );
  NOR U13294 ( .A(n15176), .B(n15174), .Z(n15175) );
  XOR U13295 ( .A(n15177), .B(n15178), .Z(n12322) );
  NOR U13296 ( .A(n15179), .B(n15177), .Z(n15178) );
  XOR U13297 ( .A(n15180), .B(n15181), .Z(n12325) );
  NOR U13298 ( .A(n15182), .B(n15180), .Z(n15181) );
  XOR U13299 ( .A(n15183), .B(n15184), .Z(n12328) );
  NOR U13300 ( .A(n15185), .B(n15183), .Z(n15184) );
  XOR U13301 ( .A(n15186), .B(n15187), .Z(n12331) );
  NOR U13302 ( .A(n15188), .B(n15186), .Z(n15187) );
  XOR U13303 ( .A(n15189), .B(n15190), .Z(n12334) );
  NOR U13304 ( .A(n15191), .B(n15189), .Z(n15190) );
  XOR U13305 ( .A(n15192), .B(n15193), .Z(n12337) );
  NOR U13306 ( .A(n15194), .B(n15192), .Z(n15193) );
  XOR U13307 ( .A(n15195), .B(n15196), .Z(n12340) );
  NOR U13308 ( .A(n15197), .B(n15195), .Z(n15196) );
  XOR U13309 ( .A(n15198), .B(n15199), .Z(n12343) );
  NOR U13310 ( .A(n15200), .B(n15198), .Z(n15199) );
  XOR U13311 ( .A(n15201), .B(n15202), .Z(n12346) );
  NOR U13312 ( .A(n15203), .B(n15201), .Z(n15202) );
  XOR U13313 ( .A(n15204), .B(n15205), .Z(n12349) );
  NOR U13314 ( .A(n15206), .B(n15204), .Z(n15205) );
  XOR U13315 ( .A(n15207), .B(n15208), .Z(n12352) );
  NOR U13316 ( .A(n15209), .B(n15207), .Z(n15208) );
  XOR U13317 ( .A(n15210), .B(n15211), .Z(n12355) );
  NOR U13318 ( .A(n15212), .B(n15210), .Z(n15211) );
  XOR U13319 ( .A(n15213), .B(n15214), .Z(n12358) );
  NOR U13320 ( .A(n15215), .B(n15213), .Z(n15214) );
  XOR U13321 ( .A(n15216), .B(n15217), .Z(n12361) );
  NOR U13322 ( .A(n15218), .B(n15216), .Z(n15217) );
  XOR U13323 ( .A(n15219), .B(n15220), .Z(n12364) );
  NOR U13324 ( .A(n15221), .B(n15219), .Z(n15220) );
  XOR U13325 ( .A(n15222), .B(n15223), .Z(n12367) );
  NOR U13326 ( .A(n15224), .B(n15222), .Z(n15223) );
  XOR U13327 ( .A(n15225), .B(n15226), .Z(n12370) );
  NOR U13328 ( .A(n15227), .B(n15225), .Z(n15226) );
  XOR U13329 ( .A(n15228), .B(n15229), .Z(n12373) );
  NOR U13330 ( .A(n15230), .B(n15228), .Z(n15229) );
  XOR U13331 ( .A(n15231), .B(n15232), .Z(n12376) );
  NOR U13332 ( .A(n15233), .B(n15231), .Z(n15232) );
  XOR U13333 ( .A(n15234), .B(n15235), .Z(n12379) );
  NOR U13334 ( .A(n15236), .B(n15234), .Z(n15235) );
  XOR U13335 ( .A(n15237), .B(n15238), .Z(n12382) );
  NOR U13336 ( .A(n15239), .B(n15237), .Z(n15238) );
  XOR U13337 ( .A(n15240), .B(n15241), .Z(n12385) );
  NOR U13338 ( .A(n15242), .B(n15240), .Z(n15241) );
  XOR U13339 ( .A(n15243), .B(n15244), .Z(n12388) );
  NOR U13340 ( .A(n15245), .B(n15243), .Z(n15244) );
  XOR U13341 ( .A(n15246), .B(n15247), .Z(n12391) );
  NOR U13342 ( .A(n15248), .B(n15246), .Z(n15247) );
  XOR U13343 ( .A(n15249), .B(n15250), .Z(n12394) );
  NOR U13344 ( .A(n15251), .B(n15249), .Z(n15250) );
  XOR U13345 ( .A(n15252), .B(n15253), .Z(n12397) );
  NOR U13346 ( .A(n15254), .B(n15252), .Z(n15253) );
  XOR U13347 ( .A(n15255), .B(n15256), .Z(n12400) );
  NOR U13348 ( .A(n15257), .B(n15255), .Z(n15256) );
  XOR U13349 ( .A(n15258), .B(n15259), .Z(n12403) );
  NOR U13350 ( .A(n15260), .B(n15258), .Z(n15259) );
  XOR U13351 ( .A(n15261), .B(n15262), .Z(n12406) );
  NOR U13352 ( .A(n15263), .B(n15261), .Z(n15262) );
  XOR U13353 ( .A(n15264), .B(n15265), .Z(n12409) );
  NOR U13354 ( .A(n15266), .B(n15264), .Z(n15265) );
  XOR U13355 ( .A(n15267), .B(n15268), .Z(n12412) );
  NOR U13356 ( .A(n15269), .B(n15267), .Z(n15268) );
  XOR U13357 ( .A(n15270), .B(n15271), .Z(n12415) );
  NOR U13358 ( .A(n15272), .B(n15270), .Z(n15271) );
  XOR U13359 ( .A(n15273), .B(n15274), .Z(n12418) );
  NOR U13360 ( .A(n15275), .B(n15273), .Z(n15274) );
  XOR U13361 ( .A(n15276), .B(n15277), .Z(n12421) );
  NOR U13362 ( .A(n15278), .B(n15276), .Z(n15277) );
  XOR U13363 ( .A(n15279), .B(n15280), .Z(n12424) );
  NOR U13364 ( .A(n15281), .B(n15279), .Z(n15280) );
  XOR U13365 ( .A(n15282), .B(n15283), .Z(n12427) );
  NOR U13366 ( .A(n15284), .B(n15282), .Z(n15283) );
  XOR U13367 ( .A(n15285), .B(n15286), .Z(n12430) );
  NOR U13368 ( .A(n15287), .B(n15285), .Z(n15286) );
  XOR U13369 ( .A(n15288), .B(n15289), .Z(n12433) );
  NOR U13370 ( .A(n15290), .B(n15288), .Z(n15289) );
  XOR U13371 ( .A(n15291), .B(n15292), .Z(n12436) );
  NOR U13372 ( .A(n15293), .B(n15291), .Z(n15292) );
  XOR U13373 ( .A(n15294), .B(n15295), .Z(n12439) );
  NOR U13374 ( .A(n15296), .B(n15294), .Z(n15295) );
  XOR U13375 ( .A(n15297), .B(n15298), .Z(n12442) );
  NOR U13376 ( .A(n15299), .B(n15297), .Z(n15298) );
  XOR U13377 ( .A(n15300), .B(n15301), .Z(n12445) );
  NOR U13378 ( .A(n15302), .B(n15300), .Z(n15301) );
  XOR U13379 ( .A(n15303), .B(n15304), .Z(n12448) );
  NOR U13380 ( .A(n15305), .B(n15303), .Z(n15304) );
  XOR U13381 ( .A(n15306), .B(n15307), .Z(n12451) );
  NOR U13382 ( .A(n15308), .B(n15306), .Z(n15307) );
  XOR U13383 ( .A(n15309), .B(n15310), .Z(n12454) );
  NOR U13384 ( .A(n15311), .B(n15309), .Z(n15310) );
  XOR U13385 ( .A(n15312), .B(n15313), .Z(n12457) );
  NOR U13386 ( .A(n15314), .B(n15312), .Z(n15313) );
  XOR U13387 ( .A(n15315), .B(n15316), .Z(n12460) );
  NOR U13388 ( .A(n15317), .B(n15315), .Z(n15316) );
  XOR U13389 ( .A(n15318), .B(n15319), .Z(n12463) );
  NOR U13390 ( .A(n15320), .B(n15318), .Z(n15319) );
  XOR U13391 ( .A(n15321), .B(n15322), .Z(n12466) );
  NOR U13392 ( .A(n15323), .B(n15321), .Z(n15322) );
  XOR U13393 ( .A(n15324), .B(n15325), .Z(n12469) );
  NOR U13394 ( .A(n15326), .B(n15324), .Z(n15325) );
  XOR U13395 ( .A(n15327), .B(n15328), .Z(n12472) );
  NOR U13396 ( .A(n15329), .B(n15327), .Z(n15328) );
  XOR U13397 ( .A(n15330), .B(n15331), .Z(n12475) );
  NOR U13398 ( .A(n15332), .B(n15330), .Z(n15331) );
  XOR U13399 ( .A(n15333), .B(n15334), .Z(n12478) );
  NOR U13400 ( .A(n15335), .B(n15333), .Z(n15334) );
  XOR U13401 ( .A(n15336), .B(n15337), .Z(n12481) );
  NOR U13402 ( .A(n15338), .B(n15336), .Z(n15337) );
  XOR U13403 ( .A(n15339), .B(n15340), .Z(n12484) );
  NOR U13404 ( .A(n15341), .B(n15339), .Z(n15340) );
  XOR U13405 ( .A(n15342), .B(n15343), .Z(n12487) );
  NOR U13406 ( .A(n15344), .B(n15342), .Z(n15343) );
  XOR U13407 ( .A(n15345), .B(n15346), .Z(n12490) );
  NOR U13408 ( .A(n15347), .B(n15345), .Z(n15346) );
  XOR U13409 ( .A(n15348), .B(n15349), .Z(n12493) );
  NOR U13410 ( .A(n15350), .B(n15348), .Z(n15349) );
  XOR U13411 ( .A(n15351), .B(n15352), .Z(n12496) );
  NOR U13412 ( .A(n15353), .B(n15351), .Z(n15352) );
  XOR U13413 ( .A(n15354), .B(n15355), .Z(n12499) );
  NOR U13414 ( .A(n15356), .B(n15354), .Z(n15355) );
  XOR U13415 ( .A(n15357), .B(n15358), .Z(n12502) );
  NOR U13416 ( .A(n15359), .B(n15357), .Z(n15358) );
  XOR U13417 ( .A(n15360), .B(n15361), .Z(n12505) );
  NOR U13418 ( .A(n15362), .B(n15360), .Z(n15361) );
  XOR U13419 ( .A(n15363), .B(n15364), .Z(n12508) );
  NOR U13420 ( .A(n15365), .B(n15363), .Z(n15364) );
  XOR U13421 ( .A(n15366), .B(n15367), .Z(n12511) );
  NOR U13422 ( .A(n15368), .B(n15366), .Z(n15367) );
  XOR U13423 ( .A(n15369), .B(n15370), .Z(n12514) );
  NOR U13424 ( .A(n15371), .B(n15369), .Z(n15370) );
  XOR U13425 ( .A(n15372), .B(n15373), .Z(n12517) );
  NOR U13426 ( .A(n15374), .B(n15372), .Z(n15373) );
  XOR U13427 ( .A(n15375), .B(n15376), .Z(n12520) );
  NOR U13428 ( .A(n15377), .B(n15375), .Z(n15376) );
  XOR U13429 ( .A(n15378), .B(n15379), .Z(n12523) );
  NOR U13430 ( .A(n15380), .B(n15378), .Z(n15379) );
  XOR U13431 ( .A(n15381), .B(n15382), .Z(n12526) );
  NOR U13432 ( .A(n15383), .B(n15381), .Z(n15382) );
  XOR U13433 ( .A(n15384), .B(n15385), .Z(n12529) );
  NOR U13434 ( .A(n15386), .B(n15384), .Z(n15385) );
  XOR U13435 ( .A(n15387), .B(n15388), .Z(n12532) );
  NOR U13436 ( .A(n15389), .B(n15387), .Z(n15388) );
  XOR U13437 ( .A(n15390), .B(n15391), .Z(n12535) );
  NOR U13438 ( .A(n15392), .B(n15390), .Z(n15391) );
  XOR U13439 ( .A(n15393), .B(n15394), .Z(n12538) );
  NOR U13440 ( .A(n15395), .B(n15393), .Z(n15394) );
  XOR U13441 ( .A(n15396), .B(n15397), .Z(n12541) );
  NOR U13442 ( .A(n15398), .B(n15396), .Z(n15397) );
  XOR U13443 ( .A(n15399), .B(n15400), .Z(n12544) );
  NOR U13444 ( .A(n15401), .B(n15399), .Z(n15400) );
  XOR U13445 ( .A(n15402), .B(n15403), .Z(n12547) );
  NOR U13446 ( .A(n15404), .B(n15402), .Z(n15403) );
  XOR U13447 ( .A(n15405), .B(n15406), .Z(n12550) );
  NOR U13448 ( .A(n15407), .B(n15405), .Z(n15406) );
  XOR U13449 ( .A(n15408), .B(n15409), .Z(n12553) );
  NOR U13450 ( .A(n15410), .B(n15408), .Z(n15409) );
  XOR U13451 ( .A(n15411), .B(n15412), .Z(n12556) );
  NOR U13452 ( .A(n15413), .B(n15411), .Z(n15412) );
  XOR U13453 ( .A(n15414), .B(n15415), .Z(n12559) );
  NOR U13454 ( .A(n15416), .B(n15414), .Z(n15415) );
  XOR U13455 ( .A(n15417), .B(n15418), .Z(n12562) );
  NOR U13456 ( .A(n15419), .B(n15417), .Z(n15418) );
  XOR U13457 ( .A(n15420), .B(n15421), .Z(n12565) );
  NOR U13458 ( .A(n15422), .B(n15420), .Z(n15421) );
  XOR U13459 ( .A(n15423), .B(n15424), .Z(n12568) );
  NOR U13460 ( .A(n15425), .B(n15423), .Z(n15424) );
  XOR U13461 ( .A(n15426), .B(n15427), .Z(n12571) );
  NOR U13462 ( .A(n15428), .B(n15426), .Z(n15427) );
  XOR U13463 ( .A(n15429), .B(n15430), .Z(n12574) );
  NOR U13464 ( .A(n15431), .B(n15429), .Z(n15430) );
  XOR U13465 ( .A(n15432), .B(n15433), .Z(n12577) );
  NOR U13466 ( .A(n15434), .B(n15432), .Z(n15433) );
  XOR U13467 ( .A(n15435), .B(n15436), .Z(n12580) );
  NOR U13468 ( .A(n15437), .B(n15435), .Z(n15436) );
  XOR U13469 ( .A(n15438), .B(n15439), .Z(n12583) );
  NOR U13470 ( .A(n15440), .B(n15438), .Z(n15439) );
  XOR U13471 ( .A(n15441), .B(n15442), .Z(n12586) );
  NOR U13472 ( .A(n15443), .B(n15441), .Z(n15442) );
  XOR U13473 ( .A(n15444), .B(n15445), .Z(n12589) );
  NOR U13474 ( .A(n15446), .B(n15444), .Z(n15445) );
  XOR U13475 ( .A(n15447), .B(n15448), .Z(n12592) );
  NOR U13476 ( .A(n15449), .B(n15447), .Z(n15448) );
  XOR U13477 ( .A(n15450), .B(n15451), .Z(n12595) );
  NOR U13478 ( .A(n15452), .B(n15450), .Z(n15451) );
  XOR U13479 ( .A(n15453), .B(n15454), .Z(n12598) );
  NOR U13480 ( .A(n15455), .B(n15453), .Z(n15454) );
  XOR U13481 ( .A(n15456), .B(n15457), .Z(n12601) );
  NOR U13482 ( .A(n15458), .B(n15456), .Z(n15457) );
  XOR U13483 ( .A(n15459), .B(n15460), .Z(n12604) );
  NOR U13484 ( .A(n15461), .B(n15459), .Z(n15460) );
  XOR U13485 ( .A(n15462), .B(n15463), .Z(n12607) );
  NOR U13486 ( .A(n15464), .B(n15462), .Z(n15463) );
  XOR U13487 ( .A(n15465), .B(n15466), .Z(n12610) );
  NOR U13488 ( .A(n15467), .B(n15465), .Z(n15466) );
  XOR U13489 ( .A(n15468), .B(n15469), .Z(n12613) );
  NOR U13490 ( .A(n15470), .B(n15468), .Z(n15469) );
  XOR U13491 ( .A(n15471), .B(n15472), .Z(n12616) );
  NOR U13492 ( .A(n15473), .B(n15471), .Z(n15472) );
  XOR U13493 ( .A(n15474), .B(n15475), .Z(n12619) );
  NOR U13494 ( .A(n15476), .B(n15474), .Z(n15475) );
  XOR U13495 ( .A(n15477), .B(n15478), .Z(n12622) );
  NOR U13496 ( .A(n15479), .B(n15477), .Z(n15478) );
  XOR U13497 ( .A(n15480), .B(n15481), .Z(n12625) );
  NOR U13498 ( .A(n15482), .B(n15480), .Z(n15481) );
  XOR U13499 ( .A(n15483), .B(n15484), .Z(n12628) );
  NOR U13500 ( .A(n15485), .B(n15483), .Z(n15484) );
  XOR U13501 ( .A(n15486), .B(n15487), .Z(n12631) );
  NOR U13502 ( .A(n15488), .B(n15486), .Z(n15487) );
  XOR U13503 ( .A(n15489), .B(n15490), .Z(n12634) );
  NOR U13504 ( .A(n15491), .B(n15489), .Z(n15490) );
  XOR U13505 ( .A(n15492), .B(n15493), .Z(n12637) );
  NOR U13506 ( .A(n15494), .B(n15492), .Z(n15493) );
  XOR U13507 ( .A(n15495), .B(n15496), .Z(n12640) );
  NOR U13508 ( .A(n15497), .B(n15495), .Z(n15496) );
  XOR U13509 ( .A(n15498), .B(n15499), .Z(n12643) );
  NOR U13510 ( .A(n15500), .B(n15498), .Z(n15499) );
  XOR U13511 ( .A(n15501), .B(n15502), .Z(n12646) );
  NOR U13512 ( .A(n15503), .B(n15501), .Z(n15502) );
  XOR U13513 ( .A(n15504), .B(n15505), .Z(n12649) );
  NOR U13514 ( .A(n15506), .B(n15504), .Z(n15505) );
  XOR U13515 ( .A(n15507), .B(n15508), .Z(n12652) );
  NOR U13516 ( .A(n15509), .B(n15507), .Z(n15508) );
  XOR U13517 ( .A(n15510), .B(n15511), .Z(n12655) );
  NOR U13518 ( .A(n15512), .B(n15510), .Z(n15511) );
  XOR U13519 ( .A(n15513), .B(n15514), .Z(n12658) );
  NOR U13520 ( .A(n15515), .B(n15513), .Z(n15514) );
  XOR U13521 ( .A(n15516), .B(n15517), .Z(n12661) );
  NOR U13522 ( .A(n15518), .B(n15516), .Z(n15517) );
  XOR U13523 ( .A(n15519), .B(n15520), .Z(n12664) );
  NOR U13524 ( .A(n15521), .B(n15519), .Z(n15520) );
  XOR U13525 ( .A(n15522), .B(n15523), .Z(n12667) );
  NOR U13526 ( .A(n15524), .B(n15522), .Z(n15523) );
  XOR U13527 ( .A(n15525), .B(n15526), .Z(n12670) );
  NOR U13528 ( .A(n15527), .B(n15525), .Z(n15526) );
  XOR U13529 ( .A(n15528), .B(n15529), .Z(n12673) );
  NOR U13530 ( .A(n15530), .B(n15528), .Z(n15529) );
  XOR U13531 ( .A(n15531), .B(n15532), .Z(n12676) );
  NOR U13532 ( .A(n15533), .B(n15531), .Z(n15532) );
  XOR U13533 ( .A(n15534), .B(n15535), .Z(n12679) );
  NOR U13534 ( .A(n15536), .B(n15534), .Z(n15535) );
  XOR U13535 ( .A(n15537), .B(n15538), .Z(n12682) );
  NOR U13536 ( .A(n15539), .B(n15537), .Z(n15538) );
  XOR U13537 ( .A(n15540), .B(n15541), .Z(n12685) );
  NOR U13538 ( .A(n15542), .B(n15540), .Z(n15541) );
  XOR U13539 ( .A(n15543), .B(n15544), .Z(n12688) );
  NOR U13540 ( .A(n15545), .B(n15543), .Z(n15544) );
  XOR U13541 ( .A(n15546), .B(n15547), .Z(n12691) );
  NOR U13542 ( .A(n15548), .B(n15546), .Z(n15547) );
  XOR U13543 ( .A(n15549), .B(n15550), .Z(n12694) );
  NOR U13544 ( .A(n15551), .B(n15549), .Z(n15550) );
  XOR U13545 ( .A(n15552), .B(n15553), .Z(n12697) );
  NOR U13546 ( .A(n15554), .B(n15552), .Z(n15553) );
  XOR U13547 ( .A(n15555), .B(n15556), .Z(n12700) );
  NOR U13548 ( .A(n15557), .B(n15555), .Z(n15556) );
  XOR U13549 ( .A(n15558), .B(n15559), .Z(n12703) );
  NOR U13550 ( .A(n15560), .B(n15558), .Z(n15559) );
  XOR U13551 ( .A(n15561), .B(n15562), .Z(n12706) );
  NOR U13552 ( .A(n15563), .B(n15561), .Z(n15562) );
  XOR U13553 ( .A(n15564), .B(n15565), .Z(n12709) );
  NOR U13554 ( .A(n15566), .B(n15564), .Z(n15565) );
  XOR U13555 ( .A(n15567), .B(n15568), .Z(n12712) );
  NOR U13556 ( .A(n15569), .B(n15567), .Z(n15568) );
  XOR U13557 ( .A(n15570), .B(n15571), .Z(n12715) );
  NOR U13558 ( .A(n15572), .B(n15570), .Z(n15571) );
  XOR U13559 ( .A(n15573), .B(n15574), .Z(n12718) );
  NOR U13560 ( .A(n15575), .B(n15573), .Z(n15574) );
  XOR U13561 ( .A(n15576), .B(n15577), .Z(n12721) );
  NOR U13562 ( .A(n15578), .B(n15576), .Z(n15577) );
  XOR U13563 ( .A(n15579), .B(n15580), .Z(n12724) );
  NOR U13564 ( .A(n15581), .B(n15579), .Z(n15580) );
  XOR U13565 ( .A(n15582), .B(n15583), .Z(n12727) );
  NOR U13566 ( .A(n15584), .B(n15582), .Z(n15583) );
  XOR U13567 ( .A(n15585), .B(n15586), .Z(n12730) );
  NOR U13568 ( .A(n15587), .B(n15585), .Z(n15586) );
  XNOR U13569 ( .A(n15588), .B(n15589), .Z(n12733) );
  NOR U13570 ( .A(n15590), .B(n15588), .Z(n15589) );
  XOR U13571 ( .A(n15591), .B(n15592), .Z(n12736) );
  AND U13572 ( .A(n119), .B(n15591), .Z(n15592) );
  XNOR U13573 ( .A(n15593), .B(n14168), .Z(n14170) );
  IV U13574 ( .A(n102), .Z(n15593) );
  XOR U13575 ( .A(n14165), .B(n14164), .Z(n102) );
  XNOR U13576 ( .A(n14162), .B(n14161), .Z(n14164) );
  XNOR U13577 ( .A(n14159), .B(n14158), .Z(n14161) );
  XNOR U13578 ( .A(n14156), .B(n14155), .Z(n14158) );
  XNOR U13579 ( .A(n14153), .B(n14152), .Z(n14155) );
  XNOR U13580 ( .A(n14150), .B(n14149), .Z(n14152) );
  XNOR U13581 ( .A(n14147), .B(n14146), .Z(n14149) );
  XNOR U13582 ( .A(n14144), .B(n14143), .Z(n14146) );
  XNOR U13583 ( .A(n14141), .B(n14140), .Z(n14143) );
  XNOR U13584 ( .A(n14138), .B(n14137), .Z(n14140) );
  XNOR U13585 ( .A(n14135), .B(n14134), .Z(n14137) );
  XNOR U13586 ( .A(n14132), .B(n14131), .Z(n14134) );
  XNOR U13587 ( .A(n14129), .B(n14128), .Z(n14131) );
  XNOR U13588 ( .A(n14126), .B(n14125), .Z(n14128) );
  XNOR U13589 ( .A(n14123), .B(n14122), .Z(n14125) );
  XNOR U13590 ( .A(n14120), .B(n14119), .Z(n14122) );
  XNOR U13591 ( .A(n14117), .B(n14116), .Z(n14119) );
  XNOR U13592 ( .A(n14114), .B(n14113), .Z(n14116) );
  XNOR U13593 ( .A(n14111), .B(n14110), .Z(n14113) );
  XNOR U13594 ( .A(n14108), .B(n14107), .Z(n14110) );
  XNOR U13595 ( .A(n14105), .B(n14104), .Z(n14107) );
  XNOR U13596 ( .A(n14102), .B(n14101), .Z(n14104) );
  XNOR U13597 ( .A(n14099), .B(n14098), .Z(n14101) );
  XNOR U13598 ( .A(n14096), .B(n14095), .Z(n14098) );
  XNOR U13599 ( .A(n14093), .B(n14092), .Z(n14095) );
  XNOR U13600 ( .A(n14090), .B(n14089), .Z(n14092) );
  XNOR U13601 ( .A(n14087), .B(n14086), .Z(n14089) );
  XNOR U13602 ( .A(n14084), .B(n14083), .Z(n14086) );
  XNOR U13603 ( .A(n14081), .B(n14080), .Z(n14083) );
  XNOR U13604 ( .A(n14078), .B(n14077), .Z(n14080) );
  XNOR U13605 ( .A(n14075), .B(n14074), .Z(n14077) );
  XNOR U13606 ( .A(n14072), .B(n14071), .Z(n14074) );
  XNOR U13607 ( .A(n14069), .B(n14068), .Z(n14071) );
  XNOR U13608 ( .A(n14066), .B(n14065), .Z(n14068) );
  XNOR U13609 ( .A(n14063), .B(n14062), .Z(n14065) );
  XNOR U13610 ( .A(n14060), .B(n14059), .Z(n14062) );
  XNOR U13611 ( .A(n14057), .B(n14056), .Z(n14059) );
  XNOR U13612 ( .A(n14054), .B(n14053), .Z(n14056) );
  XNOR U13613 ( .A(n14051), .B(n14050), .Z(n14053) );
  XNOR U13614 ( .A(n14048), .B(n14047), .Z(n14050) );
  XNOR U13615 ( .A(n14045), .B(n14044), .Z(n14047) );
  XNOR U13616 ( .A(n14042), .B(n14041), .Z(n14044) );
  XNOR U13617 ( .A(n14039), .B(n14038), .Z(n14041) );
  XNOR U13618 ( .A(n14036), .B(n14035), .Z(n14038) );
  XNOR U13619 ( .A(n14033), .B(n14032), .Z(n14035) );
  XNOR U13620 ( .A(n14030), .B(n14029), .Z(n14032) );
  XNOR U13621 ( .A(n14027), .B(n14026), .Z(n14029) );
  XNOR U13622 ( .A(n14024), .B(n14023), .Z(n14026) );
  XNOR U13623 ( .A(n14021), .B(n14020), .Z(n14023) );
  XNOR U13624 ( .A(n14018), .B(n14017), .Z(n14020) );
  XNOR U13625 ( .A(n14015), .B(n14014), .Z(n14017) );
  XNOR U13626 ( .A(n14012), .B(n14011), .Z(n14014) );
  XNOR U13627 ( .A(n14009), .B(n14008), .Z(n14011) );
  XNOR U13628 ( .A(n14006), .B(n14005), .Z(n14008) );
  XNOR U13629 ( .A(n14003), .B(n14002), .Z(n14005) );
  XNOR U13630 ( .A(n14000), .B(n13999), .Z(n14002) );
  XNOR U13631 ( .A(n13997), .B(n13996), .Z(n13999) );
  XNOR U13632 ( .A(n13994), .B(n13993), .Z(n13996) );
  XNOR U13633 ( .A(n13991), .B(n13990), .Z(n13993) );
  XNOR U13634 ( .A(n13988), .B(n13987), .Z(n13990) );
  XNOR U13635 ( .A(n13985), .B(n13984), .Z(n13987) );
  XNOR U13636 ( .A(n13982), .B(n13981), .Z(n13984) );
  XNOR U13637 ( .A(n13979), .B(n13978), .Z(n13981) );
  XNOR U13638 ( .A(n13976), .B(n13975), .Z(n13978) );
  XNOR U13639 ( .A(n13973), .B(n13972), .Z(n13975) );
  XNOR U13640 ( .A(n13970), .B(n13969), .Z(n13972) );
  XNOR U13641 ( .A(n13967), .B(n13966), .Z(n13969) );
  XNOR U13642 ( .A(n13964), .B(n13963), .Z(n13966) );
  XNOR U13643 ( .A(n13961), .B(n13960), .Z(n13963) );
  XNOR U13644 ( .A(n13958), .B(n13957), .Z(n13960) );
  XNOR U13645 ( .A(n13955), .B(n13954), .Z(n13957) );
  XNOR U13646 ( .A(n13952), .B(n13951), .Z(n13954) );
  XNOR U13647 ( .A(n13949), .B(n13948), .Z(n13951) );
  XNOR U13648 ( .A(n13946), .B(n13945), .Z(n13948) );
  XNOR U13649 ( .A(n13943), .B(n13942), .Z(n13945) );
  XNOR U13650 ( .A(n13940), .B(n13939), .Z(n13942) );
  XNOR U13651 ( .A(n13937), .B(n13936), .Z(n13939) );
  XNOR U13652 ( .A(n13934), .B(n13933), .Z(n13936) );
  XNOR U13653 ( .A(n13931), .B(n13930), .Z(n13933) );
  XNOR U13654 ( .A(n13928), .B(n13927), .Z(n13930) );
  XNOR U13655 ( .A(n13925), .B(n13924), .Z(n13927) );
  XNOR U13656 ( .A(n13922), .B(n13921), .Z(n13924) );
  XNOR U13657 ( .A(n13919), .B(n13918), .Z(n13921) );
  XNOR U13658 ( .A(n13916), .B(n13915), .Z(n13918) );
  XNOR U13659 ( .A(n13913), .B(n13912), .Z(n13915) );
  XNOR U13660 ( .A(n13910), .B(n13909), .Z(n13912) );
  XNOR U13661 ( .A(n13907), .B(n13906), .Z(n13909) );
  XNOR U13662 ( .A(n13904), .B(n13903), .Z(n13906) );
  XNOR U13663 ( .A(n13901), .B(n13900), .Z(n13903) );
  XNOR U13664 ( .A(n13898), .B(n13897), .Z(n13900) );
  XNOR U13665 ( .A(n13895), .B(n13894), .Z(n13897) );
  XNOR U13666 ( .A(n13892), .B(n13891), .Z(n13894) );
  XNOR U13667 ( .A(n13889), .B(n13888), .Z(n13891) );
  XNOR U13668 ( .A(n13886), .B(n13885), .Z(n13888) );
  XNOR U13669 ( .A(n13883), .B(n13882), .Z(n13885) );
  XNOR U13670 ( .A(n13880), .B(n13879), .Z(n13882) );
  XNOR U13671 ( .A(n13877), .B(n13876), .Z(n13879) );
  XNOR U13672 ( .A(n13874), .B(n13873), .Z(n13876) );
  XNOR U13673 ( .A(n13871), .B(n13870), .Z(n13873) );
  XNOR U13674 ( .A(n13868), .B(n13867), .Z(n13870) );
  XNOR U13675 ( .A(n13865), .B(n13864), .Z(n13867) );
  XNOR U13676 ( .A(n13862), .B(n13861), .Z(n13864) );
  XNOR U13677 ( .A(n13859), .B(n13858), .Z(n13861) );
  XNOR U13678 ( .A(n13856), .B(n13855), .Z(n13858) );
  XNOR U13679 ( .A(n13853), .B(n13852), .Z(n13855) );
  XNOR U13680 ( .A(n13850), .B(n13849), .Z(n13852) );
  XNOR U13681 ( .A(n13847), .B(n13846), .Z(n13849) );
  XNOR U13682 ( .A(n13844), .B(n13843), .Z(n13846) );
  XNOR U13683 ( .A(n13841), .B(n13840), .Z(n13843) );
  XNOR U13684 ( .A(n13838), .B(n13837), .Z(n13840) );
  XNOR U13685 ( .A(n13835), .B(n13834), .Z(n13837) );
  XNOR U13686 ( .A(n13832), .B(n13831), .Z(n13834) );
  XNOR U13687 ( .A(n13829), .B(n13828), .Z(n13831) );
  XNOR U13688 ( .A(n13826), .B(n13825), .Z(n13828) );
  XNOR U13689 ( .A(n13823), .B(n13822), .Z(n13825) );
  XNOR U13690 ( .A(n13820), .B(n13819), .Z(n13822) );
  XNOR U13691 ( .A(n13817), .B(n13816), .Z(n13819) );
  XNOR U13692 ( .A(n13814), .B(n13813), .Z(n13816) );
  XNOR U13693 ( .A(n13811), .B(n13810), .Z(n13813) );
  XNOR U13694 ( .A(n13808), .B(n13807), .Z(n13810) );
  XNOR U13695 ( .A(n13805), .B(n13804), .Z(n13807) );
  XNOR U13696 ( .A(n13802), .B(n13801), .Z(n13804) );
  XNOR U13697 ( .A(n13799), .B(n13798), .Z(n13801) );
  XNOR U13698 ( .A(n13796), .B(n13795), .Z(n13798) );
  XNOR U13699 ( .A(n13793), .B(n13792), .Z(n13795) );
  XNOR U13700 ( .A(n13790), .B(n13789), .Z(n13792) );
  XNOR U13701 ( .A(n13787), .B(n13786), .Z(n13789) );
  XNOR U13702 ( .A(n13784), .B(n13783), .Z(n13786) );
  XNOR U13703 ( .A(n13781), .B(n13780), .Z(n13783) );
  XNOR U13704 ( .A(n13778), .B(n13777), .Z(n13780) );
  XNOR U13705 ( .A(n13775), .B(n13774), .Z(n13777) );
  XNOR U13706 ( .A(n13772), .B(n13771), .Z(n13774) );
  XNOR U13707 ( .A(n13769), .B(n13768), .Z(n13771) );
  XNOR U13708 ( .A(n13766), .B(n13765), .Z(n13768) );
  XNOR U13709 ( .A(n13763), .B(n13762), .Z(n13765) );
  XNOR U13710 ( .A(n13760), .B(n13759), .Z(n13762) );
  XNOR U13711 ( .A(n13757), .B(n13756), .Z(n13759) );
  XNOR U13712 ( .A(n13754), .B(n13753), .Z(n13756) );
  XNOR U13713 ( .A(n13751), .B(n13750), .Z(n13753) );
  XNOR U13714 ( .A(n13748), .B(n13747), .Z(n13750) );
  XNOR U13715 ( .A(n13745), .B(n13744), .Z(n13747) );
  XNOR U13716 ( .A(n13742), .B(n13741), .Z(n13744) );
  XNOR U13717 ( .A(n13739), .B(n13738), .Z(n13741) );
  XNOR U13718 ( .A(n13736), .B(n13735), .Z(n13738) );
  XNOR U13719 ( .A(n13733), .B(n13732), .Z(n13735) );
  XNOR U13720 ( .A(n13730), .B(n13729), .Z(n13732) );
  XNOR U13721 ( .A(n13727), .B(n13726), .Z(n13729) );
  XNOR U13722 ( .A(n13724), .B(n13723), .Z(n13726) );
  XNOR U13723 ( .A(n13721), .B(n13720), .Z(n13723) );
  XNOR U13724 ( .A(n13718), .B(n13717), .Z(n13720) );
  XNOR U13725 ( .A(n13715), .B(n13714), .Z(n13717) );
  XNOR U13726 ( .A(n13712), .B(n13711), .Z(n13714) );
  XNOR U13727 ( .A(n13709), .B(n13708), .Z(n13711) );
  XNOR U13728 ( .A(n13706), .B(n13705), .Z(n13708) );
  XNOR U13729 ( .A(n13703), .B(n13702), .Z(n13705) );
  XNOR U13730 ( .A(n13700), .B(n13699), .Z(n13702) );
  XNOR U13731 ( .A(n13697), .B(n13696), .Z(n13699) );
  XNOR U13732 ( .A(n13694), .B(n13693), .Z(n13696) );
  XNOR U13733 ( .A(n13691), .B(n13690), .Z(n13693) );
  XNOR U13734 ( .A(n13688), .B(n13687), .Z(n13690) );
  XNOR U13735 ( .A(n13685), .B(n13684), .Z(n13687) );
  XNOR U13736 ( .A(n13682), .B(n13681), .Z(n13684) );
  XNOR U13737 ( .A(n13679), .B(n13678), .Z(n13681) );
  XNOR U13738 ( .A(n13676), .B(n13675), .Z(n13678) );
  XNOR U13739 ( .A(n13673), .B(n13672), .Z(n13675) );
  XNOR U13740 ( .A(n13670), .B(n13669), .Z(n13672) );
  XNOR U13741 ( .A(n13667), .B(n13666), .Z(n13669) );
  XNOR U13742 ( .A(n13664), .B(n13663), .Z(n13666) );
  XNOR U13743 ( .A(n13661), .B(n13660), .Z(n13663) );
  XNOR U13744 ( .A(n13658), .B(n13657), .Z(n13660) );
  XNOR U13745 ( .A(n13655), .B(n13654), .Z(n13657) );
  XNOR U13746 ( .A(n13652), .B(n13651), .Z(n13654) );
  XNOR U13747 ( .A(n13649), .B(n13648), .Z(n13651) );
  XNOR U13748 ( .A(n13646), .B(n13645), .Z(n13648) );
  XNOR U13749 ( .A(n13643), .B(n13642), .Z(n13645) );
  XNOR U13750 ( .A(n13640), .B(n13639), .Z(n13642) );
  XNOR U13751 ( .A(n13637), .B(n13636), .Z(n13639) );
  XNOR U13752 ( .A(n13634), .B(n13633), .Z(n13636) );
  XNOR U13753 ( .A(n13631), .B(n13630), .Z(n13633) );
  XNOR U13754 ( .A(n13628), .B(n13627), .Z(n13630) );
  XNOR U13755 ( .A(n13625), .B(n13624), .Z(n13627) );
  XNOR U13756 ( .A(n13622), .B(n13621), .Z(n13624) );
  XNOR U13757 ( .A(n13619), .B(n13618), .Z(n13621) );
  XNOR U13758 ( .A(n13616), .B(n13615), .Z(n13618) );
  XNOR U13759 ( .A(n13613), .B(n13612), .Z(n13615) );
  XNOR U13760 ( .A(n13610), .B(n13609), .Z(n13612) );
  XNOR U13761 ( .A(n13607), .B(n13606), .Z(n13609) );
  XNOR U13762 ( .A(n13604), .B(n13603), .Z(n13606) );
  XNOR U13763 ( .A(n13601), .B(n13600), .Z(n13603) );
  XNOR U13764 ( .A(n13598), .B(n13597), .Z(n13600) );
  XNOR U13765 ( .A(n13595), .B(n13594), .Z(n13597) );
  XNOR U13766 ( .A(n13592), .B(n13591), .Z(n13594) );
  XNOR U13767 ( .A(n13589), .B(n13588), .Z(n13591) );
  XNOR U13768 ( .A(n13586), .B(n13585), .Z(n13588) );
  XNOR U13769 ( .A(n13583), .B(n13582), .Z(n13585) );
  XNOR U13770 ( .A(n13580), .B(n13579), .Z(n13582) );
  XNOR U13771 ( .A(n13577), .B(n13576), .Z(n13579) );
  XNOR U13772 ( .A(n13574), .B(n13573), .Z(n13576) );
  XNOR U13773 ( .A(n13571), .B(n13570), .Z(n13573) );
  XNOR U13774 ( .A(n13568), .B(n13567), .Z(n13570) );
  XNOR U13775 ( .A(n13565), .B(n13564), .Z(n13567) );
  XNOR U13776 ( .A(n13562), .B(n13561), .Z(n13564) );
  XNOR U13777 ( .A(n13559), .B(n13558), .Z(n13561) );
  XNOR U13778 ( .A(n13556), .B(n13555), .Z(n13558) );
  XNOR U13779 ( .A(n13553), .B(n13552), .Z(n13555) );
  XNOR U13780 ( .A(n13550), .B(n13549), .Z(n13552) );
  XNOR U13781 ( .A(n13547), .B(n13546), .Z(n13549) );
  XNOR U13782 ( .A(n13544), .B(n13543), .Z(n13546) );
  XNOR U13783 ( .A(n13541), .B(n13540), .Z(n13543) );
  XNOR U13784 ( .A(n13538), .B(n13537), .Z(n13540) );
  XNOR U13785 ( .A(n13535), .B(n13534), .Z(n13537) );
  XNOR U13786 ( .A(n13532), .B(n13531), .Z(n13534) );
  XNOR U13787 ( .A(n13529), .B(n13528), .Z(n13531) );
  XNOR U13788 ( .A(n13526), .B(n13525), .Z(n13528) );
  XNOR U13789 ( .A(n13523), .B(n13522), .Z(n13525) );
  XNOR U13790 ( .A(n13520), .B(n13519), .Z(n13522) );
  XNOR U13791 ( .A(n13517), .B(n13516), .Z(n13519) );
  XNOR U13792 ( .A(n13514), .B(n13513), .Z(n13516) );
  XNOR U13793 ( .A(n13511), .B(n13510), .Z(n13513) );
  XNOR U13794 ( .A(n13508), .B(n13507), .Z(n13510) );
  XNOR U13795 ( .A(n13505), .B(n13504), .Z(n13507) );
  XNOR U13796 ( .A(n13502), .B(n13501), .Z(n13504) );
  XNOR U13797 ( .A(n13499), .B(n13498), .Z(n13501) );
  XNOR U13798 ( .A(n13496), .B(n13495), .Z(n13498) );
  XNOR U13799 ( .A(n13493), .B(n13492), .Z(n13495) );
  XNOR U13800 ( .A(n13490), .B(n13489), .Z(n13492) );
  XNOR U13801 ( .A(n13487), .B(n13486), .Z(n13489) );
  XNOR U13802 ( .A(n13484), .B(n13483), .Z(n13486) );
  XNOR U13803 ( .A(n13481), .B(n13480), .Z(n13483) );
  XNOR U13804 ( .A(n13478), .B(n13477), .Z(n13480) );
  XNOR U13805 ( .A(n13475), .B(n13474), .Z(n13477) );
  XNOR U13806 ( .A(n13472), .B(n13471), .Z(n13474) );
  XNOR U13807 ( .A(n13469), .B(n13468), .Z(n13471) );
  XNOR U13808 ( .A(n13466), .B(n13465), .Z(n13468) );
  XNOR U13809 ( .A(n13463), .B(n13462), .Z(n13465) );
  XNOR U13810 ( .A(n13460), .B(n13459), .Z(n13462) );
  XNOR U13811 ( .A(n13457), .B(n13456), .Z(n13459) );
  XNOR U13812 ( .A(n13454), .B(n13453), .Z(n13456) );
  XNOR U13813 ( .A(n13451), .B(n13450), .Z(n13453) );
  XNOR U13814 ( .A(n13448), .B(n13447), .Z(n13450) );
  XNOR U13815 ( .A(n13445), .B(n13444), .Z(n13447) );
  XNOR U13816 ( .A(n13442), .B(n13441), .Z(n13444) );
  XNOR U13817 ( .A(n13439), .B(n13438), .Z(n13441) );
  XNOR U13818 ( .A(n13436), .B(n13435), .Z(n13438) );
  XNOR U13819 ( .A(n13433), .B(n13432), .Z(n13435) );
  XNOR U13820 ( .A(n13430), .B(n13429), .Z(n13432) );
  XNOR U13821 ( .A(n13427), .B(n13426), .Z(n13429) );
  XNOR U13822 ( .A(n13424), .B(n13423), .Z(n13426) );
  XNOR U13823 ( .A(n13421), .B(n13420), .Z(n13423) );
  XNOR U13824 ( .A(n13418), .B(n13417), .Z(n13420) );
  XNOR U13825 ( .A(n13415), .B(n13414), .Z(n13417) );
  XNOR U13826 ( .A(n13412), .B(n13411), .Z(n13414) );
  XNOR U13827 ( .A(n13409), .B(n13408), .Z(n13411) );
  XNOR U13828 ( .A(n13406), .B(n13405), .Z(n13408) );
  XNOR U13829 ( .A(n13403), .B(n13402), .Z(n13405) );
  XNOR U13830 ( .A(n13400), .B(n13399), .Z(n13402) );
  XNOR U13831 ( .A(n13397), .B(n13396), .Z(n13399) );
  XNOR U13832 ( .A(n13394), .B(n13393), .Z(n13396) );
  XNOR U13833 ( .A(n13391), .B(n13390), .Z(n13393) );
  XNOR U13834 ( .A(n13388), .B(n13387), .Z(n13390) );
  XNOR U13835 ( .A(n13385), .B(n13384), .Z(n13387) );
  XNOR U13836 ( .A(n13382), .B(n13381), .Z(n13384) );
  XNOR U13837 ( .A(n13379), .B(n13378), .Z(n13381) );
  XNOR U13838 ( .A(n13376), .B(n13375), .Z(n13378) );
  XNOR U13839 ( .A(n13373), .B(n13372), .Z(n13375) );
  XNOR U13840 ( .A(n13370), .B(n13369), .Z(n13372) );
  XNOR U13841 ( .A(n13367), .B(n13366), .Z(n13369) );
  XNOR U13842 ( .A(n13364), .B(n13363), .Z(n13366) );
  XNOR U13843 ( .A(n13361), .B(n13360), .Z(n13363) );
  XNOR U13844 ( .A(n13358), .B(n13357), .Z(n13360) );
  XNOR U13845 ( .A(n13355), .B(n13354), .Z(n13357) );
  XNOR U13846 ( .A(n13352), .B(n13351), .Z(n13354) );
  XNOR U13847 ( .A(n13349), .B(n13348), .Z(n13351) );
  XNOR U13848 ( .A(n13346), .B(n13345), .Z(n13348) );
  XNOR U13849 ( .A(n13343), .B(n13342), .Z(n13345) );
  XNOR U13850 ( .A(n13340), .B(n13339), .Z(n13342) );
  XNOR U13851 ( .A(n13337), .B(n13336), .Z(n13339) );
  XNOR U13852 ( .A(n13334), .B(n13333), .Z(n13336) );
  XNOR U13853 ( .A(n13331), .B(n13330), .Z(n13333) );
  XNOR U13854 ( .A(n13328), .B(n13327), .Z(n13330) );
  XNOR U13855 ( .A(n13325), .B(n13324), .Z(n13327) );
  XNOR U13856 ( .A(n13322), .B(n13321), .Z(n13324) );
  XNOR U13857 ( .A(n13319), .B(n13318), .Z(n13321) );
  XNOR U13858 ( .A(n13316), .B(n13315), .Z(n13318) );
  XNOR U13859 ( .A(n13313), .B(n13312), .Z(n13315) );
  XNOR U13860 ( .A(n13310), .B(n13309), .Z(n13312) );
  XNOR U13861 ( .A(n13307), .B(n13306), .Z(n13309) );
  XNOR U13862 ( .A(n13304), .B(n13303), .Z(n13306) );
  XNOR U13863 ( .A(n13301), .B(n13300), .Z(n13303) );
  XNOR U13864 ( .A(n13298), .B(n13297), .Z(n13300) );
  XNOR U13865 ( .A(n13295), .B(n13294), .Z(n13297) );
  XNOR U13866 ( .A(n13292), .B(n13291), .Z(n13294) );
  XNOR U13867 ( .A(n13289), .B(n13288), .Z(n13291) );
  XNOR U13868 ( .A(n13286), .B(n13285), .Z(n13288) );
  XNOR U13869 ( .A(n13283), .B(n13282), .Z(n13285) );
  XNOR U13870 ( .A(n13280), .B(n13279), .Z(n13282) );
  XNOR U13871 ( .A(n13277), .B(n13276), .Z(n13279) );
  XNOR U13872 ( .A(n13274), .B(n13273), .Z(n13276) );
  XNOR U13873 ( .A(n13271), .B(n13270), .Z(n13273) );
  XNOR U13874 ( .A(n13268), .B(n13267), .Z(n13270) );
  XNOR U13875 ( .A(n13265), .B(n13264), .Z(n13267) );
  XNOR U13876 ( .A(n13262), .B(n13261), .Z(n13264) );
  XNOR U13877 ( .A(n13259), .B(n13258), .Z(n13261) );
  XNOR U13878 ( .A(n13256), .B(n13255), .Z(n13258) );
  XNOR U13879 ( .A(n13253), .B(n13252), .Z(n13255) );
  XNOR U13880 ( .A(n13250), .B(n13249), .Z(n13252) );
  XNOR U13881 ( .A(n13247), .B(n13246), .Z(n13249) );
  XNOR U13882 ( .A(n13244), .B(n13243), .Z(n13246) );
  XNOR U13883 ( .A(n13241), .B(n13240), .Z(n13243) );
  XNOR U13884 ( .A(n13238), .B(n13237), .Z(n13240) );
  XNOR U13885 ( .A(n13235), .B(n13234), .Z(n13237) );
  XNOR U13886 ( .A(n13232), .B(n13231), .Z(n13234) );
  XNOR U13887 ( .A(n13229), .B(n13228), .Z(n13231) );
  XNOR U13888 ( .A(n13226), .B(n13225), .Z(n13228) );
  XNOR U13889 ( .A(n13223), .B(n13222), .Z(n13225) );
  XNOR U13890 ( .A(n13220), .B(n13219), .Z(n13222) );
  XNOR U13891 ( .A(n13217), .B(n13216), .Z(n13219) );
  XNOR U13892 ( .A(n13214), .B(n13213), .Z(n13216) );
  XNOR U13893 ( .A(n13211), .B(n13210), .Z(n13213) );
  XNOR U13894 ( .A(n13208), .B(n13207), .Z(n13210) );
  XNOR U13895 ( .A(n13205), .B(n13204), .Z(n13207) );
  XNOR U13896 ( .A(n13202), .B(n13201), .Z(n13204) );
  XNOR U13897 ( .A(n13199), .B(n13198), .Z(n13201) );
  XNOR U13898 ( .A(n13196), .B(n13195), .Z(n13198) );
  XNOR U13899 ( .A(n13193), .B(n13192), .Z(n13195) );
  XNOR U13900 ( .A(n13190), .B(n13189), .Z(n13192) );
  XNOR U13901 ( .A(n13187), .B(n13186), .Z(n13189) );
  XNOR U13902 ( .A(n13184), .B(n13183), .Z(n13186) );
  XNOR U13903 ( .A(n13181), .B(n13180), .Z(n13183) );
  XNOR U13904 ( .A(n13178), .B(n13177), .Z(n13180) );
  XNOR U13905 ( .A(n13175), .B(n13174), .Z(n13177) );
  XNOR U13906 ( .A(n13172), .B(n13171), .Z(n13174) );
  XNOR U13907 ( .A(n13169), .B(n13168), .Z(n13171) );
  XNOR U13908 ( .A(n13166), .B(n13165), .Z(n13168) );
  XNOR U13909 ( .A(n13163), .B(n13162), .Z(n13165) );
  XNOR U13910 ( .A(n13160), .B(n13159), .Z(n13162) );
  XNOR U13911 ( .A(n13157), .B(n13156), .Z(n13159) );
  XNOR U13912 ( .A(n13154), .B(n13153), .Z(n13156) );
  XNOR U13913 ( .A(n13151), .B(n13150), .Z(n13153) );
  XNOR U13914 ( .A(n13148), .B(n13147), .Z(n13150) );
  XNOR U13915 ( .A(n13145), .B(n13144), .Z(n13147) );
  XNOR U13916 ( .A(n13142), .B(n13141), .Z(n13144) );
  XNOR U13917 ( .A(n13139), .B(n13138), .Z(n13141) );
  XNOR U13918 ( .A(n13136), .B(n13135), .Z(n13138) );
  XNOR U13919 ( .A(n13133), .B(n13132), .Z(n13135) );
  XNOR U13920 ( .A(n13130), .B(n13129), .Z(n13132) );
  XNOR U13921 ( .A(n13127), .B(n13126), .Z(n13129) );
  XNOR U13922 ( .A(n13124), .B(n13123), .Z(n13126) );
  XNOR U13923 ( .A(n13121), .B(n13120), .Z(n13123) );
  XNOR U13924 ( .A(n13118), .B(n13117), .Z(n13120) );
  XNOR U13925 ( .A(n13115), .B(n13114), .Z(n13117) );
  XNOR U13926 ( .A(n13112), .B(n13111), .Z(n13114) );
  XNOR U13927 ( .A(n13109), .B(n13108), .Z(n13111) );
  XNOR U13928 ( .A(n13106), .B(n13105), .Z(n13108) );
  XNOR U13929 ( .A(n13103), .B(n13102), .Z(n13105) );
  XNOR U13930 ( .A(n13100), .B(n13099), .Z(n13102) );
  XNOR U13931 ( .A(n13097), .B(n13096), .Z(n13099) );
  XNOR U13932 ( .A(n13094), .B(n13093), .Z(n13096) );
  XNOR U13933 ( .A(n13091), .B(n13090), .Z(n13093) );
  XNOR U13934 ( .A(n13088), .B(n13087), .Z(n13090) );
  XNOR U13935 ( .A(n13085), .B(n13084), .Z(n13087) );
  XNOR U13936 ( .A(n13082), .B(n13081), .Z(n13084) );
  XNOR U13937 ( .A(n13079), .B(n13078), .Z(n13081) );
  XNOR U13938 ( .A(n13076), .B(n13075), .Z(n13078) );
  XNOR U13939 ( .A(n13073), .B(n13072), .Z(n13075) );
  XNOR U13940 ( .A(n13070), .B(n13069), .Z(n13072) );
  XNOR U13941 ( .A(n13067), .B(n13066), .Z(n13069) );
  XNOR U13942 ( .A(n13064), .B(n13063), .Z(n13066) );
  XNOR U13943 ( .A(n13061), .B(n13060), .Z(n13063) );
  XNOR U13944 ( .A(n13058), .B(n13057), .Z(n13060) );
  XNOR U13945 ( .A(n13055), .B(n13054), .Z(n13057) );
  XNOR U13946 ( .A(n13052), .B(n13051), .Z(n13054) );
  XNOR U13947 ( .A(n13049), .B(n13048), .Z(n13051) );
  XNOR U13948 ( .A(n13046), .B(n13045), .Z(n13048) );
  XNOR U13949 ( .A(n13043), .B(n13042), .Z(n13045) );
  XNOR U13950 ( .A(n13040), .B(n13039), .Z(n13042) );
  XNOR U13951 ( .A(n13037), .B(n13036), .Z(n13039) );
  XNOR U13952 ( .A(n13034), .B(n13033), .Z(n13036) );
  XNOR U13953 ( .A(n13031), .B(n13030), .Z(n13033) );
  XNOR U13954 ( .A(n13028), .B(n13027), .Z(n13030) );
  XNOR U13955 ( .A(n13025), .B(n13024), .Z(n13027) );
  XNOR U13956 ( .A(n13022), .B(n13021), .Z(n13024) );
  XNOR U13957 ( .A(n13019), .B(n13018), .Z(n13021) );
  XNOR U13958 ( .A(n13016), .B(n13015), .Z(n13018) );
  XNOR U13959 ( .A(n13013), .B(n13012), .Z(n13015) );
  XNOR U13960 ( .A(n13010), .B(n13009), .Z(n13012) );
  XNOR U13961 ( .A(n13007), .B(n13006), .Z(n13009) );
  XNOR U13962 ( .A(n13004), .B(n13003), .Z(n13006) );
  XNOR U13963 ( .A(n13001), .B(n13000), .Z(n13003) );
  XOR U13964 ( .A(n12998), .B(n12997), .Z(n13000) );
  XOR U13965 ( .A(n12995), .B(n12994), .Z(n12997) );
  XOR U13966 ( .A(n12991), .B(n12992), .Z(n12994) );
  AND U13967 ( .A(n15594), .B(n15595), .Z(n12992) );
  XOR U13968 ( .A(n12988), .B(n12989), .Z(n12991) );
  AND U13969 ( .A(n15596), .B(n15597), .Z(n12989) );
  XOR U13970 ( .A(n12985), .B(n12986), .Z(n12988) );
  AND U13971 ( .A(n15598), .B(n15599), .Z(n12986) );
  XNOR U13972 ( .A(n12740), .B(n12983), .Z(n12985) );
  AND U13973 ( .A(n15600), .B(n15601), .Z(n12983) );
  XOR U13974 ( .A(n12742), .B(n12741), .Z(n12740) );
  AND U13975 ( .A(n15602), .B(n15603), .Z(n12741) );
  XOR U13976 ( .A(n12744), .B(n12743), .Z(n12742) );
  AND U13977 ( .A(n15604), .B(n15605), .Z(n12743) );
  XOR U13978 ( .A(n12746), .B(n12745), .Z(n12744) );
  AND U13979 ( .A(n15606), .B(n15607), .Z(n12745) );
  XOR U13980 ( .A(n12748), .B(n12747), .Z(n12746) );
  AND U13981 ( .A(n15608), .B(n15609), .Z(n12747) );
  XOR U13982 ( .A(n12750), .B(n12749), .Z(n12748) );
  AND U13983 ( .A(n15610), .B(n15611), .Z(n12749) );
  XOR U13984 ( .A(n12752), .B(n12751), .Z(n12750) );
  AND U13985 ( .A(n15612), .B(n15613), .Z(n12751) );
  XOR U13986 ( .A(n12754), .B(n12753), .Z(n12752) );
  AND U13987 ( .A(n15614), .B(n15615), .Z(n12753) );
  XOR U13988 ( .A(n12756), .B(n12755), .Z(n12754) );
  AND U13989 ( .A(n15616), .B(n15617), .Z(n12755) );
  XOR U13990 ( .A(n12758), .B(n12757), .Z(n12756) );
  AND U13991 ( .A(n15618), .B(n15619), .Z(n12757) );
  XOR U13992 ( .A(n12760), .B(n12759), .Z(n12758) );
  AND U13993 ( .A(n15620), .B(n15621), .Z(n12759) );
  XOR U13994 ( .A(n12762), .B(n12761), .Z(n12760) );
  AND U13995 ( .A(n15622), .B(n15623), .Z(n12761) );
  XOR U13996 ( .A(n12764), .B(n12763), .Z(n12762) );
  AND U13997 ( .A(n15624), .B(n15625), .Z(n12763) );
  XOR U13998 ( .A(n12766), .B(n12765), .Z(n12764) );
  AND U13999 ( .A(n15626), .B(n15627), .Z(n12765) );
  XOR U14000 ( .A(n12768), .B(n12767), .Z(n12766) );
  AND U14001 ( .A(n15628), .B(n15629), .Z(n12767) );
  XOR U14002 ( .A(n12770), .B(n12769), .Z(n12768) );
  AND U14003 ( .A(n15630), .B(n15631), .Z(n12769) );
  XOR U14004 ( .A(n12772), .B(n12771), .Z(n12770) );
  AND U14005 ( .A(n15632), .B(n15633), .Z(n12771) );
  XOR U14006 ( .A(n12774), .B(n12773), .Z(n12772) );
  AND U14007 ( .A(n15634), .B(n15635), .Z(n12773) );
  XOR U14008 ( .A(n12776), .B(n12775), .Z(n12774) );
  AND U14009 ( .A(n15636), .B(n15637), .Z(n12775) );
  XOR U14010 ( .A(n12778), .B(n12777), .Z(n12776) );
  AND U14011 ( .A(n15638), .B(n15639), .Z(n12777) );
  XOR U14012 ( .A(n12780), .B(n12779), .Z(n12778) );
  AND U14013 ( .A(n15640), .B(n15641), .Z(n12779) );
  XOR U14014 ( .A(n12782), .B(n12781), .Z(n12780) );
  AND U14015 ( .A(n15642), .B(n15643), .Z(n12781) );
  XOR U14016 ( .A(n12784), .B(n12783), .Z(n12782) );
  AND U14017 ( .A(n15644), .B(n15645), .Z(n12783) );
  XOR U14018 ( .A(n12786), .B(n12785), .Z(n12784) );
  AND U14019 ( .A(n15646), .B(n15647), .Z(n12785) );
  XOR U14020 ( .A(n12788), .B(n12787), .Z(n12786) );
  AND U14021 ( .A(n15648), .B(n15649), .Z(n12787) );
  XOR U14022 ( .A(n12790), .B(n12789), .Z(n12788) );
  AND U14023 ( .A(n15650), .B(n15651), .Z(n12789) );
  XOR U14024 ( .A(n12792), .B(n12791), .Z(n12790) );
  AND U14025 ( .A(n15652), .B(n15653), .Z(n12791) );
  XOR U14026 ( .A(n12794), .B(n12793), .Z(n12792) );
  AND U14027 ( .A(n15654), .B(n15655), .Z(n12793) );
  XOR U14028 ( .A(n12796), .B(n12795), .Z(n12794) );
  AND U14029 ( .A(n15656), .B(n15657), .Z(n12795) );
  XOR U14030 ( .A(n12798), .B(n12797), .Z(n12796) );
  AND U14031 ( .A(n15658), .B(n15659), .Z(n12797) );
  XOR U14032 ( .A(n12800), .B(n12799), .Z(n12798) );
  AND U14033 ( .A(n15660), .B(n15661), .Z(n12799) );
  XOR U14034 ( .A(n12802), .B(n12801), .Z(n12800) );
  AND U14035 ( .A(n15662), .B(n15663), .Z(n12801) );
  XOR U14036 ( .A(n12804), .B(n12803), .Z(n12802) );
  AND U14037 ( .A(n15664), .B(n15665), .Z(n12803) );
  XOR U14038 ( .A(n12806), .B(n12805), .Z(n12804) );
  AND U14039 ( .A(n15666), .B(n15667), .Z(n12805) );
  XOR U14040 ( .A(n12808), .B(n12807), .Z(n12806) );
  AND U14041 ( .A(n15668), .B(n15669), .Z(n12807) );
  XOR U14042 ( .A(n12810), .B(n12809), .Z(n12808) );
  AND U14043 ( .A(n15670), .B(n15671), .Z(n12809) );
  XOR U14044 ( .A(n12812), .B(n12811), .Z(n12810) );
  AND U14045 ( .A(n15672), .B(n15673), .Z(n12811) );
  XOR U14046 ( .A(n12814), .B(n12813), .Z(n12812) );
  AND U14047 ( .A(n15674), .B(n15675), .Z(n12813) );
  XOR U14048 ( .A(n12816), .B(n12815), .Z(n12814) );
  AND U14049 ( .A(n15676), .B(n15677), .Z(n12815) );
  XOR U14050 ( .A(n12818), .B(n12817), .Z(n12816) );
  AND U14051 ( .A(n15678), .B(n15679), .Z(n12817) );
  XOR U14052 ( .A(n12820), .B(n12819), .Z(n12818) );
  AND U14053 ( .A(n15680), .B(n15681), .Z(n12819) );
  XOR U14054 ( .A(n12822), .B(n12821), .Z(n12820) );
  AND U14055 ( .A(n15682), .B(n15683), .Z(n12821) );
  XOR U14056 ( .A(n12824), .B(n12823), .Z(n12822) );
  AND U14057 ( .A(n15684), .B(n15685), .Z(n12823) );
  XOR U14058 ( .A(n12826), .B(n12825), .Z(n12824) );
  AND U14059 ( .A(n15686), .B(n15687), .Z(n12825) );
  XOR U14060 ( .A(n12828), .B(n12827), .Z(n12826) );
  AND U14061 ( .A(n15688), .B(n15689), .Z(n12827) );
  XOR U14062 ( .A(n12830), .B(n12829), .Z(n12828) );
  AND U14063 ( .A(n15690), .B(n15691), .Z(n12829) );
  XOR U14064 ( .A(n12832), .B(n12831), .Z(n12830) );
  AND U14065 ( .A(n15692), .B(n15693), .Z(n12831) );
  XOR U14066 ( .A(n12834), .B(n12833), .Z(n12832) );
  AND U14067 ( .A(n15694), .B(n15695), .Z(n12833) );
  XOR U14068 ( .A(n12836), .B(n12835), .Z(n12834) );
  AND U14069 ( .A(n15696), .B(n15697), .Z(n12835) );
  XOR U14070 ( .A(n12838), .B(n12837), .Z(n12836) );
  AND U14071 ( .A(n15698), .B(n15699), .Z(n12837) );
  XOR U14072 ( .A(n12840), .B(n12839), .Z(n12838) );
  AND U14073 ( .A(n15700), .B(n15701), .Z(n12839) );
  XOR U14074 ( .A(n12842), .B(n12841), .Z(n12840) );
  AND U14075 ( .A(n15702), .B(n15703), .Z(n12841) );
  XOR U14076 ( .A(n12844), .B(n12843), .Z(n12842) );
  AND U14077 ( .A(n15704), .B(n15705), .Z(n12843) );
  XOR U14078 ( .A(n12846), .B(n12845), .Z(n12844) );
  AND U14079 ( .A(n15706), .B(n15707), .Z(n12845) );
  XOR U14080 ( .A(n12848), .B(n12847), .Z(n12846) );
  AND U14081 ( .A(n15708), .B(n15709), .Z(n12847) );
  XOR U14082 ( .A(n12850), .B(n12849), .Z(n12848) );
  AND U14083 ( .A(n15710), .B(n15711), .Z(n12849) );
  XOR U14084 ( .A(n12852), .B(n12851), .Z(n12850) );
  AND U14085 ( .A(n15712), .B(n15713), .Z(n12851) );
  XOR U14086 ( .A(n12854), .B(n12853), .Z(n12852) );
  AND U14087 ( .A(n15714), .B(n15715), .Z(n12853) );
  XOR U14088 ( .A(n12856), .B(n12855), .Z(n12854) );
  AND U14089 ( .A(n15716), .B(n15717), .Z(n12855) );
  XOR U14090 ( .A(n12858), .B(n12857), .Z(n12856) );
  AND U14091 ( .A(n15718), .B(n15719), .Z(n12857) );
  XOR U14092 ( .A(n12860), .B(n12859), .Z(n12858) );
  AND U14093 ( .A(n15720), .B(n15721), .Z(n12859) );
  XOR U14094 ( .A(n12862), .B(n12861), .Z(n12860) );
  AND U14095 ( .A(n15722), .B(n15723), .Z(n12861) );
  XOR U14096 ( .A(n12864), .B(n12863), .Z(n12862) );
  AND U14097 ( .A(n15724), .B(n15725), .Z(n12863) );
  XOR U14098 ( .A(n12866), .B(n12865), .Z(n12864) );
  AND U14099 ( .A(n15726), .B(n15727), .Z(n12865) );
  XOR U14100 ( .A(n12868), .B(n12867), .Z(n12866) );
  AND U14101 ( .A(n15728), .B(n15729), .Z(n12867) );
  XOR U14102 ( .A(n12870), .B(n12869), .Z(n12868) );
  AND U14103 ( .A(n15730), .B(n15731), .Z(n12869) );
  XOR U14104 ( .A(n12872), .B(n12871), .Z(n12870) );
  AND U14105 ( .A(n15732), .B(n15733), .Z(n12871) );
  XOR U14106 ( .A(n12874), .B(n12873), .Z(n12872) );
  AND U14107 ( .A(n15734), .B(n15735), .Z(n12873) );
  XOR U14108 ( .A(n12876), .B(n12875), .Z(n12874) );
  AND U14109 ( .A(n15736), .B(n15737), .Z(n12875) );
  XOR U14110 ( .A(n12885), .B(n12877), .Z(n12876) );
  AND U14111 ( .A(n15738), .B(n15739), .Z(n12877) );
  XOR U14112 ( .A(n12880), .B(n12886), .Z(n12885) );
  AND U14113 ( .A(n15740), .B(n15741), .Z(n12886) );
  XOR U14114 ( .A(n12882), .B(n12881), .Z(n12880) );
  AND U14115 ( .A(n15742), .B(n15743), .Z(n12881) );
  XOR U14116 ( .A(n12906), .B(n12883), .Z(n12882) );
  AND U14117 ( .A(n15744), .B(n15745), .Z(n12883) );
  XOR U14118 ( .A(n12901), .B(n12907), .Z(n12906) );
  AND U14119 ( .A(n15746), .B(n15747), .Z(n12907) );
  XOR U14120 ( .A(n12903), .B(n12902), .Z(n12901) );
  AND U14121 ( .A(n15748), .B(n15749), .Z(n12902) );
  XOR U14122 ( .A(n12891), .B(n12904), .Z(n12903) );
  AND U14123 ( .A(n15750), .B(n15751), .Z(n12904) );
  XOR U14124 ( .A(n12893), .B(n12892), .Z(n12891) );
  AND U14125 ( .A(n15752), .B(n15753), .Z(n12892) );
  XOR U14126 ( .A(n12895), .B(n12894), .Z(n12893) );
  AND U14127 ( .A(n15754), .B(n15755), .Z(n12894) );
  XOR U14128 ( .A(n12897), .B(n12896), .Z(n12895) );
  AND U14129 ( .A(n15756), .B(n15757), .Z(n12896) );
  XOR U14130 ( .A(n12926), .B(n12898), .Z(n12897) );
  AND U14131 ( .A(n15758), .B(n15759), .Z(n12898) );
  XOR U14132 ( .A(n12922), .B(n12927), .Z(n12926) );
  AND U14133 ( .A(n15760), .B(n15761), .Z(n12927) );
  XOR U14134 ( .A(n12924), .B(n12923), .Z(n12922) );
  AND U14135 ( .A(n15762), .B(n15763), .Z(n12923) );
  XOR U14136 ( .A(n12912), .B(n12925), .Z(n12924) );
  AND U14137 ( .A(n15764), .B(n15765), .Z(n12925) );
  XOR U14138 ( .A(n12914), .B(n12913), .Z(n12912) );
  AND U14139 ( .A(n15766), .B(n15767), .Z(n12913) );
  XOR U14140 ( .A(n12916), .B(n12915), .Z(n12914) );
  AND U14141 ( .A(n15768), .B(n15769), .Z(n12915) );
  XOR U14142 ( .A(n12918), .B(n12917), .Z(n12916) );
  AND U14143 ( .A(n15770), .B(n15771), .Z(n12917) );
  XOR U14144 ( .A(n12960), .B(n12919), .Z(n12918) );
  AND U14145 ( .A(n15772), .B(n15773), .Z(n12919) );
  XNOR U14146 ( .A(n12957), .B(n12961), .Z(n12960) );
  AND U14147 ( .A(n15774), .B(n15775), .Z(n12961) );
  XOR U14148 ( .A(n12956), .B(n12948), .Z(n12957) );
  AND U14149 ( .A(n15776), .B(n15777), .Z(n12948) );
  XNOR U14150 ( .A(n12951), .B(n12947), .Z(n12956) );
  AND U14151 ( .A(n15778), .B(n15779), .Z(n12947) );
  XOR U14152 ( .A(n12964), .B(n12952), .Z(n12951) );
  AND U14153 ( .A(n15780), .B(n15781), .Z(n12952) );
  XNOR U14154 ( .A(n12944), .B(n12965), .Z(n12964) );
  AND U14155 ( .A(n15782), .B(n15783), .Z(n12965) );
  XOR U14156 ( .A(n12943), .B(n12935), .Z(n12944) );
  AND U14157 ( .A(n15784), .B(n15785), .Z(n12935) );
  XNOR U14158 ( .A(n12938), .B(n12934), .Z(n12943) );
  AND U14159 ( .A(n15786), .B(n15787), .Z(n12934) );
  XOR U14160 ( .A(n15788), .B(n15789), .Z(n12938) );
  XOR U14161 ( .A(n15790), .B(n15791), .Z(n15789) );
  XOR U14162 ( .A(n15792), .B(n15793), .Z(n15791) );
  XNOR U14163 ( .A(n12981), .B(n12974), .Z(n15793) );
  XOR U14164 ( .A(n15794), .B(n15795), .Z(n12974) );
  XOR U14165 ( .A(n15796), .B(n15797), .Z(n15795) );
  NOR U14166 ( .A(n15798), .B(n15799), .Z(n15797) );
  NOR U14167 ( .A(n15800), .B(n15801), .Z(n15796) );
  AND U14168 ( .A(n15802), .B(n15803), .Z(n15801) );
  IV U14169 ( .A(n15804), .Z(n15800) );
  NOR U14170 ( .A(n15805), .B(n15806), .Z(n15804) );
  AND U14171 ( .A(n15798), .B(n15807), .Z(n15806) );
  AND U14172 ( .A(n15799), .B(n15808), .Z(n15805) );
  XNOR U14173 ( .A(n15809), .B(n15810), .Z(n15794) );
  AND U14174 ( .A(n15811), .B(n15812), .Z(n15810) );
  AND U14175 ( .A(n15813), .B(n15814), .Z(n15809) );
  NOR U14176 ( .A(n15815), .B(n15816), .Z(n15814) );
  IV U14177 ( .A(n15817), .Z(n15815) );
  NOR U14178 ( .A(n15818), .B(n15819), .Z(n15817) );
  NOR U14179 ( .A(n15820), .B(n15821), .Z(n15813) );
  AND U14180 ( .A(n15822), .B(n15823), .Z(n12981) );
  XOR U14181 ( .A(n12979), .B(n12980), .Z(n15792) );
  AND U14182 ( .A(n15824), .B(n15825), .Z(n12980) );
  AND U14183 ( .A(n15826), .B(n15827), .Z(n12979) );
  XOR U14184 ( .A(n15828), .B(n15829), .Z(n15790) );
  XOR U14185 ( .A(n12975), .B(n12976), .Z(n15829) );
  AND U14186 ( .A(n15830), .B(n15831), .Z(n12976) );
  AND U14187 ( .A(n15832), .B(n15833), .Z(n12975) );
  XOR U14188 ( .A(n12973), .B(n12971), .Z(n15828) );
  AND U14189 ( .A(n15834), .B(n15835), .Z(n12971) );
  AND U14190 ( .A(n15836), .B(n15837), .Z(n12973) );
  XNOR U14191 ( .A(n12982), .B(n12939), .Z(n15788) );
  AND U14192 ( .A(n15838), .B(n15839), .Z(n12939) );
  AND U14193 ( .A(n15840), .B(n15841), .Z(n12982) );
  XOR U14194 ( .A(n15842), .B(n15843), .Z(n12995) );
  AND U14195 ( .A(n15842), .B(n15844), .Z(n15843) );
  XNOR U14196 ( .A(n15845), .B(n15846), .Z(n12998) );
  AND U14197 ( .A(n15845), .B(n15847), .Z(n15846) );
  XNOR U14198 ( .A(n15848), .B(n15849), .Z(n13001) );
  AND U14199 ( .A(n15848), .B(n15850), .Z(n15849) );
  XNOR U14200 ( .A(n15851), .B(n15852), .Z(n13004) );
  AND U14201 ( .A(n15851), .B(n15853), .Z(n15852) );
  XNOR U14202 ( .A(n15854), .B(n15855), .Z(n13007) );
  AND U14203 ( .A(n15856), .B(n15854), .Z(n15855) );
  XOR U14204 ( .A(n15857), .B(n15858), .Z(n13010) );
  NOR U14205 ( .A(n15859), .B(n15857), .Z(n15858) );
  XOR U14206 ( .A(n15860), .B(n15861), .Z(n13013) );
  NOR U14207 ( .A(n15862), .B(n15860), .Z(n15861) );
  XOR U14208 ( .A(n15863), .B(n15864), .Z(n13016) );
  NOR U14209 ( .A(n15865), .B(n15863), .Z(n15864) );
  XOR U14210 ( .A(n15866), .B(n15867), .Z(n13019) );
  NOR U14211 ( .A(n15868), .B(n15866), .Z(n15867) );
  XOR U14212 ( .A(n15869), .B(n15870), .Z(n13022) );
  NOR U14213 ( .A(n15871), .B(n15869), .Z(n15870) );
  XOR U14214 ( .A(n15872), .B(n15873), .Z(n13025) );
  NOR U14215 ( .A(n15874), .B(n15872), .Z(n15873) );
  XOR U14216 ( .A(n15875), .B(n15876), .Z(n13028) );
  NOR U14217 ( .A(n15877), .B(n15875), .Z(n15876) );
  XOR U14218 ( .A(n15878), .B(n15879), .Z(n13031) );
  NOR U14219 ( .A(n15880), .B(n15878), .Z(n15879) );
  XOR U14220 ( .A(n15881), .B(n15882), .Z(n13034) );
  NOR U14221 ( .A(n15883), .B(n15881), .Z(n15882) );
  XOR U14222 ( .A(n15884), .B(n15885), .Z(n13037) );
  NOR U14223 ( .A(n15886), .B(n15884), .Z(n15885) );
  XOR U14224 ( .A(n15887), .B(n15888), .Z(n13040) );
  NOR U14225 ( .A(n15889), .B(n15887), .Z(n15888) );
  XOR U14226 ( .A(n15890), .B(n15891), .Z(n13043) );
  NOR U14227 ( .A(n15892), .B(n15890), .Z(n15891) );
  XOR U14228 ( .A(n15893), .B(n15894), .Z(n13046) );
  NOR U14229 ( .A(n15895), .B(n15893), .Z(n15894) );
  XOR U14230 ( .A(n15896), .B(n15897), .Z(n13049) );
  NOR U14231 ( .A(n15898), .B(n15896), .Z(n15897) );
  XOR U14232 ( .A(n15899), .B(n15900), .Z(n13052) );
  NOR U14233 ( .A(n15901), .B(n15899), .Z(n15900) );
  XOR U14234 ( .A(n15902), .B(n15903), .Z(n13055) );
  NOR U14235 ( .A(n15904), .B(n15902), .Z(n15903) );
  XOR U14236 ( .A(n15905), .B(n15906), .Z(n13058) );
  NOR U14237 ( .A(n15907), .B(n15905), .Z(n15906) );
  XOR U14238 ( .A(n15908), .B(n15909), .Z(n13061) );
  NOR U14239 ( .A(n15910), .B(n15908), .Z(n15909) );
  XOR U14240 ( .A(n15911), .B(n15912), .Z(n13064) );
  NOR U14241 ( .A(n15913), .B(n15911), .Z(n15912) );
  XOR U14242 ( .A(n15914), .B(n15915), .Z(n13067) );
  NOR U14243 ( .A(n15916), .B(n15914), .Z(n15915) );
  XOR U14244 ( .A(n15917), .B(n15918), .Z(n13070) );
  NOR U14245 ( .A(n15919), .B(n15917), .Z(n15918) );
  XOR U14246 ( .A(n15920), .B(n15921), .Z(n13073) );
  NOR U14247 ( .A(n15922), .B(n15920), .Z(n15921) );
  XOR U14248 ( .A(n15923), .B(n15924), .Z(n13076) );
  NOR U14249 ( .A(n15925), .B(n15923), .Z(n15924) );
  XOR U14250 ( .A(n15926), .B(n15927), .Z(n13079) );
  NOR U14251 ( .A(n15928), .B(n15926), .Z(n15927) );
  XOR U14252 ( .A(n15929), .B(n15930), .Z(n13082) );
  NOR U14253 ( .A(n15931), .B(n15929), .Z(n15930) );
  XOR U14254 ( .A(n15932), .B(n15933), .Z(n13085) );
  NOR U14255 ( .A(n15934), .B(n15932), .Z(n15933) );
  XOR U14256 ( .A(n15935), .B(n15936), .Z(n13088) );
  NOR U14257 ( .A(n15937), .B(n15935), .Z(n15936) );
  XOR U14258 ( .A(n15938), .B(n15939), .Z(n13091) );
  NOR U14259 ( .A(n15940), .B(n15938), .Z(n15939) );
  XOR U14260 ( .A(n15941), .B(n15942), .Z(n13094) );
  NOR U14261 ( .A(n15943), .B(n15941), .Z(n15942) );
  XOR U14262 ( .A(n15944), .B(n15945), .Z(n13097) );
  NOR U14263 ( .A(n15946), .B(n15944), .Z(n15945) );
  XOR U14264 ( .A(n15947), .B(n15948), .Z(n13100) );
  NOR U14265 ( .A(n15949), .B(n15947), .Z(n15948) );
  XOR U14266 ( .A(n15950), .B(n15951), .Z(n13103) );
  NOR U14267 ( .A(n15952), .B(n15950), .Z(n15951) );
  XOR U14268 ( .A(n15953), .B(n15954), .Z(n13106) );
  NOR U14269 ( .A(n15955), .B(n15953), .Z(n15954) );
  XOR U14270 ( .A(n15956), .B(n15957), .Z(n13109) );
  NOR U14271 ( .A(n15958), .B(n15956), .Z(n15957) );
  XOR U14272 ( .A(n15959), .B(n15960), .Z(n13112) );
  NOR U14273 ( .A(n15961), .B(n15959), .Z(n15960) );
  XOR U14274 ( .A(n15962), .B(n15963), .Z(n13115) );
  NOR U14275 ( .A(n15964), .B(n15962), .Z(n15963) );
  XOR U14276 ( .A(n15965), .B(n15966), .Z(n13118) );
  NOR U14277 ( .A(n15967), .B(n15965), .Z(n15966) );
  XOR U14278 ( .A(n15968), .B(n15969), .Z(n13121) );
  NOR U14279 ( .A(n15970), .B(n15968), .Z(n15969) );
  XOR U14280 ( .A(n15971), .B(n15972), .Z(n13124) );
  NOR U14281 ( .A(n15973), .B(n15971), .Z(n15972) );
  XOR U14282 ( .A(n15974), .B(n15975), .Z(n13127) );
  NOR U14283 ( .A(n15976), .B(n15974), .Z(n15975) );
  XOR U14284 ( .A(n15977), .B(n15978), .Z(n13130) );
  NOR U14285 ( .A(n15979), .B(n15977), .Z(n15978) );
  XOR U14286 ( .A(n15980), .B(n15981), .Z(n13133) );
  NOR U14287 ( .A(n15982), .B(n15980), .Z(n15981) );
  XOR U14288 ( .A(n15983), .B(n15984), .Z(n13136) );
  NOR U14289 ( .A(n15985), .B(n15983), .Z(n15984) );
  XOR U14290 ( .A(n15986), .B(n15987), .Z(n13139) );
  NOR U14291 ( .A(n15988), .B(n15986), .Z(n15987) );
  XOR U14292 ( .A(n15989), .B(n15990), .Z(n13142) );
  NOR U14293 ( .A(n15991), .B(n15989), .Z(n15990) );
  XOR U14294 ( .A(n15992), .B(n15993), .Z(n13145) );
  NOR U14295 ( .A(n15994), .B(n15992), .Z(n15993) );
  XOR U14296 ( .A(n15995), .B(n15996), .Z(n13148) );
  NOR U14297 ( .A(n15997), .B(n15995), .Z(n15996) );
  XOR U14298 ( .A(n15998), .B(n15999), .Z(n13151) );
  NOR U14299 ( .A(n16000), .B(n15998), .Z(n15999) );
  XOR U14300 ( .A(n16001), .B(n16002), .Z(n13154) );
  NOR U14301 ( .A(n16003), .B(n16001), .Z(n16002) );
  XOR U14302 ( .A(n16004), .B(n16005), .Z(n13157) );
  NOR U14303 ( .A(n16006), .B(n16004), .Z(n16005) );
  XOR U14304 ( .A(n16007), .B(n16008), .Z(n13160) );
  NOR U14305 ( .A(n16009), .B(n16007), .Z(n16008) );
  XOR U14306 ( .A(n16010), .B(n16011), .Z(n13163) );
  NOR U14307 ( .A(n16012), .B(n16010), .Z(n16011) );
  XOR U14308 ( .A(n16013), .B(n16014), .Z(n13166) );
  NOR U14309 ( .A(n16015), .B(n16013), .Z(n16014) );
  XOR U14310 ( .A(n16016), .B(n16017), .Z(n13169) );
  NOR U14311 ( .A(n16018), .B(n16016), .Z(n16017) );
  XOR U14312 ( .A(n16019), .B(n16020), .Z(n13172) );
  NOR U14313 ( .A(n16021), .B(n16019), .Z(n16020) );
  XOR U14314 ( .A(n16022), .B(n16023), .Z(n13175) );
  NOR U14315 ( .A(n16024), .B(n16022), .Z(n16023) );
  XOR U14316 ( .A(n16025), .B(n16026), .Z(n13178) );
  NOR U14317 ( .A(n16027), .B(n16025), .Z(n16026) );
  XOR U14318 ( .A(n16028), .B(n16029), .Z(n13181) );
  NOR U14319 ( .A(n16030), .B(n16028), .Z(n16029) );
  XOR U14320 ( .A(n16031), .B(n16032), .Z(n13184) );
  NOR U14321 ( .A(n16033), .B(n16031), .Z(n16032) );
  XOR U14322 ( .A(n16034), .B(n16035), .Z(n13187) );
  NOR U14323 ( .A(n16036), .B(n16034), .Z(n16035) );
  XOR U14324 ( .A(n16037), .B(n16038), .Z(n13190) );
  NOR U14325 ( .A(n16039), .B(n16037), .Z(n16038) );
  XOR U14326 ( .A(n16040), .B(n16041), .Z(n13193) );
  NOR U14327 ( .A(n16042), .B(n16040), .Z(n16041) );
  XOR U14328 ( .A(n16043), .B(n16044), .Z(n13196) );
  NOR U14329 ( .A(n16045), .B(n16043), .Z(n16044) );
  XOR U14330 ( .A(n16046), .B(n16047), .Z(n13199) );
  NOR U14331 ( .A(n16048), .B(n16046), .Z(n16047) );
  XOR U14332 ( .A(n16049), .B(n16050), .Z(n13202) );
  NOR U14333 ( .A(n16051), .B(n16049), .Z(n16050) );
  XOR U14334 ( .A(n16052), .B(n16053), .Z(n13205) );
  NOR U14335 ( .A(n16054), .B(n16052), .Z(n16053) );
  XOR U14336 ( .A(n16055), .B(n16056), .Z(n13208) );
  NOR U14337 ( .A(n16057), .B(n16055), .Z(n16056) );
  XOR U14338 ( .A(n16058), .B(n16059), .Z(n13211) );
  NOR U14339 ( .A(n16060), .B(n16058), .Z(n16059) );
  XOR U14340 ( .A(n16061), .B(n16062), .Z(n13214) );
  NOR U14341 ( .A(n16063), .B(n16061), .Z(n16062) );
  XOR U14342 ( .A(n16064), .B(n16065), .Z(n13217) );
  NOR U14343 ( .A(n16066), .B(n16064), .Z(n16065) );
  XOR U14344 ( .A(n16067), .B(n16068), .Z(n13220) );
  NOR U14345 ( .A(n16069), .B(n16067), .Z(n16068) );
  XOR U14346 ( .A(n16070), .B(n16071), .Z(n13223) );
  NOR U14347 ( .A(n16072), .B(n16070), .Z(n16071) );
  XOR U14348 ( .A(n16073), .B(n16074), .Z(n13226) );
  NOR U14349 ( .A(n16075), .B(n16073), .Z(n16074) );
  XOR U14350 ( .A(n16076), .B(n16077), .Z(n13229) );
  NOR U14351 ( .A(n16078), .B(n16076), .Z(n16077) );
  XOR U14352 ( .A(n16079), .B(n16080), .Z(n13232) );
  NOR U14353 ( .A(n16081), .B(n16079), .Z(n16080) );
  XOR U14354 ( .A(n16082), .B(n16083), .Z(n13235) );
  NOR U14355 ( .A(n16084), .B(n16082), .Z(n16083) );
  XOR U14356 ( .A(n16085), .B(n16086), .Z(n13238) );
  NOR U14357 ( .A(n16087), .B(n16085), .Z(n16086) );
  XOR U14358 ( .A(n16088), .B(n16089), .Z(n13241) );
  NOR U14359 ( .A(n16090), .B(n16088), .Z(n16089) );
  XOR U14360 ( .A(n16091), .B(n16092), .Z(n13244) );
  NOR U14361 ( .A(n16093), .B(n16091), .Z(n16092) );
  XOR U14362 ( .A(n16094), .B(n16095), .Z(n13247) );
  NOR U14363 ( .A(n16096), .B(n16094), .Z(n16095) );
  XOR U14364 ( .A(n16097), .B(n16098), .Z(n13250) );
  NOR U14365 ( .A(n16099), .B(n16097), .Z(n16098) );
  XOR U14366 ( .A(n16100), .B(n16101), .Z(n13253) );
  NOR U14367 ( .A(n16102), .B(n16100), .Z(n16101) );
  XOR U14368 ( .A(n16103), .B(n16104), .Z(n13256) );
  NOR U14369 ( .A(n16105), .B(n16103), .Z(n16104) );
  XOR U14370 ( .A(n16106), .B(n16107), .Z(n13259) );
  NOR U14371 ( .A(n16108), .B(n16106), .Z(n16107) );
  XOR U14372 ( .A(n16109), .B(n16110), .Z(n13262) );
  NOR U14373 ( .A(n16111), .B(n16109), .Z(n16110) );
  XOR U14374 ( .A(n16112), .B(n16113), .Z(n13265) );
  NOR U14375 ( .A(n16114), .B(n16112), .Z(n16113) );
  XOR U14376 ( .A(n16115), .B(n16116), .Z(n13268) );
  NOR U14377 ( .A(n16117), .B(n16115), .Z(n16116) );
  XOR U14378 ( .A(n16118), .B(n16119), .Z(n13271) );
  NOR U14379 ( .A(n16120), .B(n16118), .Z(n16119) );
  XOR U14380 ( .A(n16121), .B(n16122), .Z(n13274) );
  NOR U14381 ( .A(n16123), .B(n16121), .Z(n16122) );
  XOR U14382 ( .A(n16124), .B(n16125), .Z(n13277) );
  NOR U14383 ( .A(n16126), .B(n16124), .Z(n16125) );
  XOR U14384 ( .A(n16127), .B(n16128), .Z(n13280) );
  NOR U14385 ( .A(n16129), .B(n16127), .Z(n16128) );
  XOR U14386 ( .A(n16130), .B(n16131), .Z(n13283) );
  NOR U14387 ( .A(n16132), .B(n16130), .Z(n16131) );
  XOR U14388 ( .A(n16133), .B(n16134), .Z(n13286) );
  NOR U14389 ( .A(n16135), .B(n16133), .Z(n16134) );
  XOR U14390 ( .A(n16136), .B(n16137), .Z(n13289) );
  NOR U14391 ( .A(n16138), .B(n16136), .Z(n16137) );
  XOR U14392 ( .A(n16139), .B(n16140), .Z(n13292) );
  NOR U14393 ( .A(n16141), .B(n16139), .Z(n16140) );
  XOR U14394 ( .A(n16142), .B(n16143), .Z(n13295) );
  NOR U14395 ( .A(n16144), .B(n16142), .Z(n16143) );
  XOR U14396 ( .A(n16145), .B(n16146), .Z(n13298) );
  NOR U14397 ( .A(n16147), .B(n16145), .Z(n16146) );
  XOR U14398 ( .A(n16148), .B(n16149), .Z(n13301) );
  NOR U14399 ( .A(n16150), .B(n16148), .Z(n16149) );
  XOR U14400 ( .A(n16151), .B(n16152), .Z(n13304) );
  NOR U14401 ( .A(n16153), .B(n16151), .Z(n16152) );
  XOR U14402 ( .A(n16154), .B(n16155), .Z(n13307) );
  NOR U14403 ( .A(n16156), .B(n16154), .Z(n16155) );
  XOR U14404 ( .A(n16157), .B(n16158), .Z(n13310) );
  NOR U14405 ( .A(n16159), .B(n16157), .Z(n16158) );
  XOR U14406 ( .A(n16160), .B(n16161), .Z(n13313) );
  NOR U14407 ( .A(n16162), .B(n16160), .Z(n16161) );
  XOR U14408 ( .A(n16163), .B(n16164), .Z(n13316) );
  NOR U14409 ( .A(n16165), .B(n16163), .Z(n16164) );
  XOR U14410 ( .A(n16166), .B(n16167), .Z(n13319) );
  NOR U14411 ( .A(n16168), .B(n16166), .Z(n16167) );
  XOR U14412 ( .A(n16169), .B(n16170), .Z(n13322) );
  NOR U14413 ( .A(n16171), .B(n16169), .Z(n16170) );
  XOR U14414 ( .A(n16172), .B(n16173), .Z(n13325) );
  NOR U14415 ( .A(n16174), .B(n16172), .Z(n16173) );
  XOR U14416 ( .A(n16175), .B(n16176), .Z(n13328) );
  NOR U14417 ( .A(n16177), .B(n16175), .Z(n16176) );
  XOR U14418 ( .A(n16178), .B(n16179), .Z(n13331) );
  NOR U14419 ( .A(n16180), .B(n16178), .Z(n16179) );
  XOR U14420 ( .A(n16181), .B(n16182), .Z(n13334) );
  NOR U14421 ( .A(n16183), .B(n16181), .Z(n16182) );
  XOR U14422 ( .A(n16184), .B(n16185), .Z(n13337) );
  NOR U14423 ( .A(n16186), .B(n16184), .Z(n16185) );
  XOR U14424 ( .A(n16187), .B(n16188), .Z(n13340) );
  NOR U14425 ( .A(n16189), .B(n16187), .Z(n16188) );
  XOR U14426 ( .A(n16190), .B(n16191), .Z(n13343) );
  NOR U14427 ( .A(n16192), .B(n16190), .Z(n16191) );
  XOR U14428 ( .A(n16193), .B(n16194), .Z(n13346) );
  NOR U14429 ( .A(n16195), .B(n16193), .Z(n16194) );
  XOR U14430 ( .A(n16196), .B(n16197), .Z(n13349) );
  NOR U14431 ( .A(n16198), .B(n16196), .Z(n16197) );
  XOR U14432 ( .A(n16199), .B(n16200), .Z(n13352) );
  NOR U14433 ( .A(n16201), .B(n16199), .Z(n16200) );
  XOR U14434 ( .A(n16202), .B(n16203), .Z(n13355) );
  NOR U14435 ( .A(n16204), .B(n16202), .Z(n16203) );
  XOR U14436 ( .A(n16205), .B(n16206), .Z(n13358) );
  NOR U14437 ( .A(n16207), .B(n16205), .Z(n16206) );
  XOR U14438 ( .A(n16208), .B(n16209), .Z(n13361) );
  NOR U14439 ( .A(n16210), .B(n16208), .Z(n16209) );
  XOR U14440 ( .A(n16211), .B(n16212), .Z(n13364) );
  NOR U14441 ( .A(n16213), .B(n16211), .Z(n16212) );
  XOR U14442 ( .A(n16214), .B(n16215), .Z(n13367) );
  NOR U14443 ( .A(n16216), .B(n16214), .Z(n16215) );
  XOR U14444 ( .A(n16217), .B(n16218), .Z(n13370) );
  NOR U14445 ( .A(n16219), .B(n16217), .Z(n16218) );
  XOR U14446 ( .A(n16220), .B(n16221), .Z(n13373) );
  NOR U14447 ( .A(n16222), .B(n16220), .Z(n16221) );
  XOR U14448 ( .A(n16223), .B(n16224), .Z(n13376) );
  NOR U14449 ( .A(n16225), .B(n16223), .Z(n16224) );
  XOR U14450 ( .A(n16226), .B(n16227), .Z(n13379) );
  NOR U14451 ( .A(n16228), .B(n16226), .Z(n16227) );
  XOR U14452 ( .A(n16229), .B(n16230), .Z(n13382) );
  NOR U14453 ( .A(n16231), .B(n16229), .Z(n16230) );
  XOR U14454 ( .A(n16232), .B(n16233), .Z(n13385) );
  NOR U14455 ( .A(n16234), .B(n16232), .Z(n16233) );
  XOR U14456 ( .A(n16235), .B(n16236), .Z(n13388) );
  NOR U14457 ( .A(n16237), .B(n16235), .Z(n16236) );
  XOR U14458 ( .A(n16238), .B(n16239), .Z(n13391) );
  NOR U14459 ( .A(n16240), .B(n16238), .Z(n16239) );
  XOR U14460 ( .A(n16241), .B(n16242), .Z(n13394) );
  NOR U14461 ( .A(n16243), .B(n16241), .Z(n16242) );
  XOR U14462 ( .A(n16244), .B(n16245), .Z(n13397) );
  NOR U14463 ( .A(n16246), .B(n16244), .Z(n16245) );
  XOR U14464 ( .A(n16247), .B(n16248), .Z(n13400) );
  NOR U14465 ( .A(n16249), .B(n16247), .Z(n16248) );
  XOR U14466 ( .A(n16250), .B(n16251), .Z(n13403) );
  NOR U14467 ( .A(n16252), .B(n16250), .Z(n16251) );
  XOR U14468 ( .A(n16253), .B(n16254), .Z(n13406) );
  NOR U14469 ( .A(n16255), .B(n16253), .Z(n16254) );
  XOR U14470 ( .A(n16256), .B(n16257), .Z(n13409) );
  NOR U14471 ( .A(n16258), .B(n16256), .Z(n16257) );
  XOR U14472 ( .A(n16259), .B(n16260), .Z(n13412) );
  NOR U14473 ( .A(n16261), .B(n16259), .Z(n16260) );
  XOR U14474 ( .A(n16262), .B(n16263), .Z(n13415) );
  NOR U14475 ( .A(n16264), .B(n16262), .Z(n16263) );
  XOR U14476 ( .A(n16265), .B(n16266), .Z(n13418) );
  NOR U14477 ( .A(n16267), .B(n16265), .Z(n16266) );
  XOR U14478 ( .A(n16268), .B(n16269), .Z(n13421) );
  NOR U14479 ( .A(n16270), .B(n16268), .Z(n16269) );
  XOR U14480 ( .A(n16271), .B(n16272), .Z(n13424) );
  NOR U14481 ( .A(n16273), .B(n16271), .Z(n16272) );
  XOR U14482 ( .A(n16274), .B(n16275), .Z(n13427) );
  NOR U14483 ( .A(n16276), .B(n16274), .Z(n16275) );
  XOR U14484 ( .A(n16277), .B(n16278), .Z(n13430) );
  NOR U14485 ( .A(n16279), .B(n16277), .Z(n16278) );
  XOR U14486 ( .A(n16280), .B(n16281), .Z(n13433) );
  NOR U14487 ( .A(n16282), .B(n16280), .Z(n16281) );
  XOR U14488 ( .A(n16283), .B(n16284), .Z(n13436) );
  NOR U14489 ( .A(n16285), .B(n16283), .Z(n16284) );
  XOR U14490 ( .A(n16286), .B(n16287), .Z(n13439) );
  NOR U14491 ( .A(n16288), .B(n16286), .Z(n16287) );
  XOR U14492 ( .A(n16289), .B(n16290), .Z(n13442) );
  NOR U14493 ( .A(n16291), .B(n16289), .Z(n16290) );
  XOR U14494 ( .A(n16292), .B(n16293), .Z(n13445) );
  NOR U14495 ( .A(n16294), .B(n16292), .Z(n16293) );
  XOR U14496 ( .A(n16295), .B(n16296), .Z(n13448) );
  NOR U14497 ( .A(n16297), .B(n16295), .Z(n16296) );
  XOR U14498 ( .A(n16298), .B(n16299), .Z(n13451) );
  NOR U14499 ( .A(n16300), .B(n16298), .Z(n16299) );
  XOR U14500 ( .A(n16301), .B(n16302), .Z(n13454) );
  NOR U14501 ( .A(n16303), .B(n16301), .Z(n16302) );
  XOR U14502 ( .A(n16304), .B(n16305), .Z(n13457) );
  NOR U14503 ( .A(n16306), .B(n16304), .Z(n16305) );
  XOR U14504 ( .A(n16307), .B(n16308), .Z(n13460) );
  NOR U14505 ( .A(n16309), .B(n16307), .Z(n16308) );
  XOR U14506 ( .A(n16310), .B(n16311), .Z(n13463) );
  NOR U14507 ( .A(n16312), .B(n16310), .Z(n16311) );
  XOR U14508 ( .A(n16313), .B(n16314), .Z(n13466) );
  NOR U14509 ( .A(n16315), .B(n16313), .Z(n16314) );
  XOR U14510 ( .A(n16316), .B(n16317), .Z(n13469) );
  NOR U14511 ( .A(n16318), .B(n16316), .Z(n16317) );
  XOR U14512 ( .A(n16319), .B(n16320), .Z(n13472) );
  NOR U14513 ( .A(n16321), .B(n16319), .Z(n16320) );
  XOR U14514 ( .A(n16322), .B(n16323), .Z(n13475) );
  NOR U14515 ( .A(n16324), .B(n16322), .Z(n16323) );
  XOR U14516 ( .A(n16325), .B(n16326), .Z(n13478) );
  NOR U14517 ( .A(n16327), .B(n16325), .Z(n16326) );
  XOR U14518 ( .A(n16328), .B(n16329), .Z(n13481) );
  NOR U14519 ( .A(n16330), .B(n16328), .Z(n16329) );
  XOR U14520 ( .A(n16331), .B(n16332), .Z(n13484) );
  NOR U14521 ( .A(n16333), .B(n16331), .Z(n16332) );
  XOR U14522 ( .A(n16334), .B(n16335), .Z(n13487) );
  NOR U14523 ( .A(n16336), .B(n16334), .Z(n16335) );
  XOR U14524 ( .A(n16337), .B(n16338), .Z(n13490) );
  NOR U14525 ( .A(n16339), .B(n16337), .Z(n16338) );
  XOR U14526 ( .A(n16340), .B(n16341), .Z(n13493) );
  NOR U14527 ( .A(n16342), .B(n16340), .Z(n16341) );
  XOR U14528 ( .A(n16343), .B(n16344), .Z(n13496) );
  NOR U14529 ( .A(n16345), .B(n16343), .Z(n16344) );
  XOR U14530 ( .A(n16346), .B(n16347), .Z(n13499) );
  NOR U14531 ( .A(n16348), .B(n16346), .Z(n16347) );
  XOR U14532 ( .A(n16349), .B(n16350), .Z(n13502) );
  NOR U14533 ( .A(n16351), .B(n16349), .Z(n16350) );
  XOR U14534 ( .A(n16352), .B(n16353), .Z(n13505) );
  NOR U14535 ( .A(n16354), .B(n16352), .Z(n16353) );
  XOR U14536 ( .A(n16355), .B(n16356), .Z(n13508) );
  NOR U14537 ( .A(n16357), .B(n16355), .Z(n16356) );
  XOR U14538 ( .A(n16358), .B(n16359), .Z(n13511) );
  NOR U14539 ( .A(n16360), .B(n16358), .Z(n16359) );
  XOR U14540 ( .A(n16361), .B(n16362), .Z(n13514) );
  NOR U14541 ( .A(n16363), .B(n16361), .Z(n16362) );
  XOR U14542 ( .A(n16364), .B(n16365), .Z(n13517) );
  NOR U14543 ( .A(n16366), .B(n16364), .Z(n16365) );
  XOR U14544 ( .A(n16367), .B(n16368), .Z(n13520) );
  NOR U14545 ( .A(n16369), .B(n16367), .Z(n16368) );
  XOR U14546 ( .A(n16370), .B(n16371), .Z(n13523) );
  NOR U14547 ( .A(n16372), .B(n16370), .Z(n16371) );
  XOR U14548 ( .A(n16373), .B(n16374), .Z(n13526) );
  NOR U14549 ( .A(n16375), .B(n16373), .Z(n16374) );
  XOR U14550 ( .A(n16376), .B(n16377), .Z(n13529) );
  NOR U14551 ( .A(n16378), .B(n16376), .Z(n16377) );
  XOR U14552 ( .A(n16379), .B(n16380), .Z(n13532) );
  NOR U14553 ( .A(n16381), .B(n16379), .Z(n16380) );
  XOR U14554 ( .A(n16382), .B(n16383), .Z(n13535) );
  NOR U14555 ( .A(n16384), .B(n16382), .Z(n16383) );
  XOR U14556 ( .A(n16385), .B(n16386), .Z(n13538) );
  NOR U14557 ( .A(n16387), .B(n16385), .Z(n16386) );
  XOR U14558 ( .A(n16388), .B(n16389), .Z(n13541) );
  NOR U14559 ( .A(n16390), .B(n16388), .Z(n16389) );
  XOR U14560 ( .A(n16391), .B(n16392), .Z(n13544) );
  NOR U14561 ( .A(n16393), .B(n16391), .Z(n16392) );
  XOR U14562 ( .A(n16394), .B(n16395), .Z(n13547) );
  NOR U14563 ( .A(n16396), .B(n16394), .Z(n16395) );
  XOR U14564 ( .A(n16397), .B(n16398), .Z(n13550) );
  NOR U14565 ( .A(n16399), .B(n16397), .Z(n16398) );
  XOR U14566 ( .A(n16400), .B(n16401), .Z(n13553) );
  NOR U14567 ( .A(n16402), .B(n16400), .Z(n16401) );
  XOR U14568 ( .A(n16403), .B(n16404), .Z(n13556) );
  NOR U14569 ( .A(n16405), .B(n16403), .Z(n16404) );
  XOR U14570 ( .A(n16406), .B(n16407), .Z(n13559) );
  NOR U14571 ( .A(n16408), .B(n16406), .Z(n16407) );
  XOR U14572 ( .A(n16409), .B(n16410), .Z(n13562) );
  NOR U14573 ( .A(n16411), .B(n16409), .Z(n16410) );
  XOR U14574 ( .A(n16412), .B(n16413), .Z(n13565) );
  NOR U14575 ( .A(n16414), .B(n16412), .Z(n16413) );
  XOR U14576 ( .A(n16415), .B(n16416), .Z(n13568) );
  NOR U14577 ( .A(n16417), .B(n16415), .Z(n16416) );
  XOR U14578 ( .A(n16418), .B(n16419), .Z(n13571) );
  NOR U14579 ( .A(n16420), .B(n16418), .Z(n16419) );
  XOR U14580 ( .A(n16421), .B(n16422), .Z(n13574) );
  NOR U14581 ( .A(n16423), .B(n16421), .Z(n16422) );
  XOR U14582 ( .A(n16424), .B(n16425), .Z(n13577) );
  NOR U14583 ( .A(n16426), .B(n16424), .Z(n16425) );
  XOR U14584 ( .A(n16427), .B(n16428), .Z(n13580) );
  NOR U14585 ( .A(n16429), .B(n16427), .Z(n16428) );
  XOR U14586 ( .A(n16430), .B(n16431), .Z(n13583) );
  NOR U14587 ( .A(n16432), .B(n16430), .Z(n16431) );
  XOR U14588 ( .A(n16433), .B(n16434), .Z(n13586) );
  NOR U14589 ( .A(n16435), .B(n16433), .Z(n16434) );
  XOR U14590 ( .A(n16436), .B(n16437), .Z(n13589) );
  NOR U14591 ( .A(n16438), .B(n16436), .Z(n16437) );
  XOR U14592 ( .A(n16439), .B(n16440), .Z(n13592) );
  NOR U14593 ( .A(n16441), .B(n16439), .Z(n16440) );
  XOR U14594 ( .A(n16442), .B(n16443), .Z(n13595) );
  NOR U14595 ( .A(n16444), .B(n16442), .Z(n16443) );
  XOR U14596 ( .A(n16445), .B(n16446), .Z(n13598) );
  NOR U14597 ( .A(n16447), .B(n16445), .Z(n16446) );
  XOR U14598 ( .A(n16448), .B(n16449), .Z(n13601) );
  NOR U14599 ( .A(n16450), .B(n16448), .Z(n16449) );
  XOR U14600 ( .A(n16451), .B(n16452), .Z(n13604) );
  NOR U14601 ( .A(n16453), .B(n16451), .Z(n16452) );
  XOR U14602 ( .A(n16454), .B(n16455), .Z(n13607) );
  NOR U14603 ( .A(n16456), .B(n16454), .Z(n16455) );
  XOR U14604 ( .A(n16457), .B(n16458), .Z(n13610) );
  NOR U14605 ( .A(n16459), .B(n16457), .Z(n16458) );
  XOR U14606 ( .A(n16460), .B(n16461), .Z(n13613) );
  NOR U14607 ( .A(n16462), .B(n16460), .Z(n16461) );
  XOR U14608 ( .A(n16463), .B(n16464), .Z(n13616) );
  NOR U14609 ( .A(n16465), .B(n16463), .Z(n16464) );
  XOR U14610 ( .A(n16466), .B(n16467), .Z(n13619) );
  NOR U14611 ( .A(n16468), .B(n16466), .Z(n16467) );
  XOR U14612 ( .A(n16469), .B(n16470), .Z(n13622) );
  NOR U14613 ( .A(n16471), .B(n16469), .Z(n16470) );
  XOR U14614 ( .A(n16472), .B(n16473), .Z(n13625) );
  NOR U14615 ( .A(n16474), .B(n16472), .Z(n16473) );
  XOR U14616 ( .A(n16475), .B(n16476), .Z(n13628) );
  NOR U14617 ( .A(n16477), .B(n16475), .Z(n16476) );
  XOR U14618 ( .A(n16478), .B(n16479), .Z(n13631) );
  NOR U14619 ( .A(n16480), .B(n16478), .Z(n16479) );
  XOR U14620 ( .A(n16481), .B(n16482), .Z(n13634) );
  NOR U14621 ( .A(n16483), .B(n16481), .Z(n16482) );
  XOR U14622 ( .A(n16484), .B(n16485), .Z(n13637) );
  NOR U14623 ( .A(n16486), .B(n16484), .Z(n16485) );
  XOR U14624 ( .A(n16487), .B(n16488), .Z(n13640) );
  NOR U14625 ( .A(n16489), .B(n16487), .Z(n16488) );
  XOR U14626 ( .A(n16490), .B(n16491), .Z(n13643) );
  NOR U14627 ( .A(n16492), .B(n16490), .Z(n16491) );
  XOR U14628 ( .A(n16493), .B(n16494), .Z(n13646) );
  NOR U14629 ( .A(n16495), .B(n16493), .Z(n16494) );
  XOR U14630 ( .A(n16496), .B(n16497), .Z(n13649) );
  NOR U14631 ( .A(n16498), .B(n16496), .Z(n16497) );
  XOR U14632 ( .A(n16499), .B(n16500), .Z(n13652) );
  NOR U14633 ( .A(n16501), .B(n16499), .Z(n16500) );
  XOR U14634 ( .A(n16502), .B(n16503), .Z(n13655) );
  NOR U14635 ( .A(n16504), .B(n16502), .Z(n16503) );
  XOR U14636 ( .A(n16505), .B(n16506), .Z(n13658) );
  NOR U14637 ( .A(n16507), .B(n16505), .Z(n16506) );
  XOR U14638 ( .A(n16508), .B(n16509), .Z(n13661) );
  NOR U14639 ( .A(n16510), .B(n16508), .Z(n16509) );
  XOR U14640 ( .A(n16511), .B(n16512), .Z(n13664) );
  NOR U14641 ( .A(n16513), .B(n16511), .Z(n16512) );
  XOR U14642 ( .A(n16514), .B(n16515), .Z(n13667) );
  NOR U14643 ( .A(n16516), .B(n16514), .Z(n16515) );
  XOR U14644 ( .A(n16517), .B(n16518), .Z(n13670) );
  NOR U14645 ( .A(n16519), .B(n16517), .Z(n16518) );
  XOR U14646 ( .A(n16520), .B(n16521), .Z(n13673) );
  NOR U14647 ( .A(n16522), .B(n16520), .Z(n16521) );
  XOR U14648 ( .A(n16523), .B(n16524), .Z(n13676) );
  NOR U14649 ( .A(n16525), .B(n16523), .Z(n16524) );
  XOR U14650 ( .A(n16526), .B(n16527), .Z(n13679) );
  NOR U14651 ( .A(n16528), .B(n16526), .Z(n16527) );
  XOR U14652 ( .A(n16529), .B(n16530), .Z(n13682) );
  NOR U14653 ( .A(n16531), .B(n16529), .Z(n16530) );
  XOR U14654 ( .A(n16532), .B(n16533), .Z(n13685) );
  NOR U14655 ( .A(n16534), .B(n16532), .Z(n16533) );
  XOR U14656 ( .A(n16535), .B(n16536), .Z(n13688) );
  NOR U14657 ( .A(n16537), .B(n16535), .Z(n16536) );
  XOR U14658 ( .A(n16538), .B(n16539), .Z(n13691) );
  NOR U14659 ( .A(n16540), .B(n16538), .Z(n16539) );
  XOR U14660 ( .A(n16541), .B(n16542), .Z(n13694) );
  NOR U14661 ( .A(n16543), .B(n16541), .Z(n16542) );
  XOR U14662 ( .A(n16544), .B(n16545), .Z(n13697) );
  NOR U14663 ( .A(n16546), .B(n16544), .Z(n16545) );
  XOR U14664 ( .A(n16547), .B(n16548), .Z(n13700) );
  NOR U14665 ( .A(n16549), .B(n16547), .Z(n16548) );
  XOR U14666 ( .A(n16550), .B(n16551), .Z(n13703) );
  NOR U14667 ( .A(n16552), .B(n16550), .Z(n16551) );
  XOR U14668 ( .A(n16553), .B(n16554), .Z(n13706) );
  NOR U14669 ( .A(n16555), .B(n16553), .Z(n16554) );
  XOR U14670 ( .A(n16556), .B(n16557), .Z(n13709) );
  NOR U14671 ( .A(n16558), .B(n16556), .Z(n16557) );
  XOR U14672 ( .A(n16559), .B(n16560), .Z(n13712) );
  NOR U14673 ( .A(n16561), .B(n16559), .Z(n16560) );
  XOR U14674 ( .A(n16562), .B(n16563), .Z(n13715) );
  NOR U14675 ( .A(n16564), .B(n16562), .Z(n16563) );
  XOR U14676 ( .A(n16565), .B(n16566), .Z(n13718) );
  NOR U14677 ( .A(n16567), .B(n16565), .Z(n16566) );
  XOR U14678 ( .A(n16568), .B(n16569), .Z(n13721) );
  NOR U14679 ( .A(n16570), .B(n16568), .Z(n16569) );
  XOR U14680 ( .A(n16571), .B(n16572), .Z(n13724) );
  NOR U14681 ( .A(n16573), .B(n16571), .Z(n16572) );
  XOR U14682 ( .A(n16574), .B(n16575), .Z(n13727) );
  NOR U14683 ( .A(n16576), .B(n16574), .Z(n16575) );
  XOR U14684 ( .A(n16577), .B(n16578), .Z(n13730) );
  NOR U14685 ( .A(n16579), .B(n16577), .Z(n16578) );
  XOR U14686 ( .A(n16580), .B(n16581), .Z(n13733) );
  NOR U14687 ( .A(n16582), .B(n16580), .Z(n16581) );
  XOR U14688 ( .A(n16583), .B(n16584), .Z(n13736) );
  NOR U14689 ( .A(n16585), .B(n16583), .Z(n16584) );
  XOR U14690 ( .A(n16586), .B(n16587), .Z(n13739) );
  NOR U14691 ( .A(n16588), .B(n16586), .Z(n16587) );
  XOR U14692 ( .A(n16589), .B(n16590), .Z(n13742) );
  NOR U14693 ( .A(n16591), .B(n16589), .Z(n16590) );
  XOR U14694 ( .A(n16592), .B(n16593), .Z(n13745) );
  NOR U14695 ( .A(n16594), .B(n16592), .Z(n16593) );
  XOR U14696 ( .A(n16595), .B(n16596), .Z(n13748) );
  NOR U14697 ( .A(n16597), .B(n16595), .Z(n16596) );
  XOR U14698 ( .A(n16598), .B(n16599), .Z(n13751) );
  NOR U14699 ( .A(n16600), .B(n16598), .Z(n16599) );
  XOR U14700 ( .A(n16601), .B(n16602), .Z(n13754) );
  NOR U14701 ( .A(n16603), .B(n16601), .Z(n16602) );
  XOR U14702 ( .A(n16604), .B(n16605), .Z(n13757) );
  NOR U14703 ( .A(n16606), .B(n16604), .Z(n16605) );
  XOR U14704 ( .A(n16607), .B(n16608), .Z(n13760) );
  NOR U14705 ( .A(n16609), .B(n16607), .Z(n16608) );
  XOR U14706 ( .A(n16610), .B(n16611), .Z(n13763) );
  NOR U14707 ( .A(n16612), .B(n16610), .Z(n16611) );
  XOR U14708 ( .A(n16613), .B(n16614), .Z(n13766) );
  NOR U14709 ( .A(n16615), .B(n16613), .Z(n16614) );
  XOR U14710 ( .A(n16616), .B(n16617), .Z(n13769) );
  NOR U14711 ( .A(n16618), .B(n16616), .Z(n16617) );
  XOR U14712 ( .A(n16619), .B(n16620), .Z(n13772) );
  NOR U14713 ( .A(n16621), .B(n16619), .Z(n16620) );
  XOR U14714 ( .A(n16622), .B(n16623), .Z(n13775) );
  NOR U14715 ( .A(n16624), .B(n16622), .Z(n16623) );
  XOR U14716 ( .A(n16625), .B(n16626), .Z(n13778) );
  NOR U14717 ( .A(n16627), .B(n16625), .Z(n16626) );
  XOR U14718 ( .A(n16628), .B(n16629), .Z(n13781) );
  NOR U14719 ( .A(n16630), .B(n16628), .Z(n16629) );
  XOR U14720 ( .A(n16631), .B(n16632), .Z(n13784) );
  NOR U14721 ( .A(n16633), .B(n16631), .Z(n16632) );
  XOR U14722 ( .A(n16634), .B(n16635), .Z(n13787) );
  NOR U14723 ( .A(n16636), .B(n16634), .Z(n16635) );
  XOR U14724 ( .A(n16637), .B(n16638), .Z(n13790) );
  NOR U14725 ( .A(n16639), .B(n16637), .Z(n16638) );
  XOR U14726 ( .A(n16640), .B(n16641), .Z(n13793) );
  NOR U14727 ( .A(n16642), .B(n16640), .Z(n16641) );
  XOR U14728 ( .A(n16643), .B(n16644), .Z(n13796) );
  NOR U14729 ( .A(n16645), .B(n16643), .Z(n16644) );
  XOR U14730 ( .A(n16646), .B(n16647), .Z(n13799) );
  NOR U14731 ( .A(n16648), .B(n16646), .Z(n16647) );
  XOR U14732 ( .A(n16649), .B(n16650), .Z(n13802) );
  NOR U14733 ( .A(n16651), .B(n16649), .Z(n16650) );
  XOR U14734 ( .A(n16652), .B(n16653), .Z(n13805) );
  NOR U14735 ( .A(n16654), .B(n16652), .Z(n16653) );
  XOR U14736 ( .A(n16655), .B(n16656), .Z(n13808) );
  NOR U14737 ( .A(n16657), .B(n16655), .Z(n16656) );
  XOR U14738 ( .A(n16658), .B(n16659), .Z(n13811) );
  NOR U14739 ( .A(n16660), .B(n16658), .Z(n16659) );
  XOR U14740 ( .A(n16661), .B(n16662), .Z(n13814) );
  NOR U14741 ( .A(n16663), .B(n16661), .Z(n16662) );
  XOR U14742 ( .A(n16664), .B(n16665), .Z(n13817) );
  NOR U14743 ( .A(n16666), .B(n16664), .Z(n16665) );
  XOR U14744 ( .A(n16667), .B(n16668), .Z(n13820) );
  NOR U14745 ( .A(n16669), .B(n16667), .Z(n16668) );
  XOR U14746 ( .A(n16670), .B(n16671), .Z(n13823) );
  NOR U14747 ( .A(n16672), .B(n16670), .Z(n16671) );
  XOR U14748 ( .A(n16673), .B(n16674), .Z(n13826) );
  NOR U14749 ( .A(n16675), .B(n16673), .Z(n16674) );
  XOR U14750 ( .A(n16676), .B(n16677), .Z(n13829) );
  NOR U14751 ( .A(n16678), .B(n16676), .Z(n16677) );
  XOR U14752 ( .A(n16679), .B(n16680), .Z(n13832) );
  NOR U14753 ( .A(n16681), .B(n16679), .Z(n16680) );
  XOR U14754 ( .A(n16682), .B(n16683), .Z(n13835) );
  NOR U14755 ( .A(n16684), .B(n16682), .Z(n16683) );
  XOR U14756 ( .A(n16685), .B(n16686), .Z(n13838) );
  NOR U14757 ( .A(n16687), .B(n16685), .Z(n16686) );
  XOR U14758 ( .A(n16688), .B(n16689), .Z(n13841) );
  NOR U14759 ( .A(n16690), .B(n16688), .Z(n16689) );
  XOR U14760 ( .A(n16691), .B(n16692), .Z(n13844) );
  NOR U14761 ( .A(n16693), .B(n16691), .Z(n16692) );
  XOR U14762 ( .A(n16694), .B(n16695), .Z(n13847) );
  NOR U14763 ( .A(n16696), .B(n16694), .Z(n16695) );
  XOR U14764 ( .A(n16697), .B(n16698), .Z(n13850) );
  NOR U14765 ( .A(n16699), .B(n16697), .Z(n16698) );
  XOR U14766 ( .A(n16700), .B(n16701), .Z(n13853) );
  NOR U14767 ( .A(n16702), .B(n16700), .Z(n16701) );
  XOR U14768 ( .A(n16703), .B(n16704), .Z(n13856) );
  NOR U14769 ( .A(n16705), .B(n16703), .Z(n16704) );
  XOR U14770 ( .A(n16706), .B(n16707), .Z(n13859) );
  NOR U14771 ( .A(n16708), .B(n16706), .Z(n16707) );
  XOR U14772 ( .A(n16709), .B(n16710), .Z(n13862) );
  NOR U14773 ( .A(n16711), .B(n16709), .Z(n16710) );
  XOR U14774 ( .A(n16712), .B(n16713), .Z(n13865) );
  NOR U14775 ( .A(n16714), .B(n16712), .Z(n16713) );
  XOR U14776 ( .A(n16715), .B(n16716), .Z(n13868) );
  NOR U14777 ( .A(n16717), .B(n16715), .Z(n16716) );
  XOR U14778 ( .A(n16718), .B(n16719), .Z(n13871) );
  NOR U14779 ( .A(n16720), .B(n16718), .Z(n16719) );
  XOR U14780 ( .A(n16721), .B(n16722), .Z(n13874) );
  NOR U14781 ( .A(n16723), .B(n16721), .Z(n16722) );
  XOR U14782 ( .A(n16724), .B(n16725), .Z(n13877) );
  NOR U14783 ( .A(n16726), .B(n16724), .Z(n16725) );
  XOR U14784 ( .A(n16727), .B(n16728), .Z(n13880) );
  NOR U14785 ( .A(n16729), .B(n16727), .Z(n16728) );
  XOR U14786 ( .A(n16730), .B(n16731), .Z(n13883) );
  NOR U14787 ( .A(n16732), .B(n16730), .Z(n16731) );
  XOR U14788 ( .A(n16733), .B(n16734), .Z(n13886) );
  NOR U14789 ( .A(n16735), .B(n16733), .Z(n16734) );
  XOR U14790 ( .A(n16736), .B(n16737), .Z(n13889) );
  NOR U14791 ( .A(n16738), .B(n16736), .Z(n16737) );
  XOR U14792 ( .A(n16739), .B(n16740), .Z(n13892) );
  NOR U14793 ( .A(n16741), .B(n16739), .Z(n16740) );
  XOR U14794 ( .A(n16742), .B(n16743), .Z(n13895) );
  NOR U14795 ( .A(n16744), .B(n16742), .Z(n16743) );
  XOR U14796 ( .A(n16745), .B(n16746), .Z(n13898) );
  NOR U14797 ( .A(n16747), .B(n16745), .Z(n16746) );
  XOR U14798 ( .A(n16748), .B(n16749), .Z(n13901) );
  NOR U14799 ( .A(n16750), .B(n16748), .Z(n16749) );
  XOR U14800 ( .A(n16751), .B(n16752), .Z(n13904) );
  NOR U14801 ( .A(n16753), .B(n16751), .Z(n16752) );
  XOR U14802 ( .A(n16754), .B(n16755), .Z(n13907) );
  NOR U14803 ( .A(n16756), .B(n16754), .Z(n16755) );
  XOR U14804 ( .A(n16757), .B(n16758), .Z(n13910) );
  NOR U14805 ( .A(n16759), .B(n16757), .Z(n16758) );
  XOR U14806 ( .A(n16760), .B(n16761), .Z(n13913) );
  NOR U14807 ( .A(n16762), .B(n16760), .Z(n16761) );
  XOR U14808 ( .A(n16763), .B(n16764), .Z(n13916) );
  NOR U14809 ( .A(n16765), .B(n16763), .Z(n16764) );
  XOR U14810 ( .A(n16766), .B(n16767), .Z(n13919) );
  NOR U14811 ( .A(n16768), .B(n16766), .Z(n16767) );
  XOR U14812 ( .A(n16769), .B(n16770), .Z(n13922) );
  NOR U14813 ( .A(n16771), .B(n16769), .Z(n16770) );
  XOR U14814 ( .A(n16772), .B(n16773), .Z(n13925) );
  NOR U14815 ( .A(n16774), .B(n16772), .Z(n16773) );
  XOR U14816 ( .A(n16775), .B(n16776), .Z(n13928) );
  NOR U14817 ( .A(n16777), .B(n16775), .Z(n16776) );
  XOR U14818 ( .A(n16778), .B(n16779), .Z(n13931) );
  NOR U14819 ( .A(n16780), .B(n16778), .Z(n16779) );
  XOR U14820 ( .A(n16781), .B(n16782), .Z(n13934) );
  NOR U14821 ( .A(n16783), .B(n16781), .Z(n16782) );
  XOR U14822 ( .A(n16784), .B(n16785), .Z(n13937) );
  NOR U14823 ( .A(n16786), .B(n16784), .Z(n16785) );
  XOR U14824 ( .A(n16787), .B(n16788), .Z(n13940) );
  NOR U14825 ( .A(n16789), .B(n16787), .Z(n16788) );
  XOR U14826 ( .A(n16790), .B(n16791), .Z(n13943) );
  NOR U14827 ( .A(n16792), .B(n16790), .Z(n16791) );
  XOR U14828 ( .A(n16793), .B(n16794), .Z(n13946) );
  NOR U14829 ( .A(n16795), .B(n16793), .Z(n16794) );
  XOR U14830 ( .A(n16796), .B(n16797), .Z(n13949) );
  NOR U14831 ( .A(n16798), .B(n16796), .Z(n16797) );
  XOR U14832 ( .A(n16799), .B(n16800), .Z(n13952) );
  NOR U14833 ( .A(n16801), .B(n16799), .Z(n16800) );
  XOR U14834 ( .A(n16802), .B(n16803), .Z(n13955) );
  NOR U14835 ( .A(n16804), .B(n16802), .Z(n16803) );
  XOR U14836 ( .A(n16805), .B(n16806), .Z(n13958) );
  NOR U14837 ( .A(n16807), .B(n16805), .Z(n16806) );
  XOR U14838 ( .A(n16808), .B(n16809), .Z(n13961) );
  NOR U14839 ( .A(n16810), .B(n16808), .Z(n16809) );
  XOR U14840 ( .A(n16811), .B(n16812), .Z(n13964) );
  NOR U14841 ( .A(n16813), .B(n16811), .Z(n16812) );
  XOR U14842 ( .A(n16814), .B(n16815), .Z(n13967) );
  NOR U14843 ( .A(n16816), .B(n16814), .Z(n16815) );
  XOR U14844 ( .A(n16817), .B(n16818), .Z(n13970) );
  NOR U14845 ( .A(n16819), .B(n16817), .Z(n16818) );
  XOR U14846 ( .A(n16820), .B(n16821), .Z(n13973) );
  NOR U14847 ( .A(n16822), .B(n16820), .Z(n16821) );
  XOR U14848 ( .A(n16823), .B(n16824), .Z(n13976) );
  NOR U14849 ( .A(n16825), .B(n16823), .Z(n16824) );
  XOR U14850 ( .A(n16826), .B(n16827), .Z(n13979) );
  NOR U14851 ( .A(n16828), .B(n16826), .Z(n16827) );
  XOR U14852 ( .A(n16829), .B(n16830), .Z(n13982) );
  NOR U14853 ( .A(n16831), .B(n16829), .Z(n16830) );
  XOR U14854 ( .A(n16832), .B(n16833), .Z(n13985) );
  NOR U14855 ( .A(n16834), .B(n16832), .Z(n16833) );
  XOR U14856 ( .A(n16835), .B(n16836), .Z(n13988) );
  NOR U14857 ( .A(n16837), .B(n16835), .Z(n16836) );
  XOR U14858 ( .A(n16838), .B(n16839), .Z(n13991) );
  NOR U14859 ( .A(n16840), .B(n16838), .Z(n16839) );
  XOR U14860 ( .A(n16841), .B(n16842), .Z(n13994) );
  NOR U14861 ( .A(n16843), .B(n16841), .Z(n16842) );
  XOR U14862 ( .A(n16844), .B(n16845), .Z(n13997) );
  NOR U14863 ( .A(n16846), .B(n16844), .Z(n16845) );
  XOR U14864 ( .A(n16847), .B(n16848), .Z(n14000) );
  NOR U14865 ( .A(n16849), .B(n16847), .Z(n16848) );
  XOR U14866 ( .A(n16850), .B(n16851), .Z(n14003) );
  NOR U14867 ( .A(n16852), .B(n16850), .Z(n16851) );
  XOR U14868 ( .A(n16853), .B(n16854), .Z(n14006) );
  NOR U14869 ( .A(n16855), .B(n16853), .Z(n16854) );
  XOR U14870 ( .A(n16856), .B(n16857), .Z(n14009) );
  NOR U14871 ( .A(n16858), .B(n16856), .Z(n16857) );
  XOR U14872 ( .A(n16859), .B(n16860), .Z(n14012) );
  NOR U14873 ( .A(n16861), .B(n16859), .Z(n16860) );
  XOR U14874 ( .A(n16862), .B(n16863), .Z(n14015) );
  NOR U14875 ( .A(n16864), .B(n16862), .Z(n16863) );
  XOR U14876 ( .A(n16865), .B(n16866), .Z(n14018) );
  NOR U14877 ( .A(n16867), .B(n16865), .Z(n16866) );
  XOR U14878 ( .A(n16868), .B(n16869), .Z(n14021) );
  NOR U14879 ( .A(n16870), .B(n16868), .Z(n16869) );
  XOR U14880 ( .A(n16871), .B(n16872), .Z(n14024) );
  NOR U14881 ( .A(n16873), .B(n16871), .Z(n16872) );
  XOR U14882 ( .A(n16874), .B(n16875), .Z(n14027) );
  NOR U14883 ( .A(n16876), .B(n16874), .Z(n16875) );
  XOR U14884 ( .A(n16877), .B(n16878), .Z(n14030) );
  NOR U14885 ( .A(n16879), .B(n16877), .Z(n16878) );
  XOR U14886 ( .A(n16880), .B(n16881), .Z(n14033) );
  NOR U14887 ( .A(n16882), .B(n16880), .Z(n16881) );
  XOR U14888 ( .A(n16883), .B(n16884), .Z(n14036) );
  NOR U14889 ( .A(n16885), .B(n16883), .Z(n16884) );
  XOR U14890 ( .A(n16886), .B(n16887), .Z(n14039) );
  NOR U14891 ( .A(n16888), .B(n16886), .Z(n16887) );
  XOR U14892 ( .A(n16889), .B(n16890), .Z(n14042) );
  NOR U14893 ( .A(n16891), .B(n16889), .Z(n16890) );
  XOR U14894 ( .A(n16892), .B(n16893), .Z(n14045) );
  NOR U14895 ( .A(n16894), .B(n16892), .Z(n16893) );
  XOR U14896 ( .A(n16895), .B(n16896), .Z(n14048) );
  NOR U14897 ( .A(n16897), .B(n16895), .Z(n16896) );
  XOR U14898 ( .A(n16898), .B(n16899), .Z(n14051) );
  NOR U14899 ( .A(n16900), .B(n16898), .Z(n16899) );
  XOR U14900 ( .A(n16901), .B(n16902), .Z(n14054) );
  NOR U14901 ( .A(n16903), .B(n16901), .Z(n16902) );
  XOR U14902 ( .A(n16904), .B(n16905), .Z(n14057) );
  NOR U14903 ( .A(n16906), .B(n16904), .Z(n16905) );
  XOR U14904 ( .A(n16907), .B(n16908), .Z(n14060) );
  NOR U14905 ( .A(n16909), .B(n16907), .Z(n16908) );
  XOR U14906 ( .A(n16910), .B(n16911), .Z(n14063) );
  NOR U14907 ( .A(n16912), .B(n16910), .Z(n16911) );
  XOR U14908 ( .A(n16913), .B(n16914), .Z(n14066) );
  NOR U14909 ( .A(n16915), .B(n16913), .Z(n16914) );
  XOR U14910 ( .A(n16916), .B(n16917), .Z(n14069) );
  NOR U14911 ( .A(n16918), .B(n16916), .Z(n16917) );
  XOR U14912 ( .A(n16919), .B(n16920), .Z(n14072) );
  NOR U14913 ( .A(n16921), .B(n16919), .Z(n16920) );
  XOR U14914 ( .A(n16922), .B(n16923), .Z(n14075) );
  NOR U14915 ( .A(n16924), .B(n16922), .Z(n16923) );
  XOR U14916 ( .A(n16925), .B(n16926), .Z(n14078) );
  NOR U14917 ( .A(n16927), .B(n16925), .Z(n16926) );
  XOR U14918 ( .A(n16928), .B(n16929), .Z(n14081) );
  NOR U14919 ( .A(n16930), .B(n16928), .Z(n16929) );
  XOR U14920 ( .A(n16931), .B(n16932), .Z(n14084) );
  NOR U14921 ( .A(n16933), .B(n16931), .Z(n16932) );
  XOR U14922 ( .A(n16934), .B(n16935), .Z(n14087) );
  NOR U14923 ( .A(n16936), .B(n16934), .Z(n16935) );
  XOR U14924 ( .A(n16937), .B(n16938), .Z(n14090) );
  NOR U14925 ( .A(n16939), .B(n16937), .Z(n16938) );
  XOR U14926 ( .A(n16940), .B(n16941), .Z(n14093) );
  NOR U14927 ( .A(n16942), .B(n16940), .Z(n16941) );
  XOR U14928 ( .A(n16943), .B(n16944), .Z(n14096) );
  NOR U14929 ( .A(n16945), .B(n16943), .Z(n16944) );
  XOR U14930 ( .A(n16946), .B(n16947), .Z(n14099) );
  NOR U14931 ( .A(n16948), .B(n16946), .Z(n16947) );
  XOR U14932 ( .A(n16949), .B(n16950), .Z(n14102) );
  NOR U14933 ( .A(n16951), .B(n16949), .Z(n16950) );
  XOR U14934 ( .A(n16952), .B(n16953), .Z(n14105) );
  NOR U14935 ( .A(n16954), .B(n16952), .Z(n16953) );
  XOR U14936 ( .A(n16955), .B(n16956), .Z(n14108) );
  NOR U14937 ( .A(n16957), .B(n16955), .Z(n16956) );
  XOR U14938 ( .A(n16958), .B(n16959), .Z(n14111) );
  NOR U14939 ( .A(n16960), .B(n16958), .Z(n16959) );
  XOR U14940 ( .A(n16961), .B(n16962), .Z(n14114) );
  NOR U14941 ( .A(n16963), .B(n16961), .Z(n16962) );
  XOR U14942 ( .A(n16964), .B(n16965), .Z(n14117) );
  NOR U14943 ( .A(n16966), .B(n16964), .Z(n16965) );
  XOR U14944 ( .A(n16967), .B(n16968), .Z(n14120) );
  NOR U14945 ( .A(n16969), .B(n16967), .Z(n16968) );
  XOR U14946 ( .A(n16970), .B(n16971), .Z(n14123) );
  NOR U14947 ( .A(n16972), .B(n16970), .Z(n16971) );
  XOR U14948 ( .A(n16973), .B(n16974), .Z(n14126) );
  NOR U14949 ( .A(n16975), .B(n16973), .Z(n16974) );
  XOR U14950 ( .A(n16976), .B(n16977), .Z(n14129) );
  NOR U14951 ( .A(n16978), .B(n16976), .Z(n16977) );
  XOR U14952 ( .A(n16979), .B(n16980), .Z(n14132) );
  NOR U14953 ( .A(n16981), .B(n16979), .Z(n16980) );
  XOR U14954 ( .A(n16982), .B(n16983), .Z(n14135) );
  NOR U14955 ( .A(n16984), .B(n16982), .Z(n16983) );
  XOR U14956 ( .A(n16985), .B(n16986), .Z(n14138) );
  NOR U14957 ( .A(n16987), .B(n16985), .Z(n16986) );
  XOR U14958 ( .A(n16988), .B(n16989), .Z(n14141) );
  NOR U14959 ( .A(n16990), .B(n16988), .Z(n16989) );
  XOR U14960 ( .A(n16991), .B(n16992), .Z(n14144) );
  NOR U14961 ( .A(n16993), .B(n16991), .Z(n16992) );
  XOR U14962 ( .A(n16994), .B(n16995), .Z(n14147) );
  NOR U14963 ( .A(n16996), .B(n16994), .Z(n16995) );
  XOR U14964 ( .A(n16997), .B(n16998), .Z(n14150) );
  NOR U14965 ( .A(n16999), .B(n16997), .Z(n16998) );
  XOR U14966 ( .A(n17000), .B(n17001), .Z(n14153) );
  NOR U14967 ( .A(n17002), .B(n17000), .Z(n17001) );
  XOR U14968 ( .A(n17003), .B(n17004), .Z(n14156) );
  NOR U14969 ( .A(n17005), .B(n17003), .Z(n17004) );
  XOR U14970 ( .A(n17006), .B(n17007), .Z(n14159) );
  NOR U14971 ( .A(n17008), .B(n17006), .Z(n17007) );
  XOR U14972 ( .A(n17009), .B(n17010), .Z(n14162) );
  NOR U14973 ( .A(n17011), .B(n17009), .Z(n17010) );
  XOR U14974 ( .A(n17012), .B(n17013), .Z(n14165) );
  NOR U14975 ( .A(n117), .B(n17014), .Z(n17013) );
  XOR U14976 ( .A(n17015), .B(n17016), .Z(n14168) );
  AND U14977 ( .A(n17017), .B(n17018), .Z(n17016) );
  XOR U14978 ( .A(n17015), .B(n119), .Z(n17018) );
  XNOR U14979 ( .A(n15591), .B(n15590), .Z(n119) );
  XNOR U14980 ( .A(n15588), .B(n15587), .Z(n15590) );
  XNOR U14981 ( .A(n15585), .B(n15584), .Z(n15587) );
  XNOR U14982 ( .A(n15582), .B(n15581), .Z(n15584) );
  XNOR U14983 ( .A(n15579), .B(n15578), .Z(n15581) );
  XNOR U14984 ( .A(n15576), .B(n15575), .Z(n15578) );
  XNOR U14985 ( .A(n15573), .B(n15572), .Z(n15575) );
  XNOR U14986 ( .A(n15570), .B(n15569), .Z(n15572) );
  XNOR U14987 ( .A(n15567), .B(n15566), .Z(n15569) );
  XNOR U14988 ( .A(n15564), .B(n15563), .Z(n15566) );
  XNOR U14989 ( .A(n15561), .B(n15560), .Z(n15563) );
  XNOR U14990 ( .A(n15558), .B(n15557), .Z(n15560) );
  XNOR U14991 ( .A(n15555), .B(n15554), .Z(n15557) );
  XNOR U14992 ( .A(n15552), .B(n15551), .Z(n15554) );
  XNOR U14993 ( .A(n15549), .B(n15548), .Z(n15551) );
  XNOR U14994 ( .A(n15546), .B(n15545), .Z(n15548) );
  XNOR U14995 ( .A(n15543), .B(n15542), .Z(n15545) );
  XNOR U14996 ( .A(n15540), .B(n15539), .Z(n15542) );
  XNOR U14997 ( .A(n15537), .B(n15536), .Z(n15539) );
  XNOR U14998 ( .A(n15534), .B(n15533), .Z(n15536) );
  XNOR U14999 ( .A(n15531), .B(n15530), .Z(n15533) );
  XNOR U15000 ( .A(n15528), .B(n15527), .Z(n15530) );
  XNOR U15001 ( .A(n15525), .B(n15524), .Z(n15527) );
  XNOR U15002 ( .A(n15522), .B(n15521), .Z(n15524) );
  XNOR U15003 ( .A(n15519), .B(n15518), .Z(n15521) );
  XNOR U15004 ( .A(n15516), .B(n15515), .Z(n15518) );
  XNOR U15005 ( .A(n15513), .B(n15512), .Z(n15515) );
  XNOR U15006 ( .A(n15510), .B(n15509), .Z(n15512) );
  XNOR U15007 ( .A(n15507), .B(n15506), .Z(n15509) );
  XNOR U15008 ( .A(n15504), .B(n15503), .Z(n15506) );
  XNOR U15009 ( .A(n15501), .B(n15500), .Z(n15503) );
  XNOR U15010 ( .A(n15498), .B(n15497), .Z(n15500) );
  XNOR U15011 ( .A(n15495), .B(n15494), .Z(n15497) );
  XNOR U15012 ( .A(n15492), .B(n15491), .Z(n15494) );
  XNOR U15013 ( .A(n15489), .B(n15488), .Z(n15491) );
  XNOR U15014 ( .A(n15486), .B(n15485), .Z(n15488) );
  XNOR U15015 ( .A(n15483), .B(n15482), .Z(n15485) );
  XNOR U15016 ( .A(n15480), .B(n15479), .Z(n15482) );
  XNOR U15017 ( .A(n15477), .B(n15476), .Z(n15479) );
  XNOR U15018 ( .A(n15474), .B(n15473), .Z(n15476) );
  XNOR U15019 ( .A(n15471), .B(n15470), .Z(n15473) );
  XNOR U15020 ( .A(n15468), .B(n15467), .Z(n15470) );
  XNOR U15021 ( .A(n15465), .B(n15464), .Z(n15467) );
  XNOR U15022 ( .A(n15462), .B(n15461), .Z(n15464) );
  XNOR U15023 ( .A(n15459), .B(n15458), .Z(n15461) );
  XNOR U15024 ( .A(n15456), .B(n15455), .Z(n15458) );
  XNOR U15025 ( .A(n15453), .B(n15452), .Z(n15455) );
  XNOR U15026 ( .A(n15450), .B(n15449), .Z(n15452) );
  XNOR U15027 ( .A(n15447), .B(n15446), .Z(n15449) );
  XNOR U15028 ( .A(n15444), .B(n15443), .Z(n15446) );
  XNOR U15029 ( .A(n15441), .B(n15440), .Z(n15443) );
  XNOR U15030 ( .A(n15438), .B(n15437), .Z(n15440) );
  XNOR U15031 ( .A(n15435), .B(n15434), .Z(n15437) );
  XNOR U15032 ( .A(n15432), .B(n15431), .Z(n15434) );
  XNOR U15033 ( .A(n15429), .B(n15428), .Z(n15431) );
  XNOR U15034 ( .A(n15426), .B(n15425), .Z(n15428) );
  XNOR U15035 ( .A(n15423), .B(n15422), .Z(n15425) );
  XNOR U15036 ( .A(n15420), .B(n15419), .Z(n15422) );
  XNOR U15037 ( .A(n15417), .B(n15416), .Z(n15419) );
  XNOR U15038 ( .A(n15414), .B(n15413), .Z(n15416) );
  XNOR U15039 ( .A(n15411), .B(n15410), .Z(n15413) );
  XNOR U15040 ( .A(n15408), .B(n15407), .Z(n15410) );
  XNOR U15041 ( .A(n15405), .B(n15404), .Z(n15407) );
  XNOR U15042 ( .A(n15402), .B(n15401), .Z(n15404) );
  XNOR U15043 ( .A(n15399), .B(n15398), .Z(n15401) );
  XNOR U15044 ( .A(n15396), .B(n15395), .Z(n15398) );
  XNOR U15045 ( .A(n15393), .B(n15392), .Z(n15395) );
  XNOR U15046 ( .A(n15390), .B(n15389), .Z(n15392) );
  XNOR U15047 ( .A(n15387), .B(n15386), .Z(n15389) );
  XNOR U15048 ( .A(n15384), .B(n15383), .Z(n15386) );
  XNOR U15049 ( .A(n15381), .B(n15380), .Z(n15383) );
  XNOR U15050 ( .A(n15378), .B(n15377), .Z(n15380) );
  XNOR U15051 ( .A(n15375), .B(n15374), .Z(n15377) );
  XNOR U15052 ( .A(n15372), .B(n15371), .Z(n15374) );
  XNOR U15053 ( .A(n15369), .B(n15368), .Z(n15371) );
  XNOR U15054 ( .A(n15366), .B(n15365), .Z(n15368) );
  XNOR U15055 ( .A(n15363), .B(n15362), .Z(n15365) );
  XNOR U15056 ( .A(n15360), .B(n15359), .Z(n15362) );
  XNOR U15057 ( .A(n15357), .B(n15356), .Z(n15359) );
  XNOR U15058 ( .A(n15354), .B(n15353), .Z(n15356) );
  XNOR U15059 ( .A(n15351), .B(n15350), .Z(n15353) );
  XNOR U15060 ( .A(n15348), .B(n15347), .Z(n15350) );
  XNOR U15061 ( .A(n15345), .B(n15344), .Z(n15347) );
  XNOR U15062 ( .A(n15342), .B(n15341), .Z(n15344) );
  XNOR U15063 ( .A(n15339), .B(n15338), .Z(n15341) );
  XNOR U15064 ( .A(n15336), .B(n15335), .Z(n15338) );
  XNOR U15065 ( .A(n15333), .B(n15332), .Z(n15335) );
  XNOR U15066 ( .A(n15330), .B(n15329), .Z(n15332) );
  XNOR U15067 ( .A(n15327), .B(n15326), .Z(n15329) );
  XNOR U15068 ( .A(n15324), .B(n15323), .Z(n15326) );
  XNOR U15069 ( .A(n15321), .B(n15320), .Z(n15323) );
  XNOR U15070 ( .A(n15318), .B(n15317), .Z(n15320) );
  XNOR U15071 ( .A(n15315), .B(n15314), .Z(n15317) );
  XNOR U15072 ( .A(n15312), .B(n15311), .Z(n15314) );
  XNOR U15073 ( .A(n15309), .B(n15308), .Z(n15311) );
  XNOR U15074 ( .A(n15306), .B(n15305), .Z(n15308) );
  XNOR U15075 ( .A(n15303), .B(n15302), .Z(n15305) );
  XNOR U15076 ( .A(n15300), .B(n15299), .Z(n15302) );
  XNOR U15077 ( .A(n15297), .B(n15296), .Z(n15299) );
  XNOR U15078 ( .A(n15294), .B(n15293), .Z(n15296) );
  XNOR U15079 ( .A(n15291), .B(n15290), .Z(n15293) );
  XNOR U15080 ( .A(n15288), .B(n15287), .Z(n15290) );
  XNOR U15081 ( .A(n15285), .B(n15284), .Z(n15287) );
  XNOR U15082 ( .A(n15282), .B(n15281), .Z(n15284) );
  XNOR U15083 ( .A(n15279), .B(n15278), .Z(n15281) );
  XNOR U15084 ( .A(n15276), .B(n15275), .Z(n15278) );
  XNOR U15085 ( .A(n15273), .B(n15272), .Z(n15275) );
  XNOR U15086 ( .A(n15270), .B(n15269), .Z(n15272) );
  XNOR U15087 ( .A(n15267), .B(n15266), .Z(n15269) );
  XNOR U15088 ( .A(n15264), .B(n15263), .Z(n15266) );
  XNOR U15089 ( .A(n15261), .B(n15260), .Z(n15263) );
  XNOR U15090 ( .A(n15258), .B(n15257), .Z(n15260) );
  XNOR U15091 ( .A(n15255), .B(n15254), .Z(n15257) );
  XNOR U15092 ( .A(n15252), .B(n15251), .Z(n15254) );
  XNOR U15093 ( .A(n15249), .B(n15248), .Z(n15251) );
  XNOR U15094 ( .A(n15246), .B(n15245), .Z(n15248) );
  XNOR U15095 ( .A(n15243), .B(n15242), .Z(n15245) );
  XNOR U15096 ( .A(n15240), .B(n15239), .Z(n15242) );
  XNOR U15097 ( .A(n15237), .B(n15236), .Z(n15239) );
  XNOR U15098 ( .A(n15234), .B(n15233), .Z(n15236) );
  XNOR U15099 ( .A(n15231), .B(n15230), .Z(n15233) );
  XNOR U15100 ( .A(n15228), .B(n15227), .Z(n15230) );
  XNOR U15101 ( .A(n15225), .B(n15224), .Z(n15227) );
  XNOR U15102 ( .A(n15222), .B(n15221), .Z(n15224) );
  XNOR U15103 ( .A(n15219), .B(n15218), .Z(n15221) );
  XNOR U15104 ( .A(n15216), .B(n15215), .Z(n15218) );
  XNOR U15105 ( .A(n15213), .B(n15212), .Z(n15215) );
  XNOR U15106 ( .A(n15210), .B(n15209), .Z(n15212) );
  XNOR U15107 ( .A(n15207), .B(n15206), .Z(n15209) );
  XNOR U15108 ( .A(n15204), .B(n15203), .Z(n15206) );
  XNOR U15109 ( .A(n15201), .B(n15200), .Z(n15203) );
  XNOR U15110 ( .A(n15198), .B(n15197), .Z(n15200) );
  XNOR U15111 ( .A(n15195), .B(n15194), .Z(n15197) );
  XNOR U15112 ( .A(n15192), .B(n15191), .Z(n15194) );
  XNOR U15113 ( .A(n15189), .B(n15188), .Z(n15191) );
  XNOR U15114 ( .A(n15186), .B(n15185), .Z(n15188) );
  XNOR U15115 ( .A(n15183), .B(n15182), .Z(n15185) );
  XNOR U15116 ( .A(n15180), .B(n15179), .Z(n15182) );
  XNOR U15117 ( .A(n15177), .B(n15176), .Z(n15179) );
  XNOR U15118 ( .A(n15174), .B(n15173), .Z(n15176) );
  XNOR U15119 ( .A(n15171), .B(n15170), .Z(n15173) );
  XNOR U15120 ( .A(n15168), .B(n15167), .Z(n15170) );
  XNOR U15121 ( .A(n15165), .B(n15164), .Z(n15167) );
  XNOR U15122 ( .A(n15162), .B(n15161), .Z(n15164) );
  XNOR U15123 ( .A(n15159), .B(n15158), .Z(n15161) );
  XNOR U15124 ( .A(n15156), .B(n15155), .Z(n15158) );
  XNOR U15125 ( .A(n15153), .B(n15152), .Z(n15155) );
  XNOR U15126 ( .A(n15150), .B(n15149), .Z(n15152) );
  XNOR U15127 ( .A(n15147), .B(n15146), .Z(n15149) );
  XNOR U15128 ( .A(n15144), .B(n15143), .Z(n15146) );
  XNOR U15129 ( .A(n15141), .B(n15140), .Z(n15143) );
  XNOR U15130 ( .A(n15138), .B(n15137), .Z(n15140) );
  XNOR U15131 ( .A(n15135), .B(n15134), .Z(n15137) );
  XNOR U15132 ( .A(n15132), .B(n15131), .Z(n15134) );
  XNOR U15133 ( .A(n15129), .B(n15128), .Z(n15131) );
  XNOR U15134 ( .A(n15126), .B(n15125), .Z(n15128) );
  XNOR U15135 ( .A(n15123), .B(n15122), .Z(n15125) );
  XNOR U15136 ( .A(n15120), .B(n15119), .Z(n15122) );
  XNOR U15137 ( .A(n15117), .B(n15116), .Z(n15119) );
  XNOR U15138 ( .A(n15114), .B(n15113), .Z(n15116) );
  XNOR U15139 ( .A(n15111), .B(n15110), .Z(n15113) );
  XNOR U15140 ( .A(n15108), .B(n15107), .Z(n15110) );
  XNOR U15141 ( .A(n15105), .B(n15104), .Z(n15107) );
  XNOR U15142 ( .A(n15102), .B(n15101), .Z(n15104) );
  XNOR U15143 ( .A(n15099), .B(n15098), .Z(n15101) );
  XNOR U15144 ( .A(n15096), .B(n15095), .Z(n15098) );
  XNOR U15145 ( .A(n15093), .B(n15092), .Z(n15095) );
  XNOR U15146 ( .A(n15090), .B(n15089), .Z(n15092) );
  XNOR U15147 ( .A(n15087), .B(n15086), .Z(n15089) );
  XNOR U15148 ( .A(n15084), .B(n15083), .Z(n15086) );
  XNOR U15149 ( .A(n15081), .B(n15080), .Z(n15083) );
  XNOR U15150 ( .A(n15078), .B(n15077), .Z(n15080) );
  XNOR U15151 ( .A(n15075), .B(n15074), .Z(n15077) );
  XNOR U15152 ( .A(n15072), .B(n15071), .Z(n15074) );
  XNOR U15153 ( .A(n15069), .B(n15068), .Z(n15071) );
  XNOR U15154 ( .A(n15066), .B(n15065), .Z(n15068) );
  XNOR U15155 ( .A(n15063), .B(n15062), .Z(n15065) );
  XNOR U15156 ( .A(n15060), .B(n15059), .Z(n15062) );
  XNOR U15157 ( .A(n15057), .B(n15056), .Z(n15059) );
  XNOR U15158 ( .A(n15054), .B(n15053), .Z(n15056) );
  XNOR U15159 ( .A(n15051), .B(n15050), .Z(n15053) );
  XNOR U15160 ( .A(n15048), .B(n15047), .Z(n15050) );
  XNOR U15161 ( .A(n15045), .B(n15044), .Z(n15047) );
  XNOR U15162 ( .A(n15042), .B(n15041), .Z(n15044) );
  XNOR U15163 ( .A(n15039), .B(n15038), .Z(n15041) );
  XNOR U15164 ( .A(n15036), .B(n15035), .Z(n15038) );
  XNOR U15165 ( .A(n15033), .B(n15032), .Z(n15035) );
  XNOR U15166 ( .A(n15030), .B(n15029), .Z(n15032) );
  XNOR U15167 ( .A(n15027), .B(n15026), .Z(n15029) );
  XNOR U15168 ( .A(n15024), .B(n15023), .Z(n15026) );
  XNOR U15169 ( .A(n15021), .B(n15020), .Z(n15023) );
  XNOR U15170 ( .A(n15018), .B(n15017), .Z(n15020) );
  XNOR U15171 ( .A(n15015), .B(n15014), .Z(n15017) );
  XNOR U15172 ( .A(n15012), .B(n15011), .Z(n15014) );
  XNOR U15173 ( .A(n15009), .B(n15008), .Z(n15011) );
  XNOR U15174 ( .A(n15006), .B(n15005), .Z(n15008) );
  XNOR U15175 ( .A(n15003), .B(n15002), .Z(n15005) );
  XNOR U15176 ( .A(n15000), .B(n14999), .Z(n15002) );
  XNOR U15177 ( .A(n14997), .B(n14996), .Z(n14999) );
  XNOR U15178 ( .A(n14994), .B(n14993), .Z(n14996) );
  XNOR U15179 ( .A(n14991), .B(n14990), .Z(n14993) );
  XNOR U15180 ( .A(n14988), .B(n14987), .Z(n14990) );
  XNOR U15181 ( .A(n14985), .B(n14984), .Z(n14987) );
  XNOR U15182 ( .A(n14982), .B(n14981), .Z(n14984) );
  XNOR U15183 ( .A(n14979), .B(n14978), .Z(n14981) );
  XNOR U15184 ( .A(n14976), .B(n14975), .Z(n14978) );
  XNOR U15185 ( .A(n14973), .B(n14972), .Z(n14975) );
  XNOR U15186 ( .A(n14970), .B(n14969), .Z(n14972) );
  XNOR U15187 ( .A(n14967), .B(n14966), .Z(n14969) );
  XNOR U15188 ( .A(n14964), .B(n14963), .Z(n14966) );
  XNOR U15189 ( .A(n14961), .B(n14960), .Z(n14963) );
  XNOR U15190 ( .A(n14958), .B(n14957), .Z(n14960) );
  XNOR U15191 ( .A(n14955), .B(n14954), .Z(n14957) );
  XNOR U15192 ( .A(n14952), .B(n14951), .Z(n14954) );
  XNOR U15193 ( .A(n14949), .B(n14948), .Z(n14951) );
  XNOR U15194 ( .A(n14946), .B(n14945), .Z(n14948) );
  XNOR U15195 ( .A(n14943), .B(n14942), .Z(n14945) );
  XNOR U15196 ( .A(n14940), .B(n14939), .Z(n14942) );
  XNOR U15197 ( .A(n14937), .B(n14936), .Z(n14939) );
  XNOR U15198 ( .A(n14934), .B(n14933), .Z(n14936) );
  XNOR U15199 ( .A(n14931), .B(n14930), .Z(n14933) );
  XNOR U15200 ( .A(n14928), .B(n14927), .Z(n14930) );
  XNOR U15201 ( .A(n14925), .B(n14924), .Z(n14927) );
  XNOR U15202 ( .A(n14922), .B(n14921), .Z(n14924) );
  XNOR U15203 ( .A(n14919), .B(n14918), .Z(n14921) );
  XNOR U15204 ( .A(n14916), .B(n14915), .Z(n14918) );
  XNOR U15205 ( .A(n14913), .B(n14912), .Z(n14915) );
  XNOR U15206 ( .A(n14910), .B(n14909), .Z(n14912) );
  XNOR U15207 ( .A(n14907), .B(n14906), .Z(n14909) );
  XNOR U15208 ( .A(n14904), .B(n14903), .Z(n14906) );
  XNOR U15209 ( .A(n14901), .B(n14900), .Z(n14903) );
  XNOR U15210 ( .A(n14898), .B(n14897), .Z(n14900) );
  XNOR U15211 ( .A(n14895), .B(n14894), .Z(n14897) );
  XNOR U15212 ( .A(n14892), .B(n14891), .Z(n14894) );
  XNOR U15213 ( .A(n14889), .B(n14888), .Z(n14891) );
  XNOR U15214 ( .A(n14886), .B(n14885), .Z(n14888) );
  XNOR U15215 ( .A(n14883), .B(n14882), .Z(n14885) );
  XNOR U15216 ( .A(n14880), .B(n14879), .Z(n14882) );
  XNOR U15217 ( .A(n14877), .B(n14876), .Z(n14879) );
  XNOR U15218 ( .A(n14874), .B(n14873), .Z(n14876) );
  XNOR U15219 ( .A(n14871), .B(n14870), .Z(n14873) );
  XNOR U15220 ( .A(n14868), .B(n14867), .Z(n14870) );
  XNOR U15221 ( .A(n14865), .B(n14864), .Z(n14867) );
  XNOR U15222 ( .A(n14862), .B(n14861), .Z(n14864) );
  XNOR U15223 ( .A(n14859), .B(n14858), .Z(n14861) );
  XNOR U15224 ( .A(n14856), .B(n14855), .Z(n14858) );
  XNOR U15225 ( .A(n14853), .B(n14852), .Z(n14855) );
  XNOR U15226 ( .A(n14850), .B(n14849), .Z(n14852) );
  XNOR U15227 ( .A(n14847), .B(n14846), .Z(n14849) );
  XNOR U15228 ( .A(n14844), .B(n14843), .Z(n14846) );
  XNOR U15229 ( .A(n14841), .B(n14840), .Z(n14843) );
  XNOR U15230 ( .A(n14838), .B(n14837), .Z(n14840) );
  XNOR U15231 ( .A(n14835), .B(n14834), .Z(n14837) );
  XNOR U15232 ( .A(n14832), .B(n14831), .Z(n14834) );
  XNOR U15233 ( .A(n14829), .B(n14828), .Z(n14831) );
  XNOR U15234 ( .A(n14826), .B(n14825), .Z(n14828) );
  XNOR U15235 ( .A(n14823), .B(n14822), .Z(n14825) );
  XNOR U15236 ( .A(n14820), .B(n14819), .Z(n14822) );
  XNOR U15237 ( .A(n14817), .B(n14816), .Z(n14819) );
  XNOR U15238 ( .A(n14814), .B(n14813), .Z(n14816) );
  XNOR U15239 ( .A(n14811), .B(n14810), .Z(n14813) );
  XNOR U15240 ( .A(n14808), .B(n14807), .Z(n14810) );
  XNOR U15241 ( .A(n14805), .B(n14804), .Z(n14807) );
  XNOR U15242 ( .A(n14802), .B(n14801), .Z(n14804) );
  XNOR U15243 ( .A(n14799), .B(n14798), .Z(n14801) );
  XNOR U15244 ( .A(n14796), .B(n14795), .Z(n14798) );
  XNOR U15245 ( .A(n14793), .B(n14792), .Z(n14795) );
  XNOR U15246 ( .A(n14790), .B(n14789), .Z(n14792) );
  XNOR U15247 ( .A(n14787), .B(n14786), .Z(n14789) );
  XNOR U15248 ( .A(n14784), .B(n14783), .Z(n14786) );
  XNOR U15249 ( .A(n14781), .B(n14780), .Z(n14783) );
  XNOR U15250 ( .A(n14778), .B(n14777), .Z(n14780) );
  XNOR U15251 ( .A(n14775), .B(n14774), .Z(n14777) );
  XNOR U15252 ( .A(n14772), .B(n14771), .Z(n14774) );
  XNOR U15253 ( .A(n14769), .B(n14768), .Z(n14771) );
  XNOR U15254 ( .A(n14766), .B(n14765), .Z(n14768) );
  XNOR U15255 ( .A(n14763), .B(n14762), .Z(n14765) );
  XNOR U15256 ( .A(n14760), .B(n14759), .Z(n14762) );
  XNOR U15257 ( .A(n14757), .B(n14756), .Z(n14759) );
  XNOR U15258 ( .A(n14754), .B(n14753), .Z(n14756) );
  XNOR U15259 ( .A(n14751), .B(n14750), .Z(n14753) );
  XNOR U15260 ( .A(n14748), .B(n14747), .Z(n14750) );
  XNOR U15261 ( .A(n14745), .B(n14744), .Z(n14747) );
  XNOR U15262 ( .A(n14742), .B(n14741), .Z(n14744) );
  XNOR U15263 ( .A(n14739), .B(n14738), .Z(n14741) );
  XNOR U15264 ( .A(n14736), .B(n14735), .Z(n14738) );
  XNOR U15265 ( .A(n14733), .B(n14732), .Z(n14735) );
  XNOR U15266 ( .A(n14730), .B(n14729), .Z(n14732) );
  XNOR U15267 ( .A(n14727), .B(n14726), .Z(n14729) );
  XNOR U15268 ( .A(n14724), .B(n14723), .Z(n14726) );
  XNOR U15269 ( .A(n14721), .B(n14720), .Z(n14723) );
  XNOR U15270 ( .A(n14718), .B(n14717), .Z(n14720) );
  XNOR U15271 ( .A(n14715), .B(n14714), .Z(n14717) );
  XNOR U15272 ( .A(n14712), .B(n14711), .Z(n14714) );
  XNOR U15273 ( .A(n14709), .B(n14708), .Z(n14711) );
  XNOR U15274 ( .A(n14706), .B(n14705), .Z(n14708) );
  XNOR U15275 ( .A(n14703), .B(n14702), .Z(n14705) );
  XNOR U15276 ( .A(n14700), .B(n14699), .Z(n14702) );
  XNOR U15277 ( .A(n14697), .B(n14696), .Z(n14699) );
  XNOR U15278 ( .A(n14694), .B(n14693), .Z(n14696) );
  XNOR U15279 ( .A(n14691), .B(n14690), .Z(n14693) );
  XNOR U15280 ( .A(n14688), .B(n14687), .Z(n14690) );
  XNOR U15281 ( .A(n14685), .B(n14684), .Z(n14687) );
  XNOR U15282 ( .A(n14682), .B(n14681), .Z(n14684) );
  XNOR U15283 ( .A(n14679), .B(n14678), .Z(n14681) );
  XNOR U15284 ( .A(n14676), .B(n14675), .Z(n14678) );
  XNOR U15285 ( .A(n14673), .B(n14672), .Z(n14675) );
  XNOR U15286 ( .A(n14670), .B(n14669), .Z(n14672) );
  XNOR U15287 ( .A(n14667), .B(n14666), .Z(n14669) );
  XNOR U15288 ( .A(n14664), .B(n14663), .Z(n14666) );
  XNOR U15289 ( .A(n14661), .B(n14660), .Z(n14663) );
  XNOR U15290 ( .A(n14658), .B(n14657), .Z(n14660) );
  XNOR U15291 ( .A(n14655), .B(n14654), .Z(n14657) );
  XNOR U15292 ( .A(n14652), .B(n14651), .Z(n14654) );
  XNOR U15293 ( .A(n14649), .B(n14648), .Z(n14651) );
  XNOR U15294 ( .A(n14646), .B(n14645), .Z(n14648) );
  XNOR U15295 ( .A(n14643), .B(n14642), .Z(n14645) );
  XNOR U15296 ( .A(n14640), .B(n14639), .Z(n14642) );
  XNOR U15297 ( .A(n14637), .B(n14636), .Z(n14639) );
  XNOR U15298 ( .A(n14634), .B(n14633), .Z(n14636) );
  XNOR U15299 ( .A(n14631), .B(n14630), .Z(n14633) );
  XNOR U15300 ( .A(n14628), .B(n14627), .Z(n14630) );
  XNOR U15301 ( .A(n14625), .B(n14624), .Z(n14627) );
  XNOR U15302 ( .A(n14622), .B(n14621), .Z(n14624) );
  XNOR U15303 ( .A(n14619), .B(n14618), .Z(n14621) );
  XNOR U15304 ( .A(n14616), .B(n14615), .Z(n14618) );
  XNOR U15305 ( .A(n14613), .B(n14612), .Z(n14615) );
  XNOR U15306 ( .A(n14610), .B(n14609), .Z(n14612) );
  XNOR U15307 ( .A(n14607), .B(n14606), .Z(n14609) );
  XNOR U15308 ( .A(n14604), .B(n14603), .Z(n14606) );
  XNOR U15309 ( .A(n14601), .B(n14600), .Z(n14603) );
  XNOR U15310 ( .A(n14598), .B(n14597), .Z(n14600) );
  XNOR U15311 ( .A(n14595), .B(n14594), .Z(n14597) );
  XNOR U15312 ( .A(n14592), .B(n14591), .Z(n14594) );
  XNOR U15313 ( .A(n14589), .B(n14588), .Z(n14591) );
  XNOR U15314 ( .A(n14586), .B(n14585), .Z(n14588) );
  XNOR U15315 ( .A(n14583), .B(n14582), .Z(n14585) );
  XNOR U15316 ( .A(n14580), .B(n14579), .Z(n14582) );
  XNOR U15317 ( .A(n14577), .B(n14576), .Z(n14579) );
  XNOR U15318 ( .A(n14574), .B(n14573), .Z(n14576) );
  XNOR U15319 ( .A(n14571), .B(n14570), .Z(n14573) );
  XNOR U15320 ( .A(n14568), .B(n14567), .Z(n14570) );
  XNOR U15321 ( .A(n14565), .B(n14564), .Z(n14567) );
  XNOR U15322 ( .A(n14562), .B(n14561), .Z(n14564) );
  XNOR U15323 ( .A(n14559), .B(n14558), .Z(n14561) );
  XNOR U15324 ( .A(n14556), .B(n14555), .Z(n14558) );
  XNOR U15325 ( .A(n14553), .B(n14552), .Z(n14555) );
  XNOR U15326 ( .A(n14550), .B(n14549), .Z(n14552) );
  XNOR U15327 ( .A(n14547), .B(n14546), .Z(n14549) );
  XNOR U15328 ( .A(n14544), .B(n14543), .Z(n14546) );
  XNOR U15329 ( .A(n14541), .B(n14540), .Z(n14543) );
  XNOR U15330 ( .A(n14538), .B(n14537), .Z(n14540) );
  XNOR U15331 ( .A(n14535), .B(n14534), .Z(n14537) );
  XNOR U15332 ( .A(n14532), .B(n14531), .Z(n14534) );
  XNOR U15333 ( .A(n14529), .B(n14528), .Z(n14531) );
  XNOR U15334 ( .A(n14526), .B(n14525), .Z(n14528) );
  XNOR U15335 ( .A(n14523), .B(n14522), .Z(n14525) );
  XNOR U15336 ( .A(n14520), .B(n14519), .Z(n14522) );
  XNOR U15337 ( .A(n14517), .B(n14516), .Z(n14519) );
  XNOR U15338 ( .A(n14514), .B(n14513), .Z(n14516) );
  XNOR U15339 ( .A(n14511), .B(n14510), .Z(n14513) );
  XNOR U15340 ( .A(n14508), .B(n14507), .Z(n14510) );
  XNOR U15341 ( .A(n14505), .B(n14504), .Z(n14507) );
  XNOR U15342 ( .A(n14502), .B(n14501), .Z(n14504) );
  XNOR U15343 ( .A(n14499), .B(n14498), .Z(n14501) );
  XNOR U15344 ( .A(n14496), .B(n14495), .Z(n14498) );
  XNOR U15345 ( .A(n14493), .B(n14492), .Z(n14495) );
  XNOR U15346 ( .A(n14490), .B(n14489), .Z(n14492) );
  XNOR U15347 ( .A(n14487), .B(n14486), .Z(n14489) );
  XNOR U15348 ( .A(n14484), .B(n14483), .Z(n14486) );
  XNOR U15349 ( .A(n14481), .B(n14480), .Z(n14483) );
  XNOR U15350 ( .A(n14478), .B(n14477), .Z(n14480) );
  XNOR U15351 ( .A(n14475), .B(n14474), .Z(n14477) );
  XNOR U15352 ( .A(n14472), .B(n14471), .Z(n14474) );
  XNOR U15353 ( .A(n14469), .B(n14468), .Z(n14471) );
  XNOR U15354 ( .A(n14466), .B(n14465), .Z(n14468) );
  XNOR U15355 ( .A(n14463), .B(n14462), .Z(n14465) );
  XNOR U15356 ( .A(n14460), .B(n14459), .Z(n14462) );
  XNOR U15357 ( .A(n14457), .B(n14456), .Z(n14459) );
  XNOR U15358 ( .A(n14454), .B(n14453), .Z(n14456) );
  XNOR U15359 ( .A(n14451), .B(n14450), .Z(n14453) );
  XNOR U15360 ( .A(n14448), .B(n14447), .Z(n14450) );
  XNOR U15361 ( .A(n14445), .B(n14444), .Z(n14447) );
  XNOR U15362 ( .A(n14442), .B(n14441), .Z(n14444) );
  XNOR U15363 ( .A(n14439), .B(n14438), .Z(n14441) );
  XOR U15364 ( .A(n14436), .B(n14435), .Z(n14438) );
  XOR U15365 ( .A(n14433), .B(n14432), .Z(n14435) );
  XOR U15366 ( .A(n14429), .B(n14430), .Z(n14432) );
  AND U15367 ( .A(n17019), .B(n17020), .Z(n14430) );
  XOR U15368 ( .A(n14426), .B(n14427), .Z(n14429) );
  AND U15369 ( .A(n17021), .B(n17022), .Z(n14427) );
  XOR U15370 ( .A(n14423), .B(n14424), .Z(n14426) );
  AND U15371 ( .A(n17023), .B(n17024), .Z(n14424) );
  XNOR U15372 ( .A(n14172), .B(n14421), .Z(n14423) );
  AND U15373 ( .A(n17025), .B(n17026), .Z(n14421) );
  XOR U15374 ( .A(n14174), .B(n14173), .Z(n14172) );
  AND U15375 ( .A(n17027), .B(n17028), .Z(n14173) );
  XOR U15376 ( .A(n14176), .B(n14175), .Z(n14174) );
  AND U15377 ( .A(n17029), .B(n17030), .Z(n14175) );
  XOR U15378 ( .A(n14178), .B(n14177), .Z(n14176) );
  AND U15379 ( .A(n17031), .B(n17032), .Z(n14177) );
  XOR U15380 ( .A(n14180), .B(n14179), .Z(n14178) );
  AND U15381 ( .A(n17033), .B(n17034), .Z(n14179) );
  XOR U15382 ( .A(n14182), .B(n14181), .Z(n14180) );
  AND U15383 ( .A(n17035), .B(n17036), .Z(n14181) );
  XOR U15384 ( .A(n14184), .B(n14183), .Z(n14182) );
  AND U15385 ( .A(n17037), .B(n17038), .Z(n14183) );
  XOR U15386 ( .A(n14186), .B(n14185), .Z(n14184) );
  AND U15387 ( .A(n17039), .B(n17040), .Z(n14185) );
  XOR U15388 ( .A(n14188), .B(n14187), .Z(n14186) );
  AND U15389 ( .A(n17041), .B(n17042), .Z(n14187) );
  XOR U15390 ( .A(n14190), .B(n14189), .Z(n14188) );
  AND U15391 ( .A(n17043), .B(n17044), .Z(n14189) );
  XOR U15392 ( .A(n14192), .B(n14191), .Z(n14190) );
  AND U15393 ( .A(n17045), .B(n17046), .Z(n14191) );
  XOR U15394 ( .A(n14194), .B(n14193), .Z(n14192) );
  AND U15395 ( .A(n17047), .B(n17048), .Z(n14193) );
  XOR U15396 ( .A(n14196), .B(n14195), .Z(n14194) );
  AND U15397 ( .A(n17049), .B(n17050), .Z(n14195) );
  XOR U15398 ( .A(n14198), .B(n14197), .Z(n14196) );
  AND U15399 ( .A(n17051), .B(n17052), .Z(n14197) );
  XOR U15400 ( .A(n14200), .B(n14199), .Z(n14198) );
  AND U15401 ( .A(n17053), .B(n17054), .Z(n14199) );
  XOR U15402 ( .A(n14202), .B(n14201), .Z(n14200) );
  AND U15403 ( .A(n17055), .B(n17056), .Z(n14201) );
  XOR U15404 ( .A(n14204), .B(n14203), .Z(n14202) );
  AND U15405 ( .A(n17057), .B(n17058), .Z(n14203) );
  XOR U15406 ( .A(n14206), .B(n14205), .Z(n14204) );
  AND U15407 ( .A(n17059), .B(n17060), .Z(n14205) );
  XOR U15408 ( .A(n14208), .B(n14207), .Z(n14206) );
  AND U15409 ( .A(n17061), .B(n17062), .Z(n14207) );
  XOR U15410 ( .A(n14210), .B(n14209), .Z(n14208) );
  AND U15411 ( .A(n17063), .B(n17064), .Z(n14209) );
  XOR U15412 ( .A(n14212), .B(n14211), .Z(n14210) );
  AND U15413 ( .A(n17065), .B(n17066), .Z(n14211) );
  XOR U15414 ( .A(n14214), .B(n14213), .Z(n14212) );
  AND U15415 ( .A(n17067), .B(n17068), .Z(n14213) );
  XOR U15416 ( .A(n14216), .B(n14215), .Z(n14214) );
  AND U15417 ( .A(n17069), .B(n17070), .Z(n14215) );
  XOR U15418 ( .A(n14218), .B(n14217), .Z(n14216) );
  AND U15419 ( .A(n17071), .B(n17072), .Z(n14217) );
  XOR U15420 ( .A(n14220), .B(n14219), .Z(n14218) );
  AND U15421 ( .A(n17073), .B(n17074), .Z(n14219) );
  XOR U15422 ( .A(n14222), .B(n14221), .Z(n14220) );
  AND U15423 ( .A(n17075), .B(n17076), .Z(n14221) );
  XOR U15424 ( .A(n14224), .B(n14223), .Z(n14222) );
  AND U15425 ( .A(n17077), .B(n17078), .Z(n14223) );
  XOR U15426 ( .A(n14226), .B(n14225), .Z(n14224) );
  AND U15427 ( .A(n17079), .B(n17080), .Z(n14225) );
  XOR U15428 ( .A(n14228), .B(n14227), .Z(n14226) );
  AND U15429 ( .A(n17081), .B(n17082), .Z(n14227) );
  XOR U15430 ( .A(n14230), .B(n14229), .Z(n14228) );
  AND U15431 ( .A(n17083), .B(n17084), .Z(n14229) );
  XOR U15432 ( .A(n14232), .B(n14231), .Z(n14230) );
  AND U15433 ( .A(n17085), .B(n17086), .Z(n14231) );
  XOR U15434 ( .A(n14234), .B(n14233), .Z(n14232) );
  AND U15435 ( .A(n17087), .B(n17088), .Z(n14233) );
  XOR U15436 ( .A(n14236), .B(n14235), .Z(n14234) );
  AND U15437 ( .A(n17089), .B(n17090), .Z(n14235) );
  XOR U15438 ( .A(n14238), .B(n14237), .Z(n14236) );
  AND U15439 ( .A(n17091), .B(n17092), .Z(n14237) );
  XOR U15440 ( .A(n14240), .B(n14239), .Z(n14238) );
  AND U15441 ( .A(n17093), .B(n17094), .Z(n14239) );
  XOR U15442 ( .A(n14242), .B(n14241), .Z(n14240) );
  AND U15443 ( .A(n17095), .B(n17096), .Z(n14241) );
  XOR U15444 ( .A(n14244), .B(n14243), .Z(n14242) );
  AND U15445 ( .A(n17097), .B(n17098), .Z(n14243) );
  XOR U15446 ( .A(n14246), .B(n14245), .Z(n14244) );
  AND U15447 ( .A(n17099), .B(n17100), .Z(n14245) );
  XOR U15448 ( .A(n14248), .B(n14247), .Z(n14246) );
  AND U15449 ( .A(n17101), .B(n17102), .Z(n14247) );
  XOR U15450 ( .A(n14250), .B(n14249), .Z(n14248) );
  AND U15451 ( .A(n17103), .B(n17104), .Z(n14249) );
  XOR U15452 ( .A(n14252), .B(n14251), .Z(n14250) );
  AND U15453 ( .A(n17105), .B(n17106), .Z(n14251) );
  XOR U15454 ( .A(n14254), .B(n14253), .Z(n14252) );
  AND U15455 ( .A(n17107), .B(n17108), .Z(n14253) );
  XOR U15456 ( .A(n14256), .B(n14255), .Z(n14254) );
  AND U15457 ( .A(n17109), .B(n17110), .Z(n14255) );
  XOR U15458 ( .A(n14258), .B(n14257), .Z(n14256) );
  AND U15459 ( .A(n17111), .B(n17112), .Z(n14257) );
  XOR U15460 ( .A(n14260), .B(n14259), .Z(n14258) );
  AND U15461 ( .A(n17113), .B(n17114), .Z(n14259) );
  XOR U15462 ( .A(n14262), .B(n14261), .Z(n14260) );
  AND U15463 ( .A(n17115), .B(n17116), .Z(n14261) );
  XOR U15464 ( .A(n14264), .B(n14263), .Z(n14262) );
  AND U15465 ( .A(n17117), .B(n17118), .Z(n14263) );
  XOR U15466 ( .A(n14266), .B(n14265), .Z(n14264) );
  AND U15467 ( .A(n17119), .B(n17120), .Z(n14265) );
  XOR U15468 ( .A(n14268), .B(n14267), .Z(n14266) );
  AND U15469 ( .A(n17121), .B(n17122), .Z(n14267) );
  XOR U15470 ( .A(n14270), .B(n14269), .Z(n14268) );
  AND U15471 ( .A(n17123), .B(n17124), .Z(n14269) );
  XOR U15472 ( .A(n14272), .B(n14271), .Z(n14270) );
  AND U15473 ( .A(n17125), .B(n17126), .Z(n14271) );
  XOR U15474 ( .A(n14274), .B(n14273), .Z(n14272) );
  AND U15475 ( .A(n17127), .B(n17128), .Z(n14273) );
  XOR U15476 ( .A(n14276), .B(n14275), .Z(n14274) );
  AND U15477 ( .A(n17129), .B(n17130), .Z(n14275) );
  XOR U15478 ( .A(n14278), .B(n14277), .Z(n14276) );
  AND U15479 ( .A(n17131), .B(n17132), .Z(n14277) );
  XOR U15480 ( .A(n14280), .B(n14279), .Z(n14278) );
  AND U15481 ( .A(n17133), .B(n17134), .Z(n14279) );
  XOR U15482 ( .A(n14282), .B(n14281), .Z(n14280) );
  AND U15483 ( .A(n17135), .B(n17136), .Z(n14281) );
  XOR U15484 ( .A(n14284), .B(n14283), .Z(n14282) );
  AND U15485 ( .A(n17137), .B(n17138), .Z(n14283) );
  XOR U15486 ( .A(n14286), .B(n14285), .Z(n14284) );
  AND U15487 ( .A(n17139), .B(n17140), .Z(n14285) );
  XOR U15488 ( .A(n14288), .B(n14287), .Z(n14286) );
  AND U15489 ( .A(n17141), .B(n17142), .Z(n14287) );
  XOR U15490 ( .A(n14290), .B(n14289), .Z(n14288) );
  AND U15491 ( .A(n17143), .B(n17144), .Z(n14289) );
  XOR U15492 ( .A(n14292), .B(n14291), .Z(n14290) );
  AND U15493 ( .A(n17145), .B(n17146), .Z(n14291) );
  XOR U15494 ( .A(n14294), .B(n14293), .Z(n14292) );
  AND U15495 ( .A(n17147), .B(n17148), .Z(n14293) );
  XOR U15496 ( .A(n14296), .B(n14295), .Z(n14294) );
  AND U15497 ( .A(n17149), .B(n17150), .Z(n14295) );
  XOR U15498 ( .A(n14298), .B(n14297), .Z(n14296) );
  AND U15499 ( .A(n17151), .B(n17152), .Z(n14297) );
  XOR U15500 ( .A(n14300), .B(n14299), .Z(n14298) );
  AND U15501 ( .A(n17153), .B(n17154), .Z(n14299) );
  XOR U15502 ( .A(n14302), .B(n14301), .Z(n14300) );
  AND U15503 ( .A(n17155), .B(n17156), .Z(n14301) );
  XOR U15504 ( .A(n14304), .B(n14303), .Z(n14302) );
  AND U15505 ( .A(n17157), .B(n17158), .Z(n14303) );
  XOR U15506 ( .A(n14306), .B(n14305), .Z(n14304) );
  AND U15507 ( .A(n17159), .B(n17160), .Z(n14305) );
  XOR U15508 ( .A(n14308), .B(n14307), .Z(n14306) );
  AND U15509 ( .A(n17161), .B(n17162), .Z(n14307) );
  XOR U15510 ( .A(n14310), .B(n14309), .Z(n14308) );
  AND U15511 ( .A(n17163), .B(n17164), .Z(n14309) );
  XOR U15512 ( .A(n14312), .B(n14311), .Z(n14310) );
  AND U15513 ( .A(n17165), .B(n17166), .Z(n14311) );
  XOR U15514 ( .A(n14314), .B(n14313), .Z(n14312) );
  AND U15515 ( .A(n17167), .B(n17168), .Z(n14313) );
  XOR U15516 ( .A(n14316), .B(n14315), .Z(n14314) );
  AND U15517 ( .A(n17169), .B(n17170), .Z(n14315) );
  XOR U15518 ( .A(n14318), .B(n14317), .Z(n14316) );
  AND U15519 ( .A(n17171), .B(n17172), .Z(n14317) );
  XOR U15520 ( .A(n14320), .B(n14319), .Z(n14318) );
  AND U15521 ( .A(n17173), .B(n17174), .Z(n14319) );
  XOR U15522 ( .A(n14322), .B(n14321), .Z(n14320) );
  AND U15523 ( .A(n17175), .B(n17176), .Z(n14321) );
  XOR U15524 ( .A(n14324), .B(n14323), .Z(n14322) );
  AND U15525 ( .A(n17177), .B(n17178), .Z(n14323) );
  XOR U15526 ( .A(n14326), .B(n14325), .Z(n14324) );
  AND U15527 ( .A(n17179), .B(n17180), .Z(n14325) );
  XOR U15528 ( .A(n14328), .B(n14327), .Z(n14326) );
  AND U15529 ( .A(n17181), .B(n17182), .Z(n14327) );
  XOR U15530 ( .A(n14330), .B(n14329), .Z(n14328) );
  AND U15531 ( .A(n17183), .B(n17184), .Z(n14329) );
  XOR U15532 ( .A(n14332), .B(n14331), .Z(n14330) );
  AND U15533 ( .A(n17185), .B(n17186), .Z(n14331) );
  XOR U15534 ( .A(n14334), .B(n14333), .Z(n14332) );
  AND U15535 ( .A(n17187), .B(n17188), .Z(n14333) );
  XOR U15536 ( .A(n14336), .B(n14335), .Z(n14334) );
  AND U15537 ( .A(n17189), .B(n17190), .Z(n14335) );
  XOR U15538 ( .A(n14338), .B(n14337), .Z(n14336) );
  AND U15539 ( .A(n17191), .B(n17192), .Z(n14337) );
  XOR U15540 ( .A(n14340), .B(n14339), .Z(n14338) );
  AND U15541 ( .A(n17193), .B(n17194), .Z(n14339) );
  XOR U15542 ( .A(n14342), .B(n14341), .Z(n14340) );
  AND U15543 ( .A(n17195), .B(n17196), .Z(n14341) );
  XOR U15544 ( .A(n14344), .B(n14343), .Z(n14342) );
  AND U15545 ( .A(n17197), .B(n17198), .Z(n14343) );
  XOR U15546 ( .A(n14346), .B(n14345), .Z(n14344) );
  AND U15547 ( .A(n17199), .B(n17200), .Z(n14345) );
  XOR U15548 ( .A(n14348), .B(n14347), .Z(n14346) );
  AND U15549 ( .A(n17201), .B(n17202), .Z(n14347) );
  XOR U15550 ( .A(n14350), .B(n14349), .Z(n14348) );
  AND U15551 ( .A(n17203), .B(n17204), .Z(n14349) );
  XOR U15552 ( .A(n14352), .B(n14351), .Z(n14350) );
  AND U15553 ( .A(n17205), .B(n17206), .Z(n14351) );
  XOR U15554 ( .A(n14354), .B(n14353), .Z(n14352) );
  AND U15555 ( .A(n17207), .B(n17208), .Z(n14353) );
  XOR U15556 ( .A(n14356), .B(n14355), .Z(n14354) );
  AND U15557 ( .A(n17209), .B(n17210), .Z(n14355) );
  XOR U15558 ( .A(n14358), .B(n14357), .Z(n14356) );
  AND U15559 ( .A(n17211), .B(n17212), .Z(n14357) );
  XOR U15560 ( .A(n14360), .B(n14359), .Z(n14358) );
  AND U15561 ( .A(n17213), .B(n17214), .Z(n14359) );
  XOR U15562 ( .A(n14362), .B(n14361), .Z(n14360) );
  AND U15563 ( .A(n17215), .B(n17216), .Z(n14361) );
  XOR U15564 ( .A(n14364), .B(n14363), .Z(n14362) );
  AND U15565 ( .A(n17217), .B(n17218), .Z(n14363) );
  XOR U15566 ( .A(n14417), .B(n14365), .Z(n14364) );
  AND U15567 ( .A(n17219), .B(n17220), .Z(n14365) );
  XOR U15568 ( .A(n14419), .B(n14418), .Z(n14417) );
  AND U15569 ( .A(n17221), .B(n17222), .Z(n14418) );
  XOR U15570 ( .A(n14400), .B(n14420), .Z(n14419) );
  AND U15571 ( .A(n17223), .B(n17224), .Z(n14420) );
  XOR U15572 ( .A(n14402), .B(n14401), .Z(n14400) );
  AND U15573 ( .A(n17225), .B(n17226), .Z(n14401) );
  XOR U15574 ( .A(n14404), .B(n14403), .Z(n14402) );
  AND U15575 ( .A(n17227), .B(n17228), .Z(n14403) );
  XOR U15576 ( .A(n14408), .B(n14405), .Z(n14404) );
  AND U15577 ( .A(n17229), .B(n17230), .Z(n14405) );
  XOR U15578 ( .A(n14410), .B(n14409), .Z(n14408) );
  AND U15579 ( .A(n17231), .B(n17232), .Z(n14409) );
  XOR U15580 ( .A(n14413), .B(n14411), .Z(n14410) );
  AND U15581 ( .A(n17233), .B(n17234), .Z(n14411) );
  XOR U15582 ( .A(n14415), .B(n14414), .Z(n14413) );
  AND U15583 ( .A(n17235), .B(n17236), .Z(n14414) );
  XOR U15584 ( .A(n14380), .B(n14416), .Z(n14415) );
  AND U15585 ( .A(n17237), .B(n17238), .Z(n14416) );
  XNOR U15586 ( .A(n14387), .B(n14381), .Z(n14380) );
  AND U15587 ( .A(n17239), .B(n17240), .Z(n14381) );
  XOR U15588 ( .A(n14386), .B(n14378), .Z(n14387) );
  AND U15589 ( .A(n17241), .B(n17242), .Z(n14378) );
  XOR U15590 ( .A(n14399), .B(n14377), .Z(n14386) );
  AND U15591 ( .A(n17243), .B(n17244), .Z(n14377) );
  XNOR U15592 ( .A(n17245), .B(n17246), .Z(n14399) );
  XOR U15593 ( .A(n14397), .B(n17247), .Z(n17246) );
  XOR U15594 ( .A(n14395), .B(n14393), .Z(n17247) );
  AND U15595 ( .A(n17248), .B(n17249), .Z(n14393) );
  AND U15596 ( .A(n17250), .B(n17251), .Z(n14395) );
  AND U15597 ( .A(n17252), .B(n17253), .Z(n14397) );
  XNOR U15598 ( .A(n17254), .B(n14396), .Z(n17245) );
  XOR U15599 ( .A(n17255), .B(n17256), .Z(n14396) );
  XOR U15600 ( .A(n17257), .B(n17258), .Z(n17256) );
  AND U15601 ( .A(n17259), .B(n17260), .Z(n17258) );
  XNOR U15602 ( .A(n17261), .B(n17262), .Z(n17255) );
  NOR U15603 ( .A(n17263), .B(n17264), .Z(n17262) );
  AND U15604 ( .A(n17265), .B(n17266), .Z(n17264) );
  IV U15605 ( .A(n17267), .Z(n17263) );
  NOR U15606 ( .A(n17257), .B(n17268), .Z(n17267) );
  AND U15607 ( .A(n17269), .B(n17270), .Z(n17268) );
  NOR U15608 ( .A(n17259), .B(n17269), .Z(n17261) );
  XNOR U15609 ( .A(n14398), .B(n14376), .Z(n17254) );
  AND U15610 ( .A(n17271), .B(n17272), .Z(n14376) );
  AND U15611 ( .A(n17273), .B(n17274), .Z(n14398) );
  XOR U15612 ( .A(n17275), .B(n17276), .Z(n14433) );
  NOR U15613 ( .A(n17277), .B(n17278), .Z(n17276) );
  IV U15614 ( .A(n17275), .Z(n17277) );
  XOR U15615 ( .A(n17279), .B(n17280), .Z(n14436) );
  NOR U15616 ( .A(n17279), .B(n17281), .Z(n17280) );
  XNOR U15617 ( .A(n17282), .B(n17283), .Z(n14439) );
  AND U15618 ( .A(n17282), .B(n17284), .Z(n17283) );
  XNOR U15619 ( .A(n17285), .B(n17286), .Z(n14442) );
  AND U15620 ( .A(n17285), .B(n17287), .Z(n17286) );
  XNOR U15621 ( .A(n17288), .B(n17289), .Z(n14445) );
  AND U15622 ( .A(n17288), .B(n17290), .Z(n17289) );
  XNOR U15623 ( .A(n17291), .B(n17292), .Z(n14448) );
  AND U15624 ( .A(n17291), .B(n17293), .Z(n17292) );
  XNOR U15625 ( .A(n17294), .B(n17295), .Z(n14451) );
  AND U15626 ( .A(n17294), .B(n17296), .Z(n17295) );
  XNOR U15627 ( .A(n17297), .B(n17298), .Z(n14454) );
  AND U15628 ( .A(n17297), .B(n17299), .Z(n17298) );
  XNOR U15629 ( .A(n17300), .B(n17301), .Z(n14457) );
  AND U15630 ( .A(n17300), .B(n17302), .Z(n17301) );
  XNOR U15631 ( .A(n17303), .B(n17304), .Z(n14460) );
  AND U15632 ( .A(n17303), .B(n17305), .Z(n17304) );
  XNOR U15633 ( .A(n17306), .B(n17307), .Z(n14463) );
  AND U15634 ( .A(n17306), .B(n17308), .Z(n17307) );
  XNOR U15635 ( .A(n17309), .B(n17310), .Z(n14466) );
  AND U15636 ( .A(n17309), .B(n17311), .Z(n17310) );
  XNOR U15637 ( .A(n17312), .B(n17313), .Z(n14469) );
  AND U15638 ( .A(n17312), .B(n17314), .Z(n17313) );
  XNOR U15639 ( .A(n17315), .B(n17316), .Z(n14472) );
  AND U15640 ( .A(n17315), .B(n17317), .Z(n17316) );
  XNOR U15641 ( .A(n17318), .B(n17319), .Z(n14475) );
  AND U15642 ( .A(n17318), .B(n17320), .Z(n17319) );
  XNOR U15643 ( .A(n17321), .B(n17322), .Z(n14478) );
  AND U15644 ( .A(n17321), .B(n17323), .Z(n17322) );
  XNOR U15645 ( .A(n17324), .B(n17325), .Z(n14481) );
  AND U15646 ( .A(n17324), .B(n17326), .Z(n17325) );
  XNOR U15647 ( .A(n17327), .B(n17328), .Z(n14484) );
  AND U15648 ( .A(n17327), .B(n17329), .Z(n17328) );
  XNOR U15649 ( .A(n17330), .B(n17331), .Z(n14487) );
  AND U15650 ( .A(n17330), .B(n17332), .Z(n17331) );
  XNOR U15651 ( .A(n17333), .B(n17334), .Z(n14490) );
  AND U15652 ( .A(n17333), .B(n17335), .Z(n17334) );
  XNOR U15653 ( .A(n17336), .B(n17337), .Z(n14493) );
  AND U15654 ( .A(n17336), .B(n17338), .Z(n17337) );
  XNOR U15655 ( .A(n17339), .B(n17340), .Z(n14496) );
  AND U15656 ( .A(n17339), .B(n17341), .Z(n17340) );
  XNOR U15657 ( .A(n17342), .B(n17343), .Z(n14499) );
  AND U15658 ( .A(n17342), .B(n17344), .Z(n17343) );
  XNOR U15659 ( .A(n17345), .B(n17346), .Z(n14502) );
  AND U15660 ( .A(n17345), .B(n17347), .Z(n17346) );
  XNOR U15661 ( .A(n17348), .B(n17349), .Z(n14505) );
  AND U15662 ( .A(n17348), .B(n17350), .Z(n17349) );
  XNOR U15663 ( .A(n17351), .B(n17352), .Z(n14508) );
  AND U15664 ( .A(n17351), .B(n17353), .Z(n17352) );
  XNOR U15665 ( .A(n17354), .B(n17355), .Z(n14511) );
  AND U15666 ( .A(n17354), .B(n17356), .Z(n17355) );
  XNOR U15667 ( .A(n17357), .B(n17358), .Z(n14514) );
  AND U15668 ( .A(n17357), .B(n17359), .Z(n17358) );
  XNOR U15669 ( .A(n17360), .B(n17361), .Z(n14517) );
  AND U15670 ( .A(n17360), .B(n17362), .Z(n17361) );
  XNOR U15671 ( .A(n17363), .B(n17364), .Z(n14520) );
  AND U15672 ( .A(n17363), .B(n17365), .Z(n17364) );
  XNOR U15673 ( .A(n17366), .B(n17367), .Z(n14523) );
  AND U15674 ( .A(n17366), .B(n17368), .Z(n17367) );
  XNOR U15675 ( .A(n17369), .B(n17370), .Z(n14526) );
  AND U15676 ( .A(n17369), .B(n17371), .Z(n17370) );
  XNOR U15677 ( .A(n17372), .B(n17373), .Z(n14529) );
  AND U15678 ( .A(n17372), .B(n17374), .Z(n17373) );
  XNOR U15679 ( .A(n17375), .B(n17376), .Z(n14532) );
  AND U15680 ( .A(n17375), .B(n17377), .Z(n17376) );
  XNOR U15681 ( .A(n17378), .B(n17379), .Z(n14535) );
  AND U15682 ( .A(n17378), .B(n17380), .Z(n17379) );
  XNOR U15683 ( .A(n17381), .B(n17382), .Z(n14538) );
  AND U15684 ( .A(n17381), .B(n17383), .Z(n17382) );
  XNOR U15685 ( .A(n17384), .B(n17385), .Z(n14541) );
  AND U15686 ( .A(n17384), .B(n17386), .Z(n17385) );
  XNOR U15687 ( .A(n17387), .B(n17388), .Z(n14544) );
  AND U15688 ( .A(n17387), .B(n17389), .Z(n17388) );
  XNOR U15689 ( .A(n17390), .B(n17391), .Z(n14547) );
  AND U15690 ( .A(n17390), .B(n17392), .Z(n17391) );
  XNOR U15691 ( .A(n17393), .B(n17394), .Z(n14550) );
  AND U15692 ( .A(n17393), .B(n17395), .Z(n17394) );
  XNOR U15693 ( .A(n17396), .B(n17397), .Z(n14553) );
  AND U15694 ( .A(n17396), .B(n17398), .Z(n17397) );
  XNOR U15695 ( .A(n17399), .B(n17400), .Z(n14556) );
  AND U15696 ( .A(n17399), .B(n17401), .Z(n17400) );
  XNOR U15697 ( .A(n17402), .B(n17403), .Z(n14559) );
  AND U15698 ( .A(n17402), .B(n17404), .Z(n17403) );
  XNOR U15699 ( .A(n17405), .B(n17406), .Z(n14562) );
  AND U15700 ( .A(n17405), .B(n17407), .Z(n17406) );
  XNOR U15701 ( .A(n17408), .B(n17409), .Z(n14565) );
  AND U15702 ( .A(n17408), .B(n17410), .Z(n17409) );
  XNOR U15703 ( .A(n17411), .B(n17412), .Z(n14568) );
  AND U15704 ( .A(n17411), .B(n17413), .Z(n17412) );
  XNOR U15705 ( .A(n17414), .B(n17415), .Z(n14571) );
  AND U15706 ( .A(n17414), .B(n17416), .Z(n17415) );
  XNOR U15707 ( .A(n17417), .B(n17418), .Z(n14574) );
  AND U15708 ( .A(n17417), .B(n17419), .Z(n17418) );
  XNOR U15709 ( .A(n17420), .B(n17421), .Z(n14577) );
  AND U15710 ( .A(n17420), .B(n17422), .Z(n17421) );
  XNOR U15711 ( .A(n17423), .B(n17424), .Z(n14580) );
  AND U15712 ( .A(n17423), .B(n17425), .Z(n17424) );
  XNOR U15713 ( .A(n17426), .B(n17427), .Z(n14583) );
  AND U15714 ( .A(n17426), .B(n17428), .Z(n17427) );
  XNOR U15715 ( .A(n17429), .B(n17430), .Z(n14586) );
  AND U15716 ( .A(n17429), .B(n17431), .Z(n17430) );
  XNOR U15717 ( .A(n17432), .B(n17433), .Z(n14589) );
  AND U15718 ( .A(n17432), .B(n17434), .Z(n17433) );
  XNOR U15719 ( .A(n17435), .B(n17436), .Z(n14592) );
  AND U15720 ( .A(n17435), .B(n17437), .Z(n17436) );
  XNOR U15721 ( .A(n17438), .B(n17439), .Z(n14595) );
  AND U15722 ( .A(n17438), .B(n17440), .Z(n17439) );
  XNOR U15723 ( .A(n17441), .B(n17442), .Z(n14598) );
  AND U15724 ( .A(n17441), .B(n17443), .Z(n17442) );
  XNOR U15725 ( .A(n17444), .B(n17445), .Z(n14601) );
  AND U15726 ( .A(n17444), .B(n17446), .Z(n17445) );
  XNOR U15727 ( .A(n17447), .B(n17448), .Z(n14604) );
  AND U15728 ( .A(n17447), .B(n17449), .Z(n17448) );
  XNOR U15729 ( .A(n17450), .B(n17451), .Z(n14607) );
  AND U15730 ( .A(n17450), .B(n17452), .Z(n17451) );
  XNOR U15731 ( .A(n17453), .B(n17454), .Z(n14610) );
  AND U15732 ( .A(n17453), .B(n17455), .Z(n17454) );
  XNOR U15733 ( .A(n17456), .B(n17457), .Z(n14613) );
  AND U15734 ( .A(n17456), .B(n17458), .Z(n17457) );
  XNOR U15735 ( .A(n17459), .B(n17460), .Z(n14616) );
  AND U15736 ( .A(n17459), .B(n17461), .Z(n17460) );
  XNOR U15737 ( .A(n17462), .B(n17463), .Z(n14619) );
  AND U15738 ( .A(n17462), .B(n17464), .Z(n17463) );
  XNOR U15739 ( .A(n17465), .B(n17466), .Z(n14622) );
  AND U15740 ( .A(n17465), .B(n17467), .Z(n17466) );
  XNOR U15741 ( .A(n17468), .B(n17469), .Z(n14625) );
  AND U15742 ( .A(n17468), .B(n17470), .Z(n17469) );
  XNOR U15743 ( .A(n17471), .B(n17472), .Z(n14628) );
  AND U15744 ( .A(n17471), .B(n17473), .Z(n17472) );
  XNOR U15745 ( .A(n17474), .B(n17475), .Z(n14631) );
  AND U15746 ( .A(n17474), .B(n17476), .Z(n17475) );
  XNOR U15747 ( .A(n17477), .B(n17478), .Z(n14634) );
  AND U15748 ( .A(n17477), .B(n17479), .Z(n17478) );
  XNOR U15749 ( .A(n17480), .B(n17481), .Z(n14637) );
  AND U15750 ( .A(n17480), .B(n17482), .Z(n17481) );
  XNOR U15751 ( .A(n17483), .B(n17484), .Z(n14640) );
  AND U15752 ( .A(n17483), .B(n17485), .Z(n17484) );
  XNOR U15753 ( .A(n17486), .B(n17487), .Z(n14643) );
  AND U15754 ( .A(n17486), .B(n17488), .Z(n17487) );
  XNOR U15755 ( .A(n17489), .B(n17490), .Z(n14646) );
  AND U15756 ( .A(n17489), .B(n17491), .Z(n17490) );
  XNOR U15757 ( .A(n17492), .B(n17493), .Z(n14649) );
  AND U15758 ( .A(n17492), .B(n17494), .Z(n17493) );
  XNOR U15759 ( .A(n17495), .B(n17496), .Z(n14652) );
  AND U15760 ( .A(n17495), .B(n17497), .Z(n17496) );
  XNOR U15761 ( .A(n17498), .B(n17499), .Z(n14655) );
  AND U15762 ( .A(n17498), .B(n17500), .Z(n17499) );
  XNOR U15763 ( .A(n17501), .B(n17502), .Z(n14658) );
  AND U15764 ( .A(n17501), .B(n17503), .Z(n17502) );
  XNOR U15765 ( .A(n17504), .B(n17505), .Z(n14661) );
  AND U15766 ( .A(n17504), .B(n17506), .Z(n17505) );
  XNOR U15767 ( .A(n17507), .B(n17508), .Z(n14664) );
  AND U15768 ( .A(n17507), .B(n17509), .Z(n17508) );
  XNOR U15769 ( .A(n17510), .B(n17511), .Z(n14667) );
  AND U15770 ( .A(n17510), .B(n17512), .Z(n17511) );
  XNOR U15771 ( .A(n17513), .B(n17514), .Z(n14670) );
  AND U15772 ( .A(n17513), .B(n17515), .Z(n17514) );
  XNOR U15773 ( .A(n17516), .B(n17517), .Z(n14673) );
  AND U15774 ( .A(n17516), .B(n17518), .Z(n17517) );
  XNOR U15775 ( .A(n17519), .B(n17520), .Z(n14676) );
  AND U15776 ( .A(n17519), .B(n17521), .Z(n17520) );
  XNOR U15777 ( .A(n17522), .B(n17523), .Z(n14679) );
  AND U15778 ( .A(n17522), .B(n17524), .Z(n17523) );
  XNOR U15779 ( .A(n17525), .B(n17526), .Z(n14682) );
  AND U15780 ( .A(n17525), .B(n17527), .Z(n17526) );
  XNOR U15781 ( .A(n17528), .B(n17529), .Z(n14685) );
  AND U15782 ( .A(n17528), .B(n17530), .Z(n17529) );
  XNOR U15783 ( .A(n17531), .B(n17532), .Z(n14688) );
  AND U15784 ( .A(n17531), .B(n17533), .Z(n17532) );
  XNOR U15785 ( .A(n17534), .B(n17535), .Z(n14691) );
  AND U15786 ( .A(n17534), .B(n17536), .Z(n17535) );
  XNOR U15787 ( .A(n17537), .B(n17538), .Z(n14694) );
  AND U15788 ( .A(n17537), .B(n17539), .Z(n17538) );
  XNOR U15789 ( .A(n17540), .B(n17541), .Z(n14697) );
  AND U15790 ( .A(n17540), .B(n17542), .Z(n17541) );
  XNOR U15791 ( .A(n17543), .B(n17544), .Z(n14700) );
  AND U15792 ( .A(n17543), .B(n17545), .Z(n17544) );
  XNOR U15793 ( .A(n17546), .B(n17547), .Z(n14703) );
  AND U15794 ( .A(n17546), .B(n17548), .Z(n17547) );
  XNOR U15795 ( .A(n17549), .B(n17550), .Z(n14706) );
  AND U15796 ( .A(n17549), .B(n17551), .Z(n17550) );
  XNOR U15797 ( .A(n17552), .B(n17553), .Z(n14709) );
  AND U15798 ( .A(n17552), .B(n17554), .Z(n17553) );
  XNOR U15799 ( .A(n17555), .B(n17556), .Z(n14712) );
  AND U15800 ( .A(n17555), .B(n17557), .Z(n17556) );
  XNOR U15801 ( .A(n17558), .B(n17559), .Z(n14715) );
  AND U15802 ( .A(n17558), .B(n17560), .Z(n17559) );
  XNOR U15803 ( .A(n17561), .B(n17562), .Z(n14718) );
  AND U15804 ( .A(n17561), .B(n17563), .Z(n17562) );
  XNOR U15805 ( .A(n17564), .B(n17565), .Z(n14721) );
  AND U15806 ( .A(n17564), .B(n17566), .Z(n17565) );
  XNOR U15807 ( .A(n17567), .B(n17568), .Z(n14724) );
  AND U15808 ( .A(n17567), .B(n17569), .Z(n17568) );
  XNOR U15809 ( .A(n17570), .B(n17571), .Z(n14727) );
  AND U15810 ( .A(n17570), .B(n17572), .Z(n17571) );
  XNOR U15811 ( .A(n17573), .B(n17574), .Z(n14730) );
  AND U15812 ( .A(n17573), .B(n17575), .Z(n17574) );
  XNOR U15813 ( .A(n17576), .B(n17577), .Z(n14733) );
  AND U15814 ( .A(n17576), .B(n17578), .Z(n17577) );
  XNOR U15815 ( .A(n17579), .B(n17580), .Z(n14736) );
  AND U15816 ( .A(n17579), .B(n17581), .Z(n17580) );
  XNOR U15817 ( .A(n17582), .B(n17583), .Z(n14739) );
  AND U15818 ( .A(n17582), .B(n17584), .Z(n17583) );
  XNOR U15819 ( .A(n17585), .B(n17586), .Z(n14742) );
  AND U15820 ( .A(n17585), .B(n17587), .Z(n17586) );
  XNOR U15821 ( .A(n17588), .B(n17589), .Z(n14745) );
  AND U15822 ( .A(n17588), .B(n17590), .Z(n17589) );
  XNOR U15823 ( .A(n17591), .B(n17592), .Z(n14748) );
  AND U15824 ( .A(n17591), .B(n17593), .Z(n17592) );
  XNOR U15825 ( .A(n17594), .B(n17595), .Z(n14751) );
  AND U15826 ( .A(n17594), .B(n17596), .Z(n17595) );
  XNOR U15827 ( .A(n17597), .B(n17598), .Z(n14754) );
  AND U15828 ( .A(n17597), .B(n17599), .Z(n17598) );
  XNOR U15829 ( .A(n17600), .B(n17601), .Z(n14757) );
  AND U15830 ( .A(n17600), .B(n17602), .Z(n17601) );
  XNOR U15831 ( .A(n17603), .B(n17604), .Z(n14760) );
  AND U15832 ( .A(n17603), .B(n17605), .Z(n17604) );
  XNOR U15833 ( .A(n17606), .B(n17607), .Z(n14763) );
  AND U15834 ( .A(n17606), .B(n17608), .Z(n17607) );
  XNOR U15835 ( .A(n17609), .B(n17610), .Z(n14766) );
  AND U15836 ( .A(n17609), .B(n17611), .Z(n17610) );
  XNOR U15837 ( .A(n17612), .B(n17613), .Z(n14769) );
  AND U15838 ( .A(n17612), .B(n17614), .Z(n17613) );
  XNOR U15839 ( .A(n17615), .B(n17616), .Z(n14772) );
  AND U15840 ( .A(n17615), .B(n17617), .Z(n17616) );
  XNOR U15841 ( .A(n17618), .B(n17619), .Z(n14775) );
  AND U15842 ( .A(n17618), .B(n17620), .Z(n17619) );
  XNOR U15843 ( .A(n17621), .B(n17622), .Z(n14778) );
  AND U15844 ( .A(n17621), .B(n17623), .Z(n17622) );
  XNOR U15845 ( .A(n17624), .B(n17625), .Z(n14781) );
  AND U15846 ( .A(n17624), .B(n17626), .Z(n17625) );
  XNOR U15847 ( .A(n17627), .B(n17628), .Z(n14784) );
  AND U15848 ( .A(n17627), .B(n17629), .Z(n17628) );
  XNOR U15849 ( .A(n17630), .B(n17631), .Z(n14787) );
  AND U15850 ( .A(n17630), .B(n17632), .Z(n17631) );
  XNOR U15851 ( .A(n17633), .B(n17634), .Z(n14790) );
  AND U15852 ( .A(n17633), .B(n17635), .Z(n17634) );
  XNOR U15853 ( .A(n17636), .B(n17637), .Z(n14793) );
  AND U15854 ( .A(n17636), .B(n17638), .Z(n17637) );
  XNOR U15855 ( .A(n17639), .B(n17640), .Z(n14796) );
  AND U15856 ( .A(n17639), .B(n17641), .Z(n17640) );
  XNOR U15857 ( .A(n17642), .B(n17643), .Z(n14799) );
  AND U15858 ( .A(n17642), .B(n17644), .Z(n17643) );
  XNOR U15859 ( .A(n17645), .B(n17646), .Z(n14802) );
  AND U15860 ( .A(n17645), .B(n17647), .Z(n17646) );
  XNOR U15861 ( .A(n17648), .B(n17649), .Z(n14805) );
  AND U15862 ( .A(n17648), .B(n17650), .Z(n17649) );
  XNOR U15863 ( .A(n17651), .B(n17652), .Z(n14808) );
  AND U15864 ( .A(n17651), .B(n17653), .Z(n17652) );
  XNOR U15865 ( .A(n17654), .B(n17655), .Z(n14811) );
  AND U15866 ( .A(n17654), .B(n17656), .Z(n17655) );
  XNOR U15867 ( .A(n17657), .B(n17658), .Z(n14814) );
  AND U15868 ( .A(n17657), .B(n17659), .Z(n17658) );
  XNOR U15869 ( .A(n17660), .B(n17661), .Z(n14817) );
  AND U15870 ( .A(n17660), .B(n17662), .Z(n17661) );
  XNOR U15871 ( .A(n17663), .B(n17664), .Z(n14820) );
  AND U15872 ( .A(n17663), .B(n17665), .Z(n17664) );
  XNOR U15873 ( .A(n17666), .B(n17667), .Z(n14823) );
  AND U15874 ( .A(n17666), .B(n17668), .Z(n17667) );
  XNOR U15875 ( .A(n17669), .B(n17670), .Z(n14826) );
  AND U15876 ( .A(n17669), .B(n17671), .Z(n17670) );
  XNOR U15877 ( .A(n17672), .B(n17673), .Z(n14829) );
  AND U15878 ( .A(n17672), .B(n17674), .Z(n17673) );
  XNOR U15879 ( .A(n17675), .B(n17676), .Z(n14832) );
  AND U15880 ( .A(n17675), .B(n17677), .Z(n17676) );
  XNOR U15881 ( .A(n17678), .B(n17679), .Z(n14835) );
  AND U15882 ( .A(n17678), .B(n17680), .Z(n17679) );
  XNOR U15883 ( .A(n17681), .B(n17682), .Z(n14838) );
  AND U15884 ( .A(n17681), .B(n17683), .Z(n17682) );
  XNOR U15885 ( .A(n17684), .B(n17685), .Z(n14841) );
  AND U15886 ( .A(n17684), .B(n17686), .Z(n17685) );
  XNOR U15887 ( .A(n17687), .B(n17688), .Z(n14844) );
  AND U15888 ( .A(n17687), .B(n17689), .Z(n17688) );
  XNOR U15889 ( .A(n17690), .B(n17691), .Z(n14847) );
  AND U15890 ( .A(n17690), .B(n17692), .Z(n17691) );
  XNOR U15891 ( .A(n17693), .B(n17694), .Z(n14850) );
  AND U15892 ( .A(n17693), .B(n17695), .Z(n17694) );
  XNOR U15893 ( .A(n17696), .B(n17697), .Z(n14853) );
  AND U15894 ( .A(n17696), .B(n17698), .Z(n17697) );
  XNOR U15895 ( .A(n17699), .B(n17700), .Z(n14856) );
  AND U15896 ( .A(n17699), .B(n17701), .Z(n17700) );
  XNOR U15897 ( .A(n17702), .B(n17703), .Z(n14859) );
  AND U15898 ( .A(n17702), .B(n17704), .Z(n17703) );
  XNOR U15899 ( .A(n17705), .B(n17706), .Z(n14862) );
  AND U15900 ( .A(n17705), .B(n17707), .Z(n17706) );
  XNOR U15901 ( .A(n17708), .B(n17709), .Z(n14865) );
  AND U15902 ( .A(n17708), .B(n17710), .Z(n17709) );
  XNOR U15903 ( .A(n17711), .B(n17712), .Z(n14868) );
  AND U15904 ( .A(n17711), .B(n17713), .Z(n17712) );
  XNOR U15905 ( .A(n17714), .B(n17715), .Z(n14871) );
  AND U15906 ( .A(n17714), .B(n17716), .Z(n17715) );
  XNOR U15907 ( .A(n17717), .B(n17718), .Z(n14874) );
  AND U15908 ( .A(n17717), .B(n17719), .Z(n17718) );
  XNOR U15909 ( .A(n17720), .B(n17721), .Z(n14877) );
  AND U15910 ( .A(n17720), .B(n17722), .Z(n17721) );
  XNOR U15911 ( .A(n17723), .B(n17724), .Z(n14880) );
  AND U15912 ( .A(n17723), .B(n17725), .Z(n17724) );
  XNOR U15913 ( .A(n17726), .B(n17727), .Z(n14883) );
  AND U15914 ( .A(n17726), .B(n17728), .Z(n17727) );
  XNOR U15915 ( .A(n17729), .B(n17730), .Z(n14886) );
  AND U15916 ( .A(n17729), .B(n17731), .Z(n17730) );
  XNOR U15917 ( .A(n17732), .B(n17733), .Z(n14889) );
  AND U15918 ( .A(n17732), .B(n17734), .Z(n17733) );
  XNOR U15919 ( .A(n17735), .B(n17736), .Z(n14892) );
  AND U15920 ( .A(n17735), .B(n17737), .Z(n17736) );
  XNOR U15921 ( .A(n17738), .B(n17739), .Z(n14895) );
  AND U15922 ( .A(n17738), .B(n17740), .Z(n17739) );
  XNOR U15923 ( .A(n17741), .B(n17742), .Z(n14898) );
  AND U15924 ( .A(n17741), .B(n17743), .Z(n17742) );
  XNOR U15925 ( .A(n17744), .B(n17745), .Z(n14901) );
  AND U15926 ( .A(n17744), .B(n17746), .Z(n17745) );
  XNOR U15927 ( .A(n17747), .B(n17748), .Z(n14904) );
  AND U15928 ( .A(n17747), .B(n17749), .Z(n17748) );
  XNOR U15929 ( .A(n17750), .B(n17751), .Z(n14907) );
  AND U15930 ( .A(n17750), .B(n17752), .Z(n17751) );
  XNOR U15931 ( .A(n17753), .B(n17754), .Z(n14910) );
  AND U15932 ( .A(n17753), .B(n17755), .Z(n17754) );
  XNOR U15933 ( .A(n17756), .B(n17757), .Z(n14913) );
  AND U15934 ( .A(n17756), .B(n17758), .Z(n17757) );
  XNOR U15935 ( .A(n17759), .B(n17760), .Z(n14916) );
  AND U15936 ( .A(n17759), .B(n17761), .Z(n17760) );
  XNOR U15937 ( .A(n17762), .B(n17763), .Z(n14919) );
  AND U15938 ( .A(n17762), .B(n17764), .Z(n17763) );
  XNOR U15939 ( .A(n17765), .B(n17766), .Z(n14922) );
  AND U15940 ( .A(n17765), .B(n17767), .Z(n17766) );
  XNOR U15941 ( .A(n17768), .B(n17769), .Z(n14925) );
  AND U15942 ( .A(n17768), .B(n17770), .Z(n17769) );
  XNOR U15943 ( .A(n17771), .B(n17772), .Z(n14928) );
  AND U15944 ( .A(n17771), .B(n17773), .Z(n17772) );
  XNOR U15945 ( .A(n17774), .B(n17775), .Z(n14931) );
  AND U15946 ( .A(n17774), .B(n17776), .Z(n17775) );
  XNOR U15947 ( .A(n17777), .B(n17778), .Z(n14934) );
  AND U15948 ( .A(n17777), .B(n17779), .Z(n17778) );
  XNOR U15949 ( .A(n17780), .B(n17781), .Z(n14937) );
  AND U15950 ( .A(n17780), .B(n17782), .Z(n17781) );
  XNOR U15951 ( .A(n17783), .B(n17784), .Z(n14940) );
  AND U15952 ( .A(n17783), .B(n17785), .Z(n17784) );
  XNOR U15953 ( .A(n17786), .B(n17787), .Z(n14943) );
  AND U15954 ( .A(n17786), .B(n17788), .Z(n17787) );
  XNOR U15955 ( .A(n17789), .B(n17790), .Z(n14946) );
  AND U15956 ( .A(n17789), .B(n17791), .Z(n17790) );
  XNOR U15957 ( .A(n17792), .B(n17793), .Z(n14949) );
  AND U15958 ( .A(n17792), .B(n17794), .Z(n17793) );
  XNOR U15959 ( .A(n17795), .B(n17796), .Z(n14952) );
  AND U15960 ( .A(n17795), .B(n17797), .Z(n17796) );
  XNOR U15961 ( .A(n17798), .B(n17799), .Z(n14955) );
  AND U15962 ( .A(n17798), .B(n17800), .Z(n17799) );
  XNOR U15963 ( .A(n17801), .B(n17802), .Z(n14958) );
  AND U15964 ( .A(n17801), .B(n17803), .Z(n17802) );
  XNOR U15965 ( .A(n17804), .B(n17805), .Z(n14961) );
  AND U15966 ( .A(n17804), .B(n17806), .Z(n17805) );
  XNOR U15967 ( .A(n17807), .B(n17808), .Z(n14964) );
  AND U15968 ( .A(n17807), .B(n17809), .Z(n17808) );
  XNOR U15969 ( .A(n17810), .B(n17811), .Z(n14967) );
  AND U15970 ( .A(n17810), .B(n17812), .Z(n17811) );
  XNOR U15971 ( .A(n17813), .B(n17814), .Z(n14970) );
  AND U15972 ( .A(n17813), .B(n17815), .Z(n17814) );
  XNOR U15973 ( .A(n17816), .B(n17817), .Z(n14973) );
  AND U15974 ( .A(n17816), .B(n17818), .Z(n17817) );
  XNOR U15975 ( .A(n17819), .B(n17820), .Z(n14976) );
  AND U15976 ( .A(n17819), .B(n17821), .Z(n17820) );
  XNOR U15977 ( .A(n17822), .B(n17823), .Z(n14979) );
  AND U15978 ( .A(n17822), .B(n17824), .Z(n17823) );
  XNOR U15979 ( .A(n17825), .B(n17826), .Z(n14982) );
  AND U15980 ( .A(n17825), .B(n17827), .Z(n17826) );
  XNOR U15981 ( .A(n17828), .B(n17829), .Z(n14985) );
  AND U15982 ( .A(n17828), .B(n17830), .Z(n17829) );
  XNOR U15983 ( .A(n17831), .B(n17832), .Z(n14988) );
  AND U15984 ( .A(n17831), .B(n17833), .Z(n17832) );
  XNOR U15985 ( .A(n17834), .B(n17835), .Z(n14991) );
  AND U15986 ( .A(n17834), .B(n17836), .Z(n17835) );
  XNOR U15987 ( .A(n17837), .B(n17838), .Z(n14994) );
  AND U15988 ( .A(n17837), .B(n17839), .Z(n17838) );
  XNOR U15989 ( .A(n17840), .B(n17841), .Z(n14997) );
  AND U15990 ( .A(n17840), .B(n17842), .Z(n17841) );
  XNOR U15991 ( .A(n17843), .B(n17844), .Z(n15000) );
  AND U15992 ( .A(n17843), .B(n17845), .Z(n17844) );
  XNOR U15993 ( .A(n17846), .B(n17847), .Z(n15003) );
  AND U15994 ( .A(n17846), .B(n17848), .Z(n17847) );
  XNOR U15995 ( .A(n17849), .B(n17850), .Z(n15006) );
  AND U15996 ( .A(n17849), .B(n17851), .Z(n17850) );
  XNOR U15997 ( .A(n17852), .B(n17853), .Z(n15009) );
  AND U15998 ( .A(n17852), .B(n17854), .Z(n17853) );
  XNOR U15999 ( .A(n17855), .B(n17856), .Z(n15012) );
  AND U16000 ( .A(n17855), .B(n17857), .Z(n17856) );
  XNOR U16001 ( .A(n17858), .B(n17859), .Z(n15015) );
  AND U16002 ( .A(n17858), .B(n17860), .Z(n17859) );
  XNOR U16003 ( .A(n17861), .B(n17862), .Z(n15018) );
  AND U16004 ( .A(n17861), .B(n17863), .Z(n17862) );
  XNOR U16005 ( .A(n17864), .B(n17865), .Z(n15021) );
  AND U16006 ( .A(n17864), .B(n17866), .Z(n17865) );
  XNOR U16007 ( .A(n17867), .B(n17868), .Z(n15024) );
  AND U16008 ( .A(n17867), .B(n17869), .Z(n17868) );
  XNOR U16009 ( .A(n17870), .B(n17871), .Z(n15027) );
  AND U16010 ( .A(n17870), .B(n17872), .Z(n17871) );
  XNOR U16011 ( .A(n17873), .B(n17874), .Z(n15030) );
  AND U16012 ( .A(n17873), .B(n17875), .Z(n17874) );
  XNOR U16013 ( .A(n17876), .B(n17877), .Z(n15033) );
  AND U16014 ( .A(n17876), .B(n17878), .Z(n17877) );
  XNOR U16015 ( .A(n17879), .B(n17880), .Z(n15036) );
  AND U16016 ( .A(n17879), .B(n17881), .Z(n17880) );
  XNOR U16017 ( .A(n17882), .B(n17883), .Z(n15039) );
  AND U16018 ( .A(n17882), .B(n17884), .Z(n17883) );
  XNOR U16019 ( .A(n17885), .B(n17886), .Z(n15042) );
  AND U16020 ( .A(n17885), .B(n17887), .Z(n17886) );
  XNOR U16021 ( .A(n17888), .B(n17889), .Z(n15045) );
  AND U16022 ( .A(n17888), .B(n17890), .Z(n17889) );
  XNOR U16023 ( .A(n17891), .B(n17892), .Z(n15048) );
  AND U16024 ( .A(n17891), .B(n17893), .Z(n17892) );
  XNOR U16025 ( .A(n17894), .B(n17895), .Z(n15051) );
  AND U16026 ( .A(n17894), .B(n17896), .Z(n17895) );
  XNOR U16027 ( .A(n17897), .B(n17898), .Z(n15054) );
  AND U16028 ( .A(n17897), .B(n17899), .Z(n17898) );
  XNOR U16029 ( .A(n17900), .B(n17901), .Z(n15057) );
  AND U16030 ( .A(n17900), .B(n17902), .Z(n17901) );
  XNOR U16031 ( .A(n17903), .B(n17904), .Z(n15060) );
  AND U16032 ( .A(n17903), .B(n17905), .Z(n17904) );
  XNOR U16033 ( .A(n17906), .B(n17907), .Z(n15063) );
  AND U16034 ( .A(n17906), .B(n17908), .Z(n17907) );
  XNOR U16035 ( .A(n17909), .B(n17910), .Z(n15066) );
  AND U16036 ( .A(n17909), .B(n17911), .Z(n17910) );
  XNOR U16037 ( .A(n17912), .B(n17913), .Z(n15069) );
  AND U16038 ( .A(n17912), .B(n17914), .Z(n17913) );
  XNOR U16039 ( .A(n17915), .B(n17916), .Z(n15072) );
  AND U16040 ( .A(n17915), .B(n17917), .Z(n17916) );
  XNOR U16041 ( .A(n17918), .B(n17919), .Z(n15075) );
  AND U16042 ( .A(n17918), .B(n17920), .Z(n17919) );
  XNOR U16043 ( .A(n17921), .B(n17922), .Z(n15078) );
  AND U16044 ( .A(n17921), .B(n17923), .Z(n17922) );
  XNOR U16045 ( .A(n17924), .B(n17925), .Z(n15081) );
  AND U16046 ( .A(n17924), .B(n17926), .Z(n17925) );
  XNOR U16047 ( .A(n17927), .B(n17928), .Z(n15084) );
  AND U16048 ( .A(n17927), .B(n17929), .Z(n17928) );
  XNOR U16049 ( .A(n17930), .B(n17931), .Z(n15087) );
  AND U16050 ( .A(n17930), .B(n17932), .Z(n17931) );
  XNOR U16051 ( .A(n17933), .B(n17934), .Z(n15090) );
  AND U16052 ( .A(n17933), .B(n17935), .Z(n17934) );
  XNOR U16053 ( .A(n17936), .B(n17937), .Z(n15093) );
  AND U16054 ( .A(n17936), .B(n17938), .Z(n17937) );
  XNOR U16055 ( .A(n17939), .B(n17940), .Z(n15096) );
  AND U16056 ( .A(n17939), .B(n17941), .Z(n17940) );
  XNOR U16057 ( .A(n17942), .B(n17943), .Z(n15099) );
  AND U16058 ( .A(n17942), .B(n17944), .Z(n17943) );
  XNOR U16059 ( .A(n17945), .B(n17946), .Z(n15102) );
  AND U16060 ( .A(n17945), .B(n17947), .Z(n17946) );
  XNOR U16061 ( .A(n17948), .B(n17949), .Z(n15105) );
  AND U16062 ( .A(n17948), .B(n17950), .Z(n17949) );
  XNOR U16063 ( .A(n17951), .B(n17952), .Z(n15108) );
  AND U16064 ( .A(n17951), .B(n17953), .Z(n17952) );
  XNOR U16065 ( .A(n17954), .B(n17955), .Z(n15111) );
  AND U16066 ( .A(n17954), .B(n17956), .Z(n17955) );
  XNOR U16067 ( .A(n17957), .B(n17958), .Z(n15114) );
  AND U16068 ( .A(n17957), .B(n17959), .Z(n17958) );
  XNOR U16069 ( .A(n17960), .B(n17961), .Z(n15117) );
  AND U16070 ( .A(n17960), .B(n17962), .Z(n17961) );
  XNOR U16071 ( .A(n17963), .B(n17964), .Z(n15120) );
  AND U16072 ( .A(n17963), .B(n17965), .Z(n17964) );
  XNOR U16073 ( .A(n17966), .B(n17967), .Z(n15123) );
  AND U16074 ( .A(n17966), .B(n17968), .Z(n17967) );
  XNOR U16075 ( .A(n17969), .B(n17970), .Z(n15126) );
  AND U16076 ( .A(n17969), .B(n17971), .Z(n17970) );
  XNOR U16077 ( .A(n17972), .B(n17973), .Z(n15129) );
  AND U16078 ( .A(n17972), .B(n17974), .Z(n17973) );
  XNOR U16079 ( .A(n17975), .B(n17976), .Z(n15132) );
  AND U16080 ( .A(n17975), .B(n17977), .Z(n17976) );
  XNOR U16081 ( .A(n17978), .B(n17979), .Z(n15135) );
  AND U16082 ( .A(n17978), .B(n17980), .Z(n17979) );
  XNOR U16083 ( .A(n17981), .B(n17982), .Z(n15138) );
  AND U16084 ( .A(n17981), .B(n17983), .Z(n17982) );
  XNOR U16085 ( .A(n17984), .B(n17985), .Z(n15141) );
  AND U16086 ( .A(n17984), .B(n17986), .Z(n17985) );
  XNOR U16087 ( .A(n17987), .B(n17988), .Z(n15144) );
  AND U16088 ( .A(n17987), .B(n17989), .Z(n17988) );
  XNOR U16089 ( .A(n17990), .B(n17991), .Z(n15147) );
  AND U16090 ( .A(n17990), .B(n17992), .Z(n17991) );
  XNOR U16091 ( .A(n17993), .B(n17994), .Z(n15150) );
  AND U16092 ( .A(n17993), .B(n17995), .Z(n17994) );
  XNOR U16093 ( .A(n17996), .B(n17997), .Z(n15153) );
  AND U16094 ( .A(n17996), .B(n17998), .Z(n17997) );
  XNOR U16095 ( .A(n17999), .B(n18000), .Z(n15156) );
  AND U16096 ( .A(n17999), .B(n18001), .Z(n18000) );
  XNOR U16097 ( .A(n18002), .B(n18003), .Z(n15159) );
  AND U16098 ( .A(n18002), .B(n18004), .Z(n18003) );
  XNOR U16099 ( .A(n18005), .B(n18006), .Z(n15162) );
  AND U16100 ( .A(n18005), .B(n18007), .Z(n18006) );
  XNOR U16101 ( .A(n18008), .B(n18009), .Z(n15165) );
  AND U16102 ( .A(n18008), .B(n18010), .Z(n18009) );
  XNOR U16103 ( .A(n18011), .B(n18012), .Z(n15168) );
  AND U16104 ( .A(n18011), .B(n18013), .Z(n18012) );
  XNOR U16105 ( .A(n18014), .B(n18015), .Z(n15171) );
  AND U16106 ( .A(n18014), .B(n18016), .Z(n18015) );
  XNOR U16107 ( .A(n18017), .B(n18018), .Z(n15174) );
  AND U16108 ( .A(n18017), .B(n18019), .Z(n18018) );
  XNOR U16109 ( .A(n18020), .B(n18021), .Z(n15177) );
  AND U16110 ( .A(n18020), .B(n18022), .Z(n18021) );
  XNOR U16111 ( .A(n18023), .B(n18024), .Z(n15180) );
  AND U16112 ( .A(n18023), .B(n18025), .Z(n18024) );
  XNOR U16113 ( .A(n18026), .B(n18027), .Z(n15183) );
  AND U16114 ( .A(n18026), .B(n18028), .Z(n18027) );
  XNOR U16115 ( .A(n18029), .B(n18030), .Z(n15186) );
  AND U16116 ( .A(n18029), .B(n18031), .Z(n18030) );
  XNOR U16117 ( .A(n18032), .B(n18033), .Z(n15189) );
  AND U16118 ( .A(n18032), .B(n18034), .Z(n18033) );
  XNOR U16119 ( .A(n18035), .B(n18036), .Z(n15192) );
  AND U16120 ( .A(n18035), .B(n18037), .Z(n18036) );
  XNOR U16121 ( .A(n18038), .B(n18039), .Z(n15195) );
  AND U16122 ( .A(n18038), .B(n18040), .Z(n18039) );
  XNOR U16123 ( .A(n18041), .B(n18042), .Z(n15198) );
  AND U16124 ( .A(n18041), .B(n18043), .Z(n18042) );
  XNOR U16125 ( .A(n18044), .B(n18045), .Z(n15201) );
  AND U16126 ( .A(n18044), .B(n18046), .Z(n18045) );
  XNOR U16127 ( .A(n18047), .B(n18048), .Z(n15204) );
  AND U16128 ( .A(n18047), .B(n18049), .Z(n18048) );
  XNOR U16129 ( .A(n18050), .B(n18051), .Z(n15207) );
  AND U16130 ( .A(n18050), .B(n18052), .Z(n18051) );
  XNOR U16131 ( .A(n18053), .B(n18054), .Z(n15210) );
  AND U16132 ( .A(n18053), .B(n18055), .Z(n18054) );
  XNOR U16133 ( .A(n18056), .B(n18057), .Z(n15213) );
  AND U16134 ( .A(n18056), .B(n18058), .Z(n18057) );
  XNOR U16135 ( .A(n18059), .B(n18060), .Z(n15216) );
  AND U16136 ( .A(n18059), .B(n18061), .Z(n18060) );
  XNOR U16137 ( .A(n18062), .B(n18063), .Z(n15219) );
  AND U16138 ( .A(n18062), .B(n18064), .Z(n18063) );
  XNOR U16139 ( .A(n18065), .B(n18066), .Z(n15222) );
  AND U16140 ( .A(n18065), .B(n18067), .Z(n18066) );
  XNOR U16141 ( .A(n18068), .B(n18069), .Z(n15225) );
  AND U16142 ( .A(n18068), .B(n18070), .Z(n18069) );
  XNOR U16143 ( .A(n18071), .B(n18072), .Z(n15228) );
  AND U16144 ( .A(n18071), .B(n18073), .Z(n18072) );
  XNOR U16145 ( .A(n18074), .B(n18075), .Z(n15231) );
  AND U16146 ( .A(n18074), .B(n18076), .Z(n18075) );
  XNOR U16147 ( .A(n18077), .B(n18078), .Z(n15234) );
  AND U16148 ( .A(n18077), .B(n18079), .Z(n18078) );
  XNOR U16149 ( .A(n18080), .B(n18081), .Z(n15237) );
  AND U16150 ( .A(n18080), .B(n18082), .Z(n18081) );
  XNOR U16151 ( .A(n18083), .B(n18084), .Z(n15240) );
  AND U16152 ( .A(n18083), .B(n18085), .Z(n18084) );
  XNOR U16153 ( .A(n18086), .B(n18087), .Z(n15243) );
  AND U16154 ( .A(n18086), .B(n18088), .Z(n18087) );
  XNOR U16155 ( .A(n18089), .B(n18090), .Z(n15246) );
  AND U16156 ( .A(n18089), .B(n18091), .Z(n18090) );
  XNOR U16157 ( .A(n18092), .B(n18093), .Z(n15249) );
  AND U16158 ( .A(n18092), .B(n18094), .Z(n18093) );
  XNOR U16159 ( .A(n18095), .B(n18096), .Z(n15252) );
  AND U16160 ( .A(n18095), .B(n18097), .Z(n18096) );
  XNOR U16161 ( .A(n18098), .B(n18099), .Z(n15255) );
  AND U16162 ( .A(n18098), .B(n18100), .Z(n18099) );
  XNOR U16163 ( .A(n18101), .B(n18102), .Z(n15258) );
  AND U16164 ( .A(n18101), .B(n18103), .Z(n18102) );
  XNOR U16165 ( .A(n18104), .B(n18105), .Z(n15261) );
  AND U16166 ( .A(n18104), .B(n18106), .Z(n18105) );
  XNOR U16167 ( .A(n18107), .B(n18108), .Z(n15264) );
  AND U16168 ( .A(n18107), .B(n18109), .Z(n18108) );
  XNOR U16169 ( .A(n18110), .B(n18111), .Z(n15267) );
  AND U16170 ( .A(n18110), .B(n18112), .Z(n18111) );
  XNOR U16171 ( .A(n18113), .B(n18114), .Z(n15270) );
  AND U16172 ( .A(n18113), .B(n18115), .Z(n18114) );
  XNOR U16173 ( .A(n18116), .B(n18117), .Z(n15273) );
  AND U16174 ( .A(n18116), .B(n18118), .Z(n18117) );
  XNOR U16175 ( .A(n18119), .B(n18120), .Z(n15276) );
  AND U16176 ( .A(n18119), .B(n18121), .Z(n18120) );
  XNOR U16177 ( .A(n18122), .B(n18123), .Z(n15279) );
  AND U16178 ( .A(n18122), .B(n18124), .Z(n18123) );
  XNOR U16179 ( .A(n18125), .B(n18126), .Z(n15282) );
  AND U16180 ( .A(n18125), .B(n18127), .Z(n18126) );
  XNOR U16181 ( .A(n18128), .B(n18129), .Z(n15285) );
  AND U16182 ( .A(n18128), .B(n18130), .Z(n18129) );
  XNOR U16183 ( .A(n18131), .B(n18132), .Z(n15288) );
  AND U16184 ( .A(n18131), .B(n18133), .Z(n18132) );
  XNOR U16185 ( .A(n18134), .B(n18135), .Z(n15291) );
  AND U16186 ( .A(n18134), .B(n18136), .Z(n18135) );
  XNOR U16187 ( .A(n18137), .B(n18138), .Z(n15294) );
  AND U16188 ( .A(n18137), .B(n18139), .Z(n18138) );
  XNOR U16189 ( .A(n18140), .B(n18141), .Z(n15297) );
  AND U16190 ( .A(n18140), .B(n18142), .Z(n18141) );
  XNOR U16191 ( .A(n18143), .B(n18144), .Z(n15300) );
  AND U16192 ( .A(n18143), .B(n18145), .Z(n18144) );
  XNOR U16193 ( .A(n18146), .B(n18147), .Z(n15303) );
  AND U16194 ( .A(n18146), .B(n18148), .Z(n18147) );
  XNOR U16195 ( .A(n18149), .B(n18150), .Z(n15306) );
  AND U16196 ( .A(n18149), .B(n18151), .Z(n18150) );
  XNOR U16197 ( .A(n18152), .B(n18153), .Z(n15309) );
  AND U16198 ( .A(n18152), .B(n18154), .Z(n18153) );
  XNOR U16199 ( .A(n18155), .B(n18156), .Z(n15312) );
  AND U16200 ( .A(n18155), .B(n18157), .Z(n18156) );
  XNOR U16201 ( .A(n18158), .B(n18159), .Z(n15315) );
  AND U16202 ( .A(n18158), .B(n18160), .Z(n18159) );
  XNOR U16203 ( .A(n18161), .B(n18162), .Z(n15318) );
  AND U16204 ( .A(n18161), .B(n18163), .Z(n18162) );
  XNOR U16205 ( .A(n18164), .B(n18165), .Z(n15321) );
  AND U16206 ( .A(n18164), .B(n18166), .Z(n18165) );
  XNOR U16207 ( .A(n18167), .B(n18168), .Z(n15324) );
  AND U16208 ( .A(n18167), .B(n18169), .Z(n18168) );
  XNOR U16209 ( .A(n18170), .B(n18171), .Z(n15327) );
  AND U16210 ( .A(n18170), .B(n18172), .Z(n18171) );
  XNOR U16211 ( .A(n18173), .B(n18174), .Z(n15330) );
  AND U16212 ( .A(n18173), .B(n18175), .Z(n18174) );
  XNOR U16213 ( .A(n18176), .B(n18177), .Z(n15333) );
  AND U16214 ( .A(n18176), .B(n18178), .Z(n18177) );
  XNOR U16215 ( .A(n18179), .B(n18180), .Z(n15336) );
  AND U16216 ( .A(n18179), .B(n18181), .Z(n18180) );
  XNOR U16217 ( .A(n18182), .B(n18183), .Z(n15339) );
  AND U16218 ( .A(n18182), .B(n18184), .Z(n18183) );
  XNOR U16219 ( .A(n18185), .B(n18186), .Z(n15342) );
  AND U16220 ( .A(n18185), .B(n18187), .Z(n18186) );
  XNOR U16221 ( .A(n18188), .B(n18189), .Z(n15345) );
  AND U16222 ( .A(n18188), .B(n18190), .Z(n18189) );
  XNOR U16223 ( .A(n18191), .B(n18192), .Z(n15348) );
  AND U16224 ( .A(n18191), .B(n18193), .Z(n18192) );
  XNOR U16225 ( .A(n18194), .B(n18195), .Z(n15351) );
  AND U16226 ( .A(n18194), .B(n18196), .Z(n18195) );
  XNOR U16227 ( .A(n18197), .B(n18198), .Z(n15354) );
  AND U16228 ( .A(n18197), .B(n18199), .Z(n18198) );
  XNOR U16229 ( .A(n18200), .B(n18201), .Z(n15357) );
  AND U16230 ( .A(n18200), .B(n18202), .Z(n18201) );
  XNOR U16231 ( .A(n18203), .B(n18204), .Z(n15360) );
  AND U16232 ( .A(n18203), .B(n18205), .Z(n18204) );
  XNOR U16233 ( .A(n18206), .B(n18207), .Z(n15363) );
  AND U16234 ( .A(n18206), .B(n18208), .Z(n18207) );
  XNOR U16235 ( .A(n18209), .B(n18210), .Z(n15366) );
  AND U16236 ( .A(n18209), .B(n18211), .Z(n18210) );
  XNOR U16237 ( .A(n18212), .B(n18213), .Z(n15369) );
  AND U16238 ( .A(n18212), .B(n18214), .Z(n18213) );
  XNOR U16239 ( .A(n18215), .B(n18216), .Z(n15372) );
  AND U16240 ( .A(n18215), .B(n18217), .Z(n18216) );
  XNOR U16241 ( .A(n18218), .B(n18219), .Z(n15375) );
  AND U16242 ( .A(n18218), .B(n18220), .Z(n18219) );
  XNOR U16243 ( .A(n18221), .B(n18222), .Z(n15378) );
  AND U16244 ( .A(n18221), .B(n18223), .Z(n18222) );
  XNOR U16245 ( .A(n18224), .B(n18225), .Z(n15381) );
  AND U16246 ( .A(n18224), .B(n18226), .Z(n18225) );
  XNOR U16247 ( .A(n18227), .B(n18228), .Z(n15384) );
  AND U16248 ( .A(n18227), .B(n18229), .Z(n18228) );
  XNOR U16249 ( .A(n18230), .B(n18231), .Z(n15387) );
  AND U16250 ( .A(n18230), .B(n18232), .Z(n18231) );
  XNOR U16251 ( .A(n18233), .B(n18234), .Z(n15390) );
  AND U16252 ( .A(n18233), .B(n18235), .Z(n18234) );
  XNOR U16253 ( .A(n18236), .B(n18237), .Z(n15393) );
  AND U16254 ( .A(n18236), .B(n18238), .Z(n18237) );
  XNOR U16255 ( .A(n18239), .B(n18240), .Z(n15396) );
  AND U16256 ( .A(n18239), .B(n18241), .Z(n18240) );
  XNOR U16257 ( .A(n18242), .B(n18243), .Z(n15399) );
  AND U16258 ( .A(n18242), .B(n18244), .Z(n18243) );
  XNOR U16259 ( .A(n18245), .B(n18246), .Z(n15402) );
  AND U16260 ( .A(n18245), .B(n18247), .Z(n18246) );
  XNOR U16261 ( .A(n18248), .B(n18249), .Z(n15405) );
  AND U16262 ( .A(n18248), .B(n18250), .Z(n18249) );
  XNOR U16263 ( .A(n18251), .B(n18252), .Z(n15408) );
  AND U16264 ( .A(n18251), .B(n18253), .Z(n18252) );
  XNOR U16265 ( .A(n18254), .B(n18255), .Z(n15411) );
  AND U16266 ( .A(n18254), .B(n18256), .Z(n18255) );
  XNOR U16267 ( .A(n18257), .B(n18258), .Z(n15414) );
  AND U16268 ( .A(n18257), .B(n18259), .Z(n18258) );
  XNOR U16269 ( .A(n18260), .B(n18261), .Z(n15417) );
  AND U16270 ( .A(n18260), .B(n18262), .Z(n18261) );
  XNOR U16271 ( .A(n18263), .B(n18264), .Z(n15420) );
  AND U16272 ( .A(n18263), .B(n18265), .Z(n18264) );
  XNOR U16273 ( .A(n18266), .B(n18267), .Z(n15423) );
  AND U16274 ( .A(n18266), .B(n18268), .Z(n18267) );
  XNOR U16275 ( .A(n18269), .B(n18270), .Z(n15426) );
  AND U16276 ( .A(n18269), .B(n18271), .Z(n18270) );
  XNOR U16277 ( .A(n18272), .B(n18273), .Z(n15429) );
  AND U16278 ( .A(n18272), .B(n18274), .Z(n18273) );
  XNOR U16279 ( .A(n18275), .B(n18276), .Z(n15432) );
  AND U16280 ( .A(n18275), .B(n18277), .Z(n18276) );
  XNOR U16281 ( .A(n18278), .B(n18279), .Z(n15435) );
  AND U16282 ( .A(n18278), .B(n18280), .Z(n18279) );
  XNOR U16283 ( .A(n18281), .B(n18282), .Z(n15438) );
  AND U16284 ( .A(n18281), .B(n18283), .Z(n18282) );
  XNOR U16285 ( .A(n18284), .B(n18285), .Z(n15441) );
  AND U16286 ( .A(n18284), .B(n18286), .Z(n18285) );
  XNOR U16287 ( .A(n18287), .B(n18288), .Z(n15444) );
  AND U16288 ( .A(n18287), .B(n18289), .Z(n18288) );
  XNOR U16289 ( .A(n18290), .B(n18291), .Z(n15447) );
  AND U16290 ( .A(n18290), .B(n18292), .Z(n18291) );
  XNOR U16291 ( .A(n18293), .B(n18294), .Z(n15450) );
  AND U16292 ( .A(n18293), .B(n18295), .Z(n18294) );
  XNOR U16293 ( .A(n18296), .B(n18297), .Z(n15453) );
  AND U16294 ( .A(n18296), .B(n18298), .Z(n18297) );
  XNOR U16295 ( .A(n18299), .B(n18300), .Z(n15456) );
  AND U16296 ( .A(n18299), .B(n18301), .Z(n18300) );
  XNOR U16297 ( .A(n18302), .B(n18303), .Z(n15459) );
  AND U16298 ( .A(n18302), .B(n18304), .Z(n18303) );
  XNOR U16299 ( .A(n18305), .B(n18306), .Z(n15462) );
  AND U16300 ( .A(n18305), .B(n18307), .Z(n18306) );
  XNOR U16301 ( .A(n18308), .B(n18309), .Z(n15465) );
  AND U16302 ( .A(n18308), .B(n18310), .Z(n18309) );
  XNOR U16303 ( .A(n18311), .B(n18312), .Z(n15468) );
  AND U16304 ( .A(n18311), .B(n18313), .Z(n18312) );
  XNOR U16305 ( .A(n18314), .B(n18315), .Z(n15471) );
  AND U16306 ( .A(n18314), .B(n18316), .Z(n18315) );
  XNOR U16307 ( .A(n18317), .B(n18318), .Z(n15474) );
  AND U16308 ( .A(n18317), .B(n18319), .Z(n18318) );
  XNOR U16309 ( .A(n18320), .B(n18321), .Z(n15477) );
  AND U16310 ( .A(n18320), .B(n18322), .Z(n18321) );
  XNOR U16311 ( .A(n18323), .B(n18324), .Z(n15480) );
  AND U16312 ( .A(n18323), .B(n18325), .Z(n18324) );
  XNOR U16313 ( .A(n18326), .B(n18327), .Z(n15483) );
  AND U16314 ( .A(n18326), .B(n18328), .Z(n18327) );
  XNOR U16315 ( .A(n18329), .B(n18330), .Z(n15486) );
  AND U16316 ( .A(n18329), .B(n18331), .Z(n18330) );
  XNOR U16317 ( .A(n18332), .B(n18333), .Z(n15489) );
  AND U16318 ( .A(n18332), .B(n18334), .Z(n18333) );
  XNOR U16319 ( .A(n18335), .B(n18336), .Z(n15492) );
  AND U16320 ( .A(n18335), .B(n18337), .Z(n18336) );
  XNOR U16321 ( .A(n18338), .B(n18339), .Z(n15495) );
  AND U16322 ( .A(n18338), .B(n18340), .Z(n18339) );
  XNOR U16323 ( .A(n18341), .B(n18342), .Z(n15498) );
  AND U16324 ( .A(n18341), .B(n18343), .Z(n18342) );
  XNOR U16325 ( .A(n18344), .B(n18345), .Z(n15501) );
  AND U16326 ( .A(n18344), .B(n18346), .Z(n18345) );
  XNOR U16327 ( .A(n18347), .B(n18348), .Z(n15504) );
  AND U16328 ( .A(n18347), .B(n18349), .Z(n18348) );
  XNOR U16329 ( .A(n18350), .B(n18351), .Z(n15507) );
  AND U16330 ( .A(n18350), .B(n18352), .Z(n18351) );
  XNOR U16331 ( .A(n18353), .B(n18354), .Z(n15510) );
  AND U16332 ( .A(n18353), .B(n18355), .Z(n18354) );
  XNOR U16333 ( .A(n18356), .B(n18357), .Z(n15513) );
  AND U16334 ( .A(n18356), .B(n18358), .Z(n18357) );
  XNOR U16335 ( .A(n18359), .B(n18360), .Z(n15516) );
  AND U16336 ( .A(n18359), .B(n18361), .Z(n18360) );
  XNOR U16337 ( .A(n18362), .B(n18363), .Z(n15519) );
  AND U16338 ( .A(n18362), .B(n18364), .Z(n18363) );
  XNOR U16339 ( .A(n18365), .B(n18366), .Z(n15522) );
  AND U16340 ( .A(n18365), .B(n18367), .Z(n18366) );
  XNOR U16341 ( .A(n18368), .B(n18369), .Z(n15525) );
  AND U16342 ( .A(n18368), .B(n18370), .Z(n18369) );
  XNOR U16343 ( .A(n18371), .B(n18372), .Z(n15528) );
  AND U16344 ( .A(n18371), .B(n18373), .Z(n18372) );
  XNOR U16345 ( .A(n18374), .B(n18375), .Z(n15531) );
  AND U16346 ( .A(n18374), .B(n18376), .Z(n18375) );
  XNOR U16347 ( .A(n18377), .B(n18378), .Z(n15534) );
  AND U16348 ( .A(n18377), .B(n18379), .Z(n18378) );
  XNOR U16349 ( .A(n18380), .B(n18381), .Z(n15537) );
  AND U16350 ( .A(n18380), .B(n18382), .Z(n18381) );
  XNOR U16351 ( .A(n18383), .B(n18384), .Z(n15540) );
  AND U16352 ( .A(n18383), .B(n18385), .Z(n18384) );
  XNOR U16353 ( .A(n18386), .B(n18387), .Z(n15543) );
  AND U16354 ( .A(n18386), .B(n18388), .Z(n18387) );
  XNOR U16355 ( .A(n18389), .B(n18390), .Z(n15546) );
  AND U16356 ( .A(n18389), .B(n18391), .Z(n18390) );
  XNOR U16357 ( .A(n18392), .B(n18393), .Z(n15549) );
  AND U16358 ( .A(n18392), .B(n18394), .Z(n18393) );
  XNOR U16359 ( .A(n18395), .B(n18396), .Z(n15552) );
  AND U16360 ( .A(n18395), .B(n18397), .Z(n18396) );
  XNOR U16361 ( .A(n18398), .B(n18399), .Z(n15555) );
  AND U16362 ( .A(n18398), .B(n18400), .Z(n18399) );
  XNOR U16363 ( .A(n18401), .B(n18402), .Z(n15558) );
  AND U16364 ( .A(n18401), .B(n18403), .Z(n18402) );
  XNOR U16365 ( .A(n18404), .B(n18405), .Z(n15561) );
  AND U16366 ( .A(n18404), .B(n18406), .Z(n18405) );
  XNOR U16367 ( .A(n18407), .B(n18408), .Z(n15564) );
  AND U16368 ( .A(n18407), .B(n18409), .Z(n18408) );
  XNOR U16369 ( .A(n18410), .B(n18411), .Z(n15567) );
  AND U16370 ( .A(n18410), .B(n18412), .Z(n18411) );
  XNOR U16371 ( .A(n18413), .B(n18414), .Z(n15570) );
  AND U16372 ( .A(n18413), .B(n18415), .Z(n18414) );
  XNOR U16373 ( .A(n18416), .B(n18417), .Z(n15573) );
  AND U16374 ( .A(n18416), .B(n18418), .Z(n18417) );
  XNOR U16375 ( .A(n18419), .B(n18420), .Z(n15576) );
  AND U16376 ( .A(n18419), .B(n18421), .Z(n18420) );
  XNOR U16377 ( .A(n18422), .B(n18423), .Z(n15579) );
  AND U16378 ( .A(n18422), .B(n18424), .Z(n18423) );
  XNOR U16379 ( .A(n18425), .B(n18426), .Z(n15582) );
  AND U16380 ( .A(n18425), .B(n18427), .Z(n18426) );
  XNOR U16381 ( .A(n18428), .B(n18429), .Z(n15585) );
  AND U16382 ( .A(n18428), .B(n18430), .Z(n18429) );
  XNOR U16383 ( .A(n18431), .B(n18432), .Z(n15588) );
  AND U16384 ( .A(n18431), .B(n18433), .Z(n18432) );
  XOR U16385 ( .A(n18434), .B(n18435), .Z(n15591) );
  AND U16386 ( .A(n18434), .B(n134), .Z(n18435) );
  XNOR U16387 ( .A(n18436), .B(n17015), .Z(n17017) );
  IV U16388 ( .A(n117), .Z(n18436) );
  XOR U16389 ( .A(n17012), .B(n17011), .Z(n117) );
  XNOR U16390 ( .A(n17009), .B(n17008), .Z(n17011) );
  XNOR U16391 ( .A(n17006), .B(n17005), .Z(n17008) );
  XNOR U16392 ( .A(n17003), .B(n17002), .Z(n17005) );
  XNOR U16393 ( .A(n17000), .B(n16999), .Z(n17002) );
  XNOR U16394 ( .A(n16997), .B(n16996), .Z(n16999) );
  XNOR U16395 ( .A(n16994), .B(n16993), .Z(n16996) );
  XNOR U16396 ( .A(n16991), .B(n16990), .Z(n16993) );
  XNOR U16397 ( .A(n16988), .B(n16987), .Z(n16990) );
  XNOR U16398 ( .A(n16985), .B(n16984), .Z(n16987) );
  XNOR U16399 ( .A(n16982), .B(n16981), .Z(n16984) );
  XNOR U16400 ( .A(n16979), .B(n16978), .Z(n16981) );
  XNOR U16401 ( .A(n16976), .B(n16975), .Z(n16978) );
  XNOR U16402 ( .A(n16973), .B(n16972), .Z(n16975) );
  XNOR U16403 ( .A(n16970), .B(n16969), .Z(n16972) );
  XNOR U16404 ( .A(n16967), .B(n16966), .Z(n16969) );
  XNOR U16405 ( .A(n16964), .B(n16963), .Z(n16966) );
  XNOR U16406 ( .A(n16961), .B(n16960), .Z(n16963) );
  XNOR U16407 ( .A(n16958), .B(n16957), .Z(n16960) );
  XNOR U16408 ( .A(n16955), .B(n16954), .Z(n16957) );
  XNOR U16409 ( .A(n16952), .B(n16951), .Z(n16954) );
  XNOR U16410 ( .A(n16949), .B(n16948), .Z(n16951) );
  XNOR U16411 ( .A(n16946), .B(n16945), .Z(n16948) );
  XNOR U16412 ( .A(n16943), .B(n16942), .Z(n16945) );
  XNOR U16413 ( .A(n16940), .B(n16939), .Z(n16942) );
  XNOR U16414 ( .A(n16937), .B(n16936), .Z(n16939) );
  XNOR U16415 ( .A(n16934), .B(n16933), .Z(n16936) );
  XNOR U16416 ( .A(n16931), .B(n16930), .Z(n16933) );
  XNOR U16417 ( .A(n16928), .B(n16927), .Z(n16930) );
  XNOR U16418 ( .A(n16925), .B(n16924), .Z(n16927) );
  XNOR U16419 ( .A(n16922), .B(n16921), .Z(n16924) );
  XNOR U16420 ( .A(n16919), .B(n16918), .Z(n16921) );
  XNOR U16421 ( .A(n16916), .B(n16915), .Z(n16918) );
  XNOR U16422 ( .A(n16913), .B(n16912), .Z(n16915) );
  XNOR U16423 ( .A(n16910), .B(n16909), .Z(n16912) );
  XNOR U16424 ( .A(n16907), .B(n16906), .Z(n16909) );
  XNOR U16425 ( .A(n16904), .B(n16903), .Z(n16906) );
  XNOR U16426 ( .A(n16901), .B(n16900), .Z(n16903) );
  XNOR U16427 ( .A(n16898), .B(n16897), .Z(n16900) );
  XNOR U16428 ( .A(n16895), .B(n16894), .Z(n16897) );
  XNOR U16429 ( .A(n16892), .B(n16891), .Z(n16894) );
  XNOR U16430 ( .A(n16889), .B(n16888), .Z(n16891) );
  XNOR U16431 ( .A(n16886), .B(n16885), .Z(n16888) );
  XNOR U16432 ( .A(n16883), .B(n16882), .Z(n16885) );
  XNOR U16433 ( .A(n16880), .B(n16879), .Z(n16882) );
  XNOR U16434 ( .A(n16877), .B(n16876), .Z(n16879) );
  XNOR U16435 ( .A(n16874), .B(n16873), .Z(n16876) );
  XNOR U16436 ( .A(n16871), .B(n16870), .Z(n16873) );
  XNOR U16437 ( .A(n16868), .B(n16867), .Z(n16870) );
  XNOR U16438 ( .A(n16865), .B(n16864), .Z(n16867) );
  XNOR U16439 ( .A(n16862), .B(n16861), .Z(n16864) );
  XNOR U16440 ( .A(n16859), .B(n16858), .Z(n16861) );
  XNOR U16441 ( .A(n16856), .B(n16855), .Z(n16858) );
  XNOR U16442 ( .A(n16853), .B(n16852), .Z(n16855) );
  XNOR U16443 ( .A(n16850), .B(n16849), .Z(n16852) );
  XNOR U16444 ( .A(n16847), .B(n16846), .Z(n16849) );
  XNOR U16445 ( .A(n16844), .B(n16843), .Z(n16846) );
  XNOR U16446 ( .A(n16841), .B(n16840), .Z(n16843) );
  XNOR U16447 ( .A(n16838), .B(n16837), .Z(n16840) );
  XNOR U16448 ( .A(n16835), .B(n16834), .Z(n16837) );
  XNOR U16449 ( .A(n16832), .B(n16831), .Z(n16834) );
  XNOR U16450 ( .A(n16829), .B(n16828), .Z(n16831) );
  XNOR U16451 ( .A(n16826), .B(n16825), .Z(n16828) );
  XNOR U16452 ( .A(n16823), .B(n16822), .Z(n16825) );
  XNOR U16453 ( .A(n16820), .B(n16819), .Z(n16822) );
  XNOR U16454 ( .A(n16817), .B(n16816), .Z(n16819) );
  XNOR U16455 ( .A(n16814), .B(n16813), .Z(n16816) );
  XNOR U16456 ( .A(n16811), .B(n16810), .Z(n16813) );
  XNOR U16457 ( .A(n16808), .B(n16807), .Z(n16810) );
  XNOR U16458 ( .A(n16805), .B(n16804), .Z(n16807) );
  XNOR U16459 ( .A(n16802), .B(n16801), .Z(n16804) );
  XNOR U16460 ( .A(n16799), .B(n16798), .Z(n16801) );
  XNOR U16461 ( .A(n16796), .B(n16795), .Z(n16798) );
  XNOR U16462 ( .A(n16793), .B(n16792), .Z(n16795) );
  XNOR U16463 ( .A(n16790), .B(n16789), .Z(n16792) );
  XNOR U16464 ( .A(n16787), .B(n16786), .Z(n16789) );
  XNOR U16465 ( .A(n16784), .B(n16783), .Z(n16786) );
  XNOR U16466 ( .A(n16781), .B(n16780), .Z(n16783) );
  XNOR U16467 ( .A(n16778), .B(n16777), .Z(n16780) );
  XNOR U16468 ( .A(n16775), .B(n16774), .Z(n16777) );
  XNOR U16469 ( .A(n16772), .B(n16771), .Z(n16774) );
  XNOR U16470 ( .A(n16769), .B(n16768), .Z(n16771) );
  XNOR U16471 ( .A(n16766), .B(n16765), .Z(n16768) );
  XNOR U16472 ( .A(n16763), .B(n16762), .Z(n16765) );
  XNOR U16473 ( .A(n16760), .B(n16759), .Z(n16762) );
  XNOR U16474 ( .A(n16757), .B(n16756), .Z(n16759) );
  XNOR U16475 ( .A(n16754), .B(n16753), .Z(n16756) );
  XNOR U16476 ( .A(n16751), .B(n16750), .Z(n16753) );
  XNOR U16477 ( .A(n16748), .B(n16747), .Z(n16750) );
  XNOR U16478 ( .A(n16745), .B(n16744), .Z(n16747) );
  XNOR U16479 ( .A(n16742), .B(n16741), .Z(n16744) );
  XNOR U16480 ( .A(n16739), .B(n16738), .Z(n16741) );
  XNOR U16481 ( .A(n16736), .B(n16735), .Z(n16738) );
  XNOR U16482 ( .A(n16733), .B(n16732), .Z(n16735) );
  XNOR U16483 ( .A(n16730), .B(n16729), .Z(n16732) );
  XNOR U16484 ( .A(n16727), .B(n16726), .Z(n16729) );
  XNOR U16485 ( .A(n16724), .B(n16723), .Z(n16726) );
  XNOR U16486 ( .A(n16721), .B(n16720), .Z(n16723) );
  XNOR U16487 ( .A(n16718), .B(n16717), .Z(n16720) );
  XNOR U16488 ( .A(n16715), .B(n16714), .Z(n16717) );
  XNOR U16489 ( .A(n16712), .B(n16711), .Z(n16714) );
  XNOR U16490 ( .A(n16709), .B(n16708), .Z(n16711) );
  XNOR U16491 ( .A(n16706), .B(n16705), .Z(n16708) );
  XNOR U16492 ( .A(n16703), .B(n16702), .Z(n16705) );
  XNOR U16493 ( .A(n16700), .B(n16699), .Z(n16702) );
  XNOR U16494 ( .A(n16697), .B(n16696), .Z(n16699) );
  XNOR U16495 ( .A(n16694), .B(n16693), .Z(n16696) );
  XNOR U16496 ( .A(n16691), .B(n16690), .Z(n16693) );
  XNOR U16497 ( .A(n16688), .B(n16687), .Z(n16690) );
  XNOR U16498 ( .A(n16685), .B(n16684), .Z(n16687) );
  XNOR U16499 ( .A(n16682), .B(n16681), .Z(n16684) );
  XNOR U16500 ( .A(n16679), .B(n16678), .Z(n16681) );
  XNOR U16501 ( .A(n16676), .B(n16675), .Z(n16678) );
  XNOR U16502 ( .A(n16673), .B(n16672), .Z(n16675) );
  XNOR U16503 ( .A(n16670), .B(n16669), .Z(n16672) );
  XNOR U16504 ( .A(n16667), .B(n16666), .Z(n16669) );
  XNOR U16505 ( .A(n16664), .B(n16663), .Z(n16666) );
  XNOR U16506 ( .A(n16661), .B(n16660), .Z(n16663) );
  XNOR U16507 ( .A(n16658), .B(n16657), .Z(n16660) );
  XNOR U16508 ( .A(n16655), .B(n16654), .Z(n16657) );
  XNOR U16509 ( .A(n16652), .B(n16651), .Z(n16654) );
  XNOR U16510 ( .A(n16649), .B(n16648), .Z(n16651) );
  XNOR U16511 ( .A(n16646), .B(n16645), .Z(n16648) );
  XNOR U16512 ( .A(n16643), .B(n16642), .Z(n16645) );
  XNOR U16513 ( .A(n16640), .B(n16639), .Z(n16642) );
  XNOR U16514 ( .A(n16637), .B(n16636), .Z(n16639) );
  XNOR U16515 ( .A(n16634), .B(n16633), .Z(n16636) );
  XNOR U16516 ( .A(n16631), .B(n16630), .Z(n16633) );
  XNOR U16517 ( .A(n16628), .B(n16627), .Z(n16630) );
  XNOR U16518 ( .A(n16625), .B(n16624), .Z(n16627) );
  XNOR U16519 ( .A(n16622), .B(n16621), .Z(n16624) );
  XNOR U16520 ( .A(n16619), .B(n16618), .Z(n16621) );
  XNOR U16521 ( .A(n16616), .B(n16615), .Z(n16618) );
  XNOR U16522 ( .A(n16613), .B(n16612), .Z(n16615) );
  XNOR U16523 ( .A(n16610), .B(n16609), .Z(n16612) );
  XNOR U16524 ( .A(n16607), .B(n16606), .Z(n16609) );
  XNOR U16525 ( .A(n16604), .B(n16603), .Z(n16606) );
  XNOR U16526 ( .A(n16601), .B(n16600), .Z(n16603) );
  XNOR U16527 ( .A(n16598), .B(n16597), .Z(n16600) );
  XNOR U16528 ( .A(n16595), .B(n16594), .Z(n16597) );
  XNOR U16529 ( .A(n16592), .B(n16591), .Z(n16594) );
  XNOR U16530 ( .A(n16589), .B(n16588), .Z(n16591) );
  XNOR U16531 ( .A(n16586), .B(n16585), .Z(n16588) );
  XNOR U16532 ( .A(n16583), .B(n16582), .Z(n16585) );
  XNOR U16533 ( .A(n16580), .B(n16579), .Z(n16582) );
  XNOR U16534 ( .A(n16577), .B(n16576), .Z(n16579) );
  XNOR U16535 ( .A(n16574), .B(n16573), .Z(n16576) );
  XNOR U16536 ( .A(n16571), .B(n16570), .Z(n16573) );
  XNOR U16537 ( .A(n16568), .B(n16567), .Z(n16570) );
  XNOR U16538 ( .A(n16565), .B(n16564), .Z(n16567) );
  XNOR U16539 ( .A(n16562), .B(n16561), .Z(n16564) );
  XNOR U16540 ( .A(n16559), .B(n16558), .Z(n16561) );
  XNOR U16541 ( .A(n16556), .B(n16555), .Z(n16558) );
  XNOR U16542 ( .A(n16553), .B(n16552), .Z(n16555) );
  XNOR U16543 ( .A(n16550), .B(n16549), .Z(n16552) );
  XNOR U16544 ( .A(n16547), .B(n16546), .Z(n16549) );
  XNOR U16545 ( .A(n16544), .B(n16543), .Z(n16546) );
  XNOR U16546 ( .A(n16541), .B(n16540), .Z(n16543) );
  XNOR U16547 ( .A(n16538), .B(n16537), .Z(n16540) );
  XNOR U16548 ( .A(n16535), .B(n16534), .Z(n16537) );
  XNOR U16549 ( .A(n16532), .B(n16531), .Z(n16534) );
  XNOR U16550 ( .A(n16529), .B(n16528), .Z(n16531) );
  XNOR U16551 ( .A(n16526), .B(n16525), .Z(n16528) );
  XNOR U16552 ( .A(n16523), .B(n16522), .Z(n16525) );
  XNOR U16553 ( .A(n16520), .B(n16519), .Z(n16522) );
  XNOR U16554 ( .A(n16517), .B(n16516), .Z(n16519) );
  XNOR U16555 ( .A(n16514), .B(n16513), .Z(n16516) );
  XNOR U16556 ( .A(n16511), .B(n16510), .Z(n16513) );
  XNOR U16557 ( .A(n16508), .B(n16507), .Z(n16510) );
  XNOR U16558 ( .A(n16505), .B(n16504), .Z(n16507) );
  XNOR U16559 ( .A(n16502), .B(n16501), .Z(n16504) );
  XNOR U16560 ( .A(n16499), .B(n16498), .Z(n16501) );
  XNOR U16561 ( .A(n16496), .B(n16495), .Z(n16498) );
  XNOR U16562 ( .A(n16493), .B(n16492), .Z(n16495) );
  XNOR U16563 ( .A(n16490), .B(n16489), .Z(n16492) );
  XNOR U16564 ( .A(n16487), .B(n16486), .Z(n16489) );
  XNOR U16565 ( .A(n16484), .B(n16483), .Z(n16486) );
  XNOR U16566 ( .A(n16481), .B(n16480), .Z(n16483) );
  XNOR U16567 ( .A(n16478), .B(n16477), .Z(n16480) );
  XNOR U16568 ( .A(n16475), .B(n16474), .Z(n16477) );
  XNOR U16569 ( .A(n16472), .B(n16471), .Z(n16474) );
  XNOR U16570 ( .A(n16469), .B(n16468), .Z(n16471) );
  XNOR U16571 ( .A(n16466), .B(n16465), .Z(n16468) );
  XNOR U16572 ( .A(n16463), .B(n16462), .Z(n16465) );
  XNOR U16573 ( .A(n16460), .B(n16459), .Z(n16462) );
  XNOR U16574 ( .A(n16457), .B(n16456), .Z(n16459) );
  XNOR U16575 ( .A(n16454), .B(n16453), .Z(n16456) );
  XNOR U16576 ( .A(n16451), .B(n16450), .Z(n16453) );
  XNOR U16577 ( .A(n16448), .B(n16447), .Z(n16450) );
  XNOR U16578 ( .A(n16445), .B(n16444), .Z(n16447) );
  XNOR U16579 ( .A(n16442), .B(n16441), .Z(n16444) );
  XNOR U16580 ( .A(n16439), .B(n16438), .Z(n16441) );
  XNOR U16581 ( .A(n16436), .B(n16435), .Z(n16438) );
  XNOR U16582 ( .A(n16433), .B(n16432), .Z(n16435) );
  XNOR U16583 ( .A(n16430), .B(n16429), .Z(n16432) );
  XNOR U16584 ( .A(n16427), .B(n16426), .Z(n16429) );
  XNOR U16585 ( .A(n16424), .B(n16423), .Z(n16426) );
  XNOR U16586 ( .A(n16421), .B(n16420), .Z(n16423) );
  XNOR U16587 ( .A(n16418), .B(n16417), .Z(n16420) );
  XNOR U16588 ( .A(n16415), .B(n16414), .Z(n16417) );
  XNOR U16589 ( .A(n16412), .B(n16411), .Z(n16414) );
  XNOR U16590 ( .A(n16409), .B(n16408), .Z(n16411) );
  XNOR U16591 ( .A(n16406), .B(n16405), .Z(n16408) );
  XNOR U16592 ( .A(n16403), .B(n16402), .Z(n16405) );
  XNOR U16593 ( .A(n16400), .B(n16399), .Z(n16402) );
  XNOR U16594 ( .A(n16397), .B(n16396), .Z(n16399) );
  XNOR U16595 ( .A(n16394), .B(n16393), .Z(n16396) );
  XNOR U16596 ( .A(n16391), .B(n16390), .Z(n16393) );
  XNOR U16597 ( .A(n16388), .B(n16387), .Z(n16390) );
  XNOR U16598 ( .A(n16385), .B(n16384), .Z(n16387) );
  XNOR U16599 ( .A(n16382), .B(n16381), .Z(n16384) );
  XNOR U16600 ( .A(n16379), .B(n16378), .Z(n16381) );
  XNOR U16601 ( .A(n16376), .B(n16375), .Z(n16378) );
  XNOR U16602 ( .A(n16373), .B(n16372), .Z(n16375) );
  XNOR U16603 ( .A(n16370), .B(n16369), .Z(n16372) );
  XNOR U16604 ( .A(n16367), .B(n16366), .Z(n16369) );
  XNOR U16605 ( .A(n16364), .B(n16363), .Z(n16366) );
  XNOR U16606 ( .A(n16361), .B(n16360), .Z(n16363) );
  XNOR U16607 ( .A(n16358), .B(n16357), .Z(n16360) );
  XNOR U16608 ( .A(n16355), .B(n16354), .Z(n16357) );
  XNOR U16609 ( .A(n16352), .B(n16351), .Z(n16354) );
  XNOR U16610 ( .A(n16349), .B(n16348), .Z(n16351) );
  XNOR U16611 ( .A(n16346), .B(n16345), .Z(n16348) );
  XNOR U16612 ( .A(n16343), .B(n16342), .Z(n16345) );
  XNOR U16613 ( .A(n16340), .B(n16339), .Z(n16342) );
  XNOR U16614 ( .A(n16337), .B(n16336), .Z(n16339) );
  XNOR U16615 ( .A(n16334), .B(n16333), .Z(n16336) );
  XNOR U16616 ( .A(n16331), .B(n16330), .Z(n16333) );
  XNOR U16617 ( .A(n16328), .B(n16327), .Z(n16330) );
  XNOR U16618 ( .A(n16325), .B(n16324), .Z(n16327) );
  XNOR U16619 ( .A(n16322), .B(n16321), .Z(n16324) );
  XNOR U16620 ( .A(n16319), .B(n16318), .Z(n16321) );
  XNOR U16621 ( .A(n16316), .B(n16315), .Z(n16318) );
  XNOR U16622 ( .A(n16313), .B(n16312), .Z(n16315) );
  XNOR U16623 ( .A(n16310), .B(n16309), .Z(n16312) );
  XNOR U16624 ( .A(n16307), .B(n16306), .Z(n16309) );
  XNOR U16625 ( .A(n16304), .B(n16303), .Z(n16306) );
  XNOR U16626 ( .A(n16301), .B(n16300), .Z(n16303) );
  XNOR U16627 ( .A(n16298), .B(n16297), .Z(n16300) );
  XNOR U16628 ( .A(n16295), .B(n16294), .Z(n16297) );
  XNOR U16629 ( .A(n16292), .B(n16291), .Z(n16294) );
  XNOR U16630 ( .A(n16289), .B(n16288), .Z(n16291) );
  XNOR U16631 ( .A(n16286), .B(n16285), .Z(n16288) );
  XNOR U16632 ( .A(n16283), .B(n16282), .Z(n16285) );
  XNOR U16633 ( .A(n16280), .B(n16279), .Z(n16282) );
  XNOR U16634 ( .A(n16277), .B(n16276), .Z(n16279) );
  XNOR U16635 ( .A(n16274), .B(n16273), .Z(n16276) );
  XNOR U16636 ( .A(n16271), .B(n16270), .Z(n16273) );
  XNOR U16637 ( .A(n16268), .B(n16267), .Z(n16270) );
  XNOR U16638 ( .A(n16265), .B(n16264), .Z(n16267) );
  XNOR U16639 ( .A(n16262), .B(n16261), .Z(n16264) );
  XNOR U16640 ( .A(n16259), .B(n16258), .Z(n16261) );
  XNOR U16641 ( .A(n16256), .B(n16255), .Z(n16258) );
  XNOR U16642 ( .A(n16253), .B(n16252), .Z(n16255) );
  XNOR U16643 ( .A(n16250), .B(n16249), .Z(n16252) );
  XNOR U16644 ( .A(n16247), .B(n16246), .Z(n16249) );
  XNOR U16645 ( .A(n16244), .B(n16243), .Z(n16246) );
  XNOR U16646 ( .A(n16241), .B(n16240), .Z(n16243) );
  XNOR U16647 ( .A(n16238), .B(n16237), .Z(n16240) );
  XNOR U16648 ( .A(n16235), .B(n16234), .Z(n16237) );
  XNOR U16649 ( .A(n16232), .B(n16231), .Z(n16234) );
  XNOR U16650 ( .A(n16229), .B(n16228), .Z(n16231) );
  XNOR U16651 ( .A(n16226), .B(n16225), .Z(n16228) );
  XNOR U16652 ( .A(n16223), .B(n16222), .Z(n16225) );
  XNOR U16653 ( .A(n16220), .B(n16219), .Z(n16222) );
  XNOR U16654 ( .A(n16217), .B(n16216), .Z(n16219) );
  XNOR U16655 ( .A(n16214), .B(n16213), .Z(n16216) );
  XNOR U16656 ( .A(n16211), .B(n16210), .Z(n16213) );
  XNOR U16657 ( .A(n16208), .B(n16207), .Z(n16210) );
  XNOR U16658 ( .A(n16205), .B(n16204), .Z(n16207) );
  XNOR U16659 ( .A(n16202), .B(n16201), .Z(n16204) );
  XNOR U16660 ( .A(n16199), .B(n16198), .Z(n16201) );
  XNOR U16661 ( .A(n16196), .B(n16195), .Z(n16198) );
  XNOR U16662 ( .A(n16193), .B(n16192), .Z(n16195) );
  XNOR U16663 ( .A(n16190), .B(n16189), .Z(n16192) );
  XNOR U16664 ( .A(n16187), .B(n16186), .Z(n16189) );
  XNOR U16665 ( .A(n16184), .B(n16183), .Z(n16186) );
  XNOR U16666 ( .A(n16181), .B(n16180), .Z(n16183) );
  XNOR U16667 ( .A(n16178), .B(n16177), .Z(n16180) );
  XNOR U16668 ( .A(n16175), .B(n16174), .Z(n16177) );
  XNOR U16669 ( .A(n16172), .B(n16171), .Z(n16174) );
  XNOR U16670 ( .A(n16169), .B(n16168), .Z(n16171) );
  XNOR U16671 ( .A(n16166), .B(n16165), .Z(n16168) );
  XNOR U16672 ( .A(n16163), .B(n16162), .Z(n16165) );
  XNOR U16673 ( .A(n16160), .B(n16159), .Z(n16162) );
  XNOR U16674 ( .A(n16157), .B(n16156), .Z(n16159) );
  XNOR U16675 ( .A(n16154), .B(n16153), .Z(n16156) );
  XNOR U16676 ( .A(n16151), .B(n16150), .Z(n16153) );
  XNOR U16677 ( .A(n16148), .B(n16147), .Z(n16150) );
  XNOR U16678 ( .A(n16145), .B(n16144), .Z(n16147) );
  XNOR U16679 ( .A(n16142), .B(n16141), .Z(n16144) );
  XNOR U16680 ( .A(n16139), .B(n16138), .Z(n16141) );
  XNOR U16681 ( .A(n16136), .B(n16135), .Z(n16138) );
  XNOR U16682 ( .A(n16133), .B(n16132), .Z(n16135) );
  XNOR U16683 ( .A(n16130), .B(n16129), .Z(n16132) );
  XNOR U16684 ( .A(n16127), .B(n16126), .Z(n16129) );
  XNOR U16685 ( .A(n16124), .B(n16123), .Z(n16126) );
  XNOR U16686 ( .A(n16121), .B(n16120), .Z(n16123) );
  XNOR U16687 ( .A(n16118), .B(n16117), .Z(n16120) );
  XNOR U16688 ( .A(n16115), .B(n16114), .Z(n16117) );
  XNOR U16689 ( .A(n16112), .B(n16111), .Z(n16114) );
  XNOR U16690 ( .A(n16109), .B(n16108), .Z(n16111) );
  XNOR U16691 ( .A(n16106), .B(n16105), .Z(n16108) );
  XNOR U16692 ( .A(n16103), .B(n16102), .Z(n16105) );
  XNOR U16693 ( .A(n16100), .B(n16099), .Z(n16102) );
  XNOR U16694 ( .A(n16097), .B(n16096), .Z(n16099) );
  XNOR U16695 ( .A(n16094), .B(n16093), .Z(n16096) );
  XNOR U16696 ( .A(n16091), .B(n16090), .Z(n16093) );
  XNOR U16697 ( .A(n16088), .B(n16087), .Z(n16090) );
  XNOR U16698 ( .A(n16085), .B(n16084), .Z(n16087) );
  XNOR U16699 ( .A(n16082), .B(n16081), .Z(n16084) );
  XNOR U16700 ( .A(n16079), .B(n16078), .Z(n16081) );
  XNOR U16701 ( .A(n16076), .B(n16075), .Z(n16078) );
  XNOR U16702 ( .A(n16073), .B(n16072), .Z(n16075) );
  XNOR U16703 ( .A(n16070), .B(n16069), .Z(n16072) );
  XNOR U16704 ( .A(n16067), .B(n16066), .Z(n16069) );
  XNOR U16705 ( .A(n16064), .B(n16063), .Z(n16066) );
  XNOR U16706 ( .A(n16061), .B(n16060), .Z(n16063) );
  XNOR U16707 ( .A(n16058), .B(n16057), .Z(n16060) );
  XNOR U16708 ( .A(n16055), .B(n16054), .Z(n16057) );
  XNOR U16709 ( .A(n16052), .B(n16051), .Z(n16054) );
  XNOR U16710 ( .A(n16049), .B(n16048), .Z(n16051) );
  XNOR U16711 ( .A(n16046), .B(n16045), .Z(n16048) );
  XNOR U16712 ( .A(n16043), .B(n16042), .Z(n16045) );
  XNOR U16713 ( .A(n16040), .B(n16039), .Z(n16042) );
  XNOR U16714 ( .A(n16037), .B(n16036), .Z(n16039) );
  XNOR U16715 ( .A(n16034), .B(n16033), .Z(n16036) );
  XNOR U16716 ( .A(n16031), .B(n16030), .Z(n16033) );
  XNOR U16717 ( .A(n16028), .B(n16027), .Z(n16030) );
  XNOR U16718 ( .A(n16025), .B(n16024), .Z(n16027) );
  XNOR U16719 ( .A(n16022), .B(n16021), .Z(n16024) );
  XNOR U16720 ( .A(n16019), .B(n16018), .Z(n16021) );
  XNOR U16721 ( .A(n16016), .B(n16015), .Z(n16018) );
  XNOR U16722 ( .A(n16013), .B(n16012), .Z(n16015) );
  XNOR U16723 ( .A(n16010), .B(n16009), .Z(n16012) );
  XNOR U16724 ( .A(n16007), .B(n16006), .Z(n16009) );
  XNOR U16725 ( .A(n16004), .B(n16003), .Z(n16006) );
  XNOR U16726 ( .A(n16001), .B(n16000), .Z(n16003) );
  XNOR U16727 ( .A(n15998), .B(n15997), .Z(n16000) );
  XNOR U16728 ( .A(n15995), .B(n15994), .Z(n15997) );
  XNOR U16729 ( .A(n15992), .B(n15991), .Z(n15994) );
  XNOR U16730 ( .A(n15989), .B(n15988), .Z(n15991) );
  XNOR U16731 ( .A(n15986), .B(n15985), .Z(n15988) );
  XNOR U16732 ( .A(n15983), .B(n15982), .Z(n15985) );
  XNOR U16733 ( .A(n15980), .B(n15979), .Z(n15982) );
  XNOR U16734 ( .A(n15977), .B(n15976), .Z(n15979) );
  XNOR U16735 ( .A(n15974), .B(n15973), .Z(n15976) );
  XNOR U16736 ( .A(n15971), .B(n15970), .Z(n15973) );
  XNOR U16737 ( .A(n15968), .B(n15967), .Z(n15970) );
  XNOR U16738 ( .A(n15965), .B(n15964), .Z(n15967) );
  XNOR U16739 ( .A(n15962), .B(n15961), .Z(n15964) );
  XNOR U16740 ( .A(n15959), .B(n15958), .Z(n15961) );
  XNOR U16741 ( .A(n15956), .B(n15955), .Z(n15958) );
  XNOR U16742 ( .A(n15953), .B(n15952), .Z(n15955) );
  XNOR U16743 ( .A(n15950), .B(n15949), .Z(n15952) );
  XNOR U16744 ( .A(n15947), .B(n15946), .Z(n15949) );
  XNOR U16745 ( .A(n15944), .B(n15943), .Z(n15946) );
  XNOR U16746 ( .A(n15941), .B(n15940), .Z(n15943) );
  XNOR U16747 ( .A(n15938), .B(n15937), .Z(n15940) );
  XNOR U16748 ( .A(n15935), .B(n15934), .Z(n15937) );
  XNOR U16749 ( .A(n15932), .B(n15931), .Z(n15934) );
  XNOR U16750 ( .A(n15929), .B(n15928), .Z(n15931) );
  XNOR U16751 ( .A(n15926), .B(n15925), .Z(n15928) );
  XNOR U16752 ( .A(n15923), .B(n15922), .Z(n15925) );
  XNOR U16753 ( .A(n15920), .B(n15919), .Z(n15922) );
  XNOR U16754 ( .A(n15917), .B(n15916), .Z(n15919) );
  XNOR U16755 ( .A(n15914), .B(n15913), .Z(n15916) );
  XNOR U16756 ( .A(n15911), .B(n15910), .Z(n15913) );
  XNOR U16757 ( .A(n15908), .B(n15907), .Z(n15910) );
  XNOR U16758 ( .A(n15905), .B(n15904), .Z(n15907) );
  XNOR U16759 ( .A(n15902), .B(n15901), .Z(n15904) );
  XNOR U16760 ( .A(n15899), .B(n15898), .Z(n15901) );
  XNOR U16761 ( .A(n15896), .B(n15895), .Z(n15898) );
  XNOR U16762 ( .A(n15893), .B(n15892), .Z(n15895) );
  XNOR U16763 ( .A(n15890), .B(n15889), .Z(n15892) );
  XNOR U16764 ( .A(n15887), .B(n15886), .Z(n15889) );
  XNOR U16765 ( .A(n15884), .B(n15883), .Z(n15886) );
  XNOR U16766 ( .A(n15881), .B(n15880), .Z(n15883) );
  XNOR U16767 ( .A(n15878), .B(n15877), .Z(n15880) );
  XNOR U16768 ( .A(n15875), .B(n15874), .Z(n15877) );
  XNOR U16769 ( .A(n15872), .B(n15871), .Z(n15874) );
  XNOR U16770 ( .A(n15869), .B(n15868), .Z(n15871) );
  XNOR U16771 ( .A(n15866), .B(n15865), .Z(n15868) );
  XNOR U16772 ( .A(n15863), .B(n15862), .Z(n15865) );
  XNOR U16773 ( .A(n15860), .B(n15859), .Z(n15862) );
  XOR U16774 ( .A(n15857), .B(n15856), .Z(n15859) );
  XOR U16775 ( .A(n15854), .B(n15853), .Z(n15856) );
  XOR U16776 ( .A(n15850), .B(n15851), .Z(n15853) );
  AND U16777 ( .A(n18437), .B(n18438), .Z(n15851) );
  XOR U16778 ( .A(n15847), .B(n15848), .Z(n15850) );
  AND U16779 ( .A(n18439), .B(n18440), .Z(n15848) );
  XOR U16780 ( .A(n15844), .B(n15845), .Z(n15847) );
  AND U16781 ( .A(n18441), .B(n18442), .Z(n15845) );
  XNOR U16782 ( .A(n15594), .B(n15842), .Z(n15844) );
  AND U16783 ( .A(n18443), .B(n18444), .Z(n15842) );
  XOR U16784 ( .A(n15596), .B(n15595), .Z(n15594) );
  AND U16785 ( .A(n18445), .B(n18446), .Z(n15595) );
  XOR U16786 ( .A(n15598), .B(n15597), .Z(n15596) );
  AND U16787 ( .A(n18447), .B(n18448), .Z(n15597) );
  XOR U16788 ( .A(n15600), .B(n15599), .Z(n15598) );
  AND U16789 ( .A(n18449), .B(n18450), .Z(n15599) );
  XOR U16790 ( .A(n15602), .B(n15601), .Z(n15600) );
  AND U16791 ( .A(n18451), .B(n18452), .Z(n15601) );
  XOR U16792 ( .A(n15604), .B(n15603), .Z(n15602) );
  AND U16793 ( .A(n18453), .B(n18454), .Z(n15603) );
  XOR U16794 ( .A(n15606), .B(n15605), .Z(n15604) );
  AND U16795 ( .A(n18455), .B(n18456), .Z(n15605) );
  XOR U16796 ( .A(n15608), .B(n15607), .Z(n15606) );
  AND U16797 ( .A(n18457), .B(n18458), .Z(n15607) );
  XOR U16798 ( .A(n15610), .B(n15609), .Z(n15608) );
  AND U16799 ( .A(n18459), .B(n18460), .Z(n15609) );
  XOR U16800 ( .A(n15612), .B(n15611), .Z(n15610) );
  AND U16801 ( .A(n18461), .B(n18462), .Z(n15611) );
  XOR U16802 ( .A(n15614), .B(n15613), .Z(n15612) );
  AND U16803 ( .A(n18463), .B(n18464), .Z(n15613) );
  XOR U16804 ( .A(n15616), .B(n15615), .Z(n15614) );
  AND U16805 ( .A(n18465), .B(n18466), .Z(n15615) );
  XOR U16806 ( .A(n15618), .B(n15617), .Z(n15616) );
  AND U16807 ( .A(n18467), .B(n18468), .Z(n15617) );
  XOR U16808 ( .A(n15620), .B(n15619), .Z(n15618) );
  AND U16809 ( .A(n18469), .B(n18470), .Z(n15619) );
  XOR U16810 ( .A(n15622), .B(n15621), .Z(n15620) );
  AND U16811 ( .A(n18471), .B(n18472), .Z(n15621) );
  XOR U16812 ( .A(n15624), .B(n15623), .Z(n15622) );
  AND U16813 ( .A(n18473), .B(n18474), .Z(n15623) );
  XOR U16814 ( .A(n15626), .B(n15625), .Z(n15624) );
  AND U16815 ( .A(n18475), .B(n18476), .Z(n15625) );
  XOR U16816 ( .A(n15628), .B(n15627), .Z(n15626) );
  AND U16817 ( .A(n18477), .B(n18478), .Z(n15627) );
  XOR U16818 ( .A(n15630), .B(n15629), .Z(n15628) );
  AND U16819 ( .A(n18479), .B(n18480), .Z(n15629) );
  XOR U16820 ( .A(n15632), .B(n15631), .Z(n15630) );
  AND U16821 ( .A(n18481), .B(n18482), .Z(n15631) );
  XOR U16822 ( .A(n15634), .B(n15633), .Z(n15632) );
  AND U16823 ( .A(n18483), .B(n18484), .Z(n15633) );
  XOR U16824 ( .A(n15636), .B(n15635), .Z(n15634) );
  AND U16825 ( .A(n18485), .B(n18486), .Z(n15635) );
  XOR U16826 ( .A(n15638), .B(n15637), .Z(n15636) );
  AND U16827 ( .A(n18487), .B(n18488), .Z(n15637) );
  XOR U16828 ( .A(n15640), .B(n15639), .Z(n15638) );
  AND U16829 ( .A(n18489), .B(n18490), .Z(n15639) );
  XOR U16830 ( .A(n15642), .B(n15641), .Z(n15640) );
  AND U16831 ( .A(n18491), .B(n18492), .Z(n15641) );
  XOR U16832 ( .A(n15644), .B(n15643), .Z(n15642) );
  AND U16833 ( .A(n18493), .B(n18494), .Z(n15643) );
  XOR U16834 ( .A(n15646), .B(n15645), .Z(n15644) );
  AND U16835 ( .A(n18495), .B(n18496), .Z(n15645) );
  XOR U16836 ( .A(n15648), .B(n15647), .Z(n15646) );
  AND U16837 ( .A(n18497), .B(n18498), .Z(n15647) );
  XOR U16838 ( .A(n15650), .B(n15649), .Z(n15648) );
  AND U16839 ( .A(n18499), .B(n18500), .Z(n15649) );
  XOR U16840 ( .A(n15652), .B(n15651), .Z(n15650) );
  AND U16841 ( .A(n18501), .B(n18502), .Z(n15651) );
  XOR U16842 ( .A(n15654), .B(n15653), .Z(n15652) );
  AND U16843 ( .A(n18503), .B(n18504), .Z(n15653) );
  XOR U16844 ( .A(n15656), .B(n15655), .Z(n15654) );
  AND U16845 ( .A(n18505), .B(n18506), .Z(n15655) );
  XOR U16846 ( .A(n15658), .B(n15657), .Z(n15656) );
  AND U16847 ( .A(n18507), .B(n18508), .Z(n15657) );
  XOR U16848 ( .A(n15660), .B(n15659), .Z(n15658) );
  AND U16849 ( .A(n18509), .B(n18510), .Z(n15659) );
  XOR U16850 ( .A(n15662), .B(n15661), .Z(n15660) );
  AND U16851 ( .A(n18511), .B(n18512), .Z(n15661) );
  XOR U16852 ( .A(n15664), .B(n15663), .Z(n15662) );
  AND U16853 ( .A(n18513), .B(n18514), .Z(n15663) );
  XOR U16854 ( .A(n15666), .B(n15665), .Z(n15664) );
  AND U16855 ( .A(n18515), .B(n18516), .Z(n15665) );
  XOR U16856 ( .A(n15668), .B(n15667), .Z(n15666) );
  AND U16857 ( .A(n18517), .B(n18518), .Z(n15667) );
  XOR U16858 ( .A(n15670), .B(n15669), .Z(n15668) );
  AND U16859 ( .A(n18519), .B(n18520), .Z(n15669) );
  XOR U16860 ( .A(n15672), .B(n15671), .Z(n15670) );
  AND U16861 ( .A(n18521), .B(n18522), .Z(n15671) );
  XOR U16862 ( .A(n15674), .B(n15673), .Z(n15672) );
  AND U16863 ( .A(n18523), .B(n18524), .Z(n15673) );
  XOR U16864 ( .A(n15676), .B(n15675), .Z(n15674) );
  AND U16865 ( .A(n18525), .B(n18526), .Z(n15675) );
  XOR U16866 ( .A(n15678), .B(n15677), .Z(n15676) );
  AND U16867 ( .A(n18527), .B(n18528), .Z(n15677) );
  XOR U16868 ( .A(n15680), .B(n15679), .Z(n15678) );
  AND U16869 ( .A(n18529), .B(n18530), .Z(n15679) );
  XOR U16870 ( .A(n15682), .B(n15681), .Z(n15680) );
  AND U16871 ( .A(n18531), .B(n18532), .Z(n15681) );
  XOR U16872 ( .A(n15684), .B(n15683), .Z(n15682) );
  AND U16873 ( .A(n18533), .B(n18534), .Z(n15683) );
  XOR U16874 ( .A(n15686), .B(n15685), .Z(n15684) );
  AND U16875 ( .A(n18535), .B(n18536), .Z(n15685) );
  XOR U16876 ( .A(n15688), .B(n15687), .Z(n15686) );
  AND U16877 ( .A(n18537), .B(n18538), .Z(n15687) );
  XOR U16878 ( .A(n15690), .B(n15689), .Z(n15688) );
  AND U16879 ( .A(n18539), .B(n18540), .Z(n15689) );
  XOR U16880 ( .A(n15692), .B(n15691), .Z(n15690) );
  AND U16881 ( .A(n18541), .B(n18542), .Z(n15691) );
  XOR U16882 ( .A(n15694), .B(n15693), .Z(n15692) );
  AND U16883 ( .A(n18543), .B(n18544), .Z(n15693) );
  XOR U16884 ( .A(n15696), .B(n15695), .Z(n15694) );
  AND U16885 ( .A(n18545), .B(n18546), .Z(n15695) );
  XOR U16886 ( .A(n15698), .B(n15697), .Z(n15696) );
  AND U16887 ( .A(n18547), .B(n18548), .Z(n15697) );
  XOR U16888 ( .A(n15700), .B(n15699), .Z(n15698) );
  AND U16889 ( .A(n18549), .B(n18550), .Z(n15699) );
  XOR U16890 ( .A(n15702), .B(n15701), .Z(n15700) );
  AND U16891 ( .A(n18551), .B(n18552), .Z(n15701) );
  XOR U16892 ( .A(n15704), .B(n15703), .Z(n15702) );
  AND U16893 ( .A(n18553), .B(n18554), .Z(n15703) );
  XOR U16894 ( .A(n15706), .B(n15705), .Z(n15704) );
  AND U16895 ( .A(n18555), .B(n18556), .Z(n15705) );
  XOR U16896 ( .A(n15708), .B(n15707), .Z(n15706) );
  AND U16897 ( .A(n18557), .B(n18558), .Z(n15707) );
  XOR U16898 ( .A(n15710), .B(n15709), .Z(n15708) );
  AND U16899 ( .A(n18559), .B(n18560), .Z(n15709) );
  XOR U16900 ( .A(n15712), .B(n15711), .Z(n15710) );
  AND U16901 ( .A(n18561), .B(n18562), .Z(n15711) );
  XOR U16902 ( .A(n15714), .B(n15713), .Z(n15712) );
  AND U16903 ( .A(n18563), .B(n18564), .Z(n15713) );
  XOR U16904 ( .A(n15716), .B(n15715), .Z(n15714) );
  AND U16905 ( .A(n18565), .B(n18566), .Z(n15715) );
  XOR U16906 ( .A(n15718), .B(n15717), .Z(n15716) );
  AND U16907 ( .A(n18567), .B(n18568), .Z(n15717) );
  XOR U16908 ( .A(n15720), .B(n15719), .Z(n15718) );
  AND U16909 ( .A(n18569), .B(n18570), .Z(n15719) );
  XOR U16910 ( .A(n15722), .B(n15721), .Z(n15720) );
  AND U16911 ( .A(n18571), .B(n18572), .Z(n15721) );
  XOR U16912 ( .A(n15724), .B(n15723), .Z(n15722) );
  AND U16913 ( .A(n18573), .B(n18574), .Z(n15723) );
  XOR U16914 ( .A(n15726), .B(n15725), .Z(n15724) );
  AND U16915 ( .A(n18575), .B(n18576), .Z(n15725) );
  XOR U16916 ( .A(n15728), .B(n15727), .Z(n15726) );
  AND U16917 ( .A(n18577), .B(n18578), .Z(n15727) );
  XOR U16918 ( .A(n15730), .B(n15729), .Z(n15728) );
  AND U16919 ( .A(n18579), .B(n18580), .Z(n15729) );
  XOR U16920 ( .A(n15732), .B(n15731), .Z(n15730) );
  AND U16921 ( .A(n18581), .B(n18582), .Z(n15731) );
  XOR U16922 ( .A(n15734), .B(n15733), .Z(n15732) );
  AND U16923 ( .A(n18583), .B(n18584), .Z(n15733) );
  XOR U16924 ( .A(n15736), .B(n15735), .Z(n15734) );
  AND U16925 ( .A(n18585), .B(n18586), .Z(n15735) );
  XOR U16926 ( .A(n15738), .B(n15737), .Z(n15736) );
  AND U16927 ( .A(n18587), .B(n18588), .Z(n15737) );
  XOR U16928 ( .A(n15740), .B(n15739), .Z(n15738) );
  AND U16929 ( .A(n18589), .B(n18590), .Z(n15739) );
  XOR U16930 ( .A(n15742), .B(n15741), .Z(n15740) );
  AND U16931 ( .A(n18591), .B(n18592), .Z(n15741) );
  XOR U16932 ( .A(n15744), .B(n15743), .Z(n15742) );
  AND U16933 ( .A(n18593), .B(n18594), .Z(n15743) );
  XOR U16934 ( .A(n15746), .B(n15745), .Z(n15744) );
  AND U16935 ( .A(n18595), .B(n18596), .Z(n15745) );
  XOR U16936 ( .A(n15748), .B(n15747), .Z(n15746) );
  AND U16937 ( .A(n18597), .B(n18598), .Z(n15747) );
  XOR U16938 ( .A(n15750), .B(n15749), .Z(n15748) );
  AND U16939 ( .A(n18599), .B(n18600), .Z(n15749) );
  XOR U16940 ( .A(n15752), .B(n15751), .Z(n15750) );
  AND U16941 ( .A(n18601), .B(n18602), .Z(n15751) );
  XOR U16942 ( .A(n15754), .B(n15753), .Z(n15752) );
  AND U16943 ( .A(n18603), .B(n18604), .Z(n15753) );
  XOR U16944 ( .A(n15756), .B(n15755), .Z(n15754) );
  AND U16945 ( .A(n18605), .B(n18606), .Z(n15755) );
  XOR U16946 ( .A(n15758), .B(n15757), .Z(n15756) );
  AND U16947 ( .A(n18607), .B(n18608), .Z(n15757) );
  XOR U16948 ( .A(n15760), .B(n15759), .Z(n15758) );
  AND U16949 ( .A(n18609), .B(n18610), .Z(n15759) );
  XOR U16950 ( .A(n15762), .B(n15761), .Z(n15760) );
  AND U16951 ( .A(n18611), .B(n18612), .Z(n15761) );
  XOR U16952 ( .A(n15764), .B(n15763), .Z(n15762) );
  AND U16953 ( .A(n18613), .B(n18614), .Z(n15763) );
  XOR U16954 ( .A(n15766), .B(n15765), .Z(n15764) );
  AND U16955 ( .A(n18615), .B(n18616), .Z(n15765) );
  XOR U16956 ( .A(n15768), .B(n15767), .Z(n15766) );
  AND U16957 ( .A(n18617), .B(n18618), .Z(n15767) );
  XOR U16958 ( .A(n15770), .B(n15769), .Z(n15768) );
  AND U16959 ( .A(n18619), .B(n18620), .Z(n15769) );
  XOR U16960 ( .A(n15772), .B(n15771), .Z(n15770) );
  AND U16961 ( .A(n18621), .B(n18622), .Z(n15771) );
  XOR U16962 ( .A(n15774), .B(n15773), .Z(n15772) );
  AND U16963 ( .A(n18623), .B(n18624), .Z(n15773) );
  XOR U16964 ( .A(n15776), .B(n15775), .Z(n15774) );
  AND U16965 ( .A(n18625), .B(n18626), .Z(n15775) );
  XOR U16966 ( .A(n15778), .B(n15777), .Z(n15776) );
  AND U16967 ( .A(n18627), .B(n18628), .Z(n15777) );
  XOR U16968 ( .A(n15780), .B(n15779), .Z(n15778) );
  AND U16969 ( .A(n18629), .B(n18630), .Z(n15779) );
  XOR U16970 ( .A(n15782), .B(n15781), .Z(n15780) );
  AND U16971 ( .A(n18631), .B(n18632), .Z(n15781) );
  XOR U16972 ( .A(n15784), .B(n15783), .Z(n15782) );
  AND U16973 ( .A(n18633), .B(n18634), .Z(n15783) );
  XOR U16974 ( .A(n15786), .B(n15785), .Z(n15784) );
  AND U16975 ( .A(n18635), .B(n18636), .Z(n15785) );
  XOR U16976 ( .A(n15838), .B(n15787), .Z(n15786) );
  AND U16977 ( .A(n18637), .B(n18638), .Z(n15787) );
  XOR U16978 ( .A(n15840), .B(n15839), .Z(n15838) );
  AND U16979 ( .A(n18639), .B(n18640), .Z(n15839) );
  XOR U16980 ( .A(n15822), .B(n15841), .Z(n15840) );
  AND U16981 ( .A(n18641), .B(n18642), .Z(n15841) );
  XOR U16982 ( .A(n15824), .B(n15823), .Z(n15822) );
  AND U16983 ( .A(n18643), .B(n18644), .Z(n15823) );
  XOR U16984 ( .A(n15826), .B(n15825), .Z(n15824) );
  AND U16985 ( .A(n18645), .B(n18646), .Z(n15825) );
  XOR U16986 ( .A(n15830), .B(n15827), .Z(n15826) );
  AND U16987 ( .A(n18647), .B(n18648), .Z(n15827) );
  XOR U16988 ( .A(n15832), .B(n15831), .Z(n15830) );
  AND U16989 ( .A(n18649), .B(n18650), .Z(n15831) );
  XOR U16990 ( .A(n15834), .B(n15833), .Z(n15832) );
  AND U16991 ( .A(n18651), .B(n18652), .Z(n15833) );
  XOR U16992 ( .A(n15836), .B(n15835), .Z(n15834) );
  AND U16993 ( .A(n18653), .B(n18654), .Z(n15835) );
  XOR U16994 ( .A(n15811), .B(n15837), .Z(n15836) );
  AND U16995 ( .A(n18655), .B(n18656), .Z(n15837) );
  XNOR U16996 ( .A(n15808), .B(n15812), .Z(n15811) );
  AND U16997 ( .A(n18657), .B(n18658), .Z(n15812) );
  XOR U16998 ( .A(n15807), .B(n15799), .Z(n15808) );
  AND U16999 ( .A(n18659), .B(n18660), .Z(n15799) );
  XNOR U17000 ( .A(n15802), .B(n15798), .Z(n15807) );
  AND U17001 ( .A(n18661), .B(n18662), .Z(n15798) );
  XOR U17002 ( .A(n18663), .B(n18664), .Z(n15802) );
  XOR U17003 ( .A(n15820), .B(n18665), .Z(n18664) );
  XOR U17004 ( .A(n15818), .B(n15816), .Z(n18665) );
  AND U17005 ( .A(n18666), .B(n18667), .Z(n15816) );
  AND U17006 ( .A(n18668), .B(n18669), .Z(n15818) );
  AND U17007 ( .A(n18670), .B(n18671), .Z(n15820) );
  XNOR U17008 ( .A(n18672), .B(n15819), .Z(n18663) );
  XOR U17009 ( .A(n18673), .B(n18674), .Z(n15819) );
  XOR U17010 ( .A(n18675), .B(n18676), .Z(n18674) );
  AND U17011 ( .A(n18677), .B(n18678), .Z(n18676) );
  XNOR U17012 ( .A(n18679), .B(n18680), .Z(n18673) );
  NOR U17013 ( .A(n18681), .B(n18682), .Z(n18680) );
  AND U17014 ( .A(n18683), .B(n18684), .Z(n18682) );
  IV U17015 ( .A(n18685), .Z(n18681) );
  NOR U17016 ( .A(n18675), .B(n18686), .Z(n18685) );
  AND U17017 ( .A(n18687), .B(n18688), .Z(n18686) );
  NOR U17018 ( .A(n18677), .B(n18687), .Z(n18679) );
  XNOR U17019 ( .A(n15821), .B(n15803), .Z(n18672) );
  AND U17020 ( .A(n18689), .B(n18690), .Z(n15803) );
  AND U17021 ( .A(n18691), .B(n18692), .Z(n15821) );
  XOR U17022 ( .A(n18693), .B(n18694), .Z(n15854) );
  NOR U17023 ( .A(n18695), .B(n18696), .Z(n18694) );
  IV U17024 ( .A(n18693), .Z(n18695) );
  XOR U17025 ( .A(n18697), .B(n18698), .Z(n15857) );
  NOR U17026 ( .A(n18697), .B(n18699), .Z(n18698) );
  XNOR U17027 ( .A(n18700), .B(n18701), .Z(n15860) );
  AND U17028 ( .A(n18700), .B(n18702), .Z(n18701) );
  XNOR U17029 ( .A(n18703), .B(n18704), .Z(n15863) );
  AND U17030 ( .A(n18703), .B(n18705), .Z(n18704) );
  XNOR U17031 ( .A(n18706), .B(n18707), .Z(n15866) );
  AND U17032 ( .A(n18706), .B(n18708), .Z(n18707) );
  XNOR U17033 ( .A(n18709), .B(n18710), .Z(n15869) );
  AND U17034 ( .A(n18709), .B(n18711), .Z(n18710) );
  XNOR U17035 ( .A(n18712), .B(n18713), .Z(n15872) );
  AND U17036 ( .A(n18712), .B(n18714), .Z(n18713) );
  XNOR U17037 ( .A(n18715), .B(n18716), .Z(n15875) );
  AND U17038 ( .A(n18715), .B(n18717), .Z(n18716) );
  XNOR U17039 ( .A(n18718), .B(n18719), .Z(n15878) );
  AND U17040 ( .A(n18718), .B(n18720), .Z(n18719) );
  XNOR U17041 ( .A(n18721), .B(n18722), .Z(n15881) );
  AND U17042 ( .A(n18721), .B(n18723), .Z(n18722) );
  XNOR U17043 ( .A(n18724), .B(n18725), .Z(n15884) );
  AND U17044 ( .A(n18724), .B(n18726), .Z(n18725) );
  XNOR U17045 ( .A(n18727), .B(n18728), .Z(n15887) );
  AND U17046 ( .A(n18727), .B(n18729), .Z(n18728) );
  XNOR U17047 ( .A(n18730), .B(n18731), .Z(n15890) );
  AND U17048 ( .A(n18730), .B(n18732), .Z(n18731) );
  XNOR U17049 ( .A(n18733), .B(n18734), .Z(n15893) );
  AND U17050 ( .A(n18733), .B(n18735), .Z(n18734) );
  XNOR U17051 ( .A(n18736), .B(n18737), .Z(n15896) );
  AND U17052 ( .A(n18736), .B(n18738), .Z(n18737) );
  XNOR U17053 ( .A(n18739), .B(n18740), .Z(n15899) );
  AND U17054 ( .A(n18739), .B(n18741), .Z(n18740) );
  XNOR U17055 ( .A(n18742), .B(n18743), .Z(n15902) );
  AND U17056 ( .A(n18742), .B(n18744), .Z(n18743) );
  XNOR U17057 ( .A(n18745), .B(n18746), .Z(n15905) );
  AND U17058 ( .A(n18745), .B(n18747), .Z(n18746) );
  XNOR U17059 ( .A(n18748), .B(n18749), .Z(n15908) );
  AND U17060 ( .A(n18748), .B(n18750), .Z(n18749) );
  XNOR U17061 ( .A(n18751), .B(n18752), .Z(n15911) );
  AND U17062 ( .A(n18751), .B(n18753), .Z(n18752) );
  XNOR U17063 ( .A(n18754), .B(n18755), .Z(n15914) );
  AND U17064 ( .A(n18754), .B(n18756), .Z(n18755) );
  XNOR U17065 ( .A(n18757), .B(n18758), .Z(n15917) );
  AND U17066 ( .A(n18757), .B(n18759), .Z(n18758) );
  XNOR U17067 ( .A(n18760), .B(n18761), .Z(n15920) );
  AND U17068 ( .A(n18760), .B(n18762), .Z(n18761) );
  XNOR U17069 ( .A(n18763), .B(n18764), .Z(n15923) );
  AND U17070 ( .A(n18763), .B(n18765), .Z(n18764) );
  XNOR U17071 ( .A(n18766), .B(n18767), .Z(n15926) );
  AND U17072 ( .A(n18766), .B(n18768), .Z(n18767) );
  XNOR U17073 ( .A(n18769), .B(n18770), .Z(n15929) );
  AND U17074 ( .A(n18769), .B(n18771), .Z(n18770) );
  XNOR U17075 ( .A(n18772), .B(n18773), .Z(n15932) );
  AND U17076 ( .A(n18772), .B(n18774), .Z(n18773) );
  XNOR U17077 ( .A(n18775), .B(n18776), .Z(n15935) );
  AND U17078 ( .A(n18775), .B(n18777), .Z(n18776) );
  XNOR U17079 ( .A(n18778), .B(n18779), .Z(n15938) );
  AND U17080 ( .A(n18778), .B(n18780), .Z(n18779) );
  XNOR U17081 ( .A(n18781), .B(n18782), .Z(n15941) );
  AND U17082 ( .A(n18781), .B(n18783), .Z(n18782) );
  XNOR U17083 ( .A(n18784), .B(n18785), .Z(n15944) );
  AND U17084 ( .A(n18784), .B(n18786), .Z(n18785) );
  XNOR U17085 ( .A(n18787), .B(n18788), .Z(n15947) );
  AND U17086 ( .A(n18787), .B(n18789), .Z(n18788) );
  XNOR U17087 ( .A(n18790), .B(n18791), .Z(n15950) );
  AND U17088 ( .A(n18790), .B(n18792), .Z(n18791) );
  XNOR U17089 ( .A(n18793), .B(n18794), .Z(n15953) );
  AND U17090 ( .A(n18793), .B(n18795), .Z(n18794) );
  XNOR U17091 ( .A(n18796), .B(n18797), .Z(n15956) );
  AND U17092 ( .A(n18796), .B(n18798), .Z(n18797) );
  XNOR U17093 ( .A(n18799), .B(n18800), .Z(n15959) );
  AND U17094 ( .A(n18799), .B(n18801), .Z(n18800) );
  XNOR U17095 ( .A(n18802), .B(n18803), .Z(n15962) );
  AND U17096 ( .A(n18802), .B(n18804), .Z(n18803) );
  XNOR U17097 ( .A(n18805), .B(n18806), .Z(n15965) );
  AND U17098 ( .A(n18805), .B(n18807), .Z(n18806) );
  XNOR U17099 ( .A(n18808), .B(n18809), .Z(n15968) );
  AND U17100 ( .A(n18808), .B(n18810), .Z(n18809) );
  XNOR U17101 ( .A(n18811), .B(n18812), .Z(n15971) );
  AND U17102 ( .A(n18811), .B(n18813), .Z(n18812) );
  XNOR U17103 ( .A(n18814), .B(n18815), .Z(n15974) );
  AND U17104 ( .A(n18814), .B(n18816), .Z(n18815) );
  XNOR U17105 ( .A(n18817), .B(n18818), .Z(n15977) );
  AND U17106 ( .A(n18817), .B(n18819), .Z(n18818) );
  XNOR U17107 ( .A(n18820), .B(n18821), .Z(n15980) );
  AND U17108 ( .A(n18820), .B(n18822), .Z(n18821) );
  XNOR U17109 ( .A(n18823), .B(n18824), .Z(n15983) );
  AND U17110 ( .A(n18823), .B(n18825), .Z(n18824) );
  XNOR U17111 ( .A(n18826), .B(n18827), .Z(n15986) );
  AND U17112 ( .A(n18826), .B(n18828), .Z(n18827) );
  XNOR U17113 ( .A(n18829), .B(n18830), .Z(n15989) );
  AND U17114 ( .A(n18829), .B(n18831), .Z(n18830) );
  XNOR U17115 ( .A(n18832), .B(n18833), .Z(n15992) );
  AND U17116 ( .A(n18832), .B(n18834), .Z(n18833) );
  XNOR U17117 ( .A(n18835), .B(n18836), .Z(n15995) );
  AND U17118 ( .A(n18835), .B(n18837), .Z(n18836) );
  XNOR U17119 ( .A(n18838), .B(n18839), .Z(n15998) );
  AND U17120 ( .A(n18838), .B(n18840), .Z(n18839) );
  XNOR U17121 ( .A(n18841), .B(n18842), .Z(n16001) );
  AND U17122 ( .A(n18841), .B(n18843), .Z(n18842) );
  XNOR U17123 ( .A(n18844), .B(n18845), .Z(n16004) );
  AND U17124 ( .A(n18844), .B(n18846), .Z(n18845) );
  XNOR U17125 ( .A(n18847), .B(n18848), .Z(n16007) );
  AND U17126 ( .A(n18847), .B(n18849), .Z(n18848) );
  XNOR U17127 ( .A(n18850), .B(n18851), .Z(n16010) );
  AND U17128 ( .A(n18850), .B(n18852), .Z(n18851) );
  XNOR U17129 ( .A(n18853), .B(n18854), .Z(n16013) );
  AND U17130 ( .A(n18853), .B(n18855), .Z(n18854) );
  XNOR U17131 ( .A(n18856), .B(n18857), .Z(n16016) );
  AND U17132 ( .A(n18856), .B(n18858), .Z(n18857) );
  XNOR U17133 ( .A(n18859), .B(n18860), .Z(n16019) );
  AND U17134 ( .A(n18859), .B(n18861), .Z(n18860) );
  XNOR U17135 ( .A(n18862), .B(n18863), .Z(n16022) );
  AND U17136 ( .A(n18862), .B(n18864), .Z(n18863) );
  XNOR U17137 ( .A(n18865), .B(n18866), .Z(n16025) );
  AND U17138 ( .A(n18865), .B(n18867), .Z(n18866) );
  XNOR U17139 ( .A(n18868), .B(n18869), .Z(n16028) );
  AND U17140 ( .A(n18868), .B(n18870), .Z(n18869) );
  XNOR U17141 ( .A(n18871), .B(n18872), .Z(n16031) );
  AND U17142 ( .A(n18871), .B(n18873), .Z(n18872) );
  XNOR U17143 ( .A(n18874), .B(n18875), .Z(n16034) );
  AND U17144 ( .A(n18874), .B(n18876), .Z(n18875) );
  XNOR U17145 ( .A(n18877), .B(n18878), .Z(n16037) );
  AND U17146 ( .A(n18877), .B(n18879), .Z(n18878) );
  XNOR U17147 ( .A(n18880), .B(n18881), .Z(n16040) );
  AND U17148 ( .A(n18880), .B(n18882), .Z(n18881) );
  XNOR U17149 ( .A(n18883), .B(n18884), .Z(n16043) );
  AND U17150 ( .A(n18883), .B(n18885), .Z(n18884) );
  XNOR U17151 ( .A(n18886), .B(n18887), .Z(n16046) );
  AND U17152 ( .A(n18886), .B(n18888), .Z(n18887) );
  XNOR U17153 ( .A(n18889), .B(n18890), .Z(n16049) );
  AND U17154 ( .A(n18889), .B(n18891), .Z(n18890) );
  XNOR U17155 ( .A(n18892), .B(n18893), .Z(n16052) );
  AND U17156 ( .A(n18892), .B(n18894), .Z(n18893) );
  XNOR U17157 ( .A(n18895), .B(n18896), .Z(n16055) );
  AND U17158 ( .A(n18895), .B(n18897), .Z(n18896) );
  XNOR U17159 ( .A(n18898), .B(n18899), .Z(n16058) );
  AND U17160 ( .A(n18898), .B(n18900), .Z(n18899) );
  XNOR U17161 ( .A(n18901), .B(n18902), .Z(n16061) );
  AND U17162 ( .A(n18901), .B(n18903), .Z(n18902) );
  XNOR U17163 ( .A(n18904), .B(n18905), .Z(n16064) );
  AND U17164 ( .A(n18904), .B(n18906), .Z(n18905) );
  XNOR U17165 ( .A(n18907), .B(n18908), .Z(n16067) );
  AND U17166 ( .A(n18907), .B(n18909), .Z(n18908) );
  XNOR U17167 ( .A(n18910), .B(n18911), .Z(n16070) );
  AND U17168 ( .A(n18910), .B(n18912), .Z(n18911) );
  XNOR U17169 ( .A(n18913), .B(n18914), .Z(n16073) );
  AND U17170 ( .A(n18913), .B(n18915), .Z(n18914) );
  XNOR U17171 ( .A(n18916), .B(n18917), .Z(n16076) );
  AND U17172 ( .A(n18916), .B(n18918), .Z(n18917) );
  XNOR U17173 ( .A(n18919), .B(n18920), .Z(n16079) );
  AND U17174 ( .A(n18919), .B(n18921), .Z(n18920) );
  XNOR U17175 ( .A(n18922), .B(n18923), .Z(n16082) );
  AND U17176 ( .A(n18922), .B(n18924), .Z(n18923) );
  XNOR U17177 ( .A(n18925), .B(n18926), .Z(n16085) );
  AND U17178 ( .A(n18925), .B(n18927), .Z(n18926) );
  XNOR U17179 ( .A(n18928), .B(n18929), .Z(n16088) );
  AND U17180 ( .A(n18928), .B(n18930), .Z(n18929) );
  XNOR U17181 ( .A(n18931), .B(n18932), .Z(n16091) );
  AND U17182 ( .A(n18931), .B(n18933), .Z(n18932) );
  XNOR U17183 ( .A(n18934), .B(n18935), .Z(n16094) );
  AND U17184 ( .A(n18934), .B(n18936), .Z(n18935) );
  XNOR U17185 ( .A(n18937), .B(n18938), .Z(n16097) );
  AND U17186 ( .A(n18937), .B(n18939), .Z(n18938) );
  XNOR U17187 ( .A(n18940), .B(n18941), .Z(n16100) );
  AND U17188 ( .A(n18940), .B(n18942), .Z(n18941) );
  XNOR U17189 ( .A(n18943), .B(n18944), .Z(n16103) );
  AND U17190 ( .A(n18943), .B(n18945), .Z(n18944) );
  XNOR U17191 ( .A(n18946), .B(n18947), .Z(n16106) );
  AND U17192 ( .A(n18946), .B(n18948), .Z(n18947) );
  XNOR U17193 ( .A(n18949), .B(n18950), .Z(n16109) );
  AND U17194 ( .A(n18949), .B(n18951), .Z(n18950) );
  XNOR U17195 ( .A(n18952), .B(n18953), .Z(n16112) );
  AND U17196 ( .A(n18952), .B(n18954), .Z(n18953) );
  XNOR U17197 ( .A(n18955), .B(n18956), .Z(n16115) );
  AND U17198 ( .A(n18955), .B(n18957), .Z(n18956) );
  XNOR U17199 ( .A(n18958), .B(n18959), .Z(n16118) );
  AND U17200 ( .A(n18958), .B(n18960), .Z(n18959) );
  XNOR U17201 ( .A(n18961), .B(n18962), .Z(n16121) );
  AND U17202 ( .A(n18961), .B(n18963), .Z(n18962) );
  XNOR U17203 ( .A(n18964), .B(n18965), .Z(n16124) );
  AND U17204 ( .A(n18964), .B(n18966), .Z(n18965) );
  XNOR U17205 ( .A(n18967), .B(n18968), .Z(n16127) );
  AND U17206 ( .A(n18967), .B(n18969), .Z(n18968) );
  XNOR U17207 ( .A(n18970), .B(n18971), .Z(n16130) );
  AND U17208 ( .A(n18970), .B(n18972), .Z(n18971) );
  XNOR U17209 ( .A(n18973), .B(n18974), .Z(n16133) );
  AND U17210 ( .A(n18973), .B(n18975), .Z(n18974) );
  XNOR U17211 ( .A(n18976), .B(n18977), .Z(n16136) );
  AND U17212 ( .A(n18976), .B(n18978), .Z(n18977) );
  XNOR U17213 ( .A(n18979), .B(n18980), .Z(n16139) );
  AND U17214 ( .A(n18979), .B(n18981), .Z(n18980) );
  XNOR U17215 ( .A(n18982), .B(n18983), .Z(n16142) );
  AND U17216 ( .A(n18982), .B(n18984), .Z(n18983) );
  XNOR U17217 ( .A(n18985), .B(n18986), .Z(n16145) );
  AND U17218 ( .A(n18985), .B(n18987), .Z(n18986) );
  XNOR U17219 ( .A(n18988), .B(n18989), .Z(n16148) );
  AND U17220 ( .A(n18988), .B(n18990), .Z(n18989) );
  XNOR U17221 ( .A(n18991), .B(n18992), .Z(n16151) );
  AND U17222 ( .A(n18991), .B(n18993), .Z(n18992) );
  XNOR U17223 ( .A(n18994), .B(n18995), .Z(n16154) );
  AND U17224 ( .A(n18994), .B(n18996), .Z(n18995) );
  XNOR U17225 ( .A(n18997), .B(n18998), .Z(n16157) );
  AND U17226 ( .A(n18997), .B(n18999), .Z(n18998) );
  XNOR U17227 ( .A(n19000), .B(n19001), .Z(n16160) );
  AND U17228 ( .A(n19000), .B(n19002), .Z(n19001) );
  XNOR U17229 ( .A(n19003), .B(n19004), .Z(n16163) );
  AND U17230 ( .A(n19003), .B(n19005), .Z(n19004) );
  XNOR U17231 ( .A(n19006), .B(n19007), .Z(n16166) );
  AND U17232 ( .A(n19006), .B(n19008), .Z(n19007) );
  XNOR U17233 ( .A(n19009), .B(n19010), .Z(n16169) );
  AND U17234 ( .A(n19009), .B(n19011), .Z(n19010) );
  XNOR U17235 ( .A(n19012), .B(n19013), .Z(n16172) );
  AND U17236 ( .A(n19012), .B(n19014), .Z(n19013) );
  XNOR U17237 ( .A(n19015), .B(n19016), .Z(n16175) );
  AND U17238 ( .A(n19015), .B(n19017), .Z(n19016) );
  XNOR U17239 ( .A(n19018), .B(n19019), .Z(n16178) );
  AND U17240 ( .A(n19018), .B(n19020), .Z(n19019) );
  XNOR U17241 ( .A(n19021), .B(n19022), .Z(n16181) );
  AND U17242 ( .A(n19021), .B(n19023), .Z(n19022) );
  XNOR U17243 ( .A(n19024), .B(n19025), .Z(n16184) );
  AND U17244 ( .A(n19024), .B(n19026), .Z(n19025) );
  XNOR U17245 ( .A(n19027), .B(n19028), .Z(n16187) );
  AND U17246 ( .A(n19027), .B(n19029), .Z(n19028) );
  XNOR U17247 ( .A(n19030), .B(n19031), .Z(n16190) );
  AND U17248 ( .A(n19030), .B(n19032), .Z(n19031) );
  XNOR U17249 ( .A(n19033), .B(n19034), .Z(n16193) );
  AND U17250 ( .A(n19033), .B(n19035), .Z(n19034) );
  XNOR U17251 ( .A(n19036), .B(n19037), .Z(n16196) );
  AND U17252 ( .A(n19036), .B(n19038), .Z(n19037) );
  XNOR U17253 ( .A(n19039), .B(n19040), .Z(n16199) );
  AND U17254 ( .A(n19039), .B(n19041), .Z(n19040) );
  XNOR U17255 ( .A(n19042), .B(n19043), .Z(n16202) );
  AND U17256 ( .A(n19042), .B(n19044), .Z(n19043) );
  XNOR U17257 ( .A(n19045), .B(n19046), .Z(n16205) );
  AND U17258 ( .A(n19045), .B(n19047), .Z(n19046) );
  XNOR U17259 ( .A(n19048), .B(n19049), .Z(n16208) );
  AND U17260 ( .A(n19048), .B(n19050), .Z(n19049) );
  XNOR U17261 ( .A(n19051), .B(n19052), .Z(n16211) );
  AND U17262 ( .A(n19051), .B(n19053), .Z(n19052) );
  XNOR U17263 ( .A(n19054), .B(n19055), .Z(n16214) );
  AND U17264 ( .A(n19054), .B(n19056), .Z(n19055) );
  XNOR U17265 ( .A(n19057), .B(n19058), .Z(n16217) );
  AND U17266 ( .A(n19057), .B(n19059), .Z(n19058) );
  XNOR U17267 ( .A(n19060), .B(n19061), .Z(n16220) );
  AND U17268 ( .A(n19060), .B(n19062), .Z(n19061) );
  XNOR U17269 ( .A(n19063), .B(n19064), .Z(n16223) );
  AND U17270 ( .A(n19063), .B(n19065), .Z(n19064) );
  XNOR U17271 ( .A(n19066), .B(n19067), .Z(n16226) );
  AND U17272 ( .A(n19066), .B(n19068), .Z(n19067) );
  XNOR U17273 ( .A(n19069), .B(n19070), .Z(n16229) );
  AND U17274 ( .A(n19069), .B(n19071), .Z(n19070) );
  XNOR U17275 ( .A(n19072), .B(n19073), .Z(n16232) );
  AND U17276 ( .A(n19072), .B(n19074), .Z(n19073) );
  XNOR U17277 ( .A(n19075), .B(n19076), .Z(n16235) );
  AND U17278 ( .A(n19075), .B(n19077), .Z(n19076) );
  XNOR U17279 ( .A(n19078), .B(n19079), .Z(n16238) );
  AND U17280 ( .A(n19078), .B(n19080), .Z(n19079) );
  XNOR U17281 ( .A(n19081), .B(n19082), .Z(n16241) );
  AND U17282 ( .A(n19081), .B(n19083), .Z(n19082) );
  XNOR U17283 ( .A(n19084), .B(n19085), .Z(n16244) );
  AND U17284 ( .A(n19084), .B(n19086), .Z(n19085) );
  XNOR U17285 ( .A(n19087), .B(n19088), .Z(n16247) );
  AND U17286 ( .A(n19087), .B(n19089), .Z(n19088) );
  XNOR U17287 ( .A(n19090), .B(n19091), .Z(n16250) );
  AND U17288 ( .A(n19090), .B(n19092), .Z(n19091) );
  XNOR U17289 ( .A(n19093), .B(n19094), .Z(n16253) );
  AND U17290 ( .A(n19093), .B(n19095), .Z(n19094) );
  XNOR U17291 ( .A(n19096), .B(n19097), .Z(n16256) );
  AND U17292 ( .A(n19096), .B(n19098), .Z(n19097) );
  XNOR U17293 ( .A(n19099), .B(n19100), .Z(n16259) );
  AND U17294 ( .A(n19099), .B(n19101), .Z(n19100) );
  XNOR U17295 ( .A(n19102), .B(n19103), .Z(n16262) );
  AND U17296 ( .A(n19102), .B(n19104), .Z(n19103) );
  XNOR U17297 ( .A(n19105), .B(n19106), .Z(n16265) );
  AND U17298 ( .A(n19105), .B(n19107), .Z(n19106) );
  XNOR U17299 ( .A(n19108), .B(n19109), .Z(n16268) );
  AND U17300 ( .A(n19108), .B(n19110), .Z(n19109) );
  XNOR U17301 ( .A(n19111), .B(n19112), .Z(n16271) );
  AND U17302 ( .A(n19111), .B(n19113), .Z(n19112) );
  XNOR U17303 ( .A(n19114), .B(n19115), .Z(n16274) );
  AND U17304 ( .A(n19114), .B(n19116), .Z(n19115) );
  XNOR U17305 ( .A(n19117), .B(n19118), .Z(n16277) );
  AND U17306 ( .A(n19117), .B(n19119), .Z(n19118) );
  XNOR U17307 ( .A(n19120), .B(n19121), .Z(n16280) );
  AND U17308 ( .A(n19120), .B(n19122), .Z(n19121) );
  XNOR U17309 ( .A(n19123), .B(n19124), .Z(n16283) );
  AND U17310 ( .A(n19123), .B(n19125), .Z(n19124) );
  XNOR U17311 ( .A(n19126), .B(n19127), .Z(n16286) );
  AND U17312 ( .A(n19126), .B(n19128), .Z(n19127) );
  XNOR U17313 ( .A(n19129), .B(n19130), .Z(n16289) );
  AND U17314 ( .A(n19129), .B(n19131), .Z(n19130) );
  XNOR U17315 ( .A(n19132), .B(n19133), .Z(n16292) );
  AND U17316 ( .A(n19132), .B(n19134), .Z(n19133) );
  XNOR U17317 ( .A(n19135), .B(n19136), .Z(n16295) );
  AND U17318 ( .A(n19135), .B(n19137), .Z(n19136) );
  XNOR U17319 ( .A(n19138), .B(n19139), .Z(n16298) );
  AND U17320 ( .A(n19138), .B(n19140), .Z(n19139) );
  XNOR U17321 ( .A(n19141), .B(n19142), .Z(n16301) );
  AND U17322 ( .A(n19141), .B(n19143), .Z(n19142) );
  XNOR U17323 ( .A(n19144), .B(n19145), .Z(n16304) );
  AND U17324 ( .A(n19144), .B(n19146), .Z(n19145) );
  XNOR U17325 ( .A(n19147), .B(n19148), .Z(n16307) );
  AND U17326 ( .A(n19147), .B(n19149), .Z(n19148) );
  XNOR U17327 ( .A(n19150), .B(n19151), .Z(n16310) );
  AND U17328 ( .A(n19150), .B(n19152), .Z(n19151) );
  XNOR U17329 ( .A(n19153), .B(n19154), .Z(n16313) );
  AND U17330 ( .A(n19153), .B(n19155), .Z(n19154) );
  XNOR U17331 ( .A(n19156), .B(n19157), .Z(n16316) );
  AND U17332 ( .A(n19156), .B(n19158), .Z(n19157) );
  XNOR U17333 ( .A(n19159), .B(n19160), .Z(n16319) );
  AND U17334 ( .A(n19159), .B(n19161), .Z(n19160) );
  XNOR U17335 ( .A(n19162), .B(n19163), .Z(n16322) );
  AND U17336 ( .A(n19162), .B(n19164), .Z(n19163) );
  XNOR U17337 ( .A(n19165), .B(n19166), .Z(n16325) );
  AND U17338 ( .A(n19165), .B(n19167), .Z(n19166) );
  XNOR U17339 ( .A(n19168), .B(n19169), .Z(n16328) );
  AND U17340 ( .A(n19168), .B(n19170), .Z(n19169) );
  XNOR U17341 ( .A(n19171), .B(n19172), .Z(n16331) );
  AND U17342 ( .A(n19171), .B(n19173), .Z(n19172) );
  XNOR U17343 ( .A(n19174), .B(n19175), .Z(n16334) );
  AND U17344 ( .A(n19174), .B(n19176), .Z(n19175) );
  XNOR U17345 ( .A(n19177), .B(n19178), .Z(n16337) );
  AND U17346 ( .A(n19177), .B(n19179), .Z(n19178) );
  XNOR U17347 ( .A(n19180), .B(n19181), .Z(n16340) );
  AND U17348 ( .A(n19180), .B(n19182), .Z(n19181) );
  XNOR U17349 ( .A(n19183), .B(n19184), .Z(n16343) );
  AND U17350 ( .A(n19183), .B(n19185), .Z(n19184) );
  XNOR U17351 ( .A(n19186), .B(n19187), .Z(n16346) );
  AND U17352 ( .A(n19186), .B(n19188), .Z(n19187) );
  XNOR U17353 ( .A(n19189), .B(n19190), .Z(n16349) );
  AND U17354 ( .A(n19189), .B(n19191), .Z(n19190) );
  XNOR U17355 ( .A(n19192), .B(n19193), .Z(n16352) );
  AND U17356 ( .A(n19192), .B(n19194), .Z(n19193) );
  XNOR U17357 ( .A(n19195), .B(n19196), .Z(n16355) );
  AND U17358 ( .A(n19195), .B(n19197), .Z(n19196) );
  XNOR U17359 ( .A(n19198), .B(n19199), .Z(n16358) );
  AND U17360 ( .A(n19198), .B(n19200), .Z(n19199) );
  XNOR U17361 ( .A(n19201), .B(n19202), .Z(n16361) );
  AND U17362 ( .A(n19201), .B(n19203), .Z(n19202) );
  XNOR U17363 ( .A(n19204), .B(n19205), .Z(n16364) );
  AND U17364 ( .A(n19204), .B(n19206), .Z(n19205) );
  XNOR U17365 ( .A(n19207), .B(n19208), .Z(n16367) );
  AND U17366 ( .A(n19207), .B(n19209), .Z(n19208) );
  XNOR U17367 ( .A(n19210), .B(n19211), .Z(n16370) );
  AND U17368 ( .A(n19210), .B(n19212), .Z(n19211) );
  XNOR U17369 ( .A(n19213), .B(n19214), .Z(n16373) );
  AND U17370 ( .A(n19213), .B(n19215), .Z(n19214) );
  XNOR U17371 ( .A(n19216), .B(n19217), .Z(n16376) );
  AND U17372 ( .A(n19216), .B(n19218), .Z(n19217) );
  XNOR U17373 ( .A(n19219), .B(n19220), .Z(n16379) );
  AND U17374 ( .A(n19219), .B(n19221), .Z(n19220) );
  XNOR U17375 ( .A(n19222), .B(n19223), .Z(n16382) );
  AND U17376 ( .A(n19222), .B(n19224), .Z(n19223) );
  XNOR U17377 ( .A(n19225), .B(n19226), .Z(n16385) );
  AND U17378 ( .A(n19225), .B(n19227), .Z(n19226) );
  XNOR U17379 ( .A(n19228), .B(n19229), .Z(n16388) );
  AND U17380 ( .A(n19228), .B(n19230), .Z(n19229) );
  XNOR U17381 ( .A(n19231), .B(n19232), .Z(n16391) );
  AND U17382 ( .A(n19231), .B(n19233), .Z(n19232) );
  XNOR U17383 ( .A(n19234), .B(n19235), .Z(n16394) );
  AND U17384 ( .A(n19234), .B(n19236), .Z(n19235) );
  XNOR U17385 ( .A(n19237), .B(n19238), .Z(n16397) );
  AND U17386 ( .A(n19237), .B(n19239), .Z(n19238) );
  XNOR U17387 ( .A(n19240), .B(n19241), .Z(n16400) );
  AND U17388 ( .A(n19240), .B(n19242), .Z(n19241) );
  XNOR U17389 ( .A(n19243), .B(n19244), .Z(n16403) );
  AND U17390 ( .A(n19243), .B(n19245), .Z(n19244) );
  XNOR U17391 ( .A(n19246), .B(n19247), .Z(n16406) );
  AND U17392 ( .A(n19246), .B(n19248), .Z(n19247) );
  XNOR U17393 ( .A(n19249), .B(n19250), .Z(n16409) );
  AND U17394 ( .A(n19249), .B(n19251), .Z(n19250) );
  XNOR U17395 ( .A(n19252), .B(n19253), .Z(n16412) );
  AND U17396 ( .A(n19252), .B(n19254), .Z(n19253) );
  XNOR U17397 ( .A(n19255), .B(n19256), .Z(n16415) );
  AND U17398 ( .A(n19255), .B(n19257), .Z(n19256) );
  XNOR U17399 ( .A(n19258), .B(n19259), .Z(n16418) );
  AND U17400 ( .A(n19258), .B(n19260), .Z(n19259) );
  XNOR U17401 ( .A(n19261), .B(n19262), .Z(n16421) );
  AND U17402 ( .A(n19261), .B(n19263), .Z(n19262) );
  XNOR U17403 ( .A(n19264), .B(n19265), .Z(n16424) );
  AND U17404 ( .A(n19264), .B(n19266), .Z(n19265) );
  XNOR U17405 ( .A(n19267), .B(n19268), .Z(n16427) );
  AND U17406 ( .A(n19267), .B(n19269), .Z(n19268) );
  XNOR U17407 ( .A(n19270), .B(n19271), .Z(n16430) );
  AND U17408 ( .A(n19270), .B(n19272), .Z(n19271) );
  XNOR U17409 ( .A(n19273), .B(n19274), .Z(n16433) );
  AND U17410 ( .A(n19273), .B(n19275), .Z(n19274) );
  XNOR U17411 ( .A(n19276), .B(n19277), .Z(n16436) );
  AND U17412 ( .A(n19276), .B(n19278), .Z(n19277) );
  XNOR U17413 ( .A(n19279), .B(n19280), .Z(n16439) );
  AND U17414 ( .A(n19279), .B(n19281), .Z(n19280) );
  XNOR U17415 ( .A(n19282), .B(n19283), .Z(n16442) );
  AND U17416 ( .A(n19282), .B(n19284), .Z(n19283) );
  XNOR U17417 ( .A(n19285), .B(n19286), .Z(n16445) );
  AND U17418 ( .A(n19285), .B(n19287), .Z(n19286) );
  XNOR U17419 ( .A(n19288), .B(n19289), .Z(n16448) );
  AND U17420 ( .A(n19288), .B(n19290), .Z(n19289) );
  XNOR U17421 ( .A(n19291), .B(n19292), .Z(n16451) );
  AND U17422 ( .A(n19291), .B(n19293), .Z(n19292) );
  XNOR U17423 ( .A(n19294), .B(n19295), .Z(n16454) );
  AND U17424 ( .A(n19294), .B(n19296), .Z(n19295) );
  XNOR U17425 ( .A(n19297), .B(n19298), .Z(n16457) );
  AND U17426 ( .A(n19297), .B(n19299), .Z(n19298) );
  XNOR U17427 ( .A(n19300), .B(n19301), .Z(n16460) );
  AND U17428 ( .A(n19300), .B(n19302), .Z(n19301) );
  XNOR U17429 ( .A(n19303), .B(n19304), .Z(n16463) );
  AND U17430 ( .A(n19303), .B(n19305), .Z(n19304) );
  XNOR U17431 ( .A(n19306), .B(n19307), .Z(n16466) );
  AND U17432 ( .A(n19306), .B(n19308), .Z(n19307) );
  XNOR U17433 ( .A(n19309), .B(n19310), .Z(n16469) );
  AND U17434 ( .A(n19309), .B(n19311), .Z(n19310) );
  XNOR U17435 ( .A(n19312), .B(n19313), .Z(n16472) );
  AND U17436 ( .A(n19312), .B(n19314), .Z(n19313) );
  XNOR U17437 ( .A(n19315), .B(n19316), .Z(n16475) );
  AND U17438 ( .A(n19315), .B(n19317), .Z(n19316) );
  XNOR U17439 ( .A(n19318), .B(n19319), .Z(n16478) );
  AND U17440 ( .A(n19318), .B(n19320), .Z(n19319) );
  XNOR U17441 ( .A(n19321), .B(n19322), .Z(n16481) );
  AND U17442 ( .A(n19321), .B(n19323), .Z(n19322) );
  XNOR U17443 ( .A(n19324), .B(n19325), .Z(n16484) );
  AND U17444 ( .A(n19324), .B(n19326), .Z(n19325) );
  XNOR U17445 ( .A(n19327), .B(n19328), .Z(n16487) );
  AND U17446 ( .A(n19327), .B(n19329), .Z(n19328) );
  XNOR U17447 ( .A(n19330), .B(n19331), .Z(n16490) );
  AND U17448 ( .A(n19330), .B(n19332), .Z(n19331) );
  XNOR U17449 ( .A(n19333), .B(n19334), .Z(n16493) );
  AND U17450 ( .A(n19333), .B(n19335), .Z(n19334) );
  XNOR U17451 ( .A(n19336), .B(n19337), .Z(n16496) );
  AND U17452 ( .A(n19336), .B(n19338), .Z(n19337) );
  XNOR U17453 ( .A(n19339), .B(n19340), .Z(n16499) );
  AND U17454 ( .A(n19339), .B(n19341), .Z(n19340) );
  XNOR U17455 ( .A(n19342), .B(n19343), .Z(n16502) );
  AND U17456 ( .A(n19342), .B(n19344), .Z(n19343) );
  XNOR U17457 ( .A(n19345), .B(n19346), .Z(n16505) );
  AND U17458 ( .A(n19345), .B(n19347), .Z(n19346) );
  XNOR U17459 ( .A(n19348), .B(n19349), .Z(n16508) );
  AND U17460 ( .A(n19348), .B(n19350), .Z(n19349) );
  XNOR U17461 ( .A(n19351), .B(n19352), .Z(n16511) );
  AND U17462 ( .A(n19351), .B(n19353), .Z(n19352) );
  XNOR U17463 ( .A(n19354), .B(n19355), .Z(n16514) );
  AND U17464 ( .A(n19354), .B(n19356), .Z(n19355) );
  XNOR U17465 ( .A(n19357), .B(n19358), .Z(n16517) );
  AND U17466 ( .A(n19357), .B(n19359), .Z(n19358) );
  XNOR U17467 ( .A(n19360), .B(n19361), .Z(n16520) );
  AND U17468 ( .A(n19360), .B(n19362), .Z(n19361) );
  XNOR U17469 ( .A(n19363), .B(n19364), .Z(n16523) );
  AND U17470 ( .A(n19363), .B(n19365), .Z(n19364) );
  XNOR U17471 ( .A(n19366), .B(n19367), .Z(n16526) );
  AND U17472 ( .A(n19366), .B(n19368), .Z(n19367) );
  XNOR U17473 ( .A(n19369), .B(n19370), .Z(n16529) );
  AND U17474 ( .A(n19369), .B(n19371), .Z(n19370) );
  XNOR U17475 ( .A(n19372), .B(n19373), .Z(n16532) );
  AND U17476 ( .A(n19372), .B(n19374), .Z(n19373) );
  XNOR U17477 ( .A(n19375), .B(n19376), .Z(n16535) );
  AND U17478 ( .A(n19375), .B(n19377), .Z(n19376) );
  XNOR U17479 ( .A(n19378), .B(n19379), .Z(n16538) );
  AND U17480 ( .A(n19378), .B(n19380), .Z(n19379) );
  XNOR U17481 ( .A(n19381), .B(n19382), .Z(n16541) );
  AND U17482 ( .A(n19381), .B(n19383), .Z(n19382) );
  XNOR U17483 ( .A(n19384), .B(n19385), .Z(n16544) );
  AND U17484 ( .A(n19384), .B(n19386), .Z(n19385) );
  XNOR U17485 ( .A(n19387), .B(n19388), .Z(n16547) );
  AND U17486 ( .A(n19387), .B(n19389), .Z(n19388) );
  XNOR U17487 ( .A(n19390), .B(n19391), .Z(n16550) );
  AND U17488 ( .A(n19390), .B(n19392), .Z(n19391) );
  XNOR U17489 ( .A(n19393), .B(n19394), .Z(n16553) );
  AND U17490 ( .A(n19393), .B(n19395), .Z(n19394) );
  XNOR U17491 ( .A(n19396), .B(n19397), .Z(n16556) );
  AND U17492 ( .A(n19396), .B(n19398), .Z(n19397) );
  XNOR U17493 ( .A(n19399), .B(n19400), .Z(n16559) );
  AND U17494 ( .A(n19399), .B(n19401), .Z(n19400) );
  XNOR U17495 ( .A(n19402), .B(n19403), .Z(n16562) );
  AND U17496 ( .A(n19402), .B(n19404), .Z(n19403) );
  XNOR U17497 ( .A(n19405), .B(n19406), .Z(n16565) );
  AND U17498 ( .A(n19405), .B(n19407), .Z(n19406) );
  XNOR U17499 ( .A(n19408), .B(n19409), .Z(n16568) );
  AND U17500 ( .A(n19408), .B(n19410), .Z(n19409) );
  XNOR U17501 ( .A(n19411), .B(n19412), .Z(n16571) );
  AND U17502 ( .A(n19411), .B(n19413), .Z(n19412) );
  XNOR U17503 ( .A(n19414), .B(n19415), .Z(n16574) );
  AND U17504 ( .A(n19414), .B(n19416), .Z(n19415) );
  XNOR U17505 ( .A(n19417), .B(n19418), .Z(n16577) );
  AND U17506 ( .A(n19417), .B(n19419), .Z(n19418) );
  XNOR U17507 ( .A(n19420), .B(n19421), .Z(n16580) );
  AND U17508 ( .A(n19420), .B(n19422), .Z(n19421) );
  XNOR U17509 ( .A(n19423), .B(n19424), .Z(n16583) );
  AND U17510 ( .A(n19423), .B(n19425), .Z(n19424) );
  XNOR U17511 ( .A(n19426), .B(n19427), .Z(n16586) );
  AND U17512 ( .A(n19426), .B(n19428), .Z(n19427) );
  XNOR U17513 ( .A(n19429), .B(n19430), .Z(n16589) );
  AND U17514 ( .A(n19429), .B(n19431), .Z(n19430) );
  XNOR U17515 ( .A(n19432), .B(n19433), .Z(n16592) );
  AND U17516 ( .A(n19432), .B(n19434), .Z(n19433) );
  XNOR U17517 ( .A(n19435), .B(n19436), .Z(n16595) );
  AND U17518 ( .A(n19435), .B(n19437), .Z(n19436) );
  XNOR U17519 ( .A(n19438), .B(n19439), .Z(n16598) );
  AND U17520 ( .A(n19438), .B(n19440), .Z(n19439) );
  XNOR U17521 ( .A(n19441), .B(n19442), .Z(n16601) );
  AND U17522 ( .A(n19441), .B(n19443), .Z(n19442) );
  XNOR U17523 ( .A(n19444), .B(n19445), .Z(n16604) );
  AND U17524 ( .A(n19444), .B(n19446), .Z(n19445) );
  XNOR U17525 ( .A(n19447), .B(n19448), .Z(n16607) );
  AND U17526 ( .A(n19447), .B(n19449), .Z(n19448) );
  XNOR U17527 ( .A(n19450), .B(n19451), .Z(n16610) );
  AND U17528 ( .A(n19450), .B(n19452), .Z(n19451) );
  XNOR U17529 ( .A(n19453), .B(n19454), .Z(n16613) );
  AND U17530 ( .A(n19453), .B(n19455), .Z(n19454) );
  XNOR U17531 ( .A(n19456), .B(n19457), .Z(n16616) );
  AND U17532 ( .A(n19456), .B(n19458), .Z(n19457) );
  XNOR U17533 ( .A(n19459), .B(n19460), .Z(n16619) );
  AND U17534 ( .A(n19459), .B(n19461), .Z(n19460) );
  XNOR U17535 ( .A(n19462), .B(n19463), .Z(n16622) );
  AND U17536 ( .A(n19462), .B(n19464), .Z(n19463) );
  XNOR U17537 ( .A(n19465), .B(n19466), .Z(n16625) );
  AND U17538 ( .A(n19465), .B(n19467), .Z(n19466) );
  XNOR U17539 ( .A(n19468), .B(n19469), .Z(n16628) );
  AND U17540 ( .A(n19468), .B(n19470), .Z(n19469) );
  XNOR U17541 ( .A(n19471), .B(n19472), .Z(n16631) );
  AND U17542 ( .A(n19471), .B(n19473), .Z(n19472) );
  XNOR U17543 ( .A(n19474), .B(n19475), .Z(n16634) );
  AND U17544 ( .A(n19474), .B(n19476), .Z(n19475) );
  XNOR U17545 ( .A(n19477), .B(n19478), .Z(n16637) );
  AND U17546 ( .A(n19477), .B(n19479), .Z(n19478) );
  XNOR U17547 ( .A(n19480), .B(n19481), .Z(n16640) );
  AND U17548 ( .A(n19480), .B(n19482), .Z(n19481) );
  XNOR U17549 ( .A(n19483), .B(n19484), .Z(n16643) );
  AND U17550 ( .A(n19483), .B(n19485), .Z(n19484) );
  XNOR U17551 ( .A(n19486), .B(n19487), .Z(n16646) );
  AND U17552 ( .A(n19486), .B(n19488), .Z(n19487) );
  XNOR U17553 ( .A(n19489), .B(n19490), .Z(n16649) );
  AND U17554 ( .A(n19489), .B(n19491), .Z(n19490) );
  XNOR U17555 ( .A(n19492), .B(n19493), .Z(n16652) );
  AND U17556 ( .A(n19492), .B(n19494), .Z(n19493) );
  XNOR U17557 ( .A(n19495), .B(n19496), .Z(n16655) );
  AND U17558 ( .A(n19495), .B(n19497), .Z(n19496) );
  XNOR U17559 ( .A(n19498), .B(n19499), .Z(n16658) );
  AND U17560 ( .A(n19498), .B(n19500), .Z(n19499) );
  XNOR U17561 ( .A(n19501), .B(n19502), .Z(n16661) );
  AND U17562 ( .A(n19501), .B(n19503), .Z(n19502) );
  XNOR U17563 ( .A(n19504), .B(n19505), .Z(n16664) );
  AND U17564 ( .A(n19504), .B(n19506), .Z(n19505) );
  XNOR U17565 ( .A(n19507), .B(n19508), .Z(n16667) );
  AND U17566 ( .A(n19507), .B(n19509), .Z(n19508) );
  XNOR U17567 ( .A(n19510), .B(n19511), .Z(n16670) );
  AND U17568 ( .A(n19510), .B(n19512), .Z(n19511) );
  XNOR U17569 ( .A(n19513), .B(n19514), .Z(n16673) );
  AND U17570 ( .A(n19513), .B(n19515), .Z(n19514) );
  XNOR U17571 ( .A(n19516), .B(n19517), .Z(n16676) );
  AND U17572 ( .A(n19516), .B(n19518), .Z(n19517) );
  XNOR U17573 ( .A(n19519), .B(n19520), .Z(n16679) );
  AND U17574 ( .A(n19519), .B(n19521), .Z(n19520) );
  XNOR U17575 ( .A(n19522), .B(n19523), .Z(n16682) );
  AND U17576 ( .A(n19522), .B(n19524), .Z(n19523) );
  XNOR U17577 ( .A(n19525), .B(n19526), .Z(n16685) );
  AND U17578 ( .A(n19525), .B(n19527), .Z(n19526) );
  XNOR U17579 ( .A(n19528), .B(n19529), .Z(n16688) );
  AND U17580 ( .A(n19528), .B(n19530), .Z(n19529) );
  XNOR U17581 ( .A(n19531), .B(n19532), .Z(n16691) );
  AND U17582 ( .A(n19531), .B(n19533), .Z(n19532) );
  XNOR U17583 ( .A(n19534), .B(n19535), .Z(n16694) );
  AND U17584 ( .A(n19534), .B(n19536), .Z(n19535) );
  XNOR U17585 ( .A(n19537), .B(n19538), .Z(n16697) );
  AND U17586 ( .A(n19537), .B(n19539), .Z(n19538) );
  XNOR U17587 ( .A(n19540), .B(n19541), .Z(n16700) );
  AND U17588 ( .A(n19540), .B(n19542), .Z(n19541) );
  XNOR U17589 ( .A(n19543), .B(n19544), .Z(n16703) );
  AND U17590 ( .A(n19543), .B(n19545), .Z(n19544) );
  XNOR U17591 ( .A(n19546), .B(n19547), .Z(n16706) );
  AND U17592 ( .A(n19546), .B(n19548), .Z(n19547) );
  XNOR U17593 ( .A(n19549), .B(n19550), .Z(n16709) );
  AND U17594 ( .A(n19549), .B(n19551), .Z(n19550) );
  XNOR U17595 ( .A(n19552), .B(n19553), .Z(n16712) );
  AND U17596 ( .A(n19552), .B(n19554), .Z(n19553) );
  XNOR U17597 ( .A(n19555), .B(n19556), .Z(n16715) );
  AND U17598 ( .A(n19555), .B(n19557), .Z(n19556) );
  XNOR U17599 ( .A(n19558), .B(n19559), .Z(n16718) );
  AND U17600 ( .A(n19558), .B(n19560), .Z(n19559) );
  XNOR U17601 ( .A(n19561), .B(n19562), .Z(n16721) );
  AND U17602 ( .A(n19561), .B(n19563), .Z(n19562) );
  XNOR U17603 ( .A(n19564), .B(n19565), .Z(n16724) );
  AND U17604 ( .A(n19564), .B(n19566), .Z(n19565) );
  XNOR U17605 ( .A(n19567), .B(n19568), .Z(n16727) );
  AND U17606 ( .A(n19567), .B(n19569), .Z(n19568) );
  XNOR U17607 ( .A(n19570), .B(n19571), .Z(n16730) );
  AND U17608 ( .A(n19570), .B(n19572), .Z(n19571) );
  XNOR U17609 ( .A(n19573), .B(n19574), .Z(n16733) );
  AND U17610 ( .A(n19573), .B(n19575), .Z(n19574) );
  XNOR U17611 ( .A(n19576), .B(n19577), .Z(n16736) );
  AND U17612 ( .A(n19576), .B(n19578), .Z(n19577) );
  XNOR U17613 ( .A(n19579), .B(n19580), .Z(n16739) );
  AND U17614 ( .A(n19579), .B(n19581), .Z(n19580) );
  XNOR U17615 ( .A(n19582), .B(n19583), .Z(n16742) );
  AND U17616 ( .A(n19582), .B(n19584), .Z(n19583) );
  XNOR U17617 ( .A(n19585), .B(n19586), .Z(n16745) );
  AND U17618 ( .A(n19585), .B(n19587), .Z(n19586) );
  XNOR U17619 ( .A(n19588), .B(n19589), .Z(n16748) );
  AND U17620 ( .A(n19588), .B(n19590), .Z(n19589) );
  XNOR U17621 ( .A(n19591), .B(n19592), .Z(n16751) );
  AND U17622 ( .A(n19591), .B(n19593), .Z(n19592) );
  XNOR U17623 ( .A(n19594), .B(n19595), .Z(n16754) );
  AND U17624 ( .A(n19594), .B(n19596), .Z(n19595) );
  XNOR U17625 ( .A(n19597), .B(n19598), .Z(n16757) );
  AND U17626 ( .A(n19597), .B(n19599), .Z(n19598) );
  XNOR U17627 ( .A(n19600), .B(n19601), .Z(n16760) );
  AND U17628 ( .A(n19600), .B(n19602), .Z(n19601) );
  XNOR U17629 ( .A(n19603), .B(n19604), .Z(n16763) );
  AND U17630 ( .A(n19603), .B(n19605), .Z(n19604) );
  XNOR U17631 ( .A(n19606), .B(n19607), .Z(n16766) );
  AND U17632 ( .A(n19606), .B(n19608), .Z(n19607) );
  XNOR U17633 ( .A(n19609), .B(n19610), .Z(n16769) );
  AND U17634 ( .A(n19609), .B(n19611), .Z(n19610) );
  XNOR U17635 ( .A(n19612), .B(n19613), .Z(n16772) );
  AND U17636 ( .A(n19612), .B(n19614), .Z(n19613) );
  XNOR U17637 ( .A(n19615), .B(n19616), .Z(n16775) );
  AND U17638 ( .A(n19615), .B(n19617), .Z(n19616) );
  XNOR U17639 ( .A(n19618), .B(n19619), .Z(n16778) );
  AND U17640 ( .A(n19618), .B(n19620), .Z(n19619) );
  XNOR U17641 ( .A(n19621), .B(n19622), .Z(n16781) );
  AND U17642 ( .A(n19621), .B(n19623), .Z(n19622) );
  XNOR U17643 ( .A(n19624), .B(n19625), .Z(n16784) );
  AND U17644 ( .A(n19624), .B(n19626), .Z(n19625) );
  XNOR U17645 ( .A(n19627), .B(n19628), .Z(n16787) );
  AND U17646 ( .A(n19627), .B(n19629), .Z(n19628) );
  XNOR U17647 ( .A(n19630), .B(n19631), .Z(n16790) );
  AND U17648 ( .A(n19630), .B(n19632), .Z(n19631) );
  XNOR U17649 ( .A(n19633), .B(n19634), .Z(n16793) );
  AND U17650 ( .A(n19633), .B(n19635), .Z(n19634) );
  XNOR U17651 ( .A(n19636), .B(n19637), .Z(n16796) );
  AND U17652 ( .A(n19636), .B(n19638), .Z(n19637) );
  XNOR U17653 ( .A(n19639), .B(n19640), .Z(n16799) );
  AND U17654 ( .A(n19639), .B(n19641), .Z(n19640) );
  XNOR U17655 ( .A(n19642), .B(n19643), .Z(n16802) );
  AND U17656 ( .A(n19642), .B(n19644), .Z(n19643) );
  XNOR U17657 ( .A(n19645), .B(n19646), .Z(n16805) );
  AND U17658 ( .A(n19645), .B(n19647), .Z(n19646) );
  XNOR U17659 ( .A(n19648), .B(n19649), .Z(n16808) );
  AND U17660 ( .A(n19648), .B(n19650), .Z(n19649) );
  XNOR U17661 ( .A(n19651), .B(n19652), .Z(n16811) );
  AND U17662 ( .A(n19651), .B(n19653), .Z(n19652) );
  XNOR U17663 ( .A(n19654), .B(n19655), .Z(n16814) );
  AND U17664 ( .A(n19654), .B(n19656), .Z(n19655) );
  XNOR U17665 ( .A(n19657), .B(n19658), .Z(n16817) );
  AND U17666 ( .A(n19657), .B(n19659), .Z(n19658) );
  XNOR U17667 ( .A(n19660), .B(n19661), .Z(n16820) );
  AND U17668 ( .A(n19660), .B(n19662), .Z(n19661) );
  XNOR U17669 ( .A(n19663), .B(n19664), .Z(n16823) );
  AND U17670 ( .A(n19663), .B(n19665), .Z(n19664) );
  XNOR U17671 ( .A(n19666), .B(n19667), .Z(n16826) );
  AND U17672 ( .A(n19666), .B(n19668), .Z(n19667) );
  XNOR U17673 ( .A(n19669), .B(n19670), .Z(n16829) );
  AND U17674 ( .A(n19669), .B(n19671), .Z(n19670) );
  XNOR U17675 ( .A(n19672), .B(n19673), .Z(n16832) );
  AND U17676 ( .A(n19672), .B(n19674), .Z(n19673) );
  XNOR U17677 ( .A(n19675), .B(n19676), .Z(n16835) );
  AND U17678 ( .A(n19675), .B(n19677), .Z(n19676) );
  XNOR U17679 ( .A(n19678), .B(n19679), .Z(n16838) );
  AND U17680 ( .A(n19678), .B(n19680), .Z(n19679) );
  XNOR U17681 ( .A(n19681), .B(n19682), .Z(n16841) );
  AND U17682 ( .A(n19681), .B(n19683), .Z(n19682) );
  XNOR U17683 ( .A(n19684), .B(n19685), .Z(n16844) );
  AND U17684 ( .A(n19684), .B(n19686), .Z(n19685) );
  XNOR U17685 ( .A(n19687), .B(n19688), .Z(n16847) );
  AND U17686 ( .A(n19687), .B(n19689), .Z(n19688) );
  XNOR U17687 ( .A(n19690), .B(n19691), .Z(n16850) );
  AND U17688 ( .A(n19690), .B(n19692), .Z(n19691) );
  XNOR U17689 ( .A(n19693), .B(n19694), .Z(n16853) );
  AND U17690 ( .A(n19693), .B(n19695), .Z(n19694) );
  XNOR U17691 ( .A(n19696), .B(n19697), .Z(n16856) );
  AND U17692 ( .A(n19696), .B(n19698), .Z(n19697) );
  XNOR U17693 ( .A(n19699), .B(n19700), .Z(n16859) );
  AND U17694 ( .A(n19699), .B(n19701), .Z(n19700) );
  XNOR U17695 ( .A(n19702), .B(n19703), .Z(n16862) );
  AND U17696 ( .A(n19702), .B(n19704), .Z(n19703) );
  XNOR U17697 ( .A(n19705), .B(n19706), .Z(n16865) );
  AND U17698 ( .A(n19705), .B(n19707), .Z(n19706) );
  XNOR U17699 ( .A(n19708), .B(n19709), .Z(n16868) );
  AND U17700 ( .A(n19708), .B(n19710), .Z(n19709) );
  XNOR U17701 ( .A(n19711), .B(n19712), .Z(n16871) );
  AND U17702 ( .A(n19711), .B(n19713), .Z(n19712) );
  XNOR U17703 ( .A(n19714), .B(n19715), .Z(n16874) );
  AND U17704 ( .A(n19714), .B(n19716), .Z(n19715) );
  XNOR U17705 ( .A(n19717), .B(n19718), .Z(n16877) );
  AND U17706 ( .A(n19717), .B(n19719), .Z(n19718) );
  XNOR U17707 ( .A(n19720), .B(n19721), .Z(n16880) );
  AND U17708 ( .A(n19720), .B(n19722), .Z(n19721) );
  XNOR U17709 ( .A(n19723), .B(n19724), .Z(n16883) );
  AND U17710 ( .A(n19723), .B(n19725), .Z(n19724) );
  XNOR U17711 ( .A(n19726), .B(n19727), .Z(n16886) );
  AND U17712 ( .A(n19726), .B(n19728), .Z(n19727) );
  XNOR U17713 ( .A(n19729), .B(n19730), .Z(n16889) );
  AND U17714 ( .A(n19729), .B(n19731), .Z(n19730) );
  XNOR U17715 ( .A(n19732), .B(n19733), .Z(n16892) );
  AND U17716 ( .A(n19732), .B(n19734), .Z(n19733) );
  XNOR U17717 ( .A(n19735), .B(n19736), .Z(n16895) );
  AND U17718 ( .A(n19735), .B(n19737), .Z(n19736) );
  XNOR U17719 ( .A(n19738), .B(n19739), .Z(n16898) );
  AND U17720 ( .A(n19738), .B(n19740), .Z(n19739) );
  XNOR U17721 ( .A(n19741), .B(n19742), .Z(n16901) );
  AND U17722 ( .A(n19741), .B(n19743), .Z(n19742) );
  XNOR U17723 ( .A(n19744), .B(n19745), .Z(n16904) );
  AND U17724 ( .A(n19744), .B(n19746), .Z(n19745) );
  XNOR U17725 ( .A(n19747), .B(n19748), .Z(n16907) );
  AND U17726 ( .A(n19747), .B(n19749), .Z(n19748) );
  XNOR U17727 ( .A(n19750), .B(n19751), .Z(n16910) );
  AND U17728 ( .A(n19750), .B(n19752), .Z(n19751) );
  XNOR U17729 ( .A(n19753), .B(n19754), .Z(n16913) );
  AND U17730 ( .A(n19753), .B(n19755), .Z(n19754) );
  XNOR U17731 ( .A(n19756), .B(n19757), .Z(n16916) );
  AND U17732 ( .A(n19756), .B(n19758), .Z(n19757) );
  XNOR U17733 ( .A(n19759), .B(n19760), .Z(n16919) );
  AND U17734 ( .A(n19759), .B(n19761), .Z(n19760) );
  XNOR U17735 ( .A(n19762), .B(n19763), .Z(n16922) );
  AND U17736 ( .A(n19762), .B(n19764), .Z(n19763) );
  XNOR U17737 ( .A(n19765), .B(n19766), .Z(n16925) );
  AND U17738 ( .A(n19765), .B(n19767), .Z(n19766) );
  XNOR U17739 ( .A(n19768), .B(n19769), .Z(n16928) );
  AND U17740 ( .A(n19768), .B(n19770), .Z(n19769) );
  XNOR U17741 ( .A(n19771), .B(n19772), .Z(n16931) );
  AND U17742 ( .A(n19771), .B(n19773), .Z(n19772) );
  XNOR U17743 ( .A(n19774), .B(n19775), .Z(n16934) );
  AND U17744 ( .A(n19774), .B(n19776), .Z(n19775) );
  XNOR U17745 ( .A(n19777), .B(n19778), .Z(n16937) );
  AND U17746 ( .A(n19777), .B(n19779), .Z(n19778) );
  XNOR U17747 ( .A(n19780), .B(n19781), .Z(n16940) );
  AND U17748 ( .A(n19780), .B(n19782), .Z(n19781) );
  XNOR U17749 ( .A(n19783), .B(n19784), .Z(n16943) );
  AND U17750 ( .A(n19783), .B(n19785), .Z(n19784) );
  XNOR U17751 ( .A(n19786), .B(n19787), .Z(n16946) );
  AND U17752 ( .A(n19786), .B(n19788), .Z(n19787) );
  XNOR U17753 ( .A(n19789), .B(n19790), .Z(n16949) );
  AND U17754 ( .A(n19789), .B(n19791), .Z(n19790) );
  XNOR U17755 ( .A(n19792), .B(n19793), .Z(n16952) );
  AND U17756 ( .A(n19792), .B(n19794), .Z(n19793) );
  XNOR U17757 ( .A(n19795), .B(n19796), .Z(n16955) );
  AND U17758 ( .A(n19795), .B(n19797), .Z(n19796) );
  XNOR U17759 ( .A(n19798), .B(n19799), .Z(n16958) );
  AND U17760 ( .A(n19798), .B(n19800), .Z(n19799) );
  XNOR U17761 ( .A(n19801), .B(n19802), .Z(n16961) );
  AND U17762 ( .A(n19801), .B(n19803), .Z(n19802) );
  XNOR U17763 ( .A(n19804), .B(n19805), .Z(n16964) );
  AND U17764 ( .A(n19804), .B(n19806), .Z(n19805) );
  XNOR U17765 ( .A(n19807), .B(n19808), .Z(n16967) );
  AND U17766 ( .A(n19807), .B(n19809), .Z(n19808) );
  XNOR U17767 ( .A(n19810), .B(n19811), .Z(n16970) );
  AND U17768 ( .A(n19810), .B(n19812), .Z(n19811) );
  XNOR U17769 ( .A(n19813), .B(n19814), .Z(n16973) );
  AND U17770 ( .A(n19813), .B(n19815), .Z(n19814) );
  XNOR U17771 ( .A(n19816), .B(n19817), .Z(n16976) );
  AND U17772 ( .A(n19816), .B(n19818), .Z(n19817) );
  XNOR U17773 ( .A(n19819), .B(n19820), .Z(n16979) );
  AND U17774 ( .A(n19819), .B(n19821), .Z(n19820) );
  XNOR U17775 ( .A(n19822), .B(n19823), .Z(n16982) );
  AND U17776 ( .A(n19822), .B(n19824), .Z(n19823) );
  XNOR U17777 ( .A(n19825), .B(n19826), .Z(n16985) );
  AND U17778 ( .A(n19825), .B(n19827), .Z(n19826) );
  XNOR U17779 ( .A(n19828), .B(n19829), .Z(n16988) );
  AND U17780 ( .A(n19828), .B(n19830), .Z(n19829) );
  XNOR U17781 ( .A(n19831), .B(n19832), .Z(n16991) );
  AND U17782 ( .A(n19831), .B(n19833), .Z(n19832) );
  XNOR U17783 ( .A(n19834), .B(n19835), .Z(n16994) );
  AND U17784 ( .A(n19834), .B(n19836), .Z(n19835) );
  XNOR U17785 ( .A(n19837), .B(n19838), .Z(n16997) );
  AND U17786 ( .A(n19837), .B(n19839), .Z(n19838) );
  XNOR U17787 ( .A(n19840), .B(n19841), .Z(n17000) );
  AND U17788 ( .A(n19840), .B(n19842), .Z(n19841) );
  XNOR U17789 ( .A(n19843), .B(n19844), .Z(n17003) );
  AND U17790 ( .A(n19843), .B(n19845), .Z(n19844) );
  XNOR U17791 ( .A(n19846), .B(n19847), .Z(n17006) );
  AND U17792 ( .A(n19846), .B(n19848), .Z(n19847) );
  XNOR U17793 ( .A(n19849), .B(n19850), .Z(n17009) );
  AND U17794 ( .A(n19849), .B(n19851), .Z(n19850) );
  IV U17795 ( .A(n17014), .Z(n17012) );
  XNOR U17796 ( .A(n19852), .B(n19853), .Z(n17014) );
  AND U17797 ( .A(n19852), .B(n130), .Z(n19853) );
  XOR U17798 ( .A(n19854), .B(n19855), .Z(n17015) );
  AND U17799 ( .A(n19856), .B(n19857), .Z(n19855) );
  XOR U17800 ( .A(n134), .B(n19854), .Z(n19857) );
  XOR U17801 ( .A(n18433), .B(n18434), .Z(n134) );
  AND U17802 ( .A(n19858), .B(n19859), .Z(n18434) );
  XOR U17803 ( .A(n18430), .B(n18431), .Z(n18433) );
  AND U17804 ( .A(n19860), .B(n19861), .Z(n18431) );
  XOR U17805 ( .A(n18427), .B(n18428), .Z(n18430) );
  AND U17806 ( .A(n19862), .B(n19863), .Z(n18428) );
  XOR U17807 ( .A(n18424), .B(n18425), .Z(n18427) );
  AND U17808 ( .A(n19864), .B(n19865), .Z(n18425) );
  XOR U17809 ( .A(n18421), .B(n18422), .Z(n18424) );
  AND U17810 ( .A(n19866), .B(n19867), .Z(n18422) );
  XOR U17811 ( .A(n18418), .B(n18419), .Z(n18421) );
  AND U17812 ( .A(n19868), .B(n19869), .Z(n18419) );
  XOR U17813 ( .A(n18415), .B(n18416), .Z(n18418) );
  AND U17814 ( .A(n19870), .B(n19871), .Z(n18416) );
  XOR U17815 ( .A(n18412), .B(n18413), .Z(n18415) );
  AND U17816 ( .A(n19872), .B(n19873), .Z(n18413) );
  XOR U17817 ( .A(n18409), .B(n18410), .Z(n18412) );
  AND U17818 ( .A(n19874), .B(n19875), .Z(n18410) );
  XOR U17819 ( .A(n18406), .B(n18407), .Z(n18409) );
  AND U17820 ( .A(n19876), .B(n19877), .Z(n18407) );
  XOR U17821 ( .A(n18403), .B(n18404), .Z(n18406) );
  AND U17822 ( .A(n19878), .B(n19879), .Z(n18404) );
  XOR U17823 ( .A(n18400), .B(n18401), .Z(n18403) );
  AND U17824 ( .A(n19880), .B(n19881), .Z(n18401) );
  XOR U17825 ( .A(n18397), .B(n18398), .Z(n18400) );
  AND U17826 ( .A(n19882), .B(n19883), .Z(n18398) );
  XOR U17827 ( .A(n18394), .B(n18395), .Z(n18397) );
  AND U17828 ( .A(n19884), .B(n19885), .Z(n18395) );
  XOR U17829 ( .A(n18391), .B(n18392), .Z(n18394) );
  AND U17830 ( .A(n19886), .B(n19887), .Z(n18392) );
  XOR U17831 ( .A(n18388), .B(n18389), .Z(n18391) );
  AND U17832 ( .A(n19888), .B(n19889), .Z(n18389) );
  XOR U17833 ( .A(n18385), .B(n18386), .Z(n18388) );
  AND U17834 ( .A(n19890), .B(n19891), .Z(n18386) );
  XOR U17835 ( .A(n18382), .B(n18383), .Z(n18385) );
  AND U17836 ( .A(n19892), .B(n19893), .Z(n18383) );
  XOR U17837 ( .A(n18379), .B(n18380), .Z(n18382) );
  AND U17838 ( .A(n19894), .B(n19895), .Z(n18380) );
  XOR U17839 ( .A(n18376), .B(n18377), .Z(n18379) );
  AND U17840 ( .A(n19896), .B(n19897), .Z(n18377) );
  XOR U17841 ( .A(n18373), .B(n18374), .Z(n18376) );
  AND U17842 ( .A(n19898), .B(n19899), .Z(n18374) );
  XOR U17843 ( .A(n18370), .B(n18371), .Z(n18373) );
  AND U17844 ( .A(n19900), .B(n19901), .Z(n18371) );
  XOR U17845 ( .A(n18367), .B(n18368), .Z(n18370) );
  AND U17846 ( .A(n19902), .B(n19903), .Z(n18368) );
  XOR U17847 ( .A(n18364), .B(n18365), .Z(n18367) );
  AND U17848 ( .A(n19904), .B(n19905), .Z(n18365) );
  XOR U17849 ( .A(n18361), .B(n18362), .Z(n18364) );
  AND U17850 ( .A(n19906), .B(n19907), .Z(n18362) );
  XOR U17851 ( .A(n18358), .B(n18359), .Z(n18361) );
  AND U17852 ( .A(n19908), .B(n19909), .Z(n18359) );
  XOR U17853 ( .A(n18355), .B(n18356), .Z(n18358) );
  AND U17854 ( .A(n19910), .B(n19911), .Z(n18356) );
  XOR U17855 ( .A(n18352), .B(n18353), .Z(n18355) );
  AND U17856 ( .A(n19912), .B(n19913), .Z(n18353) );
  XOR U17857 ( .A(n18349), .B(n18350), .Z(n18352) );
  AND U17858 ( .A(n19914), .B(n19915), .Z(n18350) );
  XOR U17859 ( .A(n18346), .B(n18347), .Z(n18349) );
  AND U17860 ( .A(n19916), .B(n19917), .Z(n18347) );
  XOR U17861 ( .A(n18343), .B(n18344), .Z(n18346) );
  AND U17862 ( .A(n19918), .B(n19919), .Z(n18344) );
  XOR U17863 ( .A(n18340), .B(n18341), .Z(n18343) );
  AND U17864 ( .A(n19920), .B(n19921), .Z(n18341) );
  XOR U17865 ( .A(n18337), .B(n18338), .Z(n18340) );
  AND U17866 ( .A(n19922), .B(n19923), .Z(n18338) );
  XOR U17867 ( .A(n18334), .B(n18335), .Z(n18337) );
  AND U17868 ( .A(n19924), .B(n19925), .Z(n18335) );
  XOR U17869 ( .A(n18331), .B(n18332), .Z(n18334) );
  AND U17870 ( .A(n19926), .B(n19927), .Z(n18332) );
  XOR U17871 ( .A(n18328), .B(n18329), .Z(n18331) );
  AND U17872 ( .A(n19928), .B(n19929), .Z(n18329) );
  XOR U17873 ( .A(n18325), .B(n18326), .Z(n18328) );
  AND U17874 ( .A(n19930), .B(n19931), .Z(n18326) );
  XOR U17875 ( .A(n18322), .B(n18323), .Z(n18325) );
  AND U17876 ( .A(n19932), .B(n19933), .Z(n18323) );
  XOR U17877 ( .A(n18319), .B(n18320), .Z(n18322) );
  AND U17878 ( .A(n19934), .B(n19935), .Z(n18320) );
  XOR U17879 ( .A(n18316), .B(n18317), .Z(n18319) );
  AND U17880 ( .A(n19936), .B(n19937), .Z(n18317) );
  XOR U17881 ( .A(n18313), .B(n18314), .Z(n18316) );
  AND U17882 ( .A(n19938), .B(n19939), .Z(n18314) );
  XOR U17883 ( .A(n18310), .B(n18311), .Z(n18313) );
  AND U17884 ( .A(n19940), .B(n19941), .Z(n18311) );
  XOR U17885 ( .A(n18307), .B(n18308), .Z(n18310) );
  AND U17886 ( .A(n19942), .B(n19943), .Z(n18308) );
  XOR U17887 ( .A(n18304), .B(n18305), .Z(n18307) );
  AND U17888 ( .A(n19944), .B(n19945), .Z(n18305) );
  XOR U17889 ( .A(n18301), .B(n18302), .Z(n18304) );
  AND U17890 ( .A(n19946), .B(n19947), .Z(n18302) );
  XOR U17891 ( .A(n18298), .B(n18299), .Z(n18301) );
  AND U17892 ( .A(n19948), .B(n19949), .Z(n18299) );
  XOR U17893 ( .A(n18295), .B(n18296), .Z(n18298) );
  AND U17894 ( .A(n19950), .B(n19951), .Z(n18296) );
  XOR U17895 ( .A(n18292), .B(n18293), .Z(n18295) );
  AND U17896 ( .A(n19952), .B(n19953), .Z(n18293) );
  XOR U17897 ( .A(n18289), .B(n18290), .Z(n18292) );
  AND U17898 ( .A(n19954), .B(n19955), .Z(n18290) );
  XOR U17899 ( .A(n18286), .B(n18287), .Z(n18289) );
  AND U17900 ( .A(n19956), .B(n19957), .Z(n18287) );
  XOR U17901 ( .A(n18283), .B(n18284), .Z(n18286) );
  AND U17902 ( .A(n19958), .B(n19959), .Z(n18284) );
  XOR U17903 ( .A(n18280), .B(n18281), .Z(n18283) );
  AND U17904 ( .A(n19960), .B(n19961), .Z(n18281) );
  XOR U17905 ( .A(n18277), .B(n18278), .Z(n18280) );
  AND U17906 ( .A(n19962), .B(n19963), .Z(n18278) );
  XOR U17907 ( .A(n18274), .B(n18275), .Z(n18277) );
  AND U17908 ( .A(n19964), .B(n19965), .Z(n18275) );
  XOR U17909 ( .A(n18271), .B(n18272), .Z(n18274) );
  AND U17910 ( .A(n19966), .B(n19967), .Z(n18272) );
  XOR U17911 ( .A(n18268), .B(n18269), .Z(n18271) );
  AND U17912 ( .A(n19968), .B(n19969), .Z(n18269) );
  XOR U17913 ( .A(n18265), .B(n18266), .Z(n18268) );
  AND U17914 ( .A(n19970), .B(n19971), .Z(n18266) );
  XOR U17915 ( .A(n18262), .B(n18263), .Z(n18265) );
  AND U17916 ( .A(n19972), .B(n19973), .Z(n18263) );
  XOR U17917 ( .A(n18259), .B(n18260), .Z(n18262) );
  AND U17918 ( .A(n19974), .B(n19975), .Z(n18260) );
  XOR U17919 ( .A(n18256), .B(n18257), .Z(n18259) );
  AND U17920 ( .A(n19976), .B(n19977), .Z(n18257) );
  XOR U17921 ( .A(n18253), .B(n18254), .Z(n18256) );
  AND U17922 ( .A(n19978), .B(n19979), .Z(n18254) );
  XOR U17923 ( .A(n18250), .B(n18251), .Z(n18253) );
  AND U17924 ( .A(n19980), .B(n19981), .Z(n18251) );
  XOR U17925 ( .A(n18247), .B(n18248), .Z(n18250) );
  AND U17926 ( .A(n19982), .B(n19983), .Z(n18248) );
  XOR U17927 ( .A(n18244), .B(n18245), .Z(n18247) );
  AND U17928 ( .A(n19984), .B(n19985), .Z(n18245) );
  XOR U17929 ( .A(n18241), .B(n18242), .Z(n18244) );
  AND U17930 ( .A(n19986), .B(n19987), .Z(n18242) );
  XOR U17931 ( .A(n18238), .B(n18239), .Z(n18241) );
  AND U17932 ( .A(n19988), .B(n19989), .Z(n18239) );
  XOR U17933 ( .A(n18235), .B(n18236), .Z(n18238) );
  AND U17934 ( .A(n19990), .B(n19991), .Z(n18236) );
  XOR U17935 ( .A(n18232), .B(n18233), .Z(n18235) );
  AND U17936 ( .A(n19992), .B(n19993), .Z(n18233) );
  XOR U17937 ( .A(n18229), .B(n18230), .Z(n18232) );
  AND U17938 ( .A(n19994), .B(n19995), .Z(n18230) );
  XOR U17939 ( .A(n18226), .B(n18227), .Z(n18229) );
  AND U17940 ( .A(n19996), .B(n19997), .Z(n18227) );
  XOR U17941 ( .A(n18223), .B(n18224), .Z(n18226) );
  AND U17942 ( .A(n19998), .B(n19999), .Z(n18224) );
  XOR U17943 ( .A(n18220), .B(n18221), .Z(n18223) );
  AND U17944 ( .A(n20000), .B(n20001), .Z(n18221) );
  XOR U17945 ( .A(n18217), .B(n18218), .Z(n18220) );
  AND U17946 ( .A(n20002), .B(n20003), .Z(n18218) );
  XOR U17947 ( .A(n18214), .B(n18215), .Z(n18217) );
  AND U17948 ( .A(n20004), .B(n20005), .Z(n18215) );
  XOR U17949 ( .A(n18211), .B(n18212), .Z(n18214) );
  AND U17950 ( .A(n20006), .B(n20007), .Z(n18212) );
  XOR U17951 ( .A(n18208), .B(n18209), .Z(n18211) );
  AND U17952 ( .A(n20008), .B(n20009), .Z(n18209) );
  XOR U17953 ( .A(n18205), .B(n18206), .Z(n18208) );
  AND U17954 ( .A(n20010), .B(n20011), .Z(n18206) );
  XOR U17955 ( .A(n18202), .B(n18203), .Z(n18205) );
  AND U17956 ( .A(n20012), .B(n20013), .Z(n18203) );
  XOR U17957 ( .A(n18199), .B(n18200), .Z(n18202) );
  AND U17958 ( .A(n20014), .B(n20015), .Z(n18200) );
  XOR U17959 ( .A(n18196), .B(n18197), .Z(n18199) );
  AND U17960 ( .A(n20016), .B(n20017), .Z(n18197) );
  XOR U17961 ( .A(n18193), .B(n18194), .Z(n18196) );
  AND U17962 ( .A(n20018), .B(n20019), .Z(n18194) );
  XOR U17963 ( .A(n18190), .B(n18191), .Z(n18193) );
  AND U17964 ( .A(n20020), .B(n20021), .Z(n18191) );
  XOR U17965 ( .A(n18187), .B(n18188), .Z(n18190) );
  AND U17966 ( .A(n20022), .B(n20023), .Z(n18188) );
  XOR U17967 ( .A(n18184), .B(n18185), .Z(n18187) );
  AND U17968 ( .A(n20024), .B(n20025), .Z(n18185) );
  XOR U17969 ( .A(n18181), .B(n18182), .Z(n18184) );
  AND U17970 ( .A(n20026), .B(n20027), .Z(n18182) );
  XOR U17971 ( .A(n18178), .B(n18179), .Z(n18181) );
  AND U17972 ( .A(n20028), .B(n20029), .Z(n18179) );
  XOR U17973 ( .A(n18175), .B(n18176), .Z(n18178) );
  AND U17974 ( .A(n20030), .B(n20031), .Z(n18176) );
  XOR U17975 ( .A(n18172), .B(n18173), .Z(n18175) );
  AND U17976 ( .A(n20032), .B(n20033), .Z(n18173) );
  XOR U17977 ( .A(n18169), .B(n18170), .Z(n18172) );
  AND U17978 ( .A(n20034), .B(n20035), .Z(n18170) );
  XOR U17979 ( .A(n18166), .B(n18167), .Z(n18169) );
  AND U17980 ( .A(n20036), .B(n20037), .Z(n18167) );
  XOR U17981 ( .A(n18163), .B(n18164), .Z(n18166) );
  AND U17982 ( .A(n20038), .B(n20039), .Z(n18164) );
  XOR U17983 ( .A(n18160), .B(n18161), .Z(n18163) );
  AND U17984 ( .A(n20040), .B(n20041), .Z(n18161) );
  XOR U17985 ( .A(n18157), .B(n18158), .Z(n18160) );
  AND U17986 ( .A(n20042), .B(n20043), .Z(n18158) );
  XOR U17987 ( .A(n18154), .B(n18155), .Z(n18157) );
  AND U17988 ( .A(n20044), .B(n20045), .Z(n18155) );
  XOR U17989 ( .A(n18151), .B(n18152), .Z(n18154) );
  AND U17990 ( .A(n20046), .B(n20047), .Z(n18152) );
  XOR U17991 ( .A(n18148), .B(n18149), .Z(n18151) );
  AND U17992 ( .A(n20048), .B(n20049), .Z(n18149) );
  XOR U17993 ( .A(n18145), .B(n18146), .Z(n18148) );
  AND U17994 ( .A(n20050), .B(n20051), .Z(n18146) );
  XOR U17995 ( .A(n18142), .B(n18143), .Z(n18145) );
  AND U17996 ( .A(n20052), .B(n20053), .Z(n18143) );
  XOR U17997 ( .A(n18139), .B(n18140), .Z(n18142) );
  AND U17998 ( .A(n20054), .B(n20055), .Z(n18140) );
  XOR U17999 ( .A(n18136), .B(n18137), .Z(n18139) );
  AND U18000 ( .A(n20056), .B(n20057), .Z(n18137) );
  XOR U18001 ( .A(n18133), .B(n18134), .Z(n18136) );
  AND U18002 ( .A(n20058), .B(n20059), .Z(n18134) );
  XOR U18003 ( .A(n18130), .B(n18131), .Z(n18133) );
  AND U18004 ( .A(n20060), .B(n20061), .Z(n18131) );
  XOR U18005 ( .A(n18127), .B(n18128), .Z(n18130) );
  AND U18006 ( .A(n20062), .B(n20063), .Z(n18128) );
  XOR U18007 ( .A(n18124), .B(n18125), .Z(n18127) );
  AND U18008 ( .A(n20064), .B(n20065), .Z(n18125) );
  XOR U18009 ( .A(n18121), .B(n18122), .Z(n18124) );
  AND U18010 ( .A(n20066), .B(n20067), .Z(n18122) );
  XOR U18011 ( .A(n18118), .B(n18119), .Z(n18121) );
  AND U18012 ( .A(n20068), .B(n20069), .Z(n18119) );
  XOR U18013 ( .A(n18115), .B(n18116), .Z(n18118) );
  AND U18014 ( .A(n20070), .B(n20071), .Z(n18116) );
  XOR U18015 ( .A(n18112), .B(n18113), .Z(n18115) );
  AND U18016 ( .A(n20072), .B(n20073), .Z(n18113) );
  XOR U18017 ( .A(n18109), .B(n18110), .Z(n18112) );
  AND U18018 ( .A(n20074), .B(n20075), .Z(n18110) );
  XOR U18019 ( .A(n18106), .B(n18107), .Z(n18109) );
  AND U18020 ( .A(n20076), .B(n20077), .Z(n18107) );
  XOR U18021 ( .A(n18103), .B(n18104), .Z(n18106) );
  AND U18022 ( .A(n20078), .B(n20079), .Z(n18104) );
  XOR U18023 ( .A(n18100), .B(n18101), .Z(n18103) );
  AND U18024 ( .A(n20080), .B(n20081), .Z(n18101) );
  XOR U18025 ( .A(n18097), .B(n18098), .Z(n18100) );
  AND U18026 ( .A(n20082), .B(n20083), .Z(n18098) );
  XOR U18027 ( .A(n18094), .B(n18095), .Z(n18097) );
  AND U18028 ( .A(n20084), .B(n20085), .Z(n18095) );
  XOR U18029 ( .A(n18091), .B(n18092), .Z(n18094) );
  AND U18030 ( .A(n20086), .B(n20087), .Z(n18092) );
  XOR U18031 ( .A(n18088), .B(n18089), .Z(n18091) );
  AND U18032 ( .A(n20088), .B(n20089), .Z(n18089) );
  XOR U18033 ( .A(n18085), .B(n18086), .Z(n18088) );
  AND U18034 ( .A(n20090), .B(n20091), .Z(n18086) );
  XOR U18035 ( .A(n18082), .B(n18083), .Z(n18085) );
  AND U18036 ( .A(n20092), .B(n20093), .Z(n18083) );
  XOR U18037 ( .A(n18079), .B(n18080), .Z(n18082) );
  AND U18038 ( .A(n20094), .B(n20095), .Z(n18080) );
  XOR U18039 ( .A(n18076), .B(n18077), .Z(n18079) );
  AND U18040 ( .A(n20096), .B(n20097), .Z(n18077) );
  XOR U18041 ( .A(n18073), .B(n18074), .Z(n18076) );
  AND U18042 ( .A(n20098), .B(n20099), .Z(n18074) );
  XOR U18043 ( .A(n18070), .B(n18071), .Z(n18073) );
  AND U18044 ( .A(n20100), .B(n20101), .Z(n18071) );
  XOR U18045 ( .A(n18067), .B(n18068), .Z(n18070) );
  AND U18046 ( .A(n20102), .B(n20103), .Z(n18068) );
  XOR U18047 ( .A(n18064), .B(n18065), .Z(n18067) );
  AND U18048 ( .A(n20104), .B(n20105), .Z(n18065) );
  XOR U18049 ( .A(n18061), .B(n18062), .Z(n18064) );
  AND U18050 ( .A(n20106), .B(n20107), .Z(n18062) );
  XOR U18051 ( .A(n18058), .B(n18059), .Z(n18061) );
  AND U18052 ( .A(n20108), .B(n20109), .Z(n18059) );
  XOR U18053 ( .A(n18055), .B(n18056), .Z(n18058) );
  AND U18054 ( .A(n20110), .B(n20111), .Z(n18056) );
  XOR U18055 ( .A(n18052), .B(n18053), .Z(n18055) );
  AND U18056 ( .A(n20112), .B(n20113), .Z(n18053) );
  XOR U18057 ( .A(n18049), .B(n18050), .Z(n18052) );
  AND U18058 ( .A(n20114), .B(n20115), .Z(n18050) );
  XOR U18059 ( .A(n18046), .B(n18047), .Z(n18049) );
  AND U18060 ( .A(n20116), .B(n20117), .Z(n18047) );
  XOR U18061 ( .A(n18043), .B(n18044), .Z(n18046) );
  AND U18062 ( .A(n20118), .B(n20119), .Z(n18044) );
  XOR U18063 ( .A(n18040), .B(n18041), .Z(n18043) );
  AND U18064 ( .A(n20120), .B(n20121), .Z(n18041) );
  XOR U18065 ( .A(n18037), .B(n18038), .Z(n18040) );
  AND U18066 ( .A(n20122), .B(n20123), .Z(n18038) );
  XOR U18067 ( .A(n18034), .B(n18035), .Z(n18037) );
  AND U18068 ( .A(n20124), .B(n20125), .Z(n18035) );
  XOR U18069 ( .A(n18031), .B(n18032), .Z(n18034) );
  AND U18070 ( .A(n20126), .B(n20127), .Z(n18032) );
  XOR U18071 ( .A(n18028), .B(n18029), .Z(n18031) );
  AND U18072 ( .A(n20128), .B(n20129), .Z(n18029) );
  XOR U18073 ( .A(n18025), .B(n18026), .Z(n18028) );
  AND U18074 ( .A(n20130), .B(n20131), .Z(n18026) );
  XOR U18075 ( .A(n18022), .B(n18023), .Z(n18025) );
  AND U18076 ( .A(n20132), .B(n20133), .Z(n18023) );
  XOR U18077 ( .A(n18019), .B(n18020), .Z(n18022) );
  AND U18078 ( .A(n20134), .B(n20135), .Z(n18020) );
  XOR U18079 ( .A(n18016), .B(n18017), .Z(n18019) );
  AND U18080 ( .A(n20136), .B(n20137), .Z(n18017) );
  XOR U18081 ( .A(n18013), .B(n18014), .Z(n18016) );
  AND U18082 ( .A(n20138), .B(n20139), .Z(n18014) );
  XOR U18083 ( .A(n18010), .B(n18011), .Z(n18013) );
  AND U18084 ( .A(n20140), .B(n20141), .Z(n18011) );
  XOR U18085 ( .A(n18007), .B(n18008), .Z(n18010) );
  AND U18086 ( .A(n20142), .B(n20143), .Z(n18008) );
  XOR U18087 ( .A(n18004), .B(n18005), .Z(n18007) );
  AND U18088 ( .A(n20144), .B(n20145), .Z(n18005) );
  XOR U18089 ( .A(n18001), .B(n18002), .Z(n18004) );
  AND U18090 ( .A(n20146), .B(n20147), .Z(n18002) );
  XOR U18091 ( .A(n17998), .B(n17999), .Z(n18001) );
  AND U18092 ( .A(n20148), .B(n20149), .Z(n17999) );
  XOR U18093 ( .A(n17995), .B(n17996), .Z(n17998) );
  AND U18094 ( .A(n20150), .B(n20151), .Z(n17996) );
  XOR U18095 ( .A(n17992), .B(n17993), .Z(n17995) );
  AND U18096 ( .A(n20152), .B(n20153), .Z(n17993) );
  XOR U18097 ( .A(n17989), .B(n17990), .Z(n17992) );
  AND U18098 ( .A(n20154), .B(n20155), .Z(n17990) );
  XOR U18099 ( .A(n17986), .B(n17987), .Z(n17989) );
  AND U18100 ( .A(n20156), .B(n20157), .Z(n17987) );
  XOR U18101 ( .A(n17983), .B(n17984), .Z(n17986) );
  AND U18102 ( .A(n20158), .B(n20159), .Z(n17984) );
  XOR U18103 ( .A(n17980), .B(n17981), .Z(n17983) );
  AND U18104 ( .A(n20160), .B(n20161), .Z(n17981) );
  XOR U18105 ( .A(n17977), .B(n17978), .Z(n17980) );
  AND U18106 ( .A(n20162), .B(n20163), .Z(n17978) );
  XOR U18107 ( .A(n17974), .B(n17975), .Z(n17977) );
  AND U18108 ( .A(n20164), .B(n20165), .Z(n17975) );
  XOR U18109 ( .A(n17971), .B(n17972), .Z(n17974) );
  AND U18110 ( .A(n20166), .B(n20167), .Z(n17972) );
  XOR U18111 ( .A(n17968), .B(n17969), .Z(n17971) );
  AND U18112 ( .A(n20168), .B(n20169), .Z(n17969) );
  XOR U18113 ( .A(n17965), .B(n17966), .Z(n17968) );
  AND U18114 ( .A(n20170), .B(n20171), .Z(n17966) );
  XOR U18115 ( .A(n17962), .B(n17963), .Z(n17965) );
  AND U18116 ( .A(n20172), .B(n20173), .Z(n17963) );
  XOR U18117 ( .A(n17959), .B(n17960), .Z(n17962) );
  AND U18118 ( .A(n20174), .B(n20175), .Z(n17960) );
  XOR U18119 ( .A(n17956), .B(n17957), .Z(n17959) );
  AND U18120 ( .A(n20176), .B(n20177), .Z(n17957) );
  XOR U18121 ( .A(n17953), .B(n17954), .Z(n17956) );
  AND U18122 ( .A(n20178), .B(n20179), .Z(n17954) );
  XOR U18123 ( .A(n17950), .B(n17951), .Z(n17953) );
  AND U18124 ( .A(n20180), .B(n20181), .Z(n17951) );
  XOR U18125 ( .A(n17947), .B(n17948), .Z(n17950) );
  AND U18126 ( .A(n20182), .B(n20183), .Z(n17948) );
  XOR U18127 ( .A(n17944), .B(n17945), .Z(n17947) );
  AND U18128 ( .A(n20184), .B(n20185), .Z(n17945) );
  XOR U18129 ( .A(n17941), .B(n17942), .Z(n17944) );
  AND U18130 ( .A(n20186), .B(n20187), .Z(n17942) );
  XOR U18131 ( .A(n17938), .B(n17939), .Z(n17941) );
  AND U18132 ( .A(n20188), .B(n20189), .Z(n17939) );
  XOR U18133 ( .A(n17935), .B(n17936), .Z(n17938) );
  AND U18134 ( .A(n20190), .B(n20191), .Z(n17936) );
  XOR U18135 ( .A(n17932), .B(n17933), .Z(n17935) );
  AND U18136 ( .A(n20192), .B(n20193), .Z(n17933) );
  XOR U18137 ( .A(n17929), .B(n17930), .Z(n17932) );
  AND U18138 ( .A(n20194), .B(n20195), .Z(n17930) );
  XOR U18139 ( .A(n17926), .B(n17927), .Z(n17929) );
  AND U18140 ( .A(n20196), .B(n20197), .Z(n17927) );
  XOR U18141 ( .A(n17923), .B(n17924), .Z(n17926) );
  AND U18142 ( .A(n20198), .B(n20199), .Z(n17924) );
  XOR U18143 ( .A(n17920), .B(n17921), .Z(n17923) );
  AND U18144 ( .A(n20200), .B(n20201), .Z(n17921) );
  XOR U18145 ( .A(n17917), .B(n17918), .Z(n17920) );
  AND U18146 ( .A(n20202), .B(n20203), .Z(n17918) );
  XOR U18147 ( .A(n17914), .B(n17915), .Z(n17917) );
  AND U18148 ( .A(n20204), .B(n20205), .Z(n17915) );
  XOR U18149 ( .A(n17911), .B(n17912), .Z(n17914) );
  AND U18150 ( .A(n20206), .B(n20207), .Z(n17912) );
  XOR U18151 ( .A(n17908), .B(n17909), .Z(n17911) );
  AND U18152 ( .A(n20208), .B(n20209), .Z(n17909) );
  XOR U18153 ( .A(n17905), .B(n17906), .Z(n17908) );
  AND U18154 ( .A(n20210), .B(n20211), .Z(n17906) );
  XOR U18155 ( .A(n17902), .B(n17903), .Z(n17905) );
  AND U18156 ( .A(n20212), .B(n20213), .Z(n17903) );
  XOR U18157 ( .A(n17899), .B(n17900), .Z(n17902) );
  AND U18158 ( .A(n20214), .B(n20215), .Z(n17900) );
  XOR U18159 ( .A(n17896), .B(n17897), .Z(n17899) );
  AND U18160 ( .A(n20216), .B(n20217), .Z(n17897) );
  XOR U18161 ( .A(n17893), .B(n17894), .Z(n17896) );
  AND U18162 ( .A(n20218), .B(n20219), .Z(n17894) );
  XOR U18163 ( .A(n17890), .B(n17891), .Z(n17893) );
  AND U18164 ( .A(n20220), .B(n20221), .Z(n17891) );
  XOR U18165 ( .A(n17887), .B(n17888), .Z(n17890) );
  AND U18166 ( .A(n20222), .B(n20223), .Z(n17888) );
  XOR U18167 ( .A(n17884), .B(n17885), .Z(n17887) );
  AND U18168 ( .A(n20224), .B(n20225), .Z(n17885) );
  XOR U18169 ( .A(n17881), .B(n17882), .Z(n17884) );
  AND U18170 ( .A(n20226), .B(n20227), .Z(n17882) );
  XOR U18171 ( .A(n17878), .B(n17879), .Z(n17881) );
  AND U18172 ( .A(n20228), .B(n20229), .Z(n17879) );
  XOR U18173 ( .A(n17875), .B(n17876), .Z(n17878) );
  AND U18174 ( .A(n20230), .B(n20231), .Z(n17876) );
  XOR U18175 ( .A(n17872), .B(n17873), .Z(n17875) );
  AND U18176 ( .A(n20232), .B(n20233), .Z(n17873) );
  XOR U18177 ( .A(n17869), .B(n17870), .Z(n17872) );
  AND U18178 ( .A(n20234), .B(n20235), .Z(n17870) );
  XOR U18179 ( .A(n17866), .B(n17867), .Z(n17869) );
  AND U18180 ( .A(n20236), .B(n20237), .Z(n17867) );
  XOR U18181 ( .A(n17863), .B(n17864), .Z(n17866) );
  AND U18182 ( .A(n20238), .B(n20239), .Z(n17864) );
  XOR U18183 ( .A(n17860), .B(n17861), .Z(n17863) );
  AND U18184 ( .A(n20240), .B(n20241), .Z(n17861) );
  XOR U18185 ( .A(n17857), .B(n17858), .Z(n17860) );
  AND U18186 ( .A(n20242), .B(n20243), .Z(n17858) );
  XOR U18187 ( .A(n17854), .B(n17855), .Z(n17857) );
  AND U18188 ( .A(n20244), .B(n20245), .Z(n17855) );
  XOR U18189 ( .A(n17851), .B(n17852), .Z(n17854) );
  AND U18190 ( .A(n20246), .B(n20247), .Z(n17852) );
  XOR U18191 ( .A(n17848), .B(n17849), .Z(n17851) );
  AND U18192 ( .A(n20248), .B(n20249), .Z(n17849) );
  XOR U18193 ( .A(n17845), .B(n17846), .Z(n17848) );
  AND U18194 ( .A(n20250), .B(n20251), .Z(n17846) );
  XOR U18195 ( .A(n17842), .B(n17843), .Z(n17845) );
  AND U18196 ( .A(n20252), .B(n20253), .Z(n17843) );
  XOR U18197 ( .A(n17839), .B(n17840), .Z(n17842) );
  AND U18198 ( .A(n20254), .B(n20255), .Z(n17840) );
  XOR U18199 ( .A(n17836), .B(n17837), .Z(n17839) );
  AND U18200 ( .A(n20256), .B(n20257), .Z(n17837) );
  XOR U18201 ( .A(n17833), .B(n17834), .Z(n17836) );
  AND U18202 ( .A(n20258), .B(n20259), .Z(n17834) );
  XOR U18203 ( .A(n17830), .B(n17831), .Z(n17833) );
  AND U18204 ( .A(n20260), .B(n20261), .Z(n17831) );
  XOR U18205 ( .A(n17827), .B(n17828), .Z(n17830) );
  AND U18206 ( .A(n20262), .B(n20263), .Z(n17828) );
  XOR U18207 ( .A(n17824), .B(n17825), .Z(n17827) );
  AND U18208 ( .A(n20264), .B(n20265), .Z(n17825) );
  XOR U18209 ( .A(n17821), .B(n17822), .Z(n17824) );
  AND U18210 ( .A(n20266), .B(n20267), .Z(n17822) );
  XOR U18211 ( .A(n17818), .B(n17819), .Z(n17821) );
  AND U18212 ( .A(n20268), .B(n20269), .Z(n17819) );
  XOR U18213 ( .A(n17815), .B(n17816), .Z(n17818) );
  AND U18214 ( .A(n20270), .B(n20271), .Z(n17816) );
  XOR U18215 ( .A(n17812), .B(n17813), .Z(n17815) );
  AND U18216 ( .A(n20272), .B(n20273), .Z(n17813) );
  XOR U18217 ( .A(n17809), .B(n17810), .Z(n17812) );
  AND U18218 ( .A(n20274), .B(n20275), .Z(n17810) );
  XOR U18219 ( .A(n17806), .B(n17807), .Z(n17809) );
  AND U18220 ( .A(n20276), .B(n20277), .Z(n17807) );
  XOR U18221 ( .A(n17803), .B(n17804), .Z(n17806) );
  AND U18222 ( .A(n20278), .B(n20279), .Z(n17804) );
  XOR U18223 ( .A(n17800), .B(n17801), .Z(n17803) );
  AND U18224 ( .A(n20280), .B(n20281), .Z(n17801) );
  XOR U18225 ( .A(n17797), .B(n17798), .Z(n17800) );
  AND U18226 ( .A(n20282), .B(n20283), .Z(n17798) );
  XOR U18227 ( .A(n17794), .B(n17795), .Z(n17797) );
  AND U18228 ( .A(n20284), .B(n20285), .Z(n17795) );
  XOR U18229 ( .A(n17791), .B(n17792), .Z(n17794) );
  AND U18230 ( .A(n20286), .B(n20287), .Z(n17792) );
  XOR U18231 ( .A(n17788), .B(n17789), .Z(n17791) );
  AND U18232 ( .A(n20288), .B(n20289), .Z(n17789) );
  XOR U18233 ( .A(n17785), .B(n17786), .Z(n17788) );
  AND U18234 ( .A(n20290), .B(n20291), .Z(n17786) );
  XOR U18235 ( .A(n17782), .B(n17783), .Z(n17785) );
  AND U18236 ( .A(n20292), .B(n20293), .Z(n17783) );
  XOR U18237 ( .A(n17779), .B(n17780), .Z(n17782) );
  AND U18238 ( .A(n20294), .B(n20295), .Z(n17780) );
  XOR U18239 ( .A(n17776), .B(n17777), .Z(n17779) );
  AND U18240 ( .A(n20296), .B(n20297), .Z(n17777) );
  XOR U18241 ( .A(n17773), .B(n17774), .Z(n17776) );
  AND U18242 ( .A(n20298), .B(n20299), .Z(n17774) );
  XOR U18243 ( .A(n17770), .B(n17771), .Z(n17773) );
  AND U18244 ( .A(n20300), .B(n20301), .Z(n17771) );
  XOR U18245 ( .A(n17767), .B(n17768), .Z(n17770) );
  AND U18246 ( .A(n20302), .B(n20303), .Z(n17768) );
  XOR U18247 ( .A(n17764), .B(n17765), .Z(n17767) );
  AND U18248 ( .A(n20304), .B(n20305), .Z(n17765) );
  XOR U18249 ( .A(n17761), .B(n17762), .Z(n17764) );
  AND U18250 ( .A(n20306), .B(n20307), .Z(n17762) );
  XOR U18251 ( .A(n17758), .B(n17759), .Z(n17761) );
  AND U18252 ( .A(n20308), .B(n20309), .Z(n17759) );
  XOR U18253 ( .A(n17755), .B(n17756), .Z(n17758) );
  AND U18254 ( .A(n20310), .B(n20311), .Z(n17756) );
  XOR U18255 ( .A(n17752), .B(n17753), .Z(n17755) );
  AND U18256 ( .A(n20312), .B(n20313), .Z(n17753) );
  XOR U18257 ( .A(n17749), .B(n17750), .Z(n17752) );
  AND U18258 ( .A(n20314), .B(n20315), .Z(n17750) );
  XOR U18259 ( .A(n17746), .B(n17747), .Z(n17749) );
  AND U18260 ( .A(n20316), .B(n20317), .Z(n17747) );
  XOR U18261 ( .A(n17743), .B(n17744), .Z(n17746) );
  AND U18262 ( .A(n20318), .B(n20319), .Z(n17744) );
  XOR U18263 ( .A(n17740), .B(n17741), .Z(n17743) );
  AND U18264 ( .A(n20320), .B(n20321), .Z(n17741) );
  XOR U18265 ( .A(n17737), .B(n17738), .Z(n17740) );
  AND U18266 ( .A(n20322), .B(n20323), .Z(n17738) );
  XOR U18267 ( .A(n17734), .B(n17735), .Z(n17737) );
  AND U18268 ( .A(n20324), .B(n20325), .Z(n17735) );
  XOR U18269 ( .A(n17731), .B(n17732), .Z(n17734) );
  AND U18270 ( .A(n20326), .B(n20327), .Z(n17732) );
  XOR U18271 ( .A(n17728), .B(n17729), .Z(n17731) );
  AND U18272 ( .A(n20328), .B(n20329), .Z(n17729) );
  XOR U18273 ( .A(n17725), .B(n17726), .Z(n17728) );
  AND U18274 ( .A(n20330), .B(n20331), .Z(n17726) );
  XOR U18275 ( .A(n17722), .B(n17723), .Z(n17725) );
  AND U18276 ( .A(n20332), .B(n20333), .Z(n17723) );
  XOR U18277 ( .A(n17719), .B(n17720), .Z(n17722) );
  AND U18278 ( .A(n20334), .B(n20335), .Z(n17720) );
  XOR U18279 ( .A(n17716), .B(n17717), .Z(n17719) );
  AND U18280 ( .A(n20336), .B(n20337), .Z(n17717) );
  XOR U18281 ( .A(n17713), .B(n17714), .Z(n17716) );
  AND U18282 ( .A(n20338), .B(n20339), .Z(n17714) );
  XOR U18283 ( .A(n17710), .B(n17711), .Z(n17713) );
  AND U18284 ( .A(n20340), .B(n20341), .Z(n17711) );
  XOR U18285 ( .A(n17707), .B(n17708), .Z(n17710) );
  AND U18286 ( .A(n20342), .B(n20343), .Z(n17708) );
  XOR U18287 ( .A(n17704), .B(n17705), .Z(n17707) );
  AND U18288 ( .A(n20344), .B(n20345), .Z(n17705) );
  XOR U18289 ( .A(n17701), .B(n17702), .Z(n17704) );
  AND U18290 ( .A(n20346), .B(n20347), .Z(n17702) );
  XOR U18291 ( .A(n17698), .B(n17699), .Z(n17701) );
  AND U18292 ( .A(n20348), .B(n20349), .Z(n17699) );
  XOR U18293 ( .A(n17695), .B(n17696), .Z(n17698) );
  AND U18294 ( .A(n20350), .B(n20351), .Z(n17696) );
  XOR U18295 ( .A(n17692), .B(n17693), .Z(n17695) );
  AND U18296 ( .A(n20352), .B(n20353), .Z(n17693) );
  XOR U18297 ( .A(n17689), .B(n17690), .Z(n17692) );
  AND U18298 ( .A(n20354), .B(n20355), .Z(n17690) );
  XOR U18299 ( .A(n17686), .B(n17687), .Z(n17689) );
  AND U18300 ( .A(n20356), .B(n20357), .Z(n17687) );
  XOR U18301 ( .A(n17683), .B(n17684), .Z(n17686) );
  AND U18302 ( .A(n20358), .B(n20359), .Z(n17684) );
  XOR U18303 ( .A(n17680), .B(n17681), .Z(n17683) );
  AND U18304 ( .A(n20360), .B(n20361), .Z(n17681) );
  XOR U18305 ( .A(n17677), .B(n17678), .Z(n17680) );
  AND U18306 ( .A(n20362), .B(n20363), .Z(n17678) );
  XOR U18307 ( .A(n17674), .B(n17675), .Z(n17677) );
  AND U18308 ( .A(n20364), .B(n20365), .Z(n17675) );
  XOR U18309 ( .A(n17671), .B(n17672), .Z(n17674) );
  AND U18310 ( .A(n20366), .B(n20367), .Z(n17672) );
  XOR U18311 ( .A(n17668), .B(n17669), .Z(n17671) );
  AND U18312 ( .A(n20368), .B(n20369), .Z(n17669) );
  XOR U18313 ( .A(n17665), .B(n17666), .Z(n17668) );
  AND U18314 ( .A(n20370), .B(n20371), .Z(n17666) );
  XOR U18315 ( .A(n17662), .B(n17663), .Z(n17665) );
  AND U18316 ( .A(n20372), .B(n20373), .Z(n17663) );
  XOR U18317 ( .A(n17659), .B(n17660), .Z(n17662) );
  AND U18318 ( .A(n20374), .B(n20375), .Z(n17660) );
  XOR U18319 ( .A(n17656), .B(n17657), .Z(n17659) );
  AND U18320 ( .A(n20376), .B(n20377), .Z(n17657) );
  XOR U18321 ( .A(n17653), .B(n17654), .Z(n17656) );
  AND U18322 ( .A(n20378), .B(n20379), .Z(n17654) );
  XOR U18323 ( .A(n17650), .B(n17651), .Z(n17653) );
  AND U18324 ( .A(n20380), .B(n20381), .Z(n17651) );
  XOR U18325 ( .A(n17647), .B(n17648), .Z(n17650) );
  AND U18326 ( .A(n20382), .B(n20383), .Z(n17648) );
  XOR U18327 ( .A(n17644), .B(n17645), .Z(n17647) );
  AND U18328 ( .A(n20384), .B(n20385), .Z(n17645) );
  XOR U18329 ( .A(n17641), .B(n17642), .Z(n17644) );
  AND U18330 ( .A(n20386), .B(n20387), .Z(n17642) );
  XOR U18331 ( .A(n17638), .B(n17639), .Z(n17641) );
  AND U18332 ( .A(n20388), .B(n20389), .Z(n17639) );
  XOR U18333 ( .A(n17635), .B(n17636), .Z(n17638) );
  AND U18334 ( .A(n20390), .B(n20391), .Z(n17636) );
  XOR U18335 ( .A(n17632), .B(n17633), .Z(n17635) );
  AND U18336 ( .A(n20392), .B(n20393), .Z(n17633) );
  XOR U18337 ( .A(n17629), .B(n17630), .Z(n17632) );
  AND U18338 ( .A(n20394), .B(n20395), .Z(n17630) );
  XOR U18339 ( .A(n17626), .B(n17627), .Z(n17629) );
  AND U18340 ( .A(n20396), .B(n20397), .Z(n17627) );
  XOR U18341 ( .A(n17623), .B(n17624), .Z(n17626) );
  AND U18342 ( .A(n20398), .B(n20399), .Z(n17624) );
  XOR U18343 ( .A(n17620), .B(n17621), .Z(n17623) );
  AND U18344 ( .A(n20400), .B(n20401), .Z(n17621) );
  XOR U18345 ( .A(n17617), .B(n17618), .Z(n17620) );
  AND U18346 ( .A(n20402), .B(n20403), .Z(n17618) );
  XOR U18347 ( .A(n17614), .B(n17615), .Z(n17617) );
  AND U18348 ( .A(n20404), .B(n20405), .Z(n17615) );
  XOR U18349 ( .A(n17611), .B(n17612), .Z(n17614) );
  AND U18350 ( .A(n20406), .B(n20407), .Z(n17612) );
  XOR U18351 ( .A(n17608), .B(n17609), .Z(n17611) );
  AND U18352 ( .A(n20408), .B(n20409), .Z(n17609) );
  XOR U18353 ( .A(n17605), .B(n17606), .Z(n17608) );
  AND U18354 ( .A(n20410), .B(n20411), .Z(n17606) );
  XOR U18355 ( .A(n17602), .B(n17603), .Z(n17605) );
  AND U18356 ( .A(n20412), .B(n20413), .Z(n17603) );
  XOR U18357 ( .A(n17599), .B(n17600), .Z(n17602) );
  AND U18358 ( .A(n20414), .B(n20415), .Z(n17600) );
  XOR U18359 ( .A(n17596), .B(n17597), .Z(n17599) );
  AND U18360 ( .A(n20416), .B(n20417), .Z(n17597) );
  XOR U18361 ( .A(n17593), .B(n17594), .Z(n17596) );
  AND U18362 ( .A(n20418), .B(n20419), .Z(n17594) );
  XOR U18363 ( .A(n17590), .B(n17591), .Z(n17593) );
  AND U18364 ( .A(n20420), .B(n20421), .Z(n17591) );
  XOR U18365 ( .A(n17587), .B(n17588), .Z(n17590) );
  AND U18366 ( .A(n20422), .B(n20423), .Z(n17588) );
  XOR U18367 ( .A(n17584), .B(n17585), .Z(n17587) );
  AND U18368 ( .A(n20424), .B(n20425), .Z(n17585) );
  XOR U18369 ( .A(n17581), .B(n17582), .Z(n17584) );
  AND U18370 ( .A(n20426), .B(n20427), .Z(n17582) );
  XOR U18371 ( .A(n17578), .B(n17579), .Z(n17581) );
  AND U18372 ( .A(n20428), .B(n20429), .Z(n17579) );
  XOR U18373 ( .A(n17575), .B(n17576), .Z(n17578) );
  AND U18374 ( .A(n20430), .B(n20431), .Z(n17576) );
  XOR U18375 ( .A(n17572), .B(n17573), .Z(n17575) );
  AND U18376 ( .A(n20432), .B(n20433), .Z(n17573) );
  XOR U18377 ( .A(n17569), .B(n17570), .Z(n17572) );
  AND U18378 ( .A(n20434), .B(n20435), .Z(n17570) );
  XOR U18379 ( .A(n17566), .B(n17567), .Z(n17569) );
  AND U18380 ( .A(n20436), .B(n20437), .Z(n17567) );
  XOR U18381 ( .A(n17563), .B(n17564), .Z(n17566) );
  AND U18382 ( .A(n20438), .B(n20439), .Z(n17564) );
  XOR U18383 ( .A(n17560), .B(n17561), .Z(n17563) );
  AND U18384 ( .A(n20440), .B(n20441), .Z(n17561) );
  XOR U18385 ( .A(n17557), .B(n17558), .Z(n17560) );
  AND U18386 ( .A(n20442), .B(n20443), .Z(n17558) );
  XOR U18387 ( .A(n17554), .B(n17555), .Z(n17557) );
  AND U18388 ( .A(n20444), .B(n20445), .Z(n17555) );
  XOR U18389 ( .A(n17551), .B(n17552), .Z(n17554) );
  AND U18390 ( .A(n20446), .B(n20447), .Z(n17552) );
  XOR U18391 ( .A(n17548), .B(n17549), .Z(n17551) );
  AND U18392 ( .A(n20448), .B(n20449), .Z(n17549) );
  XOR U18393 ( .A(n17545), .B(n17546), .Z(n17548) );
  AND U18394 ( .A(n20450), .B(n20451), .Z(n17546) );
  XOR U18395 ( .A(n17542), .B(n17543), .Z(n17545) );
  AND U18396 ( .A(n20452), .B(n20453), .Z(n17543) );
  XOR U18397 ( .A(n17539), .B(n17540), .Z(n17542) );
  AND U18398 ( .A(n20454), .B(n20455), .Z(n17540) );
  XOR U18399 ( .A(n17536), .B(n17537), .Z(n17539) );
  AND U18400 ( .A(n20456), .B(n20457), .Z(n17537) );
  XOR U18401 ( .A(n17533), .B(n17534), .Z(n17536) );
  AND U18402 ( .A(n20458), .B(n20459), .Z(n17534) );
  XOR U18403 ( .A(n17530), .B(n17531), .Z(n17533) );
  AND U18404 ( .A(n20460), .B(n20461), .Z(n17531) );
  XOR U18405 ( .A(n17527), .B(n17528), .Z(n17530) );
  AND U18406 ( .A(n20462), .B(n20463), .Z(n17528) );
  XOR U18407 ( .A(n17524), .B(n17525), .Z(n17527) );
  AND U18408 ( .A(n20464), .B(n20465), .Z(n17525) );
  XOR U18409 ( .A(n17521), .B(n17522), .Z(n17524) );
  AND U18410 ( .A(n20466), .B(n20467), .Z(n17522) );
  XOR U18411 ( .A(n17518), .B(n17519), .Z(n17521) );
  AND U18412 ( .A(n20468), .B(n20469), .Z(n17519) );
  XOR U18413 ( .A(n17515), .B(n17516), .Z(n17518) );
  AND U18414 ( .A(n20470), .B(n20471), .Z(n17516) );
  XOR U18415 ( .A(n17512), .B(n17513), .Z(n17515) );
  AND U18416 ( .A(n20472), .B(n20473), .Z(n17513) );
  XOR U18417 ( .A(n17509), .B(n17510), .Z(n17512) );
  AND U18418 ( .A(n20474), .B(n20475), .Z(n17510) );
  XOR U18419 ( .A(n17506), .B(n17507), .Z(n17509) );
  AND U18420 ( .A(n20476), .B(n20477), .Z(n17507) );
  XOR U18421 ( .A(n17503), .B(n17504), .Z(n17506) );
  AND U18422 ( .A(n20478), .B(n20479), .Z(n17504) );
  XOR U18423 ( .A(n17500), .B(n17501), .Z(n17503) );
  AND U18424 ( .A(n20480), .B(n20481), .Z(n17501) );
  XOR U18425 ( .A(n17497), .B(n17498), .Z(n17500) );
  AND U18426 ( .A(n20482), .B(n20483), .Z(n17498) );
  XOR U18427 ( .A(n17494), .B(n17495), .Z(n17497) );
  AND U18428 ( .A(n20484), .B(n20485), .Z(n17495) );
  XOR U18429 ( .A(n17491), .B(n17492), .Z(n17494) );
  AND U18430 ( .A(n20486), .B(n20487), .Z(n17492) );
  XOR U18431 ( .A(n17488), .B(n17489), .Z(n17491) );
  AND U18432 ( .A(n20488), .B(n20489), .Z(n17489) );
  XOR U18433 ( .A(n17485), .B(n17486), .Z(n17488) );
  AND U18434 ( .A(n20490), .B(n20491), .Z(n17486) );
  XOR U18435 ( .A(n17482), .B(n17483), .Z(n17485) );
  AND U18436 ( .A(n20492), .B(n20493), .Z(n17483) );
  XOR U18437 ( .A(n17479), .B(n17480), .Z(n17482) );
  AND U18438 ( .A(n20494), .B(n20495), .Z(n17480) );
  XOR U18439 ( .A(n17476), .B(n17477), .Z(n17479) );
  AND U18440 ( .A(n20496), .B(n20497), .Z(n17477) );
  XOR U18441 ( .A(n17473), .B(n17474), .Z(n17476) );
  AND U18442 ( .A(n20498), .B(n20499), .Z(n17474) );
  XOR U18443 ( .A(n17470), .B(n17471), .Z(n17473) );
  AND U18444 ( .A(n20500), .B(n20501), .Z(n17471) );
  XOR U18445 ( .A(n17467), .B(n17468), .Z(n17470) );
  AND U18446 ( .A(n20502), .B(n20503), .Z(n17468) );
  XOR U18447 ( .A(n17464), .B(n17465), .Z(n17467) );
  AND U18448 ( .A(n20504), .B(n20505), .Z(n17465) );
  XOR U18449 ( .A(n17461), .B(n17462), .Z(n17464) );
  AND U18450 ( .A(n20506), .B(n20507), .Z(n17462) );
  XOR U18451 ( .A(n17458), .B(n17459), .Z(n17461) );
  AND U18452 ( .A(n20508), .B(n20509), .Z(n17459) );
  XOR U18453 ( .A(n17455), .B(n17456), .Z(n17458) );
  AND U18454 ( .A(n20510), .B(n20511), .Z(n17456) );
  XOR U18455 ( .A(n17452), .B(n17453), .Z(n17455) );
  AND U18456 ( .A(n20512), .B(n20513), .Z(n17453) );
  XOR U18457 ( .A(n17449), .B(n17450), .Z(n17452) );
  AND U18458 ( .A(n20514), .B(n20515), .Z(n17450) );
  XOR U18459 ( .A(n17446), .B(n17447), .Z(n17449) );
  AND U18460 ( .A(n20516), .B(n20517), .Z(n17447) );
  XOR U18461 ( .A(n17443), .B(n17444), .Z(n17446) );
  AND U18462 ( .A(n20518), .B(n20519), .Z(n17444) );
  XOR U18463 ( .A(n17440), .B(n17441), .Z(n17443) );
  AND U18464 ( .A(n20520), .B(n20521), .Z(n17441) );
  XOR U18465 ( .A(n17437), .B(n17438), .Z(n17440) );
  AND U18466 ( .A(n20522), .B(n20523), .Z(n17438) );
  XOR U18467 ( .A(n17434), .B(n17435), .Z(n17437) );
  AND U18468 ( .A(n20524), .B(n20525), .Z(n17435) );
  XOR U18469 ( .A(n17431), .B(n17432), .Z(n17434) );
  AND U18470 ( .A(n20526), .B(n20527), .Z(n17432) );
  XOR U18471 ( .A(n17428), .B(n17429), .Z(n17431) );
  AND U18472 ( .A(n20528), .B(n20529), .Z(n17429) );
  XOR U18473 ( .A(n17425), .B(n17426), .Z(n17428) );
  AND U18474 ( .A(n20530), .B(n20531), .Z(n17426) );
  XOR U18475 ( .A(n17422), .B(n17423), .Z(n17425) );
  AND U18476 ( .A(n20532), .B(n20533), .Z(n17423) );
  XOR U18477 ( .A(n17419), .B(n17420), .Z(n17422) );
  AND U18478 ( .A(n20534), .B(n20535), .Z(n17420) );
  XOR U18479 ( .A(n17416), .B(n17417), .Z(n17419) );
  AND U18480 ( .A(n20536), .B(n20537), .Z(n17417) );
  XOR U18481 ( .A(n17413), .B(n17414), .Z(n17416) );
  AND U18482 ( .A(n20538), .B(n20539), .Z(n17414) );
  XOR U18483 ( .A(n17410), .B(n17411), .Z(n17413) );
  AND U18484 ( .A(n20540), .B(n20541), .Z(n17411) );
  XOR U18485 ( .A(n17407), .B(n17408), .Z(n17410) );
  AND U18486 ( .A(n20542), .B(n20543), .Z(n17408) );
  XOR U18487 ( .A(n17404), .B(n17405), .Z(n17407) );
  AND U18488 ( .A(n20544), .B(n20545), .Z(n17405) );
  XOR U18489 ( .A(n17401), .B(n17402), .Z(n17404) );
  AND U18490 ( .A(n20546), .B(n20547), .Z(n17402) );
  XOR U18491 ( .A(n17398), .B(n17399), .Z(n17401) );
  AND U18492 ( .A(n20548), .B(n20549), .Z(n17399) );
  XOR U18493 ( .A(n17395), .B(n17396), .Z(n17398) );
  AND U18494 ( .A(n20550), .B(n20551), .Z(n17396) );
  XOR U18495 ( .A(n17392), .B(n17393), .Z(n17395) );
  AND U18496 ( .A(n20552), .B(n20553), .Z(n17393) );
  XOR U18497 ( .A(n17389), .B(n17390), .Z(n17392) );
  AND U18498 ( .A(n20554), .B(n20555), .Z(n17390) );
  XOR U18499 ( .A(n17386), .B(n17387), .Z(n17389) );
  AND U18500 ( .A(n20556), .B(n20557), .Z(n17387) );
  XOR U18501 ( .A(n17383), .B(n17384), .Z(n17386) );
  AND U18502 ( .A(n20558), .B(n20559), .Z(n17384) );
  XOR U18503 ( .A(n17380), .B(n17381), .Z(n17383) );
  AND U18504 ( .A(n20560), .B(n20561), .Z(n17381) );
  XOR U18505 ( .A(n17377), .B(n17378), .Z(n17380) );
  AND U18506 ( .A(n20562), .B(n20563), .Z(n17378) );
  XOR U18507 ( .A(n17374), .B(n17375), .Z(n17377) );
  AND U18508 ( .A(n20564), .B(n20565), .Z(n17375) );
  XOR U18509 ( .A(n17371), .B(n17372), .Z(n17374) );
  AND U18510 ( .A(n20566), .B(n20567), .Z(n17372) );
  XOR U18511 ( .A(n17368), .B(n17369), .Z(n17371) );
  AND U18512 ( .A(n20568), .B(n20569), .Z(n17369) );
  XOR U18513 ( .A(n17365), .B(n17366), .Z(n17368) );
  AND U18514 ( .A(n20570), .B(n20571), .Z(n17366) );
  XOR U18515 ( .A(n17362), .B(n17363), .Z(n17365) );
  AND U18516 ( .A(n20572), .B(n20573), .Z(n17363) );
  XOR U18517 ( .A(n17359), .B(n17360), .Z(n17362) );
  AND U18518 ( .A(n20574), .B(n20575), .Z(n17360) );
  XOR U18519 ( .A(n17356), .B(n17357), .Z(n17359) );
  AND U18520 ( .A(n20576), .B(n20577), .Z(n17357) );
  XOR U18521 ( .A(n17353), .B(n17354), .Z(n17356) );
  AND U18522 ( .A(n20578), .B(n20579), .Z(n17354) );
  XOR U18523 ( .A(n17350), .B(n17351), .Z(n17353) );
  AND U18524 ( .A(n20580), .B(n20581), .Z(n17351) );
  XOR U18525 ( .A(n17347), .B(n17348), .Z(n17350) );
  AND U18526 ( .A(n20582), .B(n20583), .Z(n17348) );
  XOR U18527 ( .A(n17344), .B(n17345), .Z(n17347) );
  AND U18528 ( .A(n20584), .B(n20585), .Z(n17345) );
  XOR U18529 ( .A(n17341), .B(n17342), .Z(n17344) );
  AND U18530 ( .A(n20586), .B(n20587), .Z(n17342) );
  XOR U18531 ( .A(n17338), .B(n17339), .Z(n17341) );
  AND U18532 ( .A(n20588), .B(n20589), .Z(n17339) );
  XOR U18533 ( .A(n17335), .B(n17336), .Z(n17338) );
  AND U18534 ( .A(n20590), .B(n20591), .Z(n17336) );
  XOR U18535 ( .A(n17332), .B(n17333), .Z(n17335) );
  AND U18536 ( .A(n20592), .B(n20593), .Z(n17333) );
  XOR U18537 ( .A(n17329), .B(n17330), .Z(n17332) );
  AND U18538 ( .A(n20594), .B(n20595), .Z(n17330) );
  XOR U18539 ( .A(n17326), .B(n17327), .Z(n17329) );
  AND U18540 ( .A(n20596), .B(n20597), .Z(n17327) );
  XOR U18541 ( .A(n17323), .B(n17324), .Z(n17326) );
  AND U18542 ( .A(n20598), .B(n20599), .Z(n17324) );
  XOR U18543 ( .A(n17320), .B(n17321), .Z(n17323) );
  AND U18544 ( .A(n20600), .B(n20601), .Z(n17321) );
  XOR U18545 ( .A(n17317), .B(n17318), .Z(n17320) );
  AND U18546 ( .A(n20602), .B(n20603), .Z(n17318) );
  XOR U18547 ( .A(n17314), .B(n17315), .Z(n17317) );
  AND U18548 ( .A(n20604), .B(n20605), .Z(n17315) );
  XOR U18549 ( .A(n17311), .B(n17312), .Z(n17314) );
  AND U18550 ( .A(n20606), .B(n20607), .Z(n17312) );
  XOR U18551 ( .A(n17308), .B(n17309), .Z(n17311) );
  AND U18552 ( .A(n20608), .B(n20609), .Z(n17309) );
  XOR U18553 ( .A(n17305), .B(n17306), .Z(n17308) );
  AND U18554 ( .A(n20610), .B(n20611), .Z(n17306) );
  XOR U18555 ( .A(n17302), .B(n17303), .Z(n17305) );
  AND U18556 ( .A(n20612), .B(n20613), .Z(n17303) );
  XOR U18557 ( .A(n17299), .B(n17300), .Z(n17302) );
  AND U18558 ( .A(n20614), .B(n20615), .Z(n17300) );
  XOR U18559 ( .A(n17296), .B(n17297), .Z(n17299) );
  AND U18560 ( .A(n20616), .B(n20617), .Z(n17297) );
  XOR U18561 ( .A(n17293), .B(n17294), .Z(n17296) );
  AND U18562 ( .A(n20618), .B(n20619), .Z(n17294) );
  XOR U18563 ( .A(n17290), .B(n17291), .Z(n17293) );
  AND U18564 ( .A(n20620), .B(n20621), .Z(n17291) );
  XOR U18565 ( .A(n17287), .B(n17288), .Z(n17290) );
  AND U18566 ( .A(n20622), .B(n20623), .Z(n17288) );
  XOR U18567 ( .A(n17284), .B(n17285), .Z(n17287) );
  AND U18568 ( .A(n20624), .B(n20625), .Z(n17285) );
  XNOR U18569 ( .A(n17281), .B(n17282), .Z(n17284) );
  AND U18570 ( .A(n20626), .B(n20627), .Z(n17282) );
  XOR U18571 ( .A(n20628), .B(n17279), .Z(n17281) );
  IV U18572 ( .A(n20629), .Z(n17279) );
  AND U18573 ( .A(n20630), .B(n20631), .Z(n20629) );
  IV U18574 ( .A(n17278), .Z(n20628) );
  XOR U18575 ( .A(n17019), .B(n17275), .Z(n17278) );
  AND U18576 ( .A(n20632), .B(n20633), .Z(n17275) );
  XOR U18577 ( .A(n17021), .B(n17020), .Z(n17019) );
  AND U18578 ( .A(n20634), .B(n20635), .Z(n17020) );
  XOR U18579 ( .A(n17023), .B(n17022), .Z(n17021) );
  AND U18580 ( .A(n20636), .B(n20637), .Z(n17022) );
  XOR U18581 ( .A(n17025), .B(n17024), .Z(n17023) );
  AND U18582 ( .A(n20638), .B(n20639), .Z(n17024) );
  XOR U18583 ( .A(n17027), .B(n17026), .Z(n17025) );
  AND U18584 ( .A(n20640), .B(n20641), .Z(n17026) );
  XOR U18585 ( .A(n17029), .B(n17028), .Z(n17027) );
  AND U18586 ( .A(n20642), .B(n20643), .Z(n17028) );
  XOR U18587 ( .A(n17031), .B(n17030), .Z(n17029) );
  AND U18588 ( .A(n20644), .B(n20645), .Z(n17030) );
  XOR U18589 ( .A(n17033), .B(n17032), .Z(n17031) );
  AND U18590 ( .A(n20646), .B(n20647), .Z(n17032) );
  XOR U18591 ( .A(n17035), .B(n17034), .Z(n17033) );
  AND U18592 ( .A(n20648), .B(n20649), .Z(n17034) );
  XOR U18593 ( .A(n17037), .B(n17036), .Z(n17035) );
  AND U18594 ( .A(n20650), .B(n20651), .Z(n17036) );
  XOR U18595 ( .A(n17039), .B(n17038), .Z(n17037) );
  AND U18596 ( .A(n20652), .B(n20653), .Z(n17038) );
  XOR U18597 ( .A(n17041), .B(n17040), .Z(n17039) );
  AND U18598 ( .A(n20654), .B(n20655), .Z(n17040) );
  XOR U18599 ( .A(n17043), .B(n17042), .Z(n17041) );
  AND U18600 ( .A(n20656), .B(n20657), .Z(n17042) );
  XOR U18601 ( .A(n17045), .B(n17044), .Z(n17043) );
  AND U18602 ( .A(n20658), .B(n20659), .Z(n17044) );
  XOR U18603 ( .A(n17047), .B(n17046), .Z(n17045) );
  AND U18604 ( .A(n20660), .B(n20661), .Z(n17046) );
  XOR U18605 ( .A(n17049), .B(n17048), .Z(n17047) );
  AND U18606 ( .A(n20662), .B(n20663), .Z(n17048) );
  XOR U18607 ( .A(n17051), .B(n17050), .Z(n17049) );
  AND U18608 ( .A(n20664), .B(n20665), .Z(n17050) );
  XOR U18609 ( .A(n17053), .B(n17052), .Z(n17051) );
  AND U18610 ( .A(n20666), .B(n20667), .Z(n17052) );
  XOR U18611 ( .A(n17055), .B(n17054), .Z(n17053) );
  AND U18612 ( .A(n20668), .B(n20669), .Z(n17054) );
  XOR U18613 ( .A(n17057), .B(n17056), .Z(n17055) );
  AND U18614 ( .A(n20670), .B(n20671), .Z(n17056) );
  XOR U18615 ( .A(n17059), .B(n17058), .Z(n17057) );
  AND U18616 ( .A(n20672), .B(n20673), .Z(n17058) );
  XOR U18617 ( .A(n17061), .B(n17060), .Z(n17059) );
  AND U18618 ( .A(n20674), .B(n20675), .Z(n17060) );
  XOR U18619 ( .A(n17063), .B(n17062), .Z(n17061) );
  AND U18620 ( .A(n20676), .B(n20677), .Z(n17062) );
  XOR U18621 ( .A(n17065), .B(n17064), .Z(n17063) );
  AND U18622 ( .A(n20678), .B(n20679), .Z(n17064) );
  XOR U18623 ( .A(n17067), .B(n17066), .Z(n17065) );
  AND U18624 ( .A(n20680), .B(n20681), .Z(n17066) );
  XOR U18625 ( .A(n17069), .B(n17068), .Z(n17067) );
  AND U18626 ( .A(n20682), .B(n20683), .Z(n17068) );
  XOR U18627 ( .A(n17071), .B(n17070), .Z(n17069) );
  AND U18628 ( .A(n20684), .B(n20685), .Z(n17070) );
  XOR U18629 ( .A(n17073), .B(n17072), .Z(n17071) );
  AND U18630 ( .A(n20686), .B(n20687), .Z(n17072) );
  XOR U18631 ( .A(n17075), .B(n17074), .Z(n17073) );
  AND U18632 ( .A(n20688), .B(n20689), .Z(n17074) );
  XOR U18633 ( .A(n17077), .B(n17076), .Z(n17075) );
  AND U18634 ( .A(n20690), .B(n20691), .Z(n17076) );
  XOR U18635 ( .A(n17079), .B(n17078), .Z(n17077) );
  AND U18636 ( .A(n20692), .B(n20693), .Z(n17078) );
  XOR U18637 ( .A(n17081), .B(n17080), .Z(n17079) );
  AND U18638 ( .A(n20694), .B(n20695), .Z(n17080) );
  XOR U18639 ( .A(n17083), .B(n17082), .Z(n17081) );
  AND U18640 ( .A(n20696), .B(n20697), .Z(n17082) );
  XOR U18641 ( .A(n17085), .B(n17084), .Z(n17083) );
  AND U18642 ( .A(n20698), .B(n20699), .Z(n17084) );
  XOR U18643 ( .A(n17087), .B(n17086), .Z(n17085) );
  AND U18644 ( .A(n20700), .B(n20701), .Z(n17086) );
  XOR U18645 ( .A(n17089), .B(n17088), .Z(n17087) );
  AND U18646 ( .A(n20702), .B(n20703), .Z(n17088) );
  XOR U18647 ( .A(n17091), .B(n17090), .Z(n17089) );
  AND U18648 ( .A(n20704), .B(n20705), .Z(n17090) );
  XOR U18649 ( .A(n17093), .B(n17092), .Z(n17091) );
  AND U18650 ( .A(n20706), .B(n20707), .Z(n17092) );
  XOR U18651 ( .A(n17095), .B(n17094), .Z(n17093) );
  AND U18652 ( .A(n20708), .B(n20709), .Z(n17094) );
  XOR U18653 ( .A(n17097), .B(n17096), .Z(n17095) );
  AND U18654 ( .A(n20710), .B(n20711), .Z(n17096) );
  XOR U18655 ( .A(n17099), .B(n17098), .Z(n17097) );
  AND U18656 ( .A(n20712), .B(n20713), .Z(n17098) );
  XOR U18657 ( .A(n17101), .B(n17100), .Z(n17099) );
  AND U18658 ( .A(n20714), .B(n20715), .Z(n17100) );
  XOR U18659 ( .A(n17103), .B(n17102), .Z(n17101) );
  AND U18660 ( .A(n20716), .B(n20717), .Z(n17102) );
  XOR U18661 ( .A(n17105), .B(n17104), .Z(n17103) );
  AND U18662 ( .A(n20718), .B(n20719), .Z(n17104) );
  XOR U18663 ( .A(n17107), .B(n17106), .Z(n17105) );
  AND U18664 ( .A(n20720), .B(n20721), .Z(n17106) );
  XOR U18665 ( .A(n17109), .B(n17108), .Z(n17107) );
  AND U18666 ( .A(n20722), .B(n20723), .Z(n17108) );
  XOR U18667 ( .A(n17111), .B(n17110), .Z(n17109) );
  AND U18668 ( .A(n20724), .B(n20725), .Z(n17110) );
  XOR U18669 ( .A(n17113), .B(n17112), .Z(n17111) );
  AND U18670 ( .A(n20726), .B(n20727), .Z(n17112) );
  XOR U18671 ( .A(n17115), .B(n17114), .Z(n17113) );
  AND U18672 ( .A(n20728), .B(n20729), .Z(n17114) );
  XOR U18673 ( .A(n17117), .B(n17116), .Z(n17115) );
  AND U18674 ( .A(n20730), .B(n20731), .Z(n17116) );
  XOR U18675 ( .A(n17119), .B(n17118), .Z(n17117) );
  AND U18676 ( .A(n20732), .B(n20733), .Z(n17118) );
  XOR U18677 ( .A(n17121), .B(n17120), .Z(n17119) );
  AND U18678 ( .A(n20734), .B(n20735), .Z(n17120) );
  XOR U18679 ( .A(n17123), .B(n17122), .Z(n17121) );
  AND U18680 ( .A(n20736), .B(n20737), .Z(n17122) );
  XOR U18681 ( .A(n17125), .B(n17124), .Z(n17123) );
  AND U18682 ( .A(n20738), .B(n20739), .Z(n17124) );
  XOR U18683 ( .A(n17127), .B(n17126), .Z(n17125) );
  AND U18684 ( .A(n20740), .B(n20741), .Z(n17126) );
  XOR U18685 ( .A(n17129), .B(n17128), .Z(n17127) );
  AND U18686 ( .A(n20742), .B(n20743), .Z(n17128) );
  XOR U18687 ( .A(n17131), .B(n17130), .Z(n17129) );
  AND U18688 ( .A(n20744), .B(n20745), .Z(n17130) );
  XOR U18689 ( .A(n17133), .B(n17132), .Z(n17131) );
  AND U18690 ( .A(n20746), .B(n20747), .Z(n17132) );
  XOR U18691 ( .A(n17135), .B(n17134), .Z(n17133) );
  AND U18692 ( .A(n20748), .B(n20749), .Z(n17134) );
  XOR U18693 ( .A(n17137), .B(n17136), .Z(n17135) );
  AND U18694 ( .A(n20750), .B(n20751), .Z(n17136) );
  XOR U18695 ( .A(n17139), .B(n17138), .Z(n17137) );
  AND U18696 ( .A(n20752), .B(n20753), .Z(n17138) );
  XOR U18697 ( .A(n17141), .B(n17140), .Z(n17139) );
  AND U18698 ( .A(n20754), .B(n20755), .Z(n17140) );
  XOR U18699 ( .A(n17143), .B(n17142), .Z(n17141) );
  AND U18700 ( .A(n20756), .B(n20757), .Z(n17142) );
  XOR U18701 ( .A(n17145), .B(n17144), .Z(n17143) );
  AND U18702 ( .A(n20758), .B(n20759), .Z(n17144) );
  XOR U18703 ( .A(n17147), .B(n17146), .Z(n17145) );
  AND U18704 ( .A(n20760), .B(n20761), .Z(n17146) );
  XOR U18705 ( .A(n17149), .B(n17148), .Z(n17147) );
  AND U18706 ( .A(n20762), .B(n20763), .Z(n17148) );
  XOR U18707 ( .A(n17151), .B(n17150), .Z(n17149) );
  AND U18708 ( .A(n20764), .B(n20765), .Z(n17150) );
  XOR U18709 ( .A(n17153), .B(n17152), .Z(n17151) );
  AND U18710 ( .A(n20766), .B(n20767), .Z(n17152) );
  XOR U18711 ( .A(n17155), .B(n17154), .Z(n17153) );
  AND U18712 ( .A(n20768), .B(n20769), .Z(n17154) );
  XOR U18713 ( .A(n17157), .B(n17156), .Z(n17155) );
  AND U18714 ( .A(n20770), .B(n20771), .Z(n17156) );
  XOR U18715 ( .A(n17159), .B(n17158), .Z(n17157) );
  AND U18716 ( .A(n20772), .B(n20773), .Z(n17158) );
  XOR U18717 ( .A(n17161), .B(n17160), .Z(n17159) );
  AND U18718 ( .A(n20774), .B(n20775), .Z(n17160) );
  XOR U18719 ( .A(n17163), .B(n17162), .Z(n17161) );
  AND U18720 ( .A(n20776), .B(n20777), .Z(n17162) );
  XOR U18721 ( .A(n17165), .B(n17164), .Z(n17163) );
  AND U18722 ( .A(n20778), .B(n20779), .Z(n17164) );
  XOR U18723 ( .A(n17167), .B(n17166), .Z(n17165) );
  AND U18724 ( .A(n20780), .B(n20781), .Z(n17166) );
  XOR U18725 ( .A(n17169), .B(n17168), .Z(n17167) );
  AND U18726 ( .A(n20782), .B(n20783), .Z(n17168) );
  XOR U18727 ( .A(n17171), .B(n17170), .Z(n17169) );
  AND U18728 ( .A(n20784), .B(n20785), .Z(n17170) );
  XOR U18729 ( .A(n17173), .B(n17172), .Z(n17171) );
  AND U18730 ( .A(n20786), .B(n20787), .Z(n17172) );
  XOR U18731 ( .A(n17175), .B(n17174), .Z(n17173) );
  AND U18732 ( .A(n20788), .B(n20789), .Z(n17174) );
  XOR U18733 ( .A(n17177), .B(n17176), .Z(n17175) );
  AND U18734 ( .A(n20790), .B(n20791), .Z(n17176) );
  XOR U18735 ( .A(n17179), .B(n17178), .Z(n17177) );
  AND U18736 ( .A(n20792), .B(n20793), .Z(n17178) );
  XOR U18737 ( .A(n17181), .B(n17180), .Z(n17179) );
  AND U18738 ( .A(n20794), .B(n20795), .Z(n17180) );
  XOR U18739 ( .A(n17183), .B(n17182), .Z(n17181) );
  AND U18740 ( .A(n20796), .B(n20797), .Z(n17182) );
  XOR U18741 ( .A(n17185), .B(n17184), .Z(n17183) );
  AND U18742 ( .A(n20798), .B(n20799), .Z(n17184) );
  XOR U18743 ( .A(n17187), .B(n17186), .Z(n17185) );
  AND U18744 ( .A(n20800), .B(n20801), .Z(n17186) );
  XOR U18745 ( .A(n17189), .B(n17188), .Z(n17187) );
  AND U18746 ( .A(n20802), .B(n20803), .Z(n17188) );
  XOR U18747 ( .A(n17191), .B(n17190), .Z(n17189) );
  AND U18748 ( .A(n20804), .B(n20805), .Z(n17190) );
  XOR U18749 ( .A(n17193), .B(n17192), .Z(n17191) );
  AND U18750 ( .A(n20806), .B(n20807), .Z(n17192) );
  XOR U18751 ( .A(n17195), .B(n17194), .Z(n17193) );
  AND U18752 ( .A(n20808), .B(n20809), .Z(n17194) );
  XOR U18753 ( .A(n17197), .B(n17196), .Z(n17195) );
  AND U18754 ( .A(n20810), .B(n20811), .Z(n17196) );
  XOR U18755 ( .A(n17199), .B(n17198), .Z(n17197) );
  AND U18756 ( .A(n20812), .B(n20813), .Z(n17198) );
  XOR U18757 ( .A(n17201), .B(n17200), .Z(n17199) );
  AND U18758 ( .A(n20814), .B(n20815), .Z(n17200) );
  XOR U18759 ( .A(n17203), .B(n17202), .Z(n17201) );
  AND U18760 ( .A(n20816), .B(n20817), .Z(n17202) );
  XOR U18761 ( .A(n17205), .B(n17204), .Z(n17203) );
  AND U18762 ( .A(n20818), .B(n20819), .Z(n17204) );
  XOR U18763 ( .A(n17207), .B(n17206), .Z(n17205) );
  AND U18764 ( .A(n20820), .B(n20821), .Z(n17206) );
  XOR U18765 ( .A(n17209), .B(n17208), .Z(n17207) );
  AND U18766 ( .A(n20822), .B(n20823), .Z(n17208) );
  XOR U18767 ( .A(n17211), .B(n17210), .Z(n17209) );
  AND U18768 ( .A(n20824), .B(n20825), .Z(n17210) );
  XOR U18769 ( .A(n17213), .B(n17212), .Z(n17211) );
  AND U18770 ( .A(n20826), .B(n20827), .Z(n17212) );
  XOR U18771 ( .A(n17215), .B(n17214), .Z(n17213) );
  AND U18772 ( .A(n20828), .B(n20829), .Z(n17214) );
  XOR U18773 ( .A(n17217), .B(n17216), .Z(n17215) );
  AND U18774 ( .A(n20830), .B(n20831), .Z(n17216) );
  XOR U18775 ( .A(n17219), .B(n17218), .Z(n17217) );
  AND U18776 ( .A(n20832), .B(n20833), .Z(n17218) );
  XOR U18777 ( .A(n17221), .B(n17220), .Z(n17219) );
  AND U18778 ( .A(n20834), .B(n20835), .Z(n17220) );
  XOR U18779 ( .A(n17223), .B(n17222), .Z(n17221) );
  AND U18780 ( .A(n20836), .B(n20837), .Z(n17222) );
  XOR U18781 ( .A(n17225), .B(n17224), .Z(n17223) );
  AND U18782 ( .A(n20838), .B(n20839), .Z(n17224) );
  XOR U18783 ( .A(n17227), .B(n17226), .Z(n17225) );
  AND U18784 ( .A(n20840), .B(n20841), .Z(n17226) );
  XOR U18785 ( .A(n17229), .B(n17228), .Z(n17227) );
  AND U18786 ( .A(n20842), .B(n20843), .Z(n17228) );
  XOR U18787 ( .A(n17231), .B(n17230), .Z(n17229) );
  AND U18788 ( .A(n20844), .B(n20845), .Z(n17230) );
  XOR U18789 ( .A(n17233), .B(n17232), .Z(n17231) );
  AND U18790 ( .A(n20846), .B(n20847), .Z(n17232) );
  XOR U18791 ( .A(n17235), .B(n17234), .Z(n17233) );
  AND U18792 ( .A(n20848), .B(n20849), .Z(n17234) );
  XOR U18793 ( .A(n17237), .B(n17236), .Z(n17235) );
  AND U18794 ( .A(n20850), .B(n20851), .Z(n17236) );
  XOR U18795 ( .A(n17239), .B(n17238), .Z(n17237) );
  AND U18796 ( .A(n20852), .B(n20853), .Z(n17238) );
  XOR U18797 ( .A(n17241), .B(n17240), .Z(n17239) );
  AND U18798 ( .A(n20854), .B(n20855), .Z(n17240) );
  XOR U18799 ( .A(n17243), .B(n17242), .Z(n17241) );
  AND U18800 ( .A(n20856), .B(n20857), .Z(n17242) );
  XOR U18801 ( .A(n17271), .B(n17244), .Z(n17243) );
  AND U18802 ( .A(n20858), .B(n20859), .Z(n17244) );
  XOR U18803 ( .A(n17273), .B(n17272), .Z(n17271) );
  AND U18804 ( .A(n20860), .B(n20861), .Z(n17272) );
  XOR U18805 ( .A(n17252), .B(n17274), .Z(n17273) );
  AND U18806 ( .A(n20862), .B(n20863), .Z(n17274) );
  XOR U18807 ( .A(n17248), .B(n17253), .Z(n17252) );
  AND U18808 ( .A(n20864), .B(n20865), .Z(n17253) );
  XOR U18809 ( .A(n17250), .B(n17249), .Z(n17248) );
  AND U18810 ( .A(n20866), .B(n20867), .Z(n17249) );
  XNOR U18811 ( .A(n17260), .B(n17251), .Z(n17250) );
  AND U18812 ( .A(n20868), .B(n20869), .Z(n17251) );
  XOR U18813 ( .A(n17270), .B(n17259), .Z(n17260) );
  AND U18814 ( .A(n20870), .B(n20871), .Z(n17259) );
  XNOR U18815 ( .A(n20872), .B(n17265), .Z(n17270) );
  XOR U18816 ( .A(n17266), .B(n20873), .Z(n17265) );
  AND U18817 ( .A(n20874), .B(n20875), .Z(n20873) );
  XOR U18818 ( .A(n20876), .B(n20877), .Z(n17266) );
  NOR U18819 ( .A(n20878), .B(n20879), .Z(n20877) );
  AND U18820 ( .A(n20880), .B(n20881), .Z(n20879) );
  AND U18821 ( .A(n20882), .B(n20883), .Z(n20878) );
  XNOR U18822 ( .A(n20880), .B(n20881), .Z(n20876) );
  XNOR U18823 ( .A(n17257), .B(n17269), .Z(n20872) );
  AND U18824 ( .A(n20884), .B(n20885), .Z(n17269) );
  AND U18825 ( .A(n20886), .B(n20887), .Z(n17257) );
  XNOR U18826 ( .A(n19854), .B(n130), .Z(n19856) );
  XOR U18827 ( .A(n19851), .B(n19852), .Z(n130) );
  AND U18828 ( .A(n20888), .B(n20889), .Z(n19852) );
  XOR U18829 ( .A(n19848), .B(n19849), .Z(n19851) );
  AND U18830 ( .A(n20890), .B(n20891), .Z(n19849) );
  XOR U18831 ( .A(n19845), .B(n19846), .Z(n19848) );
  AND U18832 ( .A(n20892), .B(n20893), .Z(n19846) );
  XOR U18833 ( .A(n19842), .B(n19843), .Z(n19845) );
  AND U18834 ( .A(n20894), .B(n20895), .Z(n19843) );
  XOR U18835 ( .A(n19839), .B(n19840), .Z(n19842) );
  AND U18836 ( .A(n20896), .B(n20897), .Z(n19840) );
  XOR U18837 ( .A(n19836), .B(n19837), .Z(n19839) );
  AND U18838 ( .A(n20898), .B(n20899), .Z(n19837) );
  XOR U18839 ( .A(n19833), .B(n19834), .Z(n19836) );
  AND U18840 ( .A(n20900), .B(n20901), .Z(n19834) );
  XOR U18841 ( .A(n19830), .B(n19831), .Z(n19833) );
  AND U18842 ( .A(n20902), .B(n20903), .Z(n19831) );
  XOR U18843 ( .A(n19827), .B(n19828), .Z(n19830) );
  AND U18844 ( .A(n20904), .B(n20905), .Z(n19828) );
  XOR U18845 ( .A(n19824), .B(n19825), .Z(n19827) );
  AND U18846 ( .A(n20906), .B(n20907), .Z(n19825) );
  XOR U18847 ( .A(n19821), .B(n19822), .Z(n19824) );
  AND U18848 ( .A(n20908), .B(n20909), .Z(n19822) );
  XOR U18849 ( .A(n19818), .B(n19819), .Z(n19821) );
  AND U18850 ( .A(n20910), .B(n20911), .Z(n19819) );
  XOR U18851 ( .A(n19815), .B(n19816), .Z(n19818) );
  AND U18852 ( .A(n20912), .B(n20913), .Z(n19816) );
  XOR U18853 ( .A(n19812), .B(n19813), .Z(n19815) );
  AND U18854 ( .A(n20914), .B(n20915), .Z(n19813) );
  XOR U18855 ( .A(n19809), .B(n19810), .Z(n19812) );
  AND U18856 ( .A(n20916), .B(n20917), .Z(n19810) );
  XOR U18857 ( .A(n19806), .B(n19807), .Z(n19809) );
  AND U18858 ( .A(n20918), .B(n20919), .Z(n19807) );
  XOR U18859 ( .A(n19803), .B(n19804), .Z(n19806) );
  AND U18860 ( .A(n20920), .B(n20921), .Z(n19804) );
  XOR U18861 ( .A(n19800), .B(n19801), .Z(n19803) );
  AND U18862 ( .A(n20922), .B(n20923), .Z(n19801) );
  XOR U18863 ( .A(n19797), .B(n19798), .Z(n19800) );
  AND U18864 ( .A(n20924), .B(n20925), .Z(n19798) );
  XOR U18865 ( .A(n19794), .B(n19795), .Z(n19797) );
  AND U18866 ( .A(n20926), .B(n20927), .Z(n19795) );
  XOR U18867 ( .A(n19791), .B(n19792), .Z(n19794) );
  AND U18868 ( .A(n20928), .B(n20929), .Z(n19792) );
  XOR U18869 ( .A(n19788), .B(n19789), .Z(n19791) );
  AND U18870 ( .A(n20930), .B(n20931), .Z(n19789) );
  XOR U18871 ( .A(n19785), .B(n19786), .Z(n19788) );
  AND U18872 ( .A(n20932), .B(n20933), .Z(n19786) );
  XOR U18873 ( .A(n19782), .B(n19783), .Z(n19785) );
  AND U18874 ( .A(n20934), .B(n20935), .Z(n19783) );
  XOR U18875 ( .A(n19779), .B(n19780), .Z(n19782) );
  AND U18876 ( .A(n20936), .B(n20937), .Z(n19780) );
  XOR U18877 ( .A(n19776), .B(n19777), .Z(n19779) );
  AND U18878 ( .A(n20938), .B(n20939), .Z(n19777) );
  XOR U18879 ( .A(n19773), .B(n19774), .Z(n19776) );
  AND U18880 ( .A(n20940), .B(n20941), .Z(n19774) );
  XOR U18881 ( .A(n19770), .B(n19771), .Z(n19773) );
  AND U18882 ( .A(n20942), .B(n20943), .Z(n19771) );
  XOR U18883 ( .A(n19767), .B(n19768), .Z(n19770) );
  AND U18884 ( .A(n20944), .B(n20945), .Z(n19768) );
  XOR U18885 ( .A(n19764), .B(n19765), .Z(n19767) );
  AND U18886 ( .A(n20946), .B(n20947), .Z(n19765) );
  XOR U18887 ( .A(n19761), .B(n19762), .Z(n19764) );
  AND U18888 ( .A(n20948), .B(n20949), .Z(n19762) );
  XOR U18889 ( .A(n19758), .B(n19759), .Z(n19761) );
  AND U18890 ( .A(n20950), .B(n20951), .Z(n19759) );
  XOR U18891 ( .A(n19755), .B(n19756), .Z(n19758) );
  AND U18892 ( .A(n20952), .B(n20953), .Z(n19756) );
  XOR U18893 ( .A(n19752), .B(n19753), .Z(n19755) );
  AND U18894 ( .A(n20954), .B(n20955), .Z(n19753) );
  XOR U18895 ( .A(n19749), .B(n19750), .Z(n19752) );
  AND U18896 ( .A(n20956), .B(n20957), .Z(n19750) );
  XOR U18897 ( .A(n19746), .B(n19747), .Z(n19749) );
  AND U18898 ( .A(n20958), .B(n20959), .Z(n19747) );
  XOR U18899 ( .A(n19743), .B(n19744), .Z(n19746) );
  AND U18900 ( .A(n20960), .B(n20961), .Z(n19744) );
  XOR U18901 ( .A(n19740), .B(n19741), .Z(n19743) );
  AND U18902 ( .A(n20962), .B(n20963), .Z(n19741) );
  XOR U18903 ( .A(n19737), .B(n19738), .Z(n19740) );
  AND U18904 ( .A(n20964), .B(n20965), .Z(n19738) );
  XOR U18905 ( .A(n19734), .B(n19735), .Z(n19737) );
  AND U18906 ( .A(n20966), .B(n20967), .Z(n19735) );
  XOR U18907 ( .A(n19731), .B(n19732), .Z(n19734) );
  AND U18908 ( .A(n20968), .B(n20969), .Z(n19732) );
  XOR U18909 ( .A(n19728), .B(n19729), .Z(n19731) );
  AND U18910 ( .A(n20970), .B(n20971), .Z(n19729) );
  XOR U18911 ( .A(n19725), .B(n19726), .Z(n19728) );
  AND U18912 ( .A(n20972), .B(n20973), .Z(n19726) );
  XOR U18913 ( .A(n19722), .B(n19723), .Z(n19725) );
  AND U18914 ( .A(n20974), .B(n20975), .Z(n19723) );
  XOR U18915 ( .A(n19719), .B(n19720), .Z(n19722) );
  AND U18916 ( .A(n20976), .B(n20977), .Z(n19720) );
  XOR U18917 ( .A(n19716), .B(n19717), .Z(n19719) );
  AND U18918 ( .A(n20978), .B(n20979), .Z(n19717) );
  XOR U18919 ( .A(n19713), .B(n19714), .Z(n19716) );
  AND U18920 ( .A(n20980), .B(n20981), .Z(n19714) );
  XOR U18921 ( .A(n19710), .B(n19711), .Z(n19713) );
  AND U18922 ( .A(n20982), .B(n20983), .Z(n19711) );
  XOR U18923 ( .A(n19707), .B(n19708), .Z(n19710) );
  AND U18924 ( .A(n20984), .B(n20985), .Z(n19708) );
  XOR U18925 ( .A(n19704), .B(n19705), .Z(n19707) );
  AND U18926 ( .A(n20986), .B(n20987), .Z(n19705) );
  XOR U18927 ( .A(n19701), .B(n19702), .Z(n19704) );
  AND U18928 ( .A(n20988), .B(n20989), .Z(n19702) );
  XOR U18929 ( .A(n19698), .B(n19699), .Z(n19701) );
  AND U18930 ( .A(n20990), .B(n20991), .Z(n19699) );
  XOR U18931 ( .A(n19695), .B(n19696), .Z(n19698) );
  AND U18932 ( .A(n20992), .B(n20993), .Z(n19696) );
  XOR U18933 ( .A(n19692), .B(n19693), .Z(n19695) );
  AND U18934 ( .A(n20994), .B(n20995), .Z(n19693) );
  XOR U18935 ( .A(n19689), .B(n19690), .Z(n19692) );
  AND U18936 ( .A(n20996), .B(n20997), .Z(n19690) );
  XOR U18937 ( .A(n19686), .B(n19687), .Z(n19689) );
  AND U18938 ( .A(n20998), .B(n20999), .Z(n19687) );
  XOR U18939 ( .A(n19683), .B(n19684), .Z(n19686) );
  AND U18940 ( .A(n21000), .B(n21001), .Z(n19684) );
  XOR U18941 ( .A(n19680), .B(n19681), .Z(n19683) );
  AND U18942 ( .A(n21002), .B(n21003), .Z(n19681) );
  XOR U18943 ( .A(n19677), .B(n19678), .Z(n19680) );
  AND U18944 ( .A(n21004), .B(n21005), .Z(n19678) );
  XOR U18945 ( .A(n19674), .B(n19675), .Z(n19677) );
  AND U18946 ( .A(n21006), .B(n21007), .Z(n19675) );
  XOR U18947 ( .A(n19671), .B(n19672), .Z(n19674) );
  AND U18948 ( .A(n21008), .B(n21009), .Z(n19672) );
  XOR U18949 ( .A(n19668), .B(n19669), .Z(n19671) );
  AND U18950 ( .A(n21010), .B(n21011), .Z(n19669) );
  XOR U18951 ( .A(n19665), .B(n19666), .Z(n19668) );
  AND U18952 ( .A(n21012), .B(n21013), .Z(n19666) );
  XOR U18953 ( .A(n19662), .B(n19663), .Z(n19665) );
  AND U18954 ( .A(n21014), .B(n21015), .Z(n19663) );
  XOR U18955 ( .A(n19659), .B(n19660), .Z(n19662) );
  AND U18956 ( .A(n21016), .B(n21017), .Z(n19660) );
  XOR U18957 ( .A(n19656), .B(n19657), .Z(n19659) );
  AND U18958 ( .A(n21018), .B(n21019), .Z(n19657) );
  XOR U18959 ( .A(n19653), .B(n19654), .Z(n19656) );
  AND U18960 ( .A(n21020), .B(n21021), .Z(n19654) );
  XOR U18961 ( .A(n19650), .B(n19651), .Z(n19653) );
  AND U18962 ( .A(n21022), .B(n21023), .Z(n19651) );
  XOR U18963 ( .A(n19647), .B(n19648), .Z(n19650) );
  AND U18964 ( .A(n21024), .B(n21025), .Z(n19648) );
  XOR U18965 ( .A(n19644), .B(n19645), .Z(n19647) );
  AND U18966 ( .A(n21026), .B(n21027), .Z(n19645) );
  XOR U18967 ( .A(n19641), .B(n19642), .Z(n19644) );
  AND U18968 ( .A(n21028), .B(n21029), .Z(n19642) );
  XOR U18969 ( .A(n19638), .B(n19639), .Z(n19641) );
  AND U18970 ( .A(n21030), .B(n21031), .Z(n19639) );
  XOR U18971 ( .A(n19635), .B(n19636), .Z(n19638) );
  AND U18972 ( .A(n21032), .B(n21033), .Z(n19636) );
  XOR U18973 ( .A(n19632), .B(n19633), .Z(n19635) );
  AND U18974 ( .A(n21034), .B(n21035), .Z(n19633) );
  XOR U18975 ( .A(n19629), .B(n19630), .Z(n19632) );
  AND U18976 ( .A(n21036), .B(n21037), .Z(n19630) );
  XOR U18977 ( .A(n19626), .B(n19627), .Z(n19629) );
  AND U18978 ( .A(n21038), .B(n21039), .Z(n19627) );
  XOR U18979 ( .A(n19623), .B(n19624), .Z(n19626) );
  AND U18980 ( .A(n21040), .B(n21041), .Z(n19624) );
  XOR U18981 ( .A(n19620), .B(n19621), .Z(n19623) );
  AND U18982 ( .A(n21042), .B(n21043), .Z(n19621) );
  XOR U18983 ( .A(n19617), .B(n19618), .Z(n19620) );
  AND U18984 ( .A(n21044), .B(n21045), .Z(n19618) );
  XOR U18985 ( .A(n19614), .B(n19615), .Z(n19617) );
  AND U18986 ( .A(n21046), .B(n21047), .Z(n19615) );
  XOR U18987 ( .A(n19611), .B(n19612), .Z(n19614) );
  AND U18988 ( .A(n21048), .B(n21049), .Z(n19612) );
  XOR U18989 ( .A(n19608), .B(n19609), .Z(n19611) );
  AND U18990 ( .A(n21050), .B(n21051), .Z(n19609) );
  XOR U18991 ( .A(n19605), .B(n19606), .Z(n19608) );
  AND U18992 ( .A(n21052), .B(n21053), .Z(n19606) );
  XOR U18993 ( .A(n19602), .B(n19603), .Z(n19605) );
  AND U18994 ( .A(n21054), .B(n21055), .Z(n19603) );
  XOR U18995 ( .A(n19599), .B(n19600), .Z(n19602) );
  AND U18996 ( .A(n21056), .B(n21057), .Z(n19600) );
  XOR U18997 ( .A(n19596), .B(n19597), .Z(n19599) );
  AND U18998 ( .A(n21058), .B(n21059), .Z(n19597) );
  XOR U18999 ( .A(n19593), .B(n19594), .Z(n19596) );
  AND U19000 ( .A(n21060), .B(n21061), .Z(n19594) );
  XOR U19001 ( .A(n19590), .B(n19591), .Z(n19593) );
  AND U19002 ( .A(n21062), .B(n21063), .Z(n19591) );
  XOR U19003 ( .A(n19587), .B(n19588), .Z(n19590) );
  AND U19004 ( .A(n21064), .B(n21065), .Z(n19588) );
  XOR U19005 ( .A(n19584), .B(n19585), .Z(n19587) );
  AND U19006 ( .A(n21066), .B(n21067), .Z(n19585) );
  XOR U19007 ( .A(n19581), .B(n19582), .Z(n19584) );
  AND U19008 ( .A(n21068), .B(n21069), .Z(n19582) );
  XOR U19009 ( .A(n19578), .B(n19579), .Z(n19581) );
  AND U19010 ( .A(n21070), .B(n21071), .Z(n19579) );
  XOR U19011 ( .A(n19575), .B(n19576), .Z(n19578) );
  AND U19012 ( .A(n21072), .B(n21073), .Z(n19576) );
  XOR U19013 ( .A(n19572), .B(n19573), .Z(n19575) );
  AND U19014 ( .A(n21074), .B(n21075), .Z(n19573) );
  XOR U19015 ( .A(n19569), .B(n19570), .Z(n19572) );
  AND U19016 ( .A(n21076), .B(n21077), .Z(n19570) );
  XOR U19017 ( .A(n19566), .B(n19567), .Z(n19569) );
  AND U19018 ( .A(n21078), .B(n21079), .Z(n19567) );
  XOR U19019 ( .A(n19563), .B(n19564), .Z(n19566) );
  AND U19020 ( .A(n21080), .B(n21081), .Z(n19564) );
  XOR U19021 ( .A(n19560), .B(n19561), .Z(n19563) );
  AND U19022 ( .A(n21082), .B(n21083), .Z(n19561) );
  XOR U19023 ( .A(n19557), .B(n19558), .Z(n19560) );
  AND U19024 ( .A(n21084), .B(n21085), .Z(n19558) );
  XOR U19025 ( .A(n19554), .B(n19555), .Z(n19557) );
  AND U19026 ( .A(n21086), .B(n21087), .Z(n19555) );
  XOR U19027 ( .A(n19551), .B(n19552), .Z(n19554) );
  AND U19028 ( .A(n21088), .B(n21089), .Z(n19552) );
  XOR U19029 ( .A(n19548), .B(n19549), .Z(n19551) );
  AND U19030 ( .A(n21090), .B(n21091), .Z(n19549) );
  XOR U19031 ( .A(n19545), .B(n19546), .Z(n19548) );
  AND U19032 ( .A(n21092), .B(n21093), .Z(n19546) );
  XOR U19033 ( .A(n19542), .B(n19543), .Z(n19545) );
  AND U19034 ( .A(n21094), .B(n21095), .Z(n19543) );
  XOR U19035 ( .A(n19539), .B(n19540), .Z(n19542) );
  AND U19036 ( .A(n21096), .B(n21097), .Z(n19540) );
  XOR U19037 ( .A(n19536), .B(n19537), .Z(n19539) );
  AND U19038 ( .A(n21098), .B(n21099), .Z(n19537) );
  XOR U19039 ( .A(n19533), .B(n19534), .Z(n19536) );
  AND U19040 ( .A(n21100), .B(n21101), .Z(n19534) );
  XOR U19041 ( .A(n19530), .B(n19531), .Z(n19533) );
  AND U19042 ( .A(n21102), .B(n21103), .Z(n19531) );
  XOR U19043 ( .A(n19527), .B(n19528), .Z(n19530) );
  AND U19044 ( .A(n21104), .B(n21105), .Z(n19528) );
  XOR U19045 ( .A(n19524), .B(n19525), .Z(n19527) );
  AND U19046 ( .A(n21106), .B(n21107), .Z(n19525) );
  XOR U19047 ( .A(n19521), .B(n19522), .Z(n19524) );
  AND U19048 ( .A(n21108), .B(n21109), .Z(n19522) );
  XOR U19049 ( .A(n19518), .B(n19519), .Z(n19521) );
  AND U19050 ( .A(n21110), .B(n21111), .Z(n19519) );
  XOR U19051 ( .A(n19515), .B(n19516), .Z(n19518) );
  AND U19052 ( .A(n21112), .B(n21113), .Z(n19516) );
  XOR U19053 ( .A(n19512), .B(n19513), .Z(n19515) );
  AND U19054 ( .A(n21114), .B(n21115), .Z(n19513) );
  XOR U19055 ( .A(n19509), .B(n19510), .Z(n19512) );
  AND U19056 ( .A(n21116), .B(n21117), .Z(n19510) );
  XOR U19057 ( .A(n19506), .B(n19507), .Z(n19509) );
  AND U19058 ( .A(n21118), .B(n21119), .Z(n19507) );
  XOR U19059 ( .A(n19503), .B(n19504), .Z(n19506) );
  AND U19060 ( .A(n21120), .B(n21121), .Z(n19504) );
  XOR U19061 ( .A(n19500), .B(n19501), .Z(n19503) );
  AND U19062 ( .A(n21122), .B(n21123), .Z(n19501) );
  XOR U19063 ( .A(n19497), .B(n19498), .Z(n19500) );
  AND U19064 ( .A(n21124), .B(n21125), .Z(n19498) );
  XOR U19065 ( .A(n19494), .B(n19495), .Z(n19497) );
  AND U19066 ( .A(n21126), .B(n21127), .Z(n19495) );
  XOR U19067 ( .A(n19491), .B(n19492), .Z(n19494) );
  AND U19068 ( .A(n21128), .B(n21129), .Z(n19492) );
  XOR U19069 ( .A(n19488), .B(n19489), .Z(n19491) );
  AND U19070 ( .A(n21130), .B(n21131), .Z(n19489) );
  XOR U19071 ( .A(n19485), .B(n19486), .Z(n19488) );
  AND U19072 ( .A(n21132), .B(n21133), .Z(n19486) );
  XOR U19073 ( .A(n19482), .B(n19483), .Z(n19485) );
  AND U19074 ( .A(n21134), .B(n21135), .Z(n19483) );
  XOR U19075 ( .A(n19479), .B(n19480), .Z(n19482) );
  AND U19076 ( .A(n21136), .B(n21137), .Z(n19480) );
  XOR U19077 ( .A(n19476), .B(n19477), .Z(n19479) );
  AND U19078 ( .A(n21138), .B(n21139), .Z(n19477) );
  XOR U19079 ( .A(n19473), .B(n19474), .Z(n19476) );
  AND U19080 ( .A(n21140), .B(n21141), .Z(n19474) );
  XOR U19081 ( .A(n19470), .B(n19471), .Z(n19473) );
  AND U19082 ( .A(n21142), .B(n21143), .Z(n19471) );
  XOR U19083 ( .A(n19467), .B(n19468), .Z(n19470) );
  AND U19084 ( .A(n21144), .B(n21145), .Z(n19468) );
  XOR U19085 ( .A(n19464), .B(n19465), .Z(n19467) );
  AND U19086 ( .A(n21146), .B(n21147), .Z(n19465) );
  XOR U19087 ( .A(n19461), .B(n19462), .Z(n19464) );
  AND U19088 ( .A(n21148), .B(n21149), .Z(n19462) );
  XOR U19089 ( .A(n19458), .B(n19459), .Z(n19461) );
  AND U19090 ( .A(n21150), .B(n21151), .Z(n19459) );
  XOR U19091 ( .A(n19455), .B(n19456), .Z(n19458) );
  AND U19092 ( .A(n21152), .B(n21153), .Z(n19456) );
  XOR U19093 ( .A(n19452), .B(n19453), .Z(n19455) );
  AND U19094 ( .A(n21154), .B(n21155), .Z(n19453) );
  XOR U19095 ( .A(n19449), .B(n19450), .Z(n19452) );
  AND U19096 ( .A(n21156), .B(n21157), .Z(n19450) );
  XOR U19097 ( .A(n19446), .B(n19447), .Z(n19449) );
  AND U19098 ( .A(n21158), .B(n21159), .Z(n19447) );
  XOR U19099 ( .A(n19443), .B(n19444), .Z(n19446) );
  AND U19100 ( .A(n21160), .B(n21161), .Z(n19444) );
  XOR U19101 ( .A(n19440), .B(n19441), .Z(n19443) );
  AND U19102 ( .A(n21162), .B(n21163), .Z(n19441) );
  XOR U19103 ( .A(n19437), .B(n19438), .Z(n19440) );
  AND U19104 ( .A(n21164), .B(n21165), .Z(n19438) );
  XOR U19105 ( .A(n19434), .B(n19435), .Z(n19437) );
  AND U19106 ( .A(n21166), .B(n21167), .Z(n19435) );
  XOR U19107 ( .A(n19431), .B(n19432), .Z(n19434) );
  AND U19108 ( .A(n21168), .B(n21169), .Z(n19432) );
  XOR U19109 ( .A(n19428), .B(n19429), .Z(n19431) );
  AND U19110 ( .A(n21170), .B(n21171), .Z(n19429) );
  XOR U19111 ( .A(n19425), .B(n19426), .Z(n19428) );
  AND U19112 ( .A(n21172), .B(n21173), .Z(n19426) );
  XOR U19113 ( .A(n19422), .B(n19423), .Z(n19425) );
  AND U19114 ( .A(n21174), .B(n21175), .Z(n19423) );
  XOR U19115 ( .A(n19419), .B(n19420), .Z(n19422) );
  AND U19116 ( .A(n21176), .B(n21177), .Z(n19420) );
  XOR U19117 ( .A(n19416), .B(n19417), .Z(n19419) );
  AND U19118 ( .A(n21178), .B(n21179), .Z(n19417) );
  XOR U19119 ( .A(n19413), .B(n19414), .Z(n19416) );
  AND U19120 ( .A(n21180), .B(n21181), .Z(n19414) );
  XOR U19121 ( .A(n19410), .B(n19411), .Z(n19413) );
  AND U19122 ( .A(n21182), .B(n21183), .Z(n19411) );
  XOR U19123 ( .A(n19407), .B(n19408), .Z(n19410) );
  AND U19124 ( .A(n21184), .B(n21185), .Z(n19408) );
  XOR U19125 ( .A(n19404), .B(n19405), .Z(n19407) );
  AND U19126 ( .A(n21186), .B(n21187), .Z(n19405) );
  XOR U19127 ( .A(n19401), .B(n19402), .Z(n19404) );
  AND U19128 ( .A(n21188), .B(n21189), .Z(n19402) );
  XOR U19129 ( .A(n19398), .B(n19399), .Z(n19401) );
  AND U19130 ( .A(n21190), .B(n21191), .Z(n19399) );
  XOR U19131 ( .A(n19395), .B(n19396), .Z(n19398) );
  AND U19132 ( .A(n21192), .B(n21193), .Z(n19396) );
  XOR U19133 ( .A(n19392), .B(n19393), .Z(n19395) );
  AND U19134 ( .A(n21194), .B(n21195), .Z(n19393) );
  XOR U19135 ( .A(n19389), .B(n19390), .Z(n19392) );
  AND U19136 ( .A(n21196), .B(n21197), .Z(n19390) );
  XOR U19137 ( .A(n19386), .B(n19387), .Z(n19389) );
  AND U19138 ( .A(n21198), .B(n21199), .Z(n19387) );
  XOR U19139 ( .A(n19383), .B(n19384), .Z(n19386) );
  AND U19140 ( .A(n21200), .B(n21201), .Z(n19384) );
  XOR U19141 ( .A(n19380), .B(n19381), .Z(n19383) );
  AND U19142 ( .A(n21202), .B(n21203), .Z(n19381) );
  XOR U19143 ( .A(n19377), .B(n19378), .Z(n19380) );
  AND U19144 ( .A(n21204), .B(n21205), .Z(n19378) );
  XOR U19145 ( .A(n19374), .B(n19375), .Z(n19377) );
  AND U19146 ( .A(n21206), .B(n21207), .Z(n19375) );
  XOR U19147 ( .A(n19371), .B(n19372), .Z(n19374) );
  AND U19148 ( .A(n21208), .B(n21209), .Z(n19372) );
  XOR U19149 ( .A(n19368), .B(n19369), .Z(n19371) );
  AND U19150 ( .A(n21210), .B(n21211), .Z(n19369) );
  XOR U19151 ( .A(n19365), .B(n19366), .Z(n19368) );
  AND U19152 ( .A(n21212), .B(n21213), .Z(n19366) );
  XOR U19153 ( .A(n19362), .B(n19363), .Z(n19365) );
  AND U19154 ( .A(n21214), .B(n21215), .Z(n19363) );
  XOR U19155 ( .A(n19359), .B(n19360), .Z(n19362) );
  AND U19156 ( .A(n21216), .B(n21217), .Z(n19360) );
  XOR U19157 ( .A(n19356), .B(n19357), .Z(n19359) );
  AND U19158 ( .A(n21218), .B(n21219), .Z(n19357) );
  XOR U19159 ( .A(n19353), .B(n19354), .Z(n19356) );
  AND U19160 ( .A(n21220), .B(n21221), .Z(n19354) );
  XOR U19161 ( .A(n19350), .B(n19351), .Z(n19353) );
  AND U19162 ( .A(n21222), .B(n21223), .Z(n19351) );
  XOR U19163 ( .A(n19347), .B(n19348), .Z(n19350) );
  AND U19164 ( .A(n21224), .B(n21225), .Z(n19348) );
  XOR U19165 ( .A(n19344), .B(n19345), .Z(n19347) );
  AND U19166 ( .A(n21226), .B(n21227), .Z(n19345) );
  XOR U19167 ( .A(n19341), .B(n19342), .Z(n19344) );
  AND U19168 ( .A(n21228), .B(n21229), .Z(n19342) );
  XOR U19169 ( .A(n19338), .B(n19339), .Z(n19341) );
  AND U19170 ( .A(n21230), .B(n21231), .Z(n19339) );
  XOR U19171 ( .A(n19335), .B(n19336), .Z(n19338) );
  AND U19172 ( .A(n21232), .B(n21233), .Z(n19336) );
  XOR U19173 ( .A(n19332), .B(n19333), .Z(n19335) );
  AND U19174 ( .A(n21234), .B(n21235), .Z(n19333) );
  XOR U19175 ( .A(n19329), .B(n19330), .Z(n19332) );
  AND U19176 ( .A(n21236), .B(n21237), .Z(n19330) );
  XOR U19177 ( .A(n19326), .B(n19327), .Z(n19329) );
  AND U19178 ( .A(n21238), .B(n21239), .Z(n19327) );
  XOR U19179 ( .A(n19323), .B(n19324), .Z(n19326) );
  AND U19180 ( .A(n21240), .B(n21241), .Z(n19324) );
  XOR U19181 ( .A(n19320), .B(n19321), .Z(n19323) );
  AND U19182 ( .A(n21242), .B(n21243), .Z(n19321) );
  XOR U19183 ( .A(n19317), .B(n19318), .Z(n19320) );
  AND U19184 ( .A(n21244), .B(n21245), .Z(n19318) );
  XOR U19185 ( .A(n19314), .B(n19315), .Z(n19317) );
  AND U19186 ( .A(n21246), .B(n21247), .Z(n19315) );
  XOR U19187 ( .A(n19311), .B(n19312), .Z(n19314) );
  AND U19188 ( .A(n21248), .B(n21249), .Z(n19312) );
  XOR U19189 ( .A(n19308), .B(n19309), .Z(n19311) );
  AND U19190 ( .A(n21250), .B(n21251), .Z(n19309) );
  XOR U19191 ( .A(n19305), .B(n19306), .Z(n19308) );
  AND U19192 ( .A(n21252), .B(n21253), .Z(n19306) );
  XOR U19193 ( .A(n19302), .B(n19303), .Z(n19305) );
  AND U19194 ( .A(n21254), .B(n21255), .Z(n19303) );
  XOR U19195 ( .A(n19299), .B(n19300), .Z(n19302) );
  AND U19196 ( .A(n21256), .B(n21257), .Z(n19300) );
  XOR U19197 ( .A(n19296), .B(n19297), .Z(n19299) );
  AND U19198 ( .A(n21258), .B(n21259), .Z(n19297) );
  XOR U19199 ( .A(n19293), .B(n19294), .Z(n19296) );
  AND U19200 ( .A(n21260), .B(n21261), .Z(n19294) );
  XOR U19201 ( .A(n19290), .B(n19291), .Z(n19293) );
  AND U19202 ( .A(n21262), .B(n21263), .Z(n19291) );
  XOR U19203 ( .A(n19287), .B(n19288), .Z(n19290) );
  AND U19204 ( .A(n21264), .B(n21265), .Z(n19288) );
  XOR U19205 ( .A(n19284), .B(n19285), .Z(n19287) );
  AND U19206 ( .A(n21266), .B(n21267), .Z(n19285) );
  XOR U19207 ( .A(n19281), .B(n19282), .Z(n19284) );
  AND U19208 ( .A(n21268), .B(n21269), .Z(n19282) );
  XOR U19209 ( .A(n19278), .B(n19279), .Z(n19281) );
  AND U19210 ( .A(n21270), .B(n21271), .Z(n19279) );
  XOR U19211 ( .A(n19275), .B(n19276), .Z(n19278) );
  AND U19212 ( .A(n21272), .B(n21273), .Z(n19276) );
  XOR U19213 ( .A(n19272), .B(n19273), .Z(n19275) );
  AND U19214 ( .A(n21274), .B(n21275), .Z(n19273) );
  XOR U19215 ( .A(n19269), .B(n19270), .Z(n19272) );
  AND U19216 ( .A(n21276), .B(n21277), .Z(n19270) );
  XOR U19217 ( .A(n19266), .B(n19267), .Z(n19269) );
  AND U19218 ( .A(n21278), .B(n21279), .Z(n19267) );
  XOR U19219 ( .A(n19263), .B(n19264), .Z(n19266) );
  AND U19220 ( .A(n21280), .B(n21281), .Z(n19264) );
  XOR U19221 ( .A(n19260), .B(n19261), .Z(n19263) );
  AND U19222 ( .A(n21282), .B(n21283), .Z(n19261) );
  XOR U19223 ( .A(n19257), .B(n19258), .Z(n19260) );
  AND U19224 ( .A(n21284), .B(n21285), .Z(n19258) );
  XOR U19225 ( .A(n19254), .B(n19255), .Z(n19257) );
  AND U19226 ( .A(n21286), .B(n21287), .Z(n19255) );
  XOR U19227 ( .A(n19251), .B(n19252), .Z(n19254) );
  AND U19228 ( .A(n21288), .B(n21289), .Z(n19252) );
  XOR U19229 ( .A(n19248), .B(n19249), .Z(n19251) );
  AND U19230 ( .A(n21290), .B(n21291), .Z(n19249) );
  XOR U19231 ( .A(n19245), .B(n19246), .Z(n19248) );
  AND U19232 ( .A(n21292), .B(n21293), .Z(n19246) );
  XOR U19233 ( .A(n19242), .B(n19243), .Z(n19245) );
  AND U19234 ( .A(n21294), .B(n21295), .Z(n19243) );
  XOR U19235 ( .A(n19239), .B(n19240), .Z(n19242) );
  AND U19236 ( .A(n21296), .B(n21297), .Z(n19240) );
  XOR U19237 ( .A(n19236), .B(n19237), .Z(n19239) );
  AND U19238 ( .A(n21298), .B(n21299), .Z(n19237) );
  XOR U19239 ( .A(n19233), .B(n19234), .Z(n19236) );
  AND U19240 ( .A(n21300), .B(n21301), .Z(n19234) );
  XOR U19241 ( .A(n19230), .B(n19231), .Z(n19233) );
  AND U19242 ( .A(n21302), .B(n21303), .Z(n19231) );
  XOR U19243 ( .A(n19227), .B(n19228), .Z(n19230) );
  AND U19244 ( .A(n21304), .B(n21305), .Z(n19228) );
  XOR U19245 ( .A(n19224), .B(n19225), .Z(n19227) );
  AND U19246 ( .A(n21306), .B(n21307), .Z(n19225) );
  XOR U19247 ( .A(n19221), .B(n19222), .Z(n19224) );
  AND U19248 ( .A(n21308), .B(n21309), .Z(n19222) );
  XOR U19249 ( .A(n19218), .B(n19219), .Z(n19221) );
  AND U19250 ( .A(n21310), .B(n21311), .Z(n19219) );
  XOR U19251 ( .A(n19215), .B(n19216), .Z(n19218) );
  AND U19252 ( .A(n21312), .B(n21313), .Z(n19216) );
  XOR U19253 ( .A(n19212), .B(n19213), .Z(n19215) );
  AND U19254 ( .A(n21314), .B(n21315), .Z(n19213) );
  XOR U19255 ( .A(n19209), .B(n19210), .Z(n19212) );
  AND U19256 ( .A(n21316), .B(n21317), .Z(n19210) );
  XOR U19257 ( .A(n19206), .B(n19207), .Z(n19209) );
  AND U19258 ( .A(n21318), .B(n21319), .Z(n19207) );
  XOR U19259 ( .A(n19203), .B(n19204), .Z(n19206) );
  AND U19260 ( .A(n21320), .B(n21321), .Z(n19204) );
  XOR U19261 ( .A(n19200), .B(n19201), .Z(n19203) );
  AND U19262 ( .A(n21322), .B(n21323), .Z(n19201) );
  XOR U19263 ( .A(n19197), .B(n19198), .Z(n19200) );
  AND U19264 ( .A(n21324), .B(n21325), .Z(n19198) );
  XOR U19265 ( .A(n19194), .B(n19195), .Z(n19197) );
  AND U19266 ( .A(n21326), .B(n21327), .Z(n19195) );
  XOR U19267 ( .A(n19191), .B(n19192), .Z(n19194) );
  AND U19268 ( .A(n21328), .B(n21329), .Z(n19192) );
  XOR U19269 ( .A(n19188), .B(n19189), .Z(n19191) );
  AND U19270 ( .A(n21330), .B(n21331), .Z(n19189) );
  XOR U19271 ( .A(n19185), .B(n19186), .Z(n19188) );
  AND U19272 ( .A(n21332), .B(n21333), .Z(n19186) );
  XOR U19273 ( .A(n19182), .B(n19183), .Z(n19185) );
  AND U19274 ( .A(n21334), .B(n21335), .Z(n19183) );
  XOR U19275 ( .A(n19179), .B(n19180), .Z(n19182) );
  AND U19276 ( .A(n21336), .B(n21337), .Z(n19180) );
  XOR U19277 ( .A(n19176), .B(n19177), .Z(n19179) );
  AND U19278 ( .A(n21338), .B(n21339), .Z(n19177) );
  XOR U19279 ( .A(n19173), .B(n19174), .Z(n19176) );
  AND U19280 ( .A(n21340), .B(n21341), .Z(n19174) );
  XOR U19281 ( .A(n19170), .B(n19171), .Z(n19173) );
  AND U19282 ( .A(n21342), .B(n21343), .Z(n19171) );
  XOR U19283 ( .A(n19167), .B(n19168), .Z(n19170) );
  AND U19284 ( .A(n21344), .B(n21345), .Z(n19168) );
  XOR U19285 ( .A(n19164), .B(n19165), .Z(n19167) );
  AND U19286 ( .A(n21346), .B(n21347), .Z(n19165) );
  XOR U19287 ( .A(n19161), .B(n19162), .Z(n19164) );
  AND U19288 ( .A(n21348), .B(n21349), .Z(n19162) );
  XOR U19289 ( .A(n19158), .B(n19159), .Z(n19161) );
  AND U19290 ( .A(n21350), .B(n21351), .Z(n19159) );
  XOR U19291 ( .A(n19155), .B(n19156), .Z(n19158) );
  AND U19292 ( .A(n21352), .B(n21353), .Z(n19156) );
  XOR U19293 ( .A(n19152), .B(n19153), .Z(n19155) );
  AND U19294 ( .A(n21354), .B(n21355), .Z(n19153) );
  XOR U19295 ( .A(n19149), .B(n19150), .Z(n19152) );
  AND U19296 ( .A(n21356), .B(n21357), .Z(n19150) );
  XOR U19297 ( .A(n19146), .B(n19147), .Z(n19149) );
  AND U19298 ( .A(n21358), .B(n21359), .Z(n19147) );
  XOR U19299 ( .A(n19143), .B(n19144), .Z(n19146) );
  AND U19300 ( .A(n21360), .B(n21361), .Z(n19144) );
  XOR U19301 ( .A(n19140), .B(n19141), .Z(n19143) );
  AND U19302 ( .A(n21362), .B(n21363), .Z(n19141) );
  XOR U19303 ( .A(n19137), .B(n19138), .Z(n19140) );
  AND U19304 ( .A(n21364), .B(n21365), .Z(n19138) );
  XOR U19305 ( .A(n19134), .B(n19135), .Z(n19137) );
  AND U19306 ( .A(n21366), .B(n21367), .Z(n19135) );
  XOR U19307 ( .A(n19131), .B(n19132), .Z(n19134) );
  AND U19308 ( .A(n21368), .B(n21369), .Z(n19132) );
  XOR U19309 ( .A(n19128), .B(n19129), .Z(n19131) );
  AND U19310 ( .A(n21370), .B(n21371), .Z(n19129) );
  XOR U19311 ( .A(n19125), .B(n19126), .Z(n19128) );
  AND U19312 ( .A(n21372), .B(n21373), .Z(n19126) );
  XOR U19313 ( .A(n19122), .B(n19123), .Z(n19125) );
  AND U19314 ( .A(n21374), .B(n21375), .Z(n19123) );
  XOR U19315 ( .A(n19119), .B(n19120), .Z(n19122) );
  AND U19316 ( .A(n21376), .B(n21377), .Z(n19120) );
  XOR U19317 ( .A(n19116), .B(n19117), .Z(n19119) );
  AND U19318 ( .A(n21378), .B(n21379), .Z(n19117) );
  XOR U19319 ( .A(n19113), .B(n19114), .Z(n19116) );
  AND U19320 ( .A(n21380), .B(n21381), .Z(n19114) );
  XOR U19321 ( .A(n19110), .B(n19111), .Z(n19113) );
  AND U19322 ( .A(n21382), .B(n21383), .Z(n19111) );
  XOR U19323 ( .A(n19107), .B(n19108), .Z(n19110) );
  AND U19324 ( .A(n21384), .B(n21385), .Z(n19108) );
  XOR U19325 ( .A(n19104), .B(n19105), .Z(n19107) );
  AND U19326 ( .A(n21386), .B(n21387), .Z(n19105) );
  XOR U19327 ( .A(n19101), .B(n19102), .Z(n19104) );
  AND U19328 ( .A(n21388), .B(n21389), .Z(n19102) );
  XOR U19329 ( .A(n19098), .B(n19099), .Z(n19101) );
  AND U19330 ( .A(n21390), .B(n21391), .Z(n19099) );
  XOR U19331 ( .A(n19095), .B(n19096), .Z(n19098) );
  AND U19332 ( .A(n21392), .B(n21393), .Z(n19096) );
  XOR U19333 ( .A(n19092), .B(n19093), .Z(n19095) );
  AND U19334 ( .A(n21394), .B(n21395), .Z(n19093) );
  XOR U19335 ( .A(n19089), .B(n19090), .Z(n19092) );
  AND U19336 ( .A(n21396), .B(n21397), .Z(n19090) );
  XOR U19337 ( .A(n19086), .B(n19087), .Z(n19089) );
  AND U19338 ( .A(n21398), .B(n21399), .Z(n19087) );
  XOR U19339 ( .A(n19083), .B(n19084), .Z(n19086) );
  AND U19340 ( .A(n21400), .B(n21401), .Z(n19084) );
  XOR U19341 ( .A(n19080), .B(n19081), .Z(n19083) );
  AND U19342 ( .A(n21402), .B(n21403), .Z(n19081) );
  XOR U19343 ( .A(n19077), .B(n19078), .Z(n19080) );
  AND U19344 ( .A(n21404), .B(n21405), .Z(n19078) );
  XOR U19345 ( .A(n19074), .B(n19075), .Z(n19077) );
  AND U19346 ( .A(n21406), .B(n21407), .Z(n19075) );
  XOR U19347 ( .A(n19071), .B(n19072), .Z(n19074) );
  AND U19348 ( .A(n21408), .B(n21409), .Z(n19072) );
  XOR U19349 ( .A(n19068), .B(n19069), .Z(n19071) );
  AND U19350 ( .A(n21410), .B(n21411), .Z(n19069) );
  XOR U19351 ( .A(n19065), .B(n19066), .Z(n19068) );
  AND U19352 ( .A(n21412), .B(n21413), .Z(n19066) );
  XOR U19353 ( .A(n19062), .B(n19063), .Z(n19065) );
  AND U19354 ( .A(n21414), .B(n21415), .Z(n19063) );
  XOR U19355 ( .A(n19059), .B(n19060), .Z(n19062) );
  AND U19356 ( .A(n21416), .B(n21417), .Z(n19060) );
  XOR U19357 ( .A(n19056), .B(n19057), .Z(n19059) );
  AND U19358 ( .A(n21418), .B(n21419), .Z(n19057) );
  XOR U19359 ( .A(n19053), .B(n19054), .Z(n19056) );
  AND U19360 ( .A(n21420), .B(n21421), .Z(n19054) );
  XOR U19361 ( .A(n19050), .B(n19051), .Z(n19053) );
  AND U19362 ( .A(n21422), .B(n21423), .Z(n19051) );
  XOR U19363 ( .A(n19047), .B(n19048), .Z(n19050) );
  AND U19364 ( .A(n21424), .B(n21425), .Z(n19048) );
  XOR U19365 ( .A(n19044), .B(n19045), .Z(n19047) );
  AND U19366 ( .A(n21426), .B(n21427), .Z(n19045) );
  XOR U19367 ( .A(n19041), .B(n19042), .Z(n19044) );
  AND U19368 ( .A(n21428), .B(n21429), .Z(n19042) );
  XOR U19369 ( .A(n19038), .B(n19039), .Z(n19041) );
  AND U19370 ( .A(n21430), .B(n21431), .Z(n19039) );
  XOR U19371 ( .A(n19035), .B(n19036), .Z(n19038) );
  AND U19372 ( .A(n21432), .B(n21433), .Z(n19036) );
  XOR U19373 ( .A(n19032), .B(n19033), .Z(n19035) );
  AND U19374 ( .A(n21434), .B(n21435), .Z(n19033) );
  XOR U19375 ( .A(n19029), .B(n19030), .Z(n19032) );
  AND U19376 ( .A(n21436), .B(n21437), .Z(n19030) );
  XOR U19377 ( .A(n19026), .B(n19027), .Z(n19029) );
  AND U19378 ( .A(n21438), .B(n21439), .Z(n19027) );
  XOR U19379 ( .A(n19023), .B(n19024), .Z(n19026) );
  AND U19380 ( .A(n21440), .B(n21441), .Z(n19024) );
  XOR U19381 ( .A(n19020), .B(n19021), .Z(n19023) );
  AND U19382 ( .A(n21442), .B(n21443), .Z(n19021) );
  XOR U19383 ( .A(n19017), .B(n19018), .Z(n19020) );
  AND U19384 ( .A(n21444), .B(n21445), .Z(n19018) );
  XOR U19385 ( .A(n19014), .B(n19015), .Z(n19017) );
  AND U19386 ( .A(n21446), .B(n21447), .Z(n19015) );
  XOR U19387 ( .A(n19011), .B(n19012), .Z(n19014) );
  AND U19388 ( .A(n21448), .B(n21449), .Z(n19012) );
  XOR U19389 ( .A(n19008), .B(n19009), .Z(n19011) );
  AND U19390 ( .A(n21450), .B(n21451), .Z(n19009) );
  XOR U19391 ( .A(n19005), .B(n19006), .Z(n19008) );
  AND U19392 ( .A(n21452), .B(n21453), .Z(n19006) );
  XOR U19393 ( .A(n19002), .B(n19003), .Z(n19005) );
  AND U19394 ( .A(n21454), .B(n21455), .Z(n19003) );
  XOR U19395 ( .A(n18999), .B(n19000), .Z(n19002) );
  AND U19396 ( .A(n21456), .B(n21457), .Z(n19000) );
  XOR U19397 ( .A(n18996), .B(n18997), .Z(n18999) );
  AND U19398 ( .A(n21458), .B(n21459), .Z(n18997) );
  XOR U19399 ( .A(n18993), .B(n18994), .Z(n18996) );
  AND U19400 ( .A(n21460), .B(n21461), .Z(n18994) );
  XOR U19401 ( .A(n18990), .B(n18991), .Z(n18993) );
  AND U19402 ( .A(n21462), .B(n21463), .Z(n18991) );
  XOR U19403 ( .A(n18987), .B(n18988), .Z(n18990) );
  AND U19404 ( .A(n21464), .B(n21465), .Z(n18988) );
  XOR U19405 ( .A(n18984), .B(n18985), .Z(n18987) );
  AND U19406 ( .A(n21466), .B(n21467), .Z(n18985) );
  XOR U19407 ( .A(n18981), .B(n18982), .Z(n18984) );
  AND U19408 ( .A(n21468), .B(n21469), .Z(n18982) );
  XOR U19409 ( .A(n18978), .B(n18979), .Z(n18981) );
  AND U19410 ( .A(n21470), .B(n21471), .Z(n18979) );
  XOR U19411 ( .A(n18975), .B(n18976), .Z(n18978) );
  AND U19412 ( .A(n21472), .B(n21473), .Z(n18976) );
  XOR U19413 ( .A(n18972), .B(n18973), .Z(n18975) );
  AND U19414 ( .A(n21474), .B(n21475), .Z(n18973) );
  XOR U19415 ( .A(n18969), .B(n18970), .Z(n18972) );
  AND U19416 ( .A(n21476), .B(n21477), .Z(n18970) );
  XOR U19417 ( .A(n18966), .B(n18967), .Z(n18969) );
  AND U19418 ( .A(n21478), .B(n21479), .Z(n18967) );
  XOR U19419 ( .A(n18963), .B(n18964), .Z(n18966) );
  AND U19420 ( .A(n21480), .B(n21481), .Z(n18964) );
  XOR U19421 ( .A(n18960), .B(n18961), .Z(n18963) );
  AND U19422 ( .A(n21482), .B(n21483), .Z(n18961) );
  XOR U19423 ( .A(n18957), .B(n18958), .Z(n18960) );
  AND U19424 ( .A(n21484), .B(n21485), .Z(n18958) );
  XOR U19425 ( .A(n18954), .B(n18955), .Z(n18957) );
  AND U19426 ( .A(n21486), .B(n21487), .Z(n18955) );
  XOR U19427 ( .A(n18951), .B(n18952), .Z(n18954) );
  AND U19428 ( .A(n21488), .B(n21489), .Z(n18952) );
  XOR U19429 ( .A(n18948), .B(n18949), .Z(n18951) );
  AND U19430 ( .A(n21490), .B(n21491), .Z(n18949) );
  XOR U19431 ( .A(n18945), .B(n18946), .Z(n18948) );
  AND U19432 ( .A(n21492), .B(n21493), .Z(n18946) );
  XOR U19433 ( .A(n18942), .B(n18943), .Z(n18945) );
  AND U19434 ( .A(n21494), .B(n21495), .Z(n18943) );
  XOR U19435 ( .A(n18939), .B(n18940), .Z(n18942) );
  AND U19436 ( .A(n21496), .B(n21497), .Z(n18940) );
  XOR U19437 ( .A(n18936), .B(n18937), .Z(n18939) );
  AND U19438 ( .A(n21498), .B(n21499), .Z(n18937) );
  XOR U19439 ( .A(n18933), .B(n18934), .Z(n18936) );
  AND U19440 ( .A(n21500), .B(n21501), .Z(n18934) );
  XOR U19441 ( .A(n18930), .B(n18931), .Z(n18933) );
  AND U19442 ( .A(n21502), .B(n21503), .Z(n18931) );
  XOR U19443 ( .A(n18927), .B(n18928), .Z(n18930) );
  AND U19444 ( .A(n21504), .B(n21505), .Z(n18928) );
  XOR U19445 ( .A(n18924), .B(n18925), .Z(n18927) );
  AND U19446 ( .A(n21506), .B(n21507), .Z(n18925) );
  XOR U19447 ( .A(n18921), .B(n18922), .Z(n18924) );
  AND U19448 ( .A(n21508), .B(n21509), .Z(n18922) );
  XOR U19449 ( .A(n18918), .B(n18919), .Z(n18921) );
  AND U19450 ( .A(n21510), .B(n21511), .Z(n18919) );
  XOR U19451 ( .A(n18915), .B(n18916), .Z(n18918) );
  AND U19452 ( .A(n21512), .B(n21513), .Z(n18916) );
  XOR U19453 ( .A(n18912), .B(n18913), .Z(n18915) );
  AND U19454 ( .A(n21514), .B(n21515), .Z(n18913) );
  XOR U19455 ( .A(n18909), .B(n18910), .Z(n18912) );
  AND U19456 ( .A(n21516), .B(n21517), .Z(n18910) );
  XOR U19457 ( .A(n18906), .B(n18907), .Z(n18909) );
  AND U19458 ( .A(n21518), .B(n21519), .Z(n18907) );
  XOR U19459 ( .A(n18903), .B(n18904), .Z(n18906) );
  AND U19460 ( .A(n21520), .B(n21521), .Z(n18904) );
  XOR U19461 ( .A(n18900), .B(n18901), .Z(n18903) );
  AND U19462 ( .A(n21522), .B(n21523), .Z(n18901) );
  XOR U19463 ( .A(n18897), .B(n18898), .Z(n18900) );
  AND U19464 ( .A(n21524), .B(n21525), .Z(n18898) );
  XOR U19465 ( .A(n18894), .B(n18895), .Z(n18897) );
  AND U19466 ( .A(n21526), .B(n21527), .Z(n18895) );
  XOR U19467 ( .A(n18891), .B(n18892), .Z(n18894) );
  AND U19468 ( .A(n21528), .B(n21529), .Z(n18892) );
  XOR U19469 ( .A(n18888), .B(n18889), .Z(n18891) );
  AND U19470 ( .A(n21530), .B(n21531), .Z(n18889) );
  XOR U19471 ( .A(n18885), .B(n18886), .Z(n18888) );
  AND U19472 ( .A(n21532), .B(n21533), .Z(n18886) );
  XOR U19473 ( .A(n18882), .B(n18883), .Z(n18885) );
  AND U19474 ( .A(n21534), .B(n21535), .Z(n18883) );
  XOR U19475 ( .A(n18879), .B(n18880), .Z(n18882) );
  AND U19476 ( .A(n21536), .B(n21537), .Z(n18880) );
  XOR U19477 ( .A(n18876), .B(n18877), .Z(n18879) );
  AND U19478 ( .A(n21538), .B(n21539), .Z(n18877) );
  XOR U19479 ( .A(n18873), .B(n18874), .Z(n18876) );
  AND U19480 ( .A(n21540), .B(n21541), .Z(n18874) );
  XOR U19481 ( .A(n18870), .B(n18871), .Z(n18873) );
  AND U19482 ( .A(n21542), .B(n21543), .Z(n18871) );
  XOR U19483 ( .A(n18867), .B(n18868), .Z(n18870) );
  AND U19484 ( .A(n21544), .B(n21545), .Z(n18868) );
  XOR U19485 ( .A(n18864), .B(n18865), .Z(n18867) );
  AND U19486 ( .A(n21546), .B(n21547), .Z(n18865) );
  XOR U19487 ( .A(n18861), .B(n18862), .Z(n18864) );
  AND U19488 ( .A(n21548), .B(n21549), .Z(n18862) );
  XOR U19489 ( .A(n18858), .B(n18859), .Z(n18861) );
  AND U19490 ( .A(n21550), .B(n21551), .Z(n18859) );
  XOR U19491 ( .A(n18855), .B(n18856), .Z(n18858) );
  AND U19492 ( .A(n21552), .B(n21553), .Z(n18856) );
  XOR U19493 ( .A(n18852), .B(n18853), .Z(n18855) );
  AND U19494 ( .A(n21554), .B(n21555), .Z(n18853) );
  XOR U19495 ( .A(n18849), .B(n18850), .Z(n18852) );
  AND U19496 ( .A(n21556), .B(n21557), .Z(n18850) );
  XOR U19497 ( .A(n18846), .B(n18847), .Z(n18849) );
  AND U19498 ( .A(n21558), .B(n21559), .Z(n18847) );
  XOR U19499 ( .A(n18843), .B(n18844), .Z(n18846) );
  AND U19500 ( .A(n21560), .B(n21561), .Z(n18844) );
  XOR U19501 ( .A(n18840), .B(n18841), .Z(n18843) );
  AND U19502 ( .A(n21562), .B(n21563), .Z(n18841) );
  XOR U19503 ( .A(n18837), .B(n18838), .Z(n18840) );
  AND U19504 ( .A(n21564), .B(n21565), .Z(n18838) );
  XOR U19505 ( .A(n18834), .B(n18835), .Z(n18837) );
  AND U19506 ( .A(n21566), .B(n21567), .Z(n18835) );
  XOR U19507 ( .A(n18831), .B(n18832), .Z(n18834) );
  AND U19508 ( .A(n21568), .B(n21569), .Z(n18832) );
  XOR U19509 ( .A(n18828), .B(n18829), .Z(n18831) );
  AND U19510 ( .A(n21570), .B(n21571), .Z(n18829) );
  XOR U19511 ( .A(n18825), .B(n18826), .Z(n18828) );
  AND U19512 ( .A(n21572), .B(n21573), .Z(n18826) );
  XOR U19513 ( .A(n18822), .B(n18823), .Z(n18825) );
  AND U19514 ( .A(n21574), .B(n21575), .Z(n18823) );
  XOR U19515 ( .A(n18819), .B(n18820), .Z(n18822) );
  AND U19516 ( .A(n21576), .B(n21577), .Z(n18820) );
  XOR U19517 ( .A(n18816), .B(n18817), .Z(n18819) );
  AND U19518 ( .A(n21578), .B(n21579), .Z(n18817) );
  XOR U19519 ( .A(n18813), .B(n18814), .Z(n18816) );
  AND U19520 ( .A(n21580), .B(n21581), .Z(n18814) );
  XOR U19521 ( .A(n18810), .B(n18811), .Z(n18813) );
  AND U19522 ( .A(n21582), .B(n21583), .Z(n18811) );
  XOR U19523 ( .A(n18807), .B(n18808), .Z(n18810) );
  AND U19524 ( .A(n21584), .B(n21585), .Z(n18808) );
  XOR U19525 ( .A(n18804), .B(n18805), .Z(n18807) );
  AND U19526 ( .A(n21586), .B(n21587), .Z(n18805) );
  XOR U19527 ( .A(n18801), .B(n18802), .Z(n18804) );
  AND U19528 ( .A(n21588), .B(n21589), .Z(n18802) );
  XOR U19529 ( .A(n18798), .B(n18799), .Z(n18801) );
  AND U19530 ( .A(n21590), .B(n21591), .Z(n18799) );
  XOR U19531 ( .A(n18795), .B(n18796), .Z(n18798) );
  AND U19532 ( .A(n21592), .B(n21593), .Z(n18796) );
  XOR U19533 ( .A(n18792), .B(n18793), .Z(n18795) );
  AND U19534 ( .A(n21594), .B(n21595), .Z(n18793) );
  XOR U19535 ( .A(n18789), .B(n18790), .Z(n18792) );
  AND U19536 ( .A(n21596), .B(n21597), .Z(n18790) );
  XOR U19537 ( .A(n18786), .B(n18787), .Z(n18789) );
  AND U19538 ( .A(n21598), .B(n21599), .Z(n18787) );
  XOR U19539 ( .A(n18783), .B(n18784), .Z(n18786) );
  AND U19540 ( .A(n21600), .B(n21601), .Z(n18784) );
  XOR U19541 ( .A(n18780), .B(n18781), .Z(n18783) );
  AND U19542 ( .A(n21602), .B(n21603), .Z(n18781) );
  XOR U19543 ( .A(n18777), .B(n18778), .Z(n18780) );
  AND U19544 ( .A(n21604), .B(n21605), .Z(n18778) );
  XOR U19545 ( .A(n18774), .B(n18775), .Z(n18777) );
  AND U19546 ( .A(n21606), .B(n21607), .Z(n18775) );
  XOR U19547 ( .A(n18771), .B(n18772), .Z(n18774) );
  AND U19548 ( .A(n21608), .B(n21609), .Z(n18772) );
  XOR U19549 ( .A(n18768), .B(n18769), .Z(n18771) );
  AND U19550 ( .A(n21610), .B(n21611), .Z(n18769) );
  XOR U19551 ( .A(n18765), .B(n18766), .Z(n18768) );
  AND U19552 ( .A(n21612), .B(n21613), .Z(n18766) );
  XOR U19553 ( .A(n18762), .B(n18763), .Z(n18765) );
  AND U19554 ( .A(n21614), .B(n21615), .Z(n18763) );
  XOR U19555 ( .A(n18759), .B(n18760), .Z(n18762) );
  AND U19556 ( .A(n21616), .B(n21617), .Z(n18760) );
  XOR U19557 ( .A(n18756), .B(n18757), .Z(n18759) );
  AND U19558 ( .A(n21618), .B(n21619), .Z(n18757) );
  XOR U19559 ( .A(n18753), .B(n18754), .Z(n18756) );
  AND U19560 ( .A(n21620), .B(n21621), .Z(n18754) );
  XOR U19561 ( .A(n18750), .B(n18751), .Z(n18753) );
  AND U19562 ( .A(n21622), .B(n21623), .Z(n18751) );
  XOR U19563 ( .A(n18747), .B(n18748), .Z(n18750) );
  AND U19564 ( .A(n21624), .B(n21625), .Z(n18748) );
  XOR U19565 ( .A(n18744), .B(n18745), .Z(n18747) );
  AND U19566 ( .A(n21626), .B(n21627), .Z(n18745) );
  XOR U19567 ( .A(n18741), .B(n18742), .Z(n18744) );
  AND U19568 ( .A(n21628), .B(n21629), .Z(n18742) );
  XOR U19569 ( .A(n18738), .B(n18739), .Z(n18741) );
  AND U19570 ( .A(n21630), .B(n21631), .Z(n18739) );
  XOR U19571 ( .A(n18735), .B(n18736), .Z(n18738) );
  AND U19572 ( .A(n21632), .B(n21633), .Z(n18736) );
  XOR U19573 ( .A(n18732), .B(n18733), .Z(n18735) );
  AND U19574 ( .A(n21634), .B(n21635), .Z(n18733) );
  XOR U19575 ( .A(n18729), .B(n18730), .Z(n18732) );
  AND U19576 ( .A(n21636), .B(n21637), .Z(n18730) );
  XOR U19577 ( .A(n18726), .B(n18727), .Z(n18729) );
  AND U19578 ( .A(n21638), .B(n21639), .Z(n18727) );
  XOR U19579 ( .A(n18723), .B(n18724), .Z(n18726) );
  AND U19580 ( .A(n21640), .B(n21641), .Z(n18724) );
  XOR U19581 ( .A(n18720), .B(n18721), .Z(n18723) );
  AND U19582 ( .A(n21642), .B(n21643), .Z(n18721) );
  XOR U19583 ( .A(n18717), .B(n18718), .Z(n18720) );
  AND U19584 ( .A(n21644), .B(n21645), .Z(n18718) );
  XOR U19585 ( .A(n18714), .B(n18715), .Z(n18717) );
  AND U19586 ( .A(n21646), .B(n21647), .Z(n18715) );
  XOR U19587 ( .A(n18711), .B(n18712), .Z(n18714) );
  AND U19588 ( .A(n21648), .B(n21649), .Z(n18712) );
  XOR U19589 ( .A(n18708), .B(n18709), .Z(n18711) );
  AND U19590 ( .A(n21650), .B(n21651), .Z(n18709) );
  XOR U19591 ( .A(n18705), .B(n18706), .Z(n18708) );
  AND U19592 ( .A(n21652), .B(n21653), .Z(n18706) );
  XOR U19593 ( .A(n18702), .B(n18703), .Z(n18705) );
  AND U19594 ( .A(n21654), .B(n21655), .Z(n18703) );
  XNOR U19595 ( .A(n18699), .B(n18700), .Z(n18702) );
  AND U19596 ( .A(n21656), .B(n21657), .Z(n18700) );
  XOR U19597 ( .A(n21658), .B(n18697), .Z(n18699) );
  IV U19598 ( .A(n21659), .Z(n18697) );
  AND U19599 ( .A(n21660), .B(n21661), .Z(n21659) );
  IV U19600 ( .A(n18696), .Z(n21658) );
  XOR U19601 ( .A(n18437), .B(n18693), .Z(n18696) );
  AND U19602 ( .A(n21662), .B(n21663), .Z(n18693) );
  XOR U19603 ( .A(n18439), .B(n18438), .Z(n18437) );
  AND U19604 ( .A(n21664), .B(n21665), .Z(n18438) );
  XOR U19605 ( .A(n18441), .B(n18440), .Z(n18439) );
  AND U19606 ( .A(n21666), .B(n21667), .Z(n18440) );
  XOR U19607 ( .A(n18443), .B(n18442), .Z(n18441) );
  AND U19608 ( .A(n21668), .B(n21669), .Z(n18442) );
  XOR U19609 ( .A(n18445), .B(n18444), .Z(n18443) );
  AND U19610 ( .A(n21670), .B(n21671), .Z(n18444) );
  XOR U19611 ( .A(n18447), .B(n18446), .Z(n18445) );
  AND U19612 ( .A(n21672), .B(n21673), .Z(n18446) );
  XOR U19613 ( .A(n18449), .B(n18448), .Z(n18447) );
  AND U19614 ( .A(n21674), .B(n21675), .Z(n18448) );
  XOR U19615 ( .A(n18451), .B(n18450), .Z(n18449) );
  AND U19616 ( .A(n21676), .B(n21677), .Z(n18450) );
  XOR U19617 ( .A(n18453), .B(n18452), .Z(n18451) );
  AND U19618 ( .A(n21678), .B(n21679), .Z(n18452) );
  XOR U19619 ( .A(n18455), .B(n18454), .Z(n18453) );
  AND U19620 ( .A(n21680), .B(n21681), .Z(n18454) );
  XOR U19621 ( .A(n18457), .B(n18456), .Z(n18455) );
  AND U19622 ( .A(n21682), .B(n21683), .Z(n18456) );
  XOR U19623 ( .A(n18459), .B(n18458), .Z(n18457) );
  AND U19624 ( .A(n21684), .B(n21685), .Z(n18458) );
  XOR U19625 ( .A(n18461), .B(n18460), .Z(n18459) );
  AND U19626 ( .A(n21686), .B(n21687), .Z(n18460) );
  XOR U19627 ( .A(n18463), .B(n18462), .Z(n18461) );
  AND U19628 ( .A(n21688), .B(n21689), .Z(n18462) );
  XOR U19629 ( .A(n18465), .B(n18464), .Z(n18463) );
  AND U19630 ( .A(n21690), .B(n21691), .Z(n18464) );
  XOR U19631 ( .A(n18467), .B(n18466), .Z(n18465) );
  AND U19632 ( .A(n21692), .B(n21693), .Z(n18466) );
  XOR U19633 ( .A(n18469), .B(n18468), .Z(n18467) );
  AND U19634 ( .A(n21694), .B(n21695), .Z(n18468) );
  XOR U19635 ( .A(n18471), .B(n18470), .Z(n18469) );
  AND U19636 ( .A(n21696), .B(n21697), .Z(n18470) );
  XOR U19637 ( .A(n18473), .B(n18472), .Z(n18471) );
  AND U19638 ( .A(n21698), .B(n21699), .Z(n18472) );
  XOR U19639 ( .A(n18475), .B(n18474), .Z(n18473) );
  AND U19640 ( .A(n21700), .B(n21701), .Z(n18474) );
  XOR U19641 ( .A(n18477), .B(n18476), .Z(n18475) );
  AND U19642 ( .A(n21702), .B(n21703), .Z(n18476) );
  XOR U19643 ( .A(n18479), .B(n18478), .Z(n18477) );
  AND U19644 ( .A(n21704), .B(n21705), .Z(n18478) );
  XOR U19645 ( .A(n18481), .B(n18480), .Z(n18479) );
  AND U19646 ( .A(n21706), .B(n21707), .Z(n18480) );
  XOR U19647 ( .A(n18483), .B(n18482), .Z(n18481) );
  AND U19648 ( .A(n21708), .B(n21709), .Z(n18482) );
  XOR U19649 ( .A(n18485), .B(n18484), .Z(n18483) );
  AND U19650 ( .A(n21710), .B(n21711), .Z(n18484) );
  XOR U19651 ( .A(n18487), .B(n18486), .Z(n18485) );
  AND U19652 ( .A(n21712), .B(n21713), .Z(n18486) );
  XOR U19653 ( .A(n18489), .B(n18488), .Z(n18487) );
  AND U19654 ( .A(n21714), .B(n21715), .Z(n18488) );
  XOR U19655 ( .A(n18491), .B(n18490), .Z(n18489) );
  AND U19656 ( .A(n21716), .B(n21717), .Z(n18490) );
  XOR U19657 ( .A(n18493), .B(n18492), .Z(n18491) );
  AND U19658 ( .A(n21718), .B(n21719), .Z(n18492) );
  XOR U19659 ( .A(n18495), .B(n18494), .Z(n18493) );
  AND U19660 ( .A(n21720), .B(n21721), .Z(n18494) );
  XOR U19661 ( .A(n18497), .B(n18496), .Z(n18495) );
  AND U19662 ( .A(n21722), .B(n21723), .Z(n18496) );
  XOR U19663 ( .A(n18499), .B(n18498), .Z(n18497) );
  AND U19664 ( .A(n21724), .B(n21725), .Z(n18498) );
  XOR U19665 ( .A(n18501), .B(n18500), .Z(n18499) );
  AND U19666 ( .A(n21726), .B(n21727), .Z(n18500) );
  XOR U19667 ( .A(n18503), .B(n18502), .Z(n18501) );
  AND U19668 ( .A(n21728), .B(n21729), .Z(n18502) );
  XOR U19669 ( .A(n18505), .B(n18504), .Z(n18503) );
  AND U19670 ( .A(n21730), .B(n21731), .Z(n18504) );
  XOR U19671 ( .A(n18507), .B(n18506), .Z(n18505) );
  AND U19672 ( .A(n21732), .B(n21733), .Z(n18506) );
  XOR U19673 ( .A(n18509), .B(n18508), .Z(n18507) );
  AND U19674 ( .A(n21734), .B(n21735), .Z(n18508) );
  XOR U19675 ( .A(n18511), .B(n18510), .Z(n18509) );
  AND U19676 ( .A(n21736), .B(n21737), .Z(n18510) );
  XOR U19677 ( .A(n18513), .B(n18512), .Z(n18511) );
  AND U19678 ( .A(n21738), .B(n21739), .Z(n18512) );
  XOR U19679 ( .A(n18515), .B(n18514), .Z(n18513) );
  AND U19680 ( .A(n21740), .B(n21741), .Z(n18514) );
  XOR U19681 ( .A(n18517), .B(n18516), .Z(n18515) );
  AND U19682 ( .A(n21742), .B(n21743), .Z(n18516) );
  XOR U19683 ( .A(n18519), .B(n18518), .Z(n18517) );
  AND U19684 ( .A(n21744), .B(n21745), .Z(n18518) );
  XOR U19685 ( .A(n18521), .B(n18520), .Z(n18519) );
  AND U19686 ( .A(n21746), .B(n21747), .Z(n18520) );
  XOR U19687 ( .A(n18523), .B(n18522), .Z(n18521) );
  AND U19688 ( .A(n21748), .B(n21749), .Z(n18522) );
  XOR U19689 ( .A(n18525), .B(n18524), .Z(n18523) );
  AND U19690 ( .A(n21750), .B(n21751), .Z(n18524) );
  XOR U19691 ( .A(n18527), .B(n18526), .Z(n18525) );
  AND U19692 ( .A(n21752), .B(n21753), .Z(n18526) );
  XOR U19693 ( .A(n18529), .B(n18528), .Z(n18527) );
  AND U19694 ( .A(n21754), .B(n21755), .Z(n18528) );
  XOR U19695 ( .A(n18531), .B(n18530), .Z(n18529) );
  AND U19696 ( .A(n21756), .B(n21757), .Z(n18530) );
  XOR U19697 ( .A(n18533), .B(n18532), .Z(n18531) );
  AND U19698 ( .A(n21758), .B(n21759), .Z(n18532) );
  XOR U19699 ( .A(n18535), .B(n18534), .Z(n18533) );
  AND U19700 ( .A(n21760), .B(n21761), .Z(n18534) );
  XOR U19701 ( .A(n18537), .B(n18536), .Z(n18535) );
  AND U19702 ( .A(n21762), .B(n21763), .Z(n18536) );
  XOR U19703 ( .A(n18539), .B(n18538), .Z(n18537) );
  AND U19704 ( .A(n21764), .B(n21765), .Z(n18538) );
  XOR U19705 ( .A(n18541), .B(n18540), .Z(n18539) );
  AND U19706 ( .A(n21766), .B(n21767), .Z(n18540) );
  XOR U19707 ( .A(n18543), .B(n18542), .Z(n18541) );
  AND U19708 ( .A(n21768), .B(n21769), .Z(n18542) );
  XOR U19709 ( .A(n18545), .B(n18544), .Z(n18543) );
  AND U19710 ( .A(n21770), .B(n21771), .Z(n18544) );
  XOR U19711 ( .A(n18547), .B(n18546), .Z(n18545) );
  AND U19712 ( .A(n21772), .B(n21773), .Z(n18546) );
  XOR U19713 ( .A(n18549), .B(n18548), .Z(n18547) );
  AND U19714 ( .A(n21774), .B(n21775), .Z(n18548) );
  XOR U19715 ( .A(n18551), .B(n18550), .Z(n18549) );
  AND U19716 ( .A(n21776), .B(n21777), .Z(n18550) );
  XOR U19717 ( .A(n18553), .B(n18552), .Z(n18551) );
  AND U19718 ( .A(n21778), .B(n21779), .Z(n18552) );
  XOR U19719 ( .A(n18555), .B(n18554), .Z(n18553) );
  AND U19720 ( .A(n21780), .B(n21781), .Z(n18554) );
  XOR U19721 ( .A(n18557), .B(n18556), .Z(n18555) );
  AND U19722 ( .A(n21782), .B(n21783), .Z(n18556) );
  XOR U19723 ( .A(n18559), .B(n18558), .Z(n18557) );
  AND U19724 ( .A(n21784), .B(n21785), .Z(n18558) );
  XOR U19725 ( .A(n18561), .B(n18560), .Z(n18559) );
  AND U19726 ( .A(n21786), .B(n21787), .Z(n18560) );
  XOR U19727 ( .A(n18563), .B(n18562), .Z(n18561) );
  AND U19728 ( .A(n21788), .B(n21789), .Z(n18562) );
  XOR U19729 ( .A(n18565), .B(n18564), .Z(n18563) );
  AND U19730 ( .A(n21790), .B(n21791), .Z(n18564) );
  XOR U19731 ( .A(n18567), .B(n18566), .Z(n18565) );
  AND U19732 ( .A(n21792), .B(n21793), .Z(n18566) );
  XOR U19733 ( .A(n18569), .B(n18568), .Z(n18567) );
  AND U19734 ( .A(n21794), .B(n21795), .Z(n18568) );
  XOR U19735 ( .A(n18571), .B(n18570), .Z(n18569) );
  AND U19736 ( .A(n21796), .B(n21797), .Z(n18570) );
  XOR U19737 ( .A(n18573), .B(n18572), .Z(n18571) );
  AND U19738 ( .A(n21798), .B(n21799), .Z(n18572) );
  XOR U19739 ( .A(n18575), .B(n18574), .Z(n18573) );
  AND U19740 ( .A(n21800), .B(n21801), .Z(n18574) );
  XOR U19741 ( .A(n18577), .B(n18576), .Z(n18575) );
  AND U19742 ( .A(n21802), .B(n21803), .Z(n18576) );
  XOR U19743 ( .A(n18579), .B(n18578), .Z(n18577) );
  AND U19744 ( .A(n21804), .B(n21805), .Z(n18578) );
  XOR U19745 ( .A(n18581), .B(n18580), .Z(n18579) );
  AND U19746 ( .A(n21806), .B(n21807), .Z(n18580) );
  XOR U19747 ( .A(n18583), .B(n18582), .Z(n18581) );
  AND U19748 ( .A(n21808), .B(n21809), .Z(n18582) );
  XOR U19749 ( .A(n18585), .B(n18584), .Z(n18583) );
  AND U19750 ( .A(n21810), .B(n21811), .Z(n18584) );
  XOR U19751 ( .A(n18587), .B(n18586), .Z(n18585) );
  AND U19752 ( .A(n21812), .B(n21813), .Z(n18586) );
  XOR U19753 ( .A(n18589), .B(n18588), .Z(n18587) );
  AND U19754 ( .A(n21814), .B(n21815), .Z(n18588) );
  XOR U19755 ( .A(n18591), .B(n18590), .Z(n18589) );
  AND U19756 ( .A(n21816), .B(n21817), .Z(n18590) );
  XOR U19757 ( .A(n18593), .B(n18592), .Z(n18591) );
  AND U19758 ( .A(n21818), .B(n21819), .Z(n18592) );
  XOR U19759 ( .A(n18595), .B(n18594), .Z(n18593) );
  AND U19760 ( .A(n21820), .B(n21821), .Z(n18594) );
  XOR U19761 ( .A(n18597), .B(n18596), .Z(n18595) );
  AND U19762 ( .A(n21822), .B(n21823), .Z(n18596) );
  XOR U19763 ( .A(n18599), .B(n18598), .Z(n18597) );
  AND U19764 ( .A(n21824), .B(n21825), .Z(n18598) );
  XOR U19765 ( .A(n18601), .B(n18600), .Z(n18599) );
  AND U19766 ( .A(n21826), .B(n21827), .Z(n18600) );
  XOR U19767 ( .A(n18603), .B(n18602), .Z(n18601) );
  AND U19768 ( .A(n21828), .B(n21829), .Z(n18602) );
  XOR U19769 ( .A(n18605), .B(n18604), .Z(n18603) );
  AND U19770 ( .A(n21830), .B(n21831), .Z(n18604) );
  XOR U19771 ( .A(n18607), .B(n18606), .Z(n18605) );
  AND U19772 ( .A(n21832), .B(n21833), .Z(n18606) );
  XOR U19773 ( .A(n18609), .B(n18608), .Z(n18607) );
  AND U19774 ( .A(n21834), .B(n21835), .Z(n18608) );
  XOR U19775 ( .A(n18611), .B(n18610), .Z(n18609) );
  AND U19776 ( .A(n21836), .B(n21837), .Z(n18610) );
  XOR U19777 ( .A(n18613), .B(n18612), .Z(n18611) );
  AND U19778 ( .A(n21838), .B(n21839), .Z(n18612) );
  XOR U19779 ( .A(n18615), .B(n18614), .Z(n18613) );
  AND U19780 ( .A(n21840), .B(n21841), .Z(n18614) );
  XOR U19781 ( .A(n18617), .B(n18616), .Z(n18615) );
  AND U19782 ( .A(n21842), .B(n21843), .Z(n18616) );
  XOR U19783 ( .A(n18619), .B(n18618), .Z(n18617) );
  AND U19784 ( .A(n21844), .B(n21845), .Z(n18618) );
  XOR U19785 ( .A(n18621), .B(n18620), .Z(n18619) );
  AND U19786 ( .A(n21846), .B(n21847), .Z(n18620) );
  XOR U19787 ( .A(n18623), .B(n18622), .Z(n18621) );
  AND U19788 ( .A(n21848), .B(n21849), .Z(n18622) );
  XOR U19789 ( .A(n18625), .B(n18624), .Z(n18623) );
  AND U19790 ( .A(n21850), .B(n21851), .Z(n18624) );
  XOR U19791 ( .A(n18627), .B(n18626), .Z(n18625) );
  AND U19792 ( .A(n21852), .B(n21853), .Z(n18626) );
  XOR U19793 ( .A(n18629), .B(n18628), .Z(n18627) );
  AND U19794 ( .A(n21854), .B(n21855), .Z(n18628) );
  XOR U19795 ( .A(n18631), .B(n18630), .Z(n18629) );
  AND U19796 ( .A(n21856), .B(n21857), .Z(n18630) );
  XOR U19797 ( .A(n18633), .B(n18632), .Z(n18631) );
  AND U19798 ( .A(n21858), .B(n21859), .Z(n18632) );
  XOR U19799 ( .A(n18635), .B(n18634), .Z(n18633) );
  AND U19800 ( .A(n21860), .B(n21861), .Z(n18634) );
  XOR U19801 ( .A(n18637), .B(n18636), .Z(n18635) );
  AND U19802 ( .A(n21862), .B(n21863), .Z(n18636) );
  XOR U19803 ( .A(n18639), .B(n18638), .Z(n18637) );
  AND U19804 ( .A(n21864), .B(n21865), .Z(n18638) );
  XOR U19805 ( .A(n18641), .B(n18640), .Z(n18639) );
  AND U19806 ( .A(n21866), .B(n21867), .Z(n18640) );
  XOR U19807 ( .A(n18643), .B(n18642), .Z(n18641) );
  AND U19808 ( .A(n21868), .B(n21869), .Z(n18642) );
  XOR U19809 ( .A(n18645), .B(n18644), .Z(n18643) );
  AND U19810 ( .A(n21870), .B(n21871), .Z(n18644) );
  XOR U19811 ( .A(n18647), .B(n18646), .Z(n18645) );
  AND U19812 ( .A(n21872), .B(n21873), .Z(n18646) );
  XOR U19813 ( .A(n18649), .B(n18648), .Z(n18647) );
  AND U19814 ( .A(n21874), .B(n21875), .Z(n18648) );
  XOR U19815 ( .A(n18651), .B(n18650), .Z(n18649) );
  AND U19816 ( .A(n21876), .B(n21877), .Z(n18650) );
  XOR U19817 ( .A(n18653), .B(n18652), .Z(n18651) );
  AND U19818 ( .A(n21878), .B(n21879), .Z(n18652) );
  XOR U19819 ( .A(n18655), .B(n18654), .Z(n18653) );
  AND U19820 ( .A(n21880), .B(n21881), .Z(n18654) );
  XOR U19821 ( .A(n18657), .B(n18656), .Z(n18655) );
  AND U19822 ( .A(n21882), .B(n21883), .Z(n18656) );
  XOR U19823 ( .A(n18659), .B(n18658), .Z(n18657) );
  AND U19824 ( .A(n21884), .B(n21885), .Z(n18658) );
  XOR U19825 ( .A(n18661), .B(n18660), .Z(n18659) );
  AND U19826 ( .A(n21886), .B(n21887), .Z(n18660) );
  XOR U19827 ( .A(n18689), .B(n18662), .Z(n18661) );
  AND U19828 ( .A(n21888), .B(n21889), .Z(n18662) );
  XOR U19829 ( .A(n18691), .B(n18690), .Z(n18689) );
  AND U19830 ( .A(n21890), .B(n21891), .Z(n18690) );
  XOR U19831 ( .A(n18670), .B(n18692), .Z(n18691) );
  AND U19832 ( .A(n21892), .B(n21893), .Z(n18692) );
  XOR U19833 ( .A(n18666), .B(n18671), .Z(n18670) );
  AND U19834 ( .A(n21894), .B(n21895), .Z(n18671) );
  XOR U19835 ( .A(n18668), .B(n18667), .Z(n18666) );
  AND U19836 ( .A(n21896), .B(n21897), .Z(n18667) );
  XNOR U19837 ( .A(n18678), .B(n18669), .Z(n18668) );
  AND U19838 ( .A(n21898), .B(n21899), .Z(n18669) );
  XOR U19839 ( .A(n18688), .B(n18677), .Z(n18678) );
  AND U19840 ( .A(n21900), .B(n21901), .Z(n18677) );
  XNOR U19841 ( .A(n21902), .B(n18683), .Z(n18688) );
  XOR U19842 ( .A(n18684), .B(n21903), .Z(n18683) );
  AND U19843 ( .A(n21904), .B(n21905), .Z(n21903) );
  XOR U19844 ( .A(n21906), .B(n21907), .Z(n18684) );
  NOR U19845 ( .A(n21908), .B(n21909), .Z(n21907) );
  AND U19846 ( .A(n21910), .B(n21911), .Z(n21909) );
  AND U19847 ( .A(n21912), .B(n21913), .Z(n21908) );
  XNOR U19848 ( .A(n21910), .B(n21911), .Z(n21906) );
  XNOR U19849 ( .A(n18675), .B(n18687), .Z(n21902) );
  AND U19850 ( .A(n21914), .B(n21915), .Z(n18687) );
  AND U19851 ( .A(n21916), .B(n21917), .Z(n18675) );
  AND U19852 ( .A(n143), .B(n145), .Z(n19854) );
  XOR U19853 ( .A(n19859), .B(n19858), .Z(n145) );
  NOR U19854 ( .A(n21918), .B(n21919), .Z(n19858) );
  XOR U19855 ( .A(n19861), .B(n19860), .Z(n19859) );
  NOR U19856 ( .A(n21920), .B(n21921), .Z(n19860) );
  XOR U19857 ( .A(n19863), .B(n19862), .Z(n19861) );
  NOR U19858 ( .A(n21922), .B(n21923), .Z(n19862) );
  XOR U19859 ( .A(n19865), .B(n19864), .Z(n19863) );
  NOR U19860 ( .A(n21924), .B(n21925), .Z(n19864) );
  XOR U19861 ( .A(n19867), .B(n19866), .Z(n19865) );
  NOR U19862 ( .A(n21926), .B(n21927), .Z(n19866) );
  XOR U19863 ( .A(n19869), .B(n19868), .Z(n19867) );
  NOR U19864 ( .A(n21928), .B(n21929), .Z(n19868) );
  XOR U19865 ( .A(n19871), .B(n19870), .Z(n19869) );
  NOR U19866 ( .A(n21930), .B(n21931), .Z(n19870) );
  XOR U19867 ( .A(n19873), .B(n19872), .Z(n19871) );
  NOR U19868 ( .A(n21932), .B(n21933), .Z(n19872) );
  XOR U19869 ( .A(n19875), .B(n19874), .Z(n19873) );
  NOR U19870 ( .A(n21934), .B(n21935), .Z(n19874) );
  XOR U19871 ( .A(n19877), .B(n19876), .Z(n19875) );
  NOR U19872 ( .A(n21936), .B(n21937), .Z(n19876) );
  XOR U19873 ( .A(n19879), .B(n19878), .Z(n19877) );
  NOR U19874 ( .A(n21938), .B(n21939), .Z(n19878) );
  XOR U19875 ( .A(n19881), .B(n19880), .Z(n19879) );
  NOR U19876 ( .A(n21940), .B(n21941), .Z(n19880) );
  XOR U19877 ( .A(n19883), .B(n19882), .Z(n19881) );
  NOR U19878 ( .A(n21942), .B(n21943), .Z(n19882) );
  XOR U19879 ( .A(n19885), .B(n19884), .Z(n19883) );
  NOR U19880 ( .A(n21944), .B(n21945), .Z(n19884) );
  XOR U19881 ( .A(n19887), .B(n19886), .Z(n19885) );
  NOR U19882 ( .A(n21946), .B(n21947), .Z(n19886) );
  XOR U19883 ( .A(n19889), .B(n19888), .Z(n19887) );
  NOR U19884 ( .A(n21948), .B(n21949), .Z(n19888) );
  XOR U19885 ( .A(n19891), .B(n19890), .Z(n19889) );
  NOR U19886 ( .A(n21950), .B(n21951), .Z(n19890) );
  XOR U19887 ( .A(n19893), .B(n19892), .Z(n19891) );
  NOR U19888 ( .A(n21952), .B(n21953), .Z(n19892) );
  XOR U19889 ( .A(n19895), .B(n19894), .Z(n19893) );
  NOR U19890 ( .A(n21954), .B(n21955), .Z(n19894) );
  XOR U19891 ( .A(n19897), .B(n19896), .Z(n19895) );
  NOR U19892 ( .A(n21956), .B(n21957), .Z(n19896) );
  XOR U19893 ( .A(n19899), .B(n19898), .Z(n19897) );
  NOR U19894 ( .A(n21958), .B(n21959), .Z(n19898) );
  XOR U19895 ( .A(n19901), .B(n19900), .Z(n19899) );
  NOR U19896 ( .A(n21960), .B(n21961), .Z(n19900) );
  XOR U19897 ( .A(n19903), .B(n19902), .Z(n19901) );
  NOR U19898 ( .A(n21962), .B(n21963), .Z(n19902) );
  XOR U19899 ( .A(n19905), .B(n19904), .Z(n19903) );
  NOR U19900 ( .A(n21964), .B(n21965), .Z(n19904) );
  XOR U19901 ( .A(n19907), .B(n19906), .Z(n19905) );
  NOR U19902 ( .A(n21966), .B(n21967), .Z(n19906) );
  XOR U19903 ( .A(n19909), .B(n19908), .Z(n19907) );
  NOR U19904 ( .A(n21968), .B(n21969), .Z(n19908) );
  XOR U19905 ( .A(n19911), .B(n19910), .Z(n19909) );
  NOR U19906 ( .A(n21970), .B(n21971), .Z(n19910) );
  XOR U19907 ( .A(n19913), .B(n19912), .Z(n19911) );
  NOR U19908 ( .A(n21972), .B(n21973), .Z(n19912) );
  XOR U19909 ( .A(n19915), .B(n19914), .Z(n19913) );
  NOR U19910 ( .A(n21974), .B(n21975), .Z(n19914) );
  XOR U19911 ( .A(n19917), .B(n19916), .Z(n19915) );
  NOR U19912 ( .A(n21976), .B(n21977), .Z(n19916) );
  XOR U19913 ( .A(n19919), .B(n19918), .Z(n19917) );
  NOR U19914 ( .A(n21978), .B(n21979), .Z(n19918) );
  XOR U19915 ( .A(n19921), .B(n19920), .Z(n19919) );
  NOR U19916 ( .A(n21980), .B(n21981), .Z(n19920) );
  XOR U19917 ( .A(n19923), .B(n19922), .Z(n19921) );
  NOR U19918 ( .A(n21982), .B(n21983), .Z(n19922) );
  XOR U19919 ( .A(n19925), .B(n19924), .Z(n19923) );
  NOR U19920 ( .A(n21984), .B(n21985), .Z(n19924) );
  XOR U19921 ( .A(n19927), .B(n19926), .Z(n19925) );
  NOR U19922 ( .A(n21986), .B(n21987), .Z(n19926) );
  XOR U19923 ( .A(n19929), .B(n19928), .Z(n19927) );
  NOR U19924 ( .A(n21988), .B(n21989), .Z(n19928) );
  XOR U19925 ( .A(n19931), .B(n19930), .Z(n19929) );
  NOR U19926 ( .A(n21990), .B(n21991), .Z(n19930) );
  XOR U19927 ( .A(n19933), .B(n19932), .Z(n19931) );
  NOR U19928 ( .A(n21992), .B(n21993), .Z(n19932) );
  XOR U19929 ( .A(n19935), .B(n19934), .Z(n19933) );
  NOR U19930 ( .A(n21994), .B(n21995), .Z(n19934) );
  XOR U19931 ( .A(n19937), .B(n19936), .Z(n19935) );
  NOR U19932 ( .A(n21996), .B(n21997), .Z(n19936) );
  XOR U19933 ( .A(n19939), .B(n19938), .Z(n19937) );
  NOR U19934 ( .A(n21998), .B(n21999), .Z(n19938) );
  XOR U19935 ( .A(n19941), .B(n19940), .Z(n19939) );
  NOR U19936 ( .A(n22000), .B(n22001), .Z(n19940) );
  XOR U19937 ( .A(n19943), .B(n19942), .Z(n19941) );
  NOR U19938 ( .A(n22002), .B(n22003), .Z(n19942) );
  XOR U19939 ( .A(n19945), .B(n19944), .Z(n19943) );
  NOR U19940 ( .A(n22004), .B(n22005), .Z(n19944) );
  XOR U19941 ( .A(n19947), .B(n19946), .Z(n19945) );
  NOR U19942 ( .A(n22006), .B(n22007), .Z(n19946) );
  XOR U19943 ( .A(n19949), .B(n19948), .Z(n19947) );
  NOR U19944 ( .A(n22008), .B(n22009), .Z(n19948) );
  XOR U19945 ( .A(n19951), .B(n19950), .Z(n19949) );
  NOR U19946 ( .A(n22010), .B(n22011), .Z(n19950) );
  XOR U19947 ( .A(n19953), .B(n19952), .Z(n19951) );
  NOR U19948 ( .A(n22012), .B(n22013), .Z(n19952) );
  XOR U19949 ( .A(n19955), .B(n19954), .Z(n19953) );
  NOR U19950 ( .A(n22014), .B(n22015), .Z(n19954) );
  XOR U19951 ( .A(n19957), .B(n19956), .Z(n19955) );
  NOR U19952 ( .A(n22016), .B(n22017), .Z(n19956) );
  XOR U19953 ( .A(n19959), .B(n19958), .Z(n19957) );
  NOR U19954 ( .A(n22018), .B(n22019), .Z(n19958) );
  XOR U19955 ( .A(n19961), .B(n19960), .Z(n19959) );
  NOR U19956 ( .A(n22020), .B(n22021), .Z(n19960) );
  XOR U19957 ( .A(n19963), .B(n19962), .Z(n19961) );
  NOR U19958 ( .A(n22022), .B(n22023), .Z(n19962) );
  XOR U19959 ( .A(n19965), .B(n19964), .Z(n19963) );
  NOR U19960 ( .A(n22024), .B(n22025), .Z(n19964) );
  XOR U19961 ( .A(n19967), .B(n19966), .Z(n19965) );
  NOR U19962 ( .A(n22026), .B(n22027), .Z(n19966) );
  XOR U19963 ( .A(n19969), .B(n19968), .Z(n19967) );
  NOR U19964 ( .A(n22028), .B(n22029), .Z(n19968) );
  XOR U19965 ( .A(n19971), .B(n19970), .Z(n19969) );
  NOR U19966 ( .A(n22030), .B(n22031), .Z(n19970) );
  XOR U19967 ( .A(n19973), .B(n19972), .Z(n19971) );
  NOR U19968 ( .A(n22032), .B(n22033), .Z(n19972) );
  XOR U19969 ( .A(n19975), .B(n19974), .Z(n19973) );
  NOR U19970 ( .A(n22034), .B(n22035), .Z(n19974) );
  XOR U19971 ( .A(n19977), .B(n19976), .Z(n19975) );
  NOR U19972 ( .A(n22036), .B(n22037), .Z(n19976) );
  XOR U19973 ( .A(n19979), .B(n19978), .Z(n19977) );
  NOR U19974 ( .A(n22038), .B(n22039), .Z(n19978) );
  XOR U19975 ( .A(n19981), .B(n19980), .Z(n19979) );
  NOR U19976 ( .A(n22040), .B(n22041), .Z(n19980) );
  XOR U19977 ( .A(n19983), .B(n19982), .Z(n19981) );
  NOR U19978 ( .A(n22042), .B(n22043), .Z(n19982) );
  XOR U19979 ( .A(n19985), .B(n19984), .Z(n19983) );
  NOR U19980 ( .A(n22044), .B(n22045), .Z(n19984) );
  XOR U19981 ( .A(n19987), .B(n19986), .Z(n19985) );
  NOR U19982 ( .A(n22046), .B(n22047), .Z(n19986) );
  XOR U19983 ( .A(n19989), .B(n19988), .Z(n19987) );
  NOR U19984 ( .A(n22048), .B(n22049), .Z(n19988) );
  XOR U19985 ( .A(n19991), .B(n19990), .Z(n19989) );
  NOR U19986 ( .A(n22050), .B(n22051), .Z(n19990) );
  XOR U19987 ( .A(n19993), .B(n19992), .Z(n19991) );
  NOR U19988 ( .A(n22052), .B(n22053), .Z(n19992) );
  XOR U19989 ( .A(n19995), .B(n19994), .Z(n19993) );
  NOR U19990 ( .A(n22054), .B(n22055), .Z(n19994) );
  XOR U19991 ( .A(n19997), .B(n19996), .Z(n19995) );
  NOR U19992 ( .A(n22056), .B(n22057), .Z(n19996) );
  XOR U19993 ( .A(n19999), .B(n19998), .Z(n19997) );
  NOR U19994 ( .A(n22058), .B(n22059), .Z(n19998) );
  XOR U19995 ( .A(n20001), .B(n20000), .Z(n19999) );
  NOR U19996 ( .A(n22060), .B(n22061), .Z(n20000) );
  XOR U19997 ( .A(n20003), .B(n20002), .Z(n20001) );
  NOR U19998 ( .A(n22062), .B(n22063), .Z(n20002) );
  XOR U19999 ( .A(n20005), .B(n20004), .Z(n20003) );
  NOR U20000 ( .A(n22064), .B(n22065), .Z(n20004) );
  XOR U20001 ( .A(n20007), .B(n20006), .Z(n20005) );
  NOR U20002 ( .A(n22066), .B(n22067), .Z(n20006) );
  XOR U20003 ( .A(n20009), .B(n20008), .Z(n20007) );
  NOR U20004 ( .A(n22068), .B(n22069), .Z(n20008) );
  XOR U20005 ( .A(n20011), .B(n20010), .Z(n20009) );
  NOR U20006 ( .A(n22070), .B(n22071), .Z(n20010) );
  XOR U20007 ( .A(n20013), .B(n20012), .Z(n20011) );
  NOR U20008 ( .A(n22072), .B(n22073), .Z(n20012) );
  XOR U20009 ( .A(n20015), .B(n20014), .Z(n20013) );
  NOR U20010 ( .A(n22074), .B(n22075), .Z(n20014) );
  XOR U20011 ( .A(n20017), .B(n20016), .Z(n20015) );
  NOR U20012 ( .A(n22076), .B(n22077), .Z(n20016) );
  XOR U20013 ( .A(n20019), .B(n20018), .Z(n20017) );
  NOR U20014 ( .A(n22078), .B(n22079), .Z(n20018) );
  XOR U20015 ( .A(n20021), .B(n20020), .Z(n20019) );
  NOR U20016 ( .A(n22080), .B(n22081), .Z(n20020) );
  XOR U20017 ( .A(n20023), .B(n20022), .Z(n20021) );
  NOR U20018 ( .A(n22082), .B(n22083), .Z(n20022) );
  XOR U20019 ( .A(n20025), .B(n20024), .Z(n20023) );
  NOR U20020 ( .A(n22084), .B(n22085), .Z(n20024) );
  XOR U20021 ( .A(n20027), .B(n20026), .Z(n20025) );
  NOR U20022 ( .A(n22086), .B(n22087), .Z(n20026) );
  XOR U20023 ( .A(n20029), .B(n20028), .Z(n20027) );
  NOR U20024 ( .A(n22088), .B(n22089), .Z(n20028) );
  XOR U20025 ( .A(n20031), .B(n20030), .Z(n20029) );
  NOR U20026 ( .A(n22090), .B(n22091), .Z(n20030) );
  XOR U20027 ( .A(n20033), .B(n20032), .Z(n20031) );
  NOR U20028 ( .A(n22092), .B(n22093), .Z(n20032) );
  XOR U20029 ( .A(n20035), .B(n20034), .Z(n20033) );
  NOR U20030 ( .A(n22094), .B(n22095), .Z(n20034) );
  XOR U20031 ( .A(n20037), .B(n20036), .Z(n20035) );
  NOR U20032 ( .A(n22096), .B(n22097), .Z(n20036) );
  XOR U20033 ( .A(n20039), .B(n20038), .Z(n20037) );
  NOR U20034 ( .A(n22098), .B(n22099), .Z(n20038) );
  XOR U20035 ( .A(n20041), .B(n20040), .Z(n20039) );
  NOR U20036 ( .A(n22100), .B(n22101), .Z(n20040) );
  XOR U20037 ( .A(n20043), .B(n20042), .Z(n20041) );
  NOR U20038 ( .A(n22102), .B(n22103), .Z(n20042) );
  XOR U20039 ( .A(n20045), .B(n20044), .Z(n20043) );
  NOR U20040 ( .A(n22104), .B(n22105), .Z(n20044) );
  XOR U20041 ( .A(n20047), .B(n20046), .Z(n20045) );
  NOR U20042 ( .A(n22106), .B(n22107), .Z(n20046) );
  XOR U20043 ( .A(n20049), .B(n20048), .Z(n20047) );
  NOR U20044 ( .A(n22108), .B(n22109), .Z(n20048) );
  XOR U20045 ( .A(n20051), .B(n20050), .Z(n20049) );
  NOR U20046 ( .A(n22110), .B(n22111), .Z(n20050) );
  XOR U20047 ( .A(n20053), .B(n20052), .Z(n20051) );
  NOR U20048 ( .A(n22112), .B(n22113), .Z(n20052) );
  XOR U20049 ( .A(n20055), .B(n20054), .Z(n20053) );
  NOR U20050 ( .A(n22114), .B(n22115), .Z(n20054) );
  XOR U20051 ( .A(n20057), .B(n20056), .Z(n20055) );
  NOR U20052 ( .A(n22116), .B(n22117), .Z(n20056) );
  XOR U20053 ( .A(n20059), .B(n20058), .Z(n20057) );
  NOR U20054 ( .A(n22118), .B(n22119), .Z(n20058) );
  XOR U20055 ( .A(n20061), .B(n20060), .Z(n20059) );
  NOR U20056 ( .A(n22120), .B(n22121), .Z(n20060) );
  XOR U20057 ( .A(n20063), .B(n20062), .Z(n20061) );
  NOR U20058 ( .A(n22122), .B(n22123), .Z(n20062) );
  XOR U20059 ( .A(n20065), .B(n20064), .Z(n20063) );
  NOR U20060 ( .A(n22124), .B(n22125), .Z(n20064) );
  XOR U20061 ( .A(n20067), .B(n20066), .Z(n20065) );
  NOR U20062 ( .A(n22126), .B(n22127), .Z(n20066) );
  XOR U20063 ( .A(n20069), .B(n20068), .Z(n20067) );
  NOR U20064 ( .A(n22128), .B(n22129), .Z(n20068) );
  XOR U20065 ( .A(n20071), .B(n20070), .Z(n20069) );
  NOR U20066 ( .A(n22130), .B(n22131), .Z(n20070) );
  XOR U20067 ( .A(n20073), .B(n20072), .Z(n20071) );
  NOR U20068 ( .A(n22132), .B(n22133), .Z(n20072) );
  XOR U20069 ( .A(n20075), .B(n20074), .Z(n20073) );
  NOR U20070 ( .A(n22134), .B(n22135), .Z(n20074) );
  XOR U20071 ( .A(n20077), .B(n20076), .Z(n20075) );
  NOR U20072 ( .A(n22136), .B(n22137), .Z(n20076) );
  XOR U20073 ( .A(n20079), .B(n20078), .Z(n20077) );
  NOR U20074 ( .A(n22138), .B(n22139), .Z(n20078) );
  XOR U20075 ( .A(n20081), .B(n20080), .Z(n20079) );
  NOR U20076 ( .A(n22140), .B(n22141), .Z(n20080) );
  XOR U20077 ( .A(n20083), .B(n20082), .Z(n20081) );
  NOR U20078 ( .A(n22142), .B(n22143), .Z(n20082) );
  XOR U20079 ( .A(n20085), .B(n20084), .Z(n20083) );
  NOR U20080 ( .A(n22144), .B(n22145), .Z(n20084) );
  XOR U20081 ( .A(n20087), .B(n20086), .Z(n20085) );
  NOR U20082 ( .A(n22146), .B(n22147), .Z(n20086) );
  XOR U20083 ( .A(n20089), .B(n20088), .Z(n20087) );
  NOR U20084 ( .A(n22148), .B(n22149), .Z(n20088) );
  XOR U20085 ( .A(n20091), .B(n20090), .Z(n20089) );
  NOR U20086 ( .A(n22150), .B(n22151), .Z(n20090) );
  XOR U20087 ( .A(n20093), .B(n20092), .Z(n20091) );
  NOR U20088 ( .A(n22152), .B(n22153), .Z(n20092) );
  XOR U20089 ( .A(n20095), .B(n20094), .Z(n20093) );
  NOR U20090 ( .A(n22154), .B(n22155), .Z(n20094) );
  XOR U20091 ( .A(n20097), .B(n20096), .Z(n20095) );
  NOR U20092 ( .A(n22156), .B(n22157), .Z(n20096) );
  XOR U20093 ( .A(n20099), .B(n20098), .Z(n20097) );
  NOR U20094 ( .A(n22158), .B(n22159), .Z(n20098) );
  XOR U20095 ( .A(n20101), .B(n20100), .Z(n20099) );
  NOR U20096 ( .A(n22160), .B(n22161), .Z(n20100) );
  XOR U20097 ( .A(n20103), .B(n20102), .Z(n20101) );
  NOR U20098 ( .A(n22162), .B(n22163), .Z(n20102) );
  XOR U20099 ( .A(n20105), .B(n20104), .Z(n20103) );
  NOR U20100 ( .A(n22164), .B(n22165), .Z(n20104) );
  XOR U20101 ( .A(n20107), .B(n20106), .Z(n20105) );
  NOR U20102 ( .A(n22166), .B(n22167), .Z(n20106) );
  XOR U20103 ( .A(n20109), .B(n20108), .Z(n20107) );
  NOR U20104 ( .A(n22168), .B(n22169), .Z(n20108) );
  XOR U20105 ( .A(n20111), .B(n20110), .Z(n20109) );
  NOR U20106 ( .A(n22170), .B(n22171), .Z(n20110) );
  XOR U20107 ( .A(n20113), .B(n20112), .Z(n20111) );
  NOR U20108 ( .A(n22172), .B(n22173), .Z(n20112) );
  XOR U20109 ( .A(n20115), .B(n20114), .Z(n20113) );
  NOR U20110 ( .A(n22174), .B(n22175), .Z(n20114) );
  XOR U20111 ( .A(n20117), .B(n20116), .Z(n20115) );
  NOR U20112 ( .A(n22176), .B(n22177), .Z(n20116) );
  XOR U20113 ( .A(n20119), .B(n20118), .Z(n20117) );
  NOR U20114 ( .A(n22178), .B(n22179), .Z(n20118) );
  XOR U20115 ( .A(n20121), .B(n20120), .Z(n20119) );
  NOR U20116 ( .A(n22180), .B(n22181), .Z(n20120) );
  XOR U20117 ( .A(n20123), .B(n20122), .Z(n20121) );
  NOR U20118 ( .A(n22182), .B(n22183), .Z(n20122) );
  XOR U20119 ( .A(n20125), .B(n20124), .Z(n20123) );
  NOR U20120 ( .A(n22184), .B(n22185), .Z(n20124) );
  XOR U20121 ( .A(n20127), .B(n20126), .Z(n20125) );
  NOR U20122 ( .A(n22186), .B(n22187), .Z(n20126) );
  XOR U20123 ( .A(n20129), .B(n20128), .Z(n20127) );
  NOR U20124 ( .A(n22188), .B(n22189), .Z(n20128) );
  XOR U20125 ( .A(n20131), .B(n20130), .Z(n20129) );
  NOR U20126 ( .A(n22190), .B(n22191), .Z(n20130) );
  XOR U20127 ( .A(n20133), .B(n20132), .Z(n20131) );
  NOR U20128 ( .A(n22192), .B(n22193), .Z(n20132) );
  XOR U20129 ( .A(n20135), .B(n20134), .Z(n20133) );
  NOR U20130 ( .A(n22194), .B(n22195), .Z(n20134) );
  XOR U20131 ( .A(n20137), .B(n20136), .Z(n20135) );
  NOR U20132 ( .A(n22196), .B(n22197), .Z(n20136) );
  XOR U20133 ( .A(n20139), .B(n20138), .Z(n20137) );
  NOR U20134 ( .A(n22198), .B(n22199), .Z(n20138) );
  XOR U20135 ( .A(n20141), .B(n20140), .Z(n20139) );
  NOR U20136 ( .A(n22200), .B(n22201), .Z(n20140) );
  XOR U20137 ( .A(n20143), .B(n20142), .Z(n20141) );
  NOR U20138 ( .A(n22202), .B(n22203), .Z(n20142) );
  XOR U20139 ( .A(n20145), .B(n20144), .Z(n20143) );
  NOR U20140 ( .A(n22204), .B(n22205), .Z(n20144) );
  XOR U20141 ( .A(n20147), .B(n20146), .Z(n20145) );
  NOR U20142 ( .A(n22206), .B(n22207), .Z(n20146) );
  XOR U20143 ( .A(n20149), .B(n20148), .Z(n20147) );
  NOR U20144 ( .A(n22208), .B(n22209), .Z(n20148) );
  XOR U20145 ( .A(n20151), .B(n20150), .Z(n20149) );
  NOR U20146 ( .A(n22210), .B(n22211), .Z(n20150) );
  XOR U20147 ( .A(n20153), .B(n20152), .Z(n20151) );
  NOR U20148 ( .A(n22212), .B(n22213), .Z(n20152) );
  XOR U20149 ( .A(n20155), .B(n20154), .Z(n20153) );
  NOR U20150 ( .A(n22214), .B(n22215), .Z(n20154) );
  XOR U20151 ( .A(n20157), .B(n20156), .Z(n20155) );
  NOR U20152 ( .A(n22216), .B(n22217), .Z(n20156) );
  XOR U20153 ( .A(n20159), .B(n20158), .Z(n20157) );
  NOR U20154 ( .A(n22218), .B(n22219), .Z(n20158) );
  XOR U20155 ( .A(n20161), .B(n20160), .Z(n20159) );
  NOR U20156 ( .A(n22220), .B(n22221), .Z(n20160) );
  XOR U20157 ( .A(n20163), .B(n20162), .Z(n20161) );
  NOR U20158 ( .A(n22222), .B(n22223), .Z(n20162) );
  XOR U20159 ( .A(n20165), .B(n20164), .Z(n20163) );
  NOR U20160 ( .A(n22224), .B(n22225), .Z(n20164) );
  XOR U20161 ( .A(n20167), .B(n20166), .Z(n20165) );
  NOR U20162 ( .A(n22226), .B(n22227), .Z(n20166) );
  XOR U20163 ( .A(n20169), .B(n20168), .Z(n20167) );
  NOR U20164 ( .A(n22228), .B(n22229), .Z(n20168) );
  XOR U20165 ( .A(n20171), .B(n20170), .Z(n20169) );
  NOR U20166 ( .A(n22230), .B(n22231), .Z(n20170) );
  XOR U20167 ( .A(n20173), .B(n20172), .Z(n20171) );
  NOR U20168 ( .A(n22232), .B(n22233), .Z(n20172) );
  XOR U20169 ( .A(n20175), .B(n20174), .Z(n20173) );
  NOR U20170 ( .A(n22234), .B(n22235), .Z(n20174) );
  XOR U20171 ( .A(n20177), .B(n20176), .Z(n20175) );
  NOR U20172 ( .A(n22236), .B(n22237), .Z(n20176) );
  XOR U20173 ( .A(n20179), .B(n20178), .Z(n20177) );
  NOR U20174 ( .A(n22238), .B(n22239), .Z(n20178) );
  XOR U20175 ( .A(n20181), .B(n20180), .Z(n20179) );
  NOR U20176 ( .A(n22240), .B(n22241), .Z(n20180) );
  XOR U20177 ( .A(n20183), .B(n20182), .Z(n20181) );
  NOR U20178 ( .A(n22242), .B(n22243), .Z(n20182) );
  XOR U20179 ( .A(n20185), .B(n20184), .Z(n20183) );
  NOR U20180 ( .A(n22244), .B(n22245), .Z(n20184) );
  XOR U20181 ( .A(n20187), .B(n20186), .Z(n20185) );
  NOR U20182 ( .A(n22246), .B(n22247), .Z(n20186) );
  XOR U20183 ( .A(n20189), .B(n20188), .Z(n20187) );
  NOR U20184 ( .A(n22248), .B(n22249), .Z(n20188) );
  XOR U20185 ( .A(n20191), .B(n20190), .Z(n20189) );
  NOR U20186 ( .A(n22250), .B(n22251), .Z(n20190) );
  XOR U20187 ( .A(n20193), .B(n20192), .Z(n20191) );
  NOR U20188 ( .A(n22252), .B(n22253), .Z(n20192) );
  XOR U20189 ( .A(n20195), .B(n20194), .Z(n20193) );
  NOR U20190 ( .A(n22254), .B(n22255), .Z(n20194) );
  XOR U20191 ( .A(n20197), .B(n20196), .Z(n20195) );
  NOR U20192 ( .A(n22256), .B(n22257), .Z(n20196) );
  XOR U20193 ( .A(n20199), .B(n20198), .Z(n20197) );
  NOR U20194 ( .A(n22258), .B(n22259), .Z(n20198) );
  XOR U20195 ( .A(n20201), .B(n20200), .Z(n20199) );
  NOR U20196 ( .A(n22260), .B(n22261), .Z(n20200) );
  XOR U20197 ( .A(n20203), .B(n20202), .Z(n20201) );
  NOR U20198 ( .A(n22262), .B(n22263), .Z(n20202) );
  XOR U20199 ( .A(n20205), .B(n20204), .Z(n20203) );
  NOR U20200 ( .A(n22264), .B(n22265), .Z(n20204) );
  XOR U20201 ( .A(n20207), .B(n20206), .Z(n20205) );
  NOR U20202 ( .A(n22266), .B(n22267), .Z(n20206) );
  XOR U20203 ( .A(n20209), .B(n20208), .Z(n20207) );
  NOR U20204 ( .A(n22268), .B(n22269), .Z(n20208) );
  XOR U20205 ( .A(n20211), .B(n20210), .Z(n20209) );
  NOR U20206 ( .A(n22270), .B(n22271), .Z(n20210) );
  XOR U20207 ( .A(n20213), .B(n20212), .Z(n20211) );
  NOR U20208 ( .A(n22272), .B(n22273), .Z(n20212) );
  XOR U20209 ( .A(n20215), .B(n20214), .Z(n20213) );
  NOR U20210 ( .A(n22274), .B(n22275), .Z(n20214) );
  XOR U20211 ( .A(n20217), .B(n20216), .Z(n20215) );
  NOR U20212 ( .A(n22276), .B(n22277), .Z(n20216) );
  XOR U20213 ( .A(n20219), .B(n20218), .Z(n20217) );
  NOR U20214 ( .A(n22278), .B(n22279), .Z(n20218) );
  XOR U20215 ( .A(n20221), .B(n20220), .Z(n20219) );
  NOR U20216 ( .A(n22280), .B(n22281), .Z(n20220) );
  XOR U20217 ( .A(n20223), .B(n20222), .Z(n20221) );
  NOR U20218 ( .A(n22282), .B(n22283), .Z(n20222) );
  XOR U20219 ( .A(n20225), .B(n20224), .Z(n20223) );
  NOR U20220 ( .A(n22284), .B(n22285), .Z(n20224) );
  XOR U20221 ( .A(n20227), .B(n20226), .Z(n20225) );
  NOR U20222 ( .A(n22286), .B(n22287), .Z(n20226) );
  XOR U20223 ( .A(n20229), .B(n20228), .Z(n20227) );
  NOR U20224 ( .A(n22288), .B(n22289), .Z(n20228) );
  XOR U20225 ( .A(n20231), .B(n20230), .Z(n20229) );
  NOR U20226 ( .A(n22290), .B(n22291), .Z(n20230) );
  XOR U20227 ( .A(n20233), .B(n20232), .Z(n20231) );
  NOR U20228 ( .A(n22292), .B(n22293), .Z(n20232) );
  XOR U20229 ( .A(n20235), .B(n20234), .Z(n20233) );
  NOR U20230 ( .A(n22294), .B(n22295), .Z(n20234) );
  XOR U20231 ( .A(n20237), .B(n20236), .Z(n20235) );
  NOR U20232 ( .A(n22296), .B(n22297), .Z(n20236) );
  XOR U20233 ( .A(n20239), .B(n20238), .Z(n20237) );
  NOR U20234 ( .A(n22298), .B(n22299), .Z(n20238) );
  XOR U20235 ( .A(n20241), .B(n20240), .Z(n20239) );
  NOR U20236 ( .A(n22300), .B(n22301), .Z(n20240) );
  XOR U20237 ( .A(n20243), .B(n20242), .Z(n20241) );
  NOR U20238 ( .A(n22302), .B(n22303), .Z(n20242) );
  XOR U20239 ( .A(n20245), .B(n20244), .Z(n20243) );
  NOR U20240 ( .A(n22304), .B(n22305), .Z(n20244) );
  XOR U20241 ( .A(n20247), .B(n20246), .Z(n20245) );
  NOR U20242 ( .A(n22306), .B(n22307), .Z(n20246) );
  XOR U20243 ( .A(n20249), .B(n20248), .Z(n20247) );
  NOR U20244 ( .A(n22308), .B(n22309), .Z(n20248) );
  XOR U20245 ( .A(n20251), .B(n20250), .Z(n20249) );
  NOR U20246 ( .A(n22310), .B(n22311), .Z(n20250) );
  XOR U20247 ( .A(n20253), .B(n20252), .Z(n20251) );
  NOR U20248 ( .A(n22312), .B(n22313), .Z(n20252) );
  XOR U20249 ( .A(n20255), .B(n20254), .Z(n20253) );
  NOR U20250 ( .A(n22314), .B(n22315), .Z(n20254) );
  XOR U20251 ( .A(n20257), .B(n20256), .Z(n20255) );
  NOR U20252 ( .A(n22316), .B(n22317), .Z(n20256) );
  XOR U20253 ( .A(n20259), .B(n20258), .Z(n20257) );
  NOR U20254 ( .A(n22318), .B(n22319), .Z(n20258) );
  XOR U20255 ( .A(n20261), .B(n20260), .Z(n20259) );
  NOR U20256 ( .A(n22320), .B(n22321), .Z(n20260) );
  XOR U20257 ( .A(n20263), .B(n20262), .Z(n20261) );
  NOR U20258 ( .A(n22322), .B(n22323), .Z(n20262) );
  XOR U20259 ( .A(n20265), .B(n20264), .Z(n20263) );
  NOR U20260 ( .A(n22324), .B(n22325), .Z(n20264) );
  XOR U20261 ( .A(n20267), .B(n20266), .Z(n20265) );
  NOR U20262 ( .A(n22326), .B(n22327), .Z(n20266) );
  XOR U20263 ( .A(n20269), .B(n20268), .Z(n20267) );
  NOR U20264 ( .A(n22328), .B(n22329), .Z(n20268) );
  XOR U20265 ( .A(n20271), .B(n20270), .Z(n20269) );
  NOR U20266 ( .A(n22330), .B(n22331), .Z(n20270) );
  XOR U20267 ( .A(n20273), .B(n20272), .Z(n20271) );
  NOR U20268 ( .A(n22332), .B(n22333), .Z(n20272) );
  XOR U20269 ( .A(n20275), .B(n20274), .Z(n20273) );
  NOR U20270 ( .A(n22334), .B(n22335), .Z(n20274) );
  XOR U20271 ( .A(n20277), .B(n20276), .Z(n20275) );
  NOR U20272 ( .A(n22336), .B(n22337), .Z(n20276) );
  XOR U20273 ( .A(n20279), .B(n20278), .Z(n20277) );
  NOR U20274 ( .A(n22338), .B(n22339), .Z(n20278) );
  XOR U20275 ( .A(n20281), .B(n20280), .Z(n20279) );
  NOR U20276 ( .A(n22340), .B(n22341), .Z(n20280) );
  XOR U20277 ( .A(n20283), .B(n20282), .Z(n20281) );
  NOR U20278 ( .A(n22342), .B(n22343), .Z(n20282) );
  XOR U20279 ( .A(n20285), .B(n20284), .Z(n20283) );
  NOR U20280 ( .A(n22344), .B(n22345), .Z(n20284) );
  XOR U20281 ( .A(n20287), .B(n20286), .Z(n20285) );
  NOR U20282 ( .A(n22346), .B(n22347), .Z(n20286) );
  XOR U20283 ( .A(n20289), .B(n20288), .Z(n20287) );
  NOR U20284 ( .A(n22348), .B(n22349), .Z(n20288) );
  XOR U20285 ( .A(n20291), .B(n20290), .Z(n20289) );
  NOR U20286 ( .A(n22350), .B(n22351), .Z(n20290) );
  XOR U20287 ( .A(n20293), .B(n20292), .Z(n20291) );
  NOR U20288 ( .A(n22352), .B(n22353), .Z(n20292) );
  XOR U20289 ( .A(n20295), .B(n20294), .Z(n20293) );
  NOR U20290 ( .A(n22354), .B(n22355), .Z(n20294) );
  XOR U20291 ( .A(n20297), .B(n20296), .Z(n20295) );
  NOR U20292 ( .A(n22356), .B(n22357), .Z(n20296) );
  XOR U20293 ( .A(n20299), .B(n20298), .Z(n20297) );
  NOR U20294 ( .A(n22358), .B(n22359), .Z(n20298) );
  XOR U20295 ( .A(n20301), .B(n20300), .Z(n20299) );
  NOR U20296 ( .A(n22360), .B(n22361), .Z(n20300) );
  XOR U20297 ( .A(n20303), .B(n20302), .Z(n20301) );
  NOR U20298 ( .A(n22362), .B(n22363), .Z(n20302) );
  XOR U20299 ( .A(n20305), .B(n20304), .Z(n20303) );
  NOR U20300 ( .A(n22364), .B(n22365), .Z(n20304) );
  XOR U20301 ( .A(n20307), .B(n20306), .Z(n20305) );
  NOR U20302 ( .A(n22366), .B(n22367), .Z(n20306) );
  XOR U20303 ( .A(n20309), .B(n20308), .Z(n20307) );
  NOR U20304 ( .A(n22368), .B(n22369), .Z(n20308) );
  XOR U20305 ( .A(n20311), .B(n20310), .Z(n20309) );
  NOR U20306 ( .A(n22370), .B(n22371), .Z(n20310) );
  XOR U20307 ( .A(n20313), .B(n20312), .Z(n20311) );
  NOR U20308 ( .A(n22372), .B(n22373), .Z(n20312) );
  XOR U20309 ( .A(n20315), .B(n20314), .Z(n20313) );
  NOR U20310 ( .A(n22374), .B(n22375), .Z(n20314) );
  XOR U20311 ( .A(n20317), .B(n20316), .Z(n20315) );
  NOR U20312 ( .A(n22376), .B(n22377), .Z(n20316) );
  XOR U20313 ( .A(n20319), .B(n20318), .Z(n20317) );
  NOR U20314 ( .A(n22378), .B(n22379), .Z(n20318) );
  XOR U20315 ( .A(n20321), .B(n20320), .Z(n20319) );
  NOR U20316 ( .A(n22380), .B(n22381), .Z(n20320) );
  XOR U20317 ( .A(n20323), .B(n20322), .Z(n20321) );
  NOR U20318 ( .A(n22382), .B(n22383), .Z(n20322) );
  XOR U20319 ( .A(n20325), .B(n20324), .Z(n20323) );
  NOR U20320 ( .A(n22384), .B(n22385), .Z(n20324) );
  XOR U20321 ( .A(n20327), .B(n20326), .Z(n20325) );
  NOR U20322 ( .A(n22386), .B(n22387), .Z(n20326) );
  XOR U20323 ( .A(n20329), .B(n20328), .Z(n20327) );
  NOR U20324 ( .A(n22388), .B(n22389), .Z(n20328) );
  XOR U20325 ( .A(n20331), .B(n20330), .Z(n20329) );
  NOR U20326 ( .A(n22390), .B(n22391), .Z(n20330) );
  XOR U20327 ( .A(n20333), .B(n20332), .Z(n20331) );
  NOR U20328 ( .A(n22392), .B(n22393), .Z(n20332) );
  XOR U20329 ( .A(n20335), .B(n20334), .Z(n20333) );
  NOR U20330 ( .A(n22394), .B(n22395), .Z(n20334) );
  XOR U20331 ( .A(n20337), .B(n20336), .Z(n20335) );
  NOR U20332 ( .A(n22396), .B(n22397), .Z(n20336) );
  XOR U20333 ( .A(n20339), .B(n20338), .Z(n20337) );
  NOR U20334 ( .A(n22398), .B(n22399), .Z(n20338) );
  XOR U20335 ( .A(n20341), .B(n20340), .Z(n20339) );
  NOR U20336 ( .A(n22400), .B(n22401), .Z(n20340) );
  XOR U20337 ( .A(n20343), .B(n20342), .Z(n20341) );
  NOR U20338 ( .A(n22402), .B(n22403), .Z(n20342) );
  XOR U20339 ( .A(n20345), .B(n20344), .Z(n20343) );
  NOR U20340 ( .A(n22404), .B(n22405), .Z(n20344) );
  XOR U20341 ( .A(n20347), .B(n20346), .Z(n20345) );
  NOR U20342 ( .A(n22406), .B(n22407), .Z(n20346) );
  XOR U20343 ( .A(n20349), .B(n20348), .Z(n20347) );
  NOR U20344 ( .A(n22408), .B(n22409), .Z(n20348) );
  XOR U20345 ( .A(n20351), .B(n20350), .Z(n20349) );
  NOR U20346 ( .A(n22410), .B(n22411), .Z(n20350) );
  XOR U20347 ( .A(n20353), .B(n20352), .Z(n20351) );
  NOR U20348 ( .A(n22412), .B(n22413), .Z(n20352) );
  XOR U20349 ( .A(n20355), .B(n20354), .Z(n20353) );
  NOR U20350 ( .A(n22414), .B(n22415), .Z(n20354) );
  XOR U20351 ( .A(n20357), .B(n20356), .Z(n20355) );
  NOR U20352 ( .A(n22416), .B(n22417), .Z(n20356) );
  XOR U20353 ( .A(n20359), .B(n20358), .Z(n20357) );
  NOR U20354 ( .A(n22418), .B(n22419), .Z(n20358) );
  XOR U20355 ( .A(n20361), .B(n20360), .Z(n20359) );
  NOR U20356 ( .A(n22420), .B(n22421), .Z(n20360) );
  XOR U20357 ( .A(n20363), .B(n20362), .Z(n20361) );
  NOR U20358 ( .A(n22422), .B(n22423), .Z(n20362) );
  XOR U20359 ( .A(n20365), .B(n20364), .Z(n20363) );
  NOR U20360 ( .A(n22424), .B(n22425), .Z(n20364) );
  XOR U20361 ( .A(n20367), .B(n20366), .Z(n20365) );
  NOR U20362 ( .A(n22426), .B(n22427), .Z(n20366) );
  XOR U20363 ( .A(n20369), .B(n20368), .Z(n20367) );
  NOR U20364 ( .A(n22428), .B(n22429), .Z(n20368) );
  XOR U20365 ( .A(n20371), .B(n20370), .Z(n20369) );
  NOR U20366 ( .A(n22430), .B(n22431), .Z(n20370) );
  XOR U20367 ( .A(n20373), .B(n20372), .Z(n20371) );
  NOR U20368 ( .A(n22432), .B(n22433), .Z(n20372) );
  XOR U20369 ( .A(n20375), .B(n20374), .Z(n20373) );
  NOR U20370 ( .A(n22434), .B(n22435), .Z(n20374) );
  XOR U20371 ( .A(n20377), .B(n20376), .Z(n20375) );
  NOR U20372 ( .A(n22436), .B(n22437), .Z(n20376) );
  XOR U20373 ( .A(n20379), .B(n20378), .Z(n20377) );
  NOR U20374 ( .A(n22438), .B(n22439), .Z(n20378) );
  XOR U20375 ( .A(n20381), .B(n20380), .Z(n20379) );
  NOR U20376 ( .A(n22440), .B(n22441), .Z(n20380) );
  XOR U20377 ( .A(n20383), .B(n20382), .Z(n20381) );
  NOR U20378 ( .A(n22442), .B(n22443), .Z(n20382) );
  XOR U20379 ( .A(n20385), .B(n20384), .Z(n20383) );
  NOR U20380 ( .A(n22444), .B(n22445), .Z(n20384) );
  XOR U20381 ( .A(n20387), .B(n20386), .Z(n20385) );
  NOR U20382 ( .A(n22446), .B(n22447), .Z(n20386) );
  XOR U20383 ( .A(n20389), .B(n20388), .Z(n20387) );
  NOR U20384 ( .A(n22448), .B(n22449), .Z(n20388) );
  XOR U20385 ( .A(n20391), .B(n20390), .Z(n20389) );
  NOR U20386 ( .A(n22450), .B(n22451), .Z(n20390) );
  XOR U20387 ( .A(n20393), .B(n20392), .Z(n20391) );
  NOR U20388 ( .A(n22452), .B(n22453), .Z(n20392) );
  XOR U20389 ( .A(n20395), .B(n20394), .Z(n20393) );
  NOR U20390 ( .A(n22454), .B(n22455), .Z(n20394) );
  XOR U20391 ( .A(n20397), .B(n20396), .Z(n20395) );
  NOR U20392 ( .A(n22456), .B(n22457), .Z(n20396) );
  XOR U20393 ( .A(n20399), .B(n20398), .Z(n20397) );
  NOR U20394 ( .A(n22458), .B(n22459), .Z(n20398) );
  XOR U20395 ( .A(n20401), .B(n20400), .Z(n20399) );
  NOR U20396 ( .A(n22460), .B(n22461), .Z(n20400) );
  XOR U20397 ( .A(n20403), .B(n20402), .Z(n20401) );
  NOR U20398 ( .A(n22462), .B(n22463), .Z(n20402) );
  XOR U20399 ( .A(n20405), .B(n20404), .Z(n20403) );
  NOR U20400 ( .A(n22464), .B(n22465), .Z(n20404) );
  XOR U20401 ( .A(n20407), .B(n20406), .Z(n20405) );
  NOR U20402 ( .A(n22466), .B(n22467), .Z(n20406) );
  XOR U20403 ( .A(n20409), .B(n20408), .Z(n20407) );
  NOR U20404 ( .A(n22468), .B(n22469), .Z(n20408) );
  XOR U20405 ( .A(n20411), .B(n20410), .Z(n20409) );
  NOR U20406 ( .A(n22470), .B(n22471), .Z(n20410) );
  XOR U20407 ( .A(n20413), .B(n20412), .Z(n20411) );
  NOR U20408 ( .A(n22472), .B(n22473), .Z(n20412) );
  XOR U20409 ( .A(n20415), .B(n20414), .Z(n20413) );
  NOR U20410 ( .A(n22474), .B(n22475), .Z(n20414) );
  XOR U20411 ( .A(n20417), .B(n20416), .Z(n20415) );
  NOR U20412 ( .A(n22476), .B(n22477), .Z(n20416) );
  XOR U20413 ( .A(n20419), .B(n20418), .Z(n20417) );
  NOR U20414 ( .A(n22478), .B(n22479), .Z(n20418) );
  XOR U20415 ( .A(n20421), .B(n20420), .Z(n20419) );
  NOR U20416 ( .A(n22480), .B(n22481), .Z(n20420) );
  XOR U20417 ( .A(n20423), .B(n20422), .Z(n20421) );
  NOR U20418 ( .A(n22482), .B(n22483), .Z(n20422) );
  XOR U20419 ( .A(n20425), .B(n20424), .Z(n20423) );
  NOR U20420 ( .A(n22484), .B(n22485), .Z(n20424) );
  XOR U20421 ( .A(n20427), .B(n20426), .Z(n20425) );
  NOR U20422 ( .A(n22486), .B(n22487), .Z(n20426) );
  XOR U20423 ( .A(n20429), .B(n20428), .Z(n20427) );
  NOR U20424 ( .A(n22488), .B(n22489), .Z(n20428) );
  XOR U20425 ( .A(n20431), .B(n20430), .Z(n20429) );
  NOR U20426 ( .A(n22490), .B(n22491), .Z(n20430) );
  XOR U20427 ( .A(n20433), .B(n20432), .Z(n20431) );
  NOR U20428 ( .A(n22492), .B(n22493), .Z(n20432) );
  XOR U20429 ( .A(n20435), .B(n20434), .Z(n20433) );
  NOR U20430 ( .A(n22494), .B(n22495), .Z(n20434) );
  XOR U20431 ( .A(n20437), .B(n20436), .Z(n20435) );
  NOR U20432 ( .A(n22496), .B(n22497), .Z(n20436) );
  XOR U20433 ( .A(n20439), .B(n20438), .Z(n20437) );
  NOR U20434 ( .A(n22498), .B(n22499), .Z(n20438) );
  XOR U20435 ( .A(n20441), .B(n20440), .Z(n20439) );
  NOR U20436 ( .A(n22500), .B(n22501), .Z(n20440) );
  XOR U20437 ( .A(n20443), .B(n20442), .Z(n20441) );
  NOR U20438 ( .A(n22502), .B(n22503), .Z(n20442) );
  XOR U20439 ( .A(n20445), .B(n20444), .Z(n20443) );
  NOR U20440 ( .A(n22504), .B(n22505), .Z(n20444) );
  XOR U20441 ( .A(n20447), .B(n20446), .Z(n20445) );
  NOR U20442 ( .A(n22506), .B(n22507), .Z(n20446) );
  XOR U20443 ( .A(n20449), .B(n20448), .Z(n20447) );
  NOR U20444 ( .A(n22508), .B(n22509), .Z(n20448) );
  XOR U20445 ( .A(n20451), .B(n20450), .Z(n20449) );
  NOR U20446 ( .A(n22510), .B(n22511), .Z(n20450) );
  XOR U20447 ( .A(n20453), .B(n20452), .Z(n20451) );
  NOR U20448 ( .A(n22512), .B(n22513), .Z(n20452) );
  XOR U20449 ( .A(n20455), .B(n20454), .Z(n20453) );
  NOR U20450 ( .A(n22514), .B(n22515), .Z(n20454) );
  XOR U20451 ( .A(n20457), .B(n20456), .Z(n20455) );
  NOR U20452 ( .A(n22516), .B(n22517), .Z(n20456) );
  XOR U20453 ( .A(n20459), .B(n20458), .Z(n20457) );
  NOR U20454 ( .A(n22518), .B(n22519), .Z(n20458) );
  XOR U20455 ( .A(n20461), .B(n20460), .Z(n20459) );
  NOR U20456 ( .A(n22520), .B(n22521), .Z(n20460) );
  XOR U20457 ( .A(n20463), .B(n20462), .Z(n20461) );
  NOR U20458 ( .A(n22522), .B(n22523), .Z(n20462) );
  XOR U20459 ( .A(n20465), .B(n20464), .Z(n20463) );
  NOR U20460 ( .A(n22524), .B(n22525), .Z(n20464) );
  XOR U20461 ( .A(n20467), .B(n20466), .Z(n20465) );
  NOR U20462 ( .A(n22526), .B(n22527), .Z(n20466) );
  XOR U20463 ( .A(n20469), .B(n20468), .Z(n20467) );
  NOR U20464 ( .A(n22528), .B(n22529), .Z(n20468) );
  XOR U20465 ( .A(n20471), .B(n20470), .Z(n20469) );
  NOR U20466 ( .A(n22530), .B(n22531), .Z(n20470) );
  XOR U20467 ( .A(n20473), .B(n20472), .Z(n20471) );
  NOR U20468 ( .A(n22532), .B(n22533), .Z(n20472) );
  XOR U20469 ( .A(n20475), .B(n20474), .Z(n20473) );
  NOR U20470 ( .A(n22534), .B(n22535), .Z(n20474) );
  XOR U20471 ( .A(n20477), .B(n20476), .Z(n20475) );
  NOR U20472 ( .A(n22536), .B(n22537), .Z(n20476) );
  XOR U20473 ( .A(n20479), .B(n20478), .Z(n20477) );
  NOR U20474 ( .A(n22538), .B(n22539), .Z(n20478) );
  XOR U20475 ( .A(n20481), .B(n20480), .Z(n20479) );
  NOR U20476 ( .A(n22540), .B(n22541), .Z(n20480) );
  XOR U20477 ( .A(n20483), .B(n20482), .Z(n20481) );
  NOR U20478 ( .A(n22542), .B(n22543), .Z(n20482) );
  XOR U20479 ( .A(n20485), .B(n20484), .Z(n20483) );
  NOR U20480 ( .A(n22544), .B(n22545), .Z(n20484) );
  XOR U20481 ( .A(n20487), .B(n20486), .Z(n20485) );
  NOR U20482 ( .A(n22546), .B(n22547), .Z(n20486) );
  XOR U20483 ( .A(n20489), .B(n20488), .Z(n20487) );
  NOR U20484 ( .A(n22548), .B(n22549), .Z(n20488) );
  XOR U20485 ( .A(n20491), .B(n20490), .Z(n20489) );
  NOR U20486 ( .A(n22550), .B(n22551), .Z(n20490) );
  XOR U20487 ( .A(n20493), .B(n20492), .Z(n20491) );
  NOR U20488 ( .A(n22552), .B(n22553), .Z(n20492) );
  XOR U20489 ( .A(n20495), .B(n20494), .Z(n20493) );
  NOR U20490 ( .A(n22554), .B(n22555), .Z(n20494) );
  XOR U20491 ( .A(n20497), .B(n20496), .Z(n20495) );
  NOR U20492 ( .A(n22556), .B(n22557), .Z(n20496) );
  XOR U20493 ( .A(n20499), .B(n20498), .Z(n20497) );
  NOR U20494 ( .A(n22558), .B(n22559), .Z(n20498) );
  XOR U20495 ( .A(n20501), .B(n20500), .Z(n20499) );
  NOR U20496 ( .A(n22560), .B(n22561), .Z(n20500) );
  XOR U20497 ( .A(n20503), .B(n20502), .Z(n20501) );
  NOR U20498 ( .A(n22562), .B(n22563), .Z(n20502) );
  XOR U20499 ( .A(n20505), .B(n20504), .Z(n20503) );
  NOR U20500 ( .A(n22564), .B(n22565), .Z(n20504) );
  XOR U20501 ( .A(n20507), .B(n20506), .Z(n20505) );
  NOR U20502 ( .A(n22566), .B(n22567), .Z(n20506) );
  XOR U20503 ( .A(n20509), .B(n20508), .Z(n20507) );
  NOR U20504 ( .A(n22568), .B(n22569), .Z(n20508) );
  XOR U20505 ( .A(n20511), .B(n20510), .Z(n20509) );
  NOR U20506 ( .A(n22570), .B(n22571), .Z(n20510) );
  XOR U20507 ( .A(n20513), .B(n20512), .Z(n20511) );
  NOR U20508 ( .A(n22572), .B(n22573), .Z(n20512) );
  XOR U20509 ( .A(n20515), .B(n20514), .Z(n20513) );
  NOR U20510 ( .A(n22574), .B(n22575), .Z(n20514) );
  XOR U20511 ( .A(n20517), .B(n20516), .Z(n20515) );
  NOR U20512 ( .A(n22576), .B(n22577), .Z(n20516) );
  XOR U20513 ( .A(n20519), .B(n20518), .Z(n20517) );
  NOR U20514 ( .A(n22578), .B(n22579), .Z(n20518) );
  XOR U20515 ( .A(n20521), .B(n20520), .Z(n20519) );
  NOR U20516 ( .A(n22580), .B(n22581), .Z(n20520) );
  XOR U20517 ( .A(n20523), .B(n20522), .Z(n20521) );
  NOR U20518 ( .A(n22582), .B(n22583), .Z(n20522) );
  XOR U20519 ( .A(n20525), .B(n20524), .Z(n20523) );
  NOR U20520 ( .A(n22584), .B(n22585), .Z(n20524) );
  XOR U20521 ( .A(n20527), .B(n20526), .Z(n20525) );
  NOR U20522 ( .A(n22586), .B(n22587), .Z(n20526) );
  XOR U20523 ( .A(n20529), .B(n20528), .Z(n20527) );
  NOR U20524 ( .A(n22588), .B(n22589), .Z(n20528) );
  XOR U20525 ( .A(n20531), .B(n20530), .Z(n20529) );
  NOR U20526 ( .A(n22590), .B(n22591), .Z(n20530) );
  XOR U20527 ( .A(n20533), .B(n20532), .Z(n20531) );
  NOR U20528 ( .A(n22592), .B(n22593), .Z(n20532) );
  XOR U20529 ( .A(n20535), .B(n20534), .Z(n20533) );
  NOR U20530 ( .A(n22594), .B(n22595), .Z(n20534) );
  XOR U20531 ( .A(n20537), .B(n20536), .Z(n20535) );
  NOR U20532 ( .A(n22596), .B(n22597), .Z(n20536) );
  XOR U20533 ( .A(n20539), .B(n20538), .Z(n20537) );
  NOR U20534 ( .A(n22598), .B(n22599), .Z(n20538) );
  XOR U20535 ( .A(n20541), .B(n20540), .Z(n20539) );
  NOR U20536 ( .A(n22600), .B(n22601), .Z(n20540) );
  XOR U20537 ( .A(n20543), .B(n20542), .Z(n20541) );
  NOR U20538 ( .A(n22602), .B(n22603), .Z(n20542) );
  XOR U20539 ( .A(n20545), .B(n20544), .Z(n20543) );
  NOR U20540 ( .A(n22604), .B(n22605), .Z(n20544) );
  XOR U20541 ( .A(n20547), .B(n20546), .Z(n20545) );
  NOR U20542 ( .A(n22606), .B(n22607), .Z(n20546) );
  XOR U20543 ( .A(n20549), .B(n20548), .Z(n20547) );
  NOR U20544 ( .A(n22608), .B(n22609), .Z(n20548) );
  XOR U20545 ( .A(n20551), .B(n20550), .Z(n20549) );
  NOR U20546 ( .A(n22610), .B(n22611), .Z(n20550) );
  XOR U20547 ( .A(n20553), .B(n20552), .Z(n20551) );
  NOR U20548 ( .A(n22612), .B(n22613), .Z(n20552) );
  XOR U20549 ( .A(n20555), .B(n20554), .Z(n20553) );
  NOR U20550 ( .A(n22614), .B(n22615), .Z(n20554) );
  XOR U20551 ( .A(n20557), .B(n20556), .Z(n20555) );
  NOR U20552 ( .A(n22616), .B(n22617), .Z(n20556) );
  XOR U20553 ( .A(n20559), .B(n20558), .Z(n20557) );
  NOR U20554 ( .A(n22618), .B(n22619), .Z(n20558) );
  XOR U20555 ( .A(n20561), .B(n20560), .Z(n20559) );
  NOR U20556 ( .A(n22620), .B(n22621), .Z(n20560) );
  XOR U20557 ( .A(n20563), .B(n20562), .Z(n20561) );
  NOR U20558 ( .A(n22622), .B(n22623), .Z(n20562) );
  XOR U20559 ( .A(n20565), .B(n20564), .Z(n20563) );
  NOR U20560 ( .A(n22624), .B(n22625), .Z(n20564) );
  XOR U20561 ( .A(n20567), .B(n20566), .Z(n20565) );
  NOR U20562 ( .A(n22626), .B(n22627), .Z(n20566) );
  XOR U20563 ( .A(n20569), .B(n20568), .Z(n20567) );
  NOR U20564 ( .A(n22628), .B(n22629), .Z(n20568) );
  XOR U20565 ( .A(n20571), .B(n20570), .Z(n20569) );
  NOR U20566 ( .A(n22630), .B(n22631), .Z(n20570) );
  XOR U20567 ( .A(n20573), .B(n20572), .Z(n20571) );
  NOR U20568 ( .A(n22632), .B(n22633), .Z(n20572) );
  XOR U20569 ( .A(n20575), .B(n20574), .Z(n20573) );
  NOR U20570 ( .A(n22634), .B(n22635), .Z(n20574) );
  XOR U20571 ( .A(n20577), .B(n20576), .Z(n20575) );
  NOR U20572 ( .A(n22636), .B(n22637), .Z(n20576) );
  XOR U20573 ( .A(n20579), .B(n20578), .Z(n20577) );
  NOR U20574 ( .A(n22638), .B(n22639), .Z(n20578) );
  XOR U20575 ( .A(n20581), .B(n20580), .Z(n20579) );
  NOR U20576 ( .A(n22640), .B(n22641), .Z(n20580) );
  XOR U20577 ( .A(n20583), .B(n20582), .Z(n20581) );
  NOR U20578 ( .A(n22642), .B(n22643), .Z(n20582) );
  XOR U20579 ( .A(n20585), .B(n20584), .Z(n20583) );
  NOR U20580 ( .A(n22644), .B(n22645), .Z(n20584) );
  XOR U20581 ( .A(n20587), .B(n20586), .Z(n20585) );
  NOR U20582 ( .A(n22646), .B(n22647), .Z(n20586) );
  XOR U20583 ( .A(n20589), .B(n20588), .Z(n20587) );
  NOR U20584 ( .A(n22648), .B(n22649), .Z(n20588) );
  XOR U20585 ( .A(n20591), .B(n20590), .Z(n20589) );
  NOR U20586 ( .A(n22650), .B(n22651), .Z(n20590) );
  XOR U20587 ( .A(n20593), .B(n20592), .Z(n20591) );
  NOR U20588 ( .A(n22652), .B(n22653), .Z(n20592) );
  XOR U20589 ( .A(n20595), .B(n20594), .Z(n20593) );
  NOR U20590 ( .A(n22654), .B(n22655), .Z(n20594) );
  XOR U20591 ( .A(n20597), .B(n20596), .Z(n20595) );
  NOR U20592 ( .A(n22656), .B(n22657), .Z(n20596) );
  XOR U20593 ( .A(n20599), .B(n20598), .Z(n20597) );
  NOR U20594 ( .A(n22658), .B(n22659), .Z(n20598) );
  XOR U20595 ( .A(n20601), .B(n20600), .Z(n20599) );
  NOR U20596 ( .A(n22660), .B(n22661), .Z(n20600) );
  XOR U20597 ( .A(n20603), .B(n20602), .Z(n20601) );
  NOR U20598 ( .A(n22662), .B(n22663), .Z(n20602) );
  XOR U20599 ( .A(n20605), .B(n20604), .Z(n20603) );
  NOR U20600 ( .A(n22664), .B(n22665), .Z(n20604) );
  XOR U20601 ( .A(n20607), .B(n20606), .Z(n20605) );
  NOR U20602 ( .A(n22666), .B(n22667), .Z(n20606) );
  XOR U20603 ( .A(n20609), .B(n20608), .Z(n20607) );
  NOR U20604 ( .A(n22668), .B(n22669), .Z(n20608) );
  XOR U20605 ( .A(n20611), .B(n20610), .Z(n20609) );
  NOR U20606 ( .A(n22670), .B(n22671), .Z(n20610) );
  XOR U20607 ( .A(n20613), .B(n20612), .Z(n20611) );
  NOR U20608 ( .A(n22672), .B(n22673), .Z(n20612) );
  XOR U20609 ( .A(n20615), .B(n20614), .Z(n20613) );
  NOR U20610 ( .A(n22674), .B(n22675), .Z(n20614) );
  XOR U20611 ( .A(n20617), .B(n20616), .Z(n20615) );
  NOR U20612 ( .A(n22676), .B(n22677), .Z(n20616) );
  XOR U20613 ( .A(n20619), .B(n20618), .Z(n20617) );
  NOR U20614 ( .A(n22678), .B(n22679), .Z(n20618) );
  XOR U20615 ( .A(n20621), .B(n20620), .Z(n20619) );
  NOR U20616 ( .A(n22680), .B(n22681), .Z(n20620) );
  XOR U20617 ( .A(n20623), .B(n20622), .Z(n20621) );
  NOR U20618 ( .A(n22682), .B(n22683), .Z(n20622) );
  XOR U20619 ( .A(n20625), .B(n20624), .Z(n20623) );
  NOR U20620 ( .A(n22684), .B(n22685), .Z(n20624) );
  XOR U20621 ( .A(n20627), .B(n20626), .Z(n20625) );
  NOR U20622 ( .A(n22686), .B(n22687), .Z(n20626) );
  XOR U20623 ( .A(n20631), .B(n20630), .Z(n20627) );
  NOR U20624 ( .A(n22688), .B(n22689), .Z(n20630) );
  XOR U20625 ( .A(n20633), .B(n20632), .Z(n20631) );
  NOR U20626 ( .A(n22690), .B(n22691), .Z(n20632) );
  XOR U20627 ( .A(n20635), .B(n20634), .Z(n20633) );
  NOR U20628 ( .A(n22692), .B(n22693), .Z(n20634) );
  XOR U20629 ( .A(n20637), .B(n20636), .Z(n20635) );
  NOR U20630 ( .A(n22694), .B(n22695), .Z(n20636) );
  XOR U20631 ( .A(n20639), .B(n20638), .Z(n20637) );
  NOR U20632 ( .A(n22696), .B(n22697), .Z(n20638) );
  XOR U20633 ( .A(n20641), .B(n20640), .Z(n20639) );
  NOR U20634 ( .A(n22698), .B(n22699), .Z(n20640) );
  XOR U20635 ( .A(n20643), .B(n20642), .Z(n20641) );
  NOR U20636 ( .A(n22700), .B(n22701), .Z(n20642) );
  XOR U20637 ( .A(n20645), .B(n20644), .Z(n20643) );
  NOR U20638 ( .A(n22702), .B(n22703), .Z(n20644) );
  XOR U20639 ( .A(n20647), .B(n20646), .Z(n20645) );
  NOR U20640 ( .A(n22704), .B(n22705), .Z(n20646) );
  XOR U20641 ( .A(n20649), .B(n20648), .Z(n20647) );
  NOR U20642 ( .A(n22706), .B(n22707), .Z(n20648) );
  XOR U20643 ( .A(n20651), .B(n20650), .Z(n20649) );
  NOR U20644 ( .A(n22708), .B(n22709), .Z(n20650) );
  XOR U20645 ( .A(n20653), .B(n20652), .Z(n20651) );
  NOR U20646 ( .A(n22710), .B(n22711), .Z(n20652) );
  XOR U20647 ( .A(n20655), .B(n20654), .Z(n20653) );
  NOR U20648 ( .A(n22712), .B(n22713), .Z(n20654) );
  XOR U20649 ( .A(n20657), .B(n20656), .Z(n20655) );
  NOR U20650 ( .A(n22714), .B(n22715), .Z(n20656) );
  XOR U20651 ( .A(n20659), .B(n20658), .Z(n20657) );
  NOR U20652 ( .A(n22716), .B(n22717), .Z(n20658) );
  XOR U20653 ( .A(n20661), .B(n20660), .Z(n20659) );
  NOR U20654 ( .A(n22718), .B(n22719), .Z(n20660) );
  XOR U20655 ( .A(n20663), .B(n20662), .Z(n20661) );
  NOR U20656 ( .A(n22720), .B(n22721), .Z(n20662) );
  XOR U20657 ( .A(n20665), .B(n20664), .Z(n20663) );
  NOR U20658 ( .A(n22722), .B(n22723), .Z(n20664) );
  XOR U20659 ( .A(n20667), .B(n20666), .Z(n20665) );
  NOR U20660 ( .A(n22724), .B(n22725), .Z(n20666) );
  XOR U20661 ( .A(n20669), .B(n20668), .Z(n20667) );
  NOR U20662 ( .A(n22726), .B(n22727), .Z(n20668) );
  XOR U20663 ( .A(n20671), .B(n20670), .Z(n20669) );
  NOR U20664 ( .A(n22728), .B(n22729), .Z(n20670) );
  XOR U20665 ( .A(n20673), .B(n20672), .Z(n20671) );
  NOR U20666 ( .A(n22730), .B(n22731), .Z(n20672) );
  XOR U20667 ( .A(n20675), .B(n20674), .Z(n20673) );
  NOR U20668 ( .A(n22732), .B(n22733), .Z(n20674) );
  XOR U20669 ( .A(n20677), .B(n20676), .Z(n20675) );
  NOR U20670 ( .A(n22734), .B(n22735), .Z(n20676) );
  XOR U20671 ( .A(n20679), .B(n20678), .Z(n20677) );
  NOR U20672 ( .A(n22736), .B(n22737), .Z(n20678) );
  XOR U20673 ( .A(n20681), .B(n20680), .Z(n20679) );
  NOR U20674 ( .A(n22738), .B(n22739), .Z(n20680) );
  XOR U20675 ( .A(n20683), .B(n20682), .Z(n20681) );
  NOR U20676 ( .A(n22740), .B(n22741), .Z(n20682) );
  XOR U20677 ( .A(n20685), .B(n20684), .Z(n20683) );
  NOR U20678 ( .A(n22742), .B(n22743), .Z(n20684) );
  XOR U20679 ( .A(n20687), .B(n20686), .Z(n20685) );
  NOR U20680 ( .A(n22744), .B(n22745), .Z(n20686) );
  XOR U20681 ( .A(n20689), .B(n20688), .Z(n20687) );
  NOR U20682 ( .A(n22746), .B(n22747), .Z(n20688) );
  XOR U20683 ( .A(n20691), .B(n20690), .Z(n20689) );
  NOR U20684 ( .A(n22748), .B(n22749), .Z(n20690) );
  XOR U20685 ( .A(n20693), .B(n20692), .Z(n20691) );
  NOR U20686 ( .A(n22750), .B(n22751), .Z(n20692) );
  XOR U20687 ( .A(n20695), .B(n20694), .Z(n20693) );
  NOR U20688 ( .A(n22752), .B(n22753), .Z(n20694) );
  XOR U20689 ( .A(n20697), .B(n20696), .Z(n20695) );
  NOR U20690 ( .A(n22754), .B(n22755), .Z(n20696) );
  XOR U20691 ( .A(n20699), .B(n20698), .Z(n20697) );
  NOR U20692 ( .A(n22756), .B(n22757), .Z(n20698) );
  XOR U20693 ( .A(n20701), .B(n20700), .Z(n20699) );
  NOR U20694 ( .A(n22758), .B(n22759), .Z(n20700) );
  XOR U20695 ( .A(n20703), .B(n20702), .Z(n20701) );
  NOR U20696 ( .A(n22760), .B(n22761), .Z(n20702) );
  XOR U20697 ( .A(n20705), .B(n20704), .Z(n20703) );
  NOR U20698 ( .A(n22762), .B(n22763), .Z(n20704) );
  XOR U20699 ( .A(n20707), .B(n20706), .Z(n20705) );
  NOR U20700 ( .A(n22764), .B(n22765), .Z(n20706) );
  XOR U20701 ( .A(n20709), .B(n20708), .Z(n20707) );
  NOR U20702 ( .A(n22766), .B(n22767), .Z(n20708) );
  XOR U20703 ( .A(n20711), .B(n20710), .Z(n20709) );
  NOR U20704 ( .A(n22768), .B(n22769), .Z(n20710) );
  XOR U20705 ( .A(n20713), .B(n20712), .Z(n20711) );
  NOR U20706 ( .A(n22770), .B(n22771), .Z(n20712) );
  XOR U20707 ( .A(n20715), .B(n20714), .Z(n20713) );
  NOR U20708 ( .A(n22772), .B(n22773), .Z(n20714) );
  XOR U20709 ( .A(n20717), .B(n20716), .Z(n20715) );
  NOR U20710 ( .A(n22774), .B(n22775), .Z(n20716) );
  XOR U20711 ( .A(n20719), .B(n20718), .Z(n20717) );
  NOR U20712 ( .A(n22776), .B(n22777), .Z(n20718) );
  XOR U20713 ( .A(n20721), .B(n20720), .Z(n20719) );
  NOR U20714 ( .A(n22778), .B(n22779), .Z(n20720) );
  XOR U20715 ( .A(n20723), .B(n20722), .Z(n20721) );
  NOR U20716 ( .A(n22780), .B(n22781), .Z(n20722) );
  XOR U20717 ( .A(n20725), .B(n20724), .Z(n20723) );
  NOR U20718 ( .A(n22782), .B(n22783), .Z(n20724) );
  XOR U20719 ( .A(n20727), .B(n20726), .Z(n20725) );
  NOR U20720 ( .A(n22784), .B(n22785), .Z(n20726) );
  XOR U20721 ( .A(n20729), .B(n20728), .Z(n20727) );
  NOR U20722 ( .A(n22786), .B(n22787), .Z(n20728) );
  XOR U20723 ( .A(n20731), .B(n20730), .Z(n20729) );
  NOR U20724 ( .A(n22788), .B(n22789), .Z(n20730) );
  XOR U20725 ( .A(n20733), .B(n20732), .Z(n20731) );
  NOR U20726 ( .A(n22790), .B(n22791), .Z(n20732) );
  XOR U20727 ( .A(n20735), .B(n20734), .Z(n20733) );
  NOR U20728 ( .A(n22792), .B(n22793), .Z(n20734) );
  XOR U20729 ( .A(n20737), .B(n20736), .Z(n20735) );
  NOR U20730 ( .A(n22794), .B(n22795), .Z(n20736) );
  XOR U20731 ( .A(n20739), .B(n20738), .Z(n20737) );
  NOR U20732 ( .A(n22796), .B(n22797), .Z(n20738) );
  XOR U20733 ( .A(n20741), .B(n20740), .Z(n20739) );
  NOR U20734 ( .A(n22798), .B(n22799), .Z(n20740) );
  XOR U20735 ( .A(n20743), .B(n20742), .Z(n20741) );
  NOR U20736 ( .A(n22800), .B(n22801), .Z(n20742) );
  XOR U20737 ( .A(n20745), .B(n20744), .Z(n20743) );
  NOR U20738 ( .A(n22802), .B(n22803), .Z(n20744) );
  XOR U20739 ( .A(n20747), .B(n20746), .Z(n20745) );
  NOR U20740 ( .A(n22804), .B(n22805), .Z(n20746) );
  XOR U20741 ( .A(n20749), .B(n20748), .Z(n20747) );
  NOR U20742 ( .A(n22806), .B(n22807), .Z(n20748) );
  XOR U20743 ( .A(n20751), .B(n20750), .Z(n20749) );
  NOR U20744 ( .A(n22808), .B(n22809), .Z(n20750) );
  XOR U20745 ( .A(n20753), .B(n20752), .Z(n20751) );
  NOR U20746 ( .A(n22810), .B(n22811), .Z(n20752) );
  XOR U20747 ( .A(n20755), .B(n20754), .Z(n20753) );
  NOR U20748 ( .A(n22812), .B(n22813), .Z(n20754) );
  XOR U20749 ( .A(n20757), .B(n20756), .Z(n20755) );
  NOR U20750 ( .A(n22814), .B(n22815), .Z(n20756) );
  XOR U20751 ( .A(n20759), .B(n20758), .Z(n20757) );
  NOR U20752 ( .A(n22816), .B(n22817), .Z(n20758) );
  XOR U20753 ( .A(n20761), .B(n20760), .Z(n20759) );
  NOR U20754 ( .A(n22818), .B(n22819), .Z(n20760) );
  XOR U20755 ( .A(n20763), .B(n20762), .Z(n20761) );
  NOR U20756 ( .A(n22820), .B(n22821), .Z(n20762) );
  XOR U20757 ( .A(n20765), .B(n20764), .Z(n20763) );
  NOR U20758 ( .A(n22822), .B(n22823), .Z(n20764) );
  XOR U20759 ( .A(n20767), .B(n20766), .Z(n20765) );
  NOR U20760 ( .A(n22824), .B(n22825), .Z(n20766) );
  XOR U20761 ( .A(n20769), .B(n20768), .Z(n20767) );
  NOR U20762 ( .A(n22826), .B(n22827), .Z(n20768) );
  XOR U20763 ( .A(n20771), .B(n20770), .Z(n20769) );
  NOR U20764 ( .A(n22828), .B(n22829), .Z(n20770) );
  XOR U20765 ( .A(n20773), .B(n20772), .Z(n20771) );
  NOR U20766 ( .A(n22830), .B(n22831), .Z(n20772) );
  XOR U20767 ( .A(n20775), .B(n20774), .Z(n20773) );
  NOR U20768 ( .A(n22832), .B(n22833), .Z(n20774) );
  XOR U20769 ( .A(n20777), .B(n20776), .Z(n20775) );
  NOR U20770 ( .A(n22834), .B(n22835), .Z(n20776) );
  XOR U20771 ( .A(n20779), .B(n20778), .Z(n20777) );
  NOR U20772 ( .A(n22836), .B(n22837), .Z(n20778) );
  XOR U20773 ( .A(n20781), .B(n20780), .Z(n20779) );
  NOR U20774 ( .A(n22838), .B(n22839), .Z(n20780) );
  XOR U20775 ( .A(n20783), .B(n20782), .Z(n20781) );
  NOR U20776 ( .A(n22840), .B(n22841), .Z(n20782) );
  XOR U20777 ( .A(n20785), .B(n20784), .Z(n20783) );
  NOR U20778 ( .A(n22842), .B(n22843), .Z(n20784) );
  XOR U20779 ( .A(n20787), .B(n20786), .Z(n20785) );
  NOR U20780 ( .A(n22844), .B(n22845), .Z(n20786) );
  XOR U20781 ( .A(n20789), .B(n20788), .Z(n20787) );
  NOR U20782 ( .A(n22846), .B(n22847), .Z(n20788) );
  XOR U20783 ( .A(n20791), .B(n20790), .Z(n20789) );
  NOR U20784 ( .A(n22848), .B(n22849), .Z(n20790) );
  XOR U20785 ( .A(n20793), .B(n20792), .Z(n20791) );
  NOR U20786 ( .A(n22850), .B(n22851), .Z(n20792) );
  XOR U20787 ( .A(n20795), .B(n20794), .Z(n20793) );
  NOR U20788 ( .A(n22852), .B(n22853), .Z(n20794) );
  XOR U20789 ( .A(n20797), .B(n20796), .Z(n20795) );
  NOR U20790 ( .A(n22854), .B(n22855), .Z(n20796) );
  XOR U20791 ( .A(n20799), .B(n20798), .Z(n20797) );
  NOR U20792 ( .A(n22856), .B(n22857), .Z(n20798) );
  XOR U20793 ( .A(n20801), .B(n20800), .Z(n20799) );
  NOR U20794 ( .A(n22858), .B(n22859), .Z(n20800) );
  XOR U20795 ( .A(n20803), .B(n20802), .Z(n20801) );
  NOR U20796 ( .A(n22860), .B(n22861), .Z(n20802) );
  XOR U20797 ( .A(n20805), .B(n20804), .Z(n20803) );
  NOR U20798 ( .A(n22862), .B(n22863), .Z(n20804) );
  XOR U20799 ( .A(n20807), .B(n20806), .Z(n20805) );
  NOR U20800 ( .A(n22864), .B(n22865), .Z(n20806) );
  XOR U20801 ( .A(n20809), .B(n20808), .Z(n20807) );
  NOR U20802 ( .A(n22866), .B(n22867), .Z(n20808) );
  XOR U20803 ( .A(n20811), .B(n20810), .Z(n20809) );
  NOR U20804 ( .A(n22868), .B(n22869), .Z(n20810) );
  XOR U20805 ( .A(n20813), .B(n20812), .Z(n20811) );
  NOR U20806 ( .A(n22870), .B(n22871), .Z(n20812) );
  XOR U20807 ( .A(n20815), .B(n20814), .Z(n20813) );
  NOR U20808 ( .A(n22872), .B(n22873), .Z(n20814) );
  XOR U20809 ( .A(n20817), .B(n20816), .Z(n20815) );
  NOR U20810 ( .A(n22874), .B(n22875), .Z(n20816) );
  XOR U20811 ( .A(n20819), .B(n20818), .Z(n20817) );
  NOR U20812 ( .A(n22876), .B(n22877), .Z(n20818) );
  XOR U20813 ( .A(n20821), .B(n20820), .Z(n20819) );
  NOR U20814 ( .A(n22878), .B(n22879), .Z(n20820) );
  XOR U20815 ( .A(n20823), .B(n20822), .Z(n20821) );
  NOR U20816 ( .A(n22880), .B(n22881), .Z(n20822) );
  XOR U20817 ( .A(n20825), .B(n20824), .Z(n20823) );
  NOR U20818 ( .A(n22882), .B(n22883), .Z(n20824) );
  XOR U20819 ( .A(n20827), .B(n20826), .Z(n20825) );
  NOR U20820 ( .A(n22884), .B(n22885), .Z(n20826) );
  XOR U20821 ( .A(n20829), .B(n20828), .Z(n20827) );
  NOR U20822 ( .A(n22886), .B(n22887), .Z(n20828) );
  XOR U20823 ( .A(n20831), .B(n20830), .Z(n20829) );
  NOR U20824 ( .A(n22888), .B(n22889), .Z(n20830) );
  XOR U20825 ( .A(n20833), .B(n20832), .Z(n20831) );
  NOR U20826 ( .A(n22890), .B(n22891), .Z(n20832) );
  XOR U20827 ( .A(n20835), .B(n20834), .Z(n20833) );
  NOR U20828 ( .A(n22892), .B(n22893), .Z(n20834) );
  XOR U20829 ( .A(n20837), .B(n20836), .Z(n20835) );
  NOR U20830 ( .A(n22894), .B(n22895), .Z(n20836) );
  XOR U20831 ( .A(n20839), .B(n20838), .Z(n20837) );
  NOR U20832 ( .A(n22896), .B(n22897), .Z(n20838) );
  XOR U20833 ( .A(n20841), .B(n20840), .Z(n20839) );
  NOR U20834 ( .A(n22898), .B(n22899), .Z(n20840) );
  XOR U20835 ( .A(n20843), .B(n20842), .Z(n20841) );
  NOR U20836 ( .A(n22900), .B(n22901), .Z(n20842) );
  XOR U20837 ( .A(n20845), .B(n20844), .Z(n20843) );
  NOR U20838 ( .A(n22902), .B(n22903), .Z(n20844) );
  XOR U20839 ( .A(n20847), .B(n20846), .Z(n20845) );
  NOR U20840 ( .A(n22904), .B(n22905), .Z(n20846) );
  XOR U20841 ( .A(n20849), .B(n20848), .Z(n20847) );
  NOR U20842 ( .A(n22906), .B(n22907), .Z(n20848) );
  XOR U20843 ( .A(n20851), .B(n20850), .Z(n20849) );
  NOR U20844 ( .A(n22908), .B(n22909), .Z(n20850) );
  XOR U20845 ( .A(n20853), .B(n20852), .Z(n20851) );
  NOR U20846 ( .A(n22910), .B(n22911), .Z(n20852) );
  XOR U20847 ( .A(n20855), .B(n20854), .Z(n20853) );
  NOR U20848 ( .A(n22912), .B(n22913), .Z(n20854) );
  XOR U20849 ( .A(n20857), .B(n20856), .Z(n20855) );
  NOR U20850 ( .A(n22914), .B(n22915), .Z(n20856) );
  XOR U20851 ( .A(n20859), .B(n20858), .Z(n20857) );
  NOR U20852 ( .A(n22916), .B(n22917), .Z(n20858) );
  XOR U20853 ( .A(n20861), .B(n20860), .Z(n20859) );
  NOR U20854 ( .A(n22918), .B(n22919), .Z(n20860) );
  XOR U20855 ( .A(n20863), .B(n20862), .Z(n20861) );
  NOR U20856 ( .A(n22920), .B(n22921), .Z(n20862) );
  XOR U20857 ( .A(n20865), .B(n20864), .Z(n20863) );
  NOR U20858 ( .A(n22922), .B(n22923), .Z(n20864) );
  XOR U20859 ( .A(n20867), .B(n20866), .Z(n20865) );
  NOR U20860 ( .A(n22924), .B(n22925), .Z(n20866) );
  XOR U20861 ( .A(n20869), .B(n20868), .Z(n20867) );
  NOR U20862 ( .A(n22926), .B(n22927), .Z(n20868) );
  XOR U20863 ( .A(n20871), .B(n20870), .Z(n20869) );
  NOR U20864 ( .A(n22928), .B(n22929), .Z(n20870) );
  XOR U20865 ( .A(n20885), .B(n20884), .Z(n20871) );
  NOR U20866 ( .A(n22930), .B(n22931), .Z(n20884) );
  XOR U20867 ( .A(n20887), .B(n20886), .Z(n20885) );
  NOR U20868 ( .A(n22932), .B(n22933), .Z(n20886) );
  XOR U20869 ( .A(n20875), .B(n20874), .Z(n20887) );
  NOR U20870 ( .A(n22934), .B(n22935), .Z(n20874) );
  XOR U20871 ( .A(n20882), .B(n20883), .Z(n20875) );
  XOR U20872 ( .A(n20880), .B(n20881), .Z(n20883) );
  NOR U20873 ( .A(n22936), .B(n22937), .Z(n20881) );
  NOR U20874 ( .A(n22938), .B(n22939), .Z(n20880) );
  NOR U20875 ( .A(n22940), .B(n22941), .Z(n20882) );
  XNOR U20876 ( .A(n20889), .B(n20888), .Z(n143) );
  NOR U20877 ( .A(n21918), .B(p_input[1022]), .Z(n20888) );
  XOR U20878 ( .A(n20891), .B(n20890), .Z(n20889) );
  NOR U20879 ( .A(n21920), .B(p_input[1020]), .Z(n20890) );
  XOR U20880 ( .A(n20893), .B(n20892), .Z(n20891) );
  NOR U20881 ( .A(n21922), .B(p_input[1018]), .Z(n20892) );
  XOR U20882 ( .A(n20895), .B(n20894), .Z(n20893) );
  NOR U20883 ( .A(n21924), .B(p_input[1016]), .Z(n20894) );
  XOR U20884 ( .A(n20897), .B(n20896), .Z(n20895) );
  NOR U20885 ( .A(n21926), .B(p_input[1014]), .Z(n20896) );
  XOR U20886 ( .A(n20899), .B(n20898), .Z(n20897) );
  NOR U20887 ( .A(n21928), .B(p_input[1012]), .Z(n20898) );
  XOR U20888 ( .A(n20901), .B(n20900), .Z(n20899) );
  NOR U20889 ( .A(n21930), .B(p_input[1010]), .Z(n20900) );
  XOR U20890 ( .A(n20903), .B(n20902), .Z(n20901) );
  NOR U20891 ( .A(n21932), .B(p_input[1008]), .Z(n20902) );
  XOR U20892 ( .A(n20905), .B(n20904), .Z(n20903) );
  NOR U20893 ( .A(n21934), .B(p_input[1006]), .Z(n20904) );
  XOR U20894 ( .A(n20907), .B(n20906), .Z(n20905) );
  NOR U20895 ( .A(n21936), .B(p_input[1004]), .Z(n20906) );
  XOR U20896 ( .A(n20909), .B(n20908), .Z(n20907) );
  NOR U20897 ( .A(n21938), .B(p_input[1002]), .Z(n20908) );
  XOR U20898 ( .A(n20911), .B(n20910), .Z(n20909) );
  NOR U20899 ( .A(n21940), .B(p_input[1000]), .Z(n20910) );
  XOR U20900 ( .A(n20913), .B(n20912), .Z(n20911) );
  NOR U20901 ( .A(n21942), .B(p_input[998]), .Z(n20912) );
  XOR U20902 ( .A(n20915), .B(n20914), .Z(n20913) );
  NOR U20903 ( .A(n21944), .B(p_input[996]), .Z(n20914) );
  XOR U20904 ( .A(n20917), .B(n20916), .Z(n20915) );
  NOR U20905 ( .A(n21946), .B(p_input[994]), .Z(n20916) );
  XOR U20906 ( .A(n20919), .B(n20918), .Z(n20917) );
  NOR U20907 ( .A(n21948), .B(p_input[992]), .Z(n20918) );
  XOR U20908 ( .A(n20921), .B(n20920), .Z(n20919) );
  NOR U20909 ( .A(n21950), .B(p_input[990]), .Z(n20920) );
  XOR U20910 ( .A(n20923), .B(n20922), .Z(n20921) );
  NOR U20911 ( .A(n21952), .B(p_input[988]), .Z(n20922) );
  XOR U20912 ( .A(n20925), .B(n20924), .Z(n20923) );
  NOR U20913 ( .A(n21954), .B(p_input[986]), .Z(n20924) );
  XOR U20914 ( .A(n20927), .B(n20926), .Z(n20925) );
  NOR U20915 ( .A(n21956), .B(p_input[984]), .Z(n20926) );
  XOR U20916 ( .A(n20929), .B(n20928), .Z(n20927) );
  NOR U20917 ( .A(n21958), .B(p_input[982]), .Z(n20928) );
  XOR U20918 ( .A(n20931), .B(n20930), .Z(n20929) );
  NOR U20919 ( .A(n21960), .B(p_input[980]), .Z(n20930) );
  XOR U20920 ( .A(n20933), .B(n20932), .Z(n20931) );
  NOR U20921 ( .A(n21962), .B(p_input[978]), .Z(n20932) );
  XOR U20922 ( .A(n20935), .B(n20934), .Z(n20933) );
  NOR U20923 ( .A(n21964), .B(p_input[976]), .Z(n20934) );
  XOR U20924 ( .A(n20937), .B(n20936), .Z(n20935) );
  NOR U20925 ( .A(n21966), .B(p_input[974]), .Z(n20936) );
  XOR U20926 ( .A(n20939), .B(n20938), .Z(n20937) );
  NOR U20927 ( .A(n21968), .B(p_input[972]), .Z(n20938) );
  XOR U20928 ( .A(n20941), .B(n20940), .Z(n20939) );
  NOR U20929 ( .A(n21970), .B(p_input[970]), .Z(n20940) );
  XOR U20930 ( .A(n20943), .B(n20942), .Z(n20941) );
  NOR U20931 ( .A(n21972), .B(p_input[968]), .Z(n20942) );
  XOR U20932 ( .A(n20945), .B(n20944), .Z(n20943) );
  NOR U20933 ( .A(n21974), .B(p_input[966]), .Z(n20944) );
  XOR U20934 ( .A(n20947), .B(n20946), .Z(n20945) );
  NOR U20935 ( .A(n21976), .B(p_input[964]), .Z(n20946) );
  XOR U20936 ( .A(n20949), .B(n20948), .Z(n20947) );
  NOR U20937 ( .A(n21978), .B(p_input[962]), .Z(n20948) );
  XOR U20938 ( .A(n20951), .B(n20950), .Z(n20949) );
  NOR U20939 ( .A(n21980), .B(p_input[960]), .Z(n20950) );
  XOR U20940 ( .A(n20953), .B(n20952), .Z(n20951) );
  NOR U20941 ( .A(n21982), .B(p_input[958]), .Z(n20952) );
  XOR U20942 ( .A(n20955), .B(n20954), .Z(n20953) );
  NOR U20943 ( .A(n21984), .B(p_input[956]), .Z(n20954) );
  XOR U20944 ( .A(n20957), .B(n20956), .Z(n20955) );
  NOR U20945 ( .A(n21986), .B(p_input[954]), .Z(n20956) );
  XOR U20946 ( .A(n20959), .B(n20958), .Z(n20957) );
  NOR U20947 ( .A(n21988), .B(p_input[952]), .Z(n20958) );
  XOR U20948 ( .A(n20961), .B(n20960), .Z(n20959) );
  NOR U20949 ( .A(n21990), .B(p_input[950]), .Z(n20960) );
  XOR U20950 ( .A(n20963), .B(n20962), .Z(n20961) );
  NOR U20951 ( .A(n21992), .B(p_input[948]), .Z(n20962) );
  XOR U20952 ( .A(n20965), .B(n20964), .Z(n20963) );
  NOR U20953 ( .A(n21994), .B(p_input[946]), .Z(n20964) );
  XOR U20954 ( .A(n20967), .B(n20966), .Z(n20965) );
  NOR U20955 ( .A(n21996), .B(p_input[944]), .Z(n20966) );
  XOR U20956 ( .A(n20969), .B(n20968), .Z(n20967) );
  NOR U20957 ( .A(n21998), .B(p_input[942]), .Z(n20968) );
  XOR U20958 ( .A(n20971), .B(n20970), .Z(n20969) );
  NOR U20959 ( .A(n22000), .B(p_input[940]), .Z(n20970) );
  XOR U20960 ( .A(n20973), .B(n20972), .Z(n20971) );
  NOR U20961 ( .A(n22002), .B(p_input[938]), .Z(n20972) );
  XOR U20962 ( .A(n20975), .B(n20974), .Z(n20973) );
  NOR U20963 ( .A(n22004), .B(p_input[936]), .Z(n20974) );
  XOR U20964 ( .A(n20977), .B(n20976), .Z(n20975) );
  NOR U20965 ( .A(n22006), .B(p_input[934]), .Z(n20976) );
  XOR U20966 ( .A(n20979), .B(n20978), .Z(n20977) );
  NOR U20967 ( .A(n22008), .B(p_input[932]), .Z(n20978) );
  XOR U20968 ( .A(n20981), .B(n20980), .Z(n20979) );
  NOR U20969 ( .A(n22010), .B(p_input[930]), .Z(n20980) );
  XOR U20970 ( .A(n20983), .B(n20982), .Z(n20981) );
  NOR U20971 ( .A(n22012), .B(p_input[928]), .Z(n20982) );
  XOR U20972 ( .A(n20985), .B(n20984), .Z(n20983) );
  NOR U20973 ( .A(n22014), .B(p_input[926]), .Z(n20984) );
  XOR U20974 ( .A(n20987), .B(n20986), .Z(n20985) );
  NOR U20975 ( .A(n22016), .B(p_input[924]), .Z(n20986) );
  XOR U20976 ( .A(n20989), .B(n20988), .Z(n20987) );
  NOR U20977 ( .A(n22018), .B(p_input[922]), .Z(n20988) );
  XOR U20978 ( .A(n20991), .B(n20990), .Z(n20989) );
  NOR U20979 ( .A(n22020), .B(p_input[920]), .Z(n20990) );
  XOR U20980 ( .A(n20993), .B(n20992), .Z(n20991) );
  NOR U20981 ( .A(n22022), .B(p_input[918]), .Z(n20992) );
  XOR U20982 ( .A(n20995), .B(n20994), .Z(n20993) );
  NOR U20983 ( .A(n22024), .B(p_input[916]), .Z(n20994) );
  XOR U20984 ( .A(n20997), .B(n20996), .Z(n20995) );
  NOR U20985 ( .A(n22026), .B(p_input[914]), .Z(n20996) );
  XOR U20986 ( .A(n20999), .B(n20998), .Z(n20997) );
  NOR U20987 ( .A(n22028), .B(p_input[912]), .Z(n20998) );
  XOR U20988 ( .A(n21001), .B(n21000), .Z(n20999) );
  NOR U20989 ( .A(n22030), .B(p_input[910]), .Z(n21000) );
  XOR U20990 ( .A(n21003), .B(n21002), .Z(n21001) );
  NOR U20991 ( .A(n22032), .B(p_input[908]), .Z(n21002) );
  XOR U20992 ( .A(n21005), .B(n21004), .Z(n21003) );
  NOR U20993 ( .A(n22034), .B(p_input[906]), .Z(n21004) );
  XOR U20994 ( .A(n21007), .B(n21006), .Z(n21005) );
  NOR U20995 ( .A(n22036), .B(p_input[904]), .Z(n21006) );
  XOR U20996 ( .A(n21009), .B(n21008), .Z(n21007) );
  NOR U20997 ( .A(n22038), .B(p_input[902]), .Z(n21008) );
  XOR U20998 ( .A(n21011), .B(n21010), .Z(n21009) );
  NOR U20999 ( .A(n22040), .B(p_input[900]), .Z(n21010) );
  XOR U21000 ( .A(n21013), .B(n21012), .Z(n21011) );
  NOR U21001 ( .A(n22042), .B(p_input[898]), .Z(n21012) );
  XOR U21002 ( .A(n21015), .B(n21014), .Z(n21013) );
  NOR U21003 ( .A(n22044), .B(p_input[896]), .Z(n21014) );
  XOR U21004 ( .A(n21017), .B(n21016), .Z(n21015) );
  NOR U21005 ( .A(n22046), .B(p_input[894]), .Z(n21016) );
  XOR U21006 ( .A(n21019), .B(n21018), .Z(n21017) );
  NOR U21007 ( .A(n22048), .B(p_input[892]), .Z(n21018) );
  XOR U21008 ( .A(n21021), .B(n21020), .Z(n21019) );
  NOR U21009 ( .A(n22050), .B(p_input[890]), .Z(n21020) );
  XOR U21010 ( .A(n21023), .B(n21022), .Z(n21021) );
  NOR U21011 ( .A(n22052), .B(p_input[888]), .Z(n21022) );
  XOR U21012 ( .A(n21025), .B(n21024), .Z(n21023) );
  NOR U21013 ( .A(n22054), .B(p_input[886]), .Z(n21024) );
  XOR U21014 ( .A(n21027), .B(n21026), .Z(n21025) );
  NOR U21015 ( .A(n22056), .B(p_input[884]), .Z(n21026) );
  XOR U21016 ( .A(n21029), .B(n21028), .Z(n21027) );
  NOR U21017 ( .A(n22058), .B(p_input[882]), .Z(n21028) );
  XOR U21018 ( .A(n21031), .B(n21030), .Z(n21029) );
  NOR U21019 ( .A(n22060), .B(p_input[880]), .Z(n21030) );
  XOR U21020 ( .A(n21033), .B(n21032), .Z(n21031) );
  NOR U21021 ( .A(n22062), .B(p_input[878]), .Z(n21032) );
  XOR U21022 ( .A(n21035), .B(n21034), .Z(n21033) );
  NOR U21023 ( .A(n22064), .B(p_input[876]), .Z(n21034) );
  XOR U21024 ( .A(n21037), .B(n21036), .Z(n21035) );
  NOR U21025 ( .A(n22066), .B(p_input[874]), .Z(n21036) );
  XOR U21026 ( .A(n21039), .B(n21038), .Z(n21037) );
  NOR U21027 ( .A(n22068), .B(p_input[872]), .Z(n21038) );
  XOR U21028 ( .A(n21041), .B(n21040), .Z(n21039) );
  NOR U21029 ( .A(n22070), .B(p_input[870]), .Z(n21040) );
  XOR U21030 ( .A(n21043), .B(n21042), .Z(n21041) );
  NOR U21031 ( .A(n22072), .B(p_input[868]), .Z(n21042) );
  XOR U21032 ( .A(n21045), .B(n21044), .Z(n21043) );
  NOR U21033 ( .A(n22074), .B(p_input[866]), .Z(n21044) );
  XOR U21034 ( .A(n21047), .B(n21046), .Z(n21045) );
  NOR U21035 ( .A(n22076), .B(p_input[864]), .Z(n21046) );
  XOR U21036 ( .A(n21049), .B(n21048), .Z(n21047) );
  NOR U21037 ( .A(n22078), .B(p_input[862]), .Z(n21048) );
  XOR U21038 ( .A(n21051), .B(n21050), .Z(n21049) );
  NOR U21039 ( .A(n22080), .B(p_input[860]), .Z(n21050) );
  XOR U21040 ( .A(n21053), .B(n21052), .Z(n21051) );
  NOR U21041 ( .A(n22082), .B(p_input[858]), .Z(n21052) );
  XOR U21042 ( .A(n21055), .B(n21054), .Z(n21053) );
  NOR U21043 ( .A(n22084), .B(p_input[856]), .Z(n21054) );
  XOR U21044 ( .A(n21057), .B(n21056), .Z(n21055) );
  NOR U21045 ( .A(n22086), .B(p_input[854]), .Z(n21056) );
  XOR U21046 ( .A(n21059), .B(n21058), .Z(n21057) );
  NOR U21047 ( .A(n22088), .B(p_input[852]), .Z(n21058) );
  XOR U21048 ( .A(n21061), .B(n21060), .Z(n21059) );
  NOR U21049 ( .A(n22090), .B(p_input[850]), .Z(n21060) );
  XOR U21050 ( .A(n21063), .B(n21062), .Z(n21061) );
  NOR U21051 ( .A(n22092), .B(p_input[848]), .Z(n21062) );
  XOR U21052 ( .A(n21065), .B(n21064), .Z(n21063) );
  NOR U21053 ( .A(n22094), .B(p_input[846]), .Z(n21064) );
  XOR U21054 ( .A(n21067), .B(n21066), .Z(n21065) );
  NOR U21055 ( .A(n22096), .B(p_input[844]), .Z(n21066) );
  XOR U21056 ( .A(n21069), .B(n21068), .Z(n21067) );
  NOR U21057 ( .A(n22098), .B(p_input[842]), .Z(n21068) );
  XOR U21058 ( .A(n21071), .B(n21070), .Z(n21069) );
  NOR U21059 ( .A(n22100), .B(p_input[840]), .Z(n21070) );
  XOR U21060 ( .A(n21073), .B(n21072), .Z(n21071) );
  NOR U21061 ( .A(n22102), .B(p_input[838]), .Z(n21072) );
  XOR U21062 ( .A(n21075), .B(n21074), .Z(n21073) );
  NOR U21063 ( .A(n22104), .B(p_input[836]), .Z(n21074) );
  XOR U21064 ( .A(n21077), .B(n21076), .Z(n21075) );
  NOR U21065 ( .A(n22106), .B(p_input[834]), .Z(n21076) );
  XOR U21066 ( .A(n21079), .B(n21078), .Z(n21077) );
  NOR U21067 ( .A(n22108), .B(p_input[832]), .Z(n21078) );
  XOR U21068 ( .A(n21081), .B(n21080), .Z(n21079) );
  NOR U21069 ( .A(n22110), .B(p_input[830]), .Z(n21080) );
  XOR U21070 ( .A(n21083), .B(n21082), .Z(n21081) );
  NOR U21071 ( .A(n22112), .B(p_input[828]), .Z(n21082) );
  XOR U21072 ( .A(n21085), .B(n21084), .Z(n21083) );
  NOR U21073 ( .A(n22114), .B(p_input[826]), .Z(n21084) );
  XOR U21074 ( .A(n21087), .B(n21086), .Z(n21085) );
  NOR U21075 ( .A(n22116), .B(p_input[824]), .Z(n21086) );
  XOR U21076 ( .A(n21089), .B(n21088), .Z(n21087) );
  NOR U21077 ( .A(n22118), .B(p_input[822]), .Z(n21088) );
  XOR U21078 ( .A(n21091), .B(n21090), .Z(n21089) );
  NOR U21079 ( .A(n22120), .B(p_input[820]), .Z(n21090) );
  XOR U21080 ( .A(n21093), .B(n21092), .Z(n21091) );
  NOR U21081 ( .A(n22122), .B(p_input[818]), .Z(n21092) );
  XOR U21082 ( .A(n21095), .B(n21094), .Z(n21093) );
  NOR U21083 ( .A(n22124), .B(p_input[816]), .Z(n21094) );
  XOR U21084 ( .A(n21097), .B(n21096), .Z(n21095) );
  NOR U21085 ( .A(n22126), .B(p_input[814]), .Z(n21096) );
  XOR U21086 ( .A(n21099), .B(n21098), .Z(n21097) );
  NOR U21087 ( .A(n22128), .B(p_input[812]), .Z(n21098) );
  XOR U21088 ( .A(n21101), .B(n21100), .Z(n21099) );
  NOR U21089 ( .A(n22130), .B(p_input[810]), .Z(n21100) );
  XOR U21090 ( .A(n21103), .B(n21102), .Z(n21101) );
  NOR U21091 ( .A(n22132), .B(p_input[808]), .Z(n21102) );
  XOR U21092 ( .A(n21105), .B(n21104), .Z(n21103) );
  NOR U21093 ( .A(n22134), .B(p_input[806]), .Z(n21104) );
  XOR U21094 ( .A(n21107), .B(n21106), .Z(n21105) );
  NOR U21095 ( .A(n22136), .B(p_input[804]), .Z(n21106) );
  XOR U21096 ( .A(n21109), .B(n21108), .Z(n21107) );
  NOR U21097 ( .A(n22138), .B(p_input[802]), .Z(n21108) );
  XOR U21098 ( .A(n21111), .B(n21110), .Z(n21109) );
  NOR U21099 ( .A(n22140), .B(p_input[800]), .Z(n21110) );
  XOR U21100 ( .A(n21113), .B(n21112), .Z(n21111) );
  NOR U21101 ( .A(n22142), .B(p_input[798]), .Z(n21112) );
  XOR U21102 ( .A(n21115), .B(n21114), .Z(n21113) );
  NOR U21103 ( .A(n22144), .B(p_input[796]), .Z(n21114) );
  XOR U21104 ( .A(n21117), .B(n21116), .Z(n21115) );
  NOR U21105 ( .A(n22146), .B(p_input[794]), .Z(n21116) );
  XOR U21106 ( .A(n21119), .B(n21118), .Z(n21117) );
  NOR U21107 ( .A(n22148), .B(p_input[792]), .Z(n21118) );
  XOR U21108 ( .A(n21121), .B(n21120), .Z(n21119) );
  NOR U21109 ( .A(n22150), .B(p_input[790]), .Z(n21120) );
  XOR U21110 ( .A(n21123), .B(n21122), .Z(n21121) );
  NOR U21111 ( .A(n22152), .B(p_input[788]), .Z(n21122) );
  XOR U21112 ( .A(n21125), .B(n21124), .Z(n21123) );
  NOR U21113 ( .A(n22154), .B(p_input[786]), .Z(n21124) );
  XOR U21114 ( .A(n21127), .B(n21126), .Z(n21125) );
  NOR U21115 ( .A(n22156), .B(p_input[784]), .Z(n21126) );
  XOR U21116 ( .A(n21129), .B(n21128), .Z(n21127) );
  NOR U21117 ( .A(n22158), .B(p_input[782]), .Z(n21128) );
  XOR U21118 ( .A(n21131), .B(n21130), .Z(n21129) );
  NOR U21119 ( .A(n22160), .B(p_input[780]), .Z(n21130) );
  XOR U21120 ( .A(n21133), .B(n21132), .Z(n21131) );
  NOR U21121 ( .A(n22162), .B(p_input[778]), .Z(n21132) );
  XOR U21122 ( .A(n21135), .B(n21134), .Z(n21133) );
  NOR U21123 ( .A(n22164), .B(p_input[776]), .Z(n21134) );
  XOR U21124 ( .A(n21137), .B(n21136), .Z(n21135) );
  NOR U21125 ( .A(n22166), .B(p_input[774]), .Z(n21136) );
  XOR U21126 ( .A(n21139), .B(n21138), .Z(n21137) );
  NOR U21127 ( .A(n22168), .B(p_input[772]), .Z(n21138) );
  XOR U21128 ( .A(n21141), .B(n21140), .Z(n21139) );
  NOR U21129 ( .A(n22170), .B(p_input[770]), .Z(n21140) );
  XOR U21130 ( .A(n21143), .B(n21142), .Z(n21141) );
  NOR U21131 ( .A(n22172), .B(p_input[768]), .Z(n21142) );
  XOR U21132 ( .A(n21145), .B(n21144), .Z(n21143) );
  NOR U21133 ( .A(n22174), .B(p_input[766]), .Z(n21144) );
  XOR U21134 ( .A(n21147), .B(n21146), .Z(n21145) );
  NOR U21135 ( .A(n22176), .B(p_input[764]), .Z(n21146) );
  XOR U21136 ( .A(n21149), .B(n21148), .Z(n21147) );
  NOR U21137 ( .A(n22178), .B(p_input[762]), .Z(n21148) );
  XOR U21138 ( .A(n21151), .B(n21150), .Z(n21149) );
  NOR U21139 ( .A(n22180), .B(p_input[760]), .Z(n21150) );
  XOR U21140 ( .A(n21153), .B(n21152), .Z(n21151) );
  NOR U21141 ( .A(n22182), .B(p_input[758]), .Z(n21152) );
  XOR U21142 ( .A(n21155), .B(n21154), .Z(n21153) );
  NOR U21143 ( .A(n22184), .B(p_input[756]), .Z(n21154) );
  XOR U21144 ( .A(n21157), .B(n21156), .Z(n21155) );
  NOR U21145 ( .A(n22186), .B(p_input[754]), .Z(n21156) );
  XOR U21146 ( .A(n21159), .B(n21158), .Z(n21157) );
  NOR U21147 ( .A(n22188), .B(p_input[752]), .Z(n21158) );
  XOR U21148 ( .A(n21161), .B(n21160), .Z(n21159) );
  NOR U21149 ( .A(n22190), .B(p_input[750]), .Z(n21160) );
  XOR U21150 ( .A(n21163), .B(n21162), .Z(n21161) );
  NOR U21151 ( .A(n22192), .B(p_input[748]), .Z(n21162) );
  XOR U21152 ( .A(n21165), .B(n21164), .Z(n21163) );
  NOR U21153 ( .A(n22194), .B(p_input[746]), .Z(n21164) );
  XOR U21154 ( .A(n21167), .B(n21166), .Z(n21165) );
  NOR U21155 ( .A(n22196), .B(p_input[744]), .Z(n21166) );
  XOR U21156 ( .A(n21169), .B(n21168), .Z(n21167) );
  NOR U21157 ( .A(n22198), .B(p_input[742]), .Z(n21168) );
  XOR U21158 ( .A(n21171), .B(n21170), .Z(n21169) );
  NOR U21159 ( .A(n22200), .B(p_input[740]), .Z(n21170) );
  XOR U21160 ( .A(n21173), .B(n21172), .Z(n21171) );
  NOR U21161 ( .A(n22202), .B(p_input[738]), .Z(n21172) );
  XOR U21162 ( .A(n21175), .B(n21174), .Z(n21173) );
  NOR U21163 ( .A(n22204), .B(p_input[736]), .Z(n21174) );
  XOR U21164 ( .A(n21177), .B(n21176), .Z(n21175) );
  NOR U21165 ( .A(n22206), .B(p_input[734]), .Z(n21176) );
  XOR U21166 ( .A(n21179), .B(n21178), .Z(n21177) );
  NOR U21167 ( .A(n22208), .B(p_input[732]), .Z(n21178) );
  XOR U21168 ( .A(n21181), .B(n21180), .Z(n21179) );
  NOR U21169 ( .A(n22210), .B(p_input[730]), .Z(n21180) );
  XOR U21170 ( .A(n21183), .B(n21182), .Z(n21181) );
  NOR U21171 ( .A(n22212), .B(p_input[728]), .Z(n21182) );
  XOR U21172 ( .A(n21185), .B(n21184), .Z(n21183) );
  NOR U21173 ( .A(n22214), .B(p_input[726]), .Z(n21184) );
  XOR U21174 ( .A(n21187), .B(n21186), .Z(n21185) );
  NOR U21175 ( .A(n22216), .B(p_input[724]), .Z(n21186) );
  XOR U21176 ( .A(n21189), .B(n21188), .Z(n21187) );
  NOR U21177 ( .A(n22218), .B(p_input[722]), .Z(n21188) );
  XOR U21178 ( .A(n21191), .B(n21190), .Z(n21189) );
  NOR U21179 ( .A(n22220), .B(p_input[720]), .Z(n21190) );
  XOR U21180 ( .A(n21193), .B(n21192), .Z(n21191) );
  NOR U21181 ( .A(n22222), .B(p_input[718]), .Z(n21192) );
  XOR U21182 ( .A(n21195), .B(n21194), .Z(n21193) );
  NOR U21183 ( .A(n22224), .B(p_input[716]), .Z(n21194) );
  XOR U21184 ( .A(n21197), .B(n21196), .Z(n21195) );
  NOR U21185 ( .A(n22226), .B(p_input[714]), .Z(n21196) );
  XOR U21186 ( .A(n21199), .B(n21198), .Z(n21197) );
  NOR U21187 ( .A(n22228), .B(p_input[712]), .Z(n21198) );
  XOR U21188 ( .A(n21201), .B(n21200), .Z(n21199) );
  NOR U21189 ( .A(n22230), .B(p_input[710]), .Z(n21200) );
  XOR U21190 ( .A(n21203), .B(n21202), .Z(n21201) );
  NOR U21191 ( .A(n22232), .B(p_input[708]), .Z(n21202) );
  XOR U21192 ( .A(n21205), .B(n21204), .Z(n21203) );
  NOR U21193 ( .A(n22234), .B(p_input[706]), .Z(n21204) );
  XOR U21194 ( .A(n21207), .B(n21206), .Z(n21205) );
  NOR U21195 ( .A(n22236), .B(p_input[704]), .Z(n21206) );
  XOR U21196 ( .A(n21209), .B(n21208), .Z(n21207) );
  NOR U21197 ( .A(n22238), .B(p_input[702]), .Z(n21208) );
  XOR U21198 ( .A(n21211), .B(n21210), .Z(n21209) );
  NOR U21199 ( .A(n22240), .B(p_input[700]), .Z(n21210) );
  XOR U21200 ( .A(n21213), .B(n21212), .Z(n21211) );
  NOR U21201 ( .A(n22242), .B(p_input[698]), .Z(n21212) );
  XOR U21202 ( .A(n21215), .B(n21214), .Z(n21213) );
  NOR U21203 ( .A(n22244), .B(p_input[696]), .Z(n21214) );
  XOR U21204 ( .A(n21217), .B(n21216), .Z(n21215) );
  NOR U21205 ( .A(n22246), .B(p_input[694]), .Z(n21216) );
  XOR U21206 ( .A(n21219), .B(n21218), .Z(n21217) );
  NOR U21207 ( .A(n22248), .B(p_input[692]), .Z(n21218) );
  XOR U21208 ( .A(n21221), .B(n21220), .Z(n21219) );
  NOR U21209 ( .A(n22250), .B(p_input[690]), .Z(n21220) );
  XOR U21210 ( .A(n21223), .B(n21222), .Z(n21221) );
  NOR U21211 ( .A(n22252), .B(p_input[688]), .Z(n21222) );
  XOR U21212 ( .A(n21225), .B(n21224), .Z(n21223) );
  NOR U21213 ( .A(n22254), .B(p_input[686]), .Z(n21224) );
  XOR U21214 ( .A(n21227), .B(n21226), .Z(n21225) );
  NOR U21215 ( .A(n22256), .B(p_input[684]), .Z(n21226) );
  XOR U21216 ( .A(n21229), .B(n21228), .Z(n21227) );
  NOR U21217 ( .A(n22258), .B(p_input[682]), .Z(n21228) );
  XOR U21218 ( .A(n21231), .B(n21230), .Z(n21229) );
  NOR U21219 ( .A(n22260), .B(p_input[680]), .Z(n21230) );
  XOR U21220 ( .A(n21233), .B(n21232), .Z(n21231) );
  NOR U21221 ( .A(n22262), .B(p_input[678]), .Z(n21232) );
  XOR U21222 ( .A(n21235), .B(n21234), .Z(n21233) );
  NOR U21223 ( .A(n22264), .B(p_input[676]), .Z(n21234) );
  XOR U21224 ( .A(n21237), .B(n21236), .Z(n21235) );
  NOR U21225 ( .A(n22266), .B(p_input[674]), .Z(n21236) );
  XOR U21226 ( .A(n21239), .B(n21238), .Z(n21237) );
  NOR U21227 ( .A(n22268), .B(p_input[672]), .Z(n21238) );
  XOR U21228 ( .A(n21241), .B(n21240), .Z(n21239) );
  NOR U21229 ( .A(n22270), .B(p_input[670]), .Z(n21240) );
  XOR U21230 ( .A(n21243), .B(n21242), .Z(n21241) );
  NOR U21231 ( .A(n22272), .B(p_input[668]), .Z(n21242) );
  XOR U21232 ( .A(n21245), .B(n21244), .Z(n21243) );
  NOR U21233 ( .A(n22274), .B(p_input[666]), .Z(n21244) );
  XOR U21234 ( .A(n21247), .B(n21246), .Z(n21245) );
  NOR U21235 ( .A(n22276), .B(p_input[664]), .Z(n21246) );
  XOR U21236 ( .A(n21249), .B(n21248), .Z(n21247) );
  NOR U21237 ( .A(n22278), .B(p_input[662]), .Z(n21248) );
  XOR U21238 ( .A(n21251), .B(n21250), .Z(n21249) );
  NOR U21239 ( .A(n22280), .B(p_input[660]), .Z(n21250) );
  XOR U21240 ( .A(n21253), .B(n21252), .Z(n21251) );
  NOR U21241 ( .A(n22282), .B(p_input[658]), .Z(n21252) );
  XOR U21242 ( .A(n21255), .B(n21254), .Z(n21253) );
  NOR U21243 ( .A(n22284), .B(p_input[656]), .Z(n21254) );
  XOR U21244 ( .A(n21257), .B(n21256), .Z(n21255) );
  NOR U21245 ( .A(n22286), .B(p_input[654]), .Z(n21256) );
  XOR U21246 ( .A(n21259), .B(n21258), .Z(n21257) );
  NOR U21247 ( .A(n22288), .B(p_input[652]), .Z(n21258) );
  XOR U21248 ( .A(n21261), .B(n21260), .Z(n21259) );
  NOR U21249 ( .A(n22290), .B(p_input[650]), .Z(n21260) );
  XOR U21250 ( .A(n21263), .B(n21262), .Z(n21261) );
  NOR U21251 ( .A(n22292), .B(p_input[648]), .Z(n21262) );
  XOR U21252 ( .A(n21265), .B(n21264), .Z(n21263) );
  NOR U21253 ( .A(n22294), .B(p_input[646]), .Z(n21264) );
  XOR U21254 ( .A(n21267), .B(n21266), .Z(n21265) );
  NOR U21255 ( .A(n22296), .B(p_input[644]), .Z(n21266) );
  XOR U21256 ( .A(n21269), .B(n21268), .Z(n21267) );
  NOR U21257 ( .A(n22298), .B(p_input[642]), .Z(n21268) );
  XOR U21258 ( .A(n21271), .B(n21270), .Z(n21269) );
  NOR U21259 ( .A(n22300), .B(p_input[640]), .Z(n21270) );
  XOR U21260 ( .A(n21273), .B(n21272), .Z(n21271) );
  NOR U21261 ( .A(n22302), .B(p_input[638]), .Z(n21272) );
  XOR U21262 ( .A(n21275), .B(n21274), .Z(n21273) );
  NOR U21263 ( .A(n22304), .B(p_input[636]), .Z(n21274) );
  XOR U21264 ( .A(n21277), .B(n21276), .Z(n21275) );
  NOR U21265 ( .A(n22306), .B(p_input[634]), .Z(n21276) );
  XOR U21266 ( .A(n21279), .B(n21278), .Z(n21277) );
  NOR U21267 ( .A(n22308), .B(p_input[632]), .Z(n21278) );
  XOR U21268 ( .A(n21281), .B(n21280), .Z(n21279) );
  NOR U21269 ( .A(n22310), .B(p_input[630]), .Z(n21280) );
  XOR U21270 ( .A(n21283), .B(n21282), .Z(n21281) );
  NOR U21271 ( .A(n22312), .B(p_input[628]), .Z(n21282) );
  XOR U21272 ( .A(n21285), .B(n21284), .Z(n21283) );
  NOR U21273 ( .A(n22314), .B(p_input[626]), .Z(n21284) );
  XOR U21274 ( .A(n21287), .B(n21286), .Z(n21285) );
  NOR U21275 ( .A(n22316), .B(p_input[624]), .Z(n21286) );
  XOR U21276 ( .A(n21289), .B(n21288), .Z(n21287) );
  NOR U21277 ( .A(n22318), .B(p_input[622]), .Z(n21288) );
  XOR U21278 ( .A(n21291), .B(n21290), .Z(n21289) );
  NOR U21279 ( .A(n22320), .B(p_input[620]), .Z(n21290) );
  XOR U21280 ( .A(n21293), .B(n21292), .Z(n21291) );
  NOR U21281 ( .A(n22322), .B(p_input[618]), .Z(n21292) );
  XOR U21282 ( .A(n21295), .B(n21294), .Z(n21293) );
  NOR U21283 ( .A(n22324), .B(p_input[616]), .Z(n21294) );
  XOR U21284 ( .A(n21297), .B(n21296), .Z(n21295) );
  NOR U21285 ( .A(n22326), .B(p_input[614]), .Z(n21296) );
  XOR U21286 ( .A(n21299), .B(n21298), .Z(n21297) );
  NOR U21287 ( .A(n22328), .B(p_input[612]), .Z(n21298) );
  XOR U21288 ( .A(n21301), .B(n21300), .Z(n21299) );
  NOR U21289 ( .A(n22330), .B(p_input[610]), .Z(n21300) );
  XOR U21290 ( .A(n21303), .B(n21302), .Z(n21301) );
  NOR U21291 ( .A(n22332), .B(p_input[608]), .Z(n21302) );
  XOR U21292 ( .A(n21305), .B(n21304), .Z(n21303) );
  NOR U21293 ( .A(n22334), .B(p_input[606]), .Z(n21304) );
  XOR U21294 ( .A(n21307), .B(n21306), .Z(n21305) );
  NOR U21295 ( .A(n22336), .B(p_input[604]), .Z(n21306) );
  XOR U21296 ( .A(n21309), .B(n21308), .Z(n21307) );
  NOR U21297 ( .A(n22338), .B(p_input[602]), .Z(n21308) );
  XOR U21298 ( .A(n21311), .B(n21310), .Z(n21309) );
  NOR U21299 ( .A(n22340), .B(p_input[600]), .Z(n21310) );
  XOR U21300 ( .A(n21313), .B(n21312), .Z(n21311) );
  NOR U21301 ( .A(n22342), .B(p_input[598]), .Z(n21312) );
  XOR U21302 ( .A(n21315), .B(n21314), .Z(n21313) );
  NOR U21303 ( .A(n22344), .B(p_input[596]), .Z(n21314) );
  XOR U21304 ( .A(n21317), .B(n21316), .Z(n21315) );
  NOR U21305 ( .A(n22346), .B(p_input[594]), .Z(n21316) );
  XOR U21306 ( .A(n21319), .B(n21318), .Z(n21317) );
  NOR U21307 ( .A(n22348), .B(p_input[592]), .Z(n21318) );
  XOR U21308 ( .A(n21321), .B(n21320), .Z(n21319) );
  NOR U21309 ( .A(n22350), .B(p_input[590]), .Z(n21320) );
  XOR U21310 ( .A(n21323), .B(n21322), .Z(n21321) );
  NOR U21311 ( .A(n22352), .B(p_input[588]), .Z(n21322) );
  XOR U21312 ( .A(n21325), .B(n21324), .Z(n21323) );
  NOR U21313 ( .A(n22354), .B(p_input[586]), .Z(n21324) );
  XOR U21314 ( .A(n21327), .B(n21326), .Z(n21325) );
  NOR U21315 ( .A(n22356), .B(p_input[584]), .Z(n21326) );
  XOR U21316 ( .A(n21329), .B(n21328), .Z(n21327) );
  NOR U21317 ( .A(n22358), .B(p_input[582]), .Z(n21328) );
  XOR U21318 ( .A(n21331), .B(n21330), .Z(n21329) );
  NOR U21319 ( .A(n22360), .B(p_input[580]), .Z(n21330) );
  XOR U21320 ( .A(n21333), .B(n21332), .Z(n21331) );
  NOR U21321 ( .A(n22362), .B(p_input[578]), .Z(n21332) );
  XOR U21322 ( .A(n21335), .B(n21334), .Z(n21333) );
  NOR U21323 ( .A(n22364), .B(p_input[576]), .Z(n21334) );
  XOR U21324 ( .A(n21337), .B(n21336), .Z(n21335) );
  NOR U21325 ( .A(n22366), .B(p_input[574]), .Z(n21336) );
  XOR U21326 ( .A(n21339), .B(n21338), .Z(n21337) );
  NOR U21327 ( .A(n22368), .B(p_input[572]), .Z(n21338) );
  XOR U21328 ( .A(n21341), .B(n21340), .Z(n21339) );
  NOR U21329 ( .A(n22370), .B(p_input[570]), .Z(n21340) );
  XOR U21330 ( .A(n21343), .B(n21342), .Z(n21341) );
  NOR U21331 ( .A(n22372), .B(p_input[568]), .Z(n21342) );
  XOR U21332 ( .A(n21345), .B(n21344), .Z(n21343) );
  NOR U21333 ( .A(n22374), .B(p_input[566]), .Z(n21344) );
  XOR U21334 ( .A(n21347), .B(n21346), .Z(n21345) );
  NOR U21335 ( .A(n22376), .B(p_input[564]), .Z(n21346) );
  XOR U21336 ( .A(n21349), .B(n21348), .Z(n21347) );
  NOR U21337 ( .A(n22378), .B(p_input[562]), .Z(n21348) );
  XOR U21338 ( .A(n21351), .B(n21350), .Z(n21349) );
  NOR U21339 ( .A(n22380), .B(p_input[560]), .Z(n21350) );
  XOR U21340 ( .A(n21353), .B(n21352), .Z(n21351) );
  NOR U21341 ( .A(n22382), .B(p_input[558]), .Z(n21352) );
  XOR U21342 ( .A(n21355), .B(n21354), .Z(n21353) );
  NOR U21343 ( .A(n22384), .B(p_input[556]), .Z(n21354) );
  XOR U21344 ( .A(n21357), .B(n21356), .Z(n21355) );
  NOR U21345 ( .A(n22386), .B(p_input[554]), .Z(n21356) );
  XOR U21346 ( .A(n21359), .B(n21358), .Z(n21357) );
  NOR U21347 ( .A(n22388), .B(p_input[552]), .Z(n21358) );
  XOR U21348 ( .A(n21361), .B(n21360), .Z(n21359) );
  NOR U21349 ( .A(n22390), .B(p_input[550]), .Z(n21360) );
  XOR U21350 ( .A(n21363), .B(n21362), .Z(n21361) );
  NOR U21351 ( .A(n22392), .B(p_input[548]), .Z(n21362) );
  XOR U21352 ( .A(n21365), .B(n21364), .Z(n21363) );
  NOR U21353 ( .A(n22394), .B(p_input[546]), .Z(n21364) );
  XOR U21354 ( .A(n21367), .B(n21366), .Z(n21365) );
  NOR U21355 ( .A(n22396), .B(p_input[544]), .Z(n21366) );
  XOR U21356 ( .A(n21369), .B(n21368), .Z(n21367) );
  NOR U21357 ( .A(n22398), .B(p_input[542]), .Z(n21368) );
  XOR U21358 ( .A(n21371), .B(n21370), .Z(n21369) );
  NOR U21359 ( .A(n22400), .B(p_input[540]), .Z(n21370) );
  XOR U21360 ( .A(n21373), .B(n21372), .Z(n21371) );
  NOR U21361 ( .A(n22402), .B(p_input[538]), .Z(n21372) );
  XOR U21362 ( .A(n21375), .B(n21374), .Z(n21373) );
  NOR U21363 ( .A(n22404), .B(p_input[536]), .Z(n21374) );
  XOR U21364 ( .A(n21377), .B(n21376), .Z(n21375) );
  NOR U21365 ( .A(n22406), .B(p_input[534]), .Z(n21376) );
  XOR U21366 ( .A(n21379), .B(n21378), .Z(n21377) );
  NOR U21367 ( .A(n22408), .B(p_input[532]), .Z(n21378) );
  XOR U21368 ( .A(n21381), .B(n21380), .Z(n21379) );
  NOR U21369 ( .A(n22410), .B(p_input[530]), .Z(n21380) );
  XOR U21370 ( .A(n21383), .B(n21382), .Z(n21381) );
  NOR U21371 ( .A(n22412), .B(p_input[528]), .Z(n21382) );
  XOR U21372 ( .A(n21385), .B(n21384), .Z(n21383) );
  NOR U21373 ( .A(n22414), .B(p_input[526]), .Z(n21384) );
  XOR U21374 ( .A(n21387), .B(n21386), .Z(n21385) );
  NOR U21375 ( .A(n22416), .B(p_input[524]), .Z(n21386) );
  XOR U21376 ( .A(n21389), .B(n21388), .Z(n21387) );
  NOR U21377 ( .A(n22418), .B(p_input[522]), .Z(n21388) );
  XOR U21378 ( .A(n21391), .B(n21390), .Z(n21389) );
  NOR U21379 ( .A(n22420), .B(p_input[520]), .Z(n21390) );
  XOR U21380 ( .A(n21393), .B(n21392), .Z(n21391) );
  NOR U21381 ( .A(n22422), .B(p_input[518]), .Z(n21392) );
  XOR U21382 ( .A(n21395), .B(n21394), .Z(n21393) );
  NOR U21383 ( .A(n22424), .B(p_input[516]), .Z(n21394) );
  XOR U21384 ( .A(n21397), .B(n21396), .Z(n21395) );
  NOR U21385 ( .A(n22426), .B(p_input[514]), .Z(n21396) );
  XOR U21386 ( .A(n21399), .B(n21398), .Z(n21397) );
  NOR U21387 ( .A(n22428), .B(p_input[512]), .Z(n21398) );
  XOR U21388 ( .A(n21401), .B(n21400), .Z(n21399) );
  NOR U21389 ( .A(n22430), .B(p_input[510]), .Z(n21400) );
  XOR U21390 ( .A(n21403), .B(n21402), .Z(n21401) );
  NOR U21391 ( .A(n22432), .B(p_input[508]), .Z(n21402) );
  XOR U21392 ( .A(n21405), .B(n21404), .Z(n21403) );
  NOR U21393 ( .A(n22434), .B(p_input[506]), .Z(n21404) );
  XOR U21394 ( .A(n21407), .B(n21406), .Z(n21405) );
  NOR U21395 ( .A(n22436), .B(p_input[504]), .Z(n21406) );
  XOR U21396 ( .A(n21409), .B(n21408), .Z(n21407) );
  NOR U21397 ( .A(n22438), .B(p_input[502]), .Z(n21408) );
  XOR U21398 ( .A(n21411), .B(n21410), .Z(n21409) );
  NOR U21399 ( .A(n22440), .B(p_input[500]), .Z(n21410) );
  XOR U21400 ( .A(n21413), .B(n21412), .Z(n21411) );
  NOR U21401 ( .A(n22442), .B(p_input[498]), .Z(n21412) );
  XOR U21402 ( .A(n21415), .B(n21414), .Z(n21413) );
  NOR U21403 ( .A(n22444), .B(p_input[496]), .Z(n21414) );
  XOR U21404 ( .A(n21417), .B(n21416), .Z(n21415) );
  NOR U21405 ( .A(n22446), .B(p_input[494]), .Z(n21416) );
  XOR U21406 ( .A(n21419), .B(n21418), .Z(n21417) );
  NOR U21407 ( .A(n22448), .B(p_input[492]), .Z(n21418) );
  XOR U21408 ( .A(n21421), .B(n21420), .Z(n21419) );
  NOR U21409 ( .A(n22450), .B(p_input[490]), .Z(n21420) );
  XOR U21410 ( .A(n21423), .B(n21422), .Z(n21421) );
  NOR U21411 ( .A(n22452), .B(p_input[488]), .Z(n21422) );
  XOR U21412 ( .A(n21425), .B(n21424), .Z(n21423) );
  NOR U21413 ( .A(n22454), .B(p_input[486]), .Z(n21424) );
  XOR U21414 ( .A(n21427), .B(n21426), .Z(n21425) );
  NOR U21415 ( .A(n22456), .B(p_input[484]), .Z(n21426) );
  XOR U21416 ( .A(n21429), .B(n21428), .Z(n21427) );
  NOR U21417 ( .A(n22458), .B(p_input[482]), .Z(n21428) );
  XOR U21418 ( .A(n21431), .B(n21430), .Z(n21429) );
  NOR U21419 ( .A(n22460), .B(p_input[480]), .Z(n21430) );
  XOR U21420 ( .A(n21433), .B(n21432), .Z(n21431) );
  NOR U21421 ( .A(n22462), .B(p_input[478]), .Z(n21432) );
  XOR U21422 ( .A(n21435), .B(n21434), .Z(n21433) );
  NOR U21423 ( .A(n22464), .B(p_input[476]), .Z(n21434) );
  XOR U21424 ( .A(n21437), .B(n21436), .Z(n21435) );
  NOR U21425 ( .A(n22466), .B(p_input[474]), .Z(n21436) );
  XOR U21426 ( .A(n21439), .B(n21438), .Z(n21437) );
  NOR U21427 ( .A(n22468), .B(p_input[472]), .Z(n21438) );
  XOR U21428 ( .A(n21441), .B(n21440), .Z(n21439) );
  NOR U21429 ( .A(n22470), .B(p_input[470]), .Z(n21440) );
  XOR U21430 ( .A(n21443), .B(n21442), .Z(n21441) );
  NOR U21431 ( .A(n22472), .B(p_input[468]), .Z(n21442) );
  XOR U21432 ( .A(n21445), .B(n21444), .Z(n21443) );
  NOR U21433 ( .A(n22474), .B(p_input[466]), .Z(n21444) );
  XOR U21434 ( .A(n21447), .B(n21446), .Z(n21445) );
  NOR U21435 ( .A(n22476), .B(p_input[464]), .Z(n21446) );
  XOR U21436 ( .A(n21449), .B(n21448), .Z(n21447) );
  NOR U21437 ( .A(n22478), .B(p_input[462]), .Z(n21448) );
  XOR U21438 ( .A(n21451), .B(n21450), .Z(n21449) );
  NOR U21439 ( .A(n22480), .B(p_input[460]), .Z(n21450) );
  XOR U21440 ( .A(n21453), .B(n21452), .Z(n21451) );
  NOR U21441 ( .A(n22482), .B(p_input[458]), .Z(n21452) );
  XOR U21442 ( .A(n21455), .B(n21454), .Z(n21453) );
  NOR U21443 ( .A(n22484), .B(p_input[456]), .Z(n21454) );
  XOR U21444 ( .A(n21457), .B(n21456), .Z(n21455) );
  NOR U21445 ( .A(n22486), .B(p_input[454]), .Z(n21456) );
  XOR U21446 ( .A(n21459), .B(n21458), .Z(n21457) );
  NOR U21447 ( .A(n22488), .B(p_input[452]), .Z(n21458) );
  XOR U21448 ( .A(n21461), .B(n21460), .Z(n21459) );
  NOR U21449 ( .A(n22490), .B(p_input[450]), .Z(n21460) );
  XOR U21450 ( .A(n21463), .B(n21462), .Z(n21461) );
  NOR U21451 ( .A(n22492), .B(p_input[448]), .Z(n21462) );
  XOR U21452 ( .A(n21465), .B(n21464), .Z(n21463) );
  NOR U21453 ( .A(n22494), .B(p_input[446]), .Z(n21464) );
  XOR U21454 ( .A(n21467), .B(n21466), .Z(n21465) );
  NOR U21455 ( .A(n22496), .B(p_input[444]), .Z(n21466) );
  XOR U21456 ( .A(n21469), .B(n21468), .Z(n21467) );
  NOR U21457 ( .A(n22498), .B(p_input[442]), .Z(n21468) );
  XOR U21458 ( .A(n21471), .B(n21470), .Z(n21469) );
  NOR U21459 ( .A(n22500), .B(p_input[440]), .Z(n21470) );
  XOR U21460 ( .A(n21473), .B(n21472), .Z(n21471) );
  NOR U21461 ( .A(n22502), .B(p_input[438]), .Z(n21472) );
  XOR U21462 ( .A(n21475), .B(n21474), .Z(n21473) );
  NOR U21463 ( .A(n22504), .B(p_input[436]), .Z(n21474) );
  XOR U21464 ( .A(n21477), .B(n21476), .Z(n21475) );
  NOR U21465 ( .A(n22506), .B(p_input[434]), .Z(n21476) );
  XOR U21466 ( .A(n21479), .B(n21478), .Z(n21477) );
  NOR U21467 ( .A(n22508), .B(p_input[432]), .Z(n21478) );
  XOR U21468 ( .A(n21481), .B(n21480), .Z(n21479) );
  NOR U21469 ( .A(n22510), .B(p_input[430]), .Z(n21480) );
  XOR U21470 ( .A(n21483), .B(n21482), .Z(n21481) );
  NOR U21471 ( .A(n22512), .B(p_input[428]), .Z(n21482) );
  XOR U21472 ( .A(n21485), .B(n21484), .Z(n21483) );
  NOR U21473 ( .A(n22514), .B(p_input[426]), .Z(n21484) );
  XOR U21474 ( .A(n21487), .B(n21486), .Z(n21485) );
  NOR U21475 ( .A(n22516), .B(p_input[424]), .Z(n21486) );
  XOR U21476 ( .A(n21489), .B(n21488), .Z(n21487) );
  NOR U21477 ( .A(n22518), .B(p_input[422]), .Z(n21488) );
  XOR U21478 ( .A(n21491), .B(n21490), .Z(n21489) );
  NOR U21479 ( .A(n22520), .B(p_input[420]), .Z(n21490) );
  XOR U21480 ( .A(n21493), .B(n21492), .Z(n21491) );
  NOR U21481 ( .A(n22522), .B(p_input[418]), .Z(n21492) );
  XOR U21482 ( .A(n21495), .B(n21494), .Z(n21493) );
  NOR U21483 ( .A(n22524), .B(p_input[416]), .Z(n21494) );
  XOR U21484 ( .A(n21497), .B(n21496), .Z(n21495) );
  NOR U21485 ( .A(n22526), .B(p_input[414]), .Z(n21496) );
  XOR U21486 ( .A(n21499), .B(n21498), .Z(n21497) );
  NOR U21487 ( .A(n22528), .B(p_input[412]), .Z(n21498) );
  XOR U21488 ( .A(n21501), .B(n21500), .Z(n21499) );
  NOR U21489 ( .A(n22530), .B(p_input[410]), .Z(n21500) );
  XOR U21490 ( .A(n21503), .B(n21502), .Z(n21501) );
  NOR U21491 ( .A(n22532), .B(p_input[408]), .Z(n21502) );
  XOR U21492 ( .A(n21505), .B(n21504), .Z(n21503) );
  NOR U21493 ( .A(n22534), .B(p_input[406]), .Z(n21504) );
  XOR U21494 ( .A(n21507), .B(n21506), .Z(n21505) );
  NOR U21495 ( .A(n22536), .B(p_input[404]), .Z(n21506) );
  XOR U21496 ( .A(n21509), .B(n21508), .Z(n21507) );
  NOR U21497 ( .A(n22538), .B(p_input[402]), .Z(n21508) );
  XOR U21498 ( .A(n21511), .B(n21510), .Z(n21509) );
  NOR U21499 ( .A(n22540), .B(p_input[400]), .Z(n21510) );
  XOR U21500 ( .A(n21513), .B(n21512), .Z(n21511) );
  NOR U21501 ( .A(n22542), .B(p_input[398]), .Z(n21512) );
  XOR U21502 ( .A(n21515), .B(n21514), .Z(n21513) );
  NOR U21503 ( .A(n22544), .B(p_input[396]), .Z(n21514) );
  XOR U21504 ( .A(n21517), .B(n21516), .Z(n21515) );
  NOR U21505 ( .A(n22546), .B(p_input[394]), .Z(n21516) );
  XOR U21506 ( .A(n21519), .B(n21518), .Z(n21517) );
  NOR U21507 ( .A(n22548), .B(p_input[392]), .Z(n21518) );
  XOR U21508 ( .A(n21521), .B(n21520), .Z(n21519) );
  NOR U21509 ( .A(n22550), .B(p_input[390]), .Z(n21520) );
  XOR U21510 ( .A(n21523), .B(n21522), .Z(n21521) );
  NOR U21511 ( .A(n22552), .B(p_input[388]), .Z(n21522) );
  XOR U21512 ( .A(n21525), .B(n21524), .Z(n21523) );
  NOR U21513 ( .A(n22554), .B(p_input[386]), .Z(n21524) );
  XOR U21514 ( .A(n21527), .B(n21526), .Z(n21525) );
  NOR U21515 ( .A(n22556), .B(p_input[384]), .Z(n21526) );
  XOR U21516 ( .A(n21529), .B(n21528), .Z(n21527) );
  NOR U21517 ( .A(n22558), .B(p_input[382]), .Z(n21528) );
  XOR U21518 ( .A(n21531), .B(n21530), .Z(n21529) );
  NOR U21519 ( .A(n22560), .B(p_input[380]), .Z(n21530) );
  XOR U21520 ( .A(n21533), .B(n21532), .Z(n21531) );
  NOR U21521 ( .A(n22562), .B(p_input[378]), .Z(n21532) );
  XOR U21522 ( .A(n21535), .B(n21534), .Z(n21533) );
  NOR U21523 ( .A(n22564), .B(p_input[376]), .Z(n21534) );
  XOR U21524 ( .A(n21537), .B(n21536), .Z(n21535) );
  NOR U21525 ( .A(n22566), .B(p_input[374]), .Z(n21536) );
  XOR U21526 ( .A(n21539), .B(n21538), .Z(n21537) );
  NOR U21527 ( .A(n22568), .B(p_input[372]), .Z(n21538) );
  XOR U21528 ( .A(n21541), .B(n21540), .Z(n21539) );
  NOR U21529 ( .A(n22570), .B(p_input[370]), .Z(n21540) );
  XOR U21530 ( .A(n21543), .B(n21542), .Z(n21541) );
  NOR U21531 ( .A(n22572), .B(p_input[368]), .Z(n21542) );
  XOR U21532 ( .A(n21545), .B(n21544), .Z(n21543) );
  NOR U21533 ( .A(n22574), .B(p_input[366]), .Z(n21544) );
  XOR U21534 ( .A(n21547), .B(n21546), .Z(n21545) );
  NOR U21535 ( .A(n22576), .B(p_input[364]), .Z(n21546) );
  XOR U21536 ( .A(n21549), .B(n21548), .Z(n21547) );
  NOR U21537 ( .A(n22578), .B(p_input[362]), .Z(n21548) );
  XOR U21538 ( .A(n21551), .B(n21550), .Z(n21549) );
  NOR U21539 ( .A(n22580), .B(p_input[360]), .Z(n21550) );
  XOR U21540 ( .A(n21553), .B(n21552), .Z(n21551) );
  NOR U21541 ( .A(n22582), .B(p_input[358]), .Z(n21552) );
  XOR U21542 ( .A(n21555), .B(n21554), .Z(n21553) );
  NOR U21543 ( .A(n22584), .B(p_input[356]), .Z(n21554) );
  XOR U21544 ( .A(n21557), .B(n21556), .Z(n21555) );
  NOR U21545 ( .A(n22586), .B(p_input[354]), .Z(n21556) );
  XOR U21546 ( .A(n21559), .B(n21558), .Z(n21557) );
  NOR U21547 ( .A(n22588), .B(p_input[352]), .Z(n21558) );
  XOR U21548 ( .A(n21561), .B(n21560), .Z(n21559) );
  NOR U21549 ( .A(n22590), .B(p_input[350]), .Z(n21560) );
  XOR U21550 ( .A(n21563), .B(n21562), .Z(n21561) );
  NOR U21551 ( .A(n22592), .B(p_input[348]), .Z(n21562) );
  XOR U21552 ( .A(n21565), .B(n21564), .Z(n21563) );
  NOR U21553 ( .A(n22594), .B(p_input[346]), .Z(n21564) );
  XOR U21554 ( .A(n21567), .B(n21566), .Z(n21565) );
  NOR U21555 ( .A(n22596), .B(p_input[344]), .Z(n21566) );
  XOR U21556 ( .A(n21569), .B(n21568), .Z(n21567) );
  NOR U21557 ( .A(n22598), .B(p_input[342]), .Z(n21568) );
  XOR U21558 ( .A(n21571), .B(n21570), .Z(n21569) );
  NOR U21559 ( .A(n22600), .B(p_input[340]), .Z(n21570) );
  XOR U21560 ( .A(n21573), .B(n21572), .Z(n21571) );
  NOR U21561 ( .A(n22602), .B(p_input[338]), .Z(n21572) );
  XOR U21562 ( .A(n21575), .B(n21574), .Z(n21573) );
  NOR U21563 ( .A(n22604), .B(p_input[336]), .Z(n21574) );
  XOR U21564 ( .A(n21577), .B(n21576), .Z(n21575) );
  NOR U21565 ( .A(n22606), .B(p_input[334]), .Z(n21576) );
  XOR U21566 ( .A(n21579), .B(n21578), .Z(n21577) );
  NOR U21567 ( .A(n22608), .B(p_input[332]), .Z(n21578) );
  XOR U21568 ( .A(n21581), .B(n21580), .Z(n21579) );
  NOR U21569 ( .A(n22610), .B(p_input[330]), .Z(n21580) );
  XOR U21570 ( .A(n21583), .B(n21582), .Z(n21581) );
  NOR U21571 ( .A(n22612), .B(p_input[328]), .Z(n21582) );
  XOR U21572 ( .A(n21585), .B(n21584), .Z(n21583) );
  NOR U21573 ( .A(n22614), .B(p_input[326]), .Z(n21584) );
  XOR U21574 ( .A(n21587), .B(n21586), .Z(n21585) );
  NOR U21575 ( .A(n22616), .B(p_input[324]), .Z(n21586) );
  XOR U21576 ( .A(n21589), .B(n21588), .Z(n21587) );
  NOR U21577 ( .A(n22618), .B(p_input[322]), .Z(n21588) );
  XOR U21578 ( .A(n21591), .B(n21590), .Z(n21589) );
  NOR U21579 ( .A(n22620), .B(p_input[320]), .Z(n21590) );
  XOR U21580 ( .A(n21593), .B(n21592), .Z(n21591) );
  NOR U21581 ( .A(n22622), .B(p_input[318]), .Z(n21592) );
  XOR U21582 ( .A(n21595), .B(n21594), .Z(n21593) );
  NOR U21583 ( .A(n22624), .B(p_input[316]), .Z(n21594) );
  XOR U21584 ( .A(n21597), .B(n21596), .Z(n21595) );
  NOR U21585 ( .A(n22626), .B(p_input[314]), .Z(n21596) );
  XOR U21586 ( .A(n21599), .B(n21598), .Z(n21597) );
  NOR U21587 ( .A(n22628), .B(p_input[312]), .Z(n21598) );
  XOR U21588 ( .A(n21601), .B(n21600), .Z(n21599) );
  NOR U21589 ( .A(n22630), .B(p_input[310]), .Z(n21600) );
  XOR U21590 ( .A(n21603), .B(n21602), .Z(n21601) );
  NOR U21591 ( .A(n22632), .B(p_input[308]), .Z(n21602) );
  XOR U21592 ( .A(n21605), .B(n21604), .Z(n21603) );
  NOR U21593 ( .A(n22634), .B(p_input[306]), .Z(n21604) );
  XOR U21594 ( .A(n21607), .B(n21606), .Z(n21605) );
  NOR U21595 ( .A(n22636), .B(p_input[304]), .Z(n21606) );
  XOR U21596 ( .A(n21609), .B(n21608), .Z(n21607) );
  NOR U21597 ( .A(n22638), .B(p_input[302]), .Z(n21608) );
  XOR U21598 ( .A(n21611), .B(n21610), .Z(n21609) );
  NOR U21599 ( .A(n22640), .B(p_input[300]), .Z(n21610) );
  XOR U21600 ( .A(n21613), .B(n21612), .Z(n21611) );
  NOR U21601 ( .A(n22642), .B(p_input[298]), .Z(n21612) );
  XOR U21602 ( .A(n21615), .B(n21614), .Z(n21613) );
  NOR U21603 ( .A(n22644), .B(p_input[296]), .Z(n21614) );
  XOR U21604 ( .A(n21617), .B(n21616), .Z(n21615) );
  NOR U21605 ( .A(n22646), .B(p_input[294]), .Z(n21616) );
  XOR U21606 ( .A(n21619), .B(n21618), .Z(n21617) );
  NOR U21607 ( .A(n22648), .B(p_input[292]), .Z(n21618) );
  XOR U21608 ( .A(n21621), .B(n21620), .Z(n21619) );
  NOR U21609 ( .A(n22650), .B(p_input[290]), .Z(n21620) );
  XOR U21610 ( .A(n21623), .B(n21622), .Z(n21621) );
  NOR U21611 ( .A(n22652), .B(p_input[288]), .Z(n21622) );
  XOR U21612 ( .A(n21625), .B(n21624), .Z(n21623) );
  NOR U21613 ( .A(n22654), .B(p_input[286]), .Z(n21624) );
  XOR U21614 ( .A(n21627), .B(n21626), .Z(n21625) );
  NOR U21615 ( .A(n22656), .B(p_input[284]), .Z(n21626) );
  XOR U21616 ( .A(n21629), .B(n21628), .Z(n21627) );
  NOR U21617 ( .A(n22658), .B(p_input[282]), .Z(n21628) );
  XOR U21618 ( .A(n21631), .B(n21630), .Z(n21629) );
  NOR U21619 ( .A(n22660), .B(p_input[280]), .Z(n21630) );
  XOR U21620 ( .A(n21633), .B(n21632), .Z(n21631) );
  NOR U21621 ( .A(n22662), .B(p_input[278]), .Z(n21632) );
  XOR U21622 ( .A(n21635), .B(n21634), .Z(n21633) );
  NOR U21623 ( .A(n22664), .B(p_input[276]), .Z(n21634) );
  XOR U21624 ( .A(n21637), .B(n21636), .Z(n21635) );
  NOR U21625 ( .A(n22666), .B(p_input[274]), .Z(n21636) );
  XOR U21626 ( .A(n21639), .B(n21638), .Z(n21637) );
  NOR U21627 ( .A(n22668), .B(p_input[272]), .Z(n21638) );
  XOR U21628 ( .A(n21641), .B(n21640), .Z(n21639) );
  NOR U21629 ( .A(n22670), .B(p_input[270]), .Z(n21640) );
  XOR U21630 ( .A(n21643), .B(n21642), .Z(n21641) );
  NOR U21631 ( .A(n22672), .B(p_input[268]), .Z(n21642) );
  XOR U21632 ( .A(n21645), .B(n21644), .Z(n21643) );
  NOR U21633 ( .A(n22674), .B(p_input[266]), .Z(n21644) );
  XOR U21634 ( .A(n21647), .B(n21646), .Z(n21645) );
  NOR U21635 ( .A(n22676), .B(p_input[264]), .Z(n21646) );
  XOR U21636 ( .A(n21649), .B(n21648), .Z(n21647) );
  NOR U21637 ( .A(n22678), .B(p_input[262]), .Z(n21648) );
  XOR U21638 ( .A(n21651), .B(n21650), .Z(n21649) );
  NOR U21639 ( .A(n22680), .B(p_input[260]), .Z(n21650) );
  XOR U21640 ( .A(n21653), .B(n21652), .Z(n21651) );
  NOR U21641 ( .A(n22682), .B(p_input[258]), .Z(n21652) );
  XOR U21642 ( .A(n21655), .B(n21654), .Z(n21653) );
  NOR U21643 ( .A(n22684), .B(p_input[256]), .Z(n21654) );
  XOR U21644 ( .A(n21657), .B(n21656), .Z(n21655) );
  NOR U21645 ( .A(n22686), .B(p_input[254]), .Z(n21656) );
  XOR U21646 ( .A(n21661), .B(n21660), .Z(n21657) );
  NOR U21647 ( .A(n22688), .B(p_input[252]), .Z(n21660) );
  XOR U21648 ( .A(n21663), .B(n21662), .Z(n21661) );
  NOR U21649 ( .A(n22690), .B(p_input[250]), .Z(n21662) );
  XOR U21650 ( .A(n21665), .B(n21664), .Z(n21663) );
  NOR U21651 ( .A(n22692), .B(p_input[248]), .Z(n21664) );
  XOR U21652 ( .A(n21667), .B(n21666), .Z(n21665) );
  NOR U21653 ( .A(n22694), .B(p_input[246]), .Z(n21666) );
  XOR U21654 ( .A(n21669), .B(n21668), .Z(n21667) );
  NOR U21655 ( .A(n22696), .B(p_input[244]), .Z(n21668) );
  XOR U21656 ( .A(n21671), .B(n21670), .Z(n21669) );
  NOR U21657 ( .A(n22698), .B(p_input[242]), .Z(n21670) );
  XOR U21658 ( .A(n21673), .B(n21672), .Z(n21671) );
  NOR U21659 ( .A(n22700), .B(p_input[240]), .Z(n21672) );
  XOR U21660 ( .A(n21675), .B(n21674), .Z(n21673) );
  NOR U21661 ( .A(n22702), .B(p_input[238]), .Z(n21674) );
  XOR U21662 ( .A(n21677), .B(n21676), .Z(n21675) );
  NOR U21663 ( .A(n22704), .B(p_input[236]), .Z(n21676) );
  XOR U21664 ( .A(n21679), .B(n21678), .Z(n21677) );
  NOR U21665 ( .A(n22706), .B(p_input[234]), .Z(n21678) );
  XOR U21666 ( .A(n21681), .B(n21680), .Z(n21679) );
  NOR U21667 ( .A(n22708), .B(p_input[232]), .Z(n21680) );
  XOR U21668 ( .A(n21683), .B(n21682), .Z(n21681) );
  NOR U21669 ( .A(n22710), .B(p_input[230]), .Z(n21682) );
  XOR U21670 ( .A(n21685), .B(n21684), .Z(n21683) );
  NOR U21671 ( .A(n22712), .B(p_input[228]), .Z(n21684) );
  XOR U21672 ( .A(n21687), .B(n21686), .Z(n21685) );
  NOR U21673 ( .A(n22714), .B(p_input[226]), .Z(n21686) );
  XOR U21674 ( .A(n21689), .B(n21688), .Z(n21687) );
  NOR U21675 ( .A(n22716), .B(p_input[224]), .Z(n21688) );
  XOR U21676 ( .A(n21691), .B(n21690), .Z(n21689) );
  NOR U21677 ( .A(n22718), .B(p_input[222]), .Z(n21690) );
  XOR U21678 ( .A(n21693), .B(n21692), .Z(n21691) );
  NOR U21679 ( .A(n22720), .B(p_input[220]), .Z(n21692) );
  XOR U21680 ( .A(n21695), .B(n21694), .Z(n21693) );
  NOR U21681 ( .A(n22722), .B(p_input[218]), .Z(n21694) );
  XOR U21682 ( .A(n21697), .B(n21696), .Z(n21695) );
  NOR U21683 ( .A(n22724), .B(p_input[216]), .Z(n21696) );
  XOR U21684 ( .A(n21699), .B(n21698), .Z(n21697) );
  NOR U21685 ( .A(n22726), .B(p_input[214]), .Z(n21698) );
  XOR U21686 ( .A(n21701), .B(n21700), .Z(n21699) );
  NOR U21687 ( .A(n22728), .B(p_input[212]), .Z(n21700) );
  XOR U21688 ( .A(n21703), .B(n21702), .Z(n21701) );
  NOR U21689 ( .A(n22730), .B(p_input[210]), .Z(n21702) );
  XOR U21690 ( .A(n21705), .B(n21704), .Z(n21703) );
  NOR U21691 ( .A(n22732), .B(p_input[208]), .Z(n21704) );
  XOR U21692 ( .A(n21707), .B(n21706), .Z(n21705) );
  NOR U21693 ( .A(n22734), .B(p_input[206]), .Z(n21706) );
  XOR U21694 ( .A(n21709), .B(n21708), .Z(n21707) );
  NOR U21695 ( .A(n22736), .B(p_input[204]), .Z(n21708) );
  XOR U21696 ( .A(n21711), .B(n21710), .Z(n21709) );
  NOR U21697 ( .A(n22738), .B(p_input[202]), .Z(n21710) );
  XOR U21698 ( .A(n21713), .B(n21712), .Z(n21711) );
  NOR U21699 ( .A(n22740), .B(p_input[200]), .Z(n21712) );
  XOR U21700 ( .A(n21715), .B(n21714), .Z(n21713) );
  NOR U21701 ( .A(n22742), .B(p_input[198]), .Z(n21714) );
  XOR U21702 ( .A(n21717), .B(n21716), .Z(n21715) );
  NOR U21703 ( .A(n22744), .B(p_input[196]), .Z(n21716) );
  XOR U21704 ( .A(n21719), .B(n21718), .Z(n21717) );
  NOR U21705 ( .A(n22746), .B(p_input[194]), .Z(n21718) );
  XOR U21706 ( .A(n21721), .B(n21720), .Z(n21719) );
  NOR U21707 ( .A(n22748), .B(p_input[192]), .Z(n21720) );
  XOR U21708 ( .A(n21723), .B(n21722), .Z(n21721) );
  NOR U21709 ( .A(n22750), .B(p_input[190]), .Z(n21722) );
  XOR U21710 ( .A(n21725), .B(n21724), .Z(n21723) );
  NOR U21711 ( .A(n22752), .B(p_input[188]), .Z(n21724) );
  XOR U21712 ( .A(n21727), .B(n21726), .Z(n21725) );
  NOR U21713 ( .A(n22754), .B(p_input[186]), .Z(n21726) );
  XOR U21714 ( .A(n21729), .B(n21728), .Z(n21727) );
  NOR U21715 ( .A(n22756), .B(p_input[184]), .Z(n21728) );
  XOR U21716 ( .A(n21731), .B(n21730), .Z(n21729) );
  NOR U21717 ( .A(n22758), .B(p_input[182]), .Z(n21730) );
  XOR U21718 ( .A(n21733), .B(n21732), .Z(n21731) );
  NOR U21719 ( .A(n22760), .B(p_input[180]), .Z(n21732) );
  XOR U21720 ( .A(n21735), .B(n21734), .Z(n21733) );
  NOR U21721 ( .A(n22762), .B(p_input[178]), .Z(n21734) );
  XOR U21722 ( .A(n21737), .B(n21736), .Z(n21735) );
  NOR U21723 ( .A(n22764), .B(p_input[176]), .Z(n21736) );
  XOR U21724 ( .A(n21739), .B(n21738), .Z(n21737) );
  NOR U21725 ( .A(n22766), .B(p_input[174]), .Z(n21738) );
  XOR U21726 ( .A(n21741), .B(n21740), .Z(n21739) );
  NOR U21727 ( .A(n22768), .B(p_input[172]), .Z(n21740) );
  XOR U21728 ( .A(n21743), .B(n21742), .Z(n21741) );
  NOR U21729 ( .A(n22770), .B(p_input[170]), .Z(n21742) );
  XOR U21730 ( .A(n21745), .B(n21744), .Z(n21743) );
  NOR U21731 ( .A(n22772), .B(p_input[168]), .Z(n21744) );
  XOR U21732 ( .A(n21747), .B(n21746), .Z(n21745) );
  NOR U21733 ( .A(n22774), .B(p_input[166]), .Z(n21746) );
  XOR U21734 ( .A(n21749), .B(n21748), .Z(n21747) );
  NOR U21735 ( .A(n22776), .B(p_input[164]), .Z(n21748) );
  XOR U21736 ( .A(n21751), .B(n21750), .Z(n21749) );
  NOR U21737 ( .A(n22778), .B(p_input[162]), .Z(n21750) );
  XOR U21738 ( .A(n21753), .B(n21752), .Z(n21751) );
  NOR U21739 ( .A(n22780), .B(p_input[160]), .Z(n21752) );
  XOR U21740 ( .A(n21755), .B(n21754), .Z(n21753) );
  NOR U21741 ( .A(n22782), .B(p_input[158]), .Z(n21754) );
  XOR U21742 ( .A(n21757), .B(n21756), .Z(n21755) );
  NOR U21743 ( .A(n22784), .B(p_input[156]), .Z(n21756) );
  XOR U21744 ( .A(n21759), .B(n21758), .Z(n21757) );
  NOR U21745 ( .A(n22786), .B(p_input[154]), .Z(n21758) );
  XOR U21746 ( .A(n21761), .B(n21760), .Z(n21759) );
  NOR U21747 ( .A(n22788), .B(p_input[152]), .Z(n21760) );
  XOR U21748 ( .A(n21763), .B(n21762), .Z(n21761) );
  NOR U21749 ( .A(n22790), .B(p_input[150]), .Z(n21762) );
  XOR U21750 ( .A(n21765), .B(n21764), .Z(n21763) );
  NOR U21751 ( .A(n22792), .B(p_input[148]), .Z(n21764) );
  XOR U21752 ( .A(n21767), .B(n21766), .Z(n21765) );
  NOR U21753 ( .A(n22794), .B(p_input[146]), .Z(n21766) );
  XOR U21754 ( .A(n21769), .B(n21768), .Z(n21767) );
  NOR U21755 ( .A(n22796), .B(p_input[144]), .Z(n21768) );
  XOR U21756 ( .A(n21771), .B(n21770), .Z(n21769) );
  NOR U21757 ( .A(n22798), .B(p_input[142]), .Z(n21770) );
  XOR U21758 ( .A(n21773), .B(n21772), .Z(n21771) );
  NOR U21759 ( .A(n22800), .B(p_input[140]), .Z(n21772) );
  XOR U21760 ( .A(n21775), .B(n21774), .Z(n21773) );
  NOR U21761 ( .A(n22802), .B(p_input[138]), .Z(n21774) );
  XOR U21762 ( .A(n21777), .B(n21776), .Z(n21775) );
  NOR U21763 ( .A(n22804), .B(p_input[136]), .Z(n21776) );
  XOR U21764 ( .A(n21779), .B(n21778), .Z(n21777) );
  NOR U21765 ( .A(n22806), .B(p_input[134]), .Z(n21778) );
  XOR U21766 ( .A(n21781), .B(n21780), .Z(n21779) );
  NOR U21767 ( .A(n22808), .B(p_input[132]), .Z(n21780) );
  XOR U21768 ( .A(n21783), .B(n21782), .Z(n21781) );
  NOR U21769 ( .A(n22810), .B(p_input[130]), .Z(n21782) );
  XOR U21770 ( .A(n21785), .B(n21784), .Z(n21783) );
  NOR U21771 ( .A(n22812), .B(p_input[128]), .Z(n21784) );
  XOR U21772 ( .A(n21787), .B(n21786), .Z(n21785) );
  NOR U21773 ( .A(n22814), .B(p_input[126]), .Z(n21786) );
  XOR U21774 ( .A(n21789), .B(n21788), .Z(n21787) );
  NOR U21775 ( .A(n22816), .B(p_input[124]), .Z(n21788) );
  XOR U21776 ( .A(n21791), .B(n21790), .Z(n21789) );
  NOR U21777 ( .A(n22818), .B(p_input[122]), .Z(n21790) );
  XOR U21778 ( .A(n21793), .B(n21792), .Z(n21791) );
  NOR U21779 ( .A(n22820), .B(p_input[120]), .Z(n21792) );
  XOR U21780 ( .A(n21795), .B(n21794), .Z(n21793) );
  NOR U21781 ( .A(n22822), .B(p_input[118]), .Z(n21794) );
  XOR U21782 ( .A(n21797), .B(n21796), .Z(n21795) );
  NOR U21783 ( .A(n22824), .B(p_input[116]), .Z(n21796) );
  XOR U21784 ( .A(n21799), .B(n21798), .Z(n21797) );
  NOR U21785 ( .A(n22826), .B(p_input[114]), .Z(n21798) );
  XOR U21786 ( .A(n21801), .B(n21800), .Z(n21799) );
  NOR U21787 ( .A(n22828), .B(p_input[112]), .Z(n21800) );
  XOR U21788 ( .A(n21803), .B(n21802), .Z(n21801) );
  NOR U21789 ( .A(n22830), .B(p_input[110]), .Z(n21802) );
  XOR U21790 ( .A(n21805), .B(n21804), .Z(n21803) );
  NOR U21791 ( .A(n22832), .B(p_input[108]), .Z(n21804) );
  XOR U21792 ( .A(n21807), .B(n21806), .Z(n21805) );
  NOR U21793 ( .A(n22834), .B(p_input[106]), .Z(n21806) );
  XOR U21794 ( .A(n21809), .B(n21808), .Z(n21807) );
  NOR U21795 ( .A(n22836), .B(p_input[104]), .Z(n21808) );
  XOR U21796 ( .A(n21811), .B(n21810), .Z(n21809) );
  NOR U21797 ( .A(n22838), .B(p_input[102]), .Z(n21810) );
  XOR U21798 ( .A(n21813), .B(n21812), .Z(n21811) );
  NOR U21799 ( .A(n22840), .B(p_input[100]), .Z(n21812) );
  XOR U21800 ( .A(n21815), .B(n21814), .Z(n21813) );
  NOR U21801 ( .A(n22842), .B(p_input[98]), .Z(n21814) );
  XOR U21802 ( .A(n21817), .B(n21816), .Z(n21815) );
  NOR U21803 ( .A(n22844), .B(p_input[96]), .Z(n21816) );
  XOR U21804 ( .A(n21819), .B(n21818), .Z(n21817) );
  NOR U21805 ( .A(n22846), .B(p_input[94]), .Z(n21818) );
  XOR U21806 ( .A(n21821), .B(n21820), .Z(n21819) );
  NOR U21807 ( .A(n22848), .B(p_input[92]), .Z(n21820) );
  XOR U21808 ( .A(n21823), .B(n21822), .Z(n21821) );
  NOR U21809 ( .A(n22850), .B(p_input[90]), .Z(n21822) );
  XOR U21810 ( .A(n21825), .B(n21824), .Z(n21823) );
  NOR U21811 ( .A(n22852), .B(p_input[88]), .Z(n21824) );
  XOR U21812 ( .A(n21827), .B(n21826), .Z(n21825) );
  NOR U21813 ( .A(n22854), .B(p_input[86]), .Z(n21826) );
  XOR U21814 ( .A(n21829), .B(n21828), .Z(n21827) );
  NOR U21815 ( .A(n22856), .B(p_input[84]), .Z(n21828) );
  XOR U21816 ( .A(n21831), .B(n21830), .Z(n21829) );
  NOR U21817 ( .A(n22858), .B(p_input[82]), .Z(n21830) );
  XOR U21818 ( .A(n21833), .B(n21832), .Z(n21831) );
  NOR U21819 ( .A(n22860), .B(p_input[80]), .Z(n21832) );
  XOR U21820 ( .A(n21835), .B(n21834), .Z(n21833) );
  NOR U21821 ( .A(n22862), .B(p_input[78]), .Z(n21834) );
  XOR U21822 ( .A(n21837), .B(n21836), .Z(n21835) );
  NOR U21823 ( .A(n22864), .B(p_input[76]), .Z(n21836) );
  XOR U21824 ( .A(n21839), .B(n21838), .Z(n21837) );
  NOR U21825 ( .A(n22866), .B(p_input[74]), .Z(n21838) );
  XOR U21826 ( .A(n21841), .B(n21840), .Z(n21839) );
  NOR U21827 ( .A(n22868), .B(p_input[72]), .Z(n21840) );
  XOR U21828 ( .A(n21843), .B(n21842), .Z(n21841) );
  NOR U21829 ( .A(n22870), .B(p_input[70]), .Z(n21842) );
  XOR U21830 ( .A(n21845), .B(n21844), .Z(n21843) );
  NOR U21831 ( .A(n22872), .B(p_input[68]), .Z(n21844) );
  XOR U21832 ( .A(n21847), .B(n21846), .Z(n21845) );
  NOR U21833 ( .A(n22874), .B(p_input[66]), .Z(n21846) );
  XOR U21834 ( .A(n21849), .B(n21848), .Z(n21847) );
  NOR U21835 ( .A(n22876), .B(p_input[64]), .Z(n21848) );
  XOR U21836 ( .A(n21851), .B(n21850), .Z(n21849) );
  NOR U21837 ( .A(n22878), .B(p_input[62]), .Z(n21850) );
  XOR U21838 ( .A(n21853), .B(n21852), .Z(n21851) );
  NOR U21839 ( .A(n22880), .B(p_input[60]), .Z(n21852) );
  XOR U21840 ( .A(n21855), .B(n21854), .Z(n21853) );
  NOR U21841 ( .A(n22882), .B(p_input[58]), .Z(n21854) );
  XOR U21842 ( .A(n21857), .B(n21856), .Z(n21855) );
  NOR U21843 ( .A(n22884), .B(p_input[56]), .Z(n21856) );
  XOR U21844 ( .A(n21859), .B(n21858), .Z(n21857) );
  NOR U21845 ( .A(n22886), .B(p_input[54]), .Z(n21858) );
  XOR U21846 ( .A(n21861), .B(n21860), .Z(n21859) );
  NOR U21847 ( .A(n22888), .B(p_input[52]), .Z(n21860) );
  XOR U21848 ( .A(n21863), .B(n21862), .Z(n21861) );
  NOR U21849 ( .A(n22890), .B(p_input[50]), .Z(n21862) );
  XOR U21850 ( .A(n21865), .B(n21864), .Z(n21863) );
  NOR U21851 ( .A(n22892), .B(p_input[48]), .Z(n21864) );
  XOR U21852 ( .A(n21867), .B(n21866), .Z(n21865) );
  NOR U21853 ( .A(n22894), .B(p_input[46]), .Z(n21866) );
  XOR U21854 ( .A(n21869), .B(n21868), .Z(n21867) );
  NOR U21855 ( .A(n22896), .B(p_input[44]), .Z(n21868) );
  XOR U21856 ( .A(n21871), .B(n21870), .Z(n21869) );
  NOR U21857 ( .A(n22898), .B(p_input[42]), .Z(n21870) );
  XOR U21858 ( .A(n21873), .B(n21872), .Z(n21871) );
  NOR U21859 ( .A(n22900), .B(p_input[40]), .Z(n21872) );
  XOR U21860 ( .A(n21875), .B(n21874), .Z(n21873) );
  NOR U21861 ( .A(n22902), .B(p_input[38]), .Z(n21874) );
  XOR U21862 ( .A(n21877), .B(n21876), .Z(n21875) );
  NOR U21863 ( .A(n22904), .B(p_input[36]), .Z(n21876) );
  XOR U21864 ( .A(n21879), .B(n21878), .Z(n21877) );
  NOR U21865 ( .A(n22906), .B(p_input[34]), .Z(n21878) );
  XOR U21866 ( .A(n21881), .B(n21880), .Z(n21879) );
  NOR U21867 ( .A(n22908), .B(p_input[32]), .Z(n21880) );
  XOR U21868 ( .A(n21883), .B(n21882), .Z(n21881) );
  NOR U21869 ( .A(n22910), .B(p_input[30]), .Z(n21882) );
  XOR U21870 ( .A(n21885), .B(n21884), .Z(n21883) );
  NOR U21871 ( .A(n22912), .B(p_input[28]), .Z(n21884) );
  XOR U21872 ( .A(n21887), .B(n21886), .Z(n21885) );
  NOR U21873 ( .A(n22914), .B(p_input[26]), .Z(n21886) );
  XOR U21874 ( .A(n21889), .B(n21888), .Z(n21887) );
  NOR U21875 ( .A(n22916), .B(p_input[24]), .Z(n21888) );
  XOR U21876 ( .A(n21891), .B(n21890), .Z(n21889) );
  NOR U21877 ( .A(n22918), .B(p_input[22]), .Z(n21890) );
  XOR U21878 ( .A(n21893), .B(n21892), .Z(n21891) );
  NOR U21879 ( .A(n22920), .B(p_input[20]), .Z(n21892) );
  XOR U21880 ( .A(n21895), .B(n21894), .Z(n21893) );
  NOR U21881 ( .A(n22922), .B(p_input[18]), .Z(n21894) );
  XOR U21882 ( .A(n21897), .B(n21896), .Z(n21895) );
  NOR U21883 ( .A(n22924), .B(p_input[16]), .Z(n21896) );
  XOR U21884 ( .A(n21899), .B(n21898), .Z(n21897) );
  NOR U21885 ( .A(n22926), .B(p_input[14]), .Z(n21898) );
  XOR U21886 ( .A(n21901), .B(n21900), .Z(n21899) );
  NOR U21887 ( .A(n22928), .B(p_input[12]), .Z(n21900) );
  XOR U21888 ( .A(n21915), .B(n21914), .Z(n21901) );
  NOR U21889 ( .A(n22930), .B(p_input[10]), .Z(n21914) );
  XOR U21890 ( .A(n21917), .B(n21916), .Z(n21915) );
  NOR U21891 ( .A(n22932), .B(p_input[8]), .Z(n21916) );
  XOR U21892 ( .A(n21905), .B(n21904), .Z(n21917) );
  NOR U21893 ( .A(n22934), .B(p_input[6]), .Z(n21904) );
  XOR U21894 ( .A(n21912), .B(n21913), .Z(n21905) );
  XOR U21895 ( .A(n21910), .B(n21911), .Z(n21913) );
  NOR U21896 ( .A(n22936), .B(p_input[2]), .Z(n21911) );
  NOR U21897 ( .A(n22938), .B(p_input[0]), .Z(n21910) );
  NOR U21898 ( .A(n22940), .B(p_input[4]), .Z(n21912) );
  XNOR U21899 ( .A(n22942), .B(n22943), .Z(n140) );
  AND U21900 ( .A(n1), .B(n22944), .Z(n22943) );
  XNOR U21901 ( .A(n22942), .B(n22945), .Z(n22944) );
  XNOR U21902 ( .A(n22946), .B(n22947), .Z(n1) );
  AND U21903 ( .A(n22948), .B(n22949), .Z(n22947) );
  XNOR U21904 ( .A(n22946), .B(n19), .Z(n22949) );
  XNOR U21905 ( .A(n22950), .B(n22951), .Z(n19) );
  AND U21906 ( .A(n22952), .B(n22953), .Z(n22951) );
  XOR U21907 ( .A(n34), .B(n22950), .Z(n22952) );
  XOR U21908 ( .A(n22954), .B(n22955), .Z(n22950) );
  AND U21909 ( .A(n34), .B(n22954), .Z(n22955) );
  XOR U21910 ( .A(n16), .B(n22946), .Z(n22948) );
  IV U21911 ( .A(n20), .Z(n16) );
  XOR U21912 ( .A(n22956), .B(n22957), .Z(n20) );
  AND U21913 ( .A(n22958), .B(n22959), .Z(n22957) );
  XOR U21914 ( .A(n35), .B(n22956), .Z(n22958) );
  XOR U21915 ( .A(n22960), .B(n22961), .Z(n22956) );
  NOR U21916 ( .A(n31), .B(n22962), .Z(n22961) );
  IV U21917 ( .A(n22960), .Z(n22962) );
  XOR U21918 ( .A(n22963), .B(n22964), .Z(n22946) );
  AND U21919 ( .A(n22965), .B(n22966), .Z(n22964) );
  XOR U21920 ( .A(n22963), .B(n34), .Z(n22966) );
  XOR U21921 ( .A(n22954), .B(n22953), .Z(n34) );
  XNOR U21922 ( .A(n22967), .B(n22968), .Z(n22953) );
  XOR U21923 ( .A(n22969), .B(n22970), .Z(n22968) );
  XOR U21924 ( .A(n22971), .B(n22972), .Z(n22970) );
  NOR U21925 ( .A(n22973), .B(n22974), .Z(n22971) );
  XOR U21926 ( .A(n22975), .B(n22976), .Z(n22969) );
  NOR U21927 ( .A(n22977), .B(n22978), .Z(n22976) );
  NOR U21928 ( .A(n22979), .B(n22980), .Z(n22975) );
  XOR U21929 ( .A(n22981), .B(n22982), .Z(n22967) );
  XOR U21930 ( .A(n22974), .B(n22978), .Z(n22982) );
  XNOR U21931 ( .A(n22983), .B(n22980), .Z(n22981) );
  XOR U21932 ( .A(n22984), .B(n22985), .Z(n22983) );
  XOR U21933 ( .A(n22986), .B(n22987), .Z(n22985) );
  XOR U21934 ( .A(n22988), .B(n22989), .Z(n22987) );
  XOR U21935 ( .A(n22990), .B(n22991), .Z(n22986) );
  NOR U21936 ( .A(n22992), .B(n22993), .Z(n22991) );
  AND U21937 ( .A(n22994), .B(n22972), .Z(n22990) );
  XOR U21938 ( .A(n22995), .B(n22996), .Z(n22984) );
  XOR U21939 ( .A(n22997), .B(n22998), .Z(n22996) );
  XOR U21940 ( .A(n22999), .B(n23000), .Z(n22998) );
  XOR U21941 ( .A(n23001), .B(n23002), .Z(n23000) );
  XOR U21942 ( .A(n23003), .B(n23004), .Z(n23002) );
  XOR U21943 ( .A(n23005), .B(n23006), .Z(n23004) );
  XNOR U21944 ( .A(n23007), .B(n23008), .Z(n23003) );
  XNOR U21945 ( .A(n23009), .B(n23010), .Z(n23008) );
  NOR U21946 ( .A(n23011), .B(n23006), .Z(n23009) );
  XOR U21947 ( .A(n23012), .B(n23013), .Z(n23001) );
  XOR U21948 ( .A(n23014), .B(n23015), .Z(n23013) );
  XNOR U21949 ( .A(n23016), .B(n23017), .Z(n23015) );
  XOR U21950 ( .A(n23018), .B(n23019), .Z(n23017) );
  XOR U21951 ( .A(n23020), .B(n23021), .Z(n23019) );
  XOR U21952 ( .A(n23022), .B(n23023), .Z(n23021) );
  XOR U21953 ( .A(n23024), .B(n23025), .Z(n23020) );
  XOR U21954 ( .A(n23026), .B(n23027), .Z(n23025) );
  XOR U21955 ( .A(n23028), .B(n23029), .Z(n23027) );
  XOR U21956 ( .A(n23030), .B(n23031), .Z(n23029) );
  XOR U21957 ( .A(n23032), .B(n23033), .Z(n23031) );
  XNOR U21958 ( .A(n23034), .B(n23035), .Z(n23030) );
  XNOR U21959 ( .A(n23036), .B(n23037), .Z(n23035) );
  NOR U21960 ( .A(n23038), .B(n23033), .Z(n23036) );
  XOR U21961 ( .A(n23039), .B(n23040), .Z(n23028) );
  XOR U21962 ( .A(n23041), .B(n23042), .Z(n23040) );
  XNOR U21963 ( .A(n23043), .B(n23044), .Z(n23042) );
  XOR U21964 ( .A(n23045), .B(n23046), .Z(n23044) );
  XOR U21965 ( .A(n23047), .B(n23048), .Z(n23046) );
  XOR U21966 ( .A(n23049), .B(n23050), .Z(n23048) );
  XOR U21967 ( .A(n23051), .B(n23052), .Z(n23047) );
  XOR U21968 ( .A(n23053), .B(n23054), .Z(n23052) );
  XOR U21969 ( .A(n23055), .B(n23056), .Z(n23054) );
  XOR U21970 ( .A(n23057), .B(n23058), .Z(n23056) );
  XOR U21971 ( .A(n23059), .B(n23060), .Z(n23058) );
  XNOR U21972 ( .A(n23061), .B(n23062), .Z(n23057) );
  XNOR U21973 ( .A(n23063), .B(n23064), .Z(n23062) );
  NOR U21974 ( .A(n23065), .B(n23060), .Z(n23063) );
  XOR U21975 ( .A(n23066), .B(n23067), .Z(n23055) );
  XOR U21976 ( .A(n23068), .B(n23069), .Z(n23067) );
  XNOR U21977 ( .A(n23070), .B(n23071), .Z(n23069) );
  XOR U21978 ( .A(n23072), .B(n23073), .Z(n23071) );
  XOR U21979 ( .A(n23074), .B(n23075), .Z(n23073) );
  XOR U21980 ( .A(n23076), .B(n23077), .Z(n23075) );
  XOR U21981 ( .A(n23078), .B(n23079), .Z(n23074) );
  XOR U21982 ( .A(n23080), .B(n23081), .Z(n23079) );
  XOR U21983 ( .A(n23082), .B(n23083), .Z(n23081) );
  XOR U21984 ( .A(n23084), .B(n23085), .Z(n23083) );
  XOR U21985 ( .A(n23086), .B(n23087), .Z(n23085) );
  XNOR U21986 ( .A(n23088), .B(n23089), .Z(n23084) );
  XNOR U21987 ( .A(n23090), .B(n23091), .Z(n23089) );
  NOR U21988 ( .A(n23092), .B(n23087), .Z(n23090) );
  XOR U21989 ( .A(n23093), .B(n23094), .Z(n23082) );
  XOR U21990 ( .A(n23095), .B(n23096), .Z(n23094) );
  XNOR U21991 ( .A(n23097), .B(n23098), .Z(n23096) );
  XOR U21992 ( .A(n23099), .B(n23100), .Z(n23098) );
  XOR U21993 ( .A(n23101), .B(n23102), .Z(n23100) );
  XOR U21994 ( .A(n23103), .B(n23104), .Z(n23102) );
  XOR U21995 ( .A(n23105), .B(n23106), .Z(n23101) );
  XOR U21996 ( .A(n23107), .B(n23108), .Z(n23106) );
  XOR U21997 ( .A(n23109), .B(n23110), .Z(n23108) );
  XOR U21998 ( .A(n23111), .B(n23112), .Z(n23110) );
  XOR U21999 ( .A(n23113), .B(n23114), .Z(n23112) );
  XNOR U22000 ( .A(n23115), .B(n23116), .Z(n23111) );
  XNOR U22001 ( .A(n23117), .B(n23118), .Z(n23116) );
  NOR U22002 ( .A(n23119), .B(n23114), .Z(n23117) );
  XOR U22003 ( .A(n23120), .B(n23121), .Z(n23109) );
  XOR U22004 ( .A(n23122), .B(n23123), .Z(n23121) );
  XNOR U22005 ( .A(n23124), .B(n23125), .Z(n23123) );
  XOR U22006 ( .A(n23126), .B(n23127), .Z(n23125) );
  XOR U22007 ( .A(n23128), .B(n23129), .Z(n23127) );
  XOR U22008 ( .A(n23130), .B(n23131), .Z(n23129) );
  XOR U22009 ( .A(n23132), .B(n23133), .Z(n23128) );
  XOR U22010 ( .A(n23134), .B(n23135), .Z(n23133) );
  XOR U22011 ( .A(n23136), .B(n23137), .Z(n23135) );
  XOR U22012 ( .A(n23138), .B(n23139), .Z(n23137) );
  XOR U22013 ( .A(n23140), .B(n23141), .Z(n23139) );
  XNOR U22014 ( .A(n23142), .B(n23143), .Z(n23138) );
  XNOR U22015 ( .A(n23144), .B(n23145), .Z(n23143) );
  NOR U22016 ( .A(n23146), .B(n23141), .Z(n23144) );
  XOR U22017 ( .A(n23147), .B(n23148), .Z(n23136) );
  XOR U22018 ( .A(n23149), .B(n23150), .Z(n23148) );
  XNOR U22019 ( .A(n23151), .B(n23152), .Z(n23150) );
  XOR U22020 ( .A(n23153), .B(n23154), .Z(n23152) );
  XOR U22021 ( .A(n23155), .B(n23156), .Z(n23154) );
  XOR U22022 ( .A(n23157), .B(n23158), .Z(n23156) );
  XOR U22023 ( .A(n23159), .B(n23160), .Z(n23155) );
  XOR U22024 ( .A(n23161), .B(n23162), .Z(n23160) );
  XOR U22025 ( .A(n23163), .B(n23164), .Z(n23162) );
  XOR U22026 ( .A(n23165), .B(n23166), .Z(n23164) );
  XOR U22027 ( .A(n23167), .B(n23168), .Z(n23166) );
  XNOR U22028 ( .A(n23169), .B(n23170), .Z(n23165) );
  XNOR U22029 ( .A(n23171), .B(n23172), .Z(n23170) );
  NOR U22030 ( .A(n23173), .B(n23168), .Z(n23171) );
  XOR U22031 ( .A(n23174), .B(n23175), .Z(n23163) );
  XOR U22032 ( .A(n23176), .B(n23177), .Z(n23175) );
  XNOR U22033 ( .A(n23178), .B(n23179), .Z(n23177) );
  XOR U22034 ( .A(n23180), .B(n23181), .Z(n23179) );
  XOR U22035 ( .A(n23182), .B(n23183), .Z(n23181) );
  XOR U22036 ( .A(n23184), .B(n23185), .Z(n23183) );
  XOR U22037 ( .A(n23186), .B(n23187), .Z(n23182) );
  XOR U22038 ( .A(n23188), .B(n23189), .Z(n23187) );
  XOR U22039 ( .A(n23190), .B(n23191), .Z(n23189) );
  XOR U22040 ( .A(n23192), .B(n23193), .Z(n23191) );
  XOR U22041 ( .A(n23194), .B(n23195), .Z(n23193) );
  XNOR U22042 ( .A(n23196), .B(n23197), .Z(n23192) );
  XNOR U22043 ( .A(n23198), .B(n23199), .Z(n23197) );
  NOR U22044 ( .A(n23200), .B(n23195), .Z(n23198) );
  XOR U22045 ( .A(n23201), .B(n23202), .Z(n23190) );
  XOR U22046 ( .A(n23203), .B(n23204), .Z(n23202) );
  XNOR U22047 ( .A(n23205), .B(n23206), .Z(n23204) );
  XOR U22048 ( .A(n23207), .B(n23208), .Z(n23206) );
  XOR U22049 ( .A(n23209), .B(n23210), .Z(n23208) );
  XOR U22050 ( .A(n23211), .B(n23212), .Z(n23210) );
  XOR U22051 ( .A(n23213), .B(n23214), .Z(n23209) );
  XOR U22052 ( .A(n23215), .B(n23216), .Z(n23214) );
  XOR U22053 ( .A(n23217), .B(n23218), .Z(n23216) );
  XOR U22054 ( .A(n23219), .B(n23220), .Z(n23218) );
  XOR U22055 ( .A(n23221), .B(n23222), .Z(n23220) );
  XNOR U22056 ( .A(n23223), .B(n23224), .Z(n23219) );
  XNOR U22057 ( .A(n23225), .B(n23226), .Z(n23224) );
  NOR U22058 ( .A(n23227), .B(n23222), .Z(n23225) );
  XOR U22059 ( .A(n23228), .B(n23229), .Z(n23217) );
  XOR U22060 ( .A(n23230), .B(n23231), .Z(n23229) );
  XNOR U22061 ( .A(n23232), .B(n23233), .Z(n23231) );
  XOR U22062 ( .A(n23234), .B(n23235), .Z(n23233) );
  XOR U22063 ( .A(n23236), .B(n23237), .Z(n23235) );
  XOR U22064 ( .A(n23238), .B(n23239), .Z(n23237) );
  XOR U22065 ( .A(n23240), .B(n23241), .Z(n23236) );
  XOR U22066 ( .A(n23242), .B(n23243), .Z(n23241) );
  XOR U22067 ( .A(n23244), .B(n23245), .Z(n23243) );
  XOR U22068 ( .A(n23246), .B(n23247), .Z(n23245) );
  XOR U22069 ( .A(n23248), .B(n23249), .Z(n23247) );
  XNOR U22070 ( .A(n23250), .B(n23251), .Z(n23246) );
  XNOR U22071 ( .A(n23252), .B(n23253), .Z(n23251) );
  NOR U22072 ( .A(n23254), .B(n23249), .Z(n23252) );
  XOR U22073 ( .A(n23255), .B(n23256), .Z(n23244) );
  XOR U22074 ( .A(n23257), .B(n23258), .Z(n23256) );
  XNOR U22075 ( .A(n23259), .B(n23260), .Z(n23258) );
  XOR U22076 ( .A(n23261), .B(n23262), .Z(n23260) );
  XOR U22077 ( .A(n23263), .B(n23264), .Z(n23262) );
  XOR U22078 ( .A(n23265), .B(n23266), .Z(n23264) );
  XOR U22079 ( .A(n23267), .B(n23268), .Z(n23263) );
  XOR U22080 ( .A(n23269), .B(n23270), .Z(n23268) );
  XOR U22081 ( .A(n23271), .B(n23272), .Z(n23270) );
  XOR U22082 ( .A(n23273), .B(n23274), .Z(n23272) );
  XOR U22083 ( .A(n23275), .B(n23276), .Z(n23274) );
  XNOR U22084 ( .A(n23277), .B(n23278), .Z(n23273) );
  XNOR U22085 ( .A(n23279), .B(n23280), .Z(n23278) );
  NOR U22086 ( .A(n23281), .B(n23276), .Z(n23279) );
  XOR U22087 ( .A(n23282), .B(n23283), .Z(n23271) );
  XOR U22088 ( .A(n23284), .B(n23285), .Z(n23283) );
  XNOR U22089 ( .A(n23286), .B(n23287), .Z(n23285) );
  XOR U22090 ( .A(n23288), .B(n23289), .Z(n23287) );
  XOR U22091 ( .A(n23290), .B(n23291), .Z(n23289) );
  XOR U22092 ( .A(n23292), .B(n23293), .Z(n23291) );
  XOR U22093 ( .A(n23294), .B(n23295), .Z(n23290) );
  XOR U22094 ( .A(n23296), .B(n23297), .Z(n23295) );
  XOR U22095 ( .A(n23298), .B(n23299), .Z(n23297) );
  XOR U22096 ( .A(n23300), .B(n23301), .Z(n23299) );
  XOR U22097 ( .A(n23302), .B(n23303), .Z(n23301) );
  XNOR U22098 ( .A(n23304), .B(n23305), .Z(n23300) );
  XNOR U22099 ( .A(n23306), .B(n23307), .Z(n23305) );
  NOR U22100 ( .A(n23308), .B(n23303), .Z(n23306) );
  XOR U22101 ( .A(n23309), .B(n23310), .Z(n23298) );
  XOR U22102 ( .A(n23311), .B(n23312), .Z(n23310) );
  XNOR U22103 ( .A(n23313), .B(n23314), .Z(n23312) );
  XOR U22104 ( .A(n23315), .B(n23316), .Z(n23314) );
  XOR U22105 ( .A(n23317), .B(n23318), .Z(n23316) );
  XOR U22106 ( .A(n23319), .B(n23320), .Z(n23318) );
  XOR U22107 ( .A(n23321), .B(n23322), .Z(n23317) );
  XOR U22108 ( .A(n23323), .B(n23324), .Z(n23322) );
  XOR U22109 ( .A(n23325), .B(n23326), .Z(n23324) );
  XOR U22110 ( .A(n23327), .B(n23328), .Z(n23326) );
  XOR U22111 ( .A(n23329), .B(n23330), .Z(n23328) );
  XNOR U22112 ( .A(n23331), .B(n23332), .Z(n23327) );
  XNOR U22113 ( .A(n23333), .B(n23334), .Z(n23332) );
  NOR U22114 ( .A(n23335), .B(n23330), .Z(n23333) );
  XOR U22115 ( .A(n23336), .B(n23337), .Z(n23325) );
  XOR U22116 ( .A(n23338), .B(n23339), .Z(n23337) );
  XNOR U22117 ( .A(n23340), .B(n23341), .Z(n23339) );
  XOR U22118 ( .A(n23342), .B(n23343), .Z(n23341) );
  XOR U22119 ( .A(n23344), .B(n23345), .Z(n23343) );
  XOR U22120 ( .A(n23346), .B(n23347), .Z(n23345) );
  XOR U22121 ( .A(n23348), .B(n23349), .Z(n23344) );
  XOR U22122 ( .A(n23350), .B(n23351), .Z(n23349) );
  XOR U22123 ( .A(n23352), .B(n23353), .Z(n23351) );
  XOR U22124 ( .A(n23354), .B(n23355), .Z(n23353) );
  XOR U22125 ( .A(n23356), .B(n23357), .Z(n23355) );
  XNOR U22126 ( .A(n23358), .B(n23359), .Z(n23354) );
  XNOR U22127 ( .A(n23360), .B(n23361), .Z(n23359) );
  NOR U22128 ( .A(n23362), .B(n23357), .Z(n23360) );
  XOR U22129 ( .A(n23363), .B(n23364), .Z(n23352) );
  XOR U22130 ( .A(n23365), .B(n23366), .Z(n23364) );
  XNOR U22131 ( .A(n23367), .B(n23368), .Z(n23366) );
  XOR U22132 ( .A(n23369), .B(n23370), .Z(n23368) );
  XOR U22133 ( .A(n23371), .B(n23372), .Z(n23370) );
  XOR U22134 ( .A(n23373), .B(n23374), .Z(n23372) );
  XOR U22135 ( .A(n23375), .B(n23376), .Z(n23371) );
  XOR U22136 ( .A(n23377), .B(n23378), .Z(n23376) );
  XOR U22137 ( .A(n23379), .B(n23380), .Z(n23378) );
  XOR U22138 ( .A(n23381), .B(n23382), .Z(n23380) );
  XOR U22139 ( .A(n23383), .B(n23384), .Z(n23382) );
  XNOR U22140 ( .A(n23385), .B(n23386), .Z(n23381) );
  XNOR U22141 ( .A(n23387), .B(n23388), .Z(n23386) );
  NOR U22142 ( .A(n23389), .B(n23384), .Z(n23387) );
  XOR U22143 ( .A(n23390), .B(n23391), .Z(n23379) );
  XOR U22144 ( .A(n23392), .B(n23393), .Z(n23391) );
  XNOR U22145 ( .A(n23394), .B(n23395), .Z(n23393) );
  XOR U22146 ( .A(n23396), .B(n23397), .Z(n23395) );
  XOR U22147 ( .A(n23398), .B(n23399), .Z(n23397) );
  XOR U22148 ( .A(n23400), .B(n23401), .Z(n23399) );
  XOR U22149 ( .A(n23402), .B(n23403), .Z(n23398) );
  XOR U22150 ( .A(n23404), .B(n23405), .Z(n23403) );
  XOR U22151 ( .A(n23406), .B(n23407), .Z(n23405) );
  XOR U22152 ( .A(n23408), .B(n23409), .Z(n23407) );
  XOR U22153 ( .A(n23410), .B(n23411), .Z(n23409) );
  XNOR U22154 ( .A(n23412), .B(n23413), .Z(n23408) );
  XNOR U22155 ( .A(n23414), .B(n23415), .Z(n23413) );
  NOR U22156 ( .A(n23416), .B(n23411), .Z(n23414) );
  XOR U22157 ( .A(n23417), .B(n23418), .Z(n23406) );
  XOR U22158 ( .A(n23419), .B(n23420), .Z(n23418) );
  XNOR U22159 ( .A(n23421), .B(n23422), .Z(n23420) );
  XOR U22160 ( .A(n23423), .B(n23424), .Z(n23422) );
  XOR U22161 ( .A(n23425), .B(n23426), .Z(n23424) );
  XOR U22162 ( .A(n23427), .B(n23428), .Z(n23426) );
  XOR U22163 ( .A(n23429), .B(n23430), .Z(n23425) );
  XOR U22164 ( .A(n23431), .B(n23432), .Z(n23430) );
  XOR U22165 ( .A(n23433), .B(n23434), .Z(n23432) );
  XOR U22166 ( .A(n23435), .B(n23436), .Z(n23434) );
  XOR U22167 ( .A(n23437), .B(n23438), .Z(n23436) );
  XNOR U22168 ( .A(n23439), .B(n23440), .Z(n23435) );
  XNOR U22169 ( .A(n23441), .B(n23442), .Z(n23440) );
  NOR U22170 ( .A(n23443), .B(n23438), .Z(n23441) );
  XOR U22171 ( .A(n23444), .B(n23445), .Z(n23433) );
  XOR U22172 ( .A(n23446), .B(n23447), .Z(n23445) );
  XNOR U22173 ( .A(n23448), .B(n23449), .Z(n23447) );
  XOR U22174 ( .A(n23450), .B(n23451), .Z(n23449) );
  XOR U22175 ( .A(n23452), .B(n23453), .Z(n23451) );
  XOR U22176 ( .A(n23454), .B(n23455), .Z(n23453) );
  XOR U22177 ( .A(n23456), .B(n23457), .Z(n23452) );
  XOR U22178 ( .A(n23458), .B(n23459), .Z(n23457) );
  XOR U22179 ( .A(n23460), .B(n23461), .Z(n23459) );
  XOR U22180 ( .A(n23462), .B(n23463), .Z(n23461) );
  XOR U22181 ( .A(n23464), .B(n23465), .Z(n23463) );
  XNOR U22182 ( .A(n23466), .B(n23467), .Z(n23462) );
  XNOR U22183 ( .A(n23468), .B(n23469), .Z(n23467) );
  NOR U22184 ( .A(n23470), .B(n23465), .Z(n23468) );
  XOR U22185 ( .A(n23471), .B(n23472), .Z(n23460) );
  XOR U22186 ( .A(n23473), .B(n23474), .Z(n23472) );
  XNOR U22187 ( .A(n23475), .B(n23476), .Z(n23474) );
  XOR U22188 ( .A(n23477), .B(n23478), .Z(n23476) );
  XOR U22189 ( .A(n23479), .B(n23480), .Z(n23478) );
  XOR U22190 ( .A(n23481), .B(n23482), .Z(n23480) );
  XOR U22191 ( .A(n23483), .B(n23484), .Z(n23479) );
  XOR U22192 ( .A(n23485), .B(n23486), .Z(n23484) );
  XOR U22193 ( .A(n23487), .B(n23488), .Z(n23486) );
  XOR U22194 ( .A(n23489), .B(n23490), .Z(n23488) );
  XOR U22195 ( .A(n23491), .B(n23492), .Z(n23490) );
  XNOR U22196 ( .A(n23493), .B(n23494), .Z(n23489) );
  XNOR U22197 ( .A(n23495), .B(n23496), .Z(n23494) );
  NOR U22198 ( .A(n23497), .B(n23492), .Z(n23495) );
  XOR U22199 ( .A(n23498), .B(n23499), .Z(n23487) );
  XOR U22200 ( .A(n23500), .B(n23501), .Z(n23499) );
  XNOR U22201 ( .A(n23502), .B(n23503), .Z(n23501) );
  XOR U22202 ( .A(n23504), .B(n23505), .Z(n23503) );
  XOR U22203 ( .A(n23506), .B(n23507), .Z(n23505) );
  XOR U22204 ( .A(n23508), .B(n23509), .Z(n23507) );
  XOR U22205 ( .A(n23510), .B(n23511), .Z(n23506) );
  XOR U22206 ( .A(n23512), .B(n23513), .Z(n23511) );
  XOR U22207 ( .A(n23514), .B(n23515), .Z(n23513) );
  XOR U22208 ( .A(n23516), .B(n23517), .Z(n23515) );
  XOR U22209 ( .A(n23518), .B(n23519), .Z(n23517) );
  XNOR U22210 ( .A(n23520), .B(n23521), .Z(n23516) );
  XNOR U22211 ( .A(n23522), .B(n23523), .Z(n23521) );
  NOR U22212 ( .A(n23524), .B(n23519), .Z(n23522) );
  XOR U22213 ( .A(n23525), .B(n23526), .Z(n23514) );
  XOR U22214 ( .A(n23527), .B(n23528), .Z(n23526) );
  XNOR U22215 ( .A(n23529), .B(n23530), .Z(n23528) );
  XOR U22216 ( .A(n23531), .B(n23532), .Z(n23530) );
  XOR U22217 ( .A(n23533), .B(n23534), .Z(n23532) );
  XOR U22218 ( .A(n23535), .B(n23536), .Z(n23534) );
  XOR U22219 ( .A(n23537), .B(n23538), .Z(n23533) );
  XOR U22220 ( .A(n23539), .B(n23540), .Z(n23538) );
  XOR U22221 ( .A(n23541), .B(n23542), .Z(n23540) );
  XOR U22222 ( .A(n23543), .B(n23544), .Z(n23542) );
  XOR U22223 ( .A(n23545), .B(n23546), .Z(n23544) );
  XNOR U22224 ( .A(n23547), .B(n23548), .Z(n23543) );
  XNOR U22225 ( .A(n23549), .B(n23550), .Z(n23548) );
  NOR U22226 ( .A(n23551), .B(n23546), .Z(n23549) );
  XOR U22227 ( .A(n23552), .B(n23553), .Z(n23541) );
  XOR U22228 ( .A(n23554), .B(n23555), .Z(n23553) );
  XOR U22229 ( .A(n23556), .B(n23557), .Z(n23555) );
  XOR U22230 ( .A(n23558), .B(n23559), .Z(n23554) );
  XOR U22231 ( .A(n23560), .B(n23561), .Z(n23552) );
  XOR U22232 ( .A(n23562), .B(n23563), .Z(n23561) );
  AND U22233 ( .A(n23564), .B(n23565), .Z(n23563) );
  XOR U22234 ( .A(n23566), .B(n23557), .Z(n23564) );
  XOR U22235 ( .A(n23567), .B(n23568), .Z(n23557) );
  NOR U22236 ( .A(n23566), .B(n23567), .Z(n23568) );
  NOR U22237 ( .A(n23569), .B(n23558), .Z(n23562) );
  XOR U22238 ( .A(n23570), .B(n23571), .Z(n23560) );
  NOR U22239 ( .A(n23572), .B(n23559), .Z(n23571) );
  NOR U22240 ( .A(n23573), .B(n23556), .Z(n23570) );
  XOR U22241 ( .A(n23574), .B(n23575), .Z(n23539) );
  NOR U22242 ( .A(n23576), .B(n23550), .Z(n23575) );
  NOR U22243 ( .A(n23577), .B(n23547), .Z(n23574) );
  XOR U22244 ( .A(n23578), .B(n23579), .Z(n23537) );
  XOR U22245 ( .A(n23580), .B(n23581), .Z(n23579) );
  NOR U22246 ( .A(n23582), .B(n23545), .Z(n23581) );
  NOR U22247 ( .A(n23583), .B(n23584), .Z(n23580) );
  XOR U22248 ( .A(n23585), .B(n23586), .Z(n23578) );
  NOR U22249 ( .A(n23587), .B(n23588), .Z(n23586) );
  NOR U22250 ( .A(n23589), .B(n23535), .Z(n23585) );
  XOR U22251 ( .A(n23590), .B(n23591), .Z(n23531) );
  XOR U22252 ( .A(n23584), .B(n23588), .Z(n23591) );
  XOR U22253 ( .A(n23592), .B(n23593), .Z(n23590) );
  NOR U22254 ( .A(n23594), .B(n23536), .Z(n23593) );
  NOR U22255 ( .A(n23595), .B(n23596), .Z(n23592) );
  XOR U22256 ( .A(n23597), .B(n23598), .Z(n23527) );
  XOR U22257 ( .A(n23599), .B(n23600), .Z(n23525) );
  XNOR U22258 ( .A(n23601), .B(n23596), .Z(n23600) );
  NOR U22259 ( .A(n23602), .B(n23597), .Z(n23601) );
  XOR U22260 ( .A(n23603), .B(n23604), .Z(n23599) );
  NOR U22261 ( .A(n23605), .B(n23598), .Z(n23604) );
  NOR U22262 ( .A(n23606), .B(n23529), .Z(n23603) );
  XOR U22263 ( .A(n23607), .B(n23608), .Z(n23512) );
  NOR U22264 ( .A(n23609), .B(n23523), .Z(n23608) );
  NOR U22265 ( .A(n23610), .B(n23520), .Z(n23607) );
  XOR U22266 ( .A(n23611), .B(n23612), .Z(n23510) );
  XOR U22267 ( .A(n23613), .B(n23614), .Z(n23612) );
  NOR U22268 ( .A(n23615), .B(n23518), .Z(n23614) );
  NOR U22269 ( .A(n23616), .B(n23617), .Z(n23613) );
  XOR U22270 ( .A(n23618), .B(n23619), .Z(n23611) );
  NOR U22271 ( .A(n23620), .B(n23621), .Z(n23619) );
  NOR U22272 ( .A(n23622), .B(n23508), .Z(n23618) );
  XOR U22273 ( .A(n23623), .B(n23624), .Z(n23504) );
  XOR U22274 ( .A(n23617), .B(n23621), .Z(n23624) );
  XOR U22275 ( .A(n23625), .B(n23626), .Z(n23623) );
  NOR U22276 ( .A(n23627), .B(n23509), .Z(n23626) );
  NOR U22277 ( .A(n23628), .B(n23629), .Z(n23625) );
  XOR U22278 ( .A(n23630), .B(n23631), .Z(n23500) );
  XOR U22279 ( .A(n23632), .B(n23633), .Z(n23498) );
  XNOR U22280 ( .A(n23634), .B(n23629), .Z(n23633) );
  NOR U22281 ( .A(n23635), .B(n23630), .Z(n23634) );
  XOR U22282 ( .A(n23636), .B(n23637), .Z(n23632) );
  NOR U22283 ( .A(n23638), .B(n23631), .Z(n23637) );
  NOR U22284 ( .A(n23639), .B(n23502), .Z(n23636) );
  XOR U22285 ( .A(n23640), .B(n23641), .Z(n23485) );
  NOR U22286 ( .A(n23642), .B(n23496), .Z(n23641) );
  NOR U22287 ( .A(n23643), .B(n23493), .Z(n23640) );
  XOR U22288 ( .A(n23644), .B(n23645), .Z(n23483) );
  XOR U22289 ( .A(n23646), .B(n23647), .Z(n23645) );
  NOR U22290 ( .A(n23648), .B(n23491), .Z(n23647) );
  NOR U22291 ( .A(n23649), .B(n23650), .Z(n23646) );
  XOR U22292 ( .A(n23651), .B(n23652), .Z(n23644) );
  NOR U22293 ( .A(n23653), .B(n23654), .Z(n23652) );
  NOR U22294 ( .A(n23655), .B(n23481), .Z(n23651) );
  XOR U22295 ( .A(n23656), .B(n23657), .Z(n23477) );
  XOR U22296 ( .A(n23650), .B(n23654), .Z(n23657) );
  XOR U22297 ( .A(n23658), .B(n23659), .Z(n23656) );
  NOR U22298 ( .A(n23660), .B(n23482), .Z(n23659) );
  NOR U22299 ( .A(n23661), .B(n23662), .Z(n23658) );
  XOR U22300 ( .A(n23663), .B(n23664), .Z(n23473) );
  XOR U22301 ( .A(n23665), .B(n23666), .Z(n23471) );
  XNOR U22302 ( .A(n23667), .B(n23662), .Z(n23666) );
  NOR U22303 ( .A(n23668), .B(n23663), .Z(n23667) );
  XOR U22304 ( .A(n23669), .B(n23670), .Z(n23665) );
  NOR U22305 ( .A(n23671), .B(n23664), .Z(n23670) );
  NOR U22306 ( .A(n23672), .B(n23475), .Z(n23669) );
  XOR U22307 ( .A(n23673), .B(n23674), .Z(n23458) );
  NOR U22308 ( .A(n23675), .B(n23469), .Z(n23674) );
  NOR U22309 ( .A(n23676), .B(n23466), .Z(n23673) );
  XOR U22310 ( .A(n23677), .B(n23678), .Z(n23456) );
  XOR U22311 ( .A(n23679), .B(n23680), .Z(n23678) );
  NOR U22312 ( .A(n23681), .B(n23464), .Z(n23680) );
  NOR U22313 ( .A(n23682), .B(n23683), .Z(n23679) );
  XOR U22314 ( .A(n23684), .B(n23685), .Z(n23677) );
  NOR U22315 ( .A(n23686), .B(n23687), .Z(n23685) );
  NOR U22316 ( .A(n23688), .B(n23454), .Z(n23684) );
  XOR U22317 ( .A(n23689), .B(n23690), .Z(n23450) );
  XOR U22318 ( .A(n23683), .B(n23687), .Z(n23690) );
  XOR U22319 ( .A(n23691), .B(n23692), .Z(n23689) );
  NOR U22320 ( .A(n23693), .B(n23455), .Z(n23692) );
  NOR U22321 ( .A(n23694), .B(n23695), .Z(n23691) );
  XOR U22322 ( .A(n23696), .B(n23697), .Z(n23446) );
  XOR U22323 ( .A(n23698), .B(n23699), .Z(n23444) );
  XNOR U22324 ( .A(n23700), .B(n23695), .Z(n23699) );
  NOR U22325 ( .A(n23701), .B(n23696), .Z(n23700) );
  XOR U22326 ( .A(n23702), .B(n23703), .Z(n23698) );
  NOR U22327 ( .A(n23704), .B(n23697), .Z(n23703) );
  NOR U22328 ( .A(n23705), .B(n23448), .Z(n23702) );
  XOR U22329 ( .A(n23706), .B(n23707), .Z(n23431) );
  NOR U22330 ( .A(n23708), .B(n23442), .Z(n23707) );
  NOR U22331 ( .A(n23709), .B(n23439), .Z(n23706) );
  XOR U22332 ( .A(n23710), .B(n23711), .Z(n23429) );
  XOR U22333 ( .A(n23712), .B(n23713), .Z(n23711) );
  NOR U22334 ( .A(n23714), .B(n23437), .Z(n23713) );
  NOR U22335 ( .A(n23715), .B(n23716), .Z(n23712) );
  XOR U22336 ( .A(n23717), .B(n23718), .Z(n23710) );
  NOR U22337 ( .A(n23719), .B(n23720), .Z(n23718) );
  NOR U22338 ( .A(n23721), .B(n23427), .Z(n23717) );
  XOR U22339 ( .A(n23722), .B(n23723), .Z(n23423) );
  XOR U22340 ( .A(n23716), .B(n23720), .Z(n23723) );
  XOR U22341 ( .A(n23724), .B(n23725), .Z(n23722) );
  NOR U22342 ( .A(n23726), .B(n23428), .Z(n23725) );
  NOR U22343 ( .A(n23727), .B(n23728), .Z(n23724) );
  XOR U22344 ( .A(n23729), .B(n23730), .Z(n23419) );
  XOR U22345 ( .A(n23731), .B(n23732), .Z(n23417) );
  XNOR U22346 ( .A(n23733), .B(n23728), .Z(n23732) );
  NOR U22347 ( .A(n23734), .B(n23729), .Z(n23733) );
  XOR U22348 ( .A(n23735), .B(n23736), .Z(n23731) );
  NOR U22349 ( .A(n23737), .B(n23730), .Z(n23736) );
  NOR U22350 ( .A(n23738), .B(n23421), .Z(n23735) );
  XOR U22351 ( .A(n23739), .B(n23740), .Z(n23404) );
  NOR U22352 ( .A(n23741), .B(n23415), .Z(n23740) );
  NOR U22353 ( .A(n23742), .B(n23412), .Z(n23739) );
  XOR U22354 ( .A(n23743), .B(n23744), .Z(n23402) );
  XOR U22355 ( .A(n23745), .B(n23746), .Z(n23744) );
  NOR U22356 ( .A(n23747), .B(n23410), .Z(n23746) );
  NOR U22357 ( .A(n23748), .B(n23749), .Z(n23745) );
  XOR U22358 ( .A(n23750), .B(n23751), .Z(n23743) );
  NOR U22359 ( .A(n23752), .B(n23753), .Z(n23751) );
  NOR U22360 ( .A(n23754), .B(n23400), .Z(n23750) );
  XOR U22361 ( .A(n23755), .B(n23756), .Z(n23396) );
  XOR U22362 ( .A(n23749), .B(n23753), .Z(n23756) );
  XOR U22363 ( .A(n23757), .B(n23758), .Z(n23755) );
  NOR U22364 ( .A(n23759), .B(n23401), .Z(n23758) );
  NOR U22365 ( .A(n23760), .B(n23761), .Z(n23757) );
  XOR U22366 ( .A(n23762), .B(n23763), .Z(n23392) );
  XOR U22367 ( .A(n23764), .B(n23765), .Z(n23390) );
  XNOR U22368 ( .A(n23766), .B(n23761), .Z(n23765) );
  NOR U22369 ( .A(n23767), .B(n23762), .Z(n23766) );
  XOR U22370 ( .A(n23768), .B(n23769), .Z(n23764) );
  NOR U22371 ( .A(n23770), .B(n23763), .Z(n23769) );
  NOR U22372 ( .A(n23771), .B(n23394), .Z(n23768) );
  XOR U22373 ( .A(n23772), .B(n23773), .Z(n23377) );
  NOR U22374 ( .A(n23774), .B(n23388), .Z(n23773) );
  NOR U22375 ( .A(n23775), .B(n23385), .Z(n23772) );
  XOR U22376 ( .A(n23776), .B(n23777), .Z(n23375) );
  XOR U22377 ( .A(n23778), .B(n23779), .Z(n23777) );
  NOR U22378 ( .A(n23780), .B(n23383), .Z(n23779) );
  NOR U22379 ( .A(n23781), .B(n23782), .Z(n23778) );
  XOR U22380 ( .A(n23783), .B(n23784), .Z(n23776) );
  NOR U22381 ( .A(n23785), .B(n23786), .Z(n23784) );
  NOR U22382 ( .A(n23787), .B(n23373), .Z(n23783) );
  XOR U22383 ( .A(n23788), .B(n23789), .Z(n23369) );
  XOR U22384 ( .A(n23782), .B(n23786), .Z(n23789) );
  XOR U22385 ( .A(n23790), .B(n23791), .Z(n23788) );
  NOR U22386 ( .A(n23792), .B(n23374), .Z(n23791) );
  NOR U22387 ( .A(n23793), .B(n23794), .Z(n23790) );
  XOR U22388 ( .A(n23795), .B(n23796), .Z(n23365) );
  XOR U22389 ( .A(n23797), .B(n23798), .Z(n23363) );
  XNOR U22390 ( .A(n23799), .B(n23794), .Z(n23798) );
  NOR U22391 ( .A(n23800), .B(n23795), .Z(n23799) );
  XOR U22392 ( .A(n23801), .B(n23802), .Z(n23797) );
  NOR U22393 ( .A(n23803), .B(n23796), .Z(n23802) );
  NOR U22394 ( .A(n23804), .B(n23367), .Z(n23801) );
  XOR U22395 ( .A(n23805), .B(n23806), .Z(n23350) );
  NOR U22396 ( .A(n23807), .B(n23361), .Z(n23806) );
  NOR U22397 ( .A(n23808), .B(n23358), .Z(n23805) );
  XOR U22398 ( .A(n23809), .B(n23810), .Z(n23348) );
  XOR U22399 ( .A(n23811), .B(n23812), .Z(n23810) );
  NOR U22400 ( .A(n23813), .B(n23356), .Z(n23812) );
  NOR U22401 ( .A(n23814), .B(n23815), .Z(n23811) );
  XOR U22402 ( .A(n23816), .B(n23817), .Z(n23809) );
  NOR U22403 ( .A(n23818), .B(n23819), .Z(n23817) );
  NOR U22404 ( .A(n23820), .B(n23346), .Z(n23816) );
  XOR U22405 ( .A(n23821), .B(n23822), .Z(n23342) );
  XOR U22406 ( .A(n23815), .B(n23819), .Z(n23822) );
  XOR U22407 ( .A(n23823), .B(n23824), .Z(n23821) );
  NOR U22408 ( .A(n23825), .B(n23347), .Z(n23824) );
  NOR U22409 ( .A(n23826), .B(n23827), .Z(n23823) );
  XOR U22410 ( .A(n23828), .B(n23829), .Z(n23338) );
  XOR U22411 ( .A(n23830), .B(n23831), .Z(n23336) );
  XNOR U22412 ( .A(n23832), .B(n23827), .Z(n23831) );
  NOR U22413 ( .A(n23833), .B(n23828), .Z(n23832) );
  XOR U22414 ( .A(n23834), .B(n23835), .Z(n23830) );
  NOR U22415 ( .A(n23836), .B(n23829), .Z(n23835) );
  NOR U22416 ( .A(n23837), .B(n23340), .Z(n23834) );
  XOR U22417 ( .A(n23838), .B(n23839), .Z(n23323) );
  NOR U22418 ( .A(n23840), .B(n23334), .Z(n23839) );
  NOR U22419 ( .A(n23841), .B(n23331), .Z(n23838) );
  XOR U22420 ( .A(n23842), .B(n23843), .Z(n23321) );
  XOR U22421 ( .A(n23844), .B(n23845), .Z(n23843) );
  NOR U22422 ( .A(n23846), .B(n23329), .Z(n23845) );
  NOR U22423 ( .A(n23847), .B(n23848), .Z(n23844) );
  XOR U22424 ( .A(n23849), .B(n23850), .Z(n23842) );
  NOR U22425 ( .A(n23851), .B(n23852), .Z(n23850) );
  NOR U22426 ( .A(n23853), .B(n23319), .Z(n23849) );
  XOR U22427 ( .A(n23854), .B(n23855), .Z(n23315) );
  XOR U22428 ( .A(n23848), .B(n23852), .Z(n23855) );
  XOR U22429 ( .A(n23856), .B(n23857), .Z(n23854) );
  NOR U22430 ( .A(n23858), .B(n23320), .Z(n23857) );
  NOR U22431 ( .A(n23859), .B(n23860), .Z(n23856) );
  XOR U22432 ( .A(n23861), .B(n23862), .Z(n23311) );
  XOR U22433 ( .A(n23863), .B(n23864), .Z(n23309) );
  XNOR U22434 ( .A(n23865), .B(n23860), .Z(n23864) );
  NOR U22435 ( .A(n23866), .B(n23861), .Z(n23865) );
  XOR U22436 ( .A(n23867), .B(n23868), .Z(n23863) );
  NOR U22437 ( .A(n23869), .B(n23862), .Z(n23868) );
  NOR U22438 ( .A(n23870), .B(n23313), .Z(n23867) );
  XOR U22439 ( .A(n23871), .B(n23872), .Z(n23296) );
  NOR U22440 ( .A(n23873), .B(n23307), .Z(n23872) );
  NOR U22441 ( .A(n23874), .B(n23304), .Z(n23871) );
  XOR U22442 ( .A(n23875), .B(n23876), .Z(n23294) );
  XOR U22443 ( .A(n23877), .B(n23878), .Z(n23876) );
  NOR U22444 ( .A(n23879), .B(n23302), .Z(n23878) );
  NOR U22445 ( .A(n23880), .B(n23881), .Z(n23877) );
  XOR U22446 ( .A(n23882), .B(n23883), .Z(n23875) );
  NOR U22447 ( .A(n23884), .B(n23885), .Z(n23883) );
  NOR U22448 ( .A(n23886), .B(n23292), .Z(n23882) );
  XOR U22449 ( .A(n23887), .B(n23888), .Z(n23288) );
  XOR U22450 ( .A(n23881), .B(n23885), .Z(n23888) );
  XOR U22451 ( .A(n23889), .B(n23890), .Z(n23887) );
  NOR U22452 ( .A(n23891), .B(n23293), .Z(n23890) );
  NOR U22453 ( .A(n23892), .B(n23893), .Z(n23889) );
  XOR U22454 ( .A(n23894), .B(n23895), .Z(n23284) );
  XOR U22455 ( .A(n23896), .B(n23897), .Z(n23282) );
  XNOR U22456 ( .A(n23898), .B(n23893), .Z(n23897) );
  NOR U22457 ( .A(n23899), .B(n23894), .Z(n23898) );
  XOR U22458 ( .A(n23900), .B(n23901), .Z(n23896) );
  NOR U22459 ( .A(n23902), .B(n23895), .Z(n23901) );
  NOR U22460 ( .A(n23903), .B(n23286), .Z(n23900) );
  XOR U22461 ( .A(n23904), .B(n23905), .Z(n23269) );
  NOR U22462 ( .A(n23906), .B(n23280), .Z(n23905) );
  NOR U22463 ( .A(n23907), .B(n23277), .Z(n23904) );
  XOR U22464 ( .A(n23908), .B(n23909), .Z(n23267) );
  XOR U22465 ( .A(n23910), .B(n23911), .Z(n23909) );
  NOR U22466 ( .A(n23912), .B(n23275), .Z(n23911) );
  NOR U22467 ( .A(n23913), .B(n23914), .Z(n23910) );
  XOR U22468 ( .A(n23915), .B(n23916), .Z(n23908) );
  NOR U22469 ( .A(n23917), .B(n23918), .Z(n23916) );
  NOR U22470 ( .A(n23919), .B(n23265), .Z(n23915) );
  XOR U22471 ( .A(n23920), .B(n23921), .Z(n23261) );
  XOR U22472 ( .A(n23914), .B(n23918), .Z(n23921) );
  XOR U22473 ( .A(n23922), .B(n23923), .Z(n23920) );
  NOR U22474 ( .A(n23924), .B(n23266), .Z(n23923) );
  NOR U22475 ( .A(n23925), .B(n23926), .Z(n23922) );
  XOR U22476 ( .A(n23927), .B(n23928), .Z(n23257) );
  XOR U22477 ( .A(n23929), .B(n23930), .Z(n23255) );
  XNOR U22478 ( .A(n23931), .B(n23926), .Z(n23930) );
  NOR U22479 ( .A(n23932), .B(n23927), .Z(n23931) );
  XOR U22480 ( .A(n23933), .B(n23934), .Z(n23929) );
  NOR U22481 ( .A(n23935), .B(n23928), .Z(n23934) );
  NOR U22482 ( .A(n23936), .B(n23259), .Z(n23933) );
  XOR U22483 ( .A(n23937), .B(n23938), .Z(n23242) );
  NOR U22484 ( .A(n23939), .B(n23253), .Z(n23938) );
  NOR U22485 ( .A(n23940), .B(n23250), .Z(n23937) );
  XOR U22486 ( .A(n23941), .B(n23942), .Z(n23240) );
  XOR U22487 ( .A(n23943), .B(n23944), .Z(n23942) );
  NOR U22488 ( .A(n23945), .B(n23248), .Z(n23944) );
  NOR U22489 ( .A(n23946), .B(n23947), .Z(n23943) );
  XOR U22490 ( .A(n23948), .B(n23949), .Z(n23941) );
  NOR U22491 ( .A(n23950), .B(n23951), .Z(n23949) );
  NOR U22492 ( .A(n23952), .B(n23238), .Z(n23948) );
  XOR U22493 ( .A(n23953), .B(n23954), .Z(n23234) );
  XOR U22494 ( .A(n23947), .B(n23951), .Z(n23954) );
  XOR U22495 ( .A(n23955), .B(n23956), .Z(n23953) );
  NOR U22496 ( .A(n23957), .B(n23239), .Z(n23956) );
  NOR U22497 ( .A(n23958), .B(n23959), .Z(n23955) );
  XOR U22498 ( .A(n23960), .B(n23961), .Z(n23230) );
  XOR U22499 ( .A(n23962), .B(n23963), .Z(n23228) );
  XNOR U22500 ( .A(n23964), .B(n23959), .Z(n23963) );
  NOR U22501 ( .A(n23965), .B(n23960), .Z(n23964) );
  XOR U22502 ( .A(n23966), .B(n23967), .Z(n23962) );
  NOR U22503 ( .A(n23968), .B(n23961), .Z(n23967) );
  NOR U22504 ( .A(n23969), .B(n23232), .Z(n23966) );
  XOR U22505 ( .A(n23970), .B(n23971), .Z(n23215) );
  NOR U22506 ( .A(n23972), .B(n23226), .Z(n23971) );
  NOR U22507 ( .A(n23973), .B(n23223), .Z(n23970) );
  XOR U22508 ( .A(n23974), .B(n23975), .Z(n23213) );
  XOR U22509 ( .A(n23976), .B(n23977), .Z(n23975) );
  NOR U22510 ( .A(n23978), .B(n23221), .Z(n23977) );
  NOR U22511 ( .A(n23979), .B(n23980), .Z(n23976) );
  XOR U22512 ( .A(n23981), .B(n23982), .Z(n23974) );
  NOR U22513 ( .A(n23983), .B(n23984), .Z(n23982) );
  NOR U22514 ( .A(n23985), .B(n23211), .Z(n23981) );
  XOR U22515 ( .A(n23986), .B(n23987), .Z(n23207) );
  XOR U22516 ( .A(n23980), .B(n23984), .Z(n23987) );
  XOR U22517 ( .A(n23988), .B(n23989), .Z(n23986) );
  NOR U22518 ( .A(n23990), .B(n23212), .Z(n23989) );
  NOR U22519 ( .A(n23991), .B(n23992), .Z(n23988) );
  XOR U22520 ( .A(n23993), .B(n23994), .Z(n23203) );
  XOR U22521 ( .A(n23995), .B(n23996), .Z(n23201) );
  XNOR U22522 ( .A(n23997), .B(n23992), .Z(n23996) );
  NOR U22523 ( .A(n23998), .B(n23993), .Z(n23997) );
  XOR U22524 ( .A(n23999), .B(n24000), .Z(n23995) );
  NOR U22525 ( .A(n24001), .B(n23994), .Z(n24000) );
  NOR U22526 ( .A(n24002), .B(n23205), .Z(n23999) );
  XOR U22527 ( .A(n24003), .B(n24004), .Z(n23188) );
  NOR U22528 ( .A(n24005), .B(n23199), .Z(n24004) );
  NOR U22529 ( .A(n24006), .B(n23196), .Z(n24003) );
  XOR U22530 ( .A(n24007), .B(n24008), .Z(n23186) );
  XOR U22531 ( .A(n24009), .B(n24010), .Z(n24008) );
  NOR U22532 ( .A(n24011), .B(n23194), .Z(n24010) );
  NOR U22533 ( .A(n24012), .B(n24013), .Z(n24009) );
  XOR U22534 ( .A(n24014), .B(n24015), .Z(n24007) );
  NOR U22535 ( .A(n24016), .B(n24017), .Z(n24015) );
  NOR U22536 ( .A(n24018), .B(n23184), .Z(n24014) );
  XOR U22537 ( .A(n24019), .B(n24020), .Z(n23180) );
  XOR U22538 ( .A(n24013), .B(n24017), .Z(n24020) );
  XOR U22539 ( .A(n24021), .B(n24022), .Z(n24019) );
  NOR U22540 ( .A(n24023), .B(n23185), .Z(n24022) );
  NOR U22541 ( .A(n24024), .B(n24025), .Z(n24021) );
  XOR U22542 ( .A(n24026), .B(n24027), .Z(n23176) );
  XOR U22543 ( .A(n24028), .B(n24029), .Z(n23174) );
  XNOR U22544 ( .A(n24030), .B(n24025), .Z(n24029) );
  NOR U22545 ( .A(n24031), .B(n24026), .Z(n24030) );
  XOR U22546 ( .A(n24032), .B(n24033), .Z(n24028) );
  NOR U22547 ( .A(n24034), .B(n24027), .Z(n24033) );
  NOR U22548 ( .A(n24035), .B(n23178), .Z(n24032) );
  XOR U22549 ( .A(n24036), .B(n24037), .Z(n23161) );
  NOR U22550 ( .A(n24038), .B(n23172), .Z(n24037) );
  NOR U22551 ( .A(n24039), .B(n23169), .Z(n24036) );
  XOR U22552 ( .A(n24040), .B(n24041), .Z(n23159) );
  XOR U22553 ( .A(n24042), .B(n24043), .Z(n24041) );
  NOR U22554 ( .A(n24044), .B(n23167), .Z(n24043) );
  NOR U22555 ( .A(n24045), .B(n24046), .Z(n24042) );
  XOR U22556 ( .A(n24047), .B(n24048), .Z(n24040) );
  NOR U22557 ( .A(n24049), .B(n24050), .Z(n24048) );
  NOR U22558 ( .A(n24051), .B(n23157), .Z(n24047) );
  XOR U22559 ( .A(n24052), .B(n24053), .Z(n23153) );
  XOR U22560 ( .A(n24046), .B(n24050), .Z(n24053) );
  XOR U22561 ( .A(n24054), .B(n24055), .Z(n24052) );
  NOR U22562 ( .A(n24056), .B(n23158), .Z(n24055) );
  NOR U22563 ( .A(n24057), .B(n24058), .Z(n24054) );
  XOR U22564 ( .A(n24059), .B(n24060), .Z(n23149) );
  XOR U22565 ( .A(n24061), .B(n24062), .Z(n23147) );
  XNOR U22566 ( .A(n24063), .B(n24058), .Z(n24062) );
  NOR U22567 ( .A(n24064), .B(n24059), .Z(n24063) );
  XOR U22568 ( .A(n24065), .B(n24066), .Z(n24061) );
  NOR U22569 ( .A(n24067), .B(n24060), .Z(n24066) );
  NOR U22570 ( .A(n24068), .B(n23151), .Z(n24065) );
  XOR U22571 ( .A(n24069), .B(n24070), .Z(n23134) );
  NOR U22572 ( .A(n24071), .B(n23145), .Z(n24070) );
  NOR U22573 ( .A(n24072), .B(n23142), .Z(n24069) );
  XOR U22574 ( .A(n24073), .B(n24074), .Z(n23132) );
  XOR U22575 ( .A(n24075), .B(n24076), .Z(n24074) );
  NOR U22576 ( .A(n24077), .B(n23140), .Z(n24076) );
  NOR U22577 ( .A(n24078), .B(n24079), .Z(n24075) );
  XOR U22578 ( .A(n24080), .B(n24081), .Z(n24073) );
  NOR U22579 ( .A(n24082), .B(n24083), .Z(n24081) );
  NOR U22580 ( .A(n24084), .B(n23130), .Z(n24080) );
  XOR U22581 ( .A(n24085), .B(n24086), .Z(n23126) );
  XOR U22582 ( .A(n24079), .B(n24083), .Z(n24086) );
  XOR U22583 ( .A(n24087), .B(n24088), .Z(n24085) );
  NOR U22584 ( .A(n24089), .B(n23131), .Z(n24088) );
  NOR U22585 ( .A(n24090), .B(n24091), .Z(n24087) );
  XOR U22586 ( .A(n24092), .B(n24093), .Z(n23122) );
  XOR U22587 ( .A(n24094), .B(n24095), .Z(n23120) );
  XNOR U22588 ( .A(n24096), .B(n24091), .Z(n24095) );
  NOR U22589 ( .A(n24097), .B(n24092), .Z(n24096) );
  XOR U22590 ( .A(n24098), .B(n24099), .Z(n24094) );
  NOR U22591 ( .A(n24100), .B(n24093), .Z(n24099) );
  NOR U22592 ( .A(n24101), .B(n23124), .Z(n24098) );
  XOR U22593 ( .A(n24102), .B(n24103), .Z(n23107) );
  NOR U22594 ( .A(n24104), .B(n23118), .Z(n24103) );
  NOR U22595 ( .A(n24105), .B(n23115), .Z(n24102) );
  XOR U22596 ( .A(n24106), .B(n24107), .Z(n23105) );
  XOR U22597 ( .A(n24108), .B(n24109), .Z(n24107) );
  NOR U22598 ( .A(n24110), .B(n23113), .Z(n24109) );
  NOR U22599 ( .A(n24111), .B(n24112), .Z(n24108) );
  XOR U22600 ( .A(n24113), .B(n24114), .Z(n24106) );
  NOR U22601 ( .A(n24115), .B(n24116), .Z(n24114) );
  NOR U22602 ( .A(n24117), .B(n23103), .Z(n24113) );
  XOR U22603 ( .A(n24118), .B(n24119), .Z(n23099) );
  XOR U22604 ( .A(n24112), .B(n24116), .Z(n24119) );
  XOR U22605 ( .A(n24120), .B(n24121), .Z(n24118) );
  NOR U22606 ( .A(n24122), .B(n23104), .Z(n24121) );
  NOR U22607 ( .A(n24123), .B(n24124), .Z(n24120) );
  XOR U22608 ( .A(n24125), .B(n24126), .Z(n23095) );
  XOR U22609 ( .A(n24127), .B(n24128), .Z(n23093) );
  XNOR U22610 ( .A(n24129), .B(n24124), .Z(n24128) );
  NOR U22611 ( .A(n24130), .B(n24125), .Z(n24129) );
  XOR U22612 ( .A(n24131), .B(n24132), .Z(n24127) );
  NOR U22613 ( .A(n24133), .B(n24126), .Z(n24132) );
  NOR U22614 ( .A(n24134), .B(n23097), .Z(n24131) );
  XOR U22615 ( .A(n24135), .B(n24136), .Z(n23080) );
  NOR U22616 ( .A(n24137), .B(n23091), .Z(n24136) );
  NOR U22617 ( .A(n24138), .B(n23088), .Z(n24135) );
  XOR U22618 ( .A(n24139), .B(n24140), .Z(n23078) );
  XOR U22619 ( .A(n24141), .B(n24142), .Z(n24140) );
  NOR U22620 ( .A(n24143), .B(n23086), .Z(n24142) );
  NOR U22621 ( .A(n24144), .B(n24145), .Z(n24141) );
  XOR U22622 ( .A(n24146), .B(n24147), .Z(n24139) );
  NOR U22623 ( .A(n24148), .B(n24149), .Z(n24147) );
  NOR U22624 ( .A(n24150), .B(n23076), .Z(n24146) );
  XOR U22625 ( .A(n24151), .B(n24152), .Z(n23072) );
  XOR U22626 ( .A(n24145), .B(n24149), .Z(n24152) );
  XOR U22627 ( .A(n24153), .B(n24154), .Z(n24151) );
  NOR U22628 ( .A(n24155), .B(n23077), .Z(n24154) );
  NOR U22629 ( .A(n24156), .B(n24157), .Z(n24153) );
  XOR U22630 ( .A(n24158), .B(n24159), .Z(n23068) );
  XOR U22631 ( .A(n24160), .B(n24161), .Z(n23066) );
  XNOR U22632 ( .A(n24162), .B(n24157), .Z(n24161) );
  NOR U22633 ( .A(n24163), .B(n24158), .Z(n24162) );
  XOR U22634 ( .A(n24164), .B(n24165), .Z(n24160) );
  NOR U22635 ( .A(n24166), .B(n24159), .Z(n24165) );
  NOR U22636 ( .A(n24167), .B(n23070), .Z(n24164) );
  XOR U22637 ( .A(n24168), .B(n24169), .Z(n23053) );
  NOR U22638 ( .A(n24170), .B(n23064), .Z(n24169) );
  NOR U22639 ( .A(n24171), .B(n23061), .Z(n24168) );
  XOR U22640 ( .A(n24172), .B(n24173), .Z(n23051) );
  XOR U22641 ( .A(n24174), .B(n24175), .Z(n24173) );
  NOR U22642 ( .A(n24176), .B(n23059), .Z(n24175) );
  NOR U22643 ( .A(n24177), .B(n24178), .Z(n24174) );
  XOR U22644 ( .A(n24179), .B(n24180), .Z(n24172) );
  NOR U22645 ( .A(n24181), .B(n24182), .Z(n24180) );
  NOR U22646 ( .A(n24183), .B(n23049), .Z(n24179) );
  XOR U22647 ( .A(n24184), .B(n24185), .Z(n23045) );
  XOR U22648 ( .A(n24178), .B(n24182), .Z(n24185) );
  XOR U22649 ( .A(n24186), .B(n24187), .Z(n24184) );
  NOR U22650 ( .A(n24188), .B(n23050), .Z(n24187) );
  NOR U22651 ( .A(n24189), .B(n24190), .Z(n24186) );
  XOR U22652 ( .A(n24191), .B(n24192), .Z(n23041) );
  XOR U22653 ( .A(n24193), .B(n24194), .Z(n23039) );
  XNOR U22654 ( .A(n24195), .B(n24190), .Z(n24194) );
  NOR U22655 ( .A(n24196), .B(n24191), .Z(n24195) );
  XOR U22656 ( .A(n24197), .B(n24198), .Z(n24193) );
  NOR U22657 ( .A(n24199), .B(n24192), .Z(n24198) );
  NOR U22658 ( .A(n24200), .B(n23043), .Z(n24197) );
  XOR U22659 ( .A(n24201), .B(n24202), .Z(n23026) );
  NOR U22660 ( .A(n24203), .B(n23037), .Z(n24202) );
  NOR U22661 ( .A(n24204), .B(n23034), .Z(n24201) );
  XOR U22662 ( .A(n24205), .B(n24206), .Z(n23024) );
  XOR U22663 ( .A(n24207), .B(n24208), .Z(n24206) );
  NOR U22664 ( .A(n24209), .B(n23032), .Z(n24208) );
  NOR U22665 ( .A(n24210), .B(n24211), .Z(n24207) );
  XOR U22666 ( .A(n24212), .B(n24213), .Z(n24205) );
  NOR U22667 ( .A(n24214), .B(n24215), .Z(n24213) );
  NOR U22668 ( .A(n24216), .B(n23022), .Z(n24212) );
  XOR U22669 ( .A(n24217), .B(n24218), .Z(n23018) );
  XOR U22670 ( .A(n24211), .B(n24215), .Z(n24218) );
  XOR U22671 ( .A(n24219), .B(n24220), .Z(n24217) );
  NOR U22672 ( .A(n24221), .B(n23023), .Z(n24220) );
  NOR U22673 ( .A(n24222), .B(n24223), .Z(n24219) );
  XOR U22674 ( .A(n24224), .B(n24225), .Z(n23014) );
  XOR U22675 ( .A(n24226), .B(n24227), .Z(n23012) );
  XNOR U22676 ( .A(n24228), .B(n24223), .Z(n24227) );
  NOR U22677 ( .A(n24229), .B(n24224), .Z(n24228) );
  XOR U22678 ( .A(n24230), .B(n24231), .Z(n24226) );
  NOR U22679 ( .A(n24232), .B(n24225), .Z(n24231) );
  NOR U22680 ( .A(n24233), .B(n23016), .Z(n24230) );
  XOR U22681 ( .A(n24234), .B(n24235), .Z(n22999) );
  NOR U22682 ( .A(n24236), .B(n23010), .Z(n24235) );
  NOR U22683 ( .A(n24237), .B(n23007), .Z(n24234) );
  XOR U22684 ( .A(n24238), .B(n24239), .Z(n22997) );
  XOR U22685 ( .A(n24240), .B(n24241), .Z(n24239) );
  NOR U22686 ( .A(n24242), .B(n23005), .Z(n24241) );
  NOR U22687 ( .A(n24243), .B(n22988), .Z(n24240) );
  XOR U22688 ( .A(n24244), .B(n24245), .Z(n24238) );
  NOR U22689 ( .A(n24246), .B(n22989), .Z(n24245) );
  NOR U22690 ( .A(n24247), .B(n24248), .Z(n24244) );
  XNOR U22691 ( .A(n22993), .B(n24248), .Z(n22995) );
  XNOR U22692 ( .A(n24249), .B(n24250), .Z(n22954) );
  NOR U22693 ( .A(n50), .B(n24249), .Z(n24250) );
  XOR U22694 ( .A(n31), .B(n22963), .Z(n22965) );
  IV U22695 ( .A(n35), .Z(n31) );
  XOR U22696 ( .A(n22960), .B(n22959), .Z(n35) );
  XNOR U22697 ( .A(n24251), .B(n24252), .Z(n22959) );
  XOR U22698 ( .A(n24253), .B(n24254), .Z(n24252) );
  XOR U22699 ( .A(n24255), .B(n24256), .Z(n24254) );
  AND U22700 ( .A(n24257), .B(n24256), .Z(n24255) );
  XOR U22701 ( .A(n24258), .B(n24259), .Z(n24253) );
  AND U22702 ( .A(n24260), .B(n24261), .Z(n24259) );
  NOR U22703 ( .A(n24262), .B(n24263), .Z(n24258) );
  XOR U22704 ( .A(n24264), .B(n24265), .Z(n24251) );
  XOR U22705 ( .A(n24266), .B(n24267), .Z(n24265) );
  XOR U22706 ( .A(n24268), .B(n24269), .Z(n24267) );
  XOR U22707 ( .A(n24270), .B(n24271), .Z(n24269) );
  XOR U22708 ( .A(n24272), .B(n24273), .Z(n24271) );
  AND U22709 ( .A(n24274), .B(n24273), .Z(n24272) );
  XOR U22710 ( .A(n24275), .B(n24276), .Z(n24270) );
  XOR U22711 ( .A(n24277), .B(n24278), .Z(n24276) );
  XOR U22712 ( .A(n24279), .B(n24280), .Z(n24278) );
  XNOR U22713 ( .A(n24281), .B(n24282), .Z(n24280) );
  NOR U22714 ( .A(n24283), .B(n24282), .Z(n24281) );
  XOR U22715 ( .A(n24284), .B(n24285), .Z(n24279) );
  XOR U22716 ( .A(n24286), .B(n24287), .Z(n24285) );
  XOR U22717 ( .A(n24288), .B(n24289), .Z(n24287) );
  XNOR U22718 ( .A(n24290), .B(n24291), .Z(n24289) );
  NOR U22719 ( .A(n24292), .B(n24291), .Z(n24290) );
  XOR U22720 ( .A(n24293), .B(n24294), .Z(n24288) );
  XOR U22721 ( .A(n24295), .B(n24296), .Z(n24294) );
  XOR U22722 ( .A(n24297), .B(n24298), .Z(n24296) );
  XNOR U22723 ( .A(n24299), .B(n24300), .Z(n24298) );
  NOR U22724 ( .A(n24301), .B(n24300), .Z(n24299) );
  XOR U22725 ( .A(n24302), .B(n24303), .Z(n24297) );
  XOR U22726 ( .A(n24304), .B(n24305), .Z(n24303) );
  XOR U22727 ( .A(n24306), .B(n24307), .Z(n24305) );
  XNOR U22728 ( .A(n24308), .B(n24309), .Z(n24307) );
  NOR U22729 ( .A(n24310), .B(n24309), .Z(n24308) );
  XOR U22730 ( .A(n24311), .B(n24312), .Z(n24306) );
  XOR U22731 ( .A(n24313), .B(n24314), .Z(n24312) );
  XOR U22732 ( .A(n24315), .B(n24316), .Z(n24314) );
  XNOR U22733 ( .A(n24317), .B(n24318), .Z(n24316) );
  NOR U22734 ( .A(n24319), .B(n24318), .Z(n24317) );
  XOR U22735 ( .A(n24320), .B(n24321), .Z(n24315) );
  XOR U22736 ( .A(n24322), .B(n24323), .Z(n24321) );
  XOR U22737 ( .A(n24324), .B(n24325), .Z(n24323) );
  XNOR U22738 ( .A(n24326), .B(n24327), .Z(n24325) );
  NOR U22739 ( .A(n24328), .B(n24327), .Z(n24326) );
  XOR U22740 ( .A(n24329), .B(n24330), .Z(n24324) );
  XOR U22741 ( .A(n24331), .B(n24332), .Z(n24330) );
  XOR U22742 ( .A(n24333), .B(n24334), .Z(n24332) );
  XNOR U22743 ( .A(n24335), .B(n24336), .Z(n24334) );
  NOR U22744 ( .A(n24337), .B(n24336), .Z(n24335) );
  XOR U22745 ( .A(n24338), .B(n24339), .Z(n24333) );
  XOR U22746 ( .A(n24340), .B(n24341), .Z(n24339) );
  XOR U22747 ( .A(n24342), .B(n24343), .Z(n24341) );
  XNOR U22748 ( .A(n24344), .B(n24345), .Z(n24343) );
  NOR U22749 ( .A(n24346), .B(n24345), .Z(n24344) );
  XOR U22750 ( .A(n24347), .B(n24348), .Z(n24342) );
  XOR U22751 ( .A(n24349), .B(n24350), .Z(n24348) );
  XOR U22752 ( .A(n24351), .B(n24352), .Z(n24350) );
  XNOR U22753 ( .A(n24353), .B(n24354), .Z(n24352) );
  NOR U22754 ( .A(n24355), .B(n24354), .Z(n24353) );
  XOR U22755 ( .A(n24356), .B(n24357), .Z(n24351) );
  XOR U22756 ( .A(n24358), .B(n24359), .Z(n24357) );
  XOR U22757 ( .A(n24360), .B(n24361), .Z(n24359) );
  XNOR U22758 ( .A(n24362), .B(n24363), .Z(n24361) );
  NOR U22759 ( .A(n24364), .B(n24363), .Z(n24362) );
  XOR U22760 ( .A(n24365), .B(n24366), .Z(n24360) );
  XOR U22761 ( .A(n24367), .B(n24368), .Z(n24366) );
  XOR U22762 ( .A(n24369), .B(n24370), .Z(n24368) );
  XNOR U22763 ( .A(n24371), .B(n24372), .Z(n24370) );
  NOR U22764 ( .A(n24373), .B(n24372), .Z(n24371) );
  XOR U22765 ( .A(n24374), .B(n24375), .Z(n24369) );
  XOR U22766 ( .A(n24376), .B(n24377), .Z(n24375) );
  XOR U22767 ( .A(n24378), .B(n24379), .Z(n24377) );
  XNOR U22768 ( .A(n24380), .B(n24381), .Z(n24379) );
  NOR U22769 ( .A(n24382), .B(n24381), .Z(n24380) );
  XOR U22770 ( .A(n24383), .B(n24384), .Z(n24378) );
  XOR U22771 ( .A(n24385), .B(n24386), .Z(n24384) );
  XOR U22772 ( .A(n24387), .B(n24388), .Z(n24386) );
  XNOR U22773 ( .A(n24389), .B(n24390), .Z(n24388) );
  NOR U22774 ( .A(n24391), .B(n24390), .Z(n24389) );
  XOR U22775 ( .A(n24392), .B(n24393), .Z(n24387) );
  XOR U22776 ( .A(n24394), .B(n24395), .Z(n24393) );
  XOR U22777 ( .A(n24396), .B(n24397), .Z(n24395) );
  XNOR U22778 ( .A(n24398), .B(n24399), .Z(n24397) );
  NOR U22779 ( .A(n24400), .B(n24399), .Z(n24398) );
  XOR U22780 ( .A(n24401), .B(n24402), .Z(n24396) );
  XOR U22781 ( .A(n24403), .B(n24404), .Z(n24402) );
  XOR U22782 ( .A(n24405), .B(n24406), .Z(n24404) );
  XNOR U22783 ( .A(n24407), .B(n24408), .Z(n24406) );
  NOR U22784 ( .A(n24409), .B(n24408), .Z(n24407) );
  XOR U22785 ( .A(n24410), .B(n24411), .Z(n24405) );
  XOR U22786 ( .A(n24412), .B(n24413), .Z(n24411) );
  XOR U22787 ( .A(n24414), .B(n24415), .Z(n24413) );
  XNOR U22788 ( .A(n24416), .B(n24417), .Z(n24415) );
  NOR U22789 ( .A(n24418), .B(n24417), .Z(n24416) );
  XOR U22790 ( .A(n24419), .B(n24420), .Z(n24414) );
  XOR U22791 ( .A(n24421), .B(n24422), .Z(n24420) );
  XOR U22792 ( .A(n24423), .B(n24424), .Z(n24422) );
  XNOR U22793 ( .A(n24425), .B(n24426), .Z(n24424) );
  NOR U22794 ( .A(n24427), .B(n24426), .Z(n24425) );
  XOR U22795 ( .A(n24428), .B(n24429), .Z(n24423) );
  XOR U22796 ( .A(n24430), .B(n24431), .Z(n24429) );
  XOR U22797 ( .A(n24432), .B(n24433), .Z(n24431) );
  XNOR U22798 ( .A(n24434), .B(n24435), .Z(n24433) );
  NOR U22799 ( .A(n24436), .B(n24435), .Z(n24434) );
  XOR U22800 ( .A(n24437), .B(n24438), .Z(n24432) );
  XOR U22801 ( .A(n24439), .B(n24440), .Z(n24438) );
  XOR U22802 ( .A(n24441), .B(n24442), .Z(n24440) );
  XNOR U22803 ( .A(n24443), .B(n24444), .Z(n24442) );
  NOR U22804 ( .A(n24445), .B(n24444), .Z(n24443) );
  XOR U22805 ( .A(n24446), .B(n24447), .Z(n24441) );
  XOR U22806 ( .A(n24448), .B(n24449), .Z(n24447) );
  XOR U22807 ( .A(n24450), .B(n24451), .Z(n24449) );
  XNOR U22808 ( .A(n24452), .B(n24453), .Z(n24451) );
  NOR U22809 ( .A(n24454), .B(n24453), .Z(n24452) );
  XOR U22810 ( .A(n24455), .B(n24456), .Z(n24450) );
  XOR U22811 ( .A(n24457), .B(n24458), .Z(n24456) );
  XOR U22812 ( .A(n24459), .B(n24460), .Z(n24458) );
  XNOR U22813 ( .A(n24461), .B(n24462), .Z(n24460) );
  NOR U22814 ( .A(n24463), .B(n24462), .Z(n24461) );
  XOR U22815 ( .A(n24464), .B(n24465), .Z(n24459) );
  XOR U22816 ( .A(n24466), .B(n24467), .Z(n24465) );
  XOR U22817 ( .A(n24468), .B(n24469), .Z(n24467) );
  XNOR U22818 ( .A(n24470), .B(n24471), .Z(n24469) );
  NOR U22819 ( .A(n24472), .B(n24471), .Z(n24470) );
  XOR U22820 ( .A(n24473), .B(n24474), .Z(n24468) );
  XOR U22821 ( .A(n24475), .B(n24476), .Z(n24474) );
  XOR U22822 ( .A(n24477), .B(n24478), .Z(n24476) );
  XNOR U22823 ( .A(n24479), .B(n24480), .Z(n24478) );
  NOR U22824 ( .A(n24481), .B(n24480), .Z(n24479) );
  XOR U22825 ( .A(n24482), .B(n24483), .Z(n24477) );
  XOR U22826 ( .A(n24484), .B(n24485), .Z(n24483) );
  XOR U22827 ( .A(n24486), .B(n24487), .Z(n24485) );
  XNOR U22828 ( .A(n24488), .B(n24489), .Z(n24487) );
  NOR U22829 ( .A(n24490), .B(n24489), .Z(n24488) );
  XOR U22830 ( .A(n24491), .B(n24492), .Z(n24486) );
  XOR U22831 ( .A(n24493), .B(n24494), .Z(n24492) );
  XOR U22832 ( .A(n24495), .B(n24496), .Z(n24494) );
  XNOR U22833 ( .A(n24497), .B(n24498), .Z(n24496) );
  NOR U22834 ( .A(n24499), .B(n24498), .Z(n24497) );
  XOR U22835 ( .A(n24500), .B(n24501), .Z(n24495) );
  XOR U22836 ( .A(n24502), .B(n24503), .Z(n24501) );
  XOR U22837 ( .A(n24504), .B(n24505), .Z(n24503) );
  XNOR U22838 ( .A(n24506), .B(n24507), .Z(n24505) );
  NOR U22839 ( .A(n24508), .B(n24507), .Z(n24506) );
  XOR U22840 ( .A(n24509), .B(n24510), .Z(n24504) );
  XOR U22841 ( .A(n24511), .B(n24512), .Z(n24510) );
  XOR U22842 ( .A(n24513), .B(n24514), .Z(n24512) );
  XNOR U22843 ( .A(n24515), .B(n24516), .Z(n24514) );
  NOR U22844 ( .A(n24517), .B(n24516), .Z(n24515) );
  XOR U22845 ( .A(n24518), .B(n24519), .Z(n24513) );
  XOR U22846 ( .A(n24520), .B(n24521), .Z(n24519) );
  XOR U22847 ( .A(n24522), .B(n24523), .Z(n24521) );
  XNOR U22848 ( .A(n24524), .B(n24525), .Z(n24523) );
  NOR U22849 ( .A(n24526), .B(n24525), .Z(n24524) );
  XOR U22850 ( .A(n24527), .B(n24528), .Z(n24522) );
  XOR U22851 ( .A(n24529), .B(n24530), .Z(n24528) );
  XOR U22852 ( .A(n24531), .B(n24532), .Z(n24530) );
  XNOR U22853 ( .A(n24533), .B(n24534), .Z(n24532) );
  NOR U22854 ( .A(n24535), .B(n24534), .Z(n24533) );
  XOR U22855 ( .A(n24536), .B(n24537), .Z(n24531) );
  XOR U22856 ( .A(n24538), .B(n24539), .Z(n24537) );
  XOR U22857 ( .A(n24540), .B(n24541), .Z(n24539) );
  XNOR U22858 ( .A(n24542), .B(n24543), .Z(n24541) );
  NOR U22859 ( .A(n24544), .B(n24543), .Z(n24542) );
  XOR U22860 ( .A(n24545), .B(n24546), .Z(n24540) );
  XOR U22861 ( .A(n24547), .B(n24548), .Z(n24546) );
  XOR U22862 ( .A(n24549), .B(n24550), .Z(n24548) );
  XNOR U22863 ( .A(n24551), .B(n24552), .Z(n24550) );
  NOR U22864 ( .A(n24553), .B(n24552), .Z(n24551) );
  XOR U22865 ( .A(n24554), .B(n24555), .Z(n24549) );
  XOR U22866 ( .A(n24556), .B(n24557), .Z(n24555) );
  XOR U22867 ( .A(n24558), .B(n24559), .Z(n24557) );
  XNOR U22868 ( .A(n24560), .B(n24561), .Z(n24559) );
  NOR U22869 ( .A(n24562), .B(n24561), .Z(n24560) );
  XOR U22870 ( .A(n24563), .B(n24564), .Z(n24558) );
  XOR U22871 ( .A(n24565), .B(n24566), .Z(n24564) );
  XOR U22872 ( .A(n24567), .B(n24568), .Z(n24566) );
  XNOR U22873 ( .A(n24569), .B(n24570), .Z(n24568) );
  NOR U22874 ( .A(n24571), .B(n24570), .Z(n24569) );
  XOR U22875 ( .A(n24572), .B(n24573), .Z(n24567) );
  XOR U22876 ( .A(n24574), .B(n24575), .Z(n24573) );
  XOR U22877 ( .A(n24576), .B(n24577), .Z(n24575) );
  XNOR U22878 ( .A(n24578), .B(n24579), .Z(n24577) );
  NOR U22879 ( .A(n24580), .B(n24579), .Z(n24578) );
  XOR U22880 ( .A(n24581), .B(n24582), .Z(n24576) );
  XOR U22881 ( .A(n24583), .B(n24584), .Z(n24582) );
  XOR U22882 ( .A(n24585), .B(n24586), .Z(n24584) );
  XNOR U22883 ( .A(n24587), .B(n24588), .Z(n24586) );
  NOR U22884 ( .A(n24589), .B(n24588), .Z(n24587) );
  XOR U22885 ( .A(n24590), .B(n24591), .Z(n24585) );
  XOR U22886 ( .A(n24592), .B(n24593), .Z(n24591) );
  XOR U22887 ( .A(n24594), .B(n24595), .Z(n24593) );
  XNOR U22888 ( .A(n24596), .B(n24597), .Z(n24595) );
  NOR U22889 ( .A(n24598), .B(n24597), .Z(n24596) );
  XOR U22890 ( .A(n24599), .B(n24600), .Z(n24594) );
  XOR U22891 ( .A(n24601), .B(n24602), .Z(n24600) );
  XOR U22892 ( .A(n24603), .B(n24604), .Z(n24602) );
  XNOR U22893 ( .A(n24605), .B(n24606), .Z(n24604) );
  NOR U22894 ( .A(n24607), .B(n24606), .Z(n24605) );
  XOR U22895 ( .A(n24608), .B(n24609), .Z(n24603) );
  XOR U22896 ( .A(n24610), .B(n24611), .Z(n24609) );
  XOR U22897 ( .A(n24612), .B(n24613), .Z(n24611) );
  XNOR U22898 ( .A(n24614), .B(n24615), .Z(n24613) );
  NOR U22899 ( .A(n24616), .B(n24615), .Z(n24614) );
  XOR U22900 ( .A(n24617), .B(n24618), .Z(n24612) );
  XOR U22901 ( .A(n24619), .B(n24620), .Z(n24618) );
  XOR U22902 ( .A(n24621), .B(n24622), .Z(n24620) );
  XNOR U22903 ( .A(n24623), .B(n24624), .Z(n24622) );
  NOR U22904 ( .A(n24625), .B(n24624), .Z(n24623) );
  XOR U22905 ( .A(n24626), .B(n24627), .Z(n24621) );
  XOR U22906 ( .A(n24628), .B(n24629), .Z(n24627) );
  XOR U22907 ( .A(n24630), .B(n24631), .Z(n24629) );
  XNOR U22908 ( .A(n24632), .B(n24633), .Z(n24631) );
  NOR U22909 ( .A(n24634), .B(n24633), .Z(n24632) );
  XOR U22910 ( .A(n24635), .B(n24636), .Z(n24630) );
  XOR U22911 ( .A(n24637), .B(n24638), .Z(n24636) );
  XOR U22912 ( .A(n24639), .B(n24640), .Z(n24638) );
  XNOR U22913 ( .A(n24641), .B(n24642), .Z(n24640) );
  NOR U22914 ( .A(n24643), .B(n24642), .Z(n24641) );
  XOR U22915 ( .A(n24644), .B(n24645), .Z(n24639) );
  XOR U22916 ( .A(n24646), .B(n24647), .Z(n24645) );
  XOR U22917 ( .A(n24648), .B(n24649), .Z(n24647) );
  XNOR U22918 ( .A(n24650), .B(n24651), .Z(n24649) );
  NOR U22919 ( .A(n24652), .B(n24651), .Z(n24650) );
  XOR U22920 ( .A(n24653), .B(n24654), .Z(n24648) );
  XOR U22921 ( .A(n24655), .B(n24656), .Z(n24654) );
  XOR U22922 ( .A(n24657), .B(n24658), .Z(n24656) );
  XNOR U22923 ( .A(n24659), .B(n24660), .Z(n24658) );
  NOR U22924 ( .A(n24661), .B(n24660), .Z(n24659) );
  XOR U22925 ( .A(n24662), .B(n24663), .Z(n24657) );
  XOR U22926 ( .A(n24664), .B(n24665), .Z(n24663) );
  XOR U22927 ( .A(n24666), .B(n24667), .Z(n24665) );
  XNOR U22928 ( .A(n24668), .B(n24669), .Z(n24667) );
  NOR U22929 ( .A(n24670), .B(n24669), .Z(n24668) );
  XOR U22930 ( .A(n24671), .B(n24672), .Z(n24666) );
  XOR U22931 ( .A(n24673), .B(n24674), .Z(n24672) );
  XOR U22932 ( .A(n24675), .B(n24676), .Z(n24674) );
  XNOR U22933 ( .A(n24677), .B(n24678), .Z(n24676) );
  NOR U22934 ( .A(n24679), .B(n24678), .Z(n24677) );
  XOR U22935 ( .A(n24680), .B(n24681), .Z(n24675) );
  XOR U22936 ( .A(n24682), .B(n24683), .Z(n24681) );
  XOR U22937 ( .A(n24684), .B(n24685), .Z(n24683) );
  XNOR U22938 ( .A(n24686), .B(n24687), .Z(n24685) );
  NOR U22939 ( .A(n24688), .B(n24687), .Z(n24686) );
  XOR U22940 ( .A(n24689), .B(n24690), .Z(n24684) );
  XOR U22941 ( .A(n24691), .B(n24692), .Z(n24690) );
  XOR U22942 ( .A(n24693), .B(n24694), .Z(n24692) );
  XNOR U22943 ( .A(n24695), .B(n24696), .Z(n24694) );
  NOR U22944 ( .A(n24697), .B(n24696), .Z(n24695) );
  XOR U22945 ( .A(n24698), .B(n24699), .Z(n24693) );
  XOR U22946 ( .A(n24700), .B(n24701), .Z(n24699) );
  XOR U22947 ( .A(n24702), .B(n24703), .Z(n24701) );
  XNOR U22948 ( .A(n24704), .B(n24705), .Z(n24703) );
  NOR U22949 ( .A(n24706), .B(n24705), .Z(n24704) );
  XOR U22950 ( .A(n24707), .B(n24708), .Z(n24702) );
  XOR U22951 ( .A(n24709), .B(n24710), .Z(n24708) );
  XOR U22952 ( .A(n24711), .B(n24712), .Z(n24710) );
  XNOR U22953 ( .A(n24713), .B(n24714), .Z(n24712) );
  NOR U22954 ( .A(n24715), .B(n24714), .Z(n24713) );
  XOR U22955 ( .A(n24716), .B(n24717), .Z(n24711) );
  XOR U22956 ( .A(n24718), .B(n24719), .Z(n24717) );
  XOR U22957 ( .A(n24720), .B(n24721), .Z(n24719) );
  XNOR U22958 ( .A(n24722), .B(n24723), .Z(n24721) );
  NOR U22959 ( .A(n24724), .B(n24723), .Z(n24722) );
  XOR U22960 ( .A(n24725), .B(n24726), .Z(n24720) );
  XOR U22961 ( .A(n24727), .B(n24728), .Z(n24726) );
  XOR U22962 ( .A(n24729), .B(n24730), .Z(n24728) );
  XNOR U22963 ( .A(n24731), .B(n24732), .Z(n24730) );
  NOR U22964 ( .A(n24733), .B(n24732), .Z(n24731) );
  XOR U22965 ( .A(n24734), .B(n24735), .Z(n24729) );
  XOR U22966 ( .A(n24736), .B(n24737), .Z(n24735) );
  XOR U22967 ( .A(n24738), .B(n24739), .Z(n24737) );
  XNOR U22968 ( .A(n24740), .B(n24741), .Z(n24739) );
  NOR U22969 ( .A(n24742), .B(n24741), .Z(n24740) );
  XOR U22970 ( .A(n24743), .B(n24744), .Z(n24738) );
  XOR U22971 ( .A(n24745), .B(n24746), .Z(n24744) );
  XOR U22972 ( .A(n24747), .B(n24748), .Z(n24746) );
  XNOR U22973 ( .A(n24749), .B(n24750), .Z(n24748) );
  NOR U22974 ( .A(n24751), .B(n24750), .Z(n24749) );
  XOR U22975 ( .A(n24752), .B(n24753), .Z(n24747) );
  XOR U22976 ( .A(n24754), .B(n24755), .Z(n24753) );
  XOR U22977 ( .A(n24756), .B(n24757), .Z(n24755) );
  XNOR U22978 ( .A(n24758), .B(n24759), .Z(n24757) );
  NOR U22979 ( .A(n24760), .B(n24759), .Z(n24758) );
  XOR U22980 ( .A(n24761), .B(n24762), .Z(n24756) );
  XOR U22981 ( .A(n24763), .B(n24764), .Z(n24762) );
  XOR U22982 ( .A(n24765), .B(n24766), .Z(n24764) );
  XNOR U22983 ( .A(n24767), .B(n24768), .Z(n24766) );
  NOR U22984 ( .A(n24769), .B(n24768), .Z(n24767) );
  XOR U22985 ( .A(n24770), .B(n24771), .Z(n24765) );
  XOR U22986 ( .A(n24772), .B(n24773), .Z(n24771) );
  XOR U22987 ( .A(n24774), .B(n24775), .Z(n24773) );
  XNOR U22988 ( .A(n24776), .B(n24777), .Z(n24775) );
  NOR U22989 ( .A(n24778), .B(n24777), .Z(n24776) );
  XOR U22990 ( .A(n24779), .B(n24780), .Z(n24774) );
  XOR U22991 ( .A(n24781), .B(n24782), .Z(n24780) );
  XOR U22992 ( .A(n24783), .B(n24784), .Z(n24782) );
  XNOR U22993 ( .A(n24785), .B(n24786), .Z(n24784) );
  NOR U22994 ( .A(n24787), .B(n24786), .Z(n24785) );
  XOR U22995 ( .A(n24788), .B(n24789), .Z(n24783) );
  XOR U22996 ( .A(n24790), .B(n24791), .Z(n24789) );
  XOR U22997 ( .A(n24792), .B(n24793), .Z(n24791) );
  XNOR U22998 ( .A(n24794), .B(n24795), .Z(n24793) );
  NOR U22999 ( .A(n24796), .B(n24795), .Z(n24794) );
  XOR U23000 ( .A(n24797), .B(n24798), .Z(n24792) );
  XOR U23001 ( .A(n24799), .B(n24800), .Z(n24798) );
  XOR U23002 ( .A(n24801), .B(n24802), .Z(n24800) );
  XNOR U23003 ( .A(n24803), .B(n24804), .Z(n24802) );
  NOR U23004 ( .A(n24805), .B(n24804), .Z(n24803) );
  XOR U23005 ( .A(n24806), .B(n24807), .Z(n24801) );
  XOR U23006 ( .A(n24808), .B(n24809), .Z(n24807) );
  XOR U23007 ( .A(n24810), .B(n24811), .Z(n24809) );
  XNOR U23008 ( .A(n24812), .B(n24813), .Z(n24811) );
  NOR U23009 ( .A(n24814), .B(n24813), .Z(n24812) );
  XOR U23010 ( .A(n24815), .B(n24816), .Z(n24810) );
  XOR U23011 ( .A(n24817), .B(n24818), .Z(n24816) );
  XOR U23012 ( .A(n24819), .B(n24820), .Z(n24818) );
  XOR U23013 ( .A(n24821), .B(n24822), .Z(n24817) );
  XNOR U23014 ( .A(n24823), .B(n24824), .Z(n24822) );
  XOR U23015 ( .A(n24825), .B(n24826), .Z(n24824) );
  XOR U23016 ( .A(n24827), .B(n24828), .Z(n24826) );
  XOR U23017 ( .A(n24829), .B(n24830), .Z(n24828) );
  XOR U23018 ( .A(n24831), .B(n24832), .Z(n24827) );
  XOR U23019 ( .A(n24833), .B(n24834), .Z(n24825) );
  XOR U23020 ( .A(n24835), .B(n24836), .Z(n24834) );
  AND U23021 ( .A(n24837), .B(n24838), .Z(n24836) );
  XNOR U23022 ( .A(n24839), .B(n24830), .Z(n24837) );
  XNOR U23023 ( .A(n24840), .B(n24841), .Z(n24830) );
  AND U23024 ( .A(n24839), .B(n24840), .Z(n24841) );
  NOR U23025 ( .A(n24842), .B(n24831), .Z(n24835) );
  XOR U23026 ( .A(n24843), .B(n24844), .Z(n24833) );
  NOR U23027 ( .A(n24845), .B(n24832), .Z(n24844) );
  NOR U23028 ( .A(n24846), .B(n24829), .Z(n24843) );
  XNOR U23029 ( .A(n24847), .B(n24848), .Z(n24821) );
  XNOR U23030 ( .A(n24849), .B(n24850), .Z(n24848) );
  NOR U23031 ( .A(n24851), .B(n24823), .Z(n24849) );
  XOR U23032 ( .A(n24852), .B(n24853), .Z(n24815) );
  XOR U23033 ( .A(n24854), .B(n24855), .Z(n24853) );
  NOR U23034 ( .A(n24856), .B(n24819), .Z(n24855) );
  NOR U23035 ( .A(n24857), .B(n24850), .Z(n24854) );
  XOR U23036 ( .A(n24858), .B(n24859), .Z(n24852) );
  NOR U23037 ( .A(n24860), .B(n24847), .Z(n24859) );
  NOR U23038 ( .A(n24861), .B(n24820), .Z(n24858) );
  XOR U23039 ( .A(n24862), .B(n24863), .Z(n24808) );
  XOR U23040 ( .A(n24864), .B(n24865), .Z(n24806) );
  XNOR U23041 ( .A(n24866), .B(n24867), .Z(n24865) );
  NOR U23042 ( .A(n24868), .B(n24867), .Z(n24866) );
  XOR U23043 ( .A(n24869), .B(n24870), .Z(n24864) );
  NOR U23044 ( .A(n24871), .B(n24862), .Z(n24870) );
  NOR U23045 ( .A(n24872), .B(n24863), .Z(n24869) );
  XOR U23046 ( .A(n24873), .B(n24874), .Z(n24799) );
  XOR U23047 ( .A(n24875), .B(n24876), .Z(n24797) );
  XNOR U23048 ( .A(n24877), .B(n24878), .Z(n24876) );
  NOR U23049 ( .A(n24879), .B(n24878), .Z(n24877) );
  XOR U23050 ( .A(n24880), .B(n24881), .Z(n24875) );
  NOR U23051 ( .A(n24882), .B(n24873), .Z(n24881) );
  NOR U23052 ( .A(n24883), .B(n24874), .Z(n24880) );
  XOR U23053 ( .A(n24884), .B(n24885), .Z(n24790) );
  XOR U23054 ( .A(n24886), .B(n24887), .Z(n24788) );
  XNOR U23055 ( .A(n24888), .B(n24889), .Z(n24887) );
  NOR U23056 ( .A(n24890), .B(n24889), .Z(n24888) );
  XOR U23057 ( .A(n24891), .B(n24892), .Z(n24886) );
  NOR U23058 ( .A(n24893), .B(n24884), .Z(n24892) );
  NOR U23059 ( .A(n24894), .B(n24885), .Z(n24891) );
  XOR U23060 ( .A(n24895), .B(n24896), .Z(n24781) );
  XOR U23061 ( .A(n24897), .B(n24898), .Z(n24779) );
  XNOR U23062 ( .A(n24899), .B(n24900), .Z(n24898) );
  NOR U23063 ( .A(n24901), .B(n24900), .Z(n24899) );
  XOR U23064 ( .A(n24902), .B(n24903), .Z(n24897) );
  NOR U23065 ( .A(n24904), .B(n24895), .Z(n24903) );
  NOR U23066 ( .A(n24905), .B(n24896), .Z(n24902) );
  XOR U23067 ( .A(n24906), .B(n24907), .Z(n24772) );
  XOR U23068 ( .A(n24908), .B(n24909), .Z(n24770) );
  XNOR U23069 ( .A(n24910), .B(n24911), .Z(n24909) );
  NOR U23070 ( .A(n24912), .B(n24911), .Z(n24910) );
  XOR U23071 ( .A(n24913), .B(n24914), .Z(n24908) );
  NOR U23072 ( .A(n24915), .B(n24906), .Z(n24914) );
  NOR U23073 ( .A(n24916), .B(n24907), .Z(n24913) );
  XOR U23074 ( .A(n24917), .B(n24918), .Z(n24763) );
  XOR U23075 ( .A(n24919), .B(n24920), .Z(n24761) );
  XNOR U23076 ( .A(n24921), .B(n24922), .Z(n24920) );
  NOR U23077 ( .A(n24923), .B(n24922), .Z(n24921) );
  XOR U23078 ( .A(n24924), .B(n24925), .Z(n24919) );
  NOR U23079 ( .A(n24926), .B(n24917), .Z(n24925) );
  NOR U23080 ( .A(n24927), .B(n24918), .Z(n24924) );
  XOR U23081 ( .A(n24928), .B(n24929), .Z(n24754) );
  XOR U23082 ( .A(n24930), .B(n24931), .Z(n24752) );
  XNOR U23083 ( .A(n24932), .B(n24933), .Z(n24931) );
  NOR U23084 ( .A(n24934), .B(n24933), .Z(n24932) );
  XOR U23085 ( .A(n24935), .B(n24936), .Z(n24930) );
  NOR U23086 ( .A(n24937), .B(n24928), .Z(n24936) );
  NOR U23087 ( .A(n24938), .B(n24929), .Z(n24935) );
  XOR U23088 ( .A(n24939), .B(n24940), .Z(n24745) );
  XOR U23089 ( .A(n24941), .B(n24942), .Z(n24743) );
  XNOR U23090 ( .A(n24943), .B(n24944), .Z(n24942) );
  NOR U23091 ( .A(n24945), .B(n24944), .Z(n24943) );
  XOR U23092 ( .A(n24946), .B(n24947), .Z(n24941) );
  NOR U23093 ( .A(n24948), .B(n24939), .Z(n24947) );
  NOR U23094 ( .A(n24949), .B(n24940), .Z(n24946) );
  XOR U23095 ( .A(n24950), .B(n24951), .Z(n24736) );
  XOR U23096 ( .A(n24952), .B(n24953), .Z(n24734) );
  XNOR U23097 ( .A(n24954), .B(n24955), .Z(n24953) );
  NOR U23098 ( .A(n24956), .B(n24955), .Z(n24954) );
  XOR U23099 ( .A(n24957), .B(n24958), .Z(n24952) );
  NOR U23100 ( .A(n24959), .B(n24950), .Z(n24958) );
  NOR U23101 ( .A(n24960), .B(n24951), .Z(n24957) );
  XOR U23102 ( .A(n24961), .B(n24962), .Z(n24727) );
  XOR U23103 ( .A(n24963), .B(n24964), .Z(n24725) );
  XNOR U23104 ( .A(n24965), .B(n24966), .Z(n24964) );
  NOR U23105 ( .A(n24967), .B(n24966), .Z(n24965) );
  XOR U23106 ( .A(n24968), .B(n24969), .Z(n24963) );
  NOR U23107 ( .A(n24970), .B(n24961), .Z(n24969) );
  NOR U23108 ( .A(n24971), .B(n24962), .Z(n24968) );
  XOR U23109 ( .A(n24972), .B(n24973), .Z(n24718) );
  XOR U23110 ( .A(n24974), .B(n24975), .Z(n24716) );
  XNOR U23111 ( .A(n24976), .B(n24977), .Z(n24975) );
  NOR U23112 ( .A(n24978), .B(n24977), .Z(n24976) );
  XOR U23113 ( .A(n24979), .B(n24980), .Z(n24974) );
  NOR U23114 ( .A(n24981), .B(n24972), .Z(n24980) );
  NOR U23115 ( .A(n24982), .B(n24973), .Z(n24979) );
  XOR U23116 ( .A(n24983), .B(n24984), .Z(n24709) );
  XOR U23117 ( .A(n24985), .B(n24986), .Z(n24707) );
  XNOR U23118 ( .A(n24987), .B(n24988), .Z(n24986) );
  NOR U23119 ( .A(n24989), .B(n24988), .Z(n24987) );
  XOR U23120 ( .A(n24990), .B(n24991), .Z(n24985) );
  NOR U23121 ( .A(n24992), .B(n24983), .Z(n24991) );
  NOR U23122 ( .A(n24993), .B(n24984), .Z(n24990) );
  XOR U23123 ( .A(n24994), .B(n24995), .Z(n24700) );
  XOR U23124 ( .A(n24996), .B(n24997), .Z(n24698) );
  XNOR U23125 ( .A(n24998), .B(n24999), .Z(n24997) );
  NOR U23126 ( .A(n25000), .B(n24999), .Z(n24998) );
  XOR U23127 ( .A(n25001), .B(n25002), .Z(n24996) );
  NOR U23128 ( .A(n25003), .B(n24994), .Z(n25002) );
  NOR U23129 ( .A(n25004), .B(n24995), .Z(n25001) );
  XOR U23130 ( .A(n25005), .B(n25006), .Z(n24691) );
  XOR U23131 ( .A(n25007), .B(n25008), .Z(n24689) );
  XNOR U23132 ( .A(n25009), .B(n25010), .Z(n25008) );
  NOR U23133 ( .A(n25011), .B(n25010), .Z(n25009) );
  XOR U23134 ( .A(n25012), .B(n25013), .Z(n25007) );
  NOR U23135 ( .A(n25014), .B(n25005), .Z(n25013) );
  NOR U23136 ( .A(n25015), .B(n25006), .Z(n25012) );
  XOR U23137 ( .A(n25016), .B(n25017), .Z(n24682) );
  XOR U23138 ( .A(n25018), .B(n25019), .Z(n24680) );
  XNOR U23139 ( .A(n25020), .B(n25021), .Z(n25019) );
  NOR U23140 ( .A(n25022), .B(n25021), .Z(n25020) );
  XOR U23141 ( .A(n25023), .B(n25024), .Z(n25018) );
  NOR U23142 ( .A(n25025), .B(n25016), .Z(n25024) );
  NOR U23143 ( .A(n25026), .B(n25017), .Z(n25023) );
  XOR U23144 ( .A(n25027), .B(n25028), .Z(n24673) );
  XOR U23145 ( .A(n25029), .B(n25030), .Z(n24671) );
  XNOR U23146 ( .A(n25031), .B(n25032), .Z(n25030) );
  NOR U23147 ( .A(n25033), .B(n25032), .Z(n25031) );
  XOR U23148 ( .A(n25034), .B(n25035), .Z(n25029) );
  NOR U23149 ( .A(n25036), .B(n25027), .Z(n25035) );
  NOR U23150 ( .A(n25037), .B(n25028), .Z(n25034) );
  XOR U23151 ( .A(n25038), .B(n25039), .Z(n24664) );
  XOR U23152 ( .A(n25040), .B(n25041), .Z(n24662) );
  XNOR U23153 ( .A(n25042), .B(n25043), .Z(n25041) );
  NOR U23154 ( .A(n25044), .B(n25043), .Z(n25042) );
  XOR U23155 ( .A(n25045), .B(n25046), .Z(n25040) );
  NOR U23156 ( .A(n25047), .B(n25038), .Z(n25046) );
  NOR U23157 ( .A(n25048), .B(n25039), .Z(n25045) );
  XOR U23158 ( .A(n25049), .B(n25050), .Z(n24655) );
  XOR U23159 ( .A(n25051), .B(n25052), .Z(n24653) );
  XNOR U23160 ( .A(n25053), .B(n25054), .Z(n25052) );
  NOR U23161 ( .A(n25055), .B(n25054), .Z(n25053) );
  XOR U23162 ( .A(n25056), .B(n25057), .Z(n25051) );
  NOR U23163 ( .A(n25058), .B(n25049), .Z(n25057) );
  NOR U23164 ( .A(n25059), .B(n25050), .Z(n25056) );
  XOR U23165 ( .A(n25060), .B(n25061), .Z(n24646) );
  XOR U23166 ( .A(n25062), .B(n25063), .Z(n24644) );
  XNOR U23167 ( .A(n25064), .B(n25065), .Z(n25063) );
  NOR U23168 ( .A(n25066), .B(n25065), .Z(n25064) );
  XOR U23169 ( .A(n25067), .B(n25068), .Z(n25062) );
  NOR U23170 ( .A(n25069), .B(n25060), .Z(n25068) );
  NOR U23171 ( .A(n25070), .B(n25061), .Z(n25067) );
  XOR U23172 ( .A(n25071), .B(n25072), .Z(n24637) );
  XOR U23173 ( .A(n25073), .B(n25074), .Z(n24635) );
  XNOR U23174 ( .A(n25075), .B(n25076), .Z(n25074) );
  NOR U23175 ( .A(n25077), .B(n25076), .Z(n25075) );
  XOR U23176 ( .A(n25078), .B(n25079), .Z(n25073) );
  NOR U23177 ( .A(n25080), .B(n25071), .Z(n25079) );
  NOR U23178 ( .A(n25081), .B(n25072), .Z(n25078) );
  XOR U23179 ( .A(n25082), .B(n25083), .Z(n24628) );
  XOR U23180 ( .A(n25084), .B(n25085), .Z(n24626) );
  XNOR U23181 ( .A(n25086), .B(n25087), .Z(n25085) );
  NOR U23182 ( .A(n25088), .B(n25087), .Z(n25086) );
  XOR U23183 ( .A(n25089), .B(n25090), .Z(n25084) );
  NOR U23184 ( .A(n25091), .B(n25082), .Z(n25090) );
  NOR U23185 ( .A(n25092), .B(n25083), .Z(n25089) );
  XOR U23186 ( .A(n25093), .B(n25094), .Z(n24619) );
  XOR U23187 ( .A(n25095), .B(n25096), .Z(n24617) );
  XNOR U23188 ( .A(n25097), .B(n25098), .Z(n25096) );
  NOR U23189 ( .A(n25099), .B(n25098), .Z(n25097) );
  XOR U23190 ( .A(n25100), .B(n25101), .Z(n25095) );
  NOR U23191 ( .A(n25102), .B(n25093), .Z(n25101) );
  NOR U23192 ( .A(n25103), .B(n25094), .Z(n25100) );
  XOR U23193 ( .A(n25104), .B(n25105), .Z(n24610) );
  XOR U23194 ( .A(n25106), .B(n25107), .Z(n24608) );
  XNOR U23195 ( .A(n25108), .B(n25109), .Z(n25107) );
  NOR U23196 ( .A(n25110), .B(n25109), .Z(n25108) );
  XOR U23197 ( .A(n25111), .B(n25112), .Z(n25106) );
  NOR U23198 ( .A(n25113), .B(n25104), .Z(n25112) );
  NOR U23199 ( .A(n25114), .B(n25105), .Z(n25111) );
  XOR U23200 ( .A(n25115), .B(n25116), .Z(n24601) );
  XOR U23201 ( .A(n25117), .B(n25118), .Z(n24599) );
  XNOR U23202 ( .A(n25119), .B(n25120), .Z(n25118) );
  NOR U23203 ( .A(n25121), .B(n25120), .Z(n25119) );
  XOR U23204 ( .A(n25122), .B(n25123), .Z(n25117) );
  NOR U23205 ( .A(n25124), .B(n25115), .Z(n25123) );
  NOR U23206 ( .A(n25125), .B(n25116), .Z(n25122) );
  XOR U23207 ( .A(n25126), .B(n25127), .Z(n24592) );
  XOR U23208 ( .A(n25128), .B(n25129), .Z(n24590) );
  XNOR U23209 ( .A(n25130), .B(n25131), .Z(n25129) );
  NOR U23210 ( .A(n25132), .B(n25131), .Z(n25130) );
  XOR U23211 ( .A(n25133), .B(n25134), .Z(n25128) );
  NOR U23212 ( .A(n25135), .B(n25126), .Z(n25134) );
  NOR U23213 ( .A(n25136), .B(n25127), .Z(n25133) );
  XOR U23214 ( .A(n25137), .B(n25138), .Z(n24583) );
  XOR U23215 ( .A(n25139), .B(n25140), .Z(n24581) );
  XNOR U23216 ( .A(n25141), .B(n25142), .Z(n25140) );
  NOR U23217 ( .A(n25143), .B(n25142), .Z(n25141) );
  XOR U23218 ( .A(n25144), .B(n25145), .Z(n25139) );
  NOR U23219 ( .A(n25146), .B(n25137), .Z(n25145) );
  NOR U23220 ( .A(n25147), .B(n25138), .Z(n25144) );
  XOR U23221 ( .A(n25148), .B(n25149), .Z(n24574) );
  XOR U23222 ( .A(n25150), .B(n25151), .Z(n24572) );
  XNOR U23223 ( .A(n25152), .B(n25153), .Z(n25151) );
  NOR U23224 ( .A(n25154), .B(n25153), .Z(n25152) );
  XOR U23225 ( .A(n25155), .B(n25156), .Z(n25150) );
  NOR U23226 ( .A(n25157), .B(n25148), .Z(n25156) );
  NOR U23227 ( .A(n25158), .B(n25149), .Z(n25155) );
  XOR U23228 ( .A(n25159), .B(n25160), .Z(n24565) );
  XOR U23229 ( .A(n25161), .B(n25162), .Z(n24563) );
  XNOR U23230 ( .A(n25163), .B(n25164), .Z(n25162) );
  NOR U23231 ( .A(n25165), .B(n25164), .Z(n25163) );
  XOR U23232 ( .A(n25166), .B(n25167), .Z(n25161) );
  NOR U23233 ( .A(n25168), .B(n25159), .Z(n25167) );
  NOR U23234 ( .A(n25169), .B(n25160), .Z(n25166) );
  XOR U23235 ( .A(n25170), .B(n25171), .Z(n24556) );
  XOR U23236 ( .A(n25172), .B(n25173), .Z(n24554) );
  XNOR U23237 ( .A(n25174), .B(n25175), .Z(n25173) );
  NOR U23238 ( .A(n25176), .B(n25175), .Z(n25174) );
  XOR U23239 ( .A(n25177), .B(n25178), .Z(n25172) );
  NOR U23240 ( .A(n25179), .B(n25170), .Z(n25178) );
  NOR U23241 ( .A(n25180), .B(n25171), .Z(n25177) );
  XOR U23242 ( .A(n25181), .B(n25182), .Z(n24547) );
  XOR U23243 ( .A(n25183), .B(n25184), .Z(n24545) );
  XNOR U23244 ( .A(n25185), .B(n25186), .Z(n25184) );
  NOR U23245 ( .A(n25187), .B(n25186), .Z(n25185) );
  XOR U23246 ( .A(n25188), .B(n25189), .Z(n25183) );
  NOR U23247 ( .A(n25190), .B(n25181), .Z(n25189) );
  NOR U23248 ( .A(n25191), .B(n25182), .Z(n25188) );
  XOR U23249 ( .A(n25192), .B(n25193), .Z(n24538) );
  XOR U23250 ( .A(n25194), .B(n25195), .Z(n24536) );
  XNOR U23251 ( .A(n25196), .B(n25197), .Z(n25195) );
  NOR U23252 ( .A(n25198), .B(n25197), .Z(n25196) );
  XOR U23253 ( .A(n25199), .B(n25200), .Z(n25194) );
  NOR U23254 ( .A(n25201), .B(n25192), .Z(n25200) );
  NOR U23255 ( .A(n25202), .B(n25193), .Z(n25199) );
  XOR U23256 ( .A(n25203), .B(n25204), .Z(n24529) );
  XOR U23257 ( .A(n25205), .B(n25206), .Z(n24527) );
  XNOR U23258 ( .A(n25207), .B(n25208), .Z(n25206) );
  NOR U23259 ( .A(n25209), .B(n25208), .Z(n25207) );
  XOR U23260 ( .A(n25210), .B(n25211), .Z(n25205) );
  NOR U23261 ( .A(n25212), .B(n25203), .Z(n25211) );
  NOR U23262 ( .A(n25213), .B(n25204), .Z(n25210) );
  XOR U23263 ( .A(n25214), .B(n25215), .Z(n24520) );
  XOR U23264 ( .A(n25216), .B(n25217), .Z(n24518) );
  XNOR U23265 ( .A(n25218), .B(n25219), .Z(n25217) );
  NOR U23266 ( .A(n25220), .B(n25219), .Z(n25218) );
  XOR U23267 ( .A(n25221), .B(n25222), .Z(n25216) );
  NOR U23268 ( .A(n25223), .B(n25214), .Z(n25222) );
  NOR U23269 ( .A(n25224), .B(n25215), .Z(n25221) );
  XOR U23270 ( .A(n25225), .B(n25226), .Z(n24511) );
  XOR U23271 ( .A(n25227), .B(n25228), .Z(n24509) );
  XNOR U23272 ( .A(n25229), .B(n25230), .Z(n25228) );
  NOR U23273 ( .A(n25231), .B(n25230), .Z(n25229) );
  XOR U23274 ( .A(n25232), .B(n25233), .Z(n25227) );
  NOR U23275 ( .A(n25234), .B(n25225), .Z(n25233) );
  NOR U23276 ( .A(n25235), .B(n25226), .Z(n25232) );
  XOR U23277 ( .A(n25236), .B(n25237), .Z(n24502) );
  XOR U23278 ( .A(n25238), .B(n25239), .Z(n24500) );
  XNOR U23279 ( .A(n25240), .B(n25241), .Z(n25239) );
  NOR U23280 ( .A(n25242), .B(n25241), .Z(n25240) );
  XOR U23281 ( .A(n25243), .B(n25244), .Z(n25238) );
  NOR U23282 ( .A(n25245), .B(n25236), .Z(n25244) );
  NOR U23283 ( .A(n25246), .B(n25237), .Z(n25243) );
  XOR U23284 ( .A(n25247), .B(n25248), .Z(n24493) );
  XOR U23285 ( .A(n25249), .B(n25250), .Z(n24491) );
  XNOR U23286 ( .A(n25251), .B(n25252), .Z(n25250) );
  NOR U23287 ( .A(n25253), .B(n25252), .Z(n25251) );
  XOR U23288 ( .A(n25254), .B(n25255), .Z(n25249) );
  NOR U23289 ( .A(n25256), .B(n25247), .Z(n25255) );
  NOR U23290 ( .A(n25257), .B(n25248), .Z(n25254) );
  XOR U23291 ( .A(n25258), .B(n25259), .Z(n24484) );
  XOR U23292 ( .A(n25260), .B(n25261), .Z(n24482) );
  XNOR U23293 ( .A(n25262), .B(n25263), .Z(n25261) );
  NOR U23294 ( .A(n25264), .B(n25263), .Z(n25262) );
  XOR U23295 ( .A(n25265), .B(n25266), .Z(n25260) );
  NOR U23296 ( .A(n25267), .B(n25258), .Z(n25266) );
  NOR U23297 ( .A(n25268), .B(n25259), .Z(n25265) );
  XOR U23298 ( .A(n25269), .B(n25270), .Z(n24475) );
  XOR U23299 ( .A(n25271), .B(n25272), .Z(n24473) );
  XNOR U23300 ( .A(n25273), .B(n25274), .Z(n25272) );
  NOR U23301 ( .A(n25275), .B(n25274), .Z(n25273) );
  XOR U23302 ( .A(n25276), .B(n25277), .Z(n25271) );
  NOR U23303 ( .A(n25278), .B(n25269), .Z(n25277) );
  NOR U23304 ( .A(n25279), .B(n25270), .Z(n25276) );
  XOR U23305 ( .A(n25280), .B(n25281), .Z(n24466) );
  XOR U23306 ( .A(n25282), .B(n25283), .Z(n24464) );
  XNOR U23307 ( .A(n25284), .B(n25285), .Z(n25283) );
  NOR U23308 ( .A(n25286), .B(n25285), .Z(n25284) );
  XOR U23309 ( .A(n25287), .B(n25288), .Z(n25282) );
  NOR U23310 ( .A(n25289), .B(n25280), .Z(n25288) );
  NOR U23311 ( .A(n25290), .B(n25281), .Z(n25287) );
  XOR U23312 ( .A(n25291), .B(n25292), .Z(n24457) );
  XOR U23313 ( .A(n25293), .B(n25294), .Z(n24455) );
  XNOR U23314 ( .A(n25295), .B(n25296), .Z(n25294) );
  NOR U23315 ( .A(n25297), .B(n25296), .Z(n25295) );
  XOR U23316 ( .A(n25298), .B(n25299), .Z(n25293) );
  NOR U23317 ( .A(n25300), .B(n25291), .Z(n25299) );
  NOR U23318 ( .A(n25301), .B(n25292), .Z(n25298) );
  XOR U23319 ( .A(n25302), .B(n25303), .Z(n24448) );
  XOR U23320 ( .A(n25304), .B(n25305), .Z(n24446) );
  XNOR U23321 ( .A(n25306), .B(n25307), .Z(n25305) );
  NOR U23322 ( .A(n25308), .B(n25307), .Z(n25306) );
  XOR U23323 ( .A(n25309), .B(n25310), .Z(n25304) );
  NOR U23324 ( .A(n25311), .B(n25302), .Z(n25310) );
  NOR U23325 ( .A(n25312), .B(n25303), .Z(n25309) );
  XOR U23326 ( .A(n25313), .B(n25314), .Z(n24439) );
  XOR U23327 ( .A(n25315), .B(n25316), .Z(n24437) );
  XNOR U23328 ( .A(n25317), .B(n25318), .Z(n25316) );
  NOR U23329 ( .A(n25319), .B(n25318), .Z(n25317) );
  XOR U23330 ( .A(n25320), .B(n25321), .Z(n25315) );
  NOR U23331 ( .A(n25322), .B(n25313), .Z(n25321) );
  NOR U23332 ( .A(n25323), .B(n25314), .Z(n25320) );
  XOR U23333 ( .A(n25324), .B(n25325), .Z(n24430) );
  XOR U23334 ( .A(n25326), .B(n25327), .Z(n24428) );
  XNOR U23335 ( .A(n25328), .B(n25329), .Z(n25327) );
  NOR U23336 ( .A(n25330), .B(n25329), .Z(n25328) );
  XOR U23337 ( .A(n25331), .B(n25332), .Z(n25326) );
  NOR U23338 ( .A(n25333), .B(n25324), .Z(n25332) );
  NOR U23339 ( .A(n25334), .B(n25325), .Z(n25331) );
  XOR U23340 ( .A(n25335), .B(n25336), .Z(n24421) );
  XOR U23341 ( .A(n25337), .B(n25338), .Z(n24419) );
  XNOR U23342 ( .A(n25339), .B(n25340), .Z(n25338) );
  NOR U23343 ( .A(n25341), .B(n25340), .Z(n25339) );
  XOR U23344 ( .A(n25342), .B(n25343), .Z(n25337) );
  NOR U23345 ( .A(n25344), .B(n25335), .Z(n25343) );
  NOR U23346 ( .A(n25345), .B(n25336), .Z(n25342) );
  XOR U23347 ( .A(n25346), .B(n25347), .Z(n24412) );
  XOR U23348 ( .A(n25348), .B(n25349), .Z(n24410) );
  XNOR U23349 ( .A(n25350), .B(n25351), .Z(n25349) );
  NOR U23350 ( .A(n25352), .B(n25351), .Z(n25350) );
  XOR U23351 ( .A(n25353), .B(n25354), .Z(n25348) );
  NOR U23352 ( .A(n25355), .B(n25346), .Z(n25354) );
  NOR U23353 ( .A(n25356), .B(n25347), .Z(n25353) );
  XOR U23354 ( .A(n25357), .B(n25358), .Z(n24403) );
  XOR U23355 ( .A(n25359), .B(n25360), .Z(n24401) );
  XNOR U23356 ( .A(n25361), .B(n25362), .Z(n25360) );
  NOR U23357 ( .A(n25363), .B(n25362), .Z(n25361) );
  XOR U23358 ( .A(n25364), .B(n25365), .Z(n25359) );
  NOR U23359 ( .A(n25366), .B(n25357), .Z(n25365) );
  NOR U23360 ( .A(n25367), .B(n25358), .Z(n25364) );
  XOR U23361 ( .A(n25368), .B(n25369), .Z(n24394) );
  XOR U23362 ( .A(n25370), .B(n25371), .Z(n24392) );
  XNOR U23363 ( .A(n25372), .B(n25373), .Z(n25371) );
  NOR U23364 ( .A(n25374), .B(n25373), .Z(n25372) );
  XOR U23365 ( .A(n25375), .B(n25376), .Z(n25370) );
  NOR U23366 ( .A(n25377), .B(n25368), .Z(n25376) );
  NOR U23367 ( .A(n25378), .B(n25369), .Z(n25375) );
  XOR U23368 ( .A(n25379), .B(n25380), .Z(n24385) );
  XOR U23369 ( .A(n25381), .B(n25382), .Z(n24383) );
  XNOR U23370 ( .A(n25383), .B(n25384), .Z(n25382) );
  NOR U23371 ( .A(n25385), .B(n25384), .Z(n25383) );
  XOR U23372 ( .A(n25386), .B(n25387), .Z(n25381) );
  NOR U23373 ( .A(n25388), .B(n25379), .Z(n25387) );
  NOR U23374 ( .A(n25389), .B(n25380), .Z(n25386) );
  XOR U23375 ( .A(n25390), .B(n25391), .Z(n24376) );
  XOR U23376 ( .A(n25392), .B(n25393), .Z(n24374) );
  XNOR U23377 ( .A(n25394), .B(n25395), .Z(n25393) );
  NOR U23378 ( .A(n25396), .B(n25395), .Z(n25394) );
  XOR U23379 ( .A(n25397), .B(n25398), .Z(n25392) );
  NOR U23380 ( .A(n25399), .B(n25390), .Z(n25398) );
  NOR U23381 ( .A(n25400), .B(n25391), .Z(n25397) );
  XOR U23382 ( .A(n25401), .B(n25402), .Z(n24367) );
  XOR U23383 ( .A(n25403), .B(n25404), .Z(n24365) );
  XNOR U23384 ( .A(n25405), .B(n25406), .Z(n25404) );
  NOR U23385 ( .A(n25407), .B(n25406), .Z(n25405) );
  XOR U23386 ( .A(n25408), .B(n25409), .Z(n25403) );
  NOR U23387 ( .A(n25410), .B(n25401), .Z(n25409) );
  NOR U23388 ( .A(n25411), .B(n25402), .Z(n25408) );
  XOR U23389 ( .A(n25412), .B(n25413), .Z(n24358) );
  XOR U23390 ( .A(n25414), .B(n25415), .Z(n24356) );
  XNOR U23391 ( .A(n25416), .B(n25417), .Z(n25415) );
  NOR U23392 ( .A(n25418), .B(n25417), .Z(n25416) );
  XOR U23393 ( .A(n25419), .B(n25420), .Z(n25414) );
  NOR U23394 ( .A(n25421), .B(n25412), .Z(n25420) );
  NOR U23395 ( .A(n25422), .B(n25413), .Z(n25419) );
  XOR U23396 ( .A(n25423), .B(n25424), .Z(n24349) );
  XOR U23397 ( .A(n25425), .B(n25426), .Z(n24347) );
  XNOR U23398 ( .A(n25427), .B(n25428), .Z(n25426) );
  NOR U23399 ( .A(n25429), .B(n25428), .Z(n25427) );
  XOR U23400 ( .A(n25430), .B(n25431), .Z(n25425) );
  NOR U23401 ( .A(n25432), .B(n25423), .Z(n25431) );
  NOR U23402 ( .A(n25433), .B(n25424), .Z(n25430) );
  XOR U23403 ( .A(n25434), .B(n25435), .Z(n24340) );
  XOR U23404 ( .A(n25436), .B(n25437), .Z(n24338) );
  XNOR U23405 ( .A(n25438), .B(n25439), .Z(n25437) );
  NOR U23406 ( .A(n25440), .B(n25439), .Z(n25438) );
  XOR U23407 ( .A(n25441), .B(n25442), .Z(n25436) );
  NOR U23408 ( .A(n25443), .B(n25434), .Z(n25442) );
  NOR U23409 ( .A(n25444), .B(n25435), .Z(n25441) );
  XOR U23410 ( .A(n25445), .B(n25446), .Z(n24331) );
  XOR U23411 ( .A(n25447), .B(n25448), .Z(n24329) );
  XNOR U23412 ( .A(n25449), .B(n25450), .Z(n25448) );
  NOR U23413 ( .A(n25451), .B(n25450), .Z(n25449) );
  XOR U23414 ( .A(n25452), .B(n25453), .Z(n25447) );
  NOR U23415 ( .A(n25454), .B(n25445), .Z(n25453) );
  NOR U23416 ( .A(n25455), .B(n25446), .Z(n25452) );
  XOR U23417 ( .A(n25456), .B(n25457), .Z(n24322) );
  XOR U23418 ( .A(n25458), .B(n25459), .Z(n24320) );
  XNOR U23419 ( .A(n25460), .B(n25461), .Z(n25459) );
  NOR U23420 ( .A(n25462), .B(n25461), .Z(n25460) );
  XOR U23421 ( .A(n25463), .B(n25464), .Z(n25458) );
  NOR U23422 ( .A(n25465), .B(n25456), .Z(n25464) );
  NOR U23423 ( .A(n25466), .B(n25457), .Z(n25463) );
  XOR U23424 ( .A(n25467), .B(n25468), .Z(n24313) );
  XOR U23425 ( .A(n25469), .B(n25470), .Z(n24311) );
  XNOR U23426 ( .A(n25471), .B(n25472), .Z(n25470) );
  NOR U23427 ( .A(n25473), .B(n25472), .Z(n25471) );
  XOR U23428 ( .A(n25474), .B(n25475), .Z(n25469) );
  NOR U23429 ( .A(n25476), .B(n25467), .Z(n25475) );
  NOR U23430 ( .A(n25477), .B(n25468), .Z(n25474) );
  XOR U23431 ( .A(n25478), .B(n25479), .Z(n24304) );
  XOR U23432 ( .A(n25480), .B(n25481), .Z(n24302) );
  XNOR U23433 ( .A(n25482), .B(n25483), .Z(n25481) );
  NOR U23434 ( .A(n25484), .B(n25483), .Z(n25482) );
  XOR U23435 ( .A(n25485), .B(n25486), .Z(n25480) );
  NOR U23436 ( .A(n25487), .B(n25478), .Z(n25486) );
  NOR U23437 ( .A(n25488), .B(n25479), .Z(n25485) );
  XOR U23438 ( .A(n25489), .B(n25490), .Z(n24295) );
  XOR U23439 ( .A(n25491), .B(n25492), .Z(n24293) );
  XNOR U23440 ( .A(n25493), .B(n25494), .Z(n25492) );
  NOR U23441 ( .A(n25495), .B(n25494), .Z(n25493) );
  XOR U23442 ( .A(n25496), .B(n25497), .Z(n25491) );
  NOR U23443 ( .A(n25498), .B(n25489), .Z(n25497) );
  NOR U23444 ( .A(n25499), .B(n25490), .Z(n25496) );
  XOR U23445 ( .A(n25500), .B(n25501), .Z(n24286) );
  XOR U23446 ( .A(n25502), .B(n25503), .Z(n24284) );
  XNOR U23447 ( .A(n25504), .B(n25505), .Z(n25503) );
  NOR U23448 ( .A(n25506), .B(n25505), .Z(n25504) );
  XOR U23449 ( .A(n25507), .B(n25508), .Z(n25502) );
  NOR U23450 ( .A(n25509), .B(n25500), .Z(n25508) );
  NOR U23451 ( .A(n25510), .B(n25501), .Z(n25507) );
  XOR U23452 ( .A(n25511), .B(n25512), .Z(n24277) );
  XOR U23453 ( .A(n25513), .B(n25514), .Z(n24275) );
  XNOR U23454 ( .A(n25515), .B(n25516), .Z(n25514) );
  NOR U23455 ( .A(n25517), .B(n25516), .Z(n25515) );
  XOR U23456 ( .A(n25518), .B(n25519), .Z(n25513) );
  NOR U23457 ( .A(n25520), .B(n25511), .Z(n25519) );
  NOR U23458 ( .A(n25521), .B(n25512), .Z(n25518) );
  XOR U23459 ( .A(n25522), .B(n25523), .Z(n24268) );
  XOR U23460 ( .A(n25524), .B(n25525), .Z(n24266) );
  XNOR U23461 ( .A(n25526), .B(n25527), .Z(n25525) );
  NOR U23462 ( .A(n25528), .B(n25527), .Z(n25526) );
  XOR U23463 ( .A(n25529), .B(n25530), .Z(n25524) );
  NOR U23464 ( .A(n25531), .B(n25522), .Z(n25530) );
  NOR U23465 ( .A(n25532), .B(n25523), .Z(n25529) );
  XOR U23466 ( .A(n24263), .B(n24261), .Z(n24264) );
  XOR U23467 ( .A(n25533), .B(n25534), .Z(n22960) );
  AND U23468 ( .A(n47), .B(n25533), .Z(n25534) );
  XOR U23469 ( .A(n25535), .B(n25536), .Z(n22963) );
  AND U23470 ( .A(n25537), .B(n25538), .Z(n25536) );
  XNOR U23471 ( .A(n25535), .B(n50), .Z(n25538) );
  XNOR U23472 ( .A(n24249), .B(n22979), .Z(n50) );
  XNOR U23473 ( .A(n22980), .B(n22977), .Z(n22979) );
  XNOR U23474 ( .A(n22978), .B(n22973), .Z(n22977) );
  XOR U23475 ( .A(n22974), .B(n22994), .Z(n22973) );
  XOR U23476 ( .A(n25539), .B(n22992), .Z(n22994) );
  XNOR U23477 ( .A(n22993), .B(n24247), .Z(n22992) );
  XNOR U23478 ( .A(n24248), .B(n24246), .Z(n24247) );
  XNOR U23479 ( .A(n22989), .B(n24243), .Z(n24246) );
  XNOR U23480 ( .A(n22988), .B(n23011), .Z(n24243) );
  XNOR U23481 ( .A(n23006), .B(n24242), .Z(n23011) );
  XNOR U23482 ( .A(n23005), .B(n24237), .Z(n24242) );
  XNOR U23483 ( .A(n23007), .B(n24236), .Z(n24237) );
  XNOR U23484 ( .A(n23010), .B(n24233), .Z(n24236) );
  XNOR U23485 ( .A(n23016), .B(n24232), .Z(n24233) );
  XNOR U23486 ( .A(n24225), .B(n24229), .Z(n24232) );
  XNOR U23487 ( .A(n24224), .B(n24222), .Z(n24229) );
  XNOR U23488 ( .A(n24223), .B(n24221), .Z(n24222) );
  XNOR U23489 ( .A(n23023), .B(n24216), .Z(n24221) );
  XNOR U23490 ( .A(n23022), .B(n24214), .Z(n24216) );
  XNOR U23491 ( .A(n24215), .B(n24210), .Z(n24214) );
  XNOR U23492 ( .A(n24211), .B(n23038), .Z(n24210) );
  XNOR U23493 ( .A(n23033), .B(n24209), .Z(n23038) );
  XNOR U23494 ( .A(n23032), .B(n24204), .Z(n24209) );
  XNOR U23495 ( .A(n23034), .B(n24203), .Z(n24204) );
  XNOR U23496 ( .A(n23037), .B(n24200), .Z(n24203) );
  XNOR U23497 ( .A(n23043), .B(n24199), .Z(n24200) );
  XNOR U23498 ( .A(n24192), .B(n24196), .Z(n24199) );
  XNOR U23499 ( .A(n24191), .B(n24189), .Z(n24196) );
  XNOR U23500 ( .A(n24190), .B(n24188), .Z(n24189) );
  XNOR U23501 ( .A(n23050), .B(n24183), .Z(n24188) );
  XNOR U23502 ( .A(n23049), .B(n24181), .Z(n24183) );
  XNOR U23503 ( .A(n24182), .B(n24177), .Z(n24181) );
  XNOR U23504 ( .A(n24178), .B(n23065), .Z(n24177) );
  XNOR U23505 ( .A(n23060), .B(n24176), .Z(n23065) );
  XNOR U23506 ( .A(n23059), .B(n24171), .Z(n24176) );
  XNOR U23507 ( .A(n23061), .B(n24170), .Z(n24171) );
  XNOR U23508 ( .A(n23064), .B(n24167), .Z(n24170) );
  XNOR U23509 ( .A(n23070), .B(n24166), .Z(n24167) );
  XNOR U23510 ( .A(n24159), .B(n24163), .Z(n24166) );
  XNOR U23511 ( .A(n24158), .B(n24156), .Z(n24163) );
  XNOR U23512 ( .A(n24157), .B(n24155), .Z(n24156) );
  XNOR U23513 ( .A(n23077), .B(n24150), .Z(n24155) );
  XNOR U23514 ( .A(n23076), .B(n24148), .Z(n24150) );
  XNOR U23515 ( .A(n24149), .B(n24144), .Z(n24148) );
  XNOR U23516 ( .A(n24145), .B(n23092), .Z(n24144) );
  XNOR U23517 ( .A(n23087), .B(n24143), .Z(n23092) );
  XNOR U23518 ( .A(n23086), .B(n24138), .Z(n24143) );
  XNOR U23519 ( .A(n23088), .B(n24137), .Z(n24138) );
  XNOR U23520 ( .A(n23091), .B(n24134), .Z(n24137) );
  XNOR U23521 ( .A(n23097), .B(n24133), .Z(n24134) );
  XNOR U23522 ( .A(n24126), .B(n24130), .Z(n24133) );
  XNOR U23523 ( .A(n24125), .B(n24123), .Z(n24130) );
  XNOR U23524 ( .A(n24124), .B(n24122), .Z(n24123) );
  XNOR U23525 ( .A(n23104), .B(n24117), .Z(n24122) );
  XNOR U23526 ( .A(n23103), .B(n24115), .Z(n24117) );
  XNOR U23527 ( .A(n24116), .B(n24111), .Z(n24115) );
  XNOR U23528 ( .A(n24112), .B(n23119), .Z(n24111) );
  XNOR U23529 ( .A(n23114), .B(n24110), .Z(n23119) );
  XNOR U23530 ( .A(n23113), .B(n24105), .Z(n24110) );
  XNOR U23531 ( .A(n23115), .B(n24104), .Z(n24105) );
  XNOR U23532 ( .A(n23118), .B(n24101), .Z(n24104) );
  XNOR U23533 ( .A(n23124), .B(n24100), .Z(n24101) );
  XNOR U23534 ( .A(n24093), .B(n24097), .Z(n24100) );
  XNOR U23535 ( .A(n24092), .B(n24090), .Z(n24097) );
  XNOR U23536 ( .A(n24091), .B(n24089), .Z(n24090) );
  XNOR U23537 ( .A(n23131), .B(n24084), .Z(n24089) );
  XNOR U23538 ( .A(n23130), .B(n24082), .Z(n24084) );
  XNOR U23539 ( .A(n24083), .B(n24078), .Z(n24082) );
  XNOR U23540 ( .A(n24079), .B(n23146), .Z(n24078) );
  XNOR U23541 ( .A(n23141), .B(n24077), .Z(n23146) );
  XNOR U23542 ( .A(n23140), .B(n24072), .Z(n24077) );
  XNOR U23543 ( .A(n23142), .B(n24071), .Z(n24072) );
  XNOR U23544 ( .A(n23145), .B(n24068), .Z(n24071) );
  XNOR U23545 ( .A(n23151), .B(n24067), .Z(n24068) );
  XNOR U23546 ( .A(n24060), .B(n24064), .Z(n24067) );
  XNOR U23547 ( .A(n24059), .B(n24057), .Z(n24064) );
  XNOR U23548 ( .A(n24058), .B(n24056), .Z(n24057) );
  XNOR U23549 ( .A(n23158), .B(n24051), .Z(n24056) );
  XNOR U23550 ( .A(n23157), .B(n24049), .Z(n24051) );
  XNOR U23551 ( .A(n24050), .B(n24045), .Z(n24049) );
  XNOR U23552 ( .A(n24046), .B(n23173), .Z(n24045) );
  XNOR U23553 ( .A(n23168), .B(n24044), .Z(n23173) );
  XNOR U23554 ( .A(n23167), .B(n24039), .Z(n24044) );
  XNOR U23555 ( .A(n23169), .B(n24038), .Z(n24039) );
  XNOR U23556 ( .A(n23172), .B(n24035), .Z(n24038) );
  XNOR U23557 ( .A(n23178), .B(n24034), .Z(n24035) );
  XNOR U23558 ( .A(n24027), .B(n24031), .Z(n24034) );
  XNOR U23559 ( .A(n24026), .B(n24024), .Z(n24031) );
  XNOR U23560 ( .A(n24025), .B(n24023), .Z(n24024) );
  XNOR U23561 ( .A(n23185), .B(n24018), .Z(n24023) );
  XNOR U23562 ( .A(n23184), .B(n24016), .Z(n24018) );
  XNOR U23563 ( .A(n24017), .B(n24012), .Z(n24016) );
  XNOR U23564 ( .A(n24013), .B(n23200), .Z(n24012) );
  XNOR U23565 ( .A(n23195), .B(n24011), .Z(n23200) );
  XNOR U23566 ( .A(n23194), .B(n24006), .Z(n24011) );
  XNOR U23567 ( .A(n23196), .B(n24005), .Z(n24006) );
  XNOR U23568 ( .A(n23199), .B(n24002), .Z(n24005) );
  XNOR U23569 ( .A(n23205), .B(n24001), .Z(n24002) );
  XNOR U23570 ( .A(n23994), .B(n23998), .Z(n24001) );
  XNOR U23571 ( .A(n23993), .B(n23991), .Z(n23998) );
  XNOR U23572 ( .A(n23992), .B(n23990), .Z(n23991) );
  XNOR U23573 ( .A(n23212), .B(n23985), .Z(n23990) );
  XNOR U23574 ( .A(n23211), .B(n23983), .Z(n23985) );
  XNOR U23575 ( .A(n23984), .B(n23979), .Z(n23983) );
  XNOR U23576 ( .A(n23980), .B(n23227), .Z(n23979) );
  XNOR U23577 ( .A(n23222), .B(n23978), .Z(n23227) );
  XNOR U23578 ( .A(n23221), .B(n23973), .Z(n23978) );
  XNOR U23579 ( .A(n23223), .B(n23972), .Z(n23973) );
  XNOR U23580 ( .A(n23226), .B(n23969), .Z(n23972) );
  XNOR U23581 ( .A(n23232), .B(n23968), .Z(n23969) );
  XNOR U23582 ( .A(n23961), .B(n23965), .Z(n23968) );
  XNOR U23583 ( .A(n23960), .B(n23958), .Z(n23965) );
  XNOR U23584 ( .A(n23959), .B(n23957), .Z(n23958) );
  XNOR U23585 ( .A(n23239), .B(n23952), .Z(n23957) );
  XNOR U23586 ( .A(n23238), .B(n23950), .Z(n23952) );
  XNOR U23587 ( .A(n23951), .B(n23946), .Z(n23950) );
  XNOR U23588 ( .A(n23947), .B(n23254), .Z(n23946) );
  XNOR U23589 ( .A(n23249), .B(n23945), .Z(n23254) );
  XNOR U23590 ( .A(n23248), .B(n23940), .Z(n23945) );
  XNOR U23591 ( .A(n23250), .B(n23939), .Z(n23940) );
  XNOR U23592 ( .A(n23253), .B(n23936), .Z(n23939) );
  XNOR U23593 ( .A(n23259), .B(n23935), .Z(n23936) );
  XNOR U23594 ( .A(n23928), .B(n23932), .Z(n23935) );
  XNOR U23595 ( .A(n23927), .B(n23925), .Z(n23932) );
  XNOR U23596 ( .A(n23926), .B(n23924), .Z(n23925) );
  XNOR U23597 ( .A(n23266), .B(n23919), .Z(n23924) );
  XNOR U23598 ( .A(n23265), .B(n23917), .Z(n23919) );
  XNOR U23599 ( .A(n23918), .B(n23913), .Z(n23917) );
  XNOR U23600 ( .A(n23914), .B(n23281), .Z(n23913) );
  XNOR U23601 ( .A(n23276), .B(n23912), .Z(n23281) );
  XNOR U23602 ( .A(n23275), .B(n23907), .Z(n23912) );
  XNOR U23603 ( .A(n23277), .B(n23906), .Z(n23907) );
  XNOR U23604 ( .A(n23280), .B(n23903), .Z(n23906) );
  XNOR U23605 ( .A(n23286), .B(n23902), .Z(n23903) );
  XNOR U23606 ( .A(n23895), .B(n23899), .Z(n23902) );
  XNOR U23607 ( .A(n23894), .B(n23892), .Z(n23899) );
  XNOR U23608 ( .A(n23893), .B(n23891), .Z(n23892) );
  XNOR U23609 ( .A(n23293), .B(n23886), .Z(n23891) );
  XNOR U23610 ( .A(n23292), .B(n23884), .Z(n23886) );
  XNOR U23611 ( .A(n23885), .B(n23880), .Z(n23884) );
  XNOR U23612 ( .A(n23881), .B(n23308), .Z(n23880) );
  XNOR U23613 ( .A(n23303), .B(n23879), .Z(n23308) );
  XNOR U23614 ( .A(n23302), .B(n23874), .Z(n23879) );
  XNOR U23615 ( .A(n23304), .B(n23873), .Z(n23874) );
  XNOR U23616 ( .A(n23307), .B(n23870), .Z(n23873) );
  XNOR U23617 ( .A(n23313), .B(n23869), .Z(n23870) );
  XNOR U23618 ( .A(n23862), .B(n23866), .Z(n23869) );
  XNOR U23619 ( .A(n23861), .B(n23859), .Z(n23866) );
  XNOR U23620 ( .A(n23860), .B(n23858), .Z(n23859) );
  XNOR U23621 ( .A(n23320), .B(n23853), .Z(n23858) );
  XNOR U23622 ( .A(n23319), .B(n23851), .Z(n23853) );
  XNOR U23623 ( .A(n23852), .B(n23847), .Z(n23851) );
  XNOR U23624 ( .A(n23848), .B(n23335), .Z(n23847) );
  XNOR U23625 ( .A(n23330), .B(n23846), .Z(n23335) );
  XNOR U23626 ( .A(n23329), .B(n23841), .Z(n23846) );
  XNOR U23627 ( .A(n23331), .B(n23840), .Z(n23841) );
  XNOR U23628 ( .A(n23334), .B(n23837), .Z(n23840) );
  XNOR U23629 ( .A(n23340), .B(n23836), .Z(n23837) );
  XNOR U23630 ( .A(n23829), .B(n23833), .Z(n23836) );
  XNOR U23631 ( .A(n23828), .B(n23826), .Z(n23833) );
  XNOR U23632 ( .A(n23827), .B(n23825), .Z(n23826) );
  XNOR U23633 ( .A(n23347), .B(n23820), .Z(n23825) );
  XNOR U23634 ( .A(n23346), .B(n23818), .Z(n23820) );
  XNOR U23635 ( .A(n23819), .B(n23814), .Z(n23818) );
  XNOR U23636 ( .A(n23815), .B(n23362), .Z(n23814) );
  XNOR U23637 ( .A(n23357), .B(n23813), .Z(n23362) );
  XNOR U23638 ( .A(n23356), .B(n23808), .Z(n23813) );
  XNOR U23639 ( .A(n23358), .B(n23807), .Z(n23808) );
  XNOR U23640 ( .A(n23361), .B(n23804), .Z(n23807) );
  XNOR U23641 ( .A(n23367), .B(n23803), .Z(n23804) );
  XNOR U23642 ( .A(n23796), .B(n23800), .Z(n23803) );
  XNOR U23643 ( .A(n23795), .B(n23793), .Z(n23800) );
  XNOR U23644 ( .A(n23794), .B(n23792), .Z(n23793) );
  XNOR U23645 ( .A(n23374), .B(n23787), .Z(n23792) );
  XNOR U23646 ( .A(n23373), .B(n23785), .Z(n23787) );
  XNOR U23647 ( .A(n23786), .B(n23781), .Z(n23785) );
  XNOR U23648 ( .A(n23782), .B(n23389), .Z(n23781) );
  XNOR U23649 ( .A(n23384), .B(n23780), .Z(n23389) );
  XNOR U23650 ( .A(n23383), .B(n23775), .Z(n23780) );
  XNOR U23651 ( .A(n23385), .B(n23774), .Z(n23775) );
  XNOR U23652 ( .A(n23388), .B(n23771), .Z(n23774) );
  XNOR U23653 ( .A(n23394), .B(n23770), .Z(n23771) );
  XNOR U23654 ( .A(n23763), .B(n23767), .Z(n23770) );
  XNOR U23655 ( .A(n23762), .B(n23760), .Z(n23767) );
  XNOR U23656 ( .A(n23761), .B(n23759), .Z(n23760) );
  XNOR U23657 ( .A(n23401), .B(n23754), .Z(n23759) );
  XNOR U23658 ( .A(n23400), .B(n23752), .Z(n23754) );
  XNOR U23659 ( .A(n23753), .B(n23748), .Z(n23752) );
  XNOR U23660 ( .A(n23749), .B(n23416), .Z(n23748) );
  XNOR U23661 ( .A(n23411), .B(n23747), .Z(n23416) );
  XNOR U23662 ( .A(n23410), .B(n23742), .Z(n23747) );
  XNOR U23663 ( .A(n23412), .B(n23741), .Z(n23742) );
  XNOR U23664 ( .A(n23415), .B(n23738), .Z(n23741) );
  XNOR U23665 ( .A(n23421), .B(n23737), .Z(n23738) );
  XNOR U23666 ( .A(n23730), .B(n23734), .Z(n23737) );
  XNOR U23667 ( .A(n23729), .B(n23727), .Z(n23734) );
  XNOR U23668 ( .A(n23728), .B(n23726), .Z(n23727) );
  XNOR U23669 ( .A(n23428), .B(n23721), .Z(n23726) );
  XNOR U23670 ( .A(n23427), .B(n23719), .Z(n23721) );
  XNOR U23671 ( .A(n23720), .B(n23715), .Z(n23719) );
  XNOR U23672 ( .A(n23716), .B(n23443), .Z(n23715) );
  XNOR U23673 ( .A(n23438), .B(n23714), .Z(n23443) );
  XNOR U23674 ( .A(n23437), .B(n23709), .Z(n23714) );
  XNOR U23675 ( .A(n23439), .B(n23708), .Z(n23709) );
  XNOR U23676 ( .A(n23442), .B(n23705), .Z(n23708) );
  XNOR U23677 ( .A(n23448), .B(n23704), .Z(n23705) );
  XNOR U23678 ( .A(n23697), .B(n23701), .Z(n23704) );
  XNOR U23679 ( .A(n23696), .B(n23694), .Z(n23701) );
  XNOR U23680 ( .A(n23695), .B(n23693), .Z(n23694) );
  XNOR U23681 ( .A(n23455), .B(n23688), .Z(n23693) );
  XNOR U23682 ( .A(n23454), .B(n23686), .Z(n23688) );
  XNOR U23683 ( .A(n23687), .B(n23682), .Z(n23686) );
  XNOR U23684 ( .A(n23683), .B(n23470), .Z(n23682) );
  XNOR U23685 ( .A(n23465), .B(n23681), .Z(n23470) );
  XNOR U23686 ( .A(n23464), .B(n23676), .Z(n23681) );
  XNOR U23687 ( .A(n23466), .B(n23675), .Z(n23676) );
  XNOR U23688 ( .A(n23469), .B(n23672), .Z(n23675) );
  XNOR U23689 ( .A(n23475), .B(n23671), .Z(n23672) );
  XNOR U23690 ( .A(n23664), .B(n23668), .Z(n23671) );
  XNOR U23691 ( .A(n23663), .B(n23661), .Z(n23668) );
  XNOR U23692 ( .A(n23662), .B(n23660), .Z(n23661) );
  XNOR U23693 ( .A(n23482), .B(n23655), .Z(n23660) );
  XNOR U23694 ( .A(n23481), .B(n23653), .Z(n23655) );
  XNOR U23695 ( .A(n23654), .B(n23649), .Z(n23653) );
  XNOR U23696 ( .A(n23650), .B(n23497), .Z(n23649) );
  XNOR U23697 ( .A(n23492), .B(n23648), .Z(n23497) );
  XNOR U23698 ( .A(n23491), .B(n23643), .Z(n23648) );
  XNOR U23699 ( .A(n23493), .B(n23642), .Z(n23643) );
  XNOR U23700 ( .A(n23496), .B(n23639), .Z(n23642) );
  XNOR U23701 ( .A(n23502), .B(n23638), .Z(n23639) );
  XNOR U23702 ( .A(n23631), .B(n23635), .Z(n23638) );
  XNOR U23703 ( .A(n23630), .B(n23628), .Z(n23635) );
  XNOR U23704 ( .A(n23629), .B(n23627), .Z(n23628) );
  XNOR U23705 ( .A(n23509), .B(n23622), .Z(n23627) );
  XNOR U23706 ( .A(n23508), .B(n23620), .Z(n23622) );
  XNOR U23707 ( .A(n23621), .B(n23616), .Z(n23620) );
  XNOR U23708 ( .A(n23617), .B(n23524), .Z(n23616) );
  XNOR U23709 ( .A(n23519), .B(n23615), .Z(n23524) );
  XNOR U23710 ( .A(n23518), .B(n23610), .Z(n23615) );
  XNOR U23711 ( .A(n23520), .B(n23609), .Z(n23610) );
  XNOR U23712 ( .A(n23523), .B(n23606), .Z(n23609) );
  XNOR U23713 ( .A(n23529), .B(n23605), .Z(n23606) );
  XNOR U23714 ( .A(n23598), .B(n23602), .Z(n23605) );
  XNOR U23715 ( .A(n23597), .B(n23595), .Z(n23602) );
  XNOR U23716 ( .A(n23596), .B(n23594), .Z(n23595) );
  XNOR U23717 ( .A(n23536), .B(n23589), .Z(n23594) );
  XNOR U23718 ( .A(n23535), .B(n23587), .Z(n23589) );
  XNOR U23719 ( .A(n23588), .B(n23583), .Z(n23587) );
  XNOR U23720 ( .A(n23584), .B(n23551), .Z(n23583) );
  XNOR U23721 ( .A(n23546), .B(n23582), .Z(n23551) );
  XNOR U23722 ( .A(n23545), .B(n23577), .Z(n23582) );
  XNOR U23723 ( .A(n23547), .B(n23576), .Z(n23577) );
  XNOR U23724 ( .A(n23550), .B(n23573), .Z(n23576) );
  XNOR U23725 ( .A(n23556), .B(n23572), .Z(n23573) );
  XNOR U23726 ( .A(n23559), .B(n23569), .Z(n23572) );
  XNOR U23727 ( .A(n23558), .B(n23566), .Z(n23569) );
  XOR U23728 ( .A(n23567), .B(n23565), .Z(n23566) );
  XNOR U23729 ( .A(n25540), .B(n25541), .Z(n23565) );
  XOR U23730 ( .A(n25542), .B(n25543), .Z(n25541) );
  XOR U23731 ( .A(n25544), .B(n25545), .Z(n25543) );
  NOR U23732 ( .A(n25546), .B(n25547), .Z(n25545) );
  NOR U23733 ( .A(n25548), .B(n25549), .Z(n25544) );
  NOR U23734 ( .A(n25550), .B(n25551), .Z(n25542) );
  XOR U23735 ( .A(n25552), .B(n25553), .Z(n25540) );
  XOR U23736 ( .A(n25554), .B(n25555), .Z(n25553) );
  XOR U23737 ( .A(n25556), .B(n25557), .Z(n25555) );
  XNOR U23738 ( .A(n25558), .B(n25559), .Z(n25557) );
  XOR U23739 ( .A(n25560), .B(n25561), .Z(n25559) );
  XOR U23740 ( .A(n25562), .B(n25563), .Z(n25561) );
  XOR U23741 ( .A(n25564), .B(n25565), .Z(n25563) );
  XOR U23742 ( .A(n25566), .B(n25567), .Z(n25562) );
  XOR U23743 ( .A(n25568), .B(n25569), .Z(n25567) );
  XOR U23744 ( .A(n25570), .B(n25571), .Z(n25569) );
  XOR U23745 ( .A(n25572), .B(n25573), .Z(n25571) );
  XOR U23746 ( .A(n25574), .B(n25575), .Z(n25573) );
  XNOR U23747 ( .A(n25576), .B(n25577), .Z(n25572) );
  XNOR U23748 ( .A(n25578), .B(n25579), .Z(n25577) );
  NOR U23749 ( .A(n25580), .B(n25575), .Z(n25578) );
  XOR U23750 ( .A(n25581), .B(n25582), .Z(n25570) );
  XOR U23751 ( .A(n25583), .B(n25584), .Z(n25582) );
  XNOR U23752 ( .A(n25585), .B(n25586), .Z(n25584) );
  XOR U23753 ( .A(n25587), .B(n25588), .Z(n25586) );
  XOR U23754 ( .A(n25589), .B(n25590), .Z(n25588) );
  XOR U23755 ( .A(n25591), .B(n25592), .Z(n25590) );
  XOR U23756 ( .A(n25593), .B(n25594), .Z(n25589) );
  XOR U23757 ( .A(n25595), .B(n25596), .Z(n25594) );
  XOR U23758 ( .A(n25597), .B(n25598), .Z(n25596) );
  XOR U23759 ( .A(n25599), .B(n25600), .Z(n25598) );
  XOR U23760 ( .A(n25601), .B(n25602), .Z(n25600) );
  XNOR U23761 ( .A(n25603), .B(n25604), .Z(n25599) );
  XNOR U23762 ( .A(n25605), .B(n25606), .Z(n25604) );
  NOR U23763 ( .A(n25607), .B(n25602), .Z(n25605) );
  XOR U23764 ( .A(n25608), .B(n25609), .Z(n25597) );
  XOR U23765 ( .A(n25610), .B(n25611), .Z(n25609) );
  XNOR U23766 ( .A(n25612), .B(n25613), .Z(n25611) );
  XOR U23767 ( .A(n25614), .B(n25615), .Z(n25613) );
  XOR U23768 ( .A(n25616), .B(n25617), .Z(n25615) );
  XOR U23769 ( .A(n25618), .B(n25619), .Z(n25617) );
  XOR U23770 ( .A(n25620), .B(n25621), .Z(n25616) );
  XOR U23771 ( .A(n25622), .B(n25623), .Z(n25621) );
  XOR U23772 ( .A(n25624), .B(n25625), .Z(n25623) );
  XOR U23773 ( .A(n25626), .B(n25627), .Z(n25625) );
  XOR U23774 ( .A(n25628), .B(n25629), .Z(n25627) );
  XNOR U23775 ( .A(n25630), .B(n25631), .Z(n25626) );
  XNOR U23776 ( .A(n25632), .B(n25633), .Z(n25631) );
  NOR U23777 ( .A(n25634), .B(n25629), .Z(n25632) );
  XOR U23778 ( .A(n25635), .B(n25636), .Z(n25624) );
  XOR U23779 ( .A(n25637), .B(n25638), .Z(n25636) );
  XNOR U23780 ( .A(n25639), .B(n25640), .Z(n25638) );
  XOR U23781 ( .A(n25641), .B(n25642), .Z(n25640) );
  XOR U23782 ( .A(n25643), .B(n25644), .Z(n25642) );
  XOR U23783 ( .A(n25645), .B(n25646), .Z(n25644) );
  XOR U23784 ( .A(n25647), .B(n25648), .Z(n25643) );
  XOR U23785 ( .A(n25649), .B(n25650), .Z(n25648) );
  XOR U23786 ( .A(n25651), .B(n25652), .Z(n25650) );
  XOR U23787 ( .A(n25653), .B(n25654), .Z(n25652) );
  XOR U23788 ( .A(n25655), .B(n25656), .Z(n25654) );
  XNOR U23789 ( .A(n25657), .B(n25658), .Z(n25653) );
  XNOR U23790 ( .A(n25659), .B(n25660), .Z(n25658) );
  NOR U23791 ( .A(n25661), .B(n25656), .Z(n25659) );
  XOR U23792 ( .A(n25662), .B(n25663), .Z(n25651) );
  XOR U23793 ( .A(n25664), .B(n25665), .Z(n25663) );
  XNOR U23794 ( .A(n25666), .B(n25667), .Z(n25665) );
  XOR U23795 ( .A(n25668), .B(n25669), .Z(n25667) );
  XOR U23796 ( .A(n25670), .B(n25671), .Z(n25669) );
  XOR U23797 ( .A(n25672), .B(n25673), .Z(n25671) );
  XOR U23798 ( .A(n25674), .B(n25675), .Z(n25670) );
  XOR U23799 ( .A(n25676), .B(n25677), .Z(n25675) );
  XOR U23800 ( .A(n25678), .B(n25679), .Z(n25677) );
  XOR U23801 ( .A(n25680), .B(n25681), .Z(n25679) );
  XOR U23802 ( .A(n25682), .B(n25683), .Z(n25681) );
  XNOR U23803 ( .A(n25684), .B(n25685), .Z(n25680) );
  XNOR U23804 ( .A(n25686), .B(n25687), .Z(n25685) );
  NOR U23805 ( .A(n25688), .B(n25683), .Z(n25686) );
  XOR U23806 ( .A(n25689), .B(n25690), .Z(n25678) );
  XOR U23807 ( .A(n25691), .B(n25692), .Z(n25690) );
  XNOR U23808 ( .A(n25693), .B(n25694), .Z(n25692) );
  XOR U23809 ( .A(n25695), .B(n25696), .Z(n25694) );
  XOR U23810 ( .A(n25697), .B(n25698), .Z(n25696) );
  XOR U23811 ( .A(n25699), .B(n25700), .Z(n25698) );
  XOR U23812 ( .A(n25701), .B(n25702), .Z(n25697) );
  XOR U23813 ( .A(n25703), .B(n25704), .Z(n25702) );
  XOR U23814 ( .A(n25705), .B(n25706), .Z(n25704) );
  XOR U23815 ( .A(n25707), .B(n25708), .Z(n25706) );
  XOR U23816 ( .A(n25709), .B(n25710), .Z(n25708) );
  XNOR U23817 ( .A(n25711), .B(n25712), .Z(n25707) );
  XNOR U23818 ( .A(n25713), .B(n25714), .Z(n25712) );
  NOR U23819 ( .A(n25715), .B(n25710), .Z(n25713) );
  XOR U23820 ( .A(n25716), .B(n25717), .Z(n25705) );
  XOR U23821 ( .A(n25718), .B(n25719), .Z(n25717) );
  XNOR U23822 ( .A(n25720), .B(n25721), .Z(n25719) );
  XOR U23823 ( .A(n25722), .B(n25723), .Z(n25721) );
  XOR U23824 ( .A(n25724), .B(n25725), .Z(n25723) );
  XOR U23825 ( .A(n25726), .B(n25727), .Z(n25725) );
  XOR U23826 ( .A(n25728), .B(n25729), .Z(n25724) );
  XOR U23827 ( .A(n25730), .B(n25731), .Z(n25729) );
  XOR U23828 ( .A(n25732), .B(n25733), .Z(n25731) );
  XOR U23829 ( .A(n25734), .B(n25735), .Z(n25733) );
  XOR U23830 ( .A(n25736), .B(n25737), .Z(n25735) );
  XNOR U23831 ( .A(n25738), .B(n25739), .Z(n25734) );
  XNOR U23832 ( .A(n25740), .B(n25741), .Z(n25739) );
  NOR U23833 ( .A(n25742), .B(n25737), .Z(n25740) );
  XOR U23834 ( .A(n25743), .B(n25744), .Z(n25732) );
  XOR U23835 ( .A(n25745), .B(n25746), .Z(n25744) );
  XNOR U23836 ( .A(n25747), .B(n25748), .Z(n25746) );
  XOR U23837 ( .A(n25749), .B(n25750), .Z(n25748) );
  XOR U23838 ( .A(n25751), .B(n25752), .Z(n25750) );
  XOR U23839 ( .A(n25753), .B(n25754), .Z(n25752) );
  XOR U23840 ( .A(n25755), .B(n25756), .Z(n25751) );
  XOR U23841 ( .A(n25757), .B(n25758), .Z(n25756) );
  XOR U23842 ( .A(n25759), .B(n25760), .Z(n25758) );
  XOR U23843 ( .A(n25761), .B(n25762), .Z(n25760) );
  XOR U23844 ( .A(n25763), .B(n25764), .Z(n25762) );
  XNOR U23845 ( .A(n25765), .B(n25766), .Z(n25761) );
  XNOR U23846 ( .A(n25767), .B(n25768), .Z(n25766) );
  NOR U23847 ( .A(n25769), .B(n25764), .Z(n25767) );
  XOR U23848 ( .A(n25770), .B(n25771), .Z(n25759) );
  XOR U23849 ( .A(n25772), .B(n25773), .Z(n25771) );
  XNOR U23850 ( .A(n25774), .B(n25775), .Z(n25773) );
  XOR U23851 ( .A(n25776), .B(n25777), .Z(n25775) );
  XOR U23852 ( .A(n25778), .B(n25779), .Z(n25777) );
  XOR U23853 ( .A(n25780), .B(n25781), .Z(n25779) );
  XOR U23854 ( .A(n25782), .B(n25783), .Z(n25778) );
  XOR U23855 ( .A(n25784), .B(n25785), .Z(n25783) );
  XOR U23856 ( .A(n25786), .B(n25787), .Z(n25785) );
  XOR U23857 ( .A(n25788), .B(n25789), .Z(n25787) );
  XOR U23858 ( .A(n25790), .B(n25791), .Z(n25789) );
  XNOR U23859 ( .A(n25792), .B(n25793), .Z(n25788) );
  XNOR U23860 ( .A(n25794), .B(n25795), .Z(n25793) );
  NOR U23861 ( .A(n25796), .B(n25791), .Z(n25794) );
  XOR U23862 ( .A(n25797), .B(n25798), .Z(n25786) );
  XOR U23863 ( .A(n25799), .B(n25800), .Z(n25798) );
  XNOR U23864 ( .A(n25801), .B(n25802), .Z(n25800) );
  XOR U23865 ( .A(n25803), .B(n25804), .Z(n25802) );
  XOR U23866 ( .A(n25805), .B(n25806), .Z(n25804) );
  XOR U23867 ( .A(n25807), .B(n25808), .Z(n25806) );
  XOR U23868 ( .A(n25809), .B(n25810), .Z(n25805) );
  XOR U23869 ( .A(n25811), .B(n25812), .Z(n25810) );
  XOR U23870 ( .A(n25813), .B(n25814), .Z(n25812) );
  XOR U23871 ( .A(n25815), .B(n25816), .Z(n25814) );
  XOR U23872 ( .A(n25817), .B(n25818), .Z(n25816) );
  XNOR U23873 ( .A(n25819), .B(n25820), .Z(n25815) );
  XNOR U23874 ( .A(n25821), .B(n25822), .Z(n25820) );
  NOR U23875 ( .A(n25823), .B(n25818), .Z(n25821) );
  XOR U23876 ( .A(n25824), .B(n25825), .Z(n25813) );
  XOR U23877 ( .A(n25826), .B(n25827), .Z(n25825) );
  XOR U23878 ( .A(n25828), .B(n25829), .Z(n25827) );
  XOR U23879 ( .A(n25830), .B(n25831), .Z(n25826) );
  XOR U23880 ( .A(n25832), .B(n25833), .Z(n25824) );
  XOR U23881 ( .A(n25834), .B(n25835), .Z(n25833) );
  AND U23882 ( .A(n25836), .B(n25837), .Z(n25835) );
  XOR U23883 ( .A(n25838), .B(n25829), .Z(n25836) );
  XOR U23884 ( .A(n25839), .B(n25840), .Z(n25829) );
  NOR U23885 ( .A(n25838), .B(n25839), .Z(n25840) );
  NOR U23886 ( .A(n25841), .B(n25830), .Z(n25834) );
  XOR U23887 ( .A(n25842), .B(n25843), .Z(n25832) );
  NOR U23888 ( .A(n25844), .B(n25831), .Z(n25843) );
  NOR U23889 ( .A(n25845), .B(n25828), .Z(n25842) );
  XOR U23890 ( .A(n25846), .B(n25847), .Z(n25811) );
  NOR U23891 ( .A(n25848), .B(n25822), .Z(n25847) );
  NOR U23892 ( .A(n25849), .B(n25819), .Z(n25846) );
  XOR U23893 ( .A(n25850), .B(n25851), .Z(n25809) );
  XOR U23894 ( .A(n25852), .B(n25853), .Z(n25851) );
  NOR U23895 ( .A(n25854), .B(n25817), .Z(n25853) );
  NOR U23896 ( .A(n25855), .B(n25856), .Z(n25852) );
  XOR U23897 ( .A(n25857), .B(n25858), .Z(n25850) );
  NOR U23898 ( .A(n25859), .B(n25860), .Z(n25858) );
  NOR U23899 ( .A(n25861), .B(n25807), .Z(n25857) );
  XOR U23900 ( .A(n25862), .B(n25863), .Z(n25803) );
  XOR U23901 ( .A(n25856), .B(n25860), .Z(n25863) );
  XOR U23902 ( .A(n25864), .B(n25865), .Z(n25862) );
  NOR U23903 ( .A(n25866), .B(n25808), .Z(n25865) );
  NOR U23904 ( .A(n25867), .B(n25868), .Z(n25864) );
  XOR U23905 ( .A(n25869), .B(n25870), .Z(n25799) );
  XOR U23906 ( .A(n25871), .B(n25872), .Z(n25797) );
  XNOR U23907 ( .A(n25873), .B(n25868), .Z(n25872) );
  NOR U23908 ( .A(n25874), .B(n25869), .Z(n25873) );
  XOR U23909 ( .A(n25875), .B(n25876), .Z(n25871) );
  NOR U23910 ( .A(n25877), .B(n25870), .Z(n25876) );
  NOR U23911 ( .A(n25878), .B(n25801), .Z(n25875) );
  XOR U23912 ( .A(n25879), .B(n25880), .Z(n25784) );
  NOR U23913 ( .A(n25881), .B(n25795), .Z(n25880) );
  NOR U23914 ( .A(n25882), .B(n25792), .Z(n25879) );
  XOR U23915 ( .A(n25883), .B(n25884), .Z(n25782) );
  XOR U23916 ( .A(n25885), .B(n25886), .Z(n25884) );
  NOR U23917 ( .A(n25887), .B(n25790), .Z(n25886) );
  NOR U23918 ( .A(n25888), .B(n25889), .Z(n25885) );
  XOR U23919 ( .A(n25890), .B(n25891), .Z(n25883) );
  NOR U23920 ( .A(n25892), .B(n25893), .Z(n25891) );
  NOR U23921 ( .A(n25894), .B(n25780), .Z(n25890) );
  XOR U23922 ( .A(n25895), .B(n25896), .Z(n25776) );
  XOR U23923 ( .A(n25889), .B(n25893), .Z(n25896) );
  XOR U23924 ( .A(n25897), .B(n25898), .Z(n25895) );
  NOR U23925 ( .A(n25899), .B(n25781), .Z(n25898) );
  NOR U23926 ( .A(n25900), .B(n25901), .Z(n25897) );
  XOR U23927 ( .A(n25902), .B(n25903), .Z(n25772) );
  XOR U23928 ( .A(n25904), .B(n25905), .Z(n25770) );
  XNOR U23929 ( .A(n25906), .B(n25901), .Z(n25905) );
  NOR U23930 ( .A(n25907), .B(n25902), .Z(n25906) );
  XOR U23931 ( .A(n25908), .B(n25909), .Z(n25904) );
  NOR U23932 ( .A(n25910), .B(n25903), .Z(n25909) );
  NOR U23933 ( .A(n25911), .B(n25774), .Z(n25908) );
  XOR U23934 ( .A(n25912), .B(n25913), .Z(n25757) );
  NOR U23935 ( .A(n25914), .B(n25768), .Z(n25913) );
  NOR U23936 ( .A(n25915), .B(n25765), .Z(n25912) );
  XOR U23937 ( .A(n25916), .B(n25917), .Z(n25755) );
  XOR U23938 ( .A(n25918), .B(n25919), .Z(n25917) );
  NOR U23939 ( .A(n25920), .B(n25763), .Z(n25919) );
  NOR U23940 ( .A(n25921), .B(n25922), .Z(n25918) );
  XOR U23941 ( .A(n25923), .B(n25924), .Z(n25916) );
  NOR U23942 ( .A(n25925), .B(n25926), .Z(n25924) );
  NOR U23943 ( .A(n25927), .B(n25753), .Z(n25923) );
  XOR U23944 ( .A(n25928), .B(n25929), .Z(n25749) );
  XOR U23945 ( .A(n25922), .B(n25926), .Z(n25929) );
  XOR U23946 ( .A(n25930), .B(n25931), .Z(n25928) );
  NOR U23947 ( .A(n25932), .B(n25754), .Z(n25931) );
  NOR U23948 ( .A(n25933), .B(n25934), .Z(n25930) );
  XOR U23949 ( .A(n25935), .B(n25936), .Z(n25745) );
  XOR U23950 ( .A(n25937), .B(n25938), .Z(n25743) );
  XNOR U23951 ( .A(n25939), .B(n25934), .Z(n25938) );
  NOR U23952 ( .A(n25940), .B(n25935), .Z(n25939) );
  XOR U23953 ( .A(n25941), .B(n25942), .Z(n25937) );
  NOR U23954 ( .A(n25943), .B(n25936), .Z(n25942) );
  NOR U23955 ( .A(n25944), .B(n25747), .Z(n25941) );
  XOR U23956 ( .A(n25945), .B(n25946), .Z(n25730) );
  NOR U23957 ( .A(n25947), .B(n25741), .Z(n25946) );
  NOR U23958 ( .A(n25948), .B(n25738), .Z(n25945) );
  XOR U23959 ( .A(n25949), .B(n25950), .Z(n25728) );
  XOR U23960 ( .A(n25951), .B(n25952), .Z(n25950) );
  NOR U23961 ( .A(n25953), .B(n25736), .Z(n25952) );
  NOR U23962 ( .A(n25954), .B(n25955), .Z(n25951) );
  XOR U23963 ( .A(n25956), .B(n25957), .Z(n25949) );
  NOR U23964 ( .A(n25958), .B(n25959), .Z(n25957) );
  NOR U23965 ( .A(n25960), .B(n25726), .Z(n25956) );
  XOR U23966 ( .A(n25961), .B(n25962), .Z(n25722) );
  XOR U23967 ( .A(n25955), .B(n25959), .Z(n25962) );
  XOR U23968 ( .A(n25963), .B(n25964), .Z(n25961) );
  NOR U23969 ( .A(n25965), .B(n25727), .Z(n25964) );
  NOR U23970 ( .A(n25966), .B(n25967), .Z(n25963) );
  XOR U23971 ( .A(n25968), .B(n25969), .Z(n25718) );
  XOR U23972 ( .A(n25970), .B(n25971), .Z(n25716) );
  XNOR U23973 ( .A(n25972), .B(n25967), .Z(n25971) );
  NOR U23974 ( .A(n25973), .B(n25968), .Z(n25972) );
  XOR U23975 ( .A(n25974), .B(n25975), .Z(n25970) );
  NOR U23976 ( .A(n25976), .B(n25969), .Z(n25975) );
  NOR U23977 ( .A(n25977), .B(n25720), .Z(n25974) );
  XOR U23978 ( .A(n25978), .B(n25979), .Z(n25703) );
  NOR U23979 ( .A(n25980), .B(n25714), .Z(n25979) );
  NOR U23980 ( .A(n25981), .B(n25711), .Z(n25978) );
  XOR U23981 ( .A(n25982), .B(n25983), .Z(n25701) );
  XOR U23982 ( .A(n25984), .B(n25985), .Z(n25983) );
  NOR U23983 ( .A(n25986), .B(n25709), .Z(n25985) );
  NOR U23984 ( .A(n25987), .B(n25988), .Z(n25984) );
  XOR U23985 ( .A(n25989), .B(n25990), .Z(n25982) );
  NOR U23986 ( .A(n25991), .B(n25992), .Z(n25990) );
  NOR U23987 ( .A(n25993), .B(n25699), .Z(n25989) );
  XOR U23988 ( .A(n25994), .B(n25995), .Z(n25695) );
  XOR U23989 ( .A(n25988), .B(n25992), .Z(n25995) );
  XOR U23990 ( .A(n25996), .B(n25997), .Z(n25994) );
  NOR U23991 ( .A(n25998), .B(n25700), .Z(n25997) );
  NOR U23992 ( .A(n25999), .B(n26000), .Z(n25996) );
  XOR U23993 ( .A(n26001), .B(n26002), .Z(n25691) );
  XOR U23994 ( .A(n26003), .B(n26004), .Z(n25689) );
  XNOR U23995 ( .A(n26005), .B(n26000), .Z(n26004) );
  NOR U23996 ( .A(n26006), .B(n26001), .Z(n26005) );
  XOR U23997 ( .A(n26007), .B(n26008), .Z(n26003) );
  NOR U23998 ( .A(n26009), .B(n26002), .Z(n26008) );
  NOR U23999 ( .A(n26010), .B(n25693), .Z(n26007) );
  XOR U24000 ( .A(n26011), .B(n26012), .Z(n25676) );
  NOR U24001 ( .A(n26013), .B(n25687), .Z(n26012) );
  NOR U24002 ( .A(n26014), .B(n25684), .Z(n26011) );
  XOR U24003 ( .A(n26015), .B(n26016), .Z(n25674) );
  XOR U24004 ( .A(n26017), .B(n26018), .Z(n26016) );
  NOR U24005 ( .A(n26019), .B(n25682), .Z(n26018) );
  NOR U24006 ( .A(n26020), .B(n26021), .Z(n26017) );
  XOR U24007 ( .A(n26022), .B(n26023), .Z(n26015) );
  NOR U24008 ( .A(n26024), .B(n26025), .Z(n26023) );
  NOR U24009 ( .A(n26026), .B(n25672), .Z(n26022) );
  XOR U24010 ( .A(n26027), .B(n26028), .Z(n25668) );
  XOR U24011 ( .A(n26021), .B(n26025), .Z(n26028) );
  XOR U24012 ( .A(n26029), .B(n26030), .Z(n26027) );
  NOR U24013 ( .A(n26031), .B(n25673), .Z(n26030) );
  NOR U24014 ( .A(n26032), .B(n26033), .Z(n26029) );
  XOR U24015 ( .A(n26034), .B(n26035), .Z(n25664) );
  XOR U24016 ( .A(n26036), .B(n26037), .Z(n25662) );
  XNOR U24017 ( .A(n26038), .B(n26033), .Z(n26037) );
  NOR U24018 ( .A(n26039), .B(n26034), .Z(n26038) );
  XOR U24019 ( .A(n26040), .B(n26041), .Z(n26036) );
  NOR U24020 ( .A(n26042), .B(n26035), .Z(n26041) );
  NOR U24021 ( .A(n26043), .B(n25666), .Z(n26040) );
  XOR U24022 ( .A(n26044), .B(n26045), .Z(n25649) );
  NOR U24023 ( .A(n26046), .B(n25660), .Z(n26045) );
  NOR U24024 ( .A(n26047), .B(n25657), .Z(n26044) );
  XOR U24025 ( .A(n26048), .B(n26049), .Z(n25647) );
  XOR U24026 ( .A(n26050), .B(n26051), .Z(n26049) );
  NOR U24027 ( .A(n26052), .B(n25655), .Z(n26051) );
  NOR U24028 ( .A(n26053), .B(n26054), .Z(n26050) );
  XOR U24029 ( .A(n26055), .B(n26056), .Z(n26048) );
  NOR U24030 ( .A(n26057), .B(n26058), .Z(n26056) );
  NOR U24031 ( .A(n26059), .B(n25645), .Z(n26055) );
  XOR U24032 ( .A(n26060), .B(n26061), .Z(n25641) );
  XOR U24033 ( .A(n26054), .B(n26058), .Z(n26061) );
  XOR U24034 ( .A(n26062), .B(n26063), .Z(n26060) );
  NOR U24035 ( .A(n26064), .B(n25646), .Z(n26063) );
  NOR U24036 ( .A(n26065), .B(n26066), .Z(n26062) );
  XOR U24037 ( .A(n26067), .B(n26068), .Z(n25637) );
  XOR U24038 ( .A(n26069), .B(n26070), .Z(n25635) );
  XNOR U24039 ( .A(n26071), .B(n26066), .Z(n26070) );
  NOR U24040 ( .A(n26072), .B(n26067), .Z(n26071) );
  XOR U24041 ( .A(n26073), .B(n26074), .Z(n26069) );
  NOR U24042 ( .A(n26075), .B(n26068), .Z(n26074) );
  NOR U24043 ( .A(n26076), .B(n25639), .Z(n26073) );
  XOR U24044 ( .A(n26077), .B(n26078), .Z(n25622) );
  NOR U24045 ( .A(n26079), .B(n25633), .Z(n26078) );
  NOR U24046 ( .A(n26080), .B(n25630), .Z(n26077) );
  XOR U24047 ( .A(n26081), .B(n26082), .Z(n25620) );
  XOR U24048 ( .A(n26083), .B(n26084), .Z(n26082) );
  NOR U24049 ( .A(n26085), .B(n25628), .Z(n26084) );
  NOR U24050 ( .A(n26086), .B(n26087), .Z(n26083) );
  XOR U24051 ( .A(n26088), .B(n26089), .Z(n26081) );
  NOR U24052 ( .A(n26090), .B(n26091), .Z(n26089) );
  NOR U24053 ( .A(n26092), .B(n25618), .Z(n26088) );
  XOR U24054 ( .A(n26093), .B(n26094), .Z(n25614) );
  XOR U24055 ( .A(n26087), .B(n26091), .Z(n26094) );
  XOR U24056 ( .A(n26095), .B(n26096), .Z(n26093) );
  NOR U24057 ( .A(n26097), .B(n25619), .Z(n26096) );
  NOR U24058 ( .A(n26098), .B(n26099), .Z(n26095) );
  XOR U24059 ( .A(n26100), .B(n26101), .Z(n25610) );
  XOR U24060 ( .A(n26102), .B(n26103), .Z(n25608) );
  XNOR U24061 ( .A(n26104), .B(n26099), .Z(n26103) );
  NOR U24062 ( .A(n26105), .B(n26100), .Z(n26104) );
  XOR U24063 ( .A(n26106), .B(n26107), .Z(n26102) );
  NOR U24064 ( .A(n26108), .B(n26101), .Z(n26107) );
  NOR U24065 ( .A(n26109), .B(n25612), .Z(n26106) );
  XOR U24066 ( .A(n26110), .B(n26111), .Z(n25595) );
  NOR U24067 ( .A(n26112), .B(n25606), .Z(n26111) );
  NOR U24068 ( .A(n26113), .B(n25603), .Z(n26110) );
  XOR U24069 ( .A(n26114), .B(n26115), .Z(n25593) );
  XOR U24070 ( .A(n26116), .B(n26117), .Z(n26115) );
  NOR U24071 ( .A(n26118), .B(n25601), .Z(n26117) );
  NOR U24072 ( .A(n26119), .B(n26120), .Z(n26116) );
  XOR U24073 ( .A(n26121), .B(n26122), .Z(n26114) );
  NOR U24074 ( .A(n26123), .B(n26124), .Z(n26122) );
  NOR U24075 ( .A(n26125), .B(n25591), .Z(n26121) );
  XOR U24076 ( .A(n26126), .B(n26127), .Z(n25587) );
  XOR U24077 ( .A(n26120), .B(n26124), .Z(n26127) );
  XOR U24078 ( .A(n26128), .B(n26129), .Z(n26126) );
  NOR U24079 ( .A(n26130), .B(n25592), .Z(n26129) );
  NOR U24080 ( .A(n26131), .B(n26132), .Z(n26128) );
  XOR U24081 ( .A(n26133), .B(n26134), .Z(n25583) );
  XOR U24082 ( .A(n26135), .B(n26136), .Z(n25581) );
  XNOR U24083 ( .A(n26137), .B(n26132), .Z(n26136) );
  NOR U24084 ( .A(n26138), .B(n26133), .Z(n26137) );
  XOR U24085 ( .A(n26139), .B(n26140), .Z(n26135) );
  NOR U24086 ( .A(n26141), .B(n26134), .Z(n26140) );
  NOR U24087 ( .A(n26142), .B(n25585), .Z(n26139) );
  XOR U24088 ( .A(n26143), .B(n26144), .Z(n25568) );
  NOR U24089 ( .A(n26145), .B(n25579), .Z(n26144) );
  NOR U24090 ( .A(n26146), .B(n25576), .Z(n26143) );
  XOR U24091 ( .A(n26147), .B(n26148), .Z(n25566) );
  XOR U24092 ( .A(n26149), .B(n26150), .Z(n26148) );
  NOR U24093 ( .A(n26151), .B(n25574), .Z(n26150) );
  NOR U24094 ( .A(n26152), .B(n26153), .Z(n26149) );
  XOR U24095 ( .A(n26154), .B(n26155), .Z(n26147) );
  NOR U24096 ( .A(n26156), .B(n26157), .Z(n26155) );
  NOR U24097 ( .A(n26158), .B(n25564), .Z(n26154) );
  XOR U24098 ( .A(n26159), .B(n26160), .Z(n25560) );
  XOR U24099 ( .A(n26153), .B(n26157), .Z(n26160) );
  XOR U24100 ( .A(n26161), .B(n26162), .Z(n26159) );
  NOR U24101 ( .A(n26163), .B(n25565), .Z(n26162) );
  NOR U24102 ( .A(n26164), .B(n26165), .Z(n26161) );
  XOR U24103 ( .A(n26166), .B(n26167), .Z(n25556) );
  XOR U24104 ( .A(n26168), .B(n26169), .Z(n25554) );
  XNOR U24105 ( .A(n26170), .B(n26165), .Z(n26169) );
  NOR U24106 ( .A(n26171), .B(n26166), .Z(n26170) );
  XOR U24107 ( .A(n26172), .B(n26173), .Z(n26168) );
  NOR U24108 ( .A(n26174), .B(n26167), .Z(n26173) );
  NOR U24109 ( .A(n26175), .B(n25558), .Z(n26172) );
  XOR U24110 ( .A(n26176), .B(n26177), .Z(n25552) );
  XNOR U24111 ( .A(n25547), .B(n26178), .Z(n26177) );
  XNOR U24112 ( .A(n26179), .B(n25551), .Z(n26178) );
  NOR U24113 ( .A(n26180), .B(n26181), .Z(n26179) );
  XNOR U24114 ( .A(n26181), .B(n25549), .Z(n26176) );
  XOR U24115 ( .A(n26182), .B(n26183), .Z(n23567) );
  NOR U24116 ( .A(n26184), .B(n26182), .Z(n26183) );
  XOR U24117 ( .A(n26185), .B(n26186), .Z(n23558) );
  NOR U24118 ( .A(n26187), .B(n26185), .Z(n26186) );
  XOR U24119 ( .A(n26188), .B(n26189), .Z(n23559) );
  NOR U24120 ( .A(n26190), .B(n26188), .Z(n26189) );
  XOR U24121 ( .A(n26191), .B(n26192), .Z(n23556) );
  NOR U24122 ( .A(n26193), .B(n26191), .Z(n26192) );
  XOR U24123 ( .A(n26194), .B(n26195), .Z(n23550) );
  NOR U24124 ( .A(n26196), .B(n26194), .Z(n26195) );
  XOR U24125 ( .A(n26197), .B(n26198), .Z(n23547) );
  NOR U24126 ( .A(n26199), .B(n26197), .Z(n26198) );
  XOR U24127 ( .A(n26200), .B(n26201), .Z(n23545) );
  NOR U24128 ( .A(n26202), .B(n26200), .Z(n26201) );
  XOR U24129 ( .A(n26203), .B(n26204), .Z(n23546) );
  NOR U24130 ( .A(n26205), .B(n26203), .Z(n26204) );
  XOR U24131 ( .A(n26206), .B(n26207), .Z(n23584) );
  NOR U24132 ( .A(n26208), .B(n26206), .Z(n26207) );
  XOR U24133 ( .A(n26209), .B(n26210), .Z(n23588) );
  NOR U24134 ( .A(n26211), .B(n26209), .Z(n26210) );
  XOR U24135 ( .A(n26212), .B(n26213), .Z(n23535) );
  NOR U24136 ( .A(n26214), .B(n26212), .Z(n26213) );
  XOR U24137 ( .A(n26215), .B(n26216), .Z(n23536) );
  NOR U24138 ( .A(n26217), .B(n26215), .Z(n26216) );
  XOR U24139 ( .A(n26218), .B(n26219), .Z(n23596) );
  NOR U24140 ( .A(n26220), .B(n26218), .Z(n26219) );
  XOR U24141 ( .A(n26221), .B(n26222), .Z(n23597) );
  NOR U24142 ( .A(n26223), .B(n26221), .Z(n26222) );
  XOR U24143 ( .A(n26224), .B(n26225), .Z(n23598) );
  NOR U24144 ( .A(n26226), .B(n26224), .Z(n26225) );
  XOR U24145 ( .A(n26227), .B(n26228), .Z(n23529) );
  NOR U24146 ( .A(n26229), .B(n26227), .Z(n26228) );
  XOR U24147 ( .A(n26230), .B(n26231), .Z(n23523) );
  NOR U24148 ( .A(n26232), .B(n26230), .Z(n26231) );
  XOR U24149 ( .A(n26233), .B(n26234), .Z(n23520) );
  NOR U24150 ( .A(n26235), .B(n26233), .Z(n26234) );
  XOR U24151 ( .A(n26236), .B(n26237), .Z(n23518) );
  NOR U24152 ( .A(n26238), .B(n26236), .Z(n26237) );
  XOR U24153 ( .A(n26239), .B(n26240), .Z(n23519) );
  NOR U24154 ( .A(n26241), .B(n26239), .Z(n26240) );
  XOR U24155 ( .A(n26242), .B(n26243), .Z(n23617) );
  NOR U24156 ( .A(n26244), .B(n26242), .Z(n26243) );
  XOR U24157 ( .A(n26245), .B(n26246), .Z(n23621) );
  NOR U24158 ( .A(n26247), .B(n26245), .Z(n26246) );
  XOR U24159 ( .A(n26248), .B(n26249), .Z(n23508) );
  NOR U24160 ( .A(n26250), .B(n26248), .Z(n26249) );
  XOR U24161 ( .A(n26251), .B(n26252), .Z(n23509) );
  NOR U24162 ( .A(n26253), .B(n26251), .Z(n26252) );
  XOR U24163 ( .A(n26254), .B(n26255), .Z(n23629) );
  NOR U24164 ( .A(n26256), .B(n26254), .Z(n26255) );
  XOR U24165 ( .A(n26257), .B(n26258), .Z(n23630) );
  NOR U24166 ( .A(n26259), .B(n26257), .Z(n26258) );
  XOR U24167 ( .A(n26260), .B(n26261), .Z(n23631) );
  NOR U24168 ( .A(n26262), .B(n26260), .Z(n26261) );
  XOR U24169 ( .A(n26263), .B(n26264), .Z(n23502) );
  NOR U24170 ( .A(n26265), .B(n26263), .Z(n26264) );
  XOR U24171 ( .A(n26266), .B(n26267), .Z(n23496) );
  NOR U24172 ( .A(n26268), .B(n26266), .Z(n26267) );
  XOR U24173 ( .A(n26269), .B(n26270), .Z(n23493) );
  NOR U24174 ( .A(n26271), .B(n26269), .Z(n26270) );
  XOR U24175 ( .A(n26272), .B(n26273), .Z(n23491) );
  NOR U24176 ( .A(n26274), .B(n26272), .Z(n26273) );
  XOR U24177 ( .A(n26275), .B(n26276), .Z(n23492) );
  NOR U24178 ( .A(n26277), .B(n26275), .Z(n26276) );
  XOR U24179 ( .A(n26278), .B(n26279), .Z(n23650) );
  NOR U24180 ( .A(n26280), .B(n26278), .Z(n26279) );
  XOR U24181 ( .A(n26281), .B(n26282), .Z(n23654) );
  NOR U24182 ( .A(n26283), .B(n26281), .Z(n26282) );
  XOR U24183 ( .A(n26284), .B(n26285), .Z(n23481) );
  NOR U24184 ( .A(n26286), .B(n26284), .Z(n26285) );
  XOR U24185 ( .A(n26287), .B(n26288), .Z(n23482) );
  NOR U24186 ( .A(n26289), .B(n26287), .Z(n26288) );
  XOR U24187 ( .A(n26290), .B(n26291), .Z(n23662) );
  NOR U24188 ( .A(n26292), .B(n26290), .Z(n26291) );
  XOR U24189 ( .A(n26293), .B(n26294), .Z(n23663) );
  NOR U24190 ( .A(n26295), .B(n26293), .Z(n26294) );
  XOR U24191 ( .A(n26296), .B(n26297), .Z(n23664) );
  NOR U24192 ( .A(n26298), .B(n26296), .Z(n26297) );
  XOR U24193 ( .A(n26299), .B(n26300), .Z(n23475) );
  NOR U24194 ( .A(n26301), .B(n26299), .Z(n26300) );
  XOR U24195 ( .A(n26302), .B(n26303), .Z(n23469) );
  NOR U24196 ( .A(n26304), .B(n26302), .Z(n26303) );
  XOR U24197 ( .A(n26305), .B(n26306), .Z(n23466) );
  NOR U24198 ( .A(n26307), .B(n26305), .Z(n26306) );
  XOR U24199 ( .A(n26308), .B(n26309), .Z(n23464) );
  NOR U24200 ( .A(n26310), .B(n26308), .Z(n26309) );
  XOR U24201 ( .A(n26311), .B(n26312), .Z(n23465) );
  NOR U24202 ( .A(n26313), .B(n26311), .Z(n26312) );
  XOR U24203 ( .A(n26314), .B(n26315), .Z(n23683) );
  NOR U24204 ( .A(n26316), .B(n26314), .Z(n26315) );
  XOR U24205 ( .A(n26317), .B(n26318), .Z(n23687) );
  NOR U24206 ( .A(n26319), .B(n26317), .Z(n26318) );
  XOR U24207 ( .A(n26320), .B(n26321), .Z(n23454) );
  NOR U24208 ( .A(n26322), .B(n26320), .Z(n26321) );
  XOR U24209 ( .A(n26323), .B(n26324), .Z(n23455) );
  NOR U24210 ( .A(n26325), .B(n26323), .Z(n26324) );
  XOR U24211 ( .A(n26326), .B(n26327), .Z(n23695) );
  NOR U24212 ( .A(n26328), .B(n26326), .Z(n26327) );
  XOR U24213 ( .A(n26329), .B(n26330), .Z(n23696) );
  NOR U24214 ( .A(n26331), .B(n26329), .Z(n26330) );
  XOR U24215 ( .A(n26332), .B(n26333), .Z(n23697) );
  NOR U24216 ( .A(n26334), .B(n26332), .Z(n26333) );
  XOR U24217 ( .A(n26335), .B(n26336), .Z(n23448) );
  NOR U24218 ( .A(n26337), .B(n26335), .Z(n26336) );
  XOR U24219 ( .A(n26338), .B(n26339), .Z(n23442) );
  NOR U24220 ( .A(n26340), .B(n26338), .Z(n26339) );
  XOR U24221 ( .A(n26341), .B(n26342), .Z(n23439) );
  NOR U24222 ( .A(n26343), .B(n26341), .Z(n26342) );
  XOR U24223 ( .A(n26344), .B(n26345), .Z(n23437) );
  NOR U24224 ( .A(n26346), .B(n26344), .Z(n26345) );
  XOR U24225 ( .A(n26347), .B(n26348), .Z(n23438) );
  NOR U24226 ( .A(n26349), .B(n26347), .Z(n26348) );
  XOR U24227 ( .A(n26350), .B(n26351), .Z(n23716) );
  NOR U24228 ( .A(n26352), .B(n26350), .Z(n26351) );
  XOR U24229 ( .A(n26353), .B(n26354), .Z(n23720) );
  NOR U24230 ( .A(n26355), .B(n26353), .Z(n26354) );
  XOR U24231 ( .A(n26356), .B(n26357), .Z(n23427) );
  NOR U24232 ( .A(n26358), .B(n26356), .Z(n26357) );
  XOR U24233 ( .A(n26359), .B(n26360), .Z(n23428) );
  NOR U24234 ( .A(n26361), .B(n26359), .Z(n26360) );
  XOR U24235 ( .A(n26362), .B(n26363), .Z(n23728) );
  NOR U24236 ( .A(n26364), .B(n26362), .Z(n26363) );
  XOR U24237 ( .A(n26365), .B(n26366), .Z(n23729) );
  NOR U24238 ( .A(n26367), .B(n26365), .Z(n26366) );
  XOR U24239 ( .A(n26368), .B(n26369), .Z(n23730) );
  NOR U24240 ( .A(n26370), .B(n26368), .Z(n26369) );
  XOR U24241 ( .A(n26371), .B(n26372), .Z(n23421) );
  NOR U24242 ( .A(n26373), .B(n26371), .Z(n26372) );
  XOR U24243 ( .A(n26374), .B(n26375), .Z(n23415) );
  NOR U24244 ( .A(n26376), .B(n26374), .Z(n26375) );
  XOR U24245 ( .A(n26377), .B(n26378), .Z(n23412) );
  NOR U24246 ( .A(n26379), .B(n26377), .Z(n26378) );
  XOR U24247 ( .A(n26380), .B(n26381), .Z(n23410) );
  NOR U24248 ( .A(n26382), .B(n26380), .Z(n26381) );
  XOR U24249 ( .A(n26383), .B(n26384), .Z(n23411) );
  NOR U24250 ( .A(n26385), .B(n26383), .Z(n26384) );
  XOR U24251 ( .A(n26386), .B(n26387), .Z(n23749) );
  NOR U24252 ( .A(n26388), .B(n26386), .Z(n26387) );
  XOR U24253 ( .A(n26389), .B(n26390), .Z(n23753) );
  NOR U24254 ( .A(n26391), .B(n26389), .Z(n26390) );
  XOR U24255 ( .A(n26392), .B(n26393), .Z(n23400) );
  NOR U24256 ( .A(n26394), .B(n26392), .Z(n26393) );
  XOR U24257 ( .A(n26395), .B(n26396), .Z(n23401) );
  NOR U24258 ( .A(n26397), .B(n26395), .Z(n26396) );
  XOR U24259 ( .A(n26398), .B(n26399), .Z(n23761) );
  NOR U24260 ( .A(n26400), .B(n26398), .Z(n26399) );
  XOR U24261 ( .A(n26401), .B(n26402), .Z(n23762) );
  NOR U24262 ( .A(n26403), .B(n26401), .Z(n26402) );
  XOR U24263 ( .A(n26404), .B(n26405), .Z(n23763) );
  NOR U24264 ( .A(n26406), .B(n26404), .Z(n26405) );
  XOR U24265 ( .A(n26407), .B(n26408), .Z(n23394) );
  NOR U24266 ( .A(n26409), .B(n26407), .Z(n26408) );
  XOR U24267 ( .A(n26410), .B(n26411), .Z(n23388) );
  NOR U24268 ( .A(n26412), .B(n26410), .Z(n26411) );
  XOR U24269 ( .A(n26413), .B(n26414), .Z(n23385) );
  NOR U24270 ( .A(n26415), .B(n26413), .Z(n26414) );
  XOR U24271 ( .A(n26416), .B(n26417), .Z(n23383) );
  NOR U24272 ( .A(n26418), .B(n26416), .Z(n26417) );
  XOR U24273 ( .A(n26419), .B(n26420), .Z(n23384) );
  NOR U24274 ( .A(n26421), .B(n26419), .Z(n26420) );
  XOR U24275 ( .A(n26422), .B(n26423), .Z(n23782) );
  NOR U24276 ( .A(n26424), .B(n26422), .Z(n26423) );
  XOR U24277 ( .A(n26425), .B(n26426), .Z(n23786) );
  NOR U24278 ( .A(n26427), .B(n26425), .Z(n26426) );
  XOR U24279 ( .A(n26428), .B(n26429), .Z(n23373) );
  NOR U24280 ( .A(n26430), .B(n26428), .Z(n26429) );
  XOR U24281 ( .A(n26431), .B(n26432), .Z(n23374) );
  NOR U24282 ( .A(n26433), .B(n26431), .Z(n26432) );
  XOR U24283 ( .A(n26434), .B(n26435), .Z(n23794) );
  NOR U24284 ( .A(n26436), .B(n26434), .Z(n26435) );
  XOR U24285 ( .A(n26437), .B(n26438), .Z(n23795) );
  NOR U24286 ( .A(n26439), .B(n26437), .Z(n26438) );
  XOR U24287 ( .A(n26440), .B(n26441), .Z(n23796) );
  NOR U24288 ( .A(n26442), .B(n26440), .Z(n26441) );
  XOR U24289 ( .A(n26443), .B(n26444), .Z(n23367) );
  NOR U24290 ( .A(n26445), .B(n26443), .Z(n26444) );
  XOR U24291 ( .A(n26446), .B(n26447), .Z(n23361) );
  NOR U24292 ( .A(n26448), .B(n26446), .Z(n26447) );
  XOR U24293 ( .A(n26449), .B(n26450), .Z(n23358) );
  NOR U24294 ( .A(n26451), .B(n26449), .Z(n26450) );
  XOR U24295 ( .A(n26452), .B(n26453), .Z(n23356) );
  NOR U24296 ( .A(n26454), .B(n26452), .Z(n26453) );
  XOR U24297 ( .A(n26455), .B(n26456), .Z(n23357) );
  NOR U24298 ( .A(n26457), .B(n26455), .Z(n26456) );
  XOR U24299 ( .A(n26458), .B(n26459), .Z(n23815) );
  NOR U24300 ( .A(n26460), .B(n26458), .Z(n26459) );
  XOR U24301 ( .A(n26461), .B(n26462), .Z(n23819) );
  NOR U24302 ( .A(n26463), .B(n26461), .Z(n26462) );
  XOR U24303 ( .A(n26464), .B(n26465), .Z(n23346) );
  NOR U24304 ( .A(n26466), .B(n26464), .Z(n26465) );
  XOR U24305 ( .A(n26467), .B(n26468), .Z(n23347) );
  NOR U24306 ( .A(n26469), .B(n26467), .Z(n26468) );
  XOR U24307 ( .A(n26470), .B(n26471), .Z(n23827) );
  NOR U24308 ( .A(n26472), .B(n26470), .Z(n26471) );
  XOR U24309 ( .A(n26473), .B(n26474), .Z(n23828) );
  NOR U24310 ( .A(n26475), .B(n26473), .Z(n26474) );
  XOR U24311 ( .A(n26476), .B(n26477), .Z(n23829) );
  NOR U24312 ( .A(n26478), .B(n26476), .Z(n26477) );
  XOR U24313 ( .A(n26479), .B(n26480), .Z(n23340) );
  NOR U24314 ( .A(n26481), .B(n26479), .Z(n26480) );
  XOR U24315 ( .A(n26482), .B(n26483), .Z(n23334) );
  NOR U24316 ( .A(n26484), .B(n26482), .Z(n26483) );
  XOR U24317 ( .A(n26485), .B(n26486), .Z(n23331) );
  NOR U24318 ( .A(n26487), .B(n26485), .Z(n26486) );
  XOR U24319 ( .A(n26488), .B(n26489), .Z(n23329) );
  NOR U24320 ( .A(n26490), .B(n26488), .Z(n26489) );
  XOR U24321 ( .A(n26491), .B(n26492), .Z(n23330) );
  NOR U24322 ( .A(n26493), .B(n26491), .Z(n26492) );
  XOR U24323 ( .A(n26494), .B(n26495), .Z(n23848) );
  NOR U24324 ( .A(n26496), .B(n26494), .Z(n26495) );
  XOR U24325 ( .A(n26497), .B(n26498), .Z(n23852) );
  NOR U24326 ( .A(n26499), .B(n26497), .Z(n26498) );
  XOR U24327 ( .A(n26500), .B(n26501), .Z(n23319) );
  NOR U24328 ( .A(n26502), .B(n26500), .Z(n26501) );
  XOR U24329 ( .A(n26503), .B(n26504), .Z(n23320) );
  NOR U24330 ( .A(n26505), .B(n26503), .Z(n26504) );
  XOR U24331 ( .A(n26506), .B(n26507), .Z(n23860) );
  NOR U24332 ( .A(n26508), .B(n26506), .Z(n26507) );
  XOR U24333 ( .A(n26509), .B(n26510), .Z(n23861) );
  NOR U24334 ( .A(n26511), .B(n26509), .Z(n26510) );
  XOR U24335 ( .A(n26512), .B(n26513), .Z(n23862) );
  NOR U24336 ( .A(n26514), .B(n26512), .Z(n26513) );
  XOR U24337 ( .A(n26515), .B(n26516), .Z(n23313) );
  NOR U24338 ( .A(n26517), .B(n26515), .Z(n26516) );
  XOR U24339 ( .A(n26518), .B(n26519), .Z(n23307) );
  NOR U24340 ( .A(n26520), .B(n26518), .Z(n26519) );
  XOR U24341 ( .A(n26521), .B(n26522), .Z(n23304) );
  NOR U24342 ( .A(n26523), .B(n26521), .Z(n26522) );
  XOR U24343 ( .A(n26524), .B(n26525), .Z(n23302) );
  NOR U24344 ( .A(n26526), .B(n26524), .Z(n26525) );
  XOR U24345 ( .A(n26527), .B(n26528), .Z(n23303) );
  NOR U24346 ( .A(n26529), .B(n26527), .Z(n26528) );
  XOR U24347 ( .A(n26530), .B(n26531), .Z(n23881) );
  NOR U24348 ( .A(n26532), .B(n26530), .Z(n26531) );
  XOR U24349 ( .A(n26533), .B(n26534), .Z(n23885) );
  NOR U24350 ( .A(n26535), .B(n26533), .Z(n26534) );
  XOR U24351 ( .A(n26536), .B(n26537), .Z(n23292) );
  NOR U24352 ( .A(n26538), .B(n26536), .Z(n26537) );
  XOR U24353 ( .A(n26539), .B(n26540), .Z(n23293) );
  NOR U24354 ( .A(n26541), .B(n26539), .Z(n26540) );
  XOR U24355 ( .A(n26542), .B(n26543), .Z(n23893) );
  NOR U24356 ( .A(n26544), .B(n26542), .Z(n26543) );
  XOR U24357 ( .A(n26545), .B(n26546), .Z(n23894) );
  NOR U24358 ( .A(n26547), .B(n26545), .Z(n26546) );
  XOR U24359 ( .A(n26548), .B(n26549), .Z(n23895) );
  NOR U24360 ( .A(n26550), .B(n26548), .Z(n26549) );
  XOR U24361 ( .A(n26551), .B(n26552), .Z(n23286) );
  NOR U24362 ( .A(n26553), .B(n26551), .Z(n26552) );
  XOR U24363 ( .A(n26554), .B(n26555), .Z(n23280) );
  NOR U24364 ( .A(n26556), .B(n26554), .Z(n26555) );
  XOR U24365 ( .A(n26557), .B(n26558), .Z(n23277) );
  NOR U24366 ( .A(n26559), .B(n26557), .Z(n26558) );
  XOR U24367 ( .A(n26560), .B(n26561), .Z(n23275) );
  NOR U24368 ( .A(n26562), .B(n26560), .Z(n26561) );
  XOR U24369 ( .A(n26563), .B(n26564), .Z(n23276) );
  NOR U24370 ( .A(n26565), .B(n26563), .Z(n26564) );
  XOR U24371 ( .A(n26566), .B(n26567), .Z(n23914) );
  NOR U24372 ( .A(n26568), .B(n26566), .Z(n26567) );
  XOR U24373 ( .A(n26569), .B(n26570), .Z(n23918) );
  NOR U24374 ( .A(n26571), .B(n26569), .Z(n26570) );
  XOR U24375 ( .A(n26572), .B(n26573), .Z(n23265) );
  NOR U24376 ( .A(n26574), .B(n26572), .Z(n26573) );
  XOR U24377 ( .A(n26575), .B(n26576), .Z(n23266) );
  NOR U24378 ( .A(n26577), .B(n26575), .Z(n26576) );
  XOR U24379 ( .A(n26578), .B(n26579), .Z(n23926) );
  NOR U24380 ( .A(n26580), .B(n26578), .Z(n26579) );
  XOR U24381 ( .A(n26581), .B(n26582), .Z(n23927) );
  NOR U24382 ( .A(n26583), .B(n26581), .Z(n26582) );
  XOR U24383 ( .A(n26584), .B(n26585), .Z(n23928) );
  NOR U24384 ( .A(n26586), .B(n26584), .Z(n26585) );
  XOR U24385 ( .A(n26587), .B(n26588), .Z(n23259) );
  NOR U24386 ( .A(n26589), .B(n26587), .Z(n26588) );
  XOR U24387 ( .A(n26590), .B(n26591), .Z(n23253) );
  NOR U24388 ( .A(n26592), .B(n26590), .Z(n26591) );
  XOR U24389 ( .A(n26593), .B(n26594), .Z(n23250) );
  NOR U24390 ( .A(n26595), .B(n26593), .Z(n26594) );
  XOR U24391 ( .A(n26596), .B(n26597), .Z(n23248) );
  NOR U24392 ( .A(n26598), .B(n26596), .Z(n26597) );
  XOR U24393 ( .A(n26599), .B(n26600), .Z(n23249) );
  NOR U24394 ( .A(n26601), .B(n26599), .Z(n26600) );
  XOR U24395 ( .A(n26602), .B(n26603), .Z(n23947) );
  NOR U24396 ( .A(n26604), .B(n26602), .Z(n26603) );
  XOR U24397 ( .A(n26605), .B(n26606), .Z(n23951) );
  NOR U24398 ( .A(n26607), .B(n26605), .Z(n26606) );
  XOR U24399 ( .A(n26608), .B(n26609), .Z(n23238) );
  NOR U24400 ( .A(n26610), .B(n26608), .Z(n26609) );
  XOR U24401 ( .A(n26611), .B(n26612), .Z(n23239) );
  NOR U24402 ( .A(n26613), .B(n26611), .Z(n26612) );
  XOR U24403 ( .A(n26614), .B(n26615), .Z(n23959) );
  NOR U24404 ( .A(n26616), .B(n26614), .Z(n26615) );
  XOR U24405 ( .A(n26617), .B(n26618), .Z(n23960) );
  NOR U24406 ( .A(n26619), .B(n26617), .Z(n26618) );
  XOR U24407 ( .A(n26620), .B(n26621), .Z(n23961) );
  NOR U24408 ( .A(n26622), .B(n26620), .Z(n26621) );
  XOR U24409 ( .A(n26623), .B(n26624), .Z(n23232) );
  NOR U24410 ( .A(n26625), .B(n26623), .Z(n26624) );
  XOR U24411 ( .A(n26626), .B(n26627), .Z(n23226) );
  NOR U24412 ( .A(n26628), .B(n26626), .Z(n26627) );
  XOR U24413 ( .A(n26629), .B(n26630), .Z(n23223) );
  NOR U24414 ( .A(n26631), .B(n26629), .Z(n26630) );
  XOR U24415 ( .A(n26632), .B(n26633), .Z(n23221) );
  NOR U24416 ( .A(n26634), .B(n26632), .Z(n26633) );
  XOR U24417 ( .A(n26635), .B(n26636), .Z(n23222) );
  NOR U24418 ( .A(n26637), .B(n26635), .Z(n26636) );
  XOR U24419 ( .A(n26638), .B(n26639), .Z(n23980) );
  NOR U24420 ( .A(n26640), .B(n26638), .Z(n26639) );
  XOR U24421 ( .A(n26641), .B(n26642), .Z(n23984) );
  NOR U24422 ( .A(n26643), .B(n26641), .Z(n26642) );
  XOR U24423 ( .A(n26644), .B(n26645), .Z(n23211) );
  NOR U24424 ( .A(n26646), .B(n26644), .Z(n26645) );
  XOR U24425 ( .A(n26647), .B(n26648), .Z(n23212) );
  NOR U24426 ( .A(n26649), .B(n26647), .Z(n26648) );
  XOR U24427 ( .A(n26650), .B(n26651), .Z(n23992) );
  NOR U24428 ( .A(n26652), .B(n26650), .Z(n26651) );
  XOR U24429 ( .A(n26653), .B(n26654), .Z(n23993) );
  NOR U24430 ( .A(n26655), .B(n26653), .Z(n26654) );
  XOR U24431 ( .A(n26656), .B(n26657), .Z(n23994) );
  NOR U24432 ( .A(n26658), .B(n26656), .Z(n26657) );
  XOR U24433 ( .A(n26659), .B(n26660), .Z(n23205) );
  NOR U24434 ( .A(n26661), .B(n26659), .Z(n26660) );
  XOR U24435 ( .A(n26662), .B(n26663), .Z(n23199) );
  NOR U24436 ( .A(n26664), .B(n26662), .Z(n26663) );
  XOR U24437 ( .A(n26665), .B(n26666), .Z(n23196) );
  NOR U24438 ( .A(n26667), .B(n26665), .Z(n26666) );
  XOR U24439 ( .A(n26668), .B(n26669), .Z(n23194) );
  NOR U24440 ( .A(n26670), .B(n26668), .Z(n26669) );
  XOR U24441 ( .A(n26671), .B(n26672), .Z(n23195) );
  NOR U24442 ( .A(n26673), .B(n26671), .Z(n26672) );
  XOR U24443 ( .A(n26674), .B(n26675), .Z(n24013) );
  NOR U24444 ( .A(n26676), .B(n26674), .Z(n26675) );
  XOR U24445 ( .A(n26677), .B(n26678), .Z(n24017) );
  NOR U24446 ( .A(n26679), .B(n26677), .Z(n26678) );
  XOR U24447 ( .A(n26680), .B(n26681), .Z(n23184) );
  NOR U24448 ( .A(n26682), .B(n26680), .Z(n26681) );
  XOR U24449 ( .A(n26683), .B(n26684), .Z(n23185) );
  NOR U24450 ( .A(n26685), .B(n26683), .Z(n26684) );
  XOR U24451 ( .A(n26686), .B(n26687), .Z(n24025) );
  NOR U24452 ( .A(n26688), .B(n26686), .Z(n26687) );
  XOR U24453 ( .A(n26689), .B(n26690), .Z(n24026) );
  NOR U24454 ( .A(n26691), .B(n26689), .Z(n26690) );
  XOR U24455 ( .A(n26692), .B(n26693), .Z(n24027) );
  NOR U24456 ( .A(n26694), .B(n26692), .Z(n26693) );
  XOR U24457 ( .A(n26695), .B(n26696), .Z(n23178) );
  NOR U24458 ( .A(n26697), .B(n26695), .Z(n26696) );
  XOR U24459 ( .A(n26698), .B(n26699), .Z(n23172) );
  NOR U24460 ( .A(n26700), .B(n26698), .Z(n26699) );
  XOR U24461 ( .A(n26701), .B(n26702), .Z(n23169) );
  NOR U24462 ( .A(n26703), .B(n26701), .Z(n26702) );
  XOR U24463 ( .A(n26704), .B(n26705), .Z(n23167) );
  NOR U24464 ( .A(n26706), .B(n26704), .Z(n26705) );
  XOR U24465 ( .A(n26707), .B(n26708), .Z(n23168) );
  NOR U24466 ( .A(n26709), .B(n26707), .Z(n26708) );
  XOR U24467 ( .A(n26710), .B(n26711), .Z(n24046) );
  NOR U24468 ( .A(n26712), .B(n26710), .Z(n26711) );
  XOR U24469 ( .A(n26713), .B(n26714), .Z(n24050) );
  NOR U24470 ( .A(n26715), .B(n26713), .Z(n26714) );
  XOR U24471 ( .A(n26716), .B(n26717), .Z(n23157) );
  NOR U24472 ( .A(n26718), .B(n26716), .Z(n26717) );
  XOR U24473 ( .A(n26719), .B(n26720), .Z(n23158) );
  NOR U24474 ( .A(n26721), .B(n26719), .Z(n26720) );
  XOR U24475 ( .A(n26722), .B(n26723), .Z(n24058) );
  NOR U24476 ( .A(n26724), .B(n26722), .Z(n26723) );
  XOR U24477 ( .A(n26725), .B(n26726), .Z(n24059) );
  NOR U24478 ( .A(n26727), .B(n26725), .Z(n26726) );
  XOR U24479 ( .A(n26728), .B(n26729), .Z(n24060) );
  NOR U24480 ( .A(n26730), .B(n26728), .Z(n26729) );
  XOR U24481 ( .A(n26731), .B(n26732), .Z(n23151) );
  NOR U24482 ( .A(n26733), .B(n26731), .Z(n26732) );
  XOR U24483 ( .A(n26734), .B(n26735), .Z(n23145) );
  NOR U24484 ( .A(n26736), .B(n26734), .Z(n26735) );
  XOR U24485 ( .A(n26737), .B(n26738), .Z(n23142) );
  NOR U24486 ( .A(n26739), .B(n26737), .Z(n26738) );
  XOR U24487 ( .A(n26740), .B(n26741), .Z(n23140) );
  NOR U24488 ( .A(n26742), .B(n26740), .Z(n26741) );
  XOR U24489 ( .A(n26743), .B(n26744), .Z(n23141) );
  NOR U24490 ( .A(n26745), .B(n26743), .Z(n26744) );
  XOR U24491 ( .A(n26746), .B(n26747), .Z(n24079) );
  NOR U24492 ( .A(n26748), .B(n26746), .Z(n26747) );
  XOR U24493 ( .A(n26749), .B(n26750), .Z(n24083) );
  NOR U24494 ( .A(n26751), .B(n26749), .Z(n26750) );
  XOR U24495 ( .A(n26752), .B(n26753), .Z(n23130) );
  NOR U24496 ( .A(n26754), .B(n26752), .Z(n26753) );
  XOR U24497 ( .A(n26755), .B(n26756), .Z(n23131) );
  NOR U24498 ( .A(n26757), .B(n26755), .Z(n26756) );
  XOR U24499 ( .A(n26758), .B(n26759), .Z(n24091) );
  NOR U24500 ( .A(n26760), .B(n26758), .Z(n26759) );
  XOR U24501 ( .A(n26761), .B(n26762), .Z(n24092) );
  NOR U24502 ( .A(n26763), .B(n26761), .Z(n26762) );
  XOR U24503 ( .A(n26764), .B(n26765), .Z(n24093) );
  NOR U24504 ( .A(n26766), .B(n26764), .Z(n26765) );
  XOR U24505 ( .A(n26767), .B(n26768), .Z(n23124) );
  NOR U24506 ( .A(n26769), .B(n26767), .Z(n26768) );
  XOR U24507 ( .A(n26770), .B(n26771), .Z(n23118) );
  NOR U24508 ( .A(n26772), .B(n26770), .Z(n26771) );
  XOR U24509 ( .A(n26773), .B(n26774), .Z(n23115) );
  NOR U24510 ( .A(n26775), .B(n26773), .Z(n26774) );
  XOR U24511 ( .A(n26776), .B(n26777), .Z(n23113) );
  NOR U24512 ( .A(n26778), .B(n26776), .Z(n26777) );
  XOR U24513 ( .A(n26779), .B(n26780), .Z(n23114) );
  NOR U24514 ( .A(n26781), .B(n26779), .Z(n26780) );
  XOR U24515 ( .A(n26782), .B(n26783), .Z(n24112) );
  NOR U24516 ( .A(n26784), .B(n26782), .Z(n26783) );
  XOR U24517 ( .A(n26785), .B(n26786), .Z(n24116) );
  NOR U24518 ( .A(n26787), .B(n26785), .Z(n26786) );
  XOR U24519 ( .A(n26788), .B(n26789), .Z(n23103) );
  NOR U24520 ( .A(n26790), .B(n26788), .Z(n26789) );
  XOR U24521 ( .A(n26791), .B(n26792), .Z(n23104) );
  NOR U24522 ( .A(n26793), .B(n26791), .Z(n26792) );
  XOR U24523 ( .A(n26794), .B(n26795), .Z(n24124) );
  NOR U24524 ( .A(n26796), .B(n26794), .Z(n26795) );
  XOR U24525 ( .A(n26797), .B(n26798), .Z(n24125) );
  NOR U24526 ( .A(n26799), .B(n26797), .Z(n26798) );
  XOR U24527 ( .A(n26800), .B(n26801), .Z(n24126) );
  NOR U24528 ( .A(n26802), .B(n26800), .Z(n26801) );
  XOR U24529 ( .A(n26803), .B(n26804), .Z(n23097) );
  NOR U24530 ( .A(n26805), .B(n26803), .Z(n26804) );
  XOR U24531 ( .A(n26806), .B(n26807), .Z(n23091) );
  NOR U24532 ( .A(n26808), .B(n26806), .Z(n26807) );
  XOR U24533 ( .A(n26809), .B(n26810), .Z(n23088) );
  NOR U24534 ( .A(n26811), .B(n26809), .Z(n26810) );
  XOR U24535 ( .A(n26812), .B(n26813), .Z(n23086) );
  NOR U24536 ( .A(n26814), .B(n26812), .Z(n26813) );
  XOR U24537 ( .A(n26815), .B(n26816), .Z(n23087) );
  NOR U24538 ( .A(n26817), .B(n26815), .Z(n26816) );
  XOR U24539 ( .A(n26818), .B(n26819), .Z(n24145) );
  NOR U24540 ( .A(n26820), .B(n26818), .Z(n26819) );
  XOR U24541 ( .A(n26821), .B(n26822), .Z(n24149) );
  NOR U24542 ( .A(n26823), .B(n26821), .Z(n26822) );
  XOR U24543 ( .A(n26824), .B(n26825), .Z(n23076) );
  NOR U24544 ( .A(n26826), .B(n26824), .Z(n26825) );
  XOR U24545 ( .A(n26827), .B(n26828), .Z(n23077) );
  NOR U24546 ( .A(n26829), .B(n26827), .Z(n26828) );
  XOR U24547 ( .A(n26830), .B(n26831), .Z(n24157) );
  NOR U24548 ( .A(n26832), .B(n26830), .Z(n26831) );
  XOR U24549 ( .A(n26833), .B(n26834), .Z(n24158) );
  NOR U24550 ( .A(n26835), .B(n26833), .Z(n26834) );
  XOR U24551 ( .A(n26836), .B(n26837), .Z(n24159) );
  NOR U24552 ( .A(n26838), .B(n26836), .Z(n26837) );
  XOR U24553 ( .A(n26839), .B(n26840), .Z(n23070) );
  NOR U24554 ( .A(n26841), .B(n26839), .Z(n26840) );
  XOR U24555 ( .A(n26842), .B(n26843), .Z(n23064) );
  NOR U24556 ( .A(n26844), .B(n26842), .Z(n26843) );
  XOR U24557 ( .A(n26845), .B(n26846), .Z(n23061) );
  NOR U24558 ( .A(n26847), .B(n26845), .Z(n26846) );
  XOR U24559 ( .A(n26848), .B(n26849), .Z(n23059) );
  NOR U24560 ( .A(n26850), .B(n26848), .Z(n26849) );
  XOR U24561 ( .A(n26851), .B(n26852), .Z(n23060) );
  NOR U24562 ( .A(n26853), .B(n26851), .Z(n26852) );
  XOR U24563 ( .A(n26854), .B(n26855), .Z(n24178) );
  NOR U24564 ( .A(n26856), .B(n26854), .Z(n26855) );
  XOR U24565 ( .A(n26857), .B(n26858), .Z(n24182) );
  NOR U24566 ( .A(n26859), .B(n26857), .Z(n26858) );
  XOR U24567 ( .A(n26860), .B(n26861), .Z(n23049) );
  NOR U24568 ( .A(n26862), .B(n26860), .Z(n26861) );
  XOR U24569 ( .A(n26863), .B(n26864), .Z(n23050) );
  NOR U24570 ( .A(n26865), .B(n26863), .Z(n26864) );
  XOR U24571 ( .A(n26866), .B(n26867), .Z(n24190) );
  NOR U24572 ( .A(n26868), .B(n26866), .Z(n26867) );
  XOR U24573 ( .A(n26869), .B(n26870), .Z(n24191) );
  NOR U24574 ( .A(n26871), .B(n26869), .Z(n26870) );
  XOR U24575 ( .A(n26872), .B(n26873), .Z(n24192) );
  NOR U24576 ( .A(n26874), .B(n26872), .Z(n26873) );
  XOR U24577 ( .A(n26875), .B(n26876), .Z(n23043) );
  NOR U24578 ( .A(n26877), .B(n26875), .Z(n26876) );
  XOR U24579 ( .A(n26878), .B(n26879), .Z(n23037) );
  NOR U24580 ( .A(n26880), .B(n26878), .Z(n26879) );
  XOR U24581 ( .A(n26881), .B(n26882), .Z(n23034) );
  NOR U24582 ( .A(n26883), .B(n26881), .Z(n26882) );
  XOR U24583 ( .A(n26884), .B(n26885), .Z(n23032) );
  NOR U24584 ( .A(n26886), .B(n26884), .Z(n26885) );
  XOR U24585 ( .A(n26887), .B(n26888), .Z(n23033) );
  NOR U24586 ( .A(n26889), .B(n26887), .Z(n26888) );
  XOR U24587 ( .A(n26890), .B(n26891), .Z(n24211) );
  NOR U24588 ( .A(n26892), .B(n26890), .Z(n26891) );
  XOR U24589 ( .A(n26893), .B(n26894), .Z(n24215) );
  NOR U24590 ( .A(n26895), .B(n26893), .Z(n26894) );
  XOR U24591 ( .A(n26896), .B(n26897), .Z(n23022) );
  NOR U24592 ( .A(n26898), .B(n26896), .Z(n26897) );
  XOR U24593 ( .A(n26899), .B(n26900), .Z(n23023) );
  NOR U24594 ( .A(n26901), .B(n26899), .Z(n26900) );
  XOR U24595 ( .A(n26902), .B(n26903), .Z(n24223) );
  NOR U24596 ( .A(n26904), .B(n26902), .Z(n26903) );
  XOR U24597 ( .A(n26905), .B(n26906), .Z(n24224) );
  NOR U24598 ( .A(n26907), .B(n26905), .Z(n26906) );
  XOR U24599 ( .A(n26908), .B(n26909), .Z(n24225) );
  NOR U24600 ( .A(n26910), .B(n26908), .Z(n26909) );
  XOR U24601 ( .A(n26911), .B(n26912), .Z(n23016) );
  NOR U24602 ( .A(n26913), .B(n26911), .Z(n26912) );
  XOR U24603 ( .A(n26914), .B(n26915), .Z(n23010) );
  NOR U24604 ( .A(n26916), .B(n26914), .Z(n26915) );
  XOR U24605 ( .A(n26917), .B(n26918), .Z(n23007) );
  NOR U24606 ( .A(n26919), .B(n26917), .Z(n26918) );
  XOR U24607 ( .A(n26920), .B(n26921), .Z(n23005) );
  NOR U24608 ( .A(n26922), .B(n26920), .Z(n26921) );
  XOR U24609 ( .A(n26923), .B(n26924), .Z(n23006) );
  NOR U24610 ( .A(n26925), .B(n26923), .Z(n26924) );
  XOR U24611 ( .A(n26926), .B(n26927), .Z(n22988) );
  NOR U24612 ( .A(n26928), .B(n26926), .Z(n26927) );
  XOR U24613 ( .A(n26929), .B(n26930), .Z(n22989) );
  NOR U24614 ( .A(n26931), .B(n26929), .Z(n26930) );
  XOR U24615 ( .A(n26932), .B(n26933), .Z(n24248) );
  NOR U24616 ( .A(n26934), .B(n26932), .Z(n26933) );
  XOR U24617 ( .A(n26935), .B(n26936), .Z(n22993) );
  NOR U24618 ( .A(n26937), .B(n26935), .Z(n26936) );
  IV U24619 ( .A(n22972), .Z(n25539) );
  XNOR U24620 ( .A(n26938), .B(n26939), .Z(n22972) );
  NOR U24621 ( .A(n26940), .B(n26938), .Z(n26939) );
  XOR U24622 ( .A(n26941), .B(n26942), .Z(n22974) );
  NOR U24623 ( .A(n26943), .B(n26941), .Z(n26942) );
  XOR U24624 ( .A(n26944), .B(n26945), .Z(n22978) );
  NOR U24625 ( .A(n26946), .B(n26944), .Z(n26945) );
  XNOR U24626 ( .A(n26947), .B(n26948), .Z(n22980) );
  AND U24627 ( .A(n26949), .B(n26947), .Z(n26948) );
  XNOR U24628 ( .A(n26950), .B(n26951), .Z(n24249) );
  AND U24629 ( .A(n65), .B(n26950), .Z(n26951) );
  XNOR U24630 ( .A(n47), .B(n25535), .Z(n25537) );
  XOR U24631 ( .A(n25533), .B(n24274), .Z(n47) );
  XOR U24632 ( .A(n26952), .B(n24262), .Z(n24274) );
  XOR U24633 ( .A(n24263), .B(n24260), .Z(n24262) );
  XOR U24634 ( .A(n24261), .B(n24257), .Z(n24260) );
  XNOR U24635 ( .A(n24256), .B(n24283), .Z(n24257) );
  XNOR U24636 ( .A(n24282), .B(n25532), .Z(n24283) );
  XNOR U24637 ( .A(n25523), .B(n25531), .Z(n25532) );
  XNOR U24638 ( .A(n25522), .B(n25528), .Z(n25531) );
  XNOR U24639 ( .A(n25527), .B(n24292), .Z(n25528) );
  XNOR U24640 ( .A(n24291), .B(n25521), .Z(n24292) );
  XNOR U24641 ( .A(n25512), .B(n25520), .Z(n25521) );
  XNOR U24642 ( .A(n25511), .B(n25517), .Z(n25520) );
  XNOR U24643 ( .A(n25516), .B(n24301), .Z(n25517) );
  XNOR U24644 ( .A(n24300), .B(n25510), .Z(n24301) );
  XNOR U24645 ( .A(n25501), .B(n25509), .Z(n25510) );
  XNOR U24646 ( .A(n25500), .B(n25506), .Z(n25509) );
  XNOR U24647 ( .A(n25505), .B(n24310), .Z(n25506) );
  XNOR U24648 ( .A(n24309), .B(n25499), .Z(n24310) );
  XNOR U24649 ( .A(n25490), .B(n25498), .Z(n25499) );
  XNOR U24650 ( .A(n25489), .B(n25495), .Z(n25498) );
  XNOR U24651 ( .A(n25494), .B(n24319), .Z(n25495) );
  XNOR U24652 ( .A(n24318), .B(n25488), .Z(n24319) );
  XNOR U24653 ( .A(n25479), .B(n25487), .Z(n25488) );
  XNOR U24654 ( .A(n25478), .B(n25484), .Z(n25487) );
  XNOR U24655 ( .A(n25483), .B(n24328), .Z(n25484) );
  XNOR U24656 ( .A(n24327), .B(n25477), .Z(n24328) );
  XNOR U24657 ( .A(n25468), .B(n25476), .Z(n25477) );
  XNOR U24658 ( .A(n25467), .B(n25473), .Z(n25476) );
  XNOR U24659 ( .A(n25472), .B(n24337), .Z(n25473) );
  XNOR U24660 ( .A(n24336), .B(n25466), .Z(n24337) );
  XNOR U24661 ( .A(n25457), .B(n25465), .Z(n25466) );
  XNOR U24662 ( .A(n25456), .B(n25462), .Z(n25465) );
  XNOR U24663 ( .A(n25461), .B(n24346), .Z(n25462) );
  XNOR U24664 ( .A(n24345), .B(n25455), .Z(n24346) );
  XNOR U24665 ( .A(n25446), .B(n25454), .Z(n25455) );
  XNOR U24666 ( .A(n25445), .B(n25451), .Z(n25454) );
  XNOR U24667 ( .A(n25450), .B(n24355), .Z(n25451) );
  XNOR U24668 ( .A(n24354), .B(n25444), .Z(n24355) );
  XNOR U24669 ( .A(n25435), .B(n25443), .Z(n25444) );
  XNOR U24670 ( .A(n25434), .B(n25440), .Z(n25443) );
  XNOR U24671 ( .A(n25439), .B(n24364), .Z(n25440) );
  XNOR U24672 ( .A(n24363), .B(n25433), .Z(n24364) );
  XNOR U24673 ( .A(n25424), .B(n25432), .Z(n25433) );
  XNOR U24674 ( .A(n25423), .B(n25429), .Z(n25432) );
  XNOR U24675 ( .A(n25428), .B(n24373), .Z(n25429) );
  XNOR U24676 ( .A(n24372), .B(n25422), .Z(n24373) );
  XNOR U24677 ( .A(n25413), .B(n25421), .Z(n25422) );
  XNOR U24678 ( .A(n25412), .B(n25418), .Z(n25421) );
  XNOR U24679 ( .A(n25417), .B(n24382), .Z(n25418) );
  XNOR U24680 ( .A(n24381), .B(n25411), .Z(n24382) );
  XNOR U24681 ( .A(n25402), .B(n25410), .Z(n25411) );
  XNOR U24682 ( .A(n25401), .B(n25407), .Z(n25410) );
  XNOR U24683 ( .A(n25406), .B(n24391), .Z(n25407) );
  XNOR U24684 ( .A(n24390), .B(n25400), .Z(n24391) );
  XNOR U24685 ( .A(n25391), .B(n25399), .Z(n25400) );
  XNOR U24686 ( .A(n25390), .B(n25396), .Z(n25399) );
  XNOR U24687 ( .A(n25395), .B(n24400), .Z(n25396) );
  XNOR U24688 ( .A(n24399), .B(n25389), .Z(n24400) );
  XNOR U24689 ( .A(n25380), .B(n25388), .Z(n25389) );
  XNOR U24690 ( .A(n25379), .B(n25385), .Z(n25388) );
  XNOR U24691 ( .A(n25384), .B(n24409), .Z(n25385) );
  XNOR U24692 ( .A(n24408), .B(n25378), .Z(n24409) );
  XNOR U24693 ( .A(n25369), .B(n25377), .Z(n25378) );
  XNOR U24694 ( .A(n25368), .B(n25374), .Z(n25377) );
  XNOR U24695 ( .A(n25373), .B(n24418), .Z(n25374) );
  XNOR U24696 ( .A(n24417), .B(n25367), .Z(n24418) );
  XNOR U24697 ( .A(n25358), .B(n25366), .Z(n25367) );
  XNOR U24698 ( .A(n25357), .B(n25363), .Z(n25366) );
  XNOR U24699 ( .A(n25362), .B(n24427), .Z(n25363) );
  XNOR U24700 ( .A(n24426), .B(n25356), .Z(n24427) );
  XNOR U24701 ( .A(n25347), .B(n25355), .Z(n25356) );
  XNOR U24702 ( .A(n25346), .B(n25352), .Z(n25355) );
  XNOR U24703 ( .A(n25351), .B(n24436), .Z(n25352) );
  XNOR U24704 ( .A(n24435), .B(n25345), .Z(n24436) );
  XNOR U24705 ( .A(n25336), .B(n25344), .Z(n25345) );
  XNOR U24706 ( .A(n25335), .B(n25341), .Z(n25344) );
  XNOR U24707 ( .A(n25340), .B(n24445), .Z(n25341) );
  XNOR U24708 ( .A(n24444), .B(n25334), .Z(n24445) );
  XNOR U24709 ( .A(n25325), .B(n25333), .Z(n25334) );
  XNOR U24710 ( .A(n25324), .B(n25330), .Z(n25333) );
  XNOR U24711 ( .A(n25329), .B(n24454), .Z(n25330) );
  XNOR U24712 ( .A(n24453), .B(n25323), .Z(n24454) );
  XNOR U24713 ( .A(n25314), .B(n25322), .Z(n25323) );
  XNOR U24714 ( .A(n25313), .B(n25319), .Z(n25322) );
  XNOR U24715 ( .A(n25318), .B(n24463), .Z(n25319) );
  XNOR U24716 ( .A(n24462), .B(n25312), .Z(n24463) );
  XNOR U24717 ( .A(n25303), .B(n25311), .Z(n25312) );
  XNOR U24718 ( .A(n25302), .B(n25308), .Z(n25311) );
  XNOR U24719 ( .A(n25307), .B(n24472), .Z(n25308) );
  XNOR U24720 ( .A(n24471), .B(n25301), .Z(n24472) );
  XNOR U24721 ( .A(n25292), .B(n25300), .Z(n25301) );
  XNOR U24722 ( .A(n25291), .B(n25297), .Z(n25300) );
  XNOR U24723 ( .A(n25296), .B(n24481), .Z(n25297) );
  XNOR U24724 ( .A(n24480), .B(n25290), .Z(n24481) );
  XNOR U24725 ( .A(n25281), .B(n25289), .Z(n25290) );
  XNOR U24726 ( .A(n25280), .B(n25286), .Z(n25289) );
  XNOR U24727 ( .A(n25285), .B(n24490), .Z(n25286) );
  XNOR U24728 ( .A(n24489), .B(n25279), .Z(n24490) );
  XNOR U24729 ( .A(n25270), .B(n25278), .Z(n25279) );
  XNOR U24730 ( .A(n25269), .B(n25275), .Z(n25278) );
  XNOR U24731 ( .A(n25274), .B(n24499), .Z(n25275) );
  XNOR U24732 ( .A(n24498), .B(n25268), .Z(n24499) );
  XNOR U24733 ( .A(n25259), .B(n25267), .Z(n25268) );
  XNOR U24734 ( .A(n25258), .B(n25264), .Z(n25267) );
  XNOR U24735 ( .A(n25263), .B(n24508), .Z(n25264) );
  XNOR U24736 ( .A(n24507), .B(n25257), .Z(n24508) );
  XNOR U24737 ( .A(n25248), .B(n25256), .Z(n25257) );
  XNOR U24738 ( .A(n25247), .B(n25253), .Z(n25256) );
  XNOR U24739 ( .A(n25252), .B(n24517), .Z(n25253) );
  XNOR U24740 ( .A(n24516), .B(n25246), .Z(n24517) );
  XNOR U24741 ( .A(n25237), .B(n25245), .Z(n25246) );
  XNOR U24742 ( .A(n25236), .B(n25242), .Z(n25245) );
  XNOR U24743 ( .A(n25241), .B(n24526), .Z(n25242) );
  XNOR U24744 ( .A(n24525), .B(n25235), .Z(n24526) );
  XNOR U24745 ( .A(n25226), .B(n25234), .Z(n25235) );
  XNOR U24746 ( .A(n25225), .B(n25231), .Z(n25234) );
  XNOR U24747 ( .A(n25230), .B(n24535), .Z(n25231) );
  XNOR U24748 ( .A(n24534), .B(n25224), .Z(n24535) );
  XNOR U24749 ( .A(n25215), .B(n25223), .Z(n25224) );
  XNOR U24750 ( .A(n25214), .B(n25220), .Z(n25223) );
  XNOR U24751 ( .A(n25219), .B(n24544), .Z(n25220) );
  XNOR U24752 ( .A(n24543), .B(n25213), .Z(n24544) );
  XNOR U24753 ( .A(n25204), .B(n25212), .Z(n25213) );
  XNOR U24754 ( .A(n25203), .B(n25209), .Z(n25212) );
  XNOR U24755 ( .A(n25208), .B(n24553), .Z(n25209) );
  XNOR U24756 ( .A(n24552), .B(n25202), .Z(n24553) );
  XNOR U24757 ( .A(n25193), .B(n25201), .Z(n25202) );
  XNOR U24758 ( .A(n25192), .B(n25198), .Z(n25201) );
  XNOR U24759 ( .A(n25197), .B(n24562), .Z(n25198) );
  XNOR U24760 ( .A(n24561), .B(n25191), .Z(n24562) );
  XNOR U24761 ( .A(n25182), .B(n25190), .Z(n25191) );
  XNOR U24762 ( .A(n25181), .B(n25187), .Z(n25190) );
  XNOR U24763 ( .A(n25186), .B(n24571), .Z(n25187) );
  XNOR U24764 ( .A(n24570), .B(n25180), .Z(n24571) );
  XNOR U24765 ( .A(n25171), .B(n25179), .Z(n25180) );
  XNOR U24766 ( .A(n25170), .B(n25176), .Z(n25179) );
  XNOR U24767 ( .A(n25175), .B(n24580), .Z(n25176) );
  XNOR U24768 ( .A(n24579), .B(n25169), .Z(n24580) );
  XNOR U24769 ( .A(n25160), .B(n25168), .Z(n25169) );
  XNOR U24770 ( .A(n25159), .B(n25165), .Z(n25168) );
  XNOR U24771 ( .A(n25164), .B(n24589), .Z(n25165) );
  XNOR U24772 ( .A(n24588), .B(n25158), .Z(n24589) );
  XNOR U24773 ( .A(n25149), .B(n25157), .Z(n25158) );
  XNOR U24774 ( .A(n25148), .B(n25154), .Z(n25157) );
  XNOR U24775 ( .A(n25153), .B(n24598), .Z(n25154) );
  XNOR U24776 ( .A(n24597), .B(n25147), .Z(n24598) );
  XNOR U24777 ( .A(n25138), .B(n25146), .Z(n25147) );
  XNOR U24778 ( .A(n25137), .B(n25143), .Z(n25146) );
  XNOR U24779 ( .A(n25142), .B(n24607), .Z(n25143) );
  XNOR U24780 ( .A(n24606), .B(n25136), .Z(n24607) );
  XNOR U24781 ( .A(n25127), .B(n25135), .Z(n25136) );
  XNOR U24782 ( .A(n25126), .B(n25132), .Z(n25135) );
  XNOR U24783 ( .A(n25131), .B(n24616), .Z(n25132) );
  XNOR U24784 ( .A(n24615), .B(n25125), .Z(n24616) );
  XNOR U24785 ( .A(n25116), .B(n25124), .Z(n25125) );
  XNOR U24786 ( .A(n25115), .B(n25121), .Z(n25124) );
  XNOR U24787 ( .A(n25120), .B(n24625), .Z(n25121) );
  XNOR U24788 ( .A(n24624), .B(n25114), .Z(n24625) );
  XNOR U24789 ( .A(n25105), .B(n25113), .Z(n25114) );
  XNOR U24790 ( .A(n25104), .B(n25110), .Z(n25113) );
  XNOR U24791 ( .A(n25109), .B(n24634), .Z(n25110) );
  XNOR U24792 ( .A(n24633), .B(n25103), .Z(n24634) );
  XNOR U24793 ( .A(n25094), .B(n25102), .Z(n25103) );
  XNOR U24794 ( .A(n25093), .B(n25099), .Z(n25102) );
  XNOR U24795 ( .A(n25098), .B(n24643), .Z(n25099) );
  XNOR U24796 ( .A(n24642), .B(n25092), .Z(n24643) );
  XNOR U24797 ( .A(n25083), .B(n25091), .Z(n25092) );
  XNOR U24798 ( .A(n25082), .B(n25088), .Z(n25091) );
  XNOR U24799 ( .A(n25087), .B(n24652), .Z(n25088) );
  XNOR U24800 ( .A(n24651), .B(n25081), .Z(n24652) );
  XNOR U24801 ( .A(n25072), .B(n25080), .Z(n25081) );
  XNOR U24802 ( .A(n25071), .B(n25077), .Z(n25080) );
  XNOR U24803 ( .A(n25076), .B(n24661), .Z(n25077) );
  XNOR U24804 ( .A(n24660), .B(n25070), .Z(n24661) );
  XNOR U24805 ( .A(n25061), .B(n25069), .Z(n25070) );
  XNOR U24806 ( .A(n25060), .B(n25066), .Z(n25069) );
  XNOR U24807 ( .A(n25065), .B(n24670), .Z(n25066) );
  XNOR U24808 ( .A(n24669), .B(n25059), .Z(n24670) );
  XNOR U24809 ( .A(n25050), .B(n25058), .Z(n25059) );
  XNOR U24810 ( .A(n25049), .B(n25055), .Z(n25058) );
  XNOR U24811 ( .A(n25054), .B(n24679), .Z(n25055) );
  XNOR U24812 ( .A(n24678), .B(n25048), .Z(n24679) );
  XNOR U24813 ( .A(n25039), .B(n25047), .Z(n25048) );
  XNOR U24814 ( .A(n25038), .B(n25044), .Z(n25047) );
  XNOR U24815 ( .A(n25043), .B(n24688), .Z(n25044) );
  XNOR U24816 ( .A(n24687), .B(n25037), .Z(n24688) );
  XNOR U24817 ( .A(n25028), .B(n25036), .Z(n25037) );
  XNOR U24818 ( .A(n25027), .B(n25033), .Z(n25036) );
  XNOR U24819 ( .A(n25032), .B(n24697), .Z(n25033) );
  XNOR U24820 ( .A(n24696), .B(n25026), .Z(n24697) );
  XNOR U24821 ( .A(n25017), .B(n25025), .Z(n25026) );
  XNOR U24822 ( .A(n25016), .B(n25022), .Z(n25025) );
  XNOR U24823 ( .A(n25021), .B(n24706), .Z(n25022) );
  XNOR U24824 ( .A(n24705), .B(n25015), .Z(n24706) );
  XNOR U24825 ( .A(n25006), .B(n25014), .Z(n25015) );
  XNOR U24826 ( .A(n25005), .B(n25011), .Z(n25014) );
  XNOR U24827 ( .A(n25010), .B(n24715), .Z(n25011) );
  XNOR U24828 ( .A(n24714), .B(n25004), .Z(n24715) );
  XNOR U24829 ( .A(n24995), .B(n25003), .Z(n25004) );
  XNOR U24830 ( .A(n24994), .B(n25000), .Z(n25003) );
  XNOR U24831 ( .A(n24999), .B(n24724), .Z(n25000) );
  XNOR U24832 ( .A(n24723), .B(n24993), .Z(n24724) );
  XNOR U24833 ( .A(n24984), .B(n24992), .Z(n24993) );
  XNOR U24834 ( .A(n24983), .B(n24989), .Z(n24992) );
  XNOR U24835 ( .A(n24988), .B(n24733), .Z(n24989) );
  XNOR U24836 ( .A(n24732), .B(n24982), .Z(n24733) );
  XNOR U24837 ( .A(n24973), .B(n24981), .Z(n24982) );
  XNOR U24838 ( .A(n24972), .B(n24978), .Z(n24981) );
  XNOR U24839 ( .A(n24977), .B(n24742), .Z(n24978) );
  XNOR U24840 ( .A(n24741), .B(n24971), .Z(n24742) );
  XNOR U24841 ( .A(n24962), .B(n24970), .Z(n24971) );
  XNOR U24842 ( .A(n24961), .B(n24967), .Z(n24970) );
  XNOR U24843 ( .A(n24966), .B(n24751), .Z(n24967) );
  XNOR U24844 ( .A(n24750), .B(n24960), .Z(n24751) );
  XNOR U24845 ( .A(n24951), .B(n24959), .Z(n24960) );
  XNOR U24846 ( .A(n24950), .B(n24956), .Z(n24959) );
  XNOR U24847 ( .A(n24955), .B(n24760), .Z(n24956) );
  XNOR U24848 ( .A(n24759), .B(n24949), .Z(n24760) );
  XNOR U24849 ( .A(n24940), .B(n24948), .Z(n24949) );
  XNOR U24850 ( .A(n24939), .B(n24945), .Z(n24948) );
  XNOR U24851 ( .A(n24944), .B(n24769), .Z(n24945) );
  XNOR U24852 ( .A(n24768), .B(n24938), .Z(n24769) );
  XNOR U24853 ( .A(n24929), .B(n24937), .Z(n24938) );
  XNOR U24854 ( .A(n24928), .B(n24934), .Z(n24937) );
  XNOR U24855 ( .A(n24933), .B(n24778), .Z(n24934) );
  XNOR U24856 ( .A(n24777), .B(n24927), .Z(n24778) );
  XNOR U24857 ( .A(n24918), .B(n24926), .Z(n24927) );
  XNOR U24858 ( .A(n24917), .B(n24923), .Z(n24926) );
  XNOR U24859 ( .A(n24922), .B(n24787), .Z(n24923) );
  XNOR U24860 ( .A(n24786), .B(n24916), .Z(n24787) );
  XNOR U24861 ( .A(n24907), .B(n24915), .Z(n24916) );
  XNOR U24862 ( .A(n24906), .B(n24912), .Z(n24915) );
  XNOR U24863 ( .A(n24911), .B(n24796), .Z(n24912) );
  XNOR U24864 ( .A(n24795), .B(n24905), .Z(n24796) );
  XNOR U24865 ( .A(n24896), .B(n24904), .Z(n24905) );
  XNOR U24866 ( .A(n24895), .B(n24901), .Z(n24904) );
  XNOR U24867 ( .A(n24900), .B(n24805), .Z(n24901) );
  XNOR U24868 ( .A(n24804), .B(n24894), .Z(n24805) );
  XNOR U24869 ( .A(n24885), .B(n24893), .Z(n24894) );
  XNOR U24870 ( .A(n24884), .B(n24890), .Z(n24893) );
  XNOR U24871 ( .A(n24889), .B(n24814), .Z(n24890) );
  XNOR U24872 ( .A(n24813), .B(n24883), .Z(n24814) );
  XNOR U24873 ( .A(n24874), .B(n24882), .Z(n24883) );
  XNOR U24874 ( .A(n24873), .B(n24879), .Z(n24882) );
  XNOR U24875 ( .A(n24878), .B(n24861), .Z(n24879) );
  XNOR U24876 ( .A(n24820), .B(n24872), .Z(n24861) );
  XNOR U24877 ( .A(n24863), .B(n24871), .Z(n24872) );
  XNOR U24878 ( .A(n24862), .B(n24868), .Z(n24871) );
  XNOR U24879 ( .A(n24867), .B(n24851), .Z(n24868) );
  XNOR U24880 ( .A(n24823), .B(n24860), .Z(n24851) );
  XNOR U24881 ( .A(n24847), .B(n24857), .Z(n24860) );
  XNOR U24882 ( .A(n24850), .B(n24856), .Z(n24857) );
  XNOR U24883 ( .A(n24819), .B(n24846), .Z(n24856) );
  XNOR U24884 ( .A(n24829), .B(n24845), .Z(n24846) );
  XNOR U24885 ( .A(n24832), .B(n24842), .Z(n24845) );
  XOR U24886 ( .A(n24831), .B(n24839), .Z(n24842) );
  XOR U24887 ( .A(n24840), .B(n24838), .Z(n24839) );
  XNOR U24888 ( .A(n26953), .B(n26954), .Z(n24838) );
  XOR U24889 ( .A(n26955), .B(n26956), .Z(n26954) );
  XNOR U24890 ( .A(n26957), .B(n26958), .Z(n26956) );
  NOR U24891 ( .A(n26959), .B(n26958), .Z(n26957) );
  XOR U24892 ( .A(n26960), .B(n26961), .Z(n26955) );
  NOR U24893 ( .A(n26962), .B(n26963), .Z(n26961) );
  AND U24894 ( .A(n26964), .B(n26965), .Z(n26960) );
  XOR U24895 ( .A(n26966), .B(n26967), .Z(n26953) );
  XOR U24896 ( .A(n26968), .B(n26969), .Z(n26967) );
  XOR U24897 ( .A(n26970), .B(n26971), .Z(n26969) );
  XOR U24898 ( .A(n26972), .B(n26973), .Z(n26971) );
  XNOR U24899 ( .A(n26974), .B(n26975), .Z(n26973) );
  NOR U24900 ( .A(n26976), .B(n26975), .Z(n26974) );
  XOR U24901 ( .A(n26977), .B(n26978), .Z(n26972) );
  XOR U24902 ( .A(n26979), .B(n26980), .Z(n26978) );
  XOR U24903 ( .A(n26981), .B(n26982), .Z(n26980) );
  XNOR U24904 ( .A(n26983), .B(n26984), .Z(n26982) );
  NOR U24905 ( .A(n26985), .B(n26984), .Z(n26983) );
  XOR U24906 ( .A(n26986), .B(n26987), .Z(n26981) );
  XOR U24907 ( .A(n26988), .B(n26989), .Z(n26987) );
  XOR U24908 ( .A(n26990), .B(n26991), .Z(n26989) );
  XNOR U24909 ( .A(n26992), .B(n26993), .Z(n26991) );
  NOR U24910 ( .A(n26994), .B(n26993), .Z(n26992) );
  XOR U24911 ( .A(n26995), .B(n26996), .Z(n26990) );
  XOR U24912 ( .A(n26997), .B(n26998), .Z(n26996) );
  XOR U24913 ( .A(n26999), .B(n27000), .Z(n26998) );
  XNOR U24914 ( .A(n27001), .B(n27002), .Z(n27000) );
  NOR U24915 ( .A(n27003), .B(n27002), .Z(n27001) );
  XOR U24916 ( .A(n27004), .B(n27005), .Z(n26999) );
  XOR U24917 ( .A(n27006), .B(n27007), .Z(n27005) );
  XOR U24918 ( .A(n27008), .B(n27009), .Z(n27007) );
  XNOR U24919 ( .A(n27010), .B(n27011), .Z(n27009) );
  NOR U24920 ( .A(n27012), .B(n27011), .Z(n27010) );
  XOR U24921 ( .A(n27013), .B(n27014), .Z(n27008) );
  XOR U24922 ( .A(n27015), .B(n27016), .Z(n27014) );
  XOR U24923 ( .A(n27017), .B(n27018), .Z(n27016) );
  XNOR U24924 ( .A(n27019), .B(n27020), .Z(n27018) );
  NOR U24925 ( .A(n27021), .B(n27020), .Z(n27019) );
  XOR U24926 ( .A(n27022), .B(n27023), .Z(n27017) );
  XOR U24927 ( .A(n27024), .B(n27025), .Z(n27023) );
  XOR U24928 ( .A(n27026), .B(n27027), .Z(n27025) );
  XNOR U24929 ( .A(n27028), .B(n27029), .Z(n27027) );
  NOR U24930 ( .A(n27030), .B(n27029), .Z(n27028) );
  XOR U24931 ( .A(n27031), .B(n27032), .Z(n27026) );
  XOR U24932 ( .A(n27033), .B(n27034), .Z(n27032) );
  XOR U24933 ( .A(n27035), .B(n27036), .Z(n27034) );
  XNOR U24934 ( .A(n27037), .B(n27038), .Z(n27036) );
  NOR U24935 ( .A(n27039), .B(n27038), .Z(n27037) );
  XOR U24936 ( .A(n27040), .B(n27041), .Z(n27035) );
  XOR U24937 ( .A(n27042), .B(n27043), .Z(n27041) );
  XOR U24938 ( .A(n27044), .B(n27045), .Z(n27043) );
  XNOR U24939 ( .A(n27046), .B(n27047), .Z(n27045) );
  NOR U24940 ( .A(n27048), .B(n27047), .Z(n27046) );
  XOR U24941 ( .A(n27049), .B(n27050), .Z(n27044) );
  XOR U24942 ( .A(n27051), .B(n27052), .Z(n27050) );
  XOR U24943 ( .A(n27053), .B(n27054), .Z(n27052) );
  XNOR U24944 ( .A(n27055), .B(n27056), .Z(n27054) );
  NOR U24945 ( .A(n27057), .B(n27056), .Z(n27055) );
  XOR U24946 ( .A(n27058), .B(n27059), .Z(n27053) );
  XOR U24947 ( .A(n27060), .B(n27061), .Z(n27059) );
  XOR U24948 ( .A(n27062), .B(n27063), .Z(n27061) );
  XNOR U24949 ( .A(n27064), .B(n27065), .Z(n27063) );
  NOR U24950 ( .A(n27066), .B(n27065), .Z(n27064) );
  XOR U24951 ( .A(n27067), .B(n27068), .Z(n27062) );
  XOR U24952 ( .A(n27069), .B(n27070), .Z(n27068) );
  XOR U24953 ( .A(n27071), .B(n27072), .Z(n27070) );
  XNOR U24954 ( .A(n27073), .B(n27074), .Z(n27072) );
  NOR U24955 ( .A(n27075), .B(n27074), .Z(n27073) );
  XOR U24956 ( .A(n27076), .B(n27077), .Z(n27071) );
  XOR U24957 ( .A(n27078), .B(n27079), .Z(n27077) );
  XOR U24958 ( .A(n27080), .B(n27081), .Z(n27079) );
  XNOR U24959 ( .A(n27082), .B(n27083), .Z(n27081) );
  NOR U24960 ( .A(n27084), .B(n27083), .Z(n27082) );
  XOR U24961 ( .A(n27085), .B(n27086), .Z(n27080) );
  XOR U24962 ( .A(n27087), .B(n27088), .Z(n27086) );
  XOR U24963 ( .A(n27089), .B(n27090), .Z(n27088) );
  XNOR U24964 ( .A(n27091), .B(n27092), .Z(n27090) );
  NOR U24965 ( .A(n27093), .B(n27092), .Z(n27091) );
  XOR U24966 ( .A(n27094), .B(n27095), .Z(n27089) );
  XOR U24967 ( .A(n27096), .B(n27097), .Z(n27095) );
  XOR U24968 ( .A(n27098), .B(n27099), .Z(n27097) );
  XNOR U24969 ( .A(n27100), .B(n27101), .Z(n27099) );
  NOR U24970 ( .A(n27102), .B(n27101), .Z(n27100) );
  XOR U24971 ( .A(n27103), .B(n27104), .Z(n27098) );
  XOR U24972 ( .A(n27105), .B(n27106), .Z(n27104) );
  XOR U24973 ( .A(n27107), .B(n27108), .Z(n27106) );
  XNOR U24974 ( .A(n27109), .B(n27110), .Z(n27108) );
  NOR U24975 ( .A(n27111), .B(n27110), .Z(n27109) );
  XOR U24976 ( .A(n27112), .B(n27113), .Z(n27107) );
  XOR U24977 ( .A(n27114), .B(n27115), .Z(n27113) );
  XOR U24978 ( .A(n27116), .B(n27117), .Z(n27115) );
  XNOR U24979 ( .A(n27118), .B(n27119), .Z(n27117) );
  NOR U24980 ( .A(n27120), .B(n27119), .Z(n27118) );
  XOR U24981 ( .A(n27121), .B(n27122), .Z(n27116) );
  XOR U24982 ( .A(n27123), .B(n27124), .Z(n27122) );
  XOR U24983 ( .A(n27125), .B(n27126), .Z(n27124) );
  XNOR U24984 ( .A(n27127), .B(n27128), .Z(n27126) );
  NOR U24985 ( .A(n27129), .B(n27128), .Z(n27127) );
  XOR U24986 ( .A(n27130), .B(n27131), .Z(n27125) );
  XOR U24987 ( .A(n27132), .B(n27133), .Z(n27131) );
  XOR U24988 ( .A(n27134), .B(n27135), .Z(n27133) );
  XNOR U24989 ( .A(n27136), .B(n27137), .Z(n27135) );
  NOR U24990 ( .A(n27138), .B(n27137), .Z(n27136) );
  XOR U24991 ( .A(n27139), .B(n27140), .Z(n27134) );
  XOR U24992 ( .A(n27141), .B(n27142), .Z(n27140) );
  XOR U24993 ( .A(n27143), .B(n27144), .Z(n27142) );
  XNOR U24994 ( .A(n27145), .B(n27146), .Z(n27144) );
  NOR U24995 ( .A(n27147), .B(n27146), .Z(n27145) );
  XOR U24996 ( .A(n27148), .B(n27149), .Z(n27143) );
  XOR U24997 ( .A(n27150), .B(n27151), .Z(n27149) );
  XOR U24998 ( .A(n27152), .B(n27153), .Z(n27151) );
  XNOR U24999 ( .A(n27154), .B(n27155), .Z(n27153) );
  NOR U25000 ( .A(n27156), .B(n27155), .Z(n27154) );
  XOR U25001 ( .A(n27157), .B(n27158), .Z(n27152) );
  XOR U25002 ( .A(n27159), .B(n27160), .Z(n27158) );
  XOR U25003 ( .A(n27161), .B(n27162), .Z(n27160) );
  XNOR U25004 ( .A(n27163), .B(n27164), .Z(n27162) );
  NOR U25005 ( .A(n27165), .B(n27164), .Z(n27163) );
  XOR U25006 ( .A(n27166), .B(n27167), .Z(n27161) );
  XOR U25007 ( .A(n27168), .B(n27169), .Z(n27167) );
  XOR U25008 ( .A(n27170), .B(n27171), .Z(n27169) );
  XNOR U25009 ( .A(n27172), .B(n27173), .Z(n27171) );
  NOR U25010 ( .A(n27174), .B(n27173), .Z(n27172) );
  XOR U25011 ( .A(n27175), .B(n27176), .Z(n27170) );
  XOR U25012 ( .A(n27177), .B(n27178), .Z(n27176) );
  XOR U25013 ( .A(n27179), .B(n27180), .Z(n27178) );
  XNOR U25014 ( .A(n27181), .B(n27182), .Z(n27180) );
  NOR U25015 ( .A(n27183), .B(n27182), .Z(n27181) );
  XOR U25016 ( .A(n27184), .B(n27185), .Z(n27179) );
  XOR U25017 ( .A(n27186), .B(n27187), .Z(n27185) );
  XOR U25018 ( .A(n27188), .B(n27189), .Z(n27187) );
  XNOR U25019 ( .A(n27190), .B(n27191), .Z(n27189) );
  NOR U25020 ( .A(n27192), .B(n27191), .Z(n27190) );
  XOR U25021 ( .A(n27193), .B(n27194), .Z(n27188) );
  XOR U25022 ( .A(n27195), .B(n27196), .Z(n27194) );
  XOR U25023 ( .A(n27197), .B(n27198), .Z(n27196) );
  XNOR U25024 ( .A(n27199), .B(n27200), .Z(n27198) );
  NOR U25025 ( .A(n27201), .B(n27200), .Z(n27199) );
  XOR U25026 ( .A(n27202), .B(n27203), .Z(n27197) );
  XOR U25027 ( .A(n27204), .B(n27205), .Z(n27203) );
  XOR U25028 ( .A(n27206), .B(n27207), .Z(n27205) );
  XNOR U25029 ( .A(n27208), .B(n27209), .Z(n27207) );
  NOR U25030 ( .A(n27210), .B(n27209), .Z(n27208) );
  XOR U25031 ( .A(n27211), .B(n27212), .Z(n27206) );
  XOR U25032 ( .A(n27213), .B(n27214), .Z(n27212) );
  XOR U25033 ( .A(n27215), .B(n27216), .Z(n27214) );
  XNOR U25034 ( .A(n27217), .B(n27218), .Z(n27216) );
  NOR U25035 ( .A(n27219), .B(n27218), .Z(n27217) );
  XOR U25036 ( .A(n27220), .B(n27221), .Z(n27215) );
  XOR U25037 ( .A(n27222), .B(n27223), .Z(n27221) );
  XOR U25038 ( .A(n27224), .B(n27225), .Z(n27223) );
  XNOR U25039 ( .A(n27226), .B(n27227), .Z(n27225) );
  NOR U25040 ( .A(n27228), .B(n27227), .Z(n27226) );
  XOR U25041 ( .A(n27229), .B(n27230), .Z(n27224) );
  XOR U25042 ( .A(n27231), .B(n27232), .Z(n27230) );
  XOR U25043 ( .A(n27233), .B(n27234), .Z(n27232) );
  XOR U25044 ( .A(n27235), .B(n27236), .Z(n27231) );
  XNOR U25045 ( .A(n27237), .B(n27238), .Z(n27236) );
  XOR U25046 ( .A(n27239), .B(n27240), .Z(n27238) );
  XOR U25047 ( .A(n27241), .B(n27242), .Z(n27240) );
  XNOR U25048 ( .A(n27243), .B(n27244), .Z(n27242) );
  XOR U25049 ( .A(n27245), .B(n27246), .Z(n27241) );
  XOR U25050 ( .A(n27247), .B(n27248), .Z(n27239) );
  XOR U25051 ( .A(n27249), .B(n27250), .Z(n27248) );
  AND U25052 ( .A(n27251), .B(n27252), .Z(n27250) );
  XOR U25053 ( .A(n27244), .B(n27253), .Z(n27251) );
  XOR U25054 ( .A(n27254), .B(n27255), .Z(n27244) );
  AND U25055 ( .A(n27253), .B(n27254), .Z(n27255) );
  NOR U25056 ( .A(n27256), .B(n27245), .Z(n27249) );
  XOR U25057 ( .A(n27257), .B(n27258), .Z(n27247) );
  NOR U25058 ( .A(n27259), .B(n27246), .Z(n27258) );
  NOR U25059 ( .A(n27260), .B(n27243), .Z(n27257) );
  XNOR U25060 ( .A(n27261), .B(n27262), .Z(n27235) );
  XNOR U25061 ( .A(n27263), .B(n27264), .Z(n27262) );
  NOR U25062 ( .A(n27265), .B(n27237), .Z(n27263) );
  XOR U25063 ( .A(n27266), .B(n27267), .Z(n27229) );
  XOR U25064 ( .A(n27268), .B(n27269), .Z(n27267) );
  NOR U25065 ( .A(n27270), .B(n27233), .Z(n27269) );
  NOR U25066 ( .A(n27271), .B(n27264), .Z(n27268) );
  XOR U25067 ( .A(n27272), .B(n27273), .Z(n27266) );
  NOR U25068 ( .A(n27274), .B(n27261), .Z(n27273) );
  NOR U25069 ( .A(n27275), .B(n27234), .Z(n27272) );
  XOR U25070 ( .A(n27276), .B(n27277), .Z(n27222) );
  XOR U25071 ( .A(n27278), .B(n27279), .Z(n27220) );
  XNOR U25072 ( .A(n27280), .B(n27281), .Z(n27279) );
  NOR U25073 ( .A(n27282), .B(n27281), .Z(n27280) );
  XOR U25074 ( .A(n27283), .B(n27284), .Z(n27278) );
  NOR U25075 ( .A(n27285), .B(n27276), .Z(n27284) );
  NOR U25076 ( .A(n27286), .B(n27277), .Z(n27283) );
  XOR U25077 ( .A(n27287), .B(n27288), .Z(n27213) );
  XOR U25078 ( .A(n27289), .B(n27290), .Z(n27211) );
  XNOR U25079 ( .A(n27291), .B(n27292), .Z(n27290) );
  NOR U25080 ( .A(n27293), .B(n27292), .Z(n27291) );
  XOR U25081 ( .A(n27294), .B(n27295), .Z(n27289) );
  NOR U25082 ( .A(n27296), .B(n27287), .Z(n27295) );
  NOR U25083 ( .A(n27297), .B(n27288), .Z(n27294) );
  XOR U25084 ( .A(n27298), .B(n27299), .Z(n27204) );
  XOR U25085 ( .A(n27300), .B(n27301), .Z(n27202) );
  XNOR U25086 ( .A(n27302), .B(n27303), .Z(n27301) );
  NOR U25087 ( .A(n27304), .B(n27303), .Z(n27302) );
  XOR U25088 ( .A(n27305), .B(n27306), .Z(n27300) );
  NOR U25089 ( .A(n27307), .B(n27298), .Z(n27306) );
  NOR U25090 ( .A(n27308), .B(n27299), .Z(n27305) );
  XOR U25091 ( .A(n27309), .B(n27310), .Z(n27195) );
  XOR U25092 ( .A(n27311), .B(n27312), .Z(n27193) );
  XNOR U25093 ( .A(n27313), .B(n27314), .Z(n27312) );
  NOR U25094 ( .A(n27315), .B(n27314), .Z(n27313) );
  XOR U25095 ( .A(n27316), .B(n27317), .Z(n27311) );
  NOR U25096 ( .A(n27318), .B(n27309), .Z(n27317) );
  NOR U25097 ( .A(n27319), .B(n27310), .Z(n27316) );
  XOR U25098 ( .A(n27320), .B(n27321), .Z(n27186) );
  XOR U25099 ( .A(n27322), .B(n27323), .Z(n27184) );
  XNOR U25100 ( .A(n27324), .B(n27325), .Z(n27323) );
  NOR U25101 ( .A(n27326), .B(n27325), .Z(n27324) );
  XOR U25102 ( .A(n27327), .B(n27328), .Z(n27322) );
  NOR U25103 ( .A(n27329), .B(n27320), .Z(n27328) );
  NOR U25104 ( .A(n27330), .B(n27321), .Z(n27327) );
  XOR U25105 ( .A(n27331), .B(n27332), .Z(n27177) );
  XOR U25106 ( .A(n27333), .B(n27334), .Z(n27175) );
  XNOR U25107 ( .A(n27335), .B(n27336), .Z(n27334) );
  NOR U25108 ( .A(n27337), .B(n27336), .Z(n27335) );
  XOR U25109 ( .A(n27338), .B(n27339), .Z(n27333) );
  NOR U25110 ( .A(n27340), .B(n27331), .Z(n27339) );
  NOR U25111 ( .A(n27341), .B(n27332), .Z(n27338) );
  XOR U25112 ( .A(n27342), .B(n27343), .Z(n27168) );
  XOR U25113 ( .A(n27344), .B(n27345), .Z(n27166) );
  XNOR U25114 ( .A(n27346), .B(n27347), .Z(n27345) );
  NOR U25115 ( .A(n27348), .B(n27347), .Z(n27346) );
  XOR U25116 ( .A(n27349), .B(n27350), .Z(n27344) );
  NOR U25117 ( .A(n27351), .B(n27342), .Z(n27350) );
  NOR U25118 ( .A(n27352), .B(n27343), .Z(n27349) );
  XOR U25119 ( .A(n27353), .B(n27354), .Z(n27159) );
  XOR U25120 ( .A(n27355), .B(n27356), .Z(n27157) );
  XNOR U25121 ( .A(n27357), .B(n27358), .Z(n27356) );
  NOR U25122 ( .A(n27359), .B(n27358), .Z(n27357) );
  XOR U25123 ( .A(n27360), .B(n27361), .Z(n27355) );
  NOR U25124 ( .A(n27362), .B(n27353), .Z(n27361) );
  NOR U25125 ( .A(n27363), .B(n27354), .Z(n27360) );
  XOR U25126 ( .A(n27364), .B(n27365), .Z(n27150) );
  XOR U25127 ( .A(n27366), .B(n27367), .Z(n27148) );
  XNOR U25128 ( .A(n27368), .B(n27369), .Z(n27367) );
  NOR U25129 ( .A(n27370), .B(n27369), .Z(n27368) );
  XOR U25130 ( .A(n27371), .B(n27372), .Z(n27366) );
  NOR U25131 ( .A(n27373), .B(n27364), .Z(n27372) );
  NOR U25132 ( .A(n27374), .B(n27365), .Z(n27371) );
  XOR U25133 ( .A(n27375), .B(n27376), .Z(n27141) );
  XOR U25134 ( .A(n27377), .B(n27378), .Z(n27139) );
  XNOR U25135 ( .A(n27379), .B(n27380), .Z(n27378) );
  NOR U25136 ( .A(n27381), .B(n27380), .Z(n27379) );
  XOR U25137 ( .A(n27382), .B(n27383), .Z(n27377) );
  NOR U25138 ( .A(n27384), .B(n27375), .Z(n27383) );
  NOR U25139 ( .A(n27385), .B(n27376), .Z(n27382) );
  XOR U25140 ( .A(n27386), .B(n27387), .Z(n27132) );
  XOR U25141 ( .A(n27388), .B(n27389), .Z(n27130) );
  XNOR U25142 ( .A(n27390), .B(n27391), .Z(n27389) );
  NOR U25143 ( .A(n27392), .B(n27391), .Z(n27390) );
  XOR U25144 ( .A(n27393), .B(n27394), .Z(n27388) );
  NOR U25145 ( .A(n27395), .B(n27386), .Z(n27394) );
  NOR U25146 ( .A(n27396), .B(n27387), .Z(n27393) );
  XOR U25147 ( .A(n27397), .B(n27398), .Z(n27123) );
  XOR U25148 ( .A(n27399), .B(n27400), .Z(n27121) );
  XNOR U25149 ( .A(n27401), .B(n27402), .Z(n27400) );
  NOR U25150 ( .A(n27403), .B(n27402), .Z(n27401) );
  XOR U25151 ( .A(n27404), .B(n27405), .Z(n27399) );
  NOR U25152 ( .A(n27406), .B(n27397), .Z(n27405) );
  NOR U25153 ( .A(n27407), .B(n27398), .Z(n27404) );
  XOR U25154 ( .A(n27408), .B(n27409), .Z(n27114) );
  XOR U25155 ( .A(n27410), .B(n27411), .Z(n27112) );
  XNOR U25156 ( .A(n27412), .B(n27413), .Z(n27411) );
  NOR U25157 ( .A(n27414), .B(n27413), .Z(n27412) );
  XOR U25158 ( .A(n27415), .B(n27416), .Z(n27410) );
  NOR U25159 ( .A(n27417), .B(n27408), .Z(n27416) );
  NOR U25160 ( .A(n27418), .B(n27409), .Z(n27415) );
  XOR U25161 ( .A(n27419), .B(n27420), .Z(n27105) );
  XOR U25162 ( .A(n27421), .B(n27422), .Z(n27103) );
  XNOR U25163 ( .A(n27423), .B(n27424), .Z(n27422) );
  NOR U25164 ( .A(n27425), .B(n27424), .Z(n27423) );
  XOR U25165 ( .A(n27426), .B(n27427), .Z(n27421) );
  NOR U25166 ( .A(n27428), .B(n27419), .Z(n27427) );
  NOR U25167 ( .A(n27429), .B(n27420), .Z(n27426) );
  XOR U25168 ( .A(n27430), .B(n27431), .Z(n27096) );
  XOR U25169 ( .A(n27432), .B(n27433), .Z(n27094) );
  XNOR U25170 ( .A(n27434), .B(n27435), .Z(n27433) );
  NOR U25171 ( .A(n27436), .B(n27435), .Z(n27434) );
  XOR U25172 ( .A(n27437), .B(n27438), .Z(n27432) );
  NOR U25173 ( .A(n27439), .B(n27430), .Z(n27438) );
  NOR U25174 ( .A(n27440), .B(n27431), .Z(n27437) );
  XOR U25175 ( .A(n27441), .B(n27442), .Z(n27087) );
  XOR U25176 ( .A(n27443), .B(n27444), .Z(n27085) );
  XNOR U25177 ( .A(n27445), .B(n27446), .Z(n27444) );
  NOR U25178 ( .A(n27447), .B(n27446), .Z(n27445) );
  XOR U25179 ( .A(n27448), .B(n27449), .Z(n27443) );
  NOR U25180 ( .A(n27450), .B(n27441), .Z(n27449) );
  NOR U25181 ( .A(n27451), .B(n27442), .Z(n27448) );
  XOR U25182 ( .A(n27452), .B(n27453), .Z(n27078) );
  XOR U25183 ( .A(n27454), .B(n27455), .Z(n27076) );
  XNOR U25184 ( .A(n27456), .B(n27457), .Z(n27455) );
  NOR U25185 ( .A(n27458), .B(n27457), .Z(n27456) );
  XOR U25186 ( .A(n27459), .B(n27460), .Z(n27454) );
  NOR U25187 ( .A(n27461), .B(n27452), .Z(n27460) );
  NOR U25188 ( .A(n27462), .B(n27453), .Z(n27459) );
  XOR U25189 ( .A(n27463), .B(n27464), .Z(n27069) );
  XOR U25190 ( .A(n27465), .B(n27466), .Z(n27067) );
  XNOR U25191 ( .A(n27467), .B(n27468), .Z(n27466) );
  NOR U25192 ( .A(n27469), .B(n27468), .Z(n27467) );
  XOR U25193 ( .A(n27470), .B(n27471), .Z(n27465) );
  NOR U25194 ( .A(n27472), .B(n27463), .Z(n27471) );
  NOR U25195 ( .A(n27473), .B(n27464), .Z(n27470) );
  XOR U25196 ( .A(n27474), .B(n27475), .Z(n27060) );
  XOR U25197 ( .A(n27476), .B(n27477), .Z(n27058) );
  XNOR U25198 ( .A(n27478), .B(n27479), .Z(n27477) );
  NOR U25199 ( .A(n27480), .B(n27479), .Z(n27478) );
  XOR U25200 ( .A(n27481), .B(n27482), .Z(n27476) );
  NOR U25201 ( .A(n27483), .B(n27474), .Z(n27482) );
  NOR U25202 ( .A(n27484), .B(n27475), .Z(n27481) );
  XOR U25203 ( .A(n27485), .B(n27486), .Z(n27051) );
  XOR U25204 ( .A(n27487), .B(n27488), .Z(n27049) );
  XNOR U25205 ( .A(n27489), .B(n27490), .Z(n27488) );
  NOR U25206 ( .A(n27491), .B(n27490), .Z(n27489) );
  XOR U25207 ( .A(n27492), .B(n27493), .Z(n27487) );
  NOR U25208 ( .A(n27494), .B(n27485), .Z(n27493) );
  NOR U25209 ( .A(n27495), .B(n27486), .Z(n27492) );
  XOR U25210 ( .A(n27496), .B(n27497), .Z(n27042) );
  XOR U25211 ( .A(n27498), .B(n27499), .Z(n27040) );
  XNOR U25212 ( .A(n27500), .B(n27501), .Z(n27499) );
  NOR U25213 ( .A(n27502), .B(n27501), .Z(n27500) );
  XOR U25214 ( .A(n27503), .B(n27504), .Z(n27498) );
  NOR U25215 ( .A(n27505), .B(n27496), .Z(n27504) );
  NOR U25216 ( .A(n27506), .B(n27497), .Z(n27503) );
  XOR U25217 ( .A(n27507), .B(n27508), .Z(n27033) );
  XOR U25218 ( .A(n27509), .B(n27510), .Z(n27031) );
  XNOR U25219 ( .A(n27511), .B(n27512), .Z(n27510) );
  NOR U25220 ( .A(n27513), .B(n27512), .Z(n27511) );
  XOR U25221 ( .A(n27514), .B(n27515), .Z(n27509) );
  NOR U25222 ( .A(n27516), .B(n27507), .Z(n27515) );
  NOR U25223 ( .A(n27517), .B(n27508), .Z(n27514) );
  XOR U25224 ( .A(n27518), .B(n27519), .Z(n27024) );
  XOR U25225 ( .A(n27520), .B(n27521), .Z(n27022) );
  XNOR U25226 ( .A(n27522), .B(n27523), .Z(n27521) );
  NOR U25227 ( .A(n27524), .B(n27523), .Z(n27522) );
  XOR U25228 ( .A(n27525), .B(n27526), .Z(n27520) );
  NOR U25229 ( .A(n27527), .B(n27518), .Z(n27526) );
  NOR U25230 ( .A(n27528), .B(n27519), .Z(n27525) );
  XOR U25231 ( .A(n27529), .B(n27530), .Z(n27015) );
  XOR U25232 ( .A(n27531), .B(n27532), .Z(n27013) );
  XNOR U25233 ( .A(n27533), .B(n27534), .Z(n27532) );
  NOR U25234 ( .A(n27535), .B(n27534), .Z(n27533) );
  XOR U25235 ( .A(n27536), .B(n27537), .Z(n27531) );
  NOR U25236 ( .A(n27538), .B(n27529), .Z(n27537) );
  NOR U25237 ( .A(n27539), .B(n27530), .Z(n27536) );
  XOR U25238 ( .A(n27540), .B(n27541), .Z(n27006) );
  XOR U25239 ( .A(n27542), .B(n27543), .Z(n27004) );
  XNOR U25240 ( .A(n27544), .B(n27545), .Z(n27543) );
  NOR U25241 ( .A(n27546), .B(n27545), .Z(n27544) );
  XOR U25242 ( .A(n27547), .B(n27548), .Z(n27542) );
  NOR U25243 ( .A(n27549), .B(n27540), .Z(n27548) );
  NOR U25244 ( .A(n27550), .B(n27541), .Z(n27547) );
  XOR U25245 ( .A(n27551), .B(n27552), .Z(n26997) );
  XOR U25246 ( .A(n27553), .B(n27554), .Z(n26995) );
  XNOR U25247 ( .A(n27555), .B(n27556), .Z(n27554) );
  NOR U25248 ( .A(n27557), .B(n27556), .Z(n27555) );
  XOR U25249 ( .A(n27558), .B(n27559), .Z(n27553) );
  NOR U25250 ( .A(n27560), .B(n27551), .Z(n27559) );
  NOR U25251 ( .A(n27561), .B(n27552), .Z(n27558) );
  XOR U25252 ( .A(n27562), .B(n27563), .Z(n26988) );
  XOR U25253 ( .A(n27564), .B(n27565), .Z(n26986) );
  XNOR U25254 ( .A(n27566), .B(n27567), .Z(n27565) );
  NOR U25255 ( .A(n27568), .B(n27567), .Z(n27566) );
  XOR U25256 ( .A(n27569), .B(n27570), .Z(n27564) );
  NOR U25257 ( .A(n27571), .B(n27562), .Z(n27570) );
  NOR U25258 ( .A(n27572), .B(n27563), .Z(n27569) );
  XOR U25259 ( .A(n27573), .B(n27574), .Z(n26979) );
  XOR U25260 ( .A(n27575), .B(n27576), .Z(n26977) );
  XNOR U25261 ( .A(n27577), .B(n27578), .Z(n27576) );
  NOR U25262 ( .A(n27579), .B(n27578), .Z(n27577) );
  XOR U25263 ( .A(n27580), .B(n27581), .Z(n27575) );
  NOR U25264 ( .A(n27582), .B(n27573), .Z(n27581) );
  NOR U25265 ( .A(n27583), .B(n27574), .Z(n27580) );
  XOR U25266 ( .A(n27584), .B(n27585), .Z(n26970) );
  XOR U25267 ( .A(n27586), .B(n27587), .Z(n26968) );
  XNOR U25268 ( .A(n27588), .B(n27589), .Z(n27587) );
  NOR U25269 ( .A(n27590), .B(n27589), .Z(n27588) );
  XOR U25270 ( .A(n27591), .B(n27592), .Z(n27586) );
  NOR U25271 ( .A(n27593), .B(n27584), .Z(n27592) );
  NOR U25272 ( .A(n27594), .B(n27585), .Z(n27591) );
  XOR U25273 ( .A(n26965), .B(n26963), .Z(n26966) );
  XNOR U25274 ( .A(n27595), .B(n27596), .Z(n24840) );
  NOR U25275 ( .A(n27597), .B(n27595), .Z(n27596) );
  XOR U25276 ( .A(n27598), .B(n27599), .Z(n24831) );
  NOR U25277 ( .A(n27600), .B(n27598), .Z(n27599) );
  XOR U25278 ( .A(n27601), .B(n27602), .Z(n24832) );
  NOR U25279 ( .A(n27603), .B(n27601), .Z(n27602) );
  XOR U25280 ( .A(n27604), .B(n27605), .Z(n24829) );
  NOR U25281 ( .A(n27606), .B(n27604), .Z(n27605) );
  XOR U25282 ( .A(n27607), .B(n27608), .Z(n24819) );
  NOR U25283 ( .A(n27609), .B(n27607), .Z(n27608) );
  XOR U25284 ( .A(n27610), .B(n27611), .Z(n24850) );
  NOR U25285 ( .A(n27612), .B(n27610), .Z(n27611) );
  XOR U25286 ( .A(n27613), .B(n27614), .Z(n24847) );
  NOR U25287 ( .A(n27615), .B(n27613), .Z(n27614) );
  XOR U25288 ( .A(n27616), .B(n27617), .Z(n24823) );
  NOR U25289 ( .A(n27618), .B(n27616), .Z(n27617) );
  XOR U25290 ( .A(n27619), .B(n27620), .Z(n24867) );
  NOR U25291 ( .A(n27621), .B(n27619), .Z(n27620) );
  XOR U25292 ( .A(n27622), .B(n27623), .Z(n24862) );
  NOR U25293 ( .A(n27624), .B(n27622), .Z(n27623) );
  XOR U25294 ( .A(n27625), .B(n27626), .Z(n24863) );
  NOR U25295 ( .A(n27627), .B(n27625), .Z(n27626) );
  XOR U25296 ( .A(n27628), .B(n27629), .Z(n24820) );
  NOR U25297 ( .A(n27630), .B(n27628), .Z(n27629) );
  XOR U25298 ( .A(n27631), .B(n27632), .Z(n24878) );
  NOR U25299 ( .A(n27633), .B(n27631), .Z(n27632) );
  XOR U25300 ( .A(n27634), .B(n27635), .Z(n24873) );
  NOR U25301 ( .A(n27636), .B(n27634), .Z(n27635) );
  XOR U25302 ( .A(n27637), .B(n27638), .Z(n24874) );
  NOR U25303 ( .A(n27639), .B(n27637), .Z(n27638) );
  XOR U25304 ( .A(n27640), .B(n27641), .Z(n24813) );
  NOR U25305 ( .A(n27642), .B(n27640), .Z(n27641) );
  XOR U25306 ( .A(n27643), .B(n27644), .Z(n24889) );
  NOR U25307 ( .A(n27645), .B(n27643), .Z(n27644) );
  XOR U25308 ( .A(n27646), .B(n27647), .Z(n24884) );
  NOR U25309 ( .A(n27648), .B(n27646), .Z(n27647) );
  XOR U25310 ( .A(n27649), .B(n27650), .Z(n24885) );
  NOR U25311 ( .A(n27651), .B(n27649), .Z(n27650) );
  XOR U25312 ( .A(n27652), .B(n27653), .Z(n24804) );
  NOR U25313 ( .A(n27654), .B(n27652), .Z(n27653) );
  XOR U25314 ( .A(n27655), .B(n27656), .Z(n24900) );
  NOR U25315 ( .A(n27657), .B(n27655), .Z(n27656) );
  XOR U25316 ( .A(n27658), .B(n27659), .Z(n24895) );
  NOR U25317 ( .A(n27660), .B(n27658), .Z(n27659) );
  XOR U25318 ( .A(n27661), .B(n27662), .Z(n24896) );
  NOR U25319 ( .A(n27663), .B(n27661), .Z(n27662) );
  XOR U25320 ( .A(n27664), .B(n27665), .Z(n24795) );
  NOR U25321 ( .A(n27666), .B(n27664), .Z(n27665) );
  XOR U25322 ( .A(n27667), .B(n27668), .Z(n24911) );
  NOR U25323 ( .A(n27669), .B(n27667), .Z(n27668) );
  XOR U25324 ( .A(n27670), .B(n27671), .Z(n24906) );
  NOR U25325 ( .A(n27672), .B(n27670), .Z(n27671) );
  XOR U25326 ( .A(n27673), .B(n27674), .Z(n24907) );
  NOR U25327 ( .A(n27675), .B(n27673), .Z(n27674) );
  XOR U25328 ( .A(n27676), .B(n27677), .Z(n24786) );
  NOR U25329 ( .A(n27678), .B(n27676), .Z(n27677) );
  XOR U25330 ( .A(n27679), .B(n27680), .Z(n24922) );
  NOR U25331 ( .A(n27681), .B(n27679), .Z(n27680) );
  XOR U25332 ( .A(n27682), .B(n27683), .Z(n24917) );
  NOR U25333 ( .A(n27684), .B(n27682), .Z(n27683) );
  XOR U25334 ( .A(n27685), .B(n27686), .Z(n24918) );
  NOR U25335 ( .A(n27687), .B(n27685), .Z(n27686) );
  XOR U25336 ( .A(n27688), .B(n27689), .Z(n24777) );
  NOR U25337 ( .A(n27690), .B(n27688), .Z(n27689) );
  XOR U25338 ( .A(n27691), .B(n27692), .Z(n24933) );
  NOR U25339 ( .A(n27693), .B(n27691), .Z(n27692) );
  XOR U25340 ( .A(n27694), .B(n27695), .Z(n24928) );
  NOR U25341 ( .A(n27696), .B(n27694), .Z(n27695) );
  XOR U25342 ( .A(n27697), .B(n27698), .Z(n24929) );
  NOR U25343 ( .A(n27699), .B(n27697), .Z(n27698) );
  XOR U25344 ( .A(n27700), .B(n27701), .Z(n24768) );
  NOR U25345 ( .A(n27702), .B(n27700), .Z(n27701) );
  XOR U25346 ( .A(n27703), .B(n27704), .Z(n24944) );
  NOR U25347 ( .A(n27705), .B(n27703), .Z(n27704) );
  XOR U25348 ( .A(n27706), .B(n27707), .Z(n24939) );
  NOR U25349 ( .A(n27708), .B(n27706), .Z(n27707) );
  XOR U25350 ( .A(n27709), .B(n27710), .Z(n24940) );
  NOR U25351 ( .A(n27711), .B(n27709), .Z(n27710) );
  XOR U25352 ( .A(n27712), .B(n27713), .Z(n24759) );
  NOR U25353 ( .A(n27714), .B(n27712), .Z(n27713) );
  XOR U25354 ( .A(n27715), .B(n27716), .Z(n24955) );
  NOR U25355 ( .A(n27717), .B(n27715), .Z(n27716) );
  XOR U25356 ( .A(n27718), .B(n27719), .Z(n24950) );
  NOR U25357 ( .A(n27720), .B(n27718), .Z(n27719) );
  XOR U25358 ( .A(n27721), .B(n27722), .Z(n24951) );
  NOR U25359 ( .A(n27723), .B(n27721), .Z(n27722) );
  XOR U25360 ( .A(n27724), .B(n27725), .Z(n24750) );
  NOR U25361 ( .A(n27726), .B(n27724), .Z(n27725) );
  XOR U25362 ( .A(n27727), .B(n27728), .Z(n24966) );
  NOR U25363 ( .A(n27729), .B(n27727), .Z(n27728) );
  XOR U25364 ( .A(n27730), .B(n27731), .Z(n24961) );
  NOR U25365 ( .A(n27732), .B(n27730), .Z(n27731) );
  XOR U25366 ( .A(n27733), .B(n27734), .Z(n24962) );
  NOR U25367 ( .A(n27735), .B(n27733), .Z(n27734) );
  XOR U25368 ( .A(n27736), .B(n27737), .Z(n24741) );
  NOR U25369 ( .A(n27738), .B(n27736), .Z(n27737) );
  XOR U25370 ( .A(n27739), .B(n27740), .Z(n24977) );
  NOR U25371 ( .A(n27741), .B(n27739), .Z(n27740) );
  XOR U25372 ( .A(n27742), .B(n27743), .Z(n24972) );
  NOR U25373 ( .A(n27744), .B(n27742), .Z(n27743) );
  XOR U25374 ( .A(n27745), .B(n27746), .Z(n24973) );
  NOR U25375 ( .A(n27747), .B(n27745), .Z(n27746) );
  XOR U25376 ( .A(n27748), .B(n27749), .Z(n24732) );
  NOR U25377 ( .A(n27750), .B(n27748), .Z(n27749) );
  XOR U25378 ( .A(n27751), .B(n27752), .Z(n24988) );
  NOR U25379 ( .A(n27753), .B(n27751), .Z(n27752) );
  XOR U25380 ( .A(n27754), .B(n27755), .Z(n24983) );
  NOR U25381 ( .A(n27756), .B(n27754), .Z(n27755) );
  XOR U25382 ( .A(n27757), .B(n27758), .Z(n24984) );
  NOR U25383 ( .A(n27759), .B(n27757), .Z(n27758) );
  XOR U25384 ( .A(n27760), .B(n27761), .Z(n24723) );
  NOR U25385 ( .A(n27762), .B(n27760), .Z(n27761) );
  XOR U25386 ( .A(n27763), .B(n27764), .Z(n24999) );
  NOR U25387 ( .A(n27765), .B(n27763), .Z(n27764) );
  XOR U25388 ( .A(n27766), .B(n27767), .Z(n24994) );
  NOR U25389 ( .A(n27768), .B(n27766), .Z(n27767) );
  XOR U25390 ( .A(n27769), .B(n27770), .Z(n24995) );
  NOR U25391 ( .A(n27771), .B(n27769), .Z(n27770) );
  XOR U25392 ( .A(n27772), .B(n27773), .Z(n24714) );
  NOR U25393 ( .A(n27774), .B(n27772), .Z(n27773) );
  XOR U25394 ( .A(n27775), .B(n27776), .Z(n25010) );
  NOR U25395 ( .A(n27777), .B(n27775), .Z(n27776) );
  XOR U25396 ( .A(n27778), .B(n27779), .Z(n25005) );
  NOR U25397 ( .A(n27780), .B(n27778), .Z(n27779) );
  XOR U25398 ( .A(n27781), .B(n27782), .Z(n25006) );
  NOR U25399 ( .A(n27783), .B(n27781), .Z(n27782) );
  XOR U25400 ( .A(n27784), .B(n27785), .Z(n24705) );
  NOR U25401 ( .A(n27786), .B(n27784), .Z(n27785) );
  XOR U25402 ( .A(n27787), .B(n27788), .Z(n25021) );
  NOR U25403 ( .A(n27789), .B(n27787), .Z(n27788) );
  XOR U25404 ( .A(n27790), .B(n27791), .Z(n25016) );
  NOR U25405 ( .A(n27792), .B(n27790), .Z(n27791) );
  XOR U25406 ( .A(n27793), .B(n27794), .Z(n25017) );
  NOR U25407 ( .A(n27795), .B(n27793), .Z(n27794) );
  XOR U25408 ( .A(n27796), .B(n27797), .Z(n24696) );
  NOR U25409 ( .A(n27798), .B(n27796), .Z(n27797) );
  XOR U25410 ( .A(n27799), .B(n27800), .Z(n25032) );
  NOR U25411 ( .A(n27801), .B(n27799), .Z(n27800) );
  XOR U25412 ( .A(n27802), .B(n27803), .Z(n25027) );
  NOR U25413 ( .A(n27804), .B(n27802), .Z(n27803) );
  XOR U25414 ( .A(n27805), .B(n27806), .Z(n25028) );
  NOR U25415 ( .A(n27807), .B(n27805), .Z(n27806) );
  XOR U25416 ( .A(n27808), .B(n27809), .Z(n24687) );
  NOR U25417 ( .A(n27810), .B(n27808), .Z(n27809) );
  XOR U25418 ( .A(n27811), .B(n27812), .Z(n25043) );
  NOR U25419 ( .A(n27813), .B(n27811), .Z(n27812) );
  XOR U25420 ( .A(n27814), .B(n27815), .Z(n25038) );
  NOR U25421 ( .A(n27816), .B(n27814), .Z(n27815) );
  XOR U25422 ( .A(n27817), .B(n27818), .Z(n25039) );
  NOR U25423 ( .A(n27819), .B(n27817), .Z(n27818) );
  XOR U25424 ( .A(n27820), .B(n27821), .Z(n24678) );
  NOR U25425 ( .A(n27822), .B(n27820), .Z(n27821) );
  XOR U25426 ( .A(n27823), .B(n27824), .Z(n25054) );
  NOR U25427 ( .A(n27825), .B(n27823), .Z(n27824) );
  XOR U25428 ( .A(n27826), .B(n27827), .Z(n25049) );
  NOR U25429 ( .A(n27828), .B(n27826), .Z(n27827) );
  XOR U25430 ( .A(n27829), .B(n27830), .Z(n25050) );
  NOR U25431 ( .A(n27831), .B(n27829), .Z(n27830) );
  XOR U25432 ( .A(n27832), .B(n27833), .Z(n24669) );
  NOR U25433 ( .A(n27834), .B(n27832), .Z(n27833) );
  XOR U25434 ( .A(n27835), .B(n27836), .Z(n25065) );
  NOR U25435 ( .A(n27837), .B(n27835), .Z(n27836) );
  XOR U25436 ( .A(n27838), .B(n27839), .Z(n25060) );
  NOR U25437 ( .A(n27840), .B(n27838), .Z(n27839) );
  XOR U25438 ( .A(n27841), .B(n27842), .Z(n25061) );
  NOR U25439 ( .A(n27843), .B(n27841), .Z(n27842) );
  XOR U25440 ( .A(n27844), .B(n27845), .Z(n24660) );
  NOR U25441 ( .A(n27846), .B(n27844), .Z(n27845) );
  XOR U25442 ( .A(n27847), .B(n27848), .Z(n25076) );
  NOR U25443 ( .A(n27849), .B(n27847), .Z(n27848) );
  XOR U25444 ( .A(n27850), .B(n27851), .Z(n25071) );
  NOR U25445 ( .A(n27852), .B(n27850), .Z(n27851) );
  XOR U25446 ( .A(n27853), .B(n27854), .Z(n25072) );
  NOR U25447 ( .A(n27855), .B(n27853), .Z(n27854) );
  XOR U25448 ( .A(n27856), .B(n27857), .Z(n24651) );
  NOR U25449 ( .A(n27858), .B(n27856), .Z(n27857) );
  XOR U25450 ( .A(n27859), .B(n27860), .Z(n25087) );
  NOR U25451 ( .A(n27861), .B(n27859), .Z(n27860) );
  XOR U25452 ( .A(n27862), .B(n27863), .Z(n25082) );
  NOR U25453 ( .A(n27864), .B(n27862), .Z(n27863) );
  XOR U25454 ( .A(n27865), .B(n27866), .Z(n25083) );
  NOR U25455 ( .A(n27867), .B(n27865), .Z(n27866) );
  XOR U25456 ( .A(n27868), .B(n27869), .Z(n24642) );
  NOR U25457 ( .A(n27870), .B(n27868), .Z(n27869) );
  XOR U25458 ( .A(n27871), .B(n27872), .Z(n25098) );
  NOR U25459 ( .A(n27873), .B(n27871), .Z(n27872) );
  XOR U25460 ( .A(n27874), .B(n27875), .Z(n25093) );
  NOR U25461 ( .A(n27876), .B(n27874), .Z(n27875) );
  XOR U25462 ( .A(n27877), .B(n27878), .Z(n25094) );
  NOR U25463 ( .A(n27879), .B(n27877), .Z(n27878) );
  XOR U25464 ( .A(n27880), .B(n27881), .Z(n24633) );
  NOR U25465 ( .A(n27882), .B(n27880), .Z(n27881) );
  XOR U25466 ( .A(n27883), .B(n27884), .Z(n25109) );
  NOR U25467 ( .A(n27885), .B(n27883), .Z(n27884) );
  XOR U25468 ( .A(n27886), .B(n27887), .Z(n25104) );
  NOR U25469 ( .A(n27888), .B(n27886), .Z(n27887) );
  XOR U25470 ( .A(n27889), .B(n27890), .Z(n25105) );
  NOR U25471 ( .A(n27891), .B(n27889), .Z(n27890) );
  XOR U25472 ( .A(n27892), .B(n27893), .Z(n24624) );
  NOR U25473 ( .A(n27894), .B(n27892), .Z(n27893) );
  XOR U25474 ( .A(n27895), .B(n27896), .Z(n25120) );
  NOR U25475 ( .A(n27897), .B(n27895), .Z(n27896) );
  XOR U25476 ( .A(n27898), .B(n27899), .Z(n25115) );
  NOR U25477 ( .A(n27900), .B(n27898), .Z(n27899) );
  XOR U25478 ( .A(n27901), .B(n27902), .Z(n25116) );
  NOR U25479 ( .A(n27903), .B(n27901), .Z(n27902) );
  XOR U25480 ( .A(n27904), .B(n27905), .Z(n24615) );
  NOR U25481 ( .A(n27906), .B(n27904), .Z(n27905) );
  XOR U25482 ( .A(n27907), .B(n27908), .Z(n25131) );
  NOR U25483 ( .A(n27909), .B(n27907), .Z(n27908) );
  XOR U25484 ( .A(n27910), .B(n27911), .Z(n25126) );
  NOR U25485 ( .A(n27912), .B(n27910), .Z(n27911) );
  XOR U25486 ( .A(n27913), .B(n27914), .Z(n25127) );
  NOR U25487 ( .A(n27915), .B(n27913), .Z(n27914) );
  XOR U25488 ( .A(n27916), .B(n27917), .Z(n24606) );
  NOR U25489 ( .A(n27918), .B(n27916), .Z(n27917) );
  XOR U25490 ( .A(n27919), .B(n27920), .Z(n25142) );
  NOR U25491 ( .A(n27921), .B(n27919), .Z(n27920) );
  XOR U25492 ( .A(n27922), .B(n27923), .Z(n25137) );
  NOR U25493 ( .A(n27924), .B(n27922), .Z(n27923) );
  XOR U25494 ( .A(n27925), .B(n27926), .Z(n25138) );
  NOR U25495 ( .A(n27927), .B(n27925), .Z(n27926) );
  XOR U25496 ( .A(n27928), .B(n27929), .Z(n24597) );
  NOR U25497 ( .A(n27930), .B(n27928), .Z(n27929) );
  XOR U25498 ( .A(n27931), .B(n27932), .Z(n25153) );
  NOR U25499 ( .A(n27933), .B(n27931), .Z(n27932) );
  XOR U25500 ( .A(n27934), .B(n27935), .Z(n25148) );
  NOR U25501 ( .A(n27936), .B(n27934), .Z(n27935) );
  XOR U25502 ( .A(n27937), .B(n27938), .Z(n25149) );
  NOR U25503 ( .A(n27939), .B(n27937), .Z(n27938) );
  XOR U25504 ( .A(n27940), .B(n27941), .Z(n24588) );
  NOR U25505 ( .A(n27942), .B(n27940), .Z(n27941) );
  XOR U25506 ( .A(n27943), .B(n27944), .Z(n25164) );
  NOR U25507 ( .A(n27945), .B(n27943), .Z(n27944) );
  XOR U25508 ( .A(n27946), .B(n27947), .Z(n25159) );
  NOR U25509 ( .A(n27948), .B(n27946), .Z(n27947) );
  XOR U25510 ( .A(n27949), .B(n27950), .Z(n25160) );
  NOR U25511 ( .A(n27951), .B(n27949), .Z(n27950) );
  XOR U25512 ( .A(n27952), .B(n27953), .Z(n24579) );
  NOR U25513 ( .A(n27954), .B(n27952), .Z(n27953) );
  XOR U25514 ( .A(n27955), .B(n27956), .Z(n25175) );
  NOR U25515 ( .A(n27957), .B(n27955), .Z(n27956) );
  XOR U25516 ( .A(n27958), .B(n27959), .Z(n25170) );
  NOR U25517 ( .A(n27960), .B(n27958), .Z(n27959) );
  XOR U25518 ( .A(n27961), .B(n27962), .Z(n25171) );
  NOR U25519 ( .A(n27963), .B(n27961), .Z(n27962) );
  XOR U25520 ( .A(n27964), .B(n27965), .Z(n24570) );
  NOR U25521 ( .A(n27966), .B(n27964), .Z(n27965) );
  XOR U25522 ( .A(n27967), .B(n27968), .Z(n25186) );
  NOR U25523 ( .A(n27969), .B(n27967), .Z(n27968) );
  XOR U25524 ( .A(n27970), .B(n27971), .Z(n25181) );
  NOR U25525 ( .A(n27972), .B(n27970), .Z(n27971) );
  XOR U25526 ( .A(n27973), .B(n27974), .Z(n25182) );
  NOR U25527 ( .A(n27975), .B(n27973), .Z(n27974) );
  XOR U25528 ( .A(n27976), .B(n27977), .Z(n24561) );
  NOR U25529 ( .A(n27978), .B(n27976), .Z(n27977) );
  XOR U25530 ( .A(n27979), .B(n27980), .Z(n25197) );
  NOR U25531 ( .A(n27981), .B(n27979), .Z(n27980) );
  XOR U25532 ( .A(n27982), .B(n27983), .Z(n25192) );
  NOR U25533 ( .A(n27984), .B(n27982), .Z(n27983) );
  XOR U25534 ( .A(n27985), .B(n27986), .Z(n25193) );
  NOR U25535 ( .A(n27987), .B(n27985), .Z(n27986) );
  XOR U25536 ( .A(n27988), .B(n27989), .Z(n24552) );
  NOR U25537 ( .A(n27990), .B(n27988), .Z(n27989) );
  XOR U25538 ( .A(n27991), .B(n27992), .Z(n25208) );
  NOR U25539 ( .A(n27993), .B(n27991), .Z(n27992) );
  XOR U25540 ( .A(n27994), .B(n27995), .Z(n25203) );
  NOR U25541 ( .A(n27996), .B(n27994), .Z(n27995) );
  XOR U25542 ( .A(n27997), .B(n27998), .Z(n25204) );
  NOR U25543 ( .A(n27999), .B(n27997), .Z(n27998) );
  XOR U25544 ( .A(n28000), .B(n28001), .Z(n24543) );
  NOR U25545 ( .A(n28002), .B(n28000), .Z(n28001) );
  XOR U25546 ( .A(n28003), .B(n28004), .Z(n25219) );
  NOR U25547 ( .A(n28005), .B(n28003), .Z(n28004) );
  XOR U25548 ( .A(n28006), .B(n28007), .Z(n25214) );
  NOR U25549 ( .A(n28008), .B(n28006), .Z(n28007) );
  XOR U25550 ( .A(n28009), .B(n28010), .Z(n25215) );
  NOR U25551 ( .A(n28011), .B(n28009), .Z(n28010) );
  XOR U25552 ( .A(n28012), .B(n28013), .Z(n24534) );
  NOR U25553 ( .A(n28014), .B(n28012), .Z(n28013) );
  XOR U25554 ( .A(n28015), .B(n28016), .Z(n25230) );
  NOR U25555 ( .A(n28017), .B(n28015), .Z(n28016) );
  XOR U25556 ( .A(n28018), .B(n28019), .Z(n25225) );
  NOR U25557 ( .A(n28020), .B(n28018), .Z(n28019) );
  XOR U25558 ( .A(n28021), .B(n28022), .Z(n25226) );
  NOR U25559 ( .A(n28023), .B(n28021), .Z(n28022) );
  XOR U25560 ( .A(n28024), .B(n28025), .Z(n24525) );
  NOR U25561 ( .A(n28026), .B(n28024), .Z(n28025) );
  XOR U25562 ( .A(n28027), .B(n28028), .Z(n25241) );
  NOR U25563 ( .A(n28029), .B(n28027), .Z(n28028) );
  XOR U25564 ( .A(n28030), .B(n28031), .Z(n25236) );
  NOR U25565 ( .A(n28032), .B(n28030), .Z(n28031) );
  XOR U25566 ( .A(n28033), .B(n28034), .Z(n25237) );
  NOR U25567 ( .A(n28035), .B(n28033), .Z(n28034) );
  XOR U25568 ( .A(n28036), .B(n28037), .Z(n24516) );
  NOR U25569 ( .A(n28038), .B(n28036), .Z(n28037) );
  XOR U25570 ( .A(n28039), .B(n28040), .Z(n25252) );
  NOR U25571 ( .A(n28041), .B(n28039), .Z(n28040) );
  XOR U25572 ( .A(n28042), .B(n28043), .Z(n25247) );
  NOR U25573 ( .A(n28044), .B(n28042), .Z(n28043) );
  XOR U25574 ( .A(n28045), .B(n28046), .Z(n25248) );
  NOR U25575 ( .A(n28047), .B(n28045), .Z(n28046) );
  XOR U25576 ( .A(n28048), .B(n28049), .Z(n24507) );
  NOR U25577 ( .A(n28050), .B(n28048), .Z(n28049) );
  XOR U25578 ( .A(n28051), .B(n28052), .Z(n25263) );
  NOR U25579 ( .A(n28053), .B(n28051), .Z(n28052) );
  XOR U25580 ( .A(n28054), .B(n28055), .Z(n25258) );
  NOR U25581 ( .A(n28056), .B(n28054), .Z(n28055) );
  XOR U25582 ( .A(n28057), .B(n28058), .Z(n25259) );
  NOR U25583 ( .A(n28059), .B(n28057), .Z(n28058) );
  XOR U25584 ( .A(n28060), .B(n28061), .Z(n24498) );
  NOR U25585 ( .A(n28062), .B(n28060), .Z(n28061) );
  XOR U25586 ( .A(n28063), .B(n28064), .Z(n25274) );
  NOR U25587 ( .A(n28065), .B(n28063), .Z(n28064) );
  XOR U25588 ( .A(n28066), .B(n28067), .Z(n25269) );
  NOR U25589 ( .A(n28068), .B(n28066), .Z(n28067) );
  XOR U25590 ( .A(n28069), .B(n28070), .Z(n25270) );
  NOR U25591 ( .A(n28071), .B(n28069), .Z(n28070) );
  XOR U25592 ( .A(n28072), .B(n28073), .Z(n24489) );
  NOR U25593 ( .A(n28074), .B(n28072), .Z(n28073) );
  XOR U25594 ( .A(n28075), .B(n28076), .Z(n25285) );
  NOR U25595 ( .A(n28077), .B(n28075), .Z(n28076) );
  XOR U25596 ( .A(n28078), .B(n28079), .Z(n25280) );
  NOR U25597 ( .A(n28080), .B(n28078), .Z(n28079) );
  XOR U25598 ( .A(n28081), .B(n28082), .Z(n25281) );
  NOR U25599 ( .A(n28083), .B(n28081), .Z(n28082) );
  XOR U25600 ( .A(n28084), .B(n28085), .Z(n24480) );
  NOR U25601 ( .A(n28086), .B(n28084), .Z(n28085) );
  XOR U25602 ( .A(n28087), .B(n28088), .Z(n25296) );
  NOR U25603 ( .A(n28089), .B(n28087), .Z(n28088) );
  XOR U25604 ( .A(n28090), .B(n28091), .Z(n25291) );
  NOR U25605 ( .A(n28092), .B(n28090), .Z(n28091) );
  XOR U25606 ( .A(n28093), .B(n28094), .Z(n25292) );
  NOR U25607 ( .A(n28095), .B(n28093), .Z(n28094) );
  XOR U25608 ( .A(n28096), .B(n28097), .Z(n24471) );
  NOR U25609 ( .A(n28098), .B(n28096), .Z(n28097) );
  XOR U25610 ( .A(n28099), .B(n28100), .Z(n25307) );
  NOR U25611 ( .A(n28101), .B(n28099), .Z(n28100) );
  XOR U25612 ( .A(n28102), .B(n28103), .Z(n25302) );
  NOR U25613 ( .A(n28104), .B(n28102), .Z(n28103) );
  XOR U25614 ( .A(n28105), .B(n28106), .Z(n25303) );
  NOR U25615 ( .A(n28107), .B(n28105), .Z(n28106) );
  XOR U25616 ( .A(n28108), .B(n28109), .Z(n24462) );
  NOR U25617 ( .A(n28110), .B(n28108), .Z(n28109) );
  XOR U25618 ( .A(n28111), .B(n28112), .Z(n25318) );
  NOR U25619 ( .A(n28113), .B(n28111), .Z(n28112) );
  XOR U25620 ( .A(n28114), .B(n28115), .Z(n25313) );
  NOR U25621 ( .A(n28116), .B(n28114), .Z(n28115) );
  XOR U25622 ( .A(n28117), .B(n28118), .Z(n25314) );
  NOR U25623 ( .A(n28119), .B(n28117), .Z(n28118) );
  XOR U25624 ( .A(n28120), .B(n28121), .Z(n24453) );
  NOR U25625 ( .A(n28122), .B(n28120), .Z(n28121) );
  XOR U25626 ( .A(n28123), .B(n28124), .Z(n25329) );
  NOR U25627 ( .A(n28125), .B(n28123), .Z(n28124) );
  XOR U25628 ( .A(n28126), .B(n28127), .Z(n25324) );
  NOR U25629 ( .A(n28128), .B(n28126), .Z(n28127) );
  XOR U25630 ( .A(n28129), .B(n28130), .Z(n25325) );
  NOR U25631 ( .A(n28131), .B(n28129), .Z(n28130) );
  XOR U25632 ( .A(n28132), .B(n28133), .Z(n24444) );
  NOR U25633 ( .A(n28134), .B(n28132), .Z(n28133) );
  XOR U25634 ( .A(n28135), .B(n28136), .Z(n25340) );
  NOR U25635 ( .A(n28137), .B(n28135), .Z(n28136) );
  XOR U25636 ( .A(n28138), .B(n28139), .Z(n25335) );
  NOR U25637 ( .A(n28140), .B(n28138), .Z(n28139) );
  XOR U25638 ( .A(n28141), .B(n28142), .Z(n25336) );
  NOR U25639 ( .A(n28143), .B(n28141), .Z(n28142) );
  XOR U25640 ( .A(n28144), .B(n28145), .Z(n24435) );
  NOR U25641 ( .A(n28146), .B(n28144), .Z(n28145) );
  XOR U25642 ( .A(n28147), .B(n28148), .Z(n25351) );
  NOR U25643 ( .A(n28149), .B(n28147), .Z(n28148) );
  XOR U25644 ( .A(n28150), .B(n28151), .Z(n25346) );
  NOR U25645 ( .A(n28152), .B(n28150), .Z(n28151) );
  XOR U25646 ( .A(n28153), .B(n28154), .Z(n25347) );
  NOR U25647 ( .A(n28155), .B(n28153), .Z(n28154) );
  XOR U25648 ( .A(n28156), .B(n28157), .Z(n24426) );
  NOR U25649 ( .A(n28158), .B(n28156), .Z(n28157) );
  XOR U25650 ( .A(n28159), .B(n28160), .Z(n25362) );
  NOR U25651 ( .A(n28161), .B(n28159), .Z(n28160) );
  XOR U25652 ( .A(n28162), .B(n28163), .Z(n25357) );
  NOR U25653 ( .A(n28164), .B(n28162), .Z(n28163) );
  XOR U25654 ( .A(n28165), .B(n28166), .Z(n25358) );
  NOR U25655 ( .A(n28167), .B(n28165), .Z(n28166) );
  XOR U25656 ( .A(n28168), .B(n28169), .Z(n24417) );
  NOR U25657 ( .A(n28170), .B(n28168), .Z(n28169) );
  XOR U25658 ( .A(n28171), .B(n28172), .Z(n25373) );
  NOR U25659 ( .A(n28173), .B(n28171), .Z(n28172) );
  XOR U25660 ( .A(n28174), .B(n28175), .Z(n25368) );
  NOR U25661 ( .A(n28176), .B(n28174), .Z(n28175) );
  XOR U25662 ( .A(n28177), .B(n28178), .Z(n25369) );
  NOR U25663 ( .A(n28179), .B(n28177), .Z(n28178) );
  XOR U25664 ( .A(n28180), .B(n28181), .Z(n24408) );
  NOR U25665 ( .A(n28182), .B(n28180), .Z(n28181) );
  XOR U25666 ( .A(n28183), .B(n28184), .Z(n25384) );
  NOR U25667 ( .A(n28185), .B(n28183), .Z(n28184) );
  XOR U25668 ( .A(n28186), .B(n28187), .Z(n25379) );
  NOR U25669 ( .A(n28188), .B(n28186), .Z(n28187) );
  XOR U25670 ( .A(n28189), .B(n28190), .Z(n25380) );
  NOR U25671 ( .A(n28191), .B(n28189), .Z(n28190) );
  XOR U25672 ( .A(n28192), .B(n28193), .Z(n24399) );
  NOR U25673 ( .A(n28194), .B(n28192), .Z(n28193) );
  XOR U25674 ( .A(n28195), .B(n28196), .Z(n25395) );
  NOR U25675 ( .A(n28197), .B(n28195), .Z(n28196) );
  XOR U25676 ( .A(n28198), .B(n28199), .Z(n25390) );
  NOR U25677 ( .A(n28200), .B(n28198), .Z(n28199) );
  XOR U25678 ( .A(n28201), .B(n28202), .Z(n25391) );
  NOR U25679 ( .A(n28203), .B(n28201), .Z(n28202) );
  XOR U25680 ( .A(n28204), .B(n28205), .Z(n24390) );
  NOR U25681 ( .A(n28206), .B(n28204), .Z(n28205) );
  XOR U25682 ( .A(n28207), .B(n28208), .Z(n25406) );
  NOR U25683 ( .A(n28209), .B(n28207), .Z(n28208) );
  XOR U25684 ( .A(n28210), .B(n28211), .Z(n25401) );
  NOR U25685 ( .A(n28212), .B(n28210), .Z(n28211) );
  XOR U25686 ( .A(n28213), .B(n28214), .Z(n25402) );
  NOR U25687 ( .A(n28215), .B(n28213), .Z(n28214) );
  XOR U25688 ( .A(n28216), .B(n28217), .Z(n24381) );
  NOR U25689 ( .A(n28218), .B(n28216), .Z(n28217) );
  XOR U25690 ( .A(n28219), .B(n28220), .Z(n25417) );
  NOR U25691 ( .A(n28221), .B(n28219), .Z(n28220) );
  XOR U25692 ( .A(n28222), .B(n28223), .Z(n25412) );
  NOR U25693 ( .A(n28224), .B(n28222), .Z(n28223) );
  XOR U25694 ( .A(n28225), .B(n28226), .Z(n25413) );
  NOR U25695 ( .A(n28227), .B(n28225), .Z(n28226) );
  XOR U25696 ( .A(n28228), .B(n28229), .Z(n24372) );
  NOR U25697 ( .A(n28230), .B(n28228), .Z(n28229) );
  XOR U25698 ( .A(n28231), .B(n28232), .Z(n25428) );
  NOR U25699 ( .A(n28233), .B(n28231), .Z(n28232) );
  XOR U25700 ( .A(n28234), .B(n28235), .Z(n25423) );
  NOR U25701 ( .A(n28236), .B(n28234), .Z(n28235) );
  XOR U25702 ( .A(n28237), .B(n28238), .Z(n25424) );
  NOR U25703 ( .A(n28239), .B(n28237), .Z(n28238) );
  XOR U25704 ( .A(n28240), .B(n28241), .Z(n24363) );
  NOR U25705 ( .A(n28242), .B(n28240), .Z(n28241) );
  XOR U25706 ( .A(n28243), .B(n28244), .Z(n25439) );
  NOR U25707 ( .A(n28245), .B(n28243), .Z(n28244) );
  XOR U25708 ( .A(n28246), .B(n28247), .Z(n25434) );
  NOR U25709 ( .A(n28248), .B(n28246), .Z(n28247) );
  XOR U25710 ( .A(n28249), .B(n28250), .Z(n25435) );
  NOR U25711 ( .A(n28251), .B(n28249), .Z(n28250) );
  XOR U25712 ( .A(n28252), .B(n28253), .Z(n24354) );
  NOR U25713 ( .A(n28254), .B(n28252), .Z(n28253) );
  XOR U25714 ( .A(n28255), .B(n28256), .Z(n25450) );
  NOR U25715 ( .A(n28257), .B(n28255), .Z(n28256) );
  XOR U25716 ( .A(n28258), .B(n28259), .Z(n25445) );
  NOR U25717 ( .A(n28260), .B(n28258), .Z(n28259) );
  XOR U25718 ( .A(n28261), .B(n28262), .Z(n25446) );
  NOR U25719 ( .A(n28263), .B(n28261), .Z(n28262) );
  XOR U25720 ( .A(n28264), .B(n28265), .Z(n24345) );
  NOR U25721 ( .A(n28266), .B(n28264), .Z(n28265) );
  XOR U25722 ( .A(n28267), .B(n28268), .Z(n25461) );
  NOR U25723 ( .A(n28269), .B(n28267), .Z(n28268) );
  XOR U25724 ( .A(n28270), .B(n28271), .Z(n25456) );
  NOR U25725 ( .A(n28272), .B(n28270), .Z(n28271) );
  XOR U25726 ( .A(n28273), .B(n28274), .Z(n25457) );
  NOR U25727 ( .A(n28275), .B(n28273), .Z(n28274) );
  XOR U25728 ( .A(n28276), .B(n28277), .Z(n24336) );
  NOR U25729 ( .A(n28278), .B(n28276), .Z(n28277) );
  XOR U25730 ( .A(n28279), .B(n28280), .Z(n25472) );
  NOR U25731 ( .A(n28281), .B(n28279), .Z(n28280) );
  XOR U25732 ( .A(n28282), .B(n28283), .Z(n25467) );
  NOR U25733 ( .A(n28284), .B(n28282), .Z(n28283) );
  XOR U25734 ( .A(n28285), .B(n28286), .Z(n25468) );
  NOR U25735 ( .A(n28287), .B(n28285), .Z(n28286) );
  XOR U25736 ( .A(n28288), .B(n28289), .Z(n24327) );
  NOR U25737 ( .A(n28290), .B(n28288), .Z(n28289) );
  XOR U25738 ( .A(n28291), .B(n28292), .Z(n25483) );
  NOR U25739 ( .A(n28293), .B(n28291), .Z(n28292) );
  XOR U25740 ( .A(n28294), .B(n28295), .Z(n25478) );
  NOR U25741 ( .A(n28296), .B(n28294), .Z(n28295) );
  XOR U25742 ( .A(n28297), .B(n28298), .Z(n25479) );
  NOR U25743 ( .A(n28299), .B(n28297), .Z(n28298) );
  XOR U25744 ( .A(n28300), .B(n28301), .Z(n24318) );
  NOR U25745 ( .A(n28302), .B(n28300), .Z(n28301) );
  XOR U25746 ( .A(n28303), .B(n28304), .Z(n25494) );
  NOR U25747 ( .A(n28305), .B(n28303), .Z(n28304) );
  XOR U25748 ( .A(n28306), .B(n28307), .Z(n25489) );
  NOR U25749 ( .A(n28308), .B(n28306), .Z(n28307) );
  XOR U25750 ( .A(n28309), .B(n28310), .Z(n25490) );
  NOR U25751 ( .A(n28311), .B(n28309), .Z(n28310) );
  XOR U25752 ( .A(n28312), .B(n28313), .Z(n24309) );
  NOR U25753 ( .A(n28314), .B(n28312), .Z(n28313) );
  XOR U25754 ( .A(n28315), .B(n28316), .Z(n25505) );
  NOR U25755 ( .A(n28317), .B(n28315), .Z(n28316) );
  XOR U25756 ( .A(n28318), .B(n28319), .Z(n25500) );
  NOR U25757 ( .A(n28320), .B(n28318), .Z(n28319) );
  XOR U25758 ( .A(n28321), .B(n28322), .Z(n25501) );
  NOR U25759 ( .A(n28323), .B(n28321), .Z(n28322) );
  XOR U25760 ( .A(n28324), .B(n28325), .Z(n24300) );
  NOR U25761 ( .A(n28326), .B(n28324), .Z(n28325) );
  XOR U25762 ( .A(n28327), .B(n28328), .Z(n25516) );
  NOR U25763 ( .A(n28329), .B(n28327), .Z(n28328) );
  XOR U25764 ( .A(n28330), .B(n28331), .Z(n25511) );
  NOR U25765 ( .A(n28332), .B(n28330), .Z(n28331) );
  XOR U25766 ( .A(n28333), .B(n28334), .Z(n25512) );
  NOR U25767 ( .A(n28335), .B(n28333), .Z(n28334) );
  XOR U25768 ( .A(n28336), .B(n28337), .Z(n24291) );
  NOR U25769 ( .A(n28338), .B(n28336), .Z(n28337) );
  XOR U25770 ( .A(n28339), .B(n28340), .Z(n25527) );
  NOR U25771 ( .A(n28341), .B(n28339), .Z(n28340) );
  XOR U25772 ( .A(n28342), .B(n28343), .Z(n25522) );
  NOR U25773 ( .A(n28344), .B(n28342), .Z(n28343) );
  XOR U25774 ( .A(n28345), .B(n28346), .Z(n25523) );
  NOR U25775 ( .A(n28347), .B(n28345), .Z(n28346) );
  XOR U25776 ( .A(n28348), .B(n28349), .Z(n24282) );
  NOR U25777 ( .A(n28350), .B(n28348), .Z(n28349) );
  XNOR U25778 ( .A(n28351), .B(n28352), .Z(n24256) );
  NOR U25779 ( .A(n28353), .B(n28351), .Z(n28352) );
  XNOR U25780 ( .A(n28354), .B(n28355), .Z(n24261) );
  NOR U25781 ( .A(n28356), .B(n28354), .Z(n28355) );
  XOR U25782 ( .A(n28357), .B(n28358), .Z(n24263) );
  NOR U25783 ( .A(n28359), .B(n28357), .Z(n28358) );
  IV U25784 ( .A(n24273), .Z(n26952) );
  XOR U25785 ( .A(n28360), .B(n28361), .Z(n24273) );
  AND U25786 ( .A(n28362), .B(n28360), .Z(n28361) );
  XOR U25787 ( .A(n28363), .B(n28364), .Z(n25533) );
  AND U25788 ( .A(n63), .B(n28363), .Z(n28364) );
  XOR U25789 ( .A(n28365), .B(n28366), .Z(n25535) );
  AND U25790 ( .A(n28367), .B(n28368), .Z(n28366) );
  XOR U25791 ( .A(n28365), .B(n65), .Z(n28368) );
  XOR U25792 ( .A(n26950), .B(n26949), .Z(n65) );
  XNOR U25793 ( .A(n26947), .B(n26946), .Z(n26949) );
  XNOR U25794 ( .A(n26944), .B(n26943), .Z(n26946) );
  XNOR U25795 ( .A(n26941), .B(n26940), .Z(n26943) );
  XNOR U25796 ( .A(n26938), .B(n26937), .Z(n26940) );
  XNOR U25797 ( .A(n26935), .B(n26934), .Z(n26937) );
  XNOR U25798 ( .A(n26932), .B(n26931), .Z(n26934) );
  XNOR U25799 ( .A(n26929), .B(n26928), .Z(n26931) );
  XNOR U25800 ( .A(n26926), .B(n26925), .Z(n26928) );
  XNOR U25801 ( .A(n26923), .B(n26922), .Z(n26925) );
  XNOR U25802 ( .A(n26920), .B(n26919), .Z(n26922) );
  XNOR U25803 ( .A(n26917), .B(n26916), .Z(n26919) );
  XNOR U25804 ( .A(n26914), .B(n26913), .Z(n26916) );
  XNOR U25805 ( .A(n26911), .B(n26910), .Z(n26913) );
  XNOR U25806 ( .A(n26908), .B(n26907), .Z(n26910) );
  XNOR U25807 ( .A(n26905), .B(n26904), .Z(n26907) );
  XNOR U25808 ( .A(n26902), .B(n26901), .Z(n26904) );
  XNOR U25809 ( .A(n26899), .B(n26898), .Z(n26901) );
  XNOR U25810 ( .A(n26896), .B(n26895), .Z(n26898) );
  XNOR U25811 ( .A(n26893), .B(n26892), .Z(n26895) );
  XNOR U25812 ( .A(n26890), .B(n26889), .Z(n26892) );
  XNOR U25813 ( .A(n26887), .B(n26886), .Z(n26889) );
  XNOR U25814 ( .A(n26884), .B(n26883), .Z(n26886) );
  XNOR U25815 ( .A(n26881), .B(n26880), .Z(n26883) );
  XNOR U25816 ( .A(n26878), .B(n26877), .Z(n26880) );
  XNOR U25817 ( .A(n26875), .B(n26874), .Z(n26877) );
  XNOR U25818 ( .A(n26872), .B(n26871), .Z(n26874) );
  XNOR U25819 ( .A(n26869), .B(n26868), .Z(n26871) );
  XNOR U25820 ( .A(n26866), .B(n26865), .Z(n26868) );
  XNOR U25821 ( .A(n26863), .B(n26862), .Z(n26865) );
  XNOR U25822 ( .A(n26860), .B(n26859), .Z(n26862) );
  XNOR U25823 ( .A(n26857), .B(n26856), .Z(n26859) );
  XNOR U25824 ( .A(n26854), .B(n26853), .Z(n26856) );
  XNOR U25825 ( .A(n26851), .B(n26850), .Z(n26853) );
  XNOR U25826 ( .A(n26848), .B(n26847), .Z(n26850) );
  XNOR U25827 ( .A(n26845), .B(n26844), .Z(n26847) );
  XNOR U25828 ( .A(n26842), .B(n26841), .Z(n26844) );
  XNOR U25829 ( .A(n26839), .B(n26838), .Z(n26841) );
  XNOR U25830 ( .A(n26836), .B(n26835), .Z(n26838) );
  XNOR U25831 ( .A(n26833), .B(n26832), .Z(n26835) );
  XNOR U25832 ( .A(n26830), .B(n26829), .Z(n26832) );
  XNOR U25833 ( .A(n26827), .B(n26826), .Z(n26829) );
  XNOR U25834 ( .A(n26824), .B(n26823), .Z(n26826) );
  XNOR U25835 ( .A(n26821), .B(n26820), .Z(n26823) );
  XNOR U25836 ( .A(n26818), .B(n26817), .Z(n26820) );
  XNOR U25837 ( .A(n26815), .B(n26814), .Z(n26817) );
  XNOR U25838 ( .A(n26812), .B(n26811), .Z(n26814) );
  XNOR U25839 ( .A(n26809), .B(n26808), .Z(n26811) );
  XNOR U25840 ( .A(n26806), .B(n26805), .Z(n26808) );
  XNOR U25841 ( .A(n26803), .B(n26802), .Z(n26805) );
  XNOR U25842 ( .A(n26800), .B(n26799), .Z(n26802) );
  XNOR U25843 ( .A(n26797), .B(n26796), .Z(n26799) );
  XNOR U25844 ( .A(n26794), .B(n26793), .Z(n26796) );
  XNOR U25845 ( .A(n26791), .B(n26790), .Z(n26793) );
  XNOR U25846 ( .A(n26788), .B(n26787), .Z(n26790) );
  XNOR U25847 ( .A(n26785), .B(n26784), .Z(n26787) );
  XNOR U25848 ( .A(n26782), .B(n26781), .Z(n26784) );
  XNOR U25849 ( .A(n26779), .B(n26778), .Z(n26781) );
  XNOR U25850 ( .A(n26776), .B(n26775), .Z(n26778) );
  XNOR U25851 ( .A(n26773), .B(n26772), .Z(n26775) );
  XNOR U25852 ( .A(n26770), .B(n26769), .Z(n26772) );
  XNOR U25853 ( .A(n26767), .B(n26766), .Z(n26769) );
  XNOR U25854 ( .A(n26764), .B(n26763), .Z(n26766) );
  XNOR U25855 ( .A(n26761), .B(n26760), .Z(n26763) );
  XNOR U25856 ( .A(n26758), .B(n26757), .Z(n26760) );
  XNOR U25857 ( .A(n26755), .B(n26754), .Z(n26757) );
  XNOR U25858 ( .A(n26752), .B(n26751), .Z(n26754) );
  XNOR U25859 ( .A(n26749), .B(n26748), .Z(n26751) );
  XNOR U25860 ( .A(n26746), .B(n26745), .Z(n26748) );
  XNOR U25861 ( .A(n26743), .B(n26742), .Z(n26745) );
  XNOR U25862 ( .A(n26740), .B(n26739), .Z(n26742) );
  XNOR U25863 ( .A(n26737), .B(n26736), .Z(n26739) );
  XNOR U25864 ( .A(n26734), .B(n26733), .Z(n26736) );
  XNOR U25865 ( .A(n26731), .B(n26730), .Z(n26733) );
  XNOR U25866 ( .A(n26728), .B(n26727), .Z(n26730) );
  XNOR U25867 ( .A(n26725), .B(n26724), .Z(n26727) );
  XNOR U25868 ( .A(n26722), .B(n26721), .Z(n26724) );
  XNOR U25869 ( .A(n26719), .B(n26718), .Z(n26721) );
  XNOR U25870 ( .A(n26716), .B(n26715), .Z(n26718) );
  XNOR U25871 ( .A(n26713), .B(n26712), .Z(n26715) );
  XNOR U25872 ( .A(n26710), .B(n26709), .Z(n26712) );
  XNOR U25873 ( .A(n26707), .B(n26706), .Z(n26709) );
  XNOR U25874 ( .A(n26704), .B(n26703), .Z(n26706) );
  XNOR U25875 ( .A(n26701), .B(n26700), .Z(n26703) );
  XNOR U25876 ( .A(n26698), .B(n26697), .Z(n26700) );
  XNOR U25877 ( .A(n26695), .B(n26694), .Z(n26697) );
  XNOR U25878 ( .A(n26692), .B(n26691), .Z(n26694) );
  XNOR U25879 ( .A(n26689), .B(n26688), .Z(n26691) );
  XNOR U25880 ( .A(n26686), .B(n26685), .Z(n26688) );
  XNOR U25881 ( .A(n26683), .B(n26682), .Z(n26685) );
  XNOR U25882 ( .A(n26680), .B(n26679), .Z(n26682) );
  XNOR U25883 ( .A(n26677), .B(n26676), .Z(n26679) );
  XNOR U25884 ( .A(n26674), .B(n26673), .Z(n26676) );
  XNOR U25885 ( .A(n26671), .B(n26670), .Z(n26673) );
  XNOR U25886 ( .A(n26668), .B(n26667), .Z(n26670) );
  XNOR U25887 ( .A(n26665), .B(n26664), .Z(n26667) );
  XNOR U25888 ( .A(n26662), .B(n26661), .Z(n26664) );
  XNOR U25889 ( .A(n26659), .B(n26658), .Z(n26661) );
  XNOR U25890 ( .A(n26656), .B(n26655), .Z(n26658) );
  XNOR U25891 ( .A(n26653), .B(n26652), .Z(n26655) );
  XNOR U25892 ( .A(n26650), .B(n26649), .Z(n26652) );
  XNOR U25893 ( .A(n26647), .B(n26646), .Z(n26649) );
  XNOR U25894 ( .A(n26644), .B(n26643), .Z(n26646) );
  XNOR U25895 ( .A(n26641), .B(n26640), .Z(n26643) );
  XNOR U25896 ( .A(n26638), .B(n26637), .Z(n26640) );
  XNOR U25897 ( .A(n26635), .B(n26634), .Z(n26637) );
  XNOR U25898 ( .A(n26632), .B(n26631), .Z(n26634) );
  XNOR U25899 ( .A(n26629), .B(n26628), .Z(n26631) );
  XNOR U25900 ( .A(n26626), .B(n26625), .Z(n26628) );
  XNOR U25901 ( .A(n26623), .B(n26622), .Z(n26625) );
  XNOR U25902 ( .A(n26620), .B(n26619), .Z(n26622) );
  XNOR U25903 ( .A(n26617), .B(n26616), .Z(n26619) );
  XNOR U25904 ( .A(n26614), .B(n26613), .Z(n26616) );
  XNOR U25905 ( .A(n26611), .B(n26610), .Z(n26613) );
  XNOR U25906 ( .A(n26608), .B(n26607), .Z(n26610) );
  XNOR U25907 ( .A(n26605), .B(n26604), .Z(n26607) );
  XNOR U25908 ( .A(n26602), .B(n26601), .Z(n26604) );
  XNOR U25909 ( .A(n26599), .B(n26598), .Z(n26601) );
  XNOR U25910 ( .A(n26596), .B(n26595), .Z(n26598) );
  XNOR U25911 ( .A(n26593), .B(n26592), .Z(n26595) );
  XNOR U25912 ( .A(n26590), .B(n26589), .Z(n26592) );
  XNOR U25913 ( .A(n26587), .B(n26586), .Z(n26589) );
  XNOR U25914 ( .A(n26584), .B(n26583), .Z(n26586) );
  XNOR U25915 ( .A(n26581), .B(n26580), .Z(n26583) );
  XNOR U25916 ( .A(n26578), .B(n26577), .Z(n26580) );
  XNOR U25917 ( .A(n26575), .B(n26574), .Z(n26577) );
  XNOR U25918 ( .A(n26572), .B(n26571), .Z(n26574) );
  XNOR U25919 ( .A(n26569), .B(n26568), .Z(n26571) );
  XNOR U25920 ( .A(n26566), .B(n26565), .Z(n26568) );
  XNOR U25921 ( .A(n26563), .B(n26562), .Z(n26565) );
  XNOR U25922 ( .A(n26560), .B(n26559), .Z(n26562) );
  XNOR U25923 ( .A(n26557), .B(n26556), .Z(n26559) );
  XNOR U25924 ( .A(n26554), .B(n26553), .Z(n26556) );
  XNOR U25925 ( .A(n26551), .B(n26550), .Z(n26553) );
  XNOR U25926 ( .A(n26548), .B(n26547), .Z(n26550) );
  XNOR U25927 ( .A(n26545), .B(n26544), .Z(n26547) );
  XNOR U25928 ( .A(n26542), .B(n26541), .Z(n26544) );
  XNOR U25929 ( .A(n26539), .B(n26538), .Z(n26541) );
  XNOR U25930 ( .A(n26536), .B(n26535), .Z(n26538) );
  XNOR U25931 ( .A(n26533), .B(n26532), .Z(n26535) );
  XNOR U25932 ( .A(n26530), .B(n26529), .Z(n26532) );
  XNOR U25933 ( .A(n26527), .B(n26526), .Z(n26529) );
  XNOR U25934 ( .A(n26524), .B(n26523), .Z(n26526) );
  XNOR U25935 ( .A(n26521), .B(n26520), .Z(n26523) );
  XNOR U25936 ( .A(n26518), .B(n26517), .Z(n26520) );
  XNOR U25937 ( .A(n26515), .B(n26514), .Z(n26517) );
  XNOR U25938 ( .A(n26512), .B(n26511), .Z(n26514) );
  XNOR U25939 ( .A(n26509), .B(n26508), .Z(n26511) );
  XNOR U25940 ( .A(n26506), .B(n26505), .Z(n26508) );
  XNOR U25941 ( .A(n26503), .B(n26502), .Z(n26505) );
  XNOR U25942 ( .A(n26500), .B(n26499), .Z(n26502) );
  XNOR U25943 ( .A(n26497), .B(n26496), .Z(n26499) );
  XNOR U25944 ( .A(n26494), .B(n26493), .Z(n26496) );
  XNOR U25945 ( .A(n26491), .B(n26490), .Z(n26493) );
  XNOR U25946 ( .A(n26488), .B(n26487), .Z(n26490) );
  XNOR U25947 ( .A(n26485), .B(n26484), .Z(n26487) );
  XNOR U25948 ( .A(n26482), .B(n26481), .Z(n26484) );
  XNOR U25949 ( .A(n26479), .B(n26478), .Z(n26481) );
  XNOR U25950 ( .A(n26476), .B(n26475), .Z(n26478) );
  XNOR U25951 ( .A(n26473), .B(n26472), .Z(n26475) );
  XNOR U25952 ( .A(n26470), .B(n26469), .Z(n26472) );
  XNOR U25953 ( .A(n26467), .B(n26466), .Z(n26469) );
  XNOR U25954 ( .A(n26464), .B(n26463), .Z(n26466) );
  XNOR U25955 ( .A(n26461), .B(n26460), .Z(n26463) );
  XNOR U25956 ( .A(n26458), .B(n26457), .Z(n26460) );
  XNOR U25957 ( .A(n26455), .B(n26454), .Z(n26457) );
  XNOR U25958 ( .A(n26452), .B(n26451), .Z(n26454) );
  XNOR U25959 ( .A(n26449), .B(n26448), .Z(n26451) );
  XNOR U25960 ( .A(n26446), .B(n26445), .Z(n26448) );
  XNOR U25961 ( .A(n26443), .B(n26442), .Z(n26445) );
  XNOR U25962 ( .A(n26440), .B(n26439), .Z(n26442) );
  XNOR U25963 ( .A(n26437), .B(n26436), .Z(n26439) );
  XNOR U25964 ( .A(n26434), .B(n26433), .Z(n26436) );
  XNOR U25965 ( .A(n26431), .B(n26430), .Z(n26433) );
  XNOR U25966 ( .A(n26428), .B(n26427), .Z(n26430) );
  XNOR U25967 ( .A(n26425), .B(n26424), .Z(n26427) );
  XNOR U25968 ( .A(n26422), .B(n26421), .Z(n26424) );
  XNOR U25969 ( .A(n26419), .B(n26418), .Z(n26421) );
  XNOR U25970 ( .A(n26416), .B(n26415), .Z(n26418) );
  XNOR U25971 ( .A(n26413), .B(n26412), .Z(n26415) );
  XNOR U25972 ( .A(n26410), .B(n26409), .Z(n26412) );
  XNOR U25973 ( .A(n26407), .B(n26406), .Z(n26409) );
  XNOR U25974 ( .A(n26404), .B(n26403), .Z(n26406) );
  XNOR U25975 ( .A(n26401), .B(n26400), .Z(n26403) );
  XNOR U25976 ( .A(n26398), .B(n26397), .Z(n26400) );
  XNOR U25977 ( .A(n26395), .B(n26394), .Z(n26397) );
  XNOR U25978 ( .A(n26392), .B(n26391), .Z(n26394) );
  XNOR U25979 ( .A(n26389), .B(n26388), .Z(n26391) );
  XNOR U25980 ( .A(n26386), .B(n26385), .Z(n26388) );
  XNOR U25981 ( .A(n26383), .B(n26382), .Z(n26385) );
  XNOR U25982 ( .A(n26380), .B(n26379), .Z(n26382) );
  XNOR U25983 ( .A(n26377), .B(n26376), .Z(n26379) );
  XNOR U25984 ( .A(n26374), .B(n26373), .Z(n26376) );
  XNOR U25985 ( .A(n26371), .B(n26370), .Z(n26373) );
  XNOR U25986 ( .A(n26368), .B(n26367), .Z(n26370) );
  XNOR U25987 ( .A(n26365), .B(n26364), .Z(n26367) );
  XNOR U25988 ( .A(n26362), .B(n26361), .Z(n26364) );
  XNOR U25989 ( .A(n26359), .B(n26358), .Z(n26361) );
  XNOR U25990 ( .A(n26356), .B(n26355), .Z(n26358) );
  XNOR U25991 ( .A(n26353), .B(n26352), .Z(n26355) );
  XNOR U25992 ( .A(n26350), .B(n26349), .Z(n26352) );
  XNOR U25993 ( .A(n26347), .B(n26346), .Z(n26349) );
  XNOR U25994 ( .A(n26344), .B(n26343), .Z(n26346) );
  XNOR U25995 ( .A(n26341), .B(n26340), .Z(n26343) );
  XNOR U25996 ( .A(n26338), .B(n26337), .Z(n26340) );
  XNOR U25997 ( .A(n26335), .B(n26334), .Z(n26337) );
  XNOR U25998 ( .A(n26332), .B(n26331), .Z(n26334) );
  XNOR U25999 ( .A(n26329), .B(n26328), .Z(n26331) );
  XNOR U26000 ( .A(n26326), .B(n26325), .Z(n26328) );
  XNOR U26001 ( .A(n26323), .B(n26322), .Z(n26325) );
  XNOR U26002 ( .A(n26320), .B(n26319), .Z(n26322) );
  XNOR U26003 ( .A(n26317), .B(n26316), .Z(n26319) );
  XNOR U26004 ( .A(n26314), .B(n26313), .Z(n26316) );
  XNOR U26005 ( .A(n26311), .B(n26310), .Z(n26313) );
  XNOR U26006 ( .A(n26308), .B(n26307), .Z(n26310) );
  XNOR U26007 ( .A(n26305), .B(n26304), .Z(n26307) );
  XNOR U26008 ( .A(n26302), .B(n26301), .Z(n26304) );
  XNOR U26009 ( .A(n26299), .B(n26298), .Z(n26301) );
  XNOR U26010 ( .A(n26296), .B(n26295), .Z(n26298) );
  XNOR U26011 ( .A(n26293), .B(n26292), .Z(n26295) );
  XNOR U26012 ( .A(n26290), .B(n26289), .Z(n26292) );
  XNOR U26013 ( .A(n26287), .B(n26286), .Z(n26289) );
  XNOR U26014 ( .A(n26284), .B(n26283), .Z(n26286) );
  XNOR U26015 ( .A(n26281), .B(n26280), .Z(n26283) );
  XNOR U26016 ( .A(n26278), .B(n26277), .Z(n26280) );
  XNOR U26017 ( .A(n26275), .B(n26274), .Z(n26277) );
  XNOR U26018 ( .A(n26272), .B(n26271), .Z(n26274) );
  XNOR U26019 ( .A(n26269), .B(n26268), .Z(n26271) );
  XNOR U26020 ( .A(n26266), .B(n26265), .Z(n26268) );
  XNOR U26021 ( .A(n26263), .B(n26262), .Z(n26265) );
  XNOR U26022 ( .A(n26260), .B(n26259), .Z(n26262) );
  XNOR U26023 ( .A(n26257), .B(n26256), .Z(n26259) );
  XNOR U26024 ( .A(n26254), .B(n26253), .Z(n26256) );
  XNOR U26025 ( .A(n26251), .B(n26250), .Z(n26253) );
  XNOR U26026 ( .A(n26248), .B(n26247), .Z(n26250) );
  XNOR U26027 ( .A(n26245), .B(n26244), .Z(n26247) );
  XNOR U26028 ( .A(n26242), .B(n26241), .Z(n26244) );
  XNOR U26029 ( .A(n26239), .B(n26238), .Z(n26241) );
  XNOR U26030 ( .A(n26236), .B(n26235), .Z(n26238) );
  XNOR U26031 ( .A(n26233), .B(n26232), .Z(n26235) );
  XNOR U26032 ( .A(n26230), .B(n26229), .Z(n26232) );
  XNOR U26033 ( .A(n26227), .B(n26226), .Z(n26229) );
  XNOR U26034 ( .A(n26224), .B(n26223), .Z(n26226) );
  XNOR U26035 ( .A(n26221), .B(n26220), .Z(n26223) );
  XNOR U26036 ( .A(n26218), .B(n26217), .Z(n26220) );
  XNOR U26037 ( .A(n26215), .B(n26214), .Z(n26217) );
  XNOR U26038 ( .A(n26212), .B(n26211), .Z(n26214) );
  XNOR U26039 ( .A(n26209), .B(n26208), .Z(n26211) );
  XNOR U26040 ( .A(n26206), .B(n26205), .Z(n26208) );
  XNOR U26041 ( .A(n26203), .B(n26202), .Z(n26205) );
  XNOR U26042 ( .A(n26200), .B(n26199), .Z(n26202) );
  XNOR U26043 ( .A(n26197), .B(n26196), .Z(n26199) );
  XNOR U26044 ( .A(n26194), .B(n26193), .Z(n26196) );
  XNOR U26045 ( .A(n26191), .B(n26190), .Z(n26193) );
  XNOR U26046 ( .A(n26188), .B(n26187), .Z(n26190) );
  XNOR U26047 ( .A(n26185), .B(n26184), .Z(n26187) );
  XNOR U26048 ( .A(n26182), .B(n26180), .Z(n26184) );
  XNOR U26049 ( .A(n26181), .B(n25548), .Z(n26180) );
  XNOR U26050 ( .A(n25549), .B(n25546), .Z(n25548) );
  XNOR U26051 ( .A(n25547), .B(n25550), .Z(n25546) );
  XNOR U26052 ( .A(n25551), .B(n26175), .Z(n25550) );
  XNOR U26053 ( .A(n25558), .B(n26174), .Z(n26175) );
  XNOR U26054 ( .A(n26167), .B(n26171), .Z(n26174) );
  XNOR U26055 ( .A(n26166), .B(n26164), .Z(n26171) );
  XNOR U26056 ( .A(n26165), .B(n26163), .Z(n26164) );
  XNOR U26057 ( .A(n25565), .B(n26158), .Z(n26163) );
  XNOR U26058 ( .A(n25564), .B(n26156), .Z(n26158) );
  XNOR U26059 ( .A(n26157), .B(n26152), .Z(n26156) );
  XNOR U26060 ( .A(n26153), .B(n25580), .Z(n26152) );
  XNOR U26061 ( .A(n25575), .B(n26151), .Z(n25580) );
  XNOR U26062 ( .A(n25574), .B(n26146), .Z(n26151) );
  XNOR U26063 ( .A(n25576), .B(n26145), .Z(n26146) );
  XNOR U26064 ( .A(n25579), .B(n26142), .Z(n26145) );
  XNOR U26065 ( .A(n25585), .B(n26141), .Z(n26142) );
  XNOR U26066 ( .A(n26134), .B(n26138), .Z(n26141) );
  XNOR U26067 ( .A(n26133), .B(n26131), .Z(n26138) );
  XNOR U26068 ( .A(n26132), .B(n26130), .Z(n26131) );
  XNOR U26069 ( .A(n25592), .B(n26125), .Z(n26130) );
  XNOR U26070 ( .A(n25591), .B(n26123), .Z(n26125) );
  XNOR U26071 ( .A(n26124), .B(n26119), .Z(n26123) );
  XNOR U26072 ( .A(n26120), .B(n25607), .Z(n26119) );
  XNOR U26073 ( .A(n25602), .B(n26118), .Z(n25607) );
  XNOR U26074 ( .A(n25601), .B(n26113), .Z(n26118) );
  XNOR U26075 ( .A(n25603), .B(n26112), .Z(n26113) );
  XNOR U26076 ( .A(n25606), .B(n26109), .Z(n26112) );
  XNOR U26077 ( .A(n25612), .B(n26108), .Z(n26109) );
  XNOR U26078 ( .A(n26101), .B(n26105), .Z(n26108) );
  XNOR U26079 ( .A(n26100), .B(n26098), .Z(n26105) );
  XNOR U26080 ( .A(n26099), .B(n26097), .Z(n26098) );
  XNOR U26081 ( .A(n25619), .B(n26092), .Z(n26097) );
  XNOR U26082 ( .A(n25618), .B(n26090), .Z(n26092) );
  XNOR U26083 ( .A(n26091), .B(n26086), .Z(n26090) );
  XNOR U26084 ( .A(n26087), .B(n25634), .Z(n26086) );
  XNOR U26085 ( .A(n25629), .B(n26085), .Z(n25634) );
  XNOR U26086 ( .A(n25628), .B(n26080), .Z(n26085) );
  XNOR U26087 ( .A(n25630), .B(n26079), .Z(n26080) );
  XNOR U26088 ( .A(n25633), .B(n26076), .Z(n26079) );
  XNOR U26089 ( .A(n25639), .B(n26075), .Z(n26076) );
  XNOR U26090 ( .A(n26068), .B(n26072), .Z(n26075) );
  XNOR U26091 ( .A(n26067), .B(n26065), .Z(n26072) );
  XNOR U26092 ( .A(n26066), .B(n26064), .Z(n26065) );
  XNOR U26093 ( .A(n25646), .B(n26059), .Z(n26064) );
  XNOR U26094 ( .A(n25645), .B(n26057), .Z(n26059) );
  XNOR U26095 ( .A(n26058), .B(n26053), .Z(n26057) );
  XNOR U26096 ( .A(n26054), .B(n25661), .Z(n26053) );
  XNOR U26097 ( .A(n25656), .B(n26052), .Z(n25661) );
  XNOR U26098 ( .A(n25655), .B(n26047), .Z(n26052) );
  XNOR U26099 ( .A(n25657), .B(n26046), .Z(n26047) );
  XNOR U26100 ( .A(n25660), .B(n26043), .Z(n26046) );
  XNOR U26101 ( .A(n25666), .B(n26042), .Z(n26043) );
  XNOR U26102 ( .A(n26035), .B(n26039), .Z(n26042) );
  XNOR U26103 ( .A(n26034), .B(n26032), .Z(n26039) );
  XNOR U26104 ( .A(n26033), .B(n26031), .Z(n26032) );
  XNOR U26105 ( .A(n25673), .B(n26026), .Z(n26031) );
  XNOR U26106 ( .A(n25672), .B(n26024), .Z(n26026) );
  XNOR U26107 ( .A(n26025), .B(n26020), .Z(n26024) );
  XNOR U26108 ( .A(n26021), .B(n25688), .Z(n26020) );
  XNOR U26109 ( .A(n25683), .B(n26019), .Z(n25688) );
  XNOR U26110 ( .A(n25682), .B(n26014), .Z(n26019) );
  XNOR U26111 ( .A(n25684), .B(n26013), .Z(n26014) );
  XNOR U26112 ( .A(n25687), .B(n26010), .Z(n26013) );
  XNOR U26113 ( .A(n25693), .B(n26009), .Z(n26010) );
  XNOR U26114 ( .A(n26002), .B(n26006), .Z(n26009) );
  XNOR U26115 ( .A(n26001), .B(n25999), .Z(n26006) );
  XNOR U26116 ( .A(n26000), .B(n25998), .Z(n25999) );
  XNOR U26117 ( .A(n25700), .B(n25993), .Z(n25998) );
  XNOR U26118 ( .A(n25699), .B(n25991), .Z(n25993) );
  XNOR U26119 ( .A(n25992), .B(n25987), .Z(n25991) );
  XNOR U26120 ( .A(n25988), .B(n25715), .Z(n25987) );
  XNOR U26121 ( .A(n25710), .B(n25986), .Z(n25715) );
  XNOR U26122 ( .A(n25709), .B(n25981), .Z(n25986) );
  XNOR U26123 ( .A(n25711), .B(n25980), .Z(n25981) );
  XNOR U26124 ( .A(n25714), .B(n25977), .Z(n25980) );
  XNOR U26125 ( .A(n25720), .B(n25976), .Z(n25977) );
  XNOR U26126 ( .A(n25969), .B(n25973), .Z(n25976) );
  XNOR U26127 ( .A(n25968), .B(n25966), .Z(n25973) );
  XNOR U26128 ( .A(n25967), .B(n25965), .Z(n25966) );
  XNOR U26129 ( .A(n25727), .B(n25960), .Z(n25965) );
  XNOR U26130 ( .A(n25726), .B(n25958), .Z(n25960) );
  XNOR U26131 ( .A(n25959), .B(n25954), .Z(n25958) );
  XNOR U26132 ( .A(n25955), .B(n25742), .Z(n25954) );
  XNOR U26133 ( .A(n25737), .B(n25953), .Z(n25742) );
  XNOR U26134 ( .A(n25736), .B(n25948), .Z(n25953) );
  XNOR U26135 ( .A(n25738), .B(n25947), .Z(n25948) );
  XNOR U26136 ( .A(n25741), .B(n25944), .Z(n25947) );
  XNOR U26137 ( .A(n25747), .B(n25943), .Z(n25944) );
  XNOR U26138 ( .A(n25936), .B(n25940), .Z(n25943) );
  XNOR U26139 ( .A(n25935), .B(n25933), .Z(n25940) );
  XNOR U26140 ( .A(n25934), .B(n25932), .Z(n25933) );
  XNOR U26141 ( .A(n25754), .B(n25927), .Z(n25932) );
  XNOR U26142 ( .A(n25753), .B(n25925), .Z(n25927) );
  XNOR U26143 ( .A(n25926), .B(n25921), .Z(n25925) );
  XNOR U26144 ( .A(n25922), .B(n25769), .Z(n25921) );
  XNOR U26145 ( .A(n25764), .B(n25920), .Z(n25769) );
  XNOR U26146 ( .A(n25763), .B(n25915), .Z(n25920) );
  XNOR U26147 ( .A(n25765), .B(n25914), .Z(n25915) );
  XNOR U26148 ( .A(n25768), .B(n25911), .Z(n25914) );
  XNOR U26149 ( .A(n25774), .B(n25910), .Z(n25911) );
  XNOR U26150 ( .A(n25903), .B(n25907), .Z(n25910) );
  XNOR U26151 ( .A(n25902), .B(n25900), .Z(n25907) );
  XNOR U26152 ( .A(n25901), .B(n25899), .Z(n25900) );
  XNOR U26153 ( .A(n25781), .B(n25894), .Z(n25899) );
  XNOR U26154 ( .A(n25780), .B(n25892), .Z(n25894) );
  XNOR U26155 ( .A(n25893), .B(n25888), .Z(n25892) );
  XNOR U26156 ( .A(n25889), .B(n25796), .Z(n25888) );
  XNOR U26157 ( .A(n25791), .B(n25887), .Z(n25796) );
  XNOR U26158 ( .A(n25790), .B(n25882), .Z(n25887) );
  XNOR U26159 ( .A(n25792), .B(n25881), .Z(n25882) );
  XNOR U26160 ( .A(n25795), .B(n25878), .Z(n25881) );
  XNOR U26161 ( .A(n25801), .B(n25877), .Z(n25878) );
  XNOR U26162 ( .A(n25870), .B(n25874), .Z(n25877) );
  XNOR U26163 ( .A(n25869), .B(n25867), .Z(n25874) );
  XNOR U26164 ( .A(n25868), .B(n25866), .Z(n25867) );
  XNOR U26165 ( .A(n25808), .B(n25861), .Z(n25866) );
  XNOR U26166 ( .A(n25807), .B(n25859), .Z(n25861) );
  XNOR U26167 ( .A(n25860), .B(n25855), .Z(n25859) );
  XNOR U26168 ( .A(n25856), .B(n25823), .Z(n25855) );
  XNOR U26169 ( .A(n25818), .B(n25854), .Z(n25823) );
  XNOR U26170 ( .A(n25817), .B(n25849), .Z(n25854) );
  XNOR U26171 ( .A(n25819), .B(n25848), .Z(n25849) );
  XNOR U26172 ( .A(n25822), .B(n25845), .Z(n25848) );
  XNOR U26173 ( .A(n25828), .B(n25844), .Z(n25845) );
  XNOR U26174 ( .A(n25831), .B(n25841), .Z(n25844) );
  XNOR U26175 ( .A(n25830), .B(n25838), .Z(n25841) );
  XOR U26176 ( .A(n25839), .B(n25837), .Z(n25838) );
  XNOR U26177 ( .A(n28369), .B(n28370), .Z(n25837) );
  XOR U26178 ( .A(n28371), .B(n28372), .Z(n28370) );
  XOR U26179 ( .A(n28373), .B(n28374), .Z(n28372) );
  NOR U26180 ( .A(n28375), .B(n28376), .Z(n28373) );
  XOR U26181 ( .A(n28377), .B(n28378), .Z(n28371) );
  NOR U26182 ( .A(n28379), .B(n28380), .Z(n28378) );
  AND U26183 ( .A(n28381), .B(n28382), .Z(n28377) );
  XOR U26184 ( .A(n28383), .B(n28384), .Z(n28369) );
  XOR U26185 ( .A(n28376), .B(n28380), .Z(n28384) );
  XOR U26186 ( .A(n28385), .B(n28382), .Z(n28383) );
  XOR U26187 ( .A(n28386), .B(n28387), .Z(n28385) );
  XOR U26188 ( .A(n28388), .B(n28389), .Z(n28387) );
  XOR U26189 ( .A(n28390), .B(n28391), .Z(n28389) );
  XOR U26190 ( .A(n28392), .B(n28393), .Z(n28388) );
  NOR U26191 ( .A(n28394), .B(n28395), .Z(n28393) );
  AND U26192 ( .A(n28396), .B(n28374), .Z(n28392) );
  XOR U26193 ( .A(n28397), .B(n28398), .Z(n28386) );
  XOR U26194 ( .A(n28399), .B(n28400), .Z(n28398) );
  XOR U26195 ( .A(n28401), .B(n28402), .Z(n28400) );
  XOR U26196 ( .A(n28403), .B(n28404), .Z(n28402) );
  XOR U26197 ( .A(n28405), .B(n28406), .Z(n28404) );
  XOR U26198 ( .A(n28407), .B(n28408), .Z(n28406) );
  XNOR U26199 ( .A(n28409), .B(n28410), .Z(n28405) );
  XOR U26200 ( .A(n28411), .B(n28412), .Z(n28410) );
  NOR U26201 ( .A(n28413), .B(n28408), .Z(n28411) );
  XOR U26202 ( .A(n28414), .B(n28415), .Z(n28403) );
  XOR U26203 ( .A(n28416), .B(n28417), .Z(n28415) );
  XOR U26204 ( .A(n28418), .B(n28419), .Z(n28417) );
  XOR U26205 ( .A(n28420), .B(n28421), .Z(n28419) );
  XOR U26206 ( .A(n28422), .B(n28423), .Z(n28421) );
  XOR U26207 ( .A(n28424), .B(n28425), .Z(n28423) );
  XOR U26208 ( .A(n28426), .B(n28427), .Z(n28425) );
  XOR U26209 ( .A(n28428), .B(n28429), .Z(n28427) );
  NOR U26210 ( .A(n28430), .B(n28431), .Z(n28429) );
  XOR U26211 ( .A(n28432), .B(n28433), .Z(n28426) );
  AND U26212 ( .A(n28428), .B(n28434), .Z(n28432) );
  XOR U26213 ( .A(n28435), .B(n28436), .Z(n28424) );
  XOR U26214 ( .A(n28437), .B(n28438), .Z(n28436) );
  XOR U26215 ( .A(n28439), .B(n28440), .Z(n28438) );
  XOR U26216 ( .A(n28441), .B(n28442), .Z(n28440) );
  XOR U26217 ( .A(n28443), .B(n28444), .Z(n28442) );
  XOR U26218 ( .A(n28445), .B(n28446), .Z(n28444) );
  XOR U26219 ( .A(n28447), .B(n28448), .Z(n28446) );
  XOR U26220 ( .A(n28449), .B(n28450), .Z(n28448) );
  XOR U26221 ( .A(n28451), .B(n28452), .Z(n28450) );
  AND U26222 ( .A(n28453), .B(n28454), .Z(n28452) );
  NOR U26223 ( .A(n28455), .B(n28456), .Z(n28454) );
  NOR U26224 ( .A(n28457), .B(n28458), .Z(n28453) );
  AND U26225 ( .A(n28459), .B(n28460), .Z(n28458) );
  AND U26226 ( .A(n28461), .B(n28462), .Z(n28451) );
  NOR U26227 ( .A(n28463), .B(n28464), .Z(n28462) );
  NOR U26228 ( .A(n28465), .B(n28466), .Z(n28461) );
  AND U26229 ( .A(n28467), .B(n28468), .Z(n28466) );
  XOR U26230 ( .A(n28469), .B(n28470), .Z(n28449) );
  AND U26231 ( .A(n28471), .B(n28472), .Z(n28470) );
  NOR U26232 ( .A(n28473), .B(n28474), .Z(n28472) );
  NOR U26233 ( .A(n28475), .B(n28476), .Z(n28471) );
  AND U26234 ( .A(n28477), .B(n28478), .Z(n28476) );
  AND U26235 ( .A(n28479), .B(n28480), .Z(n28469) );
  NOR U26236 ( .A(n28481), .B(n28482), .Z(n28480) );
  AND U26237 ( .A(n28474), .B(n28483), .Z(n28482) );
  AND U26238 ( .A(n28475), .B(n28484), .Z(n28481) );
  NOR U26239 ( .A(n28485), .B(n28486), .Z(n28479) );
  XOR U26240 ( .A(n28487), .B(n28488), .Z(n28486) );
  AND U26241 ( .A(n28489), .B(n28490), .Z(n28488) );
  NOR U26242 ( .A(n28491), .B(n28492), .Z(n28490) );
  NOR U26243 ( .A(n28493), .B(n28494), .Z(n28489) );
  AND U26244 ( .A(n28495), .B(n28496), .Z(n28494) );
  AND U26245 ( .A(n28497), .B(n28498), .Z(n28487) );
  NOR U26246 ( .A(n28499), .B(n28500), .Z(n28498) );
  AND U26247 ( .A(n28492), .B(n28501), .Z(n28500) );
  AND U26248 ( .A(n28493), .B(n28502), .Z(n28499) );
  NOR U26249 ( .A(n28503), .B(n28504), .Z(n28497) );
  XOR U26250 ( .A(n28505), .B(n28506), .Z(n28504) );
  AND U26251 ( .A(n28507), .B(n28508), .Z(n28506) );
  NOR U26252 ( .A(n28509), .B(n28510), .Z(n28508) );
  NOR U26253 ( .A(n28511), .B(n28512), .Z(n28507) );
  AND U26254 ( .A(n28513), .B(n28514), .Z(n28512) );
  AND U26255 ( .A(n28515), .B(n28516), .Z(n28505) );
  AND U26256 ( .A(n28517), .B(n28518), .Z(n28516) );
  IV U26257 ( .A(n28509), .Z(n28517) );
  NOR U26258 ( .A(n28511), .B(n28519), .Z(n28515) );
  AND U26259 ( .A(n28520), .B(n28521), .Z(n28519) );
  AND U26260 ( .A(n28522), .B(n28523), .Z(n28521) );
  NOR U26261 ( .A(n28524), .B(n28525), .Z(n28522) );
  NOR U26262 ( .A(n28526), .B(n28527), .Z(n28520) );
  AND U26263 ( .A(n28491), .B(n28528), .Z(n28503) );
  AND U26264 ( .A(n28473), .B(n28529), .Z(n28485) );
  XOR U26265 ( .A(n28530), .B(n28531), .Z(n28447) );
  XOR U26266 ( .A(n28532), .B(n28533), .Z(n28531) );
  NOR U26267 ( .A(n28534), .B(n28535), .Z(n28533) );
  AND U26268 ( .A(n28464), .B(n28536), .Z(n28535) );
  AND U26269 ( .A(n28465), .B(n28537), .Z(n28534) );
  NOR U26270 ( .A(n28538), .B(n28539), .Z(n28532) );
  AND U26271 ( .A(n28456), .B(n28540), .Z(n28539) );
  AND U26272 ( .A(n28457), .B(n28541), .Z(n28538) );
  XOR U26273 ( .A(n28542), .B(n28543), .Z(n28530) );
  AND U26274 ( .A(n28463), .B(n28544), .Z(n28543) );
  AND U26275 ( .A(n28455), .B(n28545), .Z(n28542) );
  AND U26276 ( .A(n28546), .B(n28547), .Z(n28445) );
  NOR U26277 ( .A(n28548), .B(n28549), .Z(n28547) );
  NOR U26278 ( .A(n28550), .B(n28551), .Z(n28546) );
  AND U26279 ( .A(n28552), .B(n28553), .Z(n28551) );
  XOR U26280 ( .A(n28554), .B(n28555), .Z(n28443) );
  AND U26281 ( .A(n28556), .B(n28557), .Z(n28555) );
  NOR U26282 ( .A(n28558), .B(n28559), .Z(n28557) );
  NOR U26283 ( .A(n28560), .B(n28561), .Z(n28556) );
  AND U26284 ( .A(n28562), .B(n28563), .Z(n28561) );
  NOR U26285 ( .A(n28564), .B(n28565), .Z(n28554) );
  AND U26286 ( .A(n28559), .B(n28566), .Z(n28565) );
  AND U26287 ( .A(n28560), .B(n28567), .Z(n28564) );
  XOR U26288 ( .A(n28568), .B(n28569), .Z(n28441) );
  XOR U26289 ( .A(n28570), .B(n28571), .Z(n28569) );
  NOR U26290 ( .A(n28572), .B(n28573), .Z(n28571) );
  AND U26291 ( .A(n28549), .B(n28574), .Z(n28573) );
  AND U26292 ( .A(n28550), .B(n28575), .Z(n28572) );
  AND U26293 ( .A(n28558), .B(n28576), .Z(n28570) );
  XOR U26294 ( .A(n28577), .B(n28578), .Z(n28568) );
  AND U26295 ( .A(n28548), .B(n28579), .Z(n28578) );
  AND U26296 ( .A(n28580), .B(n28581), .Z(n28577) );
  AND U26297 ( .A(n28582), .B(n28583), .Z(n28439) );
  NOR U26298 ( .A(n28584), .B(n28585), .Z(n28583) );
  NOR U26299 ( .A(n28586), .B(n28587), .Z(n28582) );
  AND U26300 ( .A(n28588), .B(n28589), .Z(n28587) );
  XOR U26301 ( .A(n28590), .B(n28591), .Z(n28437) );
  AND U26302 ( .A(n28592), .B(n28593), .Z(n28591) );
  NOR U26303 ( .A(n28580), .B(n28594), .Z(n28593) );
  NOR U26304 ( .A(n28595), .B(n28596), .Z(n28592) );
  AND U26305 ( .A(n28597), .B(n28598), .Z(n28596) );
  NOR U26306 ( .A(n28599), .B(n28600), .Z(n28590) );
  AND U26307 ( .A(n28594), .B(n28601), .Z(n28600) );
  AND U26308 ( .A(n28595), .B(n28602), .Z(n28599) );
  XOR U26309 ( .A(n28603), .B(n28604), .Z(n28435) );
  XOR U26310 ( .A(n28605), .B(n28606), .Z(n28604) );
  NOR U26311 ( .A(n28607), .B(n28608), .Z(n28606) );
  AND U26312 ( .A(n28585), .B(n28609), .Z(n28608) );
  AND U26313 ( .A(n28586), .B(n28610), .Z(n28607) );
  NOR U26314 ( .A(n28611), .B(n28612), .Z(n28605) );
  AND U26315 ( .A(n28613), .B(n28614), .Z(n28612) );
  AND U26316 ( .A(n28615), .B(n28616), .Z(n28611) );
  XOR U26317 ( .A(n28617), .B(n28618), .Z(n28603) );
  AND U26318 ( .A(n28584), .B(n28619), .Z(n28618) );
  AND U26319 ( .A(n28620), .B(n28621), .Z(n28617) );
  XOR U26320 ( .A(n28622), .B(n28623), .Z(n28422) );
  NOR U26321 ( .A(n28615), .B(n28624), .Z(n28623) );
  AND U26322 ( .A(n28625), .B(n28626), .Z(n28624) );
  NOR U26323 ( .A(n28620), .B(n28613), .Z(n28622) );
  XOR U26324 ( .A(n28627), .B(n28628), .Z(n28420) );
  XOR U26325 ( .A(n28629), .B(n28630), .Z(n28628) );
  AND U26326 ( .A(n28430), .B(n28631), .Z(n28630) );
  AND U26327 ( .A(n28431), .B(n28632), .Z(n28629) );
  XOR U26328 ( .A(n28633), .B(n28634), .Z(n28627) );
  AND U26329 ( .A(n28433), .B(n28635), .Z(n28634) );
  AND U26330 ( .A(n28636), .B(n28637), .Z(n28633) );
  XNOR U26331 ( .A(n28638), .B(n28639), .Z(n28416) );
  XOR U26332 ( .A(n28640), .B(n28641), .Z(n28414) );
  XOR U26333 ( .A(n28642), .B(n28636), .Z(n28641) );
  AND U26334 ( .A(n28643), .B(n28638), .Z(n28642) );
  XOR U26335 ( .A(n28644), .B(n28645), .Z(n28640) );
  AND U26336 ( .A(n28646), .B(n28647), .Z(n28645) );
  AND U26337 ( .A(n28648), .B(n28418), .Z(n28644) );
  XOR U26338 ( .A(n28649), .B(n28650), .Z(n28401) );
  AND U26339 ( .A(n28651), .B(n28412), .Z(n28650) );
  NOR U26340 ( .A(n28652), .B(n28409), .Z(n28649) );
  XOR U26341 ( .A(n28653), .B(n28654), .Z(n28399) );
  XOR U26342 ( .A(n28655), .B(n28656), .Z(n28654) );
  NOR U26343 ( .A(n28657), .B(n28407), .Z(n28656) );
  NOR U26344 ( .A(n28658), .B(n28390), .Z(n28655) );
  XOR U26345 ( .A(n28659), .B(n28660), .Z(n28653) );
  NOR U26346 ( .A(n28661), .B(n28391), .Z(n28660) );
  NOR U26347 ( .A(n28662), .B(n28663), .Z(n28659) );
  XNOR U26348 ( .A(n28395), .B(n28663), .Z(n28397) );
  XOR U26349 ( .A(n28664), .B(n28665), .Z(n25839) );
  NOR U26350 ( .A(n28666), .B(n28664), .Z(n28665) );
  XOR U26351 ( .A(n28667), .B(n28668), .Z(n25830) );
  NOR U26352 ( .A(n28669), .B(n28667), .Z(n28668) );
  XOR U26353 ( .A(n28670), .B(n28671), .Z(n25831) );
  NOR U26354 ( .A(n28672), .B(n28670), .Z(n28671) );
  XOR U26355 ( .A(n28673), .B(n28674), .Z(n25828) );
  NOR U26356 ( .A(n28675), .B(n28673), .Z(n28674) );
  XOR U26357 ( .A(n28676), .B(n28677), .Z(n25822) );
  NOR U26358 ( .A(n28678), .B(n28676), .Z(n28677) );
  XOR U26359 ( .A(n28679), .B(n28680), .Z(n25819) );
  NOR U26360 ( .A(n28681), .B(n28679), .Z(n28680) );
  XOR U26361 ( .A(n28682), .B(n28683), .Z(n25817) );
  NOR U26362 ( .A(n28684), .B(n28682), .Z(n28683) );
  XOR U26363 ( .A(n28685), .B(n28686), .Z(n25818) );
  NOR U26364 ( .A(n28687), .B(n28685), .Z(n28686) );
  XOR U26365 ( .A(n28688), .B(n28689), .Z(n25856) );
  NOR U26366 ( .A(n28690), .B(n28688), .Z(n28689) );
  XOR U26367 ( .A(n28691), .B(n28692), .Z(n25860) );
  NOR U26368 ( .A(n28693), .B(n28691), .Z(n28692) );
  XOR U26369 ( .A(n28694), .B(n28695), .Z(n25807) );
  NOR U26370 ( .A(n28696), .B(n28694), .Z(n28695) );
  XOR U26371 ( .A(n28697), .B(n28698), .Z(n25808) );
  NOR U26372 ( .A(n28699), .B(n28697), .Z(n28698) );
  XOR U26373 ( .A(n28700), .B(n28701), .Z(n25868) );
  NOR U26374 ( .A(n28702), .B(n28700), .Z(n28701) );
  XOR U26375 ( .A(n28703), .B(n28704), .Z(n25869) );
  NOR U26376 ( .A(n28705), .B(n28703), .Z(n28704) );
  XOR U26377 ( .A(n28706), .B(n28707), .Z(n25870) );
  NOR U26378 ( .A(n28708), .B(n28706), .Z(n28707) );
  XOR U26379 ( .A(n28709), .B(n28710), .Z(n25801) );
  NOR U26380 ( .A(n28711), .B(n28709), .Z(n28710) );
  XOR U26381 ( .A(n28712), .B(n28713), .Z(n25795) );
  NOR U26382 ( .A(n28714), .B(n28712), .Z(n28713) );
  XOR U26383 ( .A(n28715), .B(n28716), .Z(n25792) );
  NOR U26384 ( .A(n28717), .B(n28715), .Z(n28716) );
  XOR U26385 ( .A(n28718), .B(n28719), .Z(n25790) );
  NOR U26386 ( .A(n28720), .B(n28718), .Z(n28719) );
  XOR U26387 ( .A(n28721), .B(n28722), .Z(n25791) );
  NOR U26388 ( .A(n28723), .B(n28721), .Z(n28722) );
  XOR U26389 ( .A(n28724), .B(n28725), .Z(n25889) );
  NOR U26390 ( .A(n28726), .B(n28724), .Z(n28725) );
  XOR U26391 ( .A(n28727), .B(n28728), .Z(n25893) );
  NOR U26392 ( .A(n28729), .B(n28727), .Z(n28728) );
  XOR U26393 ( .A(n28730), .B(n28731), .Z(n25780) );
  NOR U26394 ( .A(n28732), .B(n28730), .Z(n28731) );
  XOR U26395 ( .A(n28733), .B(n28734), .Z(n25781) );
  NOR U26396 ( .A(n28735), .B(n28733), .Z(n28734) );
  XOR U26397 ( .A(n28736), .B(n28737), .Z(n25901) );
  NOR U26398 ( .A(n28738), .B(n28736), .Z(n28737) );
  XOR U26399 ( .A(n28739), .B(n28740), .Z(n25902) );
  NOR U26400 ( .A(n28741), .B(n28739), .Z(n28740) );
  XOR U26401 ( .A(n28742), .B(n28743), .Z(n25903) );
  NOR U26402 ( .A(n28744), .B(n28742), .Z(n28743) );
  XOR U26403 ( .A(n28745), .B(n28746), .Z(n25774) );
  NOR U26404 ( .A(n28747), .B(n28745), .Z(n28746) );
  XOR U26405 ( .A(n28748), .B(n28749), .Z(n25768) );
  NOR U26406 ( .A(n28750), .B(n28748), .Z(n28749) );
  XOR U26407 ( .A(n28751), .B(n28752), .Z(n25765) );
  NOR U26408 ( .A(n28753), .B(n28751), .Z(n28752) );
  XOR U26409 ( .A(n28754), .B(n28755), .Z(n25763) );
  NOR U26410 ( .A(n28756), .B(n28754), .Z(n28755) );
  XOR U26411 ( .A(n28757), .B(n28758), .Z(n25764) );
  NOR U26412 ( .A(n28759), .B(n28757), .Z(n28758) );
  XOR U26413 ( .A(n28760), .B(n28761), .Z(n25922) );
  NOR U26414 ( .A(n28762), .B(n28760), .Z(n28761) );
  XOR U26415 ( .A(n28763), .B(n28764), .Z(n25926) );
  NOR U26416 ( .A(n28765), .B(n28763), .Z(n28764) );
  XOR U26417 ( .A(n28766), .B(n28767), .Z(n25753) );
  NOR U26418 ( .A(n28768), .B(n28766), .Z(n28767) );
  XOR U26419 ( .A(n28769), .B(n28770), .Z(n25754) );
  NOR U26420 ( .A(n28771), .B(n28769), .Z(n28770) );
  XOR U26421 ( .A(n28772), .B(n28773), .Z(n25934) );
  NOR U26422 ( .A(n28774), .B(n28772), .Z(n28773) );
  XOR U26423 ( .A(n28775), .B(n28776), .Z(n25935) );
  NOR U26424 ( .A(n28777), .B(n28775), .Z(n28776) );
  XOR U26425 ( .A(n28778), .B(n28779), .Z(n25936) );
  NOR U26426 ( .A(n28780), .B(n28778), .Z(n28779) );
  XOR U26427 ( .A(n28781), .B(n28782), .Z(n25747) );
  NOR U26428 ( .A(n28783), .B(n28781), .Z(n28782) );
  XOR U26429 ( .A(n28784), .B(n28785), .Z(n25741) );
  NOR U26430 ( .A(n28786), .B(n28784), .Z(n28785) );
  XOR U26431 ( .A(n28787), .B(n28788), .Z(n25738) );
  NOR U26432 ( .A(n28789), .B(n28787), .Z(n28788) );
  XOR U26433 ( .A(n28790), .B(n28791), .Z(n25736) );
  NOR U26434 ( .A(n28792), .B(n28790), .Z(n28791) );
  XOR U26435 ( .A(n28793), .B(n28794), .Z(n25737) );
  NOR U26436 ( .A(n28795), .B(n28793), .Z(n28794) );
  XOR U26437 ( .A(n28796), .B(n28797), .Z(n25955) );
  NOR U26438 ( .A(n28798), .B(n28796), .Z(n28797) );
  XOR U26439 ( .A(n28799), .B(n28800), .Z(n25959) );
  NOR U26440 ( .A(n28801), .B(n28799), .Z(n28800) );
  XOR U26441 ( .A(n28802), .B(n28803), .Z(n25726) );
  NOR U26442 ( .A(n28804), .B(n28802), .Z(n28803) );
  XOR U26443 ( .A(n28805), .B(n28806), .Z(n25727) );
  NOR U26444 ( .A(n28807), .B(n28805), .Z(n28806) );
  XOR U26445 ( .A(n28808), .B(n28809), .Z(n25967) );
  NOR U26446 ( .A(n28810), .B(n28808), .Z(n28809) );
  XOR U26447 ( .A(n28811), .B(n28812), .Z(n25968) );
  NOR U26448 ( .A(n28813), .B(n28811), .Z(n28812) );
  XOR U26449 ( .A(n28814), .B(n28815), .Z(n25969) );
  NOR U26450 ( .A(n28816), .B(n28814), .Z(n28815) );
  XOR U26451 ( .A(n28817), .B(n28818), .Z(n25720) );
  NOR U26452 ( .A(n28819), .B(n28817), .Z(n28818) );
  XOR U26453 ( .A(n28820), .B(n28821), .Z(n25714) );
  NOR U26454 ( .A(n28822), .B(n28820), .Z(n28821) );
  XOR U26455 ( .A(n28823), .B(n28824), .Z(n25711) );
  NOR U26456 ( .A(n28825), .B(n28823), .Z(n28824) );
  XOR U26457 ( .A(n28826), .B(n28827), .Z(n25709) );
  NOR U26458 ( .A(n28828), .B(n28826), .Z(n28827) );
  XOR U26459 ( .A(n28829), .B(n28830), .Z(n25710) );
  NOR U26460 ( .A(n28831), .B(n28829), .Z(n28830) );
  XOR U26461 ( .A(n28832), .B(n28833), .Z(n25988) );
  NOR U26462 ( .A(n28834), .B(n28832), .Z(n28833) );
  XOR U26463 ( .A(n28835), .B(n28836), .Z(n25992) );
  NOR U26464 ( .A(n28837), .B(n28835), .Z(n28836) );
  XOR U26465 ( .A(n28838), .B(n28839), .Z(n25699) );
  NOR U26466 ( .A(n28840), .B(n28838), .Z(n28839) );
  XOR U26467 ( .A(n28841), .B(n28842), .Z(n25700) );
  NOR U26468 ( .A(n28843), .B(n28841), .Z(n28842) );
  XOR U26469 ( .A(n28844), .B(n28845), .Z(n26000) );
  NOR U26470 ( .A(n28846), .B(n28844), .Z(n28845) );
  XOR U26471 ( .A(n28847), .B(n28848), .Z(n26001) );
  NOR U26472 ( .A(n28849), .B(n28847), .Z(n28848) );
  XOR U26473 ( .A(n28850), .B(n28851), .Z(n26002) );
  NOR U26474 ( .A(n28852), .B(n28850), .Z(n28851) );
  XOR U26475 ( .A(n28853), .B(n28854), .Z(n25693) );
  NOR U26476 ( .A(n28855), .B(n28853), .Z(n28854) );
  XOR U26477 ( .A(n28856), .B(n28857), .Z(n25687) );
  NOR U26478 ( .A(n28858), .B(n28856), .Z(n28857) );
  XOR U26479 ( .A(n28859), .B(n28860), .Z(n25684) );
  NOR U26480 ( .A(n28861), .B(n28859), .Z(n28860) );
  XOR U26481 ( .A(n28862), .B(n28863), .Z(n25682) );
  NOR U26482 ( .A(n28864), .B(n28862), .Z(n28863) );
  XOR U26483 ( .A(n28865), .B(n28866), .Z(n25683) );
  NOR U26484 ( .A(n28867), .B(n28865), .Z(n28866) );
  XOR U26485 ( .A(n28868), .B(n28869), .Z(n26021) );
  NOR U26486 ( .A(n28870), .B(n28868), .Z(n28869) );
  XOR U26487 ( .A(n28871), .B(n28872), .Z(n26025) );
  NOR U26488 ( .A(n28873), .B(n28871), .Z(n28872) );
  XOR U26489 ( .A(n28874), .B(n28875), .Z(n25672) );
  NOR U26490 ( .A(n28876), .B(n28874), .Z(n28875) );
  XOR U26491 ( .A(n28877), .B(n28878), .Z(n25673) );
  NOR U26492 ( .A(n28879), .B(n28877), .Z(n28878) );
  XOR U26493 ( .A(n28880), .B(n28881), .Z(n26033) );
  NOR U26494 ( .A(n28882), .B(n28880), .Z(n28881) );
  XOR U26495 ( .A(n28883), .B(n28884), .Z(n26034) );
  NOR U26496 ( .A(n28885), .B(n28883), .Z(n28884) );
  XOR U26497 ( .A(n28886), .B(n28887), .Z(n26035) );
  NOR U26498 ( .A(n28888), .B(n28886), .Z(n28887) );
  XOR U26499 ( .A(n28889), .B(n28890), .Z(n25666) );
  NOR U26500 ( .A(n28891), .B(n28889), .Z(n28890) );
  XOR U26501 ( .A(n28892), .B(n28893), .Z(n25660) );
  NOR U26502 ( .A(n28894), .B(n28892), .Z(n28893) );
  XOR U26503 ( .A(n28895), .B(n28896), .Z(n25657) );
  NOR U26504 ( .A(n28897), .B(n28895), .Z(n28896) );
  XOR U26505 ( .A(n28898), .B(n28899), .Z(n25655) );
  NOR U26506 ( .A(n28900), .B(n28898), .Z(n28899) );
  XOR U26507 ( .A(n28901), .B(n28902), .Z(n25656) );
  NOR U26508 ( .A(n28903), .B(n28901), .Z(n28902) );
  XOR U26509 ( .A(n28904), .B(n28905), .Z(n26054) );
  NOR U26510 ( .A(n28906), .B(n28904), .Z(n28905) );
  XOR U26511 ( .A(n28907), .B(n28908), .Z(n26058) );
  NOR U26512 ( .A(n28909), .B(n28907), .Z(n28908) );
  XOR U26513 ( .A(n28910), .B(n28911), .Z(n25645) );
  NOR U26514 ( .A(n28912), .B(n28910), .Z(n28911) );
  XOR U26515 ( .A(n28913), .B(n28914), .Z(n25646) );
  NOR U26516 ( .A(n28915), .B(n28913), .Z(n28914) );
  XOR U26517 ( .A(n28916), .B(n28917), .Z(n26066) );
  NOR U26518 ( .A(n28918), .B(n28916), .Z(n28917) );
  XOR U26519 ( .A(n28919), .B(n28920), .Z(n26067) );
  NOR U26520 ( .A(n28921), .B(n28919), .Z(n28920) );
  XOR U26521 ( .A(n28922), .B(n28923), .Z(n26068) );
  NOR U26522 ( .A(n28924), .B(n28922), .Z(n28923) );
  XOR U26523 ( .A(n28925), .B(n28926), .Z(n25639) );
  NOR U26524 ( .A(n28927), .B(n28925), .Z(n28926) );
  XOR U26525 ( .A(n28928), .B(n28929), .Z(n25633) );
  NOR U26526 ( .A(n28930), .B(n28928), .Z(n28929) );
  XOR U26527 ( .A(n28931), .B(n28932), .Z(n25630) );
  NOR U26528 ( .A(n28933), .B(n28931), .Z(n28932) );
  XOR U26529 ( .A(n28934), .B(n28935), .Z(n25628) );
  NOR U26530 ( .A(n28936), .B(n28934), .Z(n28935) );
  XOR U26531 ( .A(n28937), .B(n28938), .Z(n25629) );
  NOR U26532 ( .A(n28939), .B(n28937), .Z(n28938) );
  XOR U26533 ( .A(n28940), .B(n28941), .Z(n26087) );
  NOR U26534 ( .A(n28942), .B(n28940), .Z(n28941) );
  XOR U26535 ( .A(n28943), .B(n28944), .Z(n26091) );
  NOR U26536 ( .A(n28945), .B(n28943), .Z(n28944) );
  XOR U26537 ( .A(n28946), .B(n28947), .Z(n25618) );
  NOR U26538 ( .A(n28948), .B(n28946), .Z(n28947) );
  XOR U26539 ( .A(n28949), .B(n28950), .Z(n25619) );
  NOR U26540 ( .A(n28951), .B(n28949), .Z(n28950) );
  XOR U26541 ( .A(n28952), .B(n28953), .Z(n26099) );
  NOR U26542 ( .A(n28954), .B(n28952), .Z(n28953) );
  XOR U26543 ( .A(n28955), .B(n28956), .Z(n26100) );
  NOR U26544 ( .A(n28957), .B(n28955), .Z(n28956) );
  XOR U26545 ( .A(n28958), .B(n28959), .Z(n26101) );
  NOR U26546 ( .A(n28960), .B(n28958), .Z(n28959) );
  XOR U26547 ( .A(n28961), .B(n28962), .Z(n25612) );
  NOR U26548 ( .A(n28963), .B(n28961), .Z(n28962) );
  XOR U26549 ( .A(n28964), .B(n28965), .Z(n25606) );
  NOR U26550 ( .A(n28966), .B(n28964), .Z(n28965) );
  XOR U26551 ( .A(n28967), .B(n28968), .Z(n25603) );
  NOR U26552 ( .A(n28969), .B(n28967), .Z(n28968) );
  XOR U26553 ( .A(n28970), .B(n28971), .Z(n25601) );
  NOR U26554 ( .A(n28972), .B(n28970), .Z(n28971) );
  XOR U26555 ( .A(n28973), .B(n28974), .Z(n25602) );
  NOR U26556 ( .A(n28975), .B(n28973), .Z(n28974) );
  XOR U26557 ( .A(n28976), .B(n28977), .Z(n26120) );
  NOR U26558 ( .A(n28978), .B(n28976), .Z(n28977) );
  XOR U26559 ( .A(n28979), .B(n28980), .Z(n26124) );
  NOR U26560 ( .A(n28981), .B(n28979), .Z(n28980) );
  XOR U26561 ( .A(n28982), .B(n28983), .Z(n25591) );
  NOR U26562 ( .A(n28984), .B(n28982), .Z(n28983) );
  XOR U26563 ( .A(n28985), .B(n28986), .Z(n25592) );
  NOR U26564 ( .A(n28987), .B(n28985), .Z(n28986) );
  XOR U26565 ( .A(n28988), .B(n28989), .Z(n26132) );
  NOR U26566 ( .A(n28990), .B(n28988), .Z(n28989) );
  XOR U26567 ( .A(n28991), .B(n28992), .Z(n26133) );
  NOR U26568 ( .A(n28993), .B(n28991), .Z(n28992) );
  XOR U26569 ( .A(n28994), .B(n28995), .Z(n26134) );
  NOR U26570 ( .A(n28996), .B(n28994), .Z(n28995) );
  XOR U26571 ( .A(n28997), .B(n28998), .Z(n25585) );
  NOR U26572 ( .A(n28999), .B(n28997), .Z(n28998) );
  XOR U26573 ( .A(n29000), .B(n29001), .Z(n25579) );
  NOR U26574 ( .A(n29002), .B(n29000), .Z(n29001) );
  XOR U26575 ( .A(n29003), .B(n29004), .Z(n25576) );
  NOR U26576 ( .A(n29005), .B(n29003), .Z(n29004) );
  XOR U26577 ( .A(n29006), .B(n29007), .Z(n25574) );
  NOR U26578 ( .A(n29008), .B(n29006), .Z(n29007) );
  XOR U26579 ( .A(n29009), .B(n29010), .Z(n25575) );
  NOR U26580 ( .A(n29011), .B(n29009), .Z(n29010) );
  XOR U26581 ( .A(n29012), .B(n29013), .Z(n26153) );
  NOR U26582 ( .A(n29014), .B(n29012), .Z(n29013) );
  XOR U26583 ( .A(n29015), .B(n29016), .Z(n26157) );
  NOR U26584 ( .A(n29017), .B(n29015), .Z(n29016) );
  XOR U26585 ( .A(n29018), .B(n29019), .Z(n25564) );
  NOR U26586 ( .A(n29020), .B(n29018), .Z(n29019) );
  XOR U26587 ( .A(n29021), .B(n29022), .Z(n25565) );
  NOR U26588 ( .A(n29023), .B(n29021), .Z(n29022) );
  XOR U26589 ( .A(n29024), .B(n29025), .Z(n26165) );
  NOR U26590 ( .A(n29026), .B(n29024), .Z(n29025) );
  XOR U26591 ( .A(n29027), .B(n29028), .Z(n26166) );
  NOR U26592 ( .A(n29029), .B(n29027), .Z(n29028) );
  XOR U26593 ( .A(n29030), .B(n29031), .Z(n26167) );
  NOR U26594 ( .A(n29032), .B(n29030), .Z(n29031) );
  XOR U26595 ( .A(n29033), .B(n29034), .Z(n25558) );
  NOR U26596 ( .A(n29035), .B(n29033), .Z(n29034) );
  XOR U26597 ( .A(n29036), .B(n29037), .Z(n25551) );
  NOR U26598 ( .A(n29038), .B(n29036), .Z(n29037) );
  XOR U26599 ( .A(n29039), .B(n29040), .Z(n25547) );
  NOR U26600 ( .A(n29041), .B(n29039), .Z(n29040) );
  XOR U26601 ( .A(n29042), .B(n29043), .Z(n25549) );
  NOR U26602 ( .A(n29044), .B(n29042), .Z(n29043) );
  XOR U26603 ( .A(n29045), .B(n29046), .Z(n26181) );
  NOR U26604 ( .A(n29047), .B(n29045), .Z(n29046) );
  XOR U26605 ( .A(n29048), .B(n29049), .Z(n26182) );
  NOR U26606 ( .A(n29050), .B(n29048), .Z(n29049) );
  XOR U26607 ( .A(n29051), .B(n29052), .Z(n26185) );
  NOR U26608 ( .A(n29053), .B(n29051), .Z(n29052) );
  XOR U26609 ( .A(n29054), .B(n29055), .Z(n26188) );
  NOR U26610 ( .A(n29056), .B(n29054), .Z(n29055) );
  XOR U26611 ( .A(n29057), .B(n29058), .Z(n26191) );
  NOR U26612 ( .A(n29059), .B(n29057), .Z(n29058) );
  XOR U26613 ( .A(n29060), .B(n29061), .Z(n26194) );
  NOR U26614 ( .A(n29062), .B(n29060), .Z(n29061) );
  XOR U26615 ( .A(n29063), .B(n29064), .Z(n26197) );
  NOR U26616 ( .A(n29065), .B(n29063), .Z(n29064) );
  XOR U26617 ( .A(n29066), .B(n29067), .Z(n26200) );
  NOR U26618 ( .A(n29068), .B(n29066), .Z(n29067) );
  XOR U26619 ( .A(n29069), .B(n29070), .Z(n26203) );
  NOR U26620 ( .A(n29071), .B(n29069), .Z(n29070) );
  XOR U26621 ( .A(n29072), .B(n29073), .Z(n26206) );
  NOR U26622 ( .A(n29074), .B(n29072), .Z(n29073) );
  XOR U26623 ( .A(n29075), .B(n29076), .Z(n26209) );
  NOR U26624 ( .A(n29077), .B(n29075), .Z(n29076) );
  XOR U26625 ( .A(n29078), .B(n29079), .Z(n26212) );
  NOR U26626 ( .A(n29080), .B(n29078), .Z(n29079) );
  XOR U26627 ( .A(n29081), .B(n29082), .Z(n26215) );
  NOR U26628 ( .A(n29083), .B(n29081), .Z(n29082) );
  XOR U26629 ( .A(n29084), .B(n29085), .Z(n26218) );
  NOR U26630 ( .A(n29086), .B(n29084), .Z(n29085) );
  XOR U26631 ( .A(n29087), .B(n29088), .Z(n26221) );
  NOR U26632 ( .A(n29089), .B(n29087), .Z(n29088) );
  XOR U26633 ( .A(n29090), .B(n29091), .Z(n26224) );
  NOR U26634 ( .A(n29092), .B(n29090), .Z(n29091) );
  XOR U26635 ( .A(n29093), .B(n29094), .Z(n26227) );
  NOR U26636 ( .A(n29095), .B(n29093), .Z(n29094) );
  XOR U26637 ( .A(n29096), .B(n29097), .Z(n26230) );
  NOR U26638 ( .A(n29098), .B(n29096), .Z(n29097) );
  XOR U26639 ( .A(n29099), .B(n29100), .Z(n26233) );
  NOR U26640 ( .A(n29101), .B(n29099), .Z(n29100) );
  XOR U26641 ( .A(n29102), .B(n29103), .Z(n26236) );
  NOR U26642 ( .A(n29104), .B(n29102), .Z(n29103) );
  XOR U26643 ( .A(n29105), .B(n29106), .Z(n26239) );
  NOR U26644 ( .A(n29107), .B(n29105), .Z(n29106) );
  XOR U26645 ( .A(n29108), .B(n29109), .Z(n26242) );
  NOR U26646 ( .A(n29110), .B(n29108), .Z(n29109) );
  XOR U26647 ( .A(n29111), .B(n29112), .Z(n26245) );
  NOR U26648 ( .A(n29113), .B(n29111), .Z(n29112) );
  XOR U26649 ( .A(n29114), .B(n29115), .Z(n26248) );
  NOR U26650 ( .A(n29116), .B(n29114), .Z(n29115) );
  XOR U26651 ( .A(n29117), .B(n29118), .Z(n26251) );
  NOR U26652 ( .A(n29119), .B(n29117), .Z(n29118) );
  XOR U26653 ( .A(n29120), .B(n29121), .Z(n26254) );
  NOR U26654 ( .A(n29122), .B(n29120), .Z(n29121) );
  XOR U26655 ( .A(n29123), .B(n29124), .Z(n26257) );
  NOR U26656 ( .A(n29125), .B(n29123), .Z(n29124) );
  XOR U26657 ( .A(n29126), .B(n29127), .Z(n26260) );
  NOR U26658 ( .A(n29128), .B(n29126), .Z(n29127) );
  XOR U26659 ( .A(n29129), .B(n29130), .Z(n26263) );
  NOR U26660 ( .A(n29131), .B(n29129), .Z(n29130) );
  XOR U26661 ( .A(n29132), .B(n29133), .Z(n26266) );
  NOR U26662 ( .A(n29134), .B(n29132), .Z(n29133) );
  XOR U26663 ( .A(n29135), .B(n29136), .Z(n26269) );
  NOR U26664 ( .A(n29137), .B(n29135), .Z(n29136) );
  XOR U26665 ( .A(n29138), .B(n29139), .Z(n26272) );
  NOR U26666 ( .A(n29140), .B(n29138), .Z(n29139) );
  XOR U26667 ( .A(n29141), .B(n29142), .Z(n26275) );
  NOR U26668 ( .A(n29143), .B(n29141), .Z(n29142) );
  XOR U26669 ( .A(n29144), .B(n29145), .Z(n26278) );
  NOR U26670 ( .A(n29146), .B(n29144), .Z(n29145) );
  XOR U26671 ( .A(n29147), .B(n29148), .Z(n26281) );
  NOR U26672 ( .A(n29149), .B(n29147), .Z(n29148) );
  XOR U26673 ( .A(n29150), .B(n29151), .Z(n26284) );
  NOR U26674 ( .A(n29152), .B(n29150), .Z(n29151) );
  XOR U26675 ( .A(n29153), .B(n29154), .Z(n26287) );
  NOR U26676 ( .A(n29155), .B(n29153), .Z(n29154) );
  XOR U26677 ( .A(n29156), .B(n29157), .Z(n26290) );
  NOR U26678 ( .A(n29158), .B(n29156), .Z(n29157) );
  XOR U26679 ( .A(n29159), .B(n29160), .Z(n26293) );
  NOR U26680 ( .A(n29161), .B(n29159), .Z(n29160) );
  XOR U26681 ( .A(n29162), .B(n29163), .Z(n26296) );
  NOR U26682 ( .A(n29164), .B(n29162), .Z(n29163) );
  XOR U26683 ( .A(n29165), .B(n29166), .Z(n26299) );
  NOR U26684 ( .A(n29167), .B(n29165), .Z(n29166) );
  XOR U26685 ( .A(n29168), .B(n29169), .Z(n26302) );
  NOR U26686 ( .A(n29170), .B(n29168), .Z(n29169) );
  XOR U26687 ( .A(n29171), .B(n29172), .Z(n26305) );
  NOR U26688 ( .A(n29173), .B(n29171), .Z(n29172) );
  XOR U26689 ( .A(n29174), .B(n29175), .Z(n26308) );
  NOR U26690 ( .A(n29176), .B(n29174), .Z(n29175) );
  XOR U26691 ( .A(n29177), .B(n29178), .Z(n26311) );
  NOR U26692 ( .A(n29179), .B(n29177), .Z(n29178) );
  XOR U26693 ( .A(n29180), .B(n29181), .Z(n26314) );
  NOR U26694 ( .A(n29182), .B(n29180), .Z(n29181) );
  XOR U26695 ( .A(n29183), .B(n29184), .Z(n26317) );
  NOR U26696 ( .A(n29185), .B(n29183), .Z(n29184) );
  XOR U26697 ( .A(n29186), .B(n29187), .Z(n26320) );
  NOR U26698 ( .A(n29188), .B(n29186), .Z(n29187) );
  XOR U26699 ( .A(n29189), .B(n29190), .Z(n26323) );
  NOR U26700 ( .A(n29191), .B(n29189), .Z(n29190) );
  XOR U26701 ( .A(n29192), .B(n29193), .Z(n26326) );
  NOR U26702 ( .A(n29194), .B(n29192), .Z(n29193) );
  XOR U26703 ( .A(n29195), .B(n29196), .Z(n26329) );
  NOR U26704 ( .A(n29197), .B(n29195), .Z(n29196) );
  XOR U26705 ( .A(n29198), .B(n29199), .Z(n26332) );
  NOR U26706 ( .A(n29200), .B(n29198), .Z(n29199) );
  XOR U26707 ( .A(n29201), .B(n29202), .Z(n26335) );
  NOR U26708 ( .A(n29203), .B(n29201), .Z(n29202) );
  XOR U26709 ( .A(n29204), .B(n29205), .Z(n26338) );
  NOR U26710 ( .A(n29206), .B(n29204), .Z(n29205) );
  XOR U26711 ( .A(n29207), .B(n29208), .Z(n26341) );
  NOR U26712 ( .A(n29209), .B(n29207), .Z(n29208) );
  XOR U26713 ( .A(n29210), .B(n29211), .Z(n26344) );
  NOR U26714 ( .A(n29212), .B(n29210), .Z(n29211) );
  XOR U26715 ( .A(n29213), .B(n29214), .Z(n26347) );
  NOR U26716 ( .A(n29215), .B(n29213), .Z(n29214) );
  XOR U26717 ( .A(n29216), .B(n29217), .Z(n26350) );
  NOR U26718 ( .A(n29218), .B(n29216), .Z(n29217) );
  XOR U26719 ( .A(n29219), .B(n29220), .Z(n26353) );
  NOR U26720 ( .A(n29221), .B(n29219), .Z(n29220) );
  XOR U26721 ( .A(n29222), .B(n29223), .Z(n26356) );
  NOR U26722 ( .A(n29224), .B(n29222), .Z(n29223) );
  XOR U26723 ( .A(n29225), .B(n29226), .Z(n26359) );
  NOR U26724 ( .A(n29227), .B(n29225), .Z(n29226) );
  XOR U26725 ( .A(n29228), .B(n29229), .Z(n26362) );
  NOR U26726 ( .A(n29230), .B(n29228), .Z(n29229) );
  XOR U26727 ( .A(n29231), .B(n29232), .Z(n26365) );
  NOR U26728 ( .A(n29233), .B(n29231), .Z(n29232) );
  XOR U26729 ( .A(n29234), .B(n29235), .Z(n26368) );
  NOR U26730 ( .A(n29236), .B(n29234), .Z(n29235) );
  XOR U26731 ( .A(n29237), .B(n29238), .Z(n26371) );
  NOR U26732 ( .A(n29239), .B(n29237), .Z(n29238) );
  XOR U26733 ( .A(n29240), .B(n29241), .Z(n26374) );
  NOR U26734 ( .A(n29242), .B(n29240), .Z(n29241) );
  XOR U26735 ( .A(n29243), .B(n29244), .Z(n26377) );
  NOR U26736 ( .A(n29245), .B(n29243), .Z(n29244) );
  XOR U26737 ( .A(n29246), .B(n29247), .Z(n26380) );
  NOR U26738 ( .A(n29248), .B(n29246), .Z(n29247) );
  XOR U26739 ( .A(n29249), .B(n29250), .Z(n26383) );
  NOR U26740 ( .A(n29251), .B(n29249), .Z(n29250) );
  XOR U26741 ( .A(n29252), .B(n29253), .Z(n26386) );
  NOR U26742 ( .A(n29254), .B(n29252), .Z(n29253) );
  XOR U26743 ( .A(n29255), .B(n29256), .Z(n26389) );
  NOR U26744 ( .A(n29257), .B(n29255), .Z(n29256) );
  XOR U26745 ( .A(n29258), .B(n29259), .Z(n26392) );
  NOR U26746 ( .A(n29260), .B(n29258), .Z(n29259) );
  XOR U26747 ( .A(n29261), .B(n29262), .Z(n26395) );
  NOR U26748 ( .A(n29263), .B(n29261), .Z(n29262) );
  XOR U26749 ( .A(n29264), .B(n29265), .Z(n26398) );
  NOR U26750 ( .A(n29266), .B(n29264), .Z(n29265) );
  XOR U26751 ( .A(n29267), .B(n29268), .Z(n26401) );
  NOR U26752 ( .A(n29269), .B(n29267), .Z(n29268) );
  XOR U26753 ( .A(n29270), .B(n29271), .Z(n26404) );
  NOR U26754 ( .A(n29272), .B(n29270), .Z(n29271) );
  XOR U26755 ( .A(n29273), .B(n29274), .Z(n26407) );
  NOR U26756 ( .A(n29275), .B(n29273), .Z(n29274) );
  XOR U26757 ( .A(n29276), .B(n29277), .Z(n26410) );
  NOR U26758 ( .A(n29278), .B(n29276), .Z(n29277) );
  XOR U26759 ( .A(n29279), .B(n29280), .Z(n26413) );
  NOR U26760 ( .A(n29281), .B(n29279), .Z(n29280) );
  XOR U26761 ( .A(n29282), .B(n29283), .Z(n26416) );
  NOR U26762 ( .A(n29284), .B(n29282), .Z(n29283) );
  XOR U26763 ( .A(n29285), .B(n29286), .Z(n26419) );
  NOR U26764 ( .A(n29287), .B(n29285), .Z(n29286) );
  XOR U26765 ( .A(n29288), .B(n29289), .Z(n26422) );
  NOR U26766 ( .A(n29290), .B(n29288), .Z(n29289) );
  XOR U26767 ( .A(n29291), .B(n29292), .Z(n26425) );
  NOR U26768 ( .A(n29293), .B(n29291), .Z(n29292) );
  XOR U26769 ( .A(n29294), .B(n29295), .Z(n26428) );
  NOR U26770 ( .A(n29296), .B(n29294), .Z(n29295) );
  XOR U26771 ( .A(n29297), .B(n29298), .Z(n26431) );
  NOR U26772 ( .A(n29299), .B(n29297), .Z(n29298) );
  XOR U26773 ( .A(n29300), .B(n29301), .Z(n26434) );
  NOR U26774 ( .A(n29302), .B(n29300), .Z(n29301) );
  XOR U26775 ( .A(n29303), .B(n29304), .Z(n26437) );
  NOR U26776 ( .A(n29305), .B(n29303), .Z(n29304) );
  XOR U26777 ( .A(n29306), .B(n29307), .Z(n26440) );
  NOR U26778 ( .A(n29308), .B(n29306), .Z(n29307) );
  XOR U26779 ( .A(n29309), .B(n29310), .Z(n26443) );
  NOR U26780 ( .A(n29311), .B(n29309), .Z(n29310) );
  XOR U26781 ( .A(n29312), .B(n29313), .Z(n26446) );
  NOR U26782 ( .A(n29314), .B(n29312), .Z(n29313) );
  XOR U26783 ( .A(n29315), .B(n29316), .Z(n26449) );
  NOR U26784 ( .A(n29317), .B(n29315), .Z(n29316) );
  XOR U26785 ( .A(n29318), .B(n29319), .Z(n26452) );
  NOR U26786 ( .A(n29320), .B(n29318), .Z(n29319) );
  XOR U26787 ( .A(n29321), .B(n29322), .Z(n26455) );
  NOR U26788 ( .A(n29323), .B(n29321), .Z(n29322) );
  XOR U26789 ( .A(n29324), .B(n29325), .Z(n26458) );
  NOR U26790 ( .A(n29326), .B(n29324), .Z(n29325) );
  XOR U26791 ( .A(n29327), .B(n29328), .Z(n26461) );
  NOR U26792 ( .A(n29329), .B(n29327), .Z(n29328) );
  XOR U26793 ( .A(n29330), .B(n29331), .Z(n26464) );
  NOR U26794 ( .A(n29332), .B(n29330), .Z(n29331) );
  XOR U26795 ( .A(n29333), .B(n29334), .Z(n26467) );
  NOR U26796 ( .A(n29335), .B(n29333), .Z(n29334) );
  XOR U26797 ( .A(n29336), .B(n29337), .Z(n26470) );
  NOR U26798 ( .A(n29338), .B(n29336), .Z(n29337) );
  XOR U26799 ( .A(n29339), .B(n29340), .Z(n26473) );
  NOR U26800 ( .A(n29341), .B(n29339), .Z(n29340) );
  XOR U26801 ( .A(n29342), .B(n29343), .Z(n26476) );
  NOR U26802 ( .A(n29344), .B(n29342), .Z(n29343) );
  XOR U26803 ( .A(n29345), .B(n29346), .Z(n26479) );
  NOR U26804 ( .A(n29347), .B(n29345), .Z(n29346) );
  XOR U26805 ( .A(n29348), .B(n29349), .Z(n26482) );
  NOR U26806 ( .A(n29350), .B(n29348), .Z(n29349) );
  XOR U26807 ( .A(n29351), .B(n29352), .Z(n26485) );
  NOR U26808 ( .A(n29353), .B(n29351), .Z(n29352) );
  XOR U26809 ( .A(n29354), .B(n29355), .Z(n26488) );
  NOR U26810 ( .A(n29356), .B(n29354), .Z(n29355) );
  XOR U26811 ( .A(n29357), .B(n29358), .Z(n26491) );
  NOR U26812 ( .A(n29359), .B(n29357), .Z(n29358) );
  XOR U26813 ( .A(n29360), .B(n29361), .Z(n26494) );
  NOR U26814 ( .A(n29362), .B(n29360), .Z(n29361) );
  XOR U26815 ( .A(n29363), .B(n29364), .Z(n26497) );
  NOR U26816 ( .A(n29365), .B(n29363), .Z(n29364) );
  XOR U26817 ( .A(n29366), .B(n29367), .Z(n26500) );
  NOR U26818 ( .A(n29368), .B(n29366), .Z(n29367) );
  XOR U26819 ( .A(n29369), .B(n29370), .Z(n26503) );
  NOR U26820 ( .A(n29371), .B(n29369), .Z(n29370) );
  XOR U26821 ( .A(n29372), .B(n29373), .Z(n26506) );
  NOR U26822 ( .A(n29374), .B(n29372), .Z(n29373) );
  XOR U26823 ( .A(n29375), .B(n29376), .Z(n26509) );
  NOR U26824 ( .A(n29377), .B(n29375), .Z(n29376) );
  XOR U26825 ( .A(n29378), .B(n29379), .Z(n26512) );
  NOR U26826 ( .A(n29380), .B(n29378), .Z(n29379) );
  XOR U26827 ( .A(n29381), .B(n29382), .Z(n26515) );
  NOR U26828 ( .A(n29383), .B(n29381), .Z(n29382) );
  XOR U26829 ( .A(n29384), .B(n29385), .Z(n26518) );
  NOR U26830 ( .A(n29386), .B(n29384), .Z(n29385) );
  XOR U26831 ( .A(n29387), .B(n29388), .Z(n26521) );
  NOR U26832 ( .A(n29389), .B(n29387), .Z(n29388) );
  XOR U26833 ( .A(n29390), .B(n29391), .Z(n26524) );
  NOR U26834 ( .A(n29392), .B(n29390), .Z(n29391) );
  XOR U26835 ( .A(n29393), .B(n29394), .Z(n26527) );
  NOR U26836 ( .A(n29395), .B(n29393), .Z(n29394) );
  XOR U26837 ( .A(n29396), .B(n29397), .Z(n26530) );
  NOR U26838 ( .A(n29398), .B(n29396), .Z(n29397) );
  XOR U26839 ( .A(n29399), .B(n29400), .Z(n26533) );
  NOR U26840 ( .A(n29401), .B(n29399), .Z(n29400) );
  XOR U26841 ( .A(n29402), .B(n29403), .Z(n26536) );
  NOR U26842 ( .A(n29404), .B(n29402), .Z(n29403) );
  XOR U26843 ( .A(n29405), .B(n29406), .Z(n26539) );
  NOR U26844 ( .A(n29407), .B(n29405), .Z(n29406) );
  XOR U26845 ( .A(n29408), .B(n29409), .Z(n26542) );
  NOR U26846 ( .A(n29410), .B(n29408), .Z(n29409) );
  XOR U26847 ( .A(n29411), .B(n29412), .Z(n26545) );
  NOR U26848 ( .A(n29413), .B(n29411), .Z(n29412) );
  XOR U26849 ( .A(n29414), .B(n29415), .Z(n26548) );
  NOR U26850 ( .A(n29416), .B(n29414), .Z(n29415) );
  XOR U26851 ( .A(n29417), .B(n29418), .Z(n26551) );
  NOR U26852 ( .A(n29419), .B(n29417), .Z(n29418) );
  XOR U26853 ( .A(n29420), .B(n29421), .Z(n26554) );
  NOR U26854 ( .A(n29422), .B(n29420), .Z(n29421) );
  XOR U26855 ( .A(n29423), .B(n29424), .Z(n26557) );
  NOR U26856 ( .A(n29425), .B(n29423), .Z(n29424) );
  XOR U26857 ( .A(n29426), .B(n29427), .Z(n26560) );
  NOR U26858 ( .A(n29428), .B(n29426), .Z(n29427) );
  XOR U26859 ( .A(n29429), .B(n29430), .Z(n26563) );
  NOR U26860 ( .A(n29431), .B(n29429), .Z(n29430) );
  XOR U26861 ( .A(n29432), .B(n29433), .Z(n26566) );
  NOR U26862 ( .A(n29434), .B(n29432), .Z(n29433) );
  XOR U26863 ( .A(n29435), .B(n29436), .Z(n26569) );
  NOR U26864 ( .A(n29437), .B(n29435), .Z(n29436) );
  XOR U26865 ( .A(n29438), .B(n29439), .Z(n26572) );
  NOR U26866 ( .A(n29440), .B(n29438), .Z(n29439) );
  XOR U26867 ( .A(n29441), .B(n29442), .Z(n26575) );
  NOR U26868 ( .A(n29443), .B(n29441), .Z(n29442) );
  XOR U26869 ( .A(n29444), .B(n29445), .Z(n26578) );
  NOR U26870 ( .A(n29446), .B(n29444), .Z(n29445) );
  XOR U26871 ( .A(n29447), .B(n29448), .Z(n26581) );
  NOR U26872 ( .A(n29449), .B(n29447), .Z(n29448) );
  XOR U26873 ( .A(n29450), .B(n29451), .Z(n26584) );
  NOR U26874 ( .A(n29452), .B(n29450), .Z(n29451) );
  XOR U26875 ( .A(n29453), .B(n29454), .Z(n26587) );
  NOR U26876 ( .A(n29455), .B(n29453), .Z(n29454) );
  XOR U26877 ( .A(n29456), .B(n29457), .Z(n26590) );
  NOR U26878 ( .A(n29458), .B(n29456), .Z(n29457) );
  XOR U26879 ( .A(n29459), .B(n29460), .Z(n26593) );
  NOR U26880 ( .A(n29461), .B(n29459), .Z(n29460) );
  XOR U26881 ( .A(n29462), .B(n29463), .Z(n26596) );
  NOR U26882 ( .A(n29464), .B(n29462), .Z(n29463) );
  XOR U26883 ( .A(n29465), .B(n29466), .Z(n26599) );
  NOR U26884 ( .A(n29467), .B(n29465), .Z(n29466) );
  XOR U26885 ( .A(n29468), .B(n29469), .Z(n26602) );
  NOR U26886 ( .A(n29470), .B(n29468), .Z(n29469) );
  XOR U26887 ( .A(n29471), .B(n29472), .Z(n26605) );
  NOR U26888 ( .A(n29473), .B(n29471), .Z(n29472) );
  XOR U26889 ( .A(n29474), .B(n29475), .Z(n26608) );
  NOR U26890 ( .A(n29476), .B(n29474), .Z(n29475) );
  XOR U26891 ( .A(n29477), .B(n29478), .Z(n26611) );
  NOR U26892 ( .A(n29479), .B(n29477), .Z(n29478) );
  XOR U26893 ( .A(n29480), .B(n29481), .Z(n26614) );
  NOR U26894 ( .A(n29482), .B(n29480), .Z(n29481) );
  XOR U26895 ( .A(n29483), .B(n29484), .Z(n26617) );
  NOR U26896 ( .A(n29485), .B(n29483), .Z(n29484) );
  XOR U26897 ( .A(n29486), .B(n29487), .Z(n26620) );
  NOR U26898 ( .A(n29488), .B(n29486), .Z(n29487) );
  XOR U26899 ( .A(n29489), .B(n29490), .Z(n26623) );
  NOR U26900 ( .A(n29491), .B(n29489), .Z(n29490) );
  XOR U26901 ( .A(n29492), .B(n29493), .Z(n26626) );
  NOR U26902 ( .A(n29494), .B(n29492), .Z(n29493) );
  XOR U26903 ( .A(n29495), .B(n29496), .Z(n26629) );
  NOR U26904 ( .A(n29497), .B(n29495), .Z(n29496) );
  XOR U26905 ( .A(n29498), .B(n29499), .Z(n26632) );
  NOR U26906 ( .A(n29500), .B(n29498), .Z(n29499) );
  XOR U26907 ( .A(n29501), .B(n29502), .Z(n26635) );
  NOR U26908 ( .A(n29503), .B(n29501), .Z(n29502) );
  XOR U26909 ( .A(n29504), .B(n29505), .Z(n26638) );
  NOR U26910 ( .A(n29506), .B(n29504), .Z(n29505) );
  XOR U26911 ( .A(n29507), .B(n29508), .Z(n26641) );
  NOR U26912 ( .A(n29509), .B(n29507), .Z(n29508) );
  XOR U26913 ( .A(n29510), .B(n29511), .Z(n26644) );
  NOR U26914 ( .A(n29512), .B(n29510), .Z(n29511) );
  XOR U26915 ( .A(n29513), .B(n29514), .Z(n26647) );
  NOR U26916 ( .A(n29515), .B(n29513), .Z(n29514) );
  XOR U26917 ( .A(n29516), .B(n29517), .Z(n26650) );
  NOR U26918 ( .A(n29518), .B(n29516), .Z(n29517) );
  XOR U26919 ( .A(n29519), .B(n29520), .Z(n26653) );
  NOR U26920 ( .A(n29521), .B(n29519), .Z(n29520) );
  XOR U26921 ( .A(n29522), .B(n29523), .Z(n26656) );
  NOR U26922 ( .A(n29524), .B(n29522), .Z(n29523) );
  XOR U26923 ( .A(n29525), .B(n29526), .Z(n26659) );
  NOR U26924 ( .A(n29527), .B(n29525), .Z(n29526) );
  XOR U26925 ( .A(n29528), .B(n29529), .Z(n26662) );
  NOR U26926 ( .A(n29530), .B(n29528), .Z(n29529) );
  XOR U26927 ( .A(n29531), .B(n29532), .Z(n26665) );
  NOR U26928 ( .A(n29533), .B(n29531), .Z(n29532) );
  XOR U26929 ( .A(n29534), .B(n29535), .Z(n26668) );
  NOR U26930 ( .A(n29536), .B(n29534), .Z(n29535) );
  XOR U26931 ( .A(n29537), .B(n29538), .Z(n26671) );
  NOR U26932 ( .A(n29539), .B(n29537), .Z(n29538) );
  XOR U26933 ( .A(n29540), .B(n29541), .Z(n26674) );
  NOR U26934 ( .A(n29542), .B(n29540), .Z(n29541) );
  XOR U26935 ( .A(n29543), .B(n29544), .Z(n26677) );
  NOR U26936 ( .A(n29545), .B(n29543), .Z(n29544) );
  XOR U26937 ( .A(n29546), .B(n29547), .Z(n26680) );
  NOR U26938 ( .A(n29548), .B(n29546), .Z(n29547) );
  XOR U26939 ( .A(n29549), .B(n29550), .Z(n26683) );
  NOR U26940 ( .A(n29551), .B(n29549), .Z(n29550) );
  XOR U26941 ( .A(n29552), .B(n29553), .Z(n26686) );
  NOR U26942 ( .A(n29554), .B(n29552), .Z(n29553) );
  XOR U26943 ( .A(n29555), .B(n29556), .Z(n26689) );
  NOR U26944 ( .A(n29557), .B(n29555), .Z(n29556) );
  XOR U26945 ( .A(n29558), .B(n29559), .Z(n26692) );
  NOR U26946 ( .A(n29560), .B(n29558), .Z(n29559) );
  XOR U26947 ( .A(n29561), .B(n29562), .Z(n26695) );
  NOR U26948 ( .A(n29563), .B(n29561), .Z(n29562) );
  XOR U26949 ( .A(n29564), .B(n29565), .Z(n26698) );
  NOR U26950 ( .A(n29566), .B(n29564), .Z(n29565) );
  XOR U26951 ( .A(n29567), .B(n29568), .Z(n26701) );
  NOR U26952 ( .A(n29569), .B(n29567), .Z(n29568) );
  XOR U26953 ( .A(n29570), .B(n29571), .Z(n26704) );
  NOR U26954 ( .A(n29572), .B(n29570), .Z(n29571) );
  XOR U26955 ( .A(n29573), .B(n29574), .Z(n26707) );
  NOR U26956 ( .A(n29575), .B(n29573), .Z(n29574) );
  XOR U26957 ( .A(n29576), .B(n29577), .Z(n26710) );
  NOR U26958 ( .A(n29578), .B(n29576), .Z(n29577) );
  XOR U26959 ( .A(n29579), .B(n29580), .Z(n26713) );
  NOR U26960 ( .A(n29581), .B(n29579), .Z(n29580) );
  XOR U26961 ( .A(n29582), .B(n29583), .Z(n26716) );
  NOR U26962 ( .A(n29584), .B(n29582), .Z(n29583) );
  XOR U26963 ( .A(n29585), .B(n29586), .Z(n26719) );
  NOR U26964 ( .A(n29587), .B(n29585), .Z(n29586) );
  XOR U26965 ( .A(n29588), .B(n29589), .Z(n26722) );
  NOR U26966 ( .A(n29590), .B(n29588), .Z(n29589) );
  XOR U26967 ( .A(n29591), .B(n29592), .Z(n26725) );
  NOR U26968 ( .A(n29593), .B(n29591), .Z(n29592) );
  XOR U26969 ( .A(n29594), .B(n29595), .Z(n26728) );
  NOR U26970 ( .A(n29596), .B(n29594), .Z(n29595) );
  XOR U26971 ( .A(n29597), .B(n29598), .Z(n26731) );
  NOR U26972 ( .A(n29599), .B(n29597), .Z(n29598) );
  XOR U26973 ( .A(n29600), .B(n29601), .Z(n26734) );
  NOR U26974 ( .A(n29602), .B(n29600), .Z(n29601) );
  XOR U26975 ( .A(n29603), .B(n29604), .Z(n26737) );
  NOR U26976 ( .A(n29605), .B(n29603), .Z(n29604) );
  XOR U26977 ( .A(n29606), .B(n29607), .Z(n26740) );
  NOR U26978 ( .A(n29608), .B(n29606), .Z(n29607) );
  XOR U26979 ( .A(n29609), .B(n29610), .Z(n26743) );
  NOR U26980 ( .A(n29611), .B(n29609), .Z(n29610) );
  XOR U26981 ( .A(n29612), .B(n29613), .Z(n26746) );
  NOR U26982 ( .A(n29614), .B(n29612), .Z(n29613) );
  XOR U26983 ( .A(n29615), .B(n29616), .Z(n26749) );
  NOR U26984 ( .A(n29617), .B(n29615), .Z(n29616) );
  XOR U26985 ( .A(n29618), .B(n29619), .Z(n26752) );
  NOR U26986 ( .A(n29620), .B(n29618), .Z(n29619) );
  XOR U26987 ( .A(n29621), .B(n29622), .Z(n26755) );
  NOR U26988 ( .A(n29623), .B(n29621), .Z(n29622) );
  XOR U26989 ( .A(n29624), .B(n29625), .Z(n26758) );
  NOR U26990 ( .A(n29626), .B(n29624), .Z(n29625) );
  XOR U26991 ( .A(n29627), .B(n29628), .Z(n26761) );
  NOR U26992 ( .A(n29629), .B(n29627), .Z(n29628) );
  XOR U26993 ( .A(n29630), .B(n29631), .Z(n26764) );
  NOR U26994 ( .A(n29632), .B(n29630), .Z(n29631) );
  XOR U26995 ( .A(n29633), .B(n29634), .Z(n26767) );
  NOR U26996 ( .A(n29635), .B(n29633), .Z(n29634) );
  XOR U26997 ( .A(n29636), .B(n29637), .Z(n26770) );
  NOR U26998 ( .A(n29638), .B(n29636), .Z(n29637) );
  XOR U26999 ( .A(n29639), .B(n29640), .Z(n26773) );
  NOR U27000 ( .A(n29641), .B(n29639), .Z(n29640) );
  XOR U27001 ( .A(n29642), .B(n29643), .Z(n26776) );
  NOR U27002 ( .A(n29644), .B(n29642), .Z(n29643) );
  XOR U27003 ( .A(n29645), .B(n29646), .Z(n26779) );
  NOR U27004 ( .A(n29647), .B(n29645), .Z(n29646) );
  XOR U27005 ( .A(n29648), .B(n29649), .Z(n26782) );
  NOR U27006 ( .A(n29650), .B(n29648), .Z(n29649) );
  XOR U27007 ( .A(n29651), .B(n29652), .Z(n26785) );
  NOR U27008 ( .A(n29653), .B(n29651), .Z(n29652) );
  XOR U27009 ( .A(n29654), .B(n29655), .Z(n26788) );
  NOR U27010 ( .A(n29656), .B(n29654), .Z(n29655) );
  XOR U27011 ( .A(n29657), .B(n29658), .Z(n26791) );
  NOR U27012 ( .A(n29659), .B(n29657), .Z(n29658) );
  XOR U27013 ( .A(n29660), .B(n29661), .Z(n26794) );
  NOR U27014 ( .A(n29662), .B(n29660), .Z(n29661) );
  XOR U27015 ( .A(n29663), .B(n29664), .Z(n26797) );
  NOR U27016 ( .A(n29665), .B(n29663), .Z(n29664) );
  XOR U27017 ( .A(n29666), .B(n29667), .Z(n26800) );
  NOR U27018 ( .A(n29668), .B(n29666), .Z(n29667) );
  XOR U27019 ( .A(n29669), .B(n29670), .Z(n26803) );
  NOR U27020 ( .A(n29671), .B(n29669), .Z(n29670) );
  XOR U27021 ( .A(n29672), .B(n29673), .Z(n26806) );
  NOR U27022 ( .A(n29674), .B(n29672), .Z(n29673) );
  XOR U27023 ( .A(n29675), .B(n29676), .Z(n26809) );
  NOR U27024 ( .A(n29677), .B(n29675), .Z(n29676) );
  XOR U27025 ( .A(n29678), .B(n29679), .Z(n26812) );
  NOR U27026 ( .A(n29680), .B(n29678), .Z(n29679) );
  XOR U27027 ( .A(n29681), .B(n29682), .Z(n26815) );
  NOR U27028 ( .A(n29683), .B(n29681), .Z(n29682) );
  XOR U27029 ( .A(n29684), .B(n29685), .Z(n26818) );
  NOR U27030 ( .A(n29686), .B(n29684), .Z(n29685) );
  XOR U27031 ( .A(n29687), .B(n29688), .Z(n26821) );
  NOR U27032 ( .A(n29689), .B(n29687), .Z(n29688) );
  XOR U27033 ( .A(n29690), .B(n29691), .Z(n26824) );
  NOR U27034 ( .A(n29692), .B(n29690), .Z(n29691) );
  XOR U27035 ( .A(n29693), .B(n29694), .Z(n26827) );
  NOR U27036 ( .A(n29695), .B(n29693), .Z(n29694) );
  XOR U27037 ( .A(n29696), .B(n29697), .Z(n26830) );
  NOR U27038 ( .A(n29698), .B(n29696), .Z(n29697) );
  XOR U27039 ( .A(n29699), .B(n29700), .Z(n26833) );
  NOR U27040 ( .A(n29701), .B(n29699), .Z(n29700) );
  XOR U27041 ( .A(n29702), .B(n29703), .Z(n26836) );
  NOR U27042 ( .A(n29704), .B(n29702), .Z(n29703) );
  XOR U27043 ( .A(n29705), .B(n29706), .Z(n26839) );
  NOR U27044 ( .A(n29707), .B(n29705), .Z(n29706) );
  XOR U27045 ( .A(n29708), .B(n29709), .Z(n26842) );
  NOR U27046 ( .A(n29710), .B(n29708), .Z(n29709) );
  XOR U27047 ( .A(n29711), .B(n29712), .Z(n26845) );
  NOR U27048 ( .A(n29713), .B(n29711), .Z(n29712) );
  XOR U27049 ( .A(n29714), .B(n29715), .Z(n26848) );
  NOR U27050 ( .A(n29716), .B(n29714), .Z(n29715) );
  XOR U27051 ( .A(n29717), .B(n29718), .Z(n26851) );
  NOR U27052 ( .A(n29719), .B(n29717), .Z(n29718) );
  XOR U27053 ( .A(n29720), .B(n29721), .Z(n26854) );
  NOR U27054 ( .A(n29722), .B(n29720), .Z(n29721) );
  XOR U27055 ( .A(n29723), .B(n29724), .Z(n26857) );
  NOR U27056 ( .A(n29725), .B(n29723), .Z(n29724) );
  XOR U27057 ( .A(n29726), .B(n29727), .Z(n26860) );
  NOR U27058 ( .A(n29728), .B(n29726), .Z(n29727) );
  XOR U27059 ( .A(n29729), .B(n29730), .Z(n26863) );
  NOR U27060 ( .A(n29731), .B(n29729), .Z(n29730) );
  XOR U27061 ( .A(n29732), .B(n29733), .Z(n26866) );
  NOR U27062 ( .A(n29734), .B(n29732), .Z(n29733) );
  XOR U27063 ( .A(n29735), .B(n29736), .Z(n26869) );
  NOR U27064 ( .A(n29737), .B(n29735), .Z(n29736) );
  XOR U27065 ( .A(n29738), .B(n29739), .Z(n26872) );
  NOR U27066 ( .A(n29740), .B(n29738), .Z(n29739) );
  XOR U27067 ( .A(n29741), .B(n29742), .Z(n26875) );
  NOR U27068 ( .A(n29743), .B(n29741), .Z(n29742) );
  XOR U27069 ( .A(n29744), .B(n29745), .Z(n26878) );
  NOR U27070 ( .A(n29746), .B(n29744), .Z(n29745) );
  XOR U27071 ( .A(n29747), .B(n29748), .Z(n26881) );
  NOR U27072 ( .A(n29749), .B(n29747), .Z(n29748) );
  XOR U27073 ( .A(n29750), .B(n29751), .Z(n26884) );
  NOR U27074 ( .A(n29752), .B(n29750), .Z(n29751) );
  XOR U27075 ( .A(n29753), .B(n29754), .Z(n26887) );
  NOR U27076 ( .A(n29755), .B(n29753), .Z(n29754) );
  XOR U27077 ( .A(n29756), .B(n29757), .Z(n26890) );
  NOR U27078 ( .A(n29758), .B(n29756), .Z(n29757) );
  XOR U27079 ( .A(n29759), .B(n29760), .Z(n26893) );
  NOR U27080 ( .A(n29761), .B(n29759), .Z(n29760) );
  XOR U27081 ( .A(n29762), .B(n29763), .Z(n26896) );
  NOR U27082 ( .A(n29764), .B(n29762), .Z(n29763) );
  XOR U27083 ( .A(n29765), .B(n29766), .Z(n26899) );
  NOR U27084 ( .A(n29767), .B(n29765), .Z(n29766) );
  XOR U27085 ( .A(n29768), .B(n29769), .Z(n26902) );
  NOR U27086 ( .A(n29770), .B(n29768), .Z(n29769) );
  XOR U27087 ( .A(n29771), .B(n29772), .Z(n26905) );
  NOR U27088 ( .A(n29773), .B(n29771), .Z(n29772) );
  XOR U27089 ( .A(n29774), .B(n29775), .Z(n26908) );
  NOR U27090 ( .A(n29776), .B(n29774), .Z(n29775) );
  XOR U27091 ( .A(n29777), .B(n29778), .Z(n26911) );
  NOR U27092 ( .A(n29779), .B(n29777), .Z(n29778) );
  XOR U27093 ( .A(n29780), .B(n29781), .Z(n26914) );
  NOR U27094 ( .A(n29782), .B(n29780), .Z(n29781) );
  XOR U27095 ( .A(n29783), .B(n29784), .Z(n26917) );
  NOR U27096 ( .A(n29785), .B(n29783), .Z(n29784) );
  XOR U27097 ( .A(n29786), .B(n29787), .Z(n26920) );
  NOR U27098 ( .A(n29788), .B(n29786), .Z(n29787) );
  XOR U27099 ( .A(n29789), .B(n29790), .Z(n26923) );
  NOR U27100 ( .A(n29791), .B(n29789), .Z(n29790) );
  XOR U27101 ( .A(n29792), .B(n29793), .Z(n26926) );
  NOR U27102 ( .A(n29794), .B(n29792), .Z(n29793) );
  XOR U27103 ( .A(n29795), .B(n29796), .Z(n26929) );
  NOR U27104 ( .A(n29797), .B(n29795), .Z(n29796) );
  XOR U27105 ( .A(n29798), .B(n29799), .Z(n26932) );
  NOR U27106 ( .A(n29800), .B(n29798), .Z(n29799) );
  XOR U27107 ( .A(n29801), .B(n29802), .Z(n26935) );
  NOR U27108 ( .A(n29803), .B(n29801), .Z(n29802) );
  XOR U27109 ( .A(n29804), .B(n29805), .Z(n26938) );
  NOR U27110 ( .A(n29806), .B(n29804), .Z(n29805) );
  XOR U27111 ( .A(n29807), .B(n29808), .Z(n26941) );
  NOR U27112 ( .A(n29809), .B(n29807), .Z(n29808) );
  XOR U27113 ( .A(n29810), .B(n29811), .Z(n26944) );
  NOR U27114 ( .A(n29812), .B(n29810), .Z(n29811) );
  XOR U27115 ( .A(n29813), .B(n29814), .Z(n26947) );
  AND U27116 ( .A(n29815), .B(n29813), .Z(n29814) );
  XOR U27117 ( .A(n29816), .B(n29817), .Z(n26950) );
  AND U27118 ( .A(n79), .B(n29816), .Z(n29817) );
  XNOR U27119 ( .A(n28365), .B(n63), .Z(n28367) );
  XOR U27120 ( .A(n28363), .B(n28362), .Z(n63) );
  XNOR U27121 ( .A(n28360), .B(n28359), .Z(n28362) );
  XNOR U27122 ( .A(n28357), .B(n28356), .Z(n28359) );
  XNOR U27123 ( .A(n28354), .B(n28353), .Z(n28356) );
  XNOR U27124 ( .A(n28351), .B(n28350), .Z(n28353) );
  XNOR U27125 ( .A(n28348), .B(n28347), .Z(n28350) );
  XNOR U27126 ( .A(n28345), .B(n28344), .Z(n28347) );
  XNOR U27127 ( .A(n28342), .B(n28341), .Z(n28344) );
  XNOR U27128 ( .A(n28339), .B(n28338), .Z(n28341) );
  XNOR U27129 ( .A(n28336), .B(n28335), .Z(n28338) );
  XNOR U27130 ( .A(n28333), .B(n28332), .Z(n28335) );
  XNOR U27131 ( .A(n28330), .B(n28329), .Z(n28332) );
  XNOR U27132 ( .A(n28327), .B(n28326), .Z(n28329) );
  XNOR U27133 ( .A(n28324), .B(n28323), .Z(n28326) );
  XNOR U27134 ( .A(n28321), .B(n28320), .Z(n28323) );
  XNOR U27135 ( .A(n28318), .B(n28317), .Z(n28320) );
  XNOR U27136 ( .A(n28315), .B(n28314), .Z(n28317) );
  XNOR U27137 ( .A(n28312), .B(n28311), .Z(n28314) );
  XNOR U27138 ( .A(n28309), .B(n28308), .Z(n28311) );
  XNOR U27139 ( .A(n28306), .B(n28305), .Z(n28308) );
  XNOR U27140 ( .A(n28303), .B(n28302), .Z(n28305) );
  XNOR U27141 ( .A(n28300), .B(n28299), .Z(n28302) );
  XNOR U27142 ( .A(n28297), .B(n28296), .Z(n28299) );
  XNOR U27143 ( .A(n28294), .B(n28293), .Z(n28296) );
  XNOR U27144 ( .A(n28291), .B(n28290), .Z(n28293) );
  XNOR U27145 ( .A(n28288), .B(n28287), .Z(n28290) );
  XNOR U27146 ( .A(n28285), .B(n28284), .Z(n28287) );
  XNOR U27147 ( .A(n28282), .B(n28281), .Z(n28284) );
  XNOR U27148 ( .A(n28279), .B(n28278), .Z(n28281) );
  XNOR U27149 ( .A(n28276), .B(n28275), .Z(n28278) );
  XNOR U27150 ( .A(n28273), .B(n28272), .Z(n28275) );
  XNOR U27151 ( .A(n28270), .B(n28269), .Z(n28272) );
  XNOR U27152 ( .A(n28267), .B(n28266), .Z(n28269) );
  XNOR U27153 ( .A(n28264), .B(n28263), .Z(n28266) );
  XNOR U27154 ( .A(n28261), .B(n28260), .Z(n28263) );
  XNOR U27155 ( .A(n28258), .B(n28257), .Z(n28260) );
  XNOR U27156 ( .A(n28255), .B(n28254), .Z(n28257) );
  XNOR U27157 ( .A(n28252), .B(n28251), .Z(n28254) );
  XNOR U27158 ( .A(n28249), .B(n28248), .Z(n28251) );
  XNOR U27159 ( .A(n28246), .B(n28245), .Z(n28248) );
  XNOR U27160 ( .A(n28243), .B(n28242), .Z(n28245) );
  XNOR U27161 ( .A(n28240), .B(n28239), .Z(n28242) );
  XNOR U27162 ( .A(n28237), .B(n28236), .Z(n28239) );
  XNOR U27163 ( .A(n28234), .B(n28233), .Z(n28236) );
  XNOR U27164 ( .A(n28231), .B(n28230), .Z(n28233) );
  XNOR U27165 ( .A(n28228), .B(n28227), .Z(n28230) );
  XNOR U27166 ( .A(n28225), .B(n28224), .Z(n28227) );
  XNOR U27167 ( .A(n28222), .B(n28221), .Z(n28224) );
  XNOR U27168 ( .A(n28219), .B(n28218), .Z(n28221) );
  XNOR U27169 ( .A(n28216), .B(n28215), .Z(n28218) );
  XNOR U27170 ( .A(n28213), .B(n28212), .Z(n28215) );
  XNOR U27171 ( .A(n28210), .B(n28209), .Z(n28212) );
  XNOR U27172 ( .A(n28207), .B(n28206), .Z(n28209) );
  XNOR U27173 ( .A(n28204), .B(n28203), .Z(n28206) );
  XNOR U27174 ( .A(n28201), .B(n28200), .Z(n28203) );
  XNOR U27175 ( .A(n28198), .B(n28197), .Z(n28200) );
  XNOR U27176 ( .A(n28195), .B(n28194), .Z(n28197) );
  XNOR U27177 ( .A(n28192), .B(n28191), .Z(n28194) );
  XNOR U27178 ( .A(n28189), .B(n28188), .Z(n28191) );
  XNOR U27179 ( .A(n28186), .B(n28185), .Z(n28188) );
  XNOR U27180 ( .A(n28183), .B(n28182), .Z(n28185) );
  XNOR U27181 ( .A(n28180), .B(n28179), .Z(n28182) );
  XNOR U27182 ( .A(n28177), .B(n28176), .Z(n28179) );
  XNOR U27183 ( .A(n28174), .B(n28173), .Z(n28176) );
  XNOR U27184 ( .A(n28171), .B(n28170), .Z(n28173) );
  XNOR U27185 ( .A(n28168), .B(n28167), .Z(n28170) );
  XNOR U27186 ( .A(n28165), .B(n28164), .Z(n28167) );
  XNOR U27187 ( .A(n28162), .B(n28161), .Z(n28164) );
  XNOR U27188 ( .A(n28159), .B(n28158), .Z(n28161) );
  XNOR U27189 ( .A(n28156), .B(n28155), .Z(n28158) );
  XNOR U27190 ( .A(n28153), .B(n28152), .Z(n28155) );
  XNOR U27191 ( .A(n28150), .B(n28149), .Z(n28152) );
  XNOR U27192 ( .A(n28147), .B(n28146), .Z(n28149) );
  XNOR U27193 ( .A(n28144), .B(n28143), .Z(n28146) );
  XNOR U27194 ( .A(n28141), .B(n28140), .Z(n28143) );
  XNOR U27195 ( .A(n28138), .B(n28137), .Z(n28140) );
  XNOR U27196 ( .A(n28135), .B(n28134), .Z(n28137) );
  XNOR U27197 ( .A(n28132), .B(n28131), .Z(n28134) );
  XNOR U27198 ( .A(n28129), .B(n28128), .Z(n28131) );
  XNOR U27199 ( .A(n28126), .B(n28125), .Z(n28128) );
  XNOR U27200 ( .A(n28123), .B(n28122), .Z(n28125) );
  XNOR U27201 ( .A(n28120), .B(n28119), .Z(n28122) );
  XNOR U27202 ( .A(n28117), .B(n28116), .Z(n28119) );
  XNOR U27203 ( .A(n28114), .B(n28113), .Z(n28116) );
  XNOR U27204 ( .A(n28111), .B(n28110), .Z(n28113) );
  XNOR U27205 ( .A(n28108), .B(n28107), .Z(n28110) );
  XNOR U27206 ( .A(n28105), .B(n28104), .Z(n28107) );
  XNOR U27207 ( .A(n28102), .B(n28101), .Z(n28104) );
  XNOR U27208 ( .A(n28099), .B(n28098), .Z(n28101) );
  XNOR U27209 ( .A(n28096), .B(n28095), .Z(n28098) );
  XNOR U27210 ( .A(n28093), .B(n28092), .Z(n28095) );
  XNOR U27211 ( .A(n28090), .B(n28089), .Z(n28092) );
  XNOR U27212 ( .A(n28087), .B(n28086), .Z(n28089) );
  XNOR U27213 ( .A(n28084), .B(n28083), .Z(n28086) );
  XNOR U27214 ( .A(n28081), .B(n28080), .Z(n28083) );
  XNOR U27215 ( .A(n28078), .B(n28077), .Z(n28080) );
  XNOR U27216 ( .A(n28075), .B(n28074), .Z(n28077) );
  XNOR U27217 ( .A(n28072), .B(n28071), .Z(n28074) );
  XNOR U27218 ( .A(n28069), .B(n28068), .Z(n28071) );
  XNOR U27219 ( .A(n28066), .B(n28065), .Z(n28068) );
  XNOR U27220 ( .A(n28063), .B(n28062), .Z(n28065) );
  XNOR U27221 ( .A(n28060), .B(n28059), .Z(n28062) );
  XNOR U27222 ( .A(n28057), .B(n28056), .Z(n28059) );
  XNOR U27223 ( .A(n28054), .B(n28053), .Z(n28056) );
  XNOR U27224 ( .A(n28051), .B(n28050), .Z(n28053) );
  XNOR U27225 ( .A(n28048), .B(n28047), .Z(n28050) );
  XNOR U27226 ( .A(n28045), .B(n28044), .Z(n28047) );
  XNOR U27227 ( .A(n28042), .B(n28041), .Z(n28044) );
  XNOR U27228 ( .A(n28039), .B(n28038), .Z(n28041) );
  XNOR U27229 ( .A(n28036), .B(n28035), .Z(n28038) );
  XNOR U27230 ( .A(n28033), .B(n28032), .Z(n28035) );
  XNOR U27231 ( .A(n28030), .B(n28029), .Z(n28032) );
  XNOR U27232 ( .A(n28027), .B(n28026), .Z(n28029) );
  XNOR U27233 ( .A(n28024), .B(n28023), .Z(n28026) );
  XNOR U27234 ( .A(n28021), .B(n28020), .Z(n28023) );
  XNOR U27235 ( .A(n28018), .B(n28017), .Z(n28020) );
  XNOR U27236 ( .A(n28015), .B(n28014), .Z(n28017) );
  XNOR U27237 ( .A(n28012), .B(n28011), .Z(n28014) );
  XNOR U27238 ( .A(n28009), .B(n28008), .Z(n28011) );
  XNOR U27239 ( .A(n28006), .B(n28005), .Z(n28008) );
  XNOR U27240 ( .A(n28003), .B(n28002), .Z(n28005) );
  XNOR U27241 ( .A(n28000), .B(n27999), .Z(n28002) );
  XNOR U27242 ( .A(n27997), .B(n27996), .Z(n27999) );
  XNOR U27243 ( .A(n27994), .B(n27993), .Z(n27996) );
  XNOR U27244 ( .A(n27991), .B(n27990), .Z(n27993) );
  XNOR U27245 ( .A(n27988), .B(n27987), .Z(n27990) );
  XNOR U27246 ( .A(n27985), .B(n27984), .Z(n27987) );
  XNOR U27247 ( .A(n27982), .B(n27981), .Z(n27984) );
  XNOR U27248 ( .A(n27979), .B(n27978), .Z(n27981) );
  XNOR U27249 ( .A(n27976), .B(n27975), .Z(n27978) );
  XNOR U27250 ( .A(n27973), .B(n27972), .Z(n27975) );
  XNOR U27251 ( .A(n27970), .B(n27969), .Z(n27972) );
  XNOR U27252 ( .A(n27967), .B(n27966), .Z(n27969) );
  XNOR U27253 ( .A(n27964), .B(n27963), .Z(n27966) );
  XNOR U27254 ( .A(n27961), .B(n27960), .Z(n27963) );
  XNOR U27255 ( .A(n27958), .B(n27957), .Z(n27960) );
  XNOR U27256 ( .A(n27955), .B(n27954), .Z(n27957) );
  XNOR U27257 ( .A(n27952), .B(n27951), .Z(n27954) );
  XNOR U27258 ( .A(n27949), .B(n27948), .Z(n27951) );
  XNOR U27259 ( .A(n27946), .B(n27945), .Z(n27948) );
  XNOR U27260 ( .A(n27943), .B(n27942), .Z(n27945) );
  XNOR U27261 ( .A(n27940), .B(n27939), .Z(n27942) );
  XNOR U27262 ( .A(n27937), .B(n27936), .Z(n27939) );
  XNOR U27263 ( .A(n27934), .B(n27933), .Z(n27936) );
  XNOR U27264 ( .A(n27931), .B(n27930), .Z(n27933) );
  XNOR U27265 ( .A(n27928), .B(n27927), .Z(n27930) );
  XNOR U27266 ( .A(n27925), .B(n27924), .Z(n27927) );
  XNOR U27267 ( .A(n27922), .B(n27921), .Z(n27924) );
  XNOR U27268 ( .A(n27919), .B(n27918), .Z(n27921) );
  XNOR U27269 ( .A(n27916), .B(n27915), .Z(n27918) );
  XNOR U27270 ( .A(n27913), .B(n27912), .Z(n27915) );
  XNOR U27271 ( .A(n27910), .B(n27909), .Z(n27912) );
  XNOR U27272 ( .A(n27907), .B(n27906), .Z(n27909) );
  XNOR U27273 ( .A(n27904), .B(n27903), .Z(n27906) );
  XNOR U27274 ( .A(n27901), .B(n27900), .Z(n27903) );
  XNOR U27275 ( .A(n27898), .B(n27897), .Z(n27900) );
  XNOR U27276 ( .A(n27895), .B(n27894), .Z(n27897) );
  XNOR U27277 ( .A(n27892), .B(n27891), .Z(n27894) );
  XNOR U27278 ( .A(n27889), .B(n27888), .Z(n27891) );
  XNOR U27279 ( .A(n27886), .B(n27885), .Z(n27888) );
  XNOR U27280 ( .A(n27883), .B(n27882), .Z(n27885) );
  XNOR U27281 ( .A(n27880), .B(n27879), .Z(n27882) );
  XNOR U27282 ( .A(n27877), .B(n27876), .Z(n27879) );
  XNOR U27283 ( .A(n27874), .B(n27873), .Z(n27876) );
  XNOR U27284 ( .A(n27871), .B(n27870), .Z(n27873) );
  XNOR U27285 ( .A(n27868), .B(n27867), .Z(n27870) );
  XNOR U27286 ( .A(n27865), .B(n27864), .Z(n27867) );
  XNOR U27287 ( .A(n27862), .B(n27861), .Z(n27864) );
  XNOR U27288 ( .A(n27859), .B(n27858), .Z(n27861) );
  XNOR U27289 ( .A(n27856), .B(n27855), .Z(n27858) );
  XNOR U27290 ( .A(n27853), .B(n27852), .Z(n27855) );
  XNOR U27291 ( .A(n27850), .B(n27849), .Z(n27852) );
  XNOR U27292 ( .A(n27847), .B(n27846), .Z(n27849) );
  XNOR U27293 ( .A(n27844), .B(n27843), .Z(n27846) );
  XNOR U27294 ( .A(n27841), .B(n27840), .Z(n27843) );
  XNOR U27295 ( .A(n27838), .B(n27837), .Z(n27840) );
  XNOR U27296 ( .A(n27835), .B(n27834), .Z(n27837) );
  XNOR U27297 ( .A(n27832), .B(n27831), .Z(n27834) );
  XNOR U27298 ( .A(n27829), .B(n27828), .Z(n27831) );
  XNOR U27299 ( .A(n27826), .B(n27825), .Z(n27828) );
  XNOR U27300 ( .A(n27823), .B(n27822), .Z(n27825) );
  XNOR U27301 ( .A(n27820), .B(n27819), .Z(n27822) );
  XNOR U27302 ( .A(n27817), .B(n27816), .Z(n27819) );
  XNOR U27303 ( .A(n27814), .B(n27813), .Z(n27816) );
  XNOR U27304 ( .A(n27811), .B(n27810), .Z(n27813) );
  XNOR U27305 ( .A(n27808), .B(n27807), .Z(n27810) );
  XNOR U27306 ( .A(n27805), .B(n27804), .Z(n27807) );
  XNOR U27307 ( .A(n27802), .B(n27801), .Z(n27804) );
  XNOR U27308 ( .A(n27799), .B(n27798), .Z(n27801) );
  XNOR U27309 ( .A(n27796), .B(n27795), .Z(n27798) );
  XNOR U27310 ( .A(n27793), .B(n27792), .Z(n27795) );
  XNOR U27311 ( .A(n27790), .B(n27789), .Z(n27792) );
  XNOR U27312 ( .A(n27787), .B(n27786), .Z(n27789) );
  XNOR U27313 ( .A(n27784), .B(n27783), .Z(n27786) );
  XNOR U27314 ( .A(n27781), .B(n27780), .Z(n27783) );
  XNOR U27315 ( .A(n27778), .B(n27777), .Z(n27780) );
  XNOR U27316 ( .A(n27775), .B(n27774), .Z(n27777) );
  XNOR U27317 ( .A(n27772), .B(n27771), .Z(n27774) );
  XNOR U27318 ( .A(n27769), .B(n27768), .Z(n27771) );
  XNOR U27319 ( .A(n27766), .B(n27765), .Z(n27768) );
  XNOR U27320 ( .A(n27763), .B(n27762), .Z(n27765) );
  XNOR U27321 ( .A(n27760), .B(n27759), .Z(n27762) );
  XNOR U27322 ( .A(n27757), .B(n27756), .Z(n27759) );
  XNOR U27323 ( .A(n27754), .B(n27753), .Z(n27756) );
  XNOR U27324 ( .A(n27751), .B(n27750), .Z(n27753) );
  XNOR U27325 ( .A(n27748), .B(n27747), .Z(n27750) );
  XNOR U27326 ( .A(n27745), .B(n27744), .Z(n27747) );
  XNOR U27327 ( .A(n27742), .B(n27741), .Z(n27744) );
  XNOR U27328 ( .A(n27739), .B(n27738), .Z(n27741) );
  XNOR U27329 ( .A(n27736), .B(n27735), .Z(n27738) );
  XNOR U27330 ( .A(n27733), .B(n27732), .Z(n27735) );
  XNOR U27331 ( .A(n27730), .B(n27729), .Z(n27732) );
  XNOR U27332 ( .A(n27727), .B(n27726), .Z(n27729) );
  XNOR U27333 ( .A(n27724), .B(n27723), .Z(n27726) );
  XNOR U27334 ( .A(n27721), .B(n27720), .Z(n27723) );
  XNOR U27335 ( .A(n27718), .B(n27717), .Z(n27720) );
  XNOR U27336 ( .A(n27715), .B(n27714), .Z(n27717) );
  XNOR U27337 ( .A(n27712), .B(n27711), .Z(n27714) );
  XNOR U27338 ( .A(n27709), .B(n27708), .Z(n27711) );
  XNOR U27339 ( .A(n27706), .B(n27705), .Z(n27708) );
  XNOR U27340 ( .A(n27703), .B(n27702), .Z(n27705) );
  XNOR U27341 ( .A(n27700), .B(n27699), .Z(n27702) );
  XNOR U27342 ( .A(n27697), .B(n27696), .Z(n27699) );
  XNOR U27343 ( .A(n27694), .B(n27693), .Z(n27696) );
  XNOR U27344 ( .A(n27691), .B(n27690), .Z(n27693) );
  XNOR U27345 ( .A(n27688), .B(n27687), .Z(n27690) );
  XNOR U27346 ( .A(n27685), .B(n27684), .Z(n27687) );
  XNOR U27347 ( .A(n27682), .B(n27681), .Z(n27684) );
  XNOR U27348 ( .A(n27679), .B(n27678), .Z(n27681) );
  XNOR U27349 ( .A(n27676), .B(n27675), .Z(n27678) );
  XNOR U27350 ( .A(n27673), .B(n27672), .Z(n27675) );
  XNOR U27351 ( .A(n27670), .B(n27669), .Z(n27672) );
  XNOR U27352 ( .A(n27667), .B(n27666), .Z(n27669) );
  XNOR U27353 ( .A(n27664), .B(n27663), .Z(n27666) );
  XNOR U27354 ( .A(n27661), .B(n27660), .Z(n27663) );
  XNOR U27355 ( .A(n27658), .B(n27657), .Z(n27660) );
  XNOR U27356 ( .A(n27655), .B(n27654), .Z(n27657) );
  XNOR U27357 ( .A(n27652), .B(n27651), .Z(n27654) );
  XNOR U27358 ( .A(n27649), .B(n27648), .Z(n27651) );
  XNOR U27359 ( .A(n27646), .B(n27645), .Z(n27648) );
  XNOR U27360 ( .A(n27643), .B(n27642), .Z(n27645) );
  XNOR U27361 ( .A(n27640), .B(n27639), .Z(n27642) );
  XNOR U27362 ( .A(n27637), .B(n27636), .Z(n27639) );
  XNOR U27363 ( .A(n27634), .B(n27633), .Z(n27636) );
  XNOR U27364 ( .A(n27631), .B(n27630), .Z(n27633) );
  XNOR U27365 ( .A(n27628), .B(n27627), .Z(n27630) );
  XNOR U27366 ( .A(n27625), .B(n27624), .Z(n27627) );
  XNOR U27367 ( .A(n27622), .B(n27621), .Z(n27624) );
  XNOR U27368 ( .A(n27619), .B(n27618), .Z(n27621) );
  XNOR U27369 ( .A(n27616), .B(n27615), .Z(n27618) );
  XNOR U27370 ( .A(n27613), .B(n27612), .Z(n27615) );
  XNOR U27371 ( .A(n27610), .B(n27609), .Z(n27612) );
  XNOR U27372 ( .A(n27607), .B(n27606), .Z(n27609) );
  XNOR U27373 ( .A(n27604), .B(n27603), .Z(n27606) );
  XNOR U27374 ( .A(n27601), .B(n27600), .Z(n27603) );
  XNOR U27375 ( .A(n27598), .B(n27597), .Z(n27600) );
  XNOR U27376 ( .A(n27595), .B(n26976), .Z(n27597) );
  XOR U27377 ( .A(n26975), .B(n26964), .Z(n26976) );
  XOR U27378 ( .A(n29818), .B(n26962), .Z(n26964) );
  XNOR U27379 ( .A(n26963), .B(n26959), .Z(n26962) );
  XNOR U27380 ( .A(n26958), .B(n26985), .Z(n26959) );
  XNOR U27381 ( .A(n26984), .B(n27594), .Z(n26985) );
  XNOR U27382 ( .A(n27585), .B(n27593), .Z(n27594) );
  XNOR U27383 ( .A(n27584), .B(n27590), .Z(n27593) );
  XNOR U27384 ( .A(n27589), .B(n26994), .Z(n27590) );
  XNOR U27385 ( .A(n26993), .B(n27583), .Z(n26994) );
  XNOR U27386 ( .A(n27574), .B(n27582), .Z(n27583) );
  XNOR U27387 ( .A(n27573), .B(n27579), .Z(n27582) );
  XNOR U27388 ( .A(n27578), .B(n27003), .Z(n27579) );
  XNOR U27389 ( .A(n27002), .B(n27572), .Z(n27003) );
  XNOR U27390 ( .A(n27563), .B(n27571), .Z(n27572) );
  XNOR U27391 ( .A(n27562), .B(n27568), .Z(n27571) );
  XNOR U27392 ( .A(n27567), .B(n27012), .Z(n27568) );
  XNOR U27393 ( .A(n27011), .B(n27561), .Z(n27012) );
  XNOR U27394 ( .A(n27552), .B(n27560), .Z(n27561) );
  XNOR U27395 ( .A(n27551), .B(n27557), .Z(n27560) );
  XNOR U27396 ( .A(n27556), .B(n27021), .Z(n27557) );
  XNOR U27397 ( .A(n27020), .B(n27550), .Z(n27021) );
  XNOR U27398 ( .A(n27541), .B(n27549), .Z(n27550) );
  XNOR U27399 ( .A(n27540), .B(n27546), .Z(n27549) );
  XNOR U27400 ( .A(n27545), .B(n27030), .Z(n27546) );
  XNOR U27401 ( .A(n27029), .B(n27539), .Z(n27030) );
  XNOR U27402 ( .A(n27530), .B(n27538), .Z(n27539) );
  XNOR U27403 ( .A(n27529), .B(n27535), .Z(n27538) );
  XNOR U27404 ( .A(n27534), .B(n27039), .Z(n27535) );
  XNOR U27405 ( .A(n27038), .B(n27528), .Z(n27039) );
  XNOR U27406 ( .A(n27519), .B(n27527), .Z(n27528) );
  XNOR U27407 ( .A(n27518), .B(n27524), .Z(n27527) );
  XNOR U27408 ( .A(n27523), .B(n27048), .Z(n27524) );
  XNOR U27409 ( .A(n27047), .B(n27517), .Z(n27048) );
  XNOR U27410 ( .A(n27508), .B(n27516), .Z(n27517) );
  XNOR U27411 ( .A(n27507), .B(n27513), .Z(n27516) );
  XNOR U27412 ( .A(n27512), .B(n27057), .Z(n27513) );
  XNOR U27413 ( .A(n27056), .B(n27506), .Z(n27057) );
  XNOR U27414 ( .A(n27497), .B(n27505), .Z(n27506) );
  XNOR U27415 ( .A(n27496), .B(n27502), .Z(n27505) );
  XNOR U27416 ( .A(n27501), .B(n27066), .Z(n27502) );
  XNOR U27417 ( .A(n27065), .B(n27495), .Z(n27066) );
  XNOR U27418 ( .A(n27486), .B(n27494), .Z(n27495) );
  XNOR U27419 ( .A(n27485), .B(n27491), .Z(n27494) );
  XNOR U27420 ( .A(n27490), .B(n27075), .Z(n27491) );
  XNOR U27421 ( .A(n27074), .B(n27484), .Z(n27075) );
  XNOR U27422 ( .A(n27475), .B(n27483), .Z(n27484) );
  XNOR U27423 ( .A(n27474), .B(n27480), .Z(n27483) );
  XNOR U27424 ( .A(n27479), .B(n27084), .Z(n27480) );
  XNOR U27425 ( .A(n27083), .B(n27473), .Z(n27084) );
  XNOR U27426 ( .A(n27464), .B(n27472), .Z(n27473) );
  XNOR U27427 ( .A(n27463), .B(n27469), .Z(n27472) );
  XNOR U27428 ( .A(n27468), .B(n27093), .Z(n27469) );
  XNOR U27429 ( .A(n27092), .B(n27462), .Z(n27093) );
  XNOR U27430 ( .A(n27453), .B(n27461), .Z(n27462) );
  XNOR U27431 ( .A(n27452), .B(n27458), .Z(n27461) );
  XNOR U27432 ( .A(n27457), .B(n27102), .Z(n27458) );
  XNOR U27433 ( .A(n27101), .B(n27451), .Z(n27102) );
  XNOR U27434 ( .A(n27442), .B(n27450), .Z(n27451) );
  XNOR U27435 ( .A(n27441), .B(n27447), .Z(n27450) );
  XNOR U27436 ( .A(n27446), .B(n27111), .Z(n27447) );
  XNOR U27437 ( .A(n27110), .B(n27440), .Z(n27111) );
  XNOR U27438 ( .A(n27431), .B(n27439), .Z(n27440) );
  XNOR U27439 ( .A(n27430), .B(n27436), .Z(n27439) );
  XNOR U27440 ( .A(n27435), .B(n27120), .Z(n27436) );
  XNOR U27441 ( .A(n27119), .B(n27429), .Z(n27120) );
  XNOR U27442 ( .A(n27420), .B(n27428), .Z(n27429) );
  XNOR U27443 ( .A(n27419), .B(n27425), .Z(n27428) );
  XNOR U27444 ( .A(n27424), .B(n27129), .Z(n27425) );
  XNOR U27445 ( .A(n27128), .B(n27418), .Z(n27129) );
  XNOR U27446 ( .A(n27409), .B(n27417), .Z(n27418) );
  XNOR U27447 ( .A(n27408), .B(n27414), .Z(n27417) );
  XNOR U27448 ( .A(n27413), .B(n27138), .Z(n27414) );
  XNOR U27449 ( .A(n27137), .B(n27407), .Z(n27138) );
  XNOR U27450 ( .A(n27398), .B(n27406), .Z(n27407) );
  XNOR U27451 ( .A(n27397), .B(n27403), .Z(n27406) );
  XNOR U27452 ( .A(n27402), .B(n27147), .Z(n27403) );
  XNOR U27453 ( .A(n27146), .B(n27396), .Z(n27147) );
  XNOR U27454 ( .A(n27387), .B(n27395), .Z(n27396) );
  XNOR U27455 ( .A(n27386), .B(n27392), .Z(n27395) );
  XNOR U27456 ( .A(n27391), .B(n27156), .Z(n27392) );
  XNOR U27457 ( .A(n27155), .B(n27385), .Z(n27156) );
  XNOR U27458 ( .A(n27376), .B(n27384), .Z(n27385) );
  XNOR U27459 ( .A(n27375), .B(n27381), .Z(n27384) );
  XNOR U27460 ( .A(n27380), .B(n27165), .Z(n27381) );
  XNOR U27461 ( .A(n27164), .B(n27374), .Z(n27165) );
  XNOR U27462 ( .A(n27365), .B(n27373), .Z(n27374) );
  XNOR U27463 ( .A(n27364), .B(n27370), .Z(n27373) );
  XNOR U27464 ( .A(n27369), .B(n27174), .Z(n27370) );
  XNOR U27465 ( .A(n27173), .B(n27363), .Z(n27174) );
  XNOR U27466 ( .A(n27354), .B(n27362), .Z(n27363) );
  XNOR U27467 ( .A(n27353), .B(n27359), .Z(n27362) );
  XNOR U27468 ( .A(n27358), .B(n27183), .Z(n27359) );
  XNOR U27469 ( .A(n27182), .B(n27352), .Z(n27183) );
  XNOR U27470 ( .A(n27343), .B(n27351), .Z(n27352) );
  XNOR U27471 ( .A(n27342), .B(n27348), .Z(n27351) );
  XNOR U27472 ( .A(n27347), .B(n27192), .Z(n27348) );
  XNOR U27473 ( .A(n27191), .B(n27341), .Z(n27192) );
  XNOR U27474 ( .A(n27332), .B(n27340), .Z(n27341) );
  XNOR U27475 ( .A(n27331), .B(n27337), .Z(n27340) );
  XNOR U27476 ( .A(n27336), .B(n27201), .Z(n27337) );
  XNOR U27477 ( .A(n27200), .B(n27330), .Z(n27201) );
  XNOR U27478 ( .A(n27321), .B(n27329), .Z(n27330) );
  XNOR U27479 ( .A(n27320), .B(n27326), .Z(n27329) );
  XNOR U27480 ( .A(n27325), .B(n27210), .Z(n27326) );
  XNOR U27481 ( .A(n27209), .B(n27319), .Z(n27210) );
  XNOR U27482 ( .A(n27310), .B(n27318), .Z(n27319) );
  XNOR U27483 ( .A(n27309), .B(n27315), .Z(n27318) );
  XNOR U27484 ( .A(n27314), .B(n27219), .Z(n27315) );
  XNOR U27485 ( .A(n27218), .B(n27308), .Z(n27219) );
  XNOR U27486 ( .A(n27299), .B(n27307), .Z(n27308) );
  XNOR U27487 ( .A(n27298), .B(n27304), .Z(n27307) );
  XNOR U27488 ( .A(n27303), .B(n27228), .Z(n27304) );
  XNOR U27489 ( .A(n27227), .B(n27297), .Z(n27228) );
  XNOR U27490 ( .A(n27288), .B(n27296), .Z(n27297) );
  XNOR U27491 ( .A(n27287), .B(n27293), .Z(n27296) );
  XNOR U27492 ( .A(n27292), .B(n27275), .Z(n27293) );
  XNOR U27493 ( .A(n27234), .B(n27286), .Z(n27275) );
  XNOR U27494 ( .A(n27277), .B(n27285), .Z(n27286) );
  XNOR U27495 ( .A(n27276), .B(n27282), .Z(n27285) );
  XNOR U27496 ( .A(n27281), .B(n27265), .Z(n27282) );
  XNOR U27497 ( .A(n27237), .B(n27274), .Z(n27265) );
  XNOR U27498 ( .A(n27261), .B(n27271), .Z(n27274) );
  XNOR U27499 ( .A(n27264), .B(n27270), .Z(n27271) );
  XNOR U27500 ( .A(n27233), .B(n27260), .Z(n27270) );
  XNOR U27501 ( .A(n27243), .B(n27259), .Z(n27260) );
  XNOR U27502 ( .A(n27246), .B(n27256), .Z(n27259) );
  XOR U27503 ( .A(n27245), .B(n27253), .Z(n27256) );
  XOR U27504 ( .A(n27254), .B(n27252), .Z(n27253) );
  XOR U27505 ( .A(n29819), .B(n29820), .Z(n27252) );
  XOR U27506 ( .A(n29821), .B(n29822), .Z(n29820) );
  XNOR U27507 ( .A(n29823), .B(n29824), .Z(n29822) );
  NOR U27508 ( .A(n29825), .B(n29824), .Z(n29823) );
  XOR U27509 ( .A(n29826), .B(n29827), .Z(n29821) );
  NOR U27510 ( .A(n29828), .B(n29829), .Z(n29827) );
  NOR U27511 ( .A(n29830), .B(n29831), .Z(n29826) );
  XOR U27512 ( .A(n29832), .B(n29833), .Z(n29819) );
  XOR U27513 ( .A(n29834), .B(n29835), .Z(n29833) );
  XOR U27514 ( .A(n29836), .B(n29837), .Z(n29835) );
  XOR U27515 ( .A(n29838), .B(n29839), .Z(n29837) );
  XOR U27516 ( .A(n29840), .B(n29841), .Z(n29839) );
  AND U27517 ( .A(n29842), .B(n29841), .Z(n29840) );
  XOR U27518 ( .A(n29843), .B(n29844), .Z(n29838) );
  XOR U27519 ( .A(n29845), .B(n29846), .Z(n29844) );
  XOR U27520 ( .A(n29847), .B(n29848), .Z(n29846) );
  XNOR U27521 ( .A(n29849), .B(n29850), .Z(n29848) );
  NOR U27522 ( .A(n29851), .B(n29850), .Z(n29849) );
  XOR U27523 ( .A(n29852), .B(n29853), .Z(n29847) );
  XOR U27524 ( .A(n29854), .B(n29855), .Z(n29853) );
  XNOR U27525 ( .A(n29856), .B(n29857), .Z(n29855) );
  XOR U27526 ( .A(n29858), .B(n29859), .Z(n29854) );
  XOR U27527 ( .A(n29860), .B(n29861), .Z(n29859) );
  XOR U27528 ( .A(n29862), .B(n29863), .Z(n29861) );
  XOR U27529 ( .A(n29864), .B(n29865), .Z(n29863) );
  XOR U27530 ( .A(n29866), .B(n29867), .Z(n29865) );
  XOR U27531 ( .A(n29868), .B(n29869), .Z(n29867) );
  XOR U27532 ( .A(n29870), .B(n29871), .Z(n29869) );
  XOR U27533 ( .A(n29872), .B(n29873), .Z(n29871) );
  XOR U27534 ( .A(n29874), .B(n29875), .Z(n29873) );
  XOR U27535 ( .A(n29876), .B(n29877), .Z(n29875) );
  XOR U27536 ( .A(n29878), .B(n29879), .Z(n29877) );
  XOR U27537 ( .A(n29880), .B(n29881), .Z(n29879) );
  XOR U27538 ( .A(n29882), .B(n29883), .Z(n29881) );
  XOR U27539 ( .A(n29884), .B(n29885), .Z(n29883) );
  XOR U27540 ( .A(n29886), .B(n29887), .Z(n29885) );
  XOR U27541 ( .A(n29888), .B(n29889), .Z(n29887) );
  XOR U27542 ( .A(n29890), .B(n29891), .Z(n29889) );
  AND U27543 ( .A(n29892), .B(n29893), .Z(n29891) );
  AND U27544 ( .A(n29894), .B(n29895), .Z(n29890) );
  XOR U27545 ( .A(n29896), .B(n29897), .Z(n29888) );
  AND U27546 ( .A(n29898), .B(n29899), .Z(n29897) );
  NOR U27547 ( .A(n29900), .B(n29901), .Z(n29899) );
  IV U27548 ( .A(n29902), .Z(n29900) );
  NOR U27549 ( .A(n29903), .B(n29904), .Z(n29902) );
  AND U27550 ( .A(n29905), .B(n29906), .Z(n29898) );
  NOR U27551 ( .A(n29907), .B(n29908), .Z(n29905) );
  NOR U27552 ( .A(n29909), .B(n29910), .Z(n29896) );
  XOR U27553 ( .A(n29911), .B(n29912), .Z(n29886) );
  XOR U27554 ( .A(n29913), .B(n29914), .Z(n29912) );
  NOR U27555 ( .A(n29915), .B(n29916), .Z(n29914) );
  AND U27556 ( .A(n29917), .B(n29918), .Z(n29916) );
  IV U27557 ( .A(n29919), .Z(n29915) );
  NOR U27558 ( .A(n29920), .B(n29921), .Z(n29919) );
  AND U27559 ( .A(n29909), .B(n29922), .Z(n29921) );
  AND U27560 ( .A(n29910), .B(n29923), .Z(n29920) );
  NOR U27561 ( .A(n29924), .B(n29925), .Z(n29913) );
  XOR U27562 ( .A(n29926), .B(n29927), .Z(n29911) );
  NOR U27563 ( .A(n29928), .B(n29929), .Z(n29927) );
  AND U27564 ( .A(n29930), .B(n29931), .Z(n29929) );
  IV U27565 ( .A(n29932), .Z(n29928) );
  NOR U27566 ( .A(n29933), .B(n29934), .Z(n29932) );
  AND U27567 ( .A(n29924), .B(n29935), .Z(n29934) );
  AND U27568 ( .A(n29925), .B(n29936), .Z(n29933) );
  NOR U27569 ( .A(n29937), .B(n29938), .Z(n29926) );
  AND U27570 ( .A(n29939), .B(n29940), .Z(n29884) );
  XOR U27571 ( .A(n29941), .B(n29942), .Z(n29882) );
  AND U27572 ( .A(n29943), .B(n29944), .Z(n29942) );
  NOR U27573 ( .A(n29945), .B(n29946), .Z(n29941) );
  AND U27574 ( .A(n29947), .B(n29948), .Z(n29946) );
  IV U27575 ( .A(n29949), .Z(n29945) );
  NOR U27576 ( .A(n29950), .B(n29951), .Z(n29949) );
  AND U27577 ( .A(n29937), .B(n29952), .Z(n29951) );
  AND U27578 ( .A(n29938), .B(n29953), .Z(n29950) );
  XOR U27579 ( .A(n29954), .B(n29955), .Z(n29880) );
  XOR U27580 ( .A(n29956), .B(n29957), .Z(n29955) );
  NOR U27581 ( .A(n29958), .B(n29959), .Z(n29957) );
  NOR U27582 ( .A(n29960), .B(n29961), .Z(n29956) );
  AND U27583 ( .A(n29962), .B(n29963), .Z(n29961) );
  IV U27584 ( .A(n29964), .Z(n29960) );
  NOR U27585 ( .A(n29965), .B(n29966), .Z(n29964) );
  AND U27586 ( .A(n29958), .B(n29967), .Z(n29966) );
  AND U27587 ( .A(n29959), .B(n29968), .Z(n29965) );
  XOR U27588 ( .A(n29969), .B(n29970), .Z(n29954) );
  NOR U27589 ( .A(n29971), .B(n29972), .Z(n29970) );
  NOR U27590 ( .A(n29973), .B(n29974), .Z(n29969) );
  AND U27591 ( .A(n29975), .B(n29976), .Z(n29974) );
  IV U27592 ( .A(n29977), .Z(n29973) );
  NOR U27593 ( .A(n29978), .B(n29979), .Z(n29977) );
  AND U27594 ( .A(n29971), .B(n29980), .Z(n29979) );
  AND U27595 ( .A(n29972), .B(n29981), .Z(n29978) );
  AND U27596 ( .A(n29982), .B(n29983), .Z(n29878) );
  XOR U27597 ( .A(n29984), .B(n29985), .Z(n29876) );
  AND U27598 ( .A(n29986), .B(n29987), .Z(n29985) );
  AND U27599 ( .A(n29988), .B(n29989), .Z(n29984) );
  XOR U27600 ( .A(n29990), .B(n29991), .Z(n29874) );
  XOR U27601 ( .A(n29992), .B(n29993), .Z(n29991) );
  NOR U27602 ( .A(n29994), .B(n29995), .Z(n29993) );
  NOR U27603 ( .A(n29996), .B(n29997), .Z(n29992) );
  AND U27604 ( .A(n29998), .B(n29999), .Z(n29997) );
  IV U27605 ( .A(n30000), .Z(n29996) );
  NOR U27606 ( .A(n30001), .B(n30002), .Z(n30000) );
  AND U27607 ( .A(n29994), .B(n30003), .Z(n30002) );
  AND U27608 ( .A(n29995), .B(n30004), .Z(n30001) );
  XOR U27609 ( .A(n30005), .B(n30006), .Z(n29990) );
  NOR U27610 ( .A(n30007), .B(n30008), .Z(n30006) );
  NOR U27611 ( .A(n30009), .B(n30010), .Z(n30005) );
  AND U27612 ( .A(n30011), .B(n30012), .Z(n30010) );
  IV U27613 ( .A(n30013), .Z(n30009) );
  NOR U27614 ( .A(n30014), .B(n30015), .Z(n30013) );
  AND U27615 ( .A(n30007), .B(n30016), .Z(n30015) );
  AND U27616 ( .A(n30008), .B(n30017), .Z(n30014) );
  AND U27617 ( .A(n30018), .B(n30019), .Z(n29872) );
  XOR U27618 ( .A(n30020), .B(n30021), .Z(n29870) );
  AND U27619 ( .A(n30022), .B(n30023), .Z(n30021) );
  NOR U27620 ( .A(n30024), .B(n30025), .Z(n30020) );
  XOR U27621 ( .A(n30026), .B(n30027), .Z(n29868) );
  XOR U27622 ( .A(n30028), .B(n30029), .Z(n30027) );
  NOR U27623 ( .A(n30030), .B(n30031), .Z(n30029) );
  AND U27624 ( .A(n30032), .B(n30033), .Z(n30031) );
  IV U27625 ( .A(n30034), .Z(n30030) );
  NOR U27626 ( .A(n30035), .B(n30036), .Z(n30034) );
  AND U27627 ( .A(n30024), .B(n30037), .Z(n30036) );
  AND U27628 ( .A(n30025), .B(n30038), .Z(n30035) );
  NOR U27629 ( .A(n30039), .B(n30040), .Z(n30028) );
  XOR U27630 ( .A(n30041), .B(n30042), .Z(n30026) );
  NOR U27631 ( .A(n30043), .B(n30044), .Z(n30042) );
  AND U27632 ( .A(n30045), .B(n30046), .Z(n30044) );
  IV U27633 ( .A(n30047), .Z(n30043) );
  NOR U27634 ( .A(n30048), .B(n30049), .Z(n30047) );
  AND U27635 ( .A(n30039), .B(n30050), .Z(n30049) );
  AND U27636 ( .A(n30040), .B(n30051), .Z(n30048) );
  NOR U27637 ( .A(n30052), .B(n30053), .Z(n30041) );
  NOR U27638 ( .A(n30054), .B(n30055), .Z(n29866) );
  AND U27639 ( .A(n30056), .B(n30057), .Z(n30055) );
  IV U27640 ( .A(n30058), .Z(n30054) );
  NOR U27641 ( .A(n30059), .B(n30060), .Z(n30058) );
  AND U27642 ( .A(n30052), .B(n30061), .Z(n30060) );
  AND U27643 ( .A(n30053), .B(n30062), .Z(n30059) );
  XOR U27644 ( .A(n30063), .B(n30064), .Z(n29864) );
  NOR U27645 ( .A(n30065), .B(n30066), .Z(n30064) );
  AND U27646 ( .A(n30067), .B(n30068), .Z(n30063) );
  XOR U27647 ( .A(n30069), .B(n30070), .Z(n29862) );
  XOR U27648 ( .A(n30071), .B(n30072), .Z(n30070) );
  AND U27649 ( .A(n30065), .B(n30073), .Z(n30071) );
  XOR U27650 ( .A(n30074), .B(n30075), .Z(n30069) );
  AND U27651 ( .A(n30066), .B(n30076), .Z(n30075) );
  AND U27652 ( .A(n30072), .B(n30077), .Z(n30074) );
  XOR U27653 ( .A(n30078), .B(n30079), .Z(n29858) );
  XOR U27654 ( .A(n30080), .B(n30081), .Z(n30079) );
  AND U27655 ( .A(n30082), .B(n29860), .Z(n30080) );
  XOR U27656 ( .A(n30083), .B(n30084), .Z(n29852) );
  XOR U27657 ( .A(n30085), .B(n30086), .Z(n30084) );
  AND U27658 ( .A(n29856), .B(n30087), .Z(n30086) );
  AND U27659 ( .A(n30088), .B(n30081), .Z(n30085) );
  XOR U27660 ( .A(n30089), .B(n30090), .Z(n30083) );
  AND U27661 ( .A(n30091), .B(n30078), .Z(n30090) );
  NOR U27662 ( .A(n30092), .B(n29857), .Z(n30089) );
  XOR U27663 ( .A(n30093), .B(n30094), .Z(n29845) );
  XOR U27664 ( .A(n30095), .B(n30096), .Z(n29843) );
  XOR U27665 ( .A(n30097), .B(n30098), .Z(n30096) );
  AND U27666 ( .A(n30099), .B(n30098), .Z(n30097) );
  XOR U27667 ( .A(n30100), .B(n30101), .Z(n30095) );
  NOR U27668 ( .A(n30102), .B(n30093), .Z(n30101) );
  NOR U27669 ( .A(n30103), .B(n30094), .Z(n30100) );
  XOR U27670 ( .A(n30104), .B(n30105), .Z(n29836) );
  XOR U27671 ( .A(n30106), .B(n30107), .Z(n29834) );
  XNOR U27672 ( .A(n30108), .B(n30109), .Z(n30107) );
  NOR U27673 ( .A(n30110), .B(n30109), .Z(n30108) );
  XOR U27674 ( .A(n30111), .B(n30112), .Z(n30106) );
  NOR U27675 ( .A(n30113), .B(n30104), .Z(n30112) );
  NOR U27676 ( .A(n30114), .B(n30105), .Z(n30111) );
  XNOR U27677 ( .A(n29831), .B(n29829), .Z(n29832) );
  XNOR U27678 ( .A(n30115), .B(n30116), .Z(n27254) );
  NOR U27679 ( .A(n30117), .B(n30115), .Z(n30116) );
  XOR U27680 ( .A(n30118), .B(n30119), .Z(n27245) );
  NOR U27681 ( .A(n30120), .B(n30118), .Z(n30119) );
  XOR U27682 ( .A(n30121), .B(n30122), .Z(n27246) );
  NOR U27683 ( .A(n30123), .B(n30121), .Z(n30122) );
  XOR U27684 ( .A(n30124), .B(n30125), .Z(n27243) );
  NOR U27685 ( .A(n30126), .B(n30124), .Z(n30125) );
  XOR U27686 ( .A(n30127), .B(n30128), .Z(n27233) );
  NOR U27687 ( .A(n30129), .B(n30127), .Z(n30128) );
  XOR U27688 ( .A(n30130), .B(n30131), .Z(n27264) );
  NOR U27689 ( .A(n30132), .B(n30130), .Z(n30131) );
  XOR U27690 ( .A(n30133), .B(n30134), .Z(n27261) );
  NOR U27691 ( .A(n30135), .B(n30133), .Z(n30134) );
  XOR U27692 ( .A(n30136), .B(n30137), .Z(n27237) );
  NOR U27693 ( .A(n30138), .B(n30136), .Z(n30137) );
  XOR U27694 ( .A(n30139), .B(n30140), .Z(n27281) );
  NOR U27695 ( .A(n30141), .B(n30139), .Z(n30140) );
  XOR U27696 ( .A(n30142), .B(n30143), .Z(n27276) );
  NOR U27697 ( .A(n30144), .B(n30142), .Z(n30143) );
  XOR U27698 ( .A(n30145), .B(n30146), .Z(n27277) );
  NOR U27699 ( .A(n30147), .B(n30145), .Z(n30146) );
  XOR U27700 ( .A(n30148), .B(n30149), .Z(n27234) );
  NOR U27701 ( .A(n30150), .B(n30148), .Z(n30149) );
  XOR U27702 ( .A(n30151), .B(n30152), .Z(n27292) );
  NOR U27703 ( .A(n30153), .B(n30151), .Z(n30152) );
  XOR U27704 ( .A(n30154), .B(n30155), .Z(n27287) );
  NOR U27705 ( .A(n30156), .B(n30154), .Z(n30155) );
  XOR U27706 ( .A(n30157), .B(n30158), .Z(n27288) );
  NOR U27707 ( .A(n30159), .B(n30157), .Z(n30158) );
  XOR U27708 ( .A(n30160), .B(n30161), .Z(n27227) );
  NOR U27709 ( .A(n30162), .B(n30160), .Z(n30161) );
  XOR U27710 ( .A(n30163), .B(n30164), .Z(n27303) );
  NOR U27711 ( .A(n30165), .B(n30163), .Z(n30164) );
  XOR U27712 ( .A(n30166), .B(n30167), .Z(n27298) );
  NOR U27713 ( .A(n30168), .B(n30166), .Z(n30167) );
  XOR U27714 ( .A(n30169), .B(n30170), .Z(n27299) );
  NOR U27715 ( .A(n30171), .B(n30169), .Z(n30170) );
  XOR U27716 ( .A(n30172), .B(n30173), .Z(n27218) );
  NOR U27717 ( .A(n30174), .B(n30172), .Z(n30173) );
  XOR U27718 ( .A(n30175), .B(n30176), .Z(n27314) );
  NOR U27719 ( .A(n30177), .B(n30175), .Z(n30176) );
  XOR U27720 ( .A(n30178), .B(n30179), .Z(n27309) );
  NOR U27721 ( .A(n30180), .B(n30178), .Z(n30179) );
  XOR U27722 ( .A(n30181), .B(n30182), .Z(n27310) );
  NOR U27723 ( .A(n30183), .B(n30181), .Z(n30182) );
  XOR U27724 ( .A(n30184), .B(n30185), .Z(n27209) );
  NOR U27725 ( .A(n30186), .B(n30184), .Z(n30185) );
  XOR U27726 ( .A(n30187), .B(n30188), .Z(n27325) );
  NOR U27727 ( .A(n30189), .B(n30187), .Z(n30188) );
  XOR U27728 ( .A(n30190), .B(n30191), .Z(n27320) );
  NOR U27729 ( .A(n30192), .B(n30190), .Z(n30191) );
  XOR U27730 ( .A(n30193), .B(n30194), .Z(n27321) );
  NOR U27731 ( .A(n30195), .B(n30193), .Z(n30194) );
  XOR U27732 ( .A(n30196), .B(n30197), .Z(n27200) );
  NOR U27733 ( .A(n30198), .B(n30196), .Z(n30197) );
  XOR U27734 ( .A(n30199), .B(n30200), .Z(n27336) );
  NOR U27735 ( .A(n30201), .B(n30199), .Z(n30200) );
  XOR U27736 ( .A(n30202), .B(n30203), .Z(n27331) );
  NOR U27737 ( .A(n30204), .B(n30202), .Z(n30203) );
  XOR U27738 ( .A(n30205), .B(n30206), .Z(n27332) );
  NOR U27739 ( .A(n30207), .B(n30205), .Z(n30206) );
  XOR U27740 ( .A(n30208), .B(n30209), .Z(n27191) );
  NOR U27741 ( .A(n30210), .B(n30208), .Z(n30209) );
  XOR U27742 ( .A(n30211), .B(n30212), .Z(n27347) );
  NOR U27743 ( .A(n30213), .B(n30211), .Z(n30212) );
  XOR U27744 ( .A(n30214), .B(n30215), .Z(n27342) );
  NOR U27745 ( .A(n30216), .B(n30214), .Z(n30215) );
  XOR U27746 ( .A(n30217), .B(n30218), .Z(n27343) );
  NOR U27747 ( .A(n30219), .B(n30217), .Z(n30218) );
  XOR U27748 ( .A(n30220), .B(n30221), .Z(n27182) );
  NOR U27749 ( .A(n30222), .B(n30220), .Z(n30221) );
  XOR U27750 ( .A(n30223), .B(n30224), .Z(n27358) );
  NOR U27751 ( .A(n30225), .B(n30223), .Z(n30224) );
  XOR U27752 ( .A(n30226), .B(n30227), .Z(n27353) );
  NOR U27753 ( .A(n30228), .B(n30226), .Z(n30227) );
  XOR U27754 ( .A(n30229), .B(n30230), .Z(n27354) );
  NOR U27755 ( .A(n30231), .B(n30229), .Z(n30230) );
  XOR U27756 ( .A(n30232), .B(n30233), .Z(n27173) );
  NOR U27757 ( .A(n30234), .B(n30232), .Z(n30233) );
  XOR U27758 ( .A(n30235), .B(n30236), .Z(n27369) );
  NOR U27759 ( .A(n30237), .B(n30235), .Z(n30236) );
  XOR U27760 ( .A(n30238), .B(n30239), .Z(n27364) );
  NOR U27761 ( .A(n30240), .B(n30238), .Z(n30239) );
  XOR U27762 ( .A(n30241), .B(n30242), .Z(n27365) );
  NOR U27763 ( .A(n30243), .B(n30241), .Z(n30242) );
  XOR U27764 ( .A(n30244), .B(n30245), .Z(n27164) );
  NOR U27765 ( .A(n30246), .B(n30244), .Z(n30245) );
  XOR U27766 ( .A(n30247), .B(n30248), .Z(n27380) );
  NOR U27767 ( .A(n30249), .B(n30247), .Z(n30248) );
  XOR U27768 ( .A(n30250), .B(n30251), .Z(n27375) );
  NOR U27769 ( .A(n30252), .B(n30250), .Z(n30251) );
  XOR U27770 ( .A(n30253), .B(n30254), .Z(n27376) );
  NOR U27771 ( .A(n30255), .B(n30253), .Z(n30254) );
  XOR U27772 ( .A(n30256), .B(n30257), .Z(n27155) );
  NOR U27773 ( .A(n30258), .B(n30256), .Z(n30257) );
  XOR U27774 ( .A(n30259), .B(n30260), .Z(n27391) );
  NOR U27775 ( .A(n30261), .B(n30259), .Z(n30260) );
  XOR U27776 ( .A(n30262), .B(n30263), .Z(n27386) );
  NOR U27777 ( .A(n30264), .B(n30262), .Z(n30263) );
  XOR U27778 ( .A(n30265), .B(n30266), .Z(n27387) );
  NOR U27779 ( .A(n30267), .B(n30265), .Z(n30266) );
  XOR U27780 ( .A(n30268), .B(n30269), .Z(n27146) );
  NOR U27781 ( .A(n30270), .B(n30268), .Z(n30269) );
  XOR U27782 ( .A(n30271), .B(n30272), .Z(n27402) );
  NOR U27783 ( .A(n30273), .B(n30271), .Z(n30272) );
  XOR U27784 ( .A(n30274), .B(n30275), .Z(n27397) );
  NOR U27785 ( .A(n30276), .B(n30274), .Z(n30275) );
  XOR U27786 ( .A(n30277), .B(n30278), .Z(n27398) );
  NOR U27787 ( .A(n30279), .B(n30277), .Z(n30278) );
  XOR U27788 ( .A(n30280), .B(n30281), .Z(n27137) );
  NOR U27789 ( .A(n30282), .B(n30280), .Z(n30281) );
  XOR U27790 ( .A(n30283), .B(n30284), .Z(n27413) );
  NOR U27791 ( .A(n30285), .B(n30283), .Z(n30284) );
  XOR U27792 ( .A(n30286), .B(n30287), .Z(n27408) );
  NOR U27793 ( .A(n30288), .B(n30286), .Z(n30287) );
  XOR U27794 ( .A(n30289), .B(n30290), .Z(n27409) );
  NOR U27795 ( .A(n30291), .B(n30289), .Z(n30290) );
  XOR U27796 ( .A(n30292), .B(n30293), .Z(n27128) );
  NOR U27797 ( .A(n30294), .B(n30292), .Z(n30293) );
  XOR U27798 ( .A(n30295), .B(n30296), .Z(n27424) );
  NOR U27799 ( .A(n30297), .B(n30295), .Z(n30296) );
  XOR U27800 ( .A(n30298), .B(n30299), .Z(n27419) );
  NOR U27801 ( .A(n30300), .B(n30298), .Z(n30299) );
  XOR U27802 ( .A(n30301), .B(n30302), .Z(n27420) );
  NOR U27803 ( .A(n30303), .B(n30301), .Z(n30302) );
  XOR U27804 ( .A(n30304), .B(n30305), .Z(n27119) );
  NOR U27805 ( .A(n30306), .B(n30304), .Z(n30305) );
  XOR U27806 ( .A(n30307), .B(n30308), .Z(n27435) );
  NOR U27807 ( .A(n30309), .B(n30307), .Z(n30308) );
  XOR U27808 ( .A(n30310), .B(n30311), .Z(n27430) );
  NOR U27809 ( .A(n30312), .B(n30310), .Z(n30311) );
  XOR U27810 ( .A(n30313), .B(n30314), .Z(n27431) );
  NOR U27811 ( .A(n30315), .B(n30313), .Z(n30314) );
  XOR U27812 ( .A(n30316), .B(n30317), .Z(n27110) );
  NOR U27813 ( .A(n30318), .B(n30316), .Z(n30317) );
  XOR U27814 ( .A(n30319), .B(n30320), .Z(n27446) );
  NOR U27815 ( .A(n30321), .B(n30319), .Z(n30320) );
  XOR U27816 ( .A(n30322), .B(n30323), .Z(n27441) );
  NOR U27817 ( .A(n30324), .B(n30322), .Z(n30323) );
  XOR U27818 ( .A(n30325), .B(n30326), .Z(n27442) );
  NOR U27819 ( .A(n30327), .B(n30325), .Z(n30326) );
  XOR U27820 ( .A(n30328), .B(n30329), .Z(n27101) );
  NOR U27821 ( .A(n30330), .B(n30328), .Z(n30329) );
  XOR U27822 ( .A(n30331), .B(n30332), .Z(n27457) );
  NOR U27823 ( .A(n30333), .B(n30331), .Z(n30332) );
  XOR U27824 ( .A(n30334), .B(n30335), .Z(n27452) );
  NOR U27825 ( .A(n30336), .B(n30334), .Z(n30335) );
  XOR U27826 ( .A(n30337), .B(n30338), .Z(n27453) );
  NOR U27827 ( .A(n30339), .B(n30337), .Z(n30338) );
  XOR U27828 ( .A(n30340), .B(n30341), .Z(n27092) );
  NOR U27829 ( .A(n30342), .B(n30340), .Z(n30341) );
  XOR U27830 ( .A(n30343), .B(n30344), .Z(n27468) );
  NOR U27831 ( .A(n30345), .B(n30343), .Z(n30344) );
  XOR U27832 ( .A(n30346), .B(n30347), .Z(n27463) );
  NOR U27833 ( .A(n30348), .B(n30346), .Z(n30347) );
  XOR U27834 ( .A(n30349), .B(n30350), .Z(n27464) );
  NOR U27835 ( .A(n30351), .B(n30349), .Z(n30350) );
  XOR U27836 ( .A(n30352), .B(n30353), .Z(n27083) );
  NOR U27837 ( .A(n30354), .B(n30352), .Z(n30353) );
  XOR U27838 ( .A(n30355), .B(n30356), .Z(n27479) );
  NOR U27839 ( .A(n30357), .B(n30355), .Z(n30356) );
  XOR U27840 ( .A(n30358), .B(n30359), .Z(n27474) );
  NOR U27841 ( .A(n30360), .B(n30358), .Z(n30359) );
  XOR U27842 ( .A(n30361), .B(n30362), .Z(n27475) );
  NOR U27843 ( .A(n30363), .B(n30361), .Z(n30362) );
  XOR U27844 ( .A(n30364), .B(n30365), .Z(n27074) );
  NOR U27845 ( .A(n30366), .B(n30364), .Z(n30365) );
  XOR U27846 ( .A(n30367), .B(n30368), .Z(n27490) );
  NOR U27847 ( .A(n30369), .B(n30367), .Z(n30368) );
  XOR U27848 ( .A(n30370), .B(n30371), .Z(n27485) );
  NOR U27849 ( .A(n30372), .B(n30370), .Z(n30371) );
  XOR U27850 ( .A(n30373), .B(n30374), .Z(n27486) );
  NOR U27851 ( .A(n30375), .B(n30373), .Z(n30374) );
  XOR U27852 ( .A(n30376), .B(n30377), .Z(n27065) );
  NOR U27853 ( .A(n30378), .B(n30376), .Z(n30377) );
  XOR U27854 ( .A(n30379), .B(n30380), .Z(n27501) );
  NOR U27855 ( .A(n30381), .B(n30379), .Z(n30380) );
  XOR U27856 ( .A(n30382), .B(n30383), .Z(n27496) );
  NOR U27857 ( .A(n30384), .B(n30382), .Z(n30383) );
  XOR U27858 ( .A(n30385), .B(n30386), .Z(n27497) );
  NOR U27859 ( .A(n30387), .B(n30385), .Z(n30386) );
  XOR U27860 ( .A(n30388), .B(n30389), .Z(n27056) );
  NOR U27861 ( .A(n30390), .B(n30388), .Z(n30389) );
  XOR U27862 ( .A(n30391), .B(n30392), .Z(n27512) );
  NOR U27863 ( .A(n30393), .B(n30391), .Z(n30392) );
  XOR U27864 ( .A(n30394), .B(n30395), .Z(n27507) );
  NOR U27865 ( .A(n30396), .B(n30394), .Z(n30395) );
  XOR U27866 ( .A(n30397), .B(n30398), .Z(n27508) );
  NOR U27867 ( .A(n30399), .B(n30397), .Z(n30398) );
  XOR U27868 ( .A(n30400), .B(n30401), .Z(n27047) );
  NOR U27869 ( .A(n30402), .B(n30400), .Z(n30401) );
  XOR U27870 ( .A(n30403), .B(n30404), .Z(n27523) );
  NOR U27871 ( .A(n30405), .B(n30403), .Z(n30404) );
  XOR U27872 ( .A(n30406), .B(n30407), .Z(n27518) );
  NOR U27873 ( .A(n30408), .B(n30406), .Z(n30407) );
  XOR U27874 ( .A(n30409), .B(n30410), .Z(n27519) );
  NOR U27875 ( .A(n30411), .B(n30409), .Z(n30410) );
  XOR U27876 ( .A(n30412), .B(n30413), .Z(n27038) );
  NOR U27877 ( .A(n30414), .B(n30412), .Z(n30413) );
  XOR U27878 ( .A(n30415), .B(n30416), .Z(n27534) );
  NOR U27879 ( .A(n30417), .B(n30415), .Z(n30416) );
  XOR U27880 ( .A(n30418), .B(n30419), .Z(n27529) );
  NOR U27881 ( .A(n30420), .B(n30418), .Z(n30419) );
  XOR U27882 ( .A(n30421), .B(n30422), .Z(n27530) );
  NOR U27883 ( .A(n30423), .B(n30421), .Z(n30422) );
  XOR U27884 ( .A(n30424), .B(n30425), .Z(n27029) );
  NOR U27885 ( .A(n30426), .B(n30424), .Z(n30425) );
  XOR U27886 ( .A(n30427), .B(n30428), .Z(n27545) );
  NOR U27887 ( .A(n30429), .B(n30427), .Z(n30428) );
  XOR U27888 ( .A(n30430), .B(n30431), .Z(n27540) );
  NOR U27889 ( .A(n30432), .B(n30430), .Z(n30431) );
  XOR U27890 ( .A(n30433), .B(n30434), .Z(n27541) );
  NOR U27891 ( .A(n30435), .B(n30433), .Z(n30434) );
  XOR U27892 ( .A(n30436), .B(n30437), .Z(n27020) );
  NOR U27893 ( .A(n30438), .B(n30436), .Z(n30437) );
  XOR U27894 ( .A(n30439), .B(n30440), .Z(n27556) );
  NOR U27895 ( .A(n30441), .B(n30439), .Z(n30440) );
  XOR U27896 ( .A(n30442), .B(n30443), .Z(n27551) );
  NOR U27897 ( .A(n30444), .B(n30442), .Z(n30443) );
  XOR U27898 ( .A(n30445), .B(n30446), .Z(n27552) );
  NOR U27899 ( .A(n30447), .B(n30445), .Z(n30446) );
  XOR U27900 ( .A(n30448), .B(n30449), .Z(n27011) );
  NOR U27901 ( .A(n30450), .B(n30448), .Z(n30449) );
  XOR U27902 ( .A(n30451), .B(n30452), .Z(n27567) );
  NOR U27903 ( .A(n30453), .B(n30451), .Z(n30452) );
  XOR U27904 ( .A(n30454), .B(n30455), .Z(n27562) );
  NOR U27905 ( .A(n30456), .B(n30454), .Z(n30455) );
  XOR U27906 ( .A(n30457), .B(n30458), .Z(n27563) );
  NOR U27907 ( .A(n30459), .B(n30457), .Z(n30458) );
  XOR U27908 ( .A(n30460), .B(n30461), .Z(n27002) );
  NOR U27909 ( .A(n30462), .B(n30460), .Z(n30461) );
  XOR U27910 ( .A(n30463), .B(n30464), .Z(n27578) );
  NOR U27911 ( .A(n30465), .B(n30463), .Z(n30464) );
  XOR U27912 ( .A(n30466), .B(n30467), .Z(n27573) );
  NOR U27913 ( .A(n30468), .B(n30466), .Z(n30467) );
  XOR U27914 ( .A(n30469), .B(n30470), .Z(n27574) );
  NOR U27915 ( .A(n30471), .B(n30469), .Z(n30470) );
  XOR U27916 ( .A(n30472), .B(n30473), .Z(n26993) );
  NOR U27917 ( .A(n30474), .B(n30472), .Z(n30473) );
  XOR U27918 ( .A(n30475), .B(n30476), .Z(n27589) );
  NOR U27919 ( .A(n30477), .B(n30475), .Z(n30476) );
  XOR U27920 ( .A(n30478), .B(n30479), .Z(n27584) );
  NOR U27921 ( .A(n30480), .B(n30478), .Z(n30479) );
  XOR U27922 ( .A(n30481), .B(n30482), .Z(n27585) );
  NOR U27923 ( .A(n30483), .B(n30481), .Z(n30482) );
  XOR U27924 ( .A(n30484), .B(n30485), .Z(n26984) );
  NOR U27925 ( .A(n30486), .B(n30484), .Z(n30485) );
  XOR U27926 ( .A(n30487), .B(n30488), .Z(n26958) );
  NOR U27927 ( .A(n30489), .B(n30487), .Z(n30488) );
  XOR U27928 ( .A(n30490), .B(n30491), .Z(n26963) );
  NOR U27929 ( .A(n30492), .B(n30490), .Z(n30491) );
  IV U27930 ( .A(n26965), .Z(n29818) );
  XNOR U27931 ( .A(n30493), .B(n30494), .Z(n26965) );
  NOR U27932 ( .A(n30495), .B(n30493), .Z(n30494) );
  XOR U27933 ( .A(n30496), .B(n30497), .Z(n26975) );
  NOR U27934 ( .A(n30498), .B(n30496), .Z(n30497) );
  XOR U27935 ( .A(n30499), .B(n30500), .Z(n27595) );
  NOR U27936 ( .A(n30501), .B(n30499), .Z(n30500) );
  XOR U27937 ( .A(n30502), .B(n30503), .Z(n27598) );
  NOR U27938 ( .A(n30504), .B(n30502), .Z(n30503) );
  XOR U27939 ( .A(n30505), .B(n30506), .Z(n27601) );
  NOR U27940 ( .A(n30507), .B(n30505), .Z(n30506) );
  XOR U27941 ( .A(n30508), .B(n30509), .Z(n27604) );
  NOR U27942 ( .A(n30510), .B(n30508), .Z(n30509) );
  XOR U27943 ( .A(n30511), .B(n30512), .Z(n27607) );
  NOR U27944 ( .A(n30513), .B(n30511), .Z(n30512) );
  XOR U27945 ( .A(n30514), .B(n30515), .Z(n27610) );
  NOR U27946 ( .A(n30516), .B(n30514), .Z(n30515) );
  XOR U27947 ( .A(n30517), .B(n30518), .Z(n27613) );
  NOR U27948 ( .A(n30519), .B(n30517), .Z(n30518) );
  XOR U27949 ( .A(n30520), .B(n30521), .Z(n27616) );
  NOR U27950 ( .A(n30522), .B(n30520), .Z(n30521) );
  XOR U27951 ( .A(n30523), .B(n30524), .Z(n27619) );
  NOR U27952 ( .A(n30525), .B(n30523), .Z(n30524) );
  XOR U27953 ( .A(n30526), .B(n30527), .Z(n27622) );
  NOR U27954 ( .A(n30528), .B(n30526), .Z(n30527) );
  XOR U27955 ( .A(n30529), .B(n30530), .Z(n27625) );
  NOR U27956 ( .A(n30531), .B(n30529), .Z(n30530) );
  XOR U27957 ( .A(n30532), .B(n30533), .Z(n27628) );
  NOR U27958 ( .A(n30534), .B(n30532), .Z(n30533) );
  XOR U27959 ( .A(n30535), .B(n30536), .Z(n27631) );
  NOR U27960 ( .A(n30537), .B(n30535), .Z(n30536) );
  XOR U27961 ( .A(n30538), .B(n30539), .Z(n27634) );
  NOR U27962 ( .A(n30540), .B(n30538), .Z(n30539) );
  XOR U27963 ( .A(n30541), .B(n30542), .Z(n27637) );
  NOR U27964 ( .A(n30543), .B(n30541), .Z(n30542) );
  XOR U27965 ( .A(n30544), .B(n30545), .Z(n27640) );
  NOR U27966 ( .A(n30546), .B(n30544), .Z(n30545) );
  XOR U27967 ( .A(n30547), .B(n30548), .Z(n27643) );
  NOR U27968 ( .A(n30549), .B(n30547), .Z(n30548) );
  XOR U27969 ( .A(n30550), .B(n30551), .Z(n27646) );
  NOR U27970 ( .A(n30552), .B(n30550), .Z(n30551) );
  XOR U27971 ( .A(n30553), .B(n30554), .Z(n27649) );
  NOR U27972 ( .A(n30555), .B(n30553), .Z(n30554) );
  XOR U27973 ( .A(n30556), .B(n30557), .Z(n27652) );
  NOR U27974 ( .A(n30558), .B(n30556), .Z(n30557) );
  XOR U27975 ( .A(n30559), .B(n30560), .Z(n27655) );
  NOR U27976 ( .A(n30561), .B(n30559), .Z(n30560) );
  XOR U27977 ( .A(n30562), .B(n30563), .Z(n27658) );
  NOR U27978 ( .A(n30564), .B(n30562), .Z(n30563) );
  XOR U27979 ( .A(n30565), .B(n30566), .Z(n27661) );
  NOR U27980 ( .A(n30567), .B(n30565), .Z(n30566) );
  XOR U27981 ( .A(n30568), .B(n30569), .Z(n27664) );
  NOR U27982 ( .A(n30570), .B(n30568), .Z(n30569) );
  XOR U27983 ( .A(n30571), .B(n30572), .Z(n27667) );
  NOR U27984 ( .A(n30573), .B(n30571), .Z(n30572) );
  XOR U27985 ( .A(n30574), .B(n30575), .Z(n27670) );
  NOR U27986 ( .A(n30576), .B(n30574), .Z(n30575) );
  XOR U27987 ( .A(n30577), .B(n30578), .Z(n27673) );
  NOR U27988 ( .A(n30579), .B(n30577), .Z(n30578) );
  XOR U27989 ( .A(n30580), .B(n30581), .Z(n27676) );
  NOR U27990 ( .A(n30582), .B(n30580), .Z(n30581) );
  XOR U27991 ( .A(n30583), .B(n30584), .Z(n27679) );
  NOR U27992 ( .A(n30585), .B(n30583), .Z(n30584) );
  XOR U27993 ( .A(n30586), .B(n30587), .Z(n27682) );
  NOR U27994 ( .A(n30588), .B(n30586), .Z(n30587) );
  XOR U27995 ( .A(n30589), .B(n30590), .Z(n27685) );
  NOR U27996 ( .A(n30591), .B(n30589), .Z(n30590) );
  XOR U27997 ( .A(n30592), .B(n30593), .Z(n27688) );
  NOR U27998 ( .A(n30594), .B(n30592), .Z(n30593) );
  XOR U27999 ( .A(n30595), .B(n30596), .Z(n27691) );
  NOR U28000 ( .A(n30597), .B(n30595), .Z(n30596) );
  XOR U28001 ( .A(n30598), .B(n30599), .Z(n27694) );
  NOR U28002 ( .A(n30600), .B(n30598), .Z(n30599) );
  XOR U28003 ( .A(n30601), .B(n30602), .Z(n27697) );
  NOR U28004 ( .A(n30603), .B(n30601), .Z(n30602) );
  XOR U28005 ( .A(n30604), .B(n30605), .Z(n27700) );
  NOR U28006 ( .A(n30606), .B(n30604), .Z(n30605) );
  XOR U28007 ( .A(n30607), .B(n30608), .Z(n27703) );
  NOR U28008 ( .A(n30609), .B(n30607), .Z(n30608) );
  XOR U28009 ( .A(n30610), .B(n30611), .Z(n27706) );
  NOR U28010 ( .A(n30612), .B(n30610), .Z(n30611) );
  XOR U28011 ( .A(n30613), .B(n30614), .Z(n27709) );
  NOR U28012 ( .A(n30615), .B(n30613), .Z(n30614) );
  XOR U28013 ( .A(n30616), .B(n30617), .Z(n27712) );
  NOR U28014 ( .A(n30618), .B(n30616), .Z(n30617) );
  XOR U28015 ( .A(n30619), .B(n30620), .Z(n27715) );
  NOR U28016 ( .A(n30621), .B(n30619), .Z(n30620) );
  XOR U28017 ( .A(n30622), .B(n30623), .Z(n27718) );
  NOR U28018 ( .A(n30624), .B(n30622), .Z(n30623) );
  XOR U28019 ( .A(n30625), .B(n30626), .Z(n27721) );
  NOR U28020 ( .A(n30627), .B(n30625), .Z(n30626) );
  XOR U28021 ( .A(n30628), .B(n30629), .Z(n27724) );
  NOR U28022 ( .A(n30630), .B(n30628), .Z(n30629) );
  XOR U28023 ( .A(n30631), .B(n30632), .Z(n27727) );
  NOR U28024 ( .A(n30633), .B(n30631), .Z(n30632) );
  XOR U28025 ( .A(n30634), .B(n30635), .Z(n27730) );
  NOR U28026 ( .A(n30636), .B(n30634), .Z(n30635) );
  XOR U28027 ( .A(n30637), .B(n30638), .Z(n27733) );
  NOR U28028 ( .A(n30639), .B(n30637), .Z(n30638) );
  XOR U28029 ( .A(n30640), .B(n30641), .Z(n27736) );
  NOR U28030 ( .A(n30642), .B(n30640), .Z(n30641) );
  XOR U28031 ( .A(n30643), .B(n30644), .Z(n27739) );
  NOR U28032 ( .A(n30645), .B(n30643), .Z(n30644) );
  XOR U28033 ( .A(n30646), .B(n30647), .Z(n27742) );
  NOR U28034 ( .A(n30648), .B(n30646), .Z(n30647) );
  XOR U28035 ( .A(n30649), .B(n30650), .Z(n27745) );
  NOR U28036 ( .A(n30651), .B(n30649), .Z(n30650) );
  XOR U28037 ( .A(n30652), .B(n30653), .Z(n27748) );
  NOR U28038 ( .A(n30654), .B(n30652), .Z(n30653) );
  XOR U28039 ( .A(n30655), .B(n30656), .Z(n27751) );
  NOR U28040 ( .A(n30657), .B(n30655), .Z(n30656) );
  XOR U28041 ( .A(n30658), .B(n30659), .Z(n27754) );
  NOR U28042 ( .A(n30660), .B(n30658), .Z(n30659) );
  XOR U28043 ( .A(n30661), .B(n30662), .Z(n27757) );
  NOR U28044 ( .A(n30663), .B(n30661), .Z(n30662) );
  XOR U28045 ( .A(n30664), .B(n30665), .Z(n27760) );
  NOR U28046 ( .A(n30666), .B(n30664), .Z(n30665) );
  XOR U28047 ( .A(n30667), .B(n30668), .Z(n27763) );
  NOR U28048 ( .A(n30669), .B(n30667), .Z(n30668) );
  XOR U28049 ( .A(n30670), .B(n30671), .Z(n27766) );
  NOR U28050 ( .A(n30672), .B(n30670), .Z(n30671) );
  XOR U28051 ( .A(n30673), .B(n30674), .Z(n27769) );
  NOR U28052 ( .A(n30675), .B(n30673), .Z(n30674) );
  XOR U28053 ( .A(n30676), .B(n30677), .Z(n27772) );
  NOR U28054 ( .A(n30678), .B(n30676), .Z(n30677) );
  XOR U28055 ( .A(n30679), .B(n30680), .Z(n27775) );
  NOR U28056 ( .A(n30681), .B(n30679), .Z(n30680) );
  XOR U28057 ( .A(n30682), .B(n30683), .Z(n27778) );
  NOR U28058 ( .A(n30684), .B(n30682), .Z(n30683) );
  XOR U28059 ( .A(n30685), .B(n30686), .Z(n27781) );
  NOR U28060 ( .A(n30687), .B(n30685), .Z(n30686) );
  XOR U28061 ( .A(n30688), .B(n30689), .Z(n27784) );
  NOR U28062 ( .A(n30690), .B(n30688), .Z(n30689) );
  XOR U28063 ( .A(n30691), .B(n30692), .Z(n27787) );
  NOR U28064 ( .A(n30693), .B(n30691), .Z(n30692) );
  XOR U28065 ( .A(n30694), .B(n30695), .Z(n27790) );
  NOR U28066 ( .A(n30696), .B(n30694), .Z(n30695) );
  XOR U28067 ( .A(n30697), .B(n30698), .Z(n27793) );
  NOR U28068 ( .A(n30699), .B(n30697), .Z(n30698) );
  XOR U28069 ( .A(n30700), .B(n30701), .Z(n27796) );
  NOR U28070 ( .A(n30702), .B(n30700), .Z(n30701) );
  XOR U28071 ( .A(n30703), .B(n30704), .Z(n27799) );
  NOR U28072 ( .A(n30705), .B(n30703), .Z(n30704) );
  XOR U28073 ( .A(n30706), .B(n30707), .Z(n27802) );
  NOR U28074 ( .A(n30708), .B(n30706), .Z(n30707) );
  XOR U28075 ( .A(n30709), .B(n30710), .Z(n27805) );
  NOR U28076 ( .A(n30711), .B(n30709), .Z(n30710) );
  XOR U28077 ( .A(n30712), .B(n30713), .Z(n27808) );
  NOR U28078 ( .A(n30714), .B(n30712), .Z(n30713) );
  XOR U28079 ( .A(n30715), .B(n30716), .Z(n27811) );
  NOR U28080 ( .A(n30717), .B(n30715), .Z(n30716) );
  XOR U28081 ( .A(n30718), .B(n30719), .Z(n27814) );
  NOR U28082 ( .A(n30720), .B(n30718), .Z(n30719) );
  XOR U28083 ( .A(n30721), .B(n30722), .Z(n27817) );
  NOR U28084 ( .A(n30723), .B(n30721), .Z(n30722) );
  XOR U28085 ( .A(n30724), .B(n30725), .Z(n27820) );
  NOR U28086 ( .A(n30726), .B(n30724), .Z(n30725) );
  XOR U28087 ( .A(n30727), .B(n30728), .Z(n27823) );
  NOR U28088 ( .A(n30729), .B(n30727), .Z(n30728) );
  XOR U28089 ( .A(n30730), .B(n30731), .Z(n27826) );
  NOR U28090 ( .A(n30732), .B(n30730), .Z(n30731) );
  XOR U28091 ( .A(n30733), .B(n30734), .Z(n27829) );
  NOR U28092 ( .A(n30735), .B(n30733), .Z(n30734) );
  XOR U28093 ( .A(n30736), .B(n30737), .Z(n27832) );
  NOR U28094 ( .A(n30738), .B(n30736), .Z(n30737) );
  XOR U28095 ( .A(n30739), .B(n30740), .Z(n27835) );
  NOR U28096 ( .A(n30741), .B(n30739), .Z(n30740) );
  XOR U28097 ( .A(n30742), .B(n30743), .Z(n27838) );
  NOR U28098 ( .A(n30744), .B(n30742), .Z(n30743) );
  XOR U28099 ( .A(n30745), .B(n30746), .Z(n27841) );
  NOR U28100 ( .A(n30747), .B(n30745), .Z(n30746) );
  XOR U28101 ( .A(n30748), .B(n30749), .Z(n27844) );
  NOR U28102 ( .A(n30750), .B(n30748), .Z(n30749) );
  XOR U28103 ( .A(n30751), .B(n30752), .Z(n27847) );
  NOR U28104 ( .A(n30753), .B(n30751), .Z(n30752) );
  XOR U28105 ( .A(n30754), .B(n30755), .Z(n27850) );
  NOR U28106 ( .A(n30756), .B(n30754), .Z(n30755) );
  XOR U28107 ( .A(n30757), .B(n30758), .Z(n27853) );
  NOR U28108 ( .A(n30759), .B(n30757), .Z(n30758) );
  XOR U28109 ( .A(n30760), .B(n30761), .Z(n27856) );
  NOR U28110 ( .A(n30762), .B(n30760), .Z(n30761) );
  XOR U28111 ( .A(n30763), .B(n30764), .Z(n27859) );
  NOR U28112 ( .A(n30765), .B(n30763), .Z(n30764) );
  XOR U28113 ( .A(n30766), .B(n30767), .Z(n27862) );
  NOR U28114 ( .A(n30768), .B(n30766), .Z(n30767) );
  XOR U28115 ( .A(n30769), .B(n30770), .Z(n27865) );
  NOR U28116 ( .A(n30771), .B(n30769), .Z(n30770) );
  XOR U28117 ( .A(n30772), .B(n30773), .Z(n27868) );
  NOR U28118 ( .A(n30774), .B(n30772), .Z(n30773) );
  XOR U28119 ( .A(n30775), .B(n30776), .Z(n27871) );
  NOR U28120 ( .A(n30777), .B(n30775), .Z(n30776) );
  XOR U28121 ( .A(n30778), .B(n30779), .Z(n27874) );
  NOR U28122 ( .A(n30780), .B(n30778), .Z(n30779) );
  XOR U28123 ( .A(n30781), .B(n30782), .Z(n27877) );
  NOR U28124 ( .A(n30783), .B(n30781), .Z(n30782) );
  XOR U28125 ( .A(n30784), .B(n30785), .Z(n27880) );
  NOR U28126 ( .A(n30786), .B(n30784), .Z(n30785) );
  XOR U28127 ( .A(n30787), .B(n30788), .Z(n27883) );
  NOR U28128 ( .A(n30789), .B(n30787), .Z(n30788) );
  XOR U28129 ( .A(n30790), .B(n30791), .Z(n27886) );
  NOR U28130 ( .A(n30792), .B(n30790), .Z(n30791) );
  XOR U28131 ( .A(n30793), .B(n30794), .Z(n27889) );
  NOR U28132 ( .A(n30795), .B(n30793), .Z(n30794) );
  XOR U28133 ( .A(n30796), .B(n30797), .Z(n27892) );
  NOR U28134 ( .A(n30798), .B(n30796), .Z(n30797) );
  XOR U28135 ( .A(n30799), .B(n30800), .Z(n27895) );
  NOR U28136 ( .A(n30801), .B(n30799), .Z(n30800) );
  XOR U28137 ( .A(n30802), .B(n30803), .Z(n27898) );
  NOR U28138 ( .A(n30804), .B(n30802), .Z(n30803) );
  XOR U28139 ( .A(n30805), .B(n30806), .Z(n27901) );
  NOR U28140 ( .A(n30807), .B(n30805), .Z(n30806) );
  XOR U28141 ( .A(n30808), .B(n30809), .Z(n27904) );
  NOR U28142 ( .A(n30810), .B(n30808), .Z(n30809) );
  XOR U28143 ( .A(n30811), .B(n30812), .Z(n27907) );
  NOR U28144 ( .A(n30813), .B(n30811), .Z(n30812) );
  XOR U28145 ( .A(n30814), .B(n30815), .Z(n27910) );
  NOR U28146 ( .A(n30816), .B(n30814), .Z(n30815) );
  XOR U28147 ( .A(n30817), .B(n30818), .Z(n27913) );
  NOR U28148 ( .A(n30819), .B(n30817), .Z(n30818) );
  XOR U28149 ( .A(n30820), .B(n30821), .Z(n27916) );
  NOR U28150 ( .A(n30822), .B(n30820), .Z(n30821) );
  XOR U28151 ( .A(n30823), .B(n30824), .Z(n27919) );
  NOR U28152 ( .A(n30825), .B(n30823), .Z(n30824) );
  XOR U28153 ( .A(n30826), .B(n30827), .Z(n27922) );
  NOR U28154 ( .A(n30828), .B(n30826), .Z(n30827) );
  XOR U28155 ( .A(n30829), .B(n30830), .Z(n27925) );
  NOR U28156 ( .A(n30831), .B(n30829), .Z(n30830) );
  XOR U28157 ( .A(n30832), .B(n30833), .Z(n27928) );
  NOR U28158 ( .A(n30834), .B(n30832), .Z(n30833) );
  XOR U28159 ( .A(n30835), .B(n30836), .Z(n27931) );
  NOR U28160 ( .A(n30837), .B(n30835), .Z(n30836) );
  XOR U28161 ( .A(n30838), .B(n30839), .Z(n27934) );
  NOR U28162 ( .A(n30840), .B(n30838), .Z(n30839) );
  XOR U28163 ( .A(n30841), .B(n30842), .Z(n27937) );
  NOR U28164 ( .A(n30843), .B(n30841), .Z(n30842) );
  XOR U28165 ( .A(n30844), .B(n30845), .Z(n27940) );
  NOR U28166 ( .A(n30846), .B(n30844), .Z(n30845) );
  XOR U28167 ( .A(n30847), .B(n30848), .Z(n27943) );
  NOR U28168 ( .A(n30849), .B(n30847), .Z(n30848) );
  XOR U28169 ( .A(n30850), .B(n30851), .Z(n27946) );
  NOR U28170 ( .A(n30852), .B(n30850), .Z(n30851) );
  XOR U28171 ( .A(n30853), .B(n30854), .Z(n27949) );
  NOR U28172 ( .A(n30855), .B(n30853), .Z(n30854) );
  XOR U28173 ( .A(n30856), .B(n30857), .Z(n27952) );
  NOR U28174 ( .A(n30858), .B(n30856), .Z(n30857) );
  XOR U28175 ( .A(n30859), .B(n30860), .Z(n27955) );
  NOR U28176 ( .A(n30861), .B(n30859), .Z(n30860) );
  XOR U28177 ( .A(n30862), .B(n30863), .Z(n27958) );
  NOR U28178 ( .A(n30864), .B(n30862), .Z(n30863) );
  XOR U28179 ( .A(n30865), .B(n30866), .Z(n27961) );
  NOR U28180 ( .A(n30867), .B(n30865), .Z(n30866) );
  XOR U28181 ( .A(n30868), .B(n30869), .Z(n27964) );
  NOR U28182 ( .A(n30870), .B(n30868), .Z(n30869) );
  XOR U28183 ( .A(n30871), .B(n30872), .Z(n27967) );
  NOR U28184 ( .A(n30873), .B(n30871), .Z(n30872) );
  XOR U28185 ( .A(n30874), .B(n30875), .Z(n27970) );
  NOR U28186 ( .A(n30876), .B(n30874), .Z(n30875) );
  XOR U28187 ( .A(n30877), .B(n30878), .Z(n27973) );
  NOR U28188 ( .A(n30879), .B(n30877), .Z(n30878) );
  XOR U28189 ( .A(n30880), .B(n30881), .Z(n27976) );
  NOR U28190 ( .A(n30882), .B(n30880), .Z(n30881) );
  XOR U28191 ( .A(n30883), .B(n30884), .Z(n27979) );
  NOR U28192 ( .A(n30885), .B(n30883), .Z(n30884) );
  XOR U28193 ( .A(n30886), .B(n30887), .Z(n27982) );
  NOR U28194 ( .A(n30888), .B(n30886), .Z(n30887) );
  XOR U28195 ( .A(n30889), .B(n30890), .Z(n27985) );
  NOR U28196 ( .A(n30891), .B(n30889), .Z(n30890) );
  XOR U28197 ( .A(n30892), .B(n30893), .Z(n27988) );
  NOR U28198 ( .A(n30894), .B(n30892), .Z(n30893) );
  XOR U28199 ( .A(n30895), .B(n30896), .Z(n27991) );
  NOR U28200 ( .A(n30897), .B(n30895), .Z(n30896) );
  XOR U28201 ( .A(n30898), .B(n30899), .Z(n27994) );
  NOR U28202 ( .A(n30900), .B(n30898), .Z(n30899) );
  XOR U28203 ( .A(n30901), .B(n30902), .Z(n27997) );
  NOR U28204 ( .A(n30903), .B(n30901), .Z(n30902) );
  XOR U28205 ( .A(n30904), .B(n30905), .Z(n28000) );
  NOR U28206 ( .A(n30906), .B(n30904), .Z(n30905) );
  XOR U28207 ( .A(n30907), .B(n30908), .Z(n28003) );
  NOR U28208 ( .A(n30909), .B(n30907), .Z(n30908) );
  XOR U28209 ( .A(n30910), .B(n30911), .Z(n28006) );
  NOR U28210 ( .A(n30912), .B(n30910), .Z(n30911) );
  XOR U28211 ( .A(n30913), .B(n30914), .Z(n28009) );
  NOR U28212 ( .A(n30915), .B(n30913), .Z(n30914) );
  XOR U28213 ( .A(n30916), .B(n30917), .Z(n28012) );
  NOR U28214 ( .A(n30918), .B(n30916), .Z(n30917) );
  XOR U28215 ( .A(n30919), .B(n30920), .Z(n28015) );
  NOR U28216 ( .A(n30921), .B(n30919), .Z(n30920) );
  XOR U28217 ( .A(n30922), .B(n30923), .Z(n28018) );
  NOR U28218 ( .A(n30924), .B(n30922), .Z(n30923) );
  XOR U28219 ( .A(n30925), .B(n30926), .Z(n28021) );
  NOR U28220 ( .A(n30927), .B(n30925), .Z(n30926) );
  XOR U28221 ( .A(n30928), .B(n30929), .Z(n28024) );
  NOR U28222 ( .A(n30930), .B(n30928), .Z(n30929) );
  XOR U28223 ( .A(n30931), .B(n30932), .Z(n28027) );
  NOR U28224 ( .A(n30933), .B(n30931), .Z(n30932) );
  XOR U28225 ( .A(n30934), .B(n30935), .Z(n28030) );
  NOR U28226 ( .A(n30936), .B(n30934), .Z(n30935) );
  XOR U28227 ( .A(n30937), .B(n30938), .Z(n28033) );
  NOR U28228 ( .A(n30939), .B(n30937), .Z(n30938) );
  XOR U28229 ( .A(n30940), .B(n30941), .Z(n28036) );
  NOR U28230 ( .A(n30942), .B(n30940), .Z(n30941) );
  XOR U28231 ( .A(n30943), .B(n30944), .Z(n28039) );
  NOR U28232 ( .A(n30945), .B(n30943), .Z(n30944) );
  XOR U28233 ( .A(n30946), .B(n30947), .Z(n28042) );
  NOR U28234 ( .A(n30948), .B(n30946), .Z(n30947) );
  XOR U28235 ( .A(n30949), .B(n30950), .Z(n28045) );
  NOR U28236 ( .A(n30951), .B(n30949), .Z(n30950) );
  XOR U28237 ( .A(n30952), .B(n30953), .Z(n28048) );
  NOR U28238 ( .A(n30954), .B(n30952), .Z(n30953) );
  XOR U28239 ( .A(n30955), .B(n30956), .Z(n28051) );
  NOR U28240 ( .A(n30957), .B(n30955), .Z(n30956) );
  XOR U28241 ( .A(n30958), .B(n30959), .Z(n28054) );
  NOR U28242 ( .A(n30960), .B(n30958), .Z(n30959) );
  XOR U28243 ( .A(n30961), .B(n30962), .Z(n28057) );
  NOR U28244 ( .A(n30963), .B(n30961), .Z(n30962) );
  XOR U28245 ( .A(n30964), .B(n30965), .Z(n28060) );
  NOR U28246 ( .A(n30966), .B(n30964), .Z(n30965) );
  XOR U28247 ( .A(n30967), .B(n30968), .Z(n28063) );
  NOR U28248 ( .A(n30969), .B(n30967), .Z(n30968) );
  XOR U28249 ( .A(n30970), .B(n30971), .Z(n28066) );
  NOR U28250 ( .A(n30972), .B(n30970), .Z(n30971) );
  XOR U28251 ( .A(n30973), .B(n30974), .Z(n28069) );
  NOR U28252 ( .A(n30975), .B(n30973), .Z(n30974) );
  XOR U28253 ( .A(n30976), .B(n30977), .Z(n28072) );
  NOR U28254 ( .A(n30978), .B(n30976), .Z(n30977) );
  XOR U28255 ( .A(n30979), .B(n30980), .Z(n28075) );
  NOR U28256 ( .A(n30981), .B(n30979), .Z(n30980) );
  XOR U28257 ( .A(n30982), .B(n30983), .Z(n28078) );
  NOR U28258 ( .A(n30984), .B(n30982), .Z(n30983) );
  XOR U28259 ( .A(n30985), .B(n30986), .Z(n28081) );
  NOR U28260 ( .A(n30987), .B(n30985), .Z(n30986) );
  XOR U28261 ( .A(n30988), .B(n30989), .Z(n28084) );
  NOR U28262 ( .A(n30990), .B(n30988), .Z(n30989) );
  XOR U28263 ( .A(n30991), .B(n30992), .Z(n28087) );
  NOR U28264 ( .A(n30993), .B(n30991), .Z(n30992) );
  XOR U28265 ( .A(n30994), .B(n30995), .Z(n28090) );
  NOR U28266 ( .A(n30996), .B(n30994), .Z(n30995) );
  XOR U28267 ( .A(n30997), .B(n30998), .Z(n28093) );
  NOR U28268 ( .A(n30999), .B(n30997), .Z(n30998) );
  XOR U28269 ( .A(n31000), .B(n31001), .Z(n28096) );
  NOR U28270 ( .A(n31002), .B(n31000), .Z(n31001) );
  XOR U28271 ( .A(n31003), .B(n31004), .Z(n28099) );
  NOR U28272 ( .A(n31005), .B(n31003), .Z(n31004) );
  XOR U28273 ( .A(n31006), .B(n31007), .Z(n28102) );
  NOR U28274 ( .A(n31008), .B(n31006), .Z(n31007) );
  XOR U28275 ( .A(n31009), .B(n31010), .Z(n28105) );
  NOR U28276 ( .A(n31011), .B(n31009), .Z(n31010) );
  XOR U28277 ( .A(n31012), .B(n31013), .Z(n28108) );
  NOR U28278 ( .A(n31014), .B(n31012), .Z(n31013) );
  XOR U28279 ( .A(n31015), .B(n31016), .Z(n28111) );
  NOR U28280 ( .A(n31017), .B(n31015), .Z(n31016) );
  XOR U28281 ( .A(n31018), .B(n31019), .Z(n28114) );
  NOR U28282 ( .A(n31020), .B(n31018), .Z(n31019) );
  XOR U28283 ( .A(n31021), .B(n31022), .Z(n28117) );
  NOR U28284 ( .A(n31023), .B(n31021), .Z(n31022) );
  XOR U28285 ( .A(n31024), .B(n31025), .Z(n28120) );
  NOR U28286 ( .A(n31026), .B(n31024), .Z(n31025) );
  XOR U28287 ( .A(n31027), .B(n31028), .Z(n28123) );
  NOR U28288 ( .A(n31029), .B(n31027), .Z(n31028) );
  XOR U28289 ( .A(n31030), .B(n31031), .Z(n28126) );
  NOR U28290 ( .A(n31032), .B(n31030), .Z(n31031) );
  XOR U28291 ( .A(n31033), .B(n31034), .Z(n28129) );
  NOR U28292 ( .A(n31035), .B(n31033), .Z(n31034) );
  XOR U28293 ( .A(n31036), .B(n31037), .Z(n28132) );
  NOR U28294 ( .A(n31038), .B(n31036), .Z(n31037) );
  XOR U28295 ( .A(n31039), .B(n31040), .Z(n28135) );
  NOR U28296 ( .A(n31041), .B(n31039), .Z(n31040) );
  XOR U28297 ( .A(n31042), .B(n31043), .Z(n28138) );
  NOR U28298 ( .A(n31044), .B(n31042), .Z(n31043) );
  XOR U28299 ( .A(n31045), .B(n31046), .Z(n28141) );
  NOR U28300 ( .A(n31047), .B(n31045), .Z(n31046) );
  XOR U28301 ( .A(n31048), .B(n31049), .Z(n28144) );
  NOR U28302 ( .A(n31050), .B(n31048), .Z(n31049) );
  XOR U28303 ( .A(n31051), .B(n31052), .Z(n28147) );
  NOR U28304 ( .A(n31053), .B(n31051), .Z(n31052) );
  XOR U28305 ( .A(n31054), .B(n31055), .Z(n28150) );
  NOR U28306 ( .A(n31056), .B(n31054), .Z(n31055) );
  XOR U28307 ( .A(n31057), .B(n31058), .Z(n28153) );
  NOR U28308 ( .A(n31059), .B(n31057), .Z(n31058) );
  XOR U28309 ( .A(n31060), .B(n31061), .Z(n28156) );
  NOR U28310 ( .A(n31062), .B(n31060), .Z(n31061) );
  XOR U28311 ( .A(n31063), .B(n31064), .Z(n28159) );
  NOR U28312 ( .A(n31065), .B(n31063), .Z(n31064) );
  XOR U28313 ( .A(n31066), .B(n31067), .Z(n28162) );
  NOR U28314 ( .A(n31068), .B(n31066), .Z(n31067) );
  XOR U28315 ( .A(n31069), .B(n31070), .Z(n28165) );
  NOR U28316 ( .A(n31071), .B(n31069), .Z(n31070) );
  XOR U28317 ( .A(n31072), .B(n31073), .Z(n28168) );
  NOR U28318 ( .A(n31074), .B(n31072), .Z(n31073) );
  XOR U28319 ( .A(n31075), .B(n31076), .Z(n28171) );
  NOR U28320 ( .A(n31077), .B(n31075), .Z(n31076) );
  XOR U28321 ( .A(n31078), .B(n31079), .Z(n28174) );
  NOR U28322 ( .A(n31080), .B(n31078), .Z(n31079) );
  XOR U28323 ( .A(n31081), .B(n31082), .Z(n28177) );
  NOR U28324 ( .A(n31083), .B(n31081), .Z(n31082) );
  XOR U28325 ( .A(n31084), .B(n31085), .Z(n28180) );
  NOR U28326 ( .A(n31086), .B(n31084), .Z(n31085) );
  XOR U28327 ( .A(n31087), .B(n31088), .Z(n28183) );
  NOR U28328 ( .A(n31089), .B(n31087), .Z(n31088) );
  XOR U28329 ( .A(n31090), .B(n31091), .Z(n28186) );
  NOR U28330 ( .A(n31092), .B(n31090), .Z(n31091) );
  XOR U28331 ( .A(n31093), .B(n31094), .Z(n28189) );
  NOR U28332 ( .A(n31095), .B(n31093), .Z(n31094) );
  XOR U28333 ( .A(n31096), .B(n31097), .Z(n28192) );
  NOR U28334 ( .A(n31098), .B(n31096), .Z(n31097) );
  XOR U28335 ( .A(n31099), .B(n31100), .Z(n28195) );
  NOR U28336 ( .A(n31101), .B(n31099), .Z(n31100) );
  XOR U28337 ( .A(n31102), .B(n31103), .Z(n28198) );
  NOR U28338 ( .A(n31104), .B(n31102), .Z(n31103) );
  XOR U28339 ( .A(n31105), .B(n31106), .Z(n28201) );
  NOR U28340 ( .A(n31107), .B(n31105), .Z(n31106) );
  XOR U28341 ( .A(n31108), .B(n31109), .Z(n28204) );
  NOR U28342 ( .A(n31110), .B(n31108), .Z(n31109) );
  XOR U28343 ( .A(n31111), .B(n31112), .Z(n28207) );
  NOR U28344 ( .A(n31113), .B(n31111), .Z(n31112) );
  XOR U28345 ( .A(n31114), .B(n31115), .Z(n28210) );
  NOR U28346 ( .A(n31116), .B(n31114), .Z(n31115) );
  XOR U28347 ( .A(n31117), .B(n31118), .Z(n28213) );
  NOR U28348 ( .A(n31119), .B(n31117), .Z(n31118) );
  XOR U28349 ( .A(n31120), .B(n31121), .Z(n28216) );
  NOR U28350 ( .A(n31122), .B(n31120), .Z(n31121) );
  XOR U28351 ( .A(n31123), .B(n31124), .Z(n28219) );
  NOR U28352 ( .A(n31125), .B(n31123), .Z(n31124) );
  XOR U28353 ( .A(n31126), .B(n31127), .Z(n28222) );
  NOR U28354 ( .A(n31128), .B(n31126), .Z(n31127) );
  XOR U28355 ( .A(n31129), .B(n31130), .Z(n28225) );
  NOR U28356 ( .A(n31131), .B(n31129), .Z(n31130) );
  XOR U28357 ( .A(n31132), .B(n31133), .Z(n28228) );
  NOR U28358 ( .A(n31134), .B(n31132), .Z(n31133) );
  XOR U28359 ( .A(n31135), .B(n31136), .Z(n28231) );
  NOR U28360 ( .A(n31137), .B(n31135), .Z(n31136) );
  XOR U28361 ( .A(n31138), .B(n31139), .Z(n28234) );
  NOR U28362 ( .A(n31140), .B(n31138), .Z(n31139) );
  XOR U28363 ( .A(n31141), .B(n31142), .Z(n28237) );
  NOR U28364 ( .A(n31143), .B(n31141), .Z(n31142) );
  XOR U28365 ( .A(n31144), .B(n31145), .Z(n28240) );
  NOR U28366 ( .A(n31146), .B(n31144), .Z(n31145) );
  XOR U28367 ( .A(n31147), .B(n31148), .Z(n28243) );
  NOR U28368 ( .A(n31149), .B(n31147), .Z(n31148) );
  XOR U28369 ( .A(n31150), .B(n31151), .Z(n28246) );
  NOR U28370 ( .A(n31152), .B(n31150), .Z(n31151) );
  XOR U28371 ( .A(n31153), .B(n31154), .Z(n28249) );
  NOR U28372 ( .A(n31155), .B(n31153), .Z(n31154) );
  XOR U28373 ( .A(n31156), .B(n31157), .Z(n28252) );
  NOR U28374 ( .A(n31158), .B(n31156), .Z(n31157) );
  XOR U28375 ( .A(n31159), .B(n31160), .Z(n28255) );
  NOR U28376 ( .A(n31161), .B(n31159), .Z(n31160) );
  XOR U28377 ( .A(n31162), .B(n31163), .Z(n28258) );
  NOR U28378 ( .A(n31164), .B(n31162), .Z(n31163) );
  XOR U28379 ( .A(n31165), .B(n31166), .Z(n28261) );
  NOR U28380 ( .A(n31167), .B(n31165), .Z(n31166) );
  XOR U28381 ( .A(n31168), .B(n31169), .Z(n28264) );
  NOR U28382 ( .A(n31170), .B(n31168), .Z(n31169) );
  XOR U28383 ( .A(n31171), .B(n31172), .Z(n28267) );
  NOR U28384 ( .A(n31173), .B(n31171), .Z(n31172) );
  XOR U28385 ( .A(n31174), .B(n31175), .Z(n28270) );
  NOR U28386 ( .A(n31176), .B(n31174), .Z(n31175) );
  XOR U28387 ( .A(n31177), .B(n31178), .Z(n28273) );
  NOR U28388 ( .A(n31179), .B(n31177), .Z(n31178) );
  XOR U28389 ( .A(n31180), .B(n31181), .Z(n28276) );
  NOR U28390 ( .A(n31182), .B(n31180), .Z(n31181) );
  XOR U28391 ( .A(n31183), .B(n31184), .Z(n28279) );
  NOR U28392 ( .A(n31185), .B(n31183), .Z(n31184) );
  XOR U28393 ( .A(n31186), .B(n31187), .Z(n28282) );
  NOR U28394 ( .A(n31188), .B(n31186), .Z(n31187) );
  XOR U28395 ( .A(n31189), .B(n31190), .Z(n28285) );
  NOR U28396 ( .A(n31191), .B(n31189), .Z(n31190) );
  XOR U28397 ( .A(n31192), .B(n31193), .Z(n28288) );
  NOR U28398 ( .A(n31194), .B(n31192), .Z(n31193) );
  XOR U28399 ( .A(n31195), .B(n31196), .Z(n28291) );
  NOR U28400 ( .A(n31197), .B(n31195), .Z(n31196) );
  XOR U28401 ( .A(n31198), .B(n31199), .Z(n28294) );
  NOR U28402 ( .A(n31200), .B(n31198), .Z(n31199) );
  XOR U28403 ( .A(n31201), .B(n31202), .Z(n28297) );
  NOR U28404 ( .A(n31203), .B(n31201), .Z(n31202) );
  XOR U28405 ( .A(n31204), .B(n31205), .Z(n28300) );
  NOR U28406 ( .A(n31206), .B(n31204), .Z(n31205) );
  XOR U28407 ( .A(n31207), .B(n31208), .Z(n28303) );
  NOR U28408 ( .A(n31209), .B(n31207), .Z(n31208) );
  XOR U28409 ( .A(n31210), .B(n31211), .Z(n28306) );
  NOR U28410 ( .A(n31212), .B(n31210), .Z(n31211) );
  XOR U28411 ( .A(n31213), .B(n31214), .Z(n28309) );
  NOR U28412 ( .A(n31215), .B(n31213), .Z(n31214) );
  XOR U28413 ( .A(n31216), .B(n31217), .Z(n28312) );
  NOR U28414 ( .A(n31218), .B(n31216), .Z(n31217) );
  XOR U28415 ( .A(n31219), .B(n31220), .Z(n28315) );
  NOR U28416 ( .A(n31221), .B(n31219), .Z(n31220) );
  XOR U28417 ( .A(n31222), .B(n31223), .Z(n28318) );
  NOR U28418 ( .A(n31224), .B(n31222), .Z(n31223) );
  XOR U28419 ( .A(n31225), .B(n31226), .Z(n28321) );
  NOR U28420 ( .A(n31227), .B(n31225), .Z(n31226) );
  XOR U28421 ( .A(n31228), .B(n31229), .Z(n28324) );
  NOR U28422 ( .A(n31230), .B(n31228), .Z(n31229) );
  XOR U28423 ( .A(n31231), .B(n31232), .Z(n28327) );
  NOR U28424 ( .A(n31233), .B(n31231), .Z(n31232) );
  XOR U28425 ( .A(n31234), .B(n31235), .Z(n28330) );
  NOR U28426 ( .A(n31236), .B(n31234), .Z(n31235) );
  XOR U28427 ( .A(n31237), .B(n31238), .Z(n28333) );
  NOR U28428 ( .A(n31239), .B(n31237), .Z(n31238) );
  XOR U28429 ( .A(n31240), .B(n31241), .Z(n28336) );
  NOR U28430 ( .A(n31242), .B(n31240), .Z(n31241) );
  XOR U28431 ( .A(n31243), .B(n31244), .Z(n28339) );
  NOR U28432 ( .A(n31245), .B(n31243), .Z(n31244) );
  XOR U28433 ( .A(n31246), .B(n31247), .Z(n28342) );
  NOR U28434 ( .A(n31248), .B(n31246), .Z(n31247) );
  XOR U28435 ( .A(n31249), .B(n31250), .Z(n28345) );
  NOR U28436 ( .A(n31251), .B(n31249), .Z(n31250) );
  XOR U28437 ( .A(n31252), .B(n31253), .Z(n28348) );
  NOR U28438 ( .A(n31254), .B(n31252), .Z(n31253) );
  XOR U28439 ( .A(n31255), .B(n31256), .Z(n28351) );
  NOR U28440 ( .A(n31257), .B(n31255), .Z(n31256) );
  XOR U28441 ( .A(n31258), .B(n31259), .Z(n28354) );
  NOR U28442 ( .A(n31260), .B(n31258), .Z(n31259) );
  XOR U28443 ( .A(n31261), .B(n31262), .Z(n28357) );
  NOR U28444 ( .A(n31263), .B(n31261), .Z(n31262) );
  XNOR U28445 ( .A(n31264), .B(n31265), .Z(n28360) );
  NOR U28446 ( .A(n31266), .B(n31264), .Z(n31265) );
  XOR U28447 ( .A(n31267), .B(n31268), .Z(n28363) );
  NOR U28448 ( .A(n76), .B(n31269), .Z(n31268) );
  IV U28449 ( .A(n31267), .Z(n31269) );
  XOR U28450 ( .A(n31270), .B(n31271), .Z(n28365) );
  AND U28451 ( .A(n31272), .B(n31273), .Z(n31271) );
  XOR U28452 ( .A(n31270), .B(n79), .Z(n31273) );
  XOR U28453 ( .A(n29816), .B(n29815), .Z(n79) );
  XNOR U28454 ( .A(n29813), .B(n29812), .Z(n29815) );
  XNOR U28455 ( .A(n29810), .B(n29809), .Z(n29812) );
  XNOR U28456 ( .A(n29807), .B(n29806), .Z(n29809) );
  XNOR U28457 ( .A(n29804), .B(n29803), .Z(n29806) );
  XNOR U28458 ( .A(n29801), .B(n29800), .Z(n29803) );
  XNOR U28459 ( .A(n29798), .B(n29797), .Z(n29800) );
  XNOR U28460 ( .A(n29795), .B(n29794), .Z(n29797) );
  XNOR U28461 ( .A(n29792), .B(n29791), .Z(n29794) );
  XNOR U28462 ( .A(n29789), .B(n29788), .Z(n29791) );
  XNOR U28463 ( .A(n29786), .B(n29785), .Z(n29788) );
  XNOR U28464 ( .A(n29783), .B(n29782), .Z(n29785) );
  XNOR U28465 ( .A(n29780), .B(n29779), .Z(n29782) );
  XNOR U28466 ( .A(n29777), .B(n29776), .Z(n29779) );
  XNOR U28467 ( .A(n29774), .B(n29773), .Z(n29776) );
  XNOR U28468 ( .A(n29771), .B(n29770), .Z(n29773) );
  XNOR U28469 ( .A(n29768), .B(n29767), .Z(n29770) );
  XNOR U28470 ( .A(n29765), .B(n29764), .Z(n29767) );
  XNOR U28471 ( .A(n29762), .B(n29761), .Z(n29764) );
  XNOR U28472 ( .A(n29759), .B(n29758), .Z(n29761) );
  XNOR U28473 ( .A(n29756), .B(n29755), .Z(n29758) );
  XNOR U28474 ( .A(n29753), .B(n29752), .Z(n29755) );
  XNOR U28475 ( .A(n29750), .B(n29749), .Z(n29752) );
  XNOR U28476 ( .A(n29747), .B(n29746), .Z(n29749) );
  XNOR U28477 ( .A(n29744), .B(n29743), .Z(n29746) );
  XNOR U28478 ( .A(n29741), .B(n29740), .Z(n29743) );
  XNOR U28479 ( .A(n29738), .B(n29737), .Z(n29740) );
  XNOR U28480 ( .A(n29735), .B(n29734), .Z(n29737) );
  XNOR U28481 ( .A(n29732), .B(n29731), .Z(n29734) );
  XNOR U28482 ( .A(n29729), .B(n29728), .Z(n29731) );
  XNOR U28483 ( .A(n29726), .B(n29725), .Z(n29728) );
  XNOR U28484 ( .A(n29723), .B(n29722), .Z(n29725) );
  XNOR U28485 ( .A(n29720), .B(n29719), .Z(n29722) );
  XNOR U28486 ( .A(n29717), .B(n29716), .Z(n29719) );
  XNOR U28487 ( .A(n29714), .B(n29713), .Z(n29716) );
  XNOR U28488 ( .A(n29711), .B(n29710), .Z(n29713) );
  XNOR U28489 ( .A(n29708), .B(n29707), .Z(n29710) );
  XNOR U28490 ( .A(n29705), .B(n29704), .Z(n29707) );
  XNOR U28491 ( .A(n29702), .B(n29701), .Z(n29704) );
  XNOR U28492 ( .A(n29699), .B(n29698), .Z(n29701) );
  XNOR U28493 ( .A(n29696), .B(n29695), .Z(n29698) );
  XNOR U28494 ( .A(n29693), .B(n29692), .Z(n29695) );
  XNOR U28495 ( .A(n29690), .B(n29689), .Z(n29692) );
  XNOR U28496 ( .A(n29687), .B(n29686), .Z(n29689) );
  XNOR U28497 ( .A(n29684), .B(n29683), .Z(n29686) );
  XNOR U28498 ( .A(n29681), .B(n29680), .Z(n29683) );
  XNOR U28499 ( .A(n29678), .B(n29677), .Z(n29680) );
  XNOR U28500 ( .A(n29675), .B(n29674), .Z(n29677) );
  XNOR U28501 ( .A(n29672), .B(n29671), .Z(n29674) );
  XNOR U28502 ( .A(n29669), .B(n29668), .Z(n29671) );
  XNOR U28503 ( .A(n29666), .B(n29665), .Z(n29668) );
  XNOR U28504 ( .A(n29663), .B(n29662), .Z(n29665) );
  XNOR U28505 ( .A(n29660), .B(n29659), .Z(n29662) );
  XNOR U28506 ( .A(n29657), .B(n29656), .Z(n29659) );
  XNOR U28507 ( .A(n29654), .B(n29653), .Z(n29656) );
  XNOR U28508 ( .A(n29651), .B(n29650), .Z(n29653) );
  XNOR U28509 ( .A(n29648), .B(n29647), .Z(n29650) );
  XNOR U28510 ( .A(n29645), .B(n29644), .Z(n29647) );
  XNOR U28511 ( .A(n29642), .B(n29641), .Z(n29644) );
  XNOR U28512 ( .A(n29639), .B(n29638), .Z(n29641) );
  XNOR U28513 ( .A(n29636), .B(n29635), .Z(n29638) );
  XNOR U28514 ( .A(n29633), .B(n29632), .Z(n29635) );
  XNOR U28515 ( .A(n29630), .B(n29629), .Z(n29632) );
  XNOR U28516 ( .A(n29627), .B(n29626), .Z(n29629) );
  XNOR U28517 ( .A(n29624), .B(n29623), .Z(n29626) );
  XNOR U28518 ( .A(n29621), .B(n29620), .Z(n29623) );
  XNOR U28519 ( .A(n29618), .B(n29617), .Z(n29620) );
  XNOR U28520 ( .A(n29615), .B(n29614), .Z(n29617) );
  XNOR U28521 ( .A(n29612), .B(n29611), .Z(n29614) );
  XNOR U28522 ( .A(n29609), .B(n29608), .Z(n29611) );
  XNOR U28523 ( .A(n29606), .B(n29605), .Z(n29608) );
  XNOR U28524 ( .A(n29603), .B(n29602), .Z(n29605) );
  XNOR U28525 ( .A(n29600), .B(n29599), .Z(n29602) );
  XNOR U28526 ( .A(n29597), .B(n29596), .Z(n29599) );
  XNOR U28527 ( .A(n29594), .B(n29593), .Z(n29596) );
  XNOR U28528 ( .A(n29591), .B(n29590), .Z(n29593) );
  XNOR U28529 ( .A(n29588), .B(n29587), .Z(n29590) );
  XNOR U28530 ( .A(n29585), .B(n29584), .Z(n29587) );
  XNOR U28531 ( .A(n29582), .B(n29581), .Z(n29584) );
  XNOR U28532 ( .A(n29579), .B(n29578), .Z(n29581) );
  XNOR U28533 ( .A(n29576), .B(n29575), .Z(n29578) );
  XNOR U28534 ( .A(n29573), .B(n29572), .Z(n29575) );
  XNOR U28535 ( .A(n29570), .B(n29569), .Z(n29572) );
  XNOR U28536 ( .A(n29567), .B(n29566), .Z(n29569) );
  XNOR U28537 ( .A(n29564), .B(n29563), .Z(n29566) );
  XNOR U28538 ( .A(n29561), .B(n29560), .Z(n29563) );
  XNOR U28539 ( .A(n29558), .B(n29557), .Z(n29560) );
  XNOR U28540 ( .A(n29555), .B(n29554), .Z(n29557) );
  XNOR U28541 ( .A(n29552), .B(n29551), .Z(n29554) );
  XNOR U28542 ( .A(n29549), .B(n29548), .Z(n29551) );
  XNOR U28543 ( .A(n29546), .B(n29545), .Z(n29548) );
  XNOR U28544 ( .A(n29543), .B(n29542), .Z(n29545) );
  XNOR U28545 ( .A(n29540), .B(n29539), .Z(n29542) );
  XNOR U28546 ( .A(n29537), .B(n29536), .Z(n29539) );
  XNOR U28547 ( .A(n29534), .B(n29533), .Z(n29536) );
  XNOR U28548 ( .A(n29531), .B(n29530), .Z(n29533) );
  XNOR U28549 ( .A(n29528), .B(n29527), .Z(n29530) );
  XNOR U28550 ( .A(n29525), .B(n29524), .Z(n29527) );
  XNOR U28551 ( .A(n29522), .B(n29521), .Z(n29524) );
  XNOR U28552 ( .A(n29519), .B(n29518), .Z(n29521) );
  XNOR U28553 ( .A(n29516), .B(n29515), .Z(n29518) );
  XNOR U28554 ( .A(n29513), .B(n29512), .Z(n29515) );
  XNOR U28555 ( .A(n29510), .B(n29509), .Z(n29512) );
  XNOR U28556 ( .A(n29507), .B(n29506), .Z(n29509) );
  XNOR U28557 ( .A(n29504), .B(n29503), .Z(n29506) );
  XNOR U28558 ( .A(n29501), .B(n29500), .Z(n29503) );
  XNOR U28559 ( .A(n29498), .B(n29497), .Z(n29500) );
  XNOR U28560 ( .A(n29495), .B(n29494), .Z(n29497) );
  XNOR U28561 ( .A(n29492), .B(n29491), .Z(n29494) );
  XNOR U28562 ( .A(n29489), .B(n29488), .Z(n29491) );
  XNOR U28563 ( .A(n29486), .B(n29485), .Z(n29488) );
  XNOR U28564 ( .A(n29483), .B(n29482), .Z(n29485) );
  XNOR U28565 ( .A(n29480), .B(n29479), .Z(n29482) );
  XNOR U28566 ( .A(n29477), .B(n29476), .Z(n29479) );
  XNOR U28567 ( .A(n29474), .B(n29473), .Z(n29476) );
  XNOR U28568 ( .A(n29471), .B(n29470), .Z(n29473) );
  XNOR U28569 ( .A(n29468), .B(n29467), .Z(n29470) );
  XNOR U28570 ( .A(n29465), .B(n29464), .Z(n29467) );
  XNOR U28571 ( .A(n29462), .B(n29461), .Z(n29464) );
  XNOR U28572 ( .A(n29459), .B(n29458), .Z(n29461) );
  XNOR U28573 ( .A(n29456), .B(n29455), .Z(n29458) );
  XNOR U28574 ( .A(n29453), .B(n29452), .Z(n29455) );
  XNOR U28575 ( .A(n29450), .B(n29449), .Z(n29452) );
  XNOR U28576 ( .A(n29447), .B(n29446), .Z(n29449) );
  XNOR U28577 ( .A(n29444), .B(n29443), .Z(n29446) );
  XNOR U28578 ( .A(n29441), .B(n29440), .Z(n29443) );
  XNOR U28579 ( .A(n29438), .B(n29437), .Z(n29440) );
  XNOR U28580 ( .A(n29435), .B(n29434), .Z(n29437) );
  XNOR U28581 ( .A(n29432), .B(n29431), .Z(n29434) );
  XNOR U28582 ( .A(n29429), .B(n29428), .Z(n29431) );
  XNOR U28583 ( .A(n29426), .B(n29425), .Z(n29428) );
  XNOR U28584 ( .A(n29423), .B(n29422), .Z(n29425) );
  XNOR U28585 ( .A(n29420), .B(n29419), .Z(n29422) );
  XNOR U28586 ( .A(n29417), .B(n29416), .Z(n29419) );
  XNOR U28587 ( .A(n29414), .B(n29413), .Z(n29416) );
  XNOR U28588 ( .A(n29411), .B(n29410), .Z(n29413) );
  XNOR U28589 ( .A(n29408), .B(n29407), .Z(n29410) );
  XNOR U28590 ( .A(n29405), .B(n29404), .Z(n29407) );
  XNOR U28591 ( .A(n29402), .B(n29401), .Z(n29404) );
  XNOR U28592 ( .A(n29399), .B(n29398), .Z(n29401) );
  XNOR U28593 ( .A(n29396), .B(n29395), .Z(n29398) );
  XNOR U28594 ( .A(n29393), .B(n29392), .Z(n29395) );
  XNOR U28595 ( .A(n29390), .B(n29389), .Z(n29392) );
  XNOR U28596 ( .A(n29387), .B(n29386), .Z(n29389) );
  XNOR U28597 ( .A(n29384), .B(n29383), .Z(n29386) );
  XNOR U28598 ( .A(n29381), .B(n29380), .Z(n29383) );
  XNOR U28599 ( .A(n29378), .B(n29377), .Z(n29380) );
  XNOR U28600 ( .A(n29375), .B(n29374), .Z(n29377) );
  XNOR U28601 ( .A(n29372), .B(n29371), .Z(n29374) );
  XNOR U28602 ( .A(n29369), .B(n29368), .Z(n29371) );
  XNOR U28603 ( .A(n29366), .B(n29365), .Z(n29368) );
  XNOR U28604 ( .A(n29363), .B(n29362), .Z(n29365) );
  XNOR U28605 ( .A(n29360), .B(n29359), .Z(n29362) );
  XNOR U28606 ( .A(n29357), .B(n29356), .Z(n29359) );
  XNOR U28607 ( .A(n29354), .B(n29353), .Z(n29356) );
  XNOR U28608 ( .A(n29351), .B(n29350), .Z(n29353) );
  XNOR U28609 ( .A(n29348), .B(n29347), .Z(n29350) );
  XNOR U28610 ( .A(n29345), .B(n29344), .Z(n29347) );
  XNOR U28611 ( .A(n29342), .B(n29341), .Z(n29344) );
  XNOR U28612 ( .A(n29339), .B(n29338), .Z(n29341) );
  XNOR U28613 ( .A(n29336), .B(n29335), .Z(n29338) );
  XNOR U28614 ( .A(n29333), .B(n29332), .Z(n29335) );
  XNOR U28615 ( .A(n29330), .B(n29329), .Z(n29332) );
  XNOR U28616 ( .A(n29327), .B(n29326), .Z(n29329) );
  XNOR U28617 ( .A(n29324), .B(n29323), .Z(n29326) );
  XNOR U28618 ( .A(n29321), .B(n29320), .Z(n29323) );
  XNOR U28619 ( .A(n29318), .B(n29317), .Z(n29320) );
  XNOR U28620 ( .A(n29315), .B(n29314), .Z(n29317) );
  XNOR U28621 ( .A(n29312), .B(n29311), .Z(n29314) );
  XNOR U28622 ( .A(n29309), .B(n29308), .Z(n29311) );
  XNOR U28623 ( .A(n29306), .B(n29305), .Z(n29308) );
  XNOR U28624 ( .A(n29303), .B(n29302), .Z(n29305) );
  XNOR U28625 ( .A(n29300), .B(n29299), .Z(n29302) );
  XNOR U28626 ( .A(n29297), .B(n29296), .Z(n29299) );
  XNOR U28627 ( .A(n29294), .B(n29293), .Z(n29296) );
  XNOR U28628 ( .A(n29291), .B(n29290), .Z(n29293) );
  XNOR U28629 ( .A(n29288), .B(n29287), .Z(n29290) );
  XNOR U28630 ( .A(n29285), .B(n29284), .Z(n29287) );
  XNOR U28631 ( .A(n29282), .B(n29281), .Z(n29284) );
  XNOR U28632 ( .A(n29279), .B(n29278), .Z(n29281) );
  XNOR U28633 ( .A(n29276), .B(n29275), .Z(n29278) );
  XNOR U28634 ( .A(n29273), .B(n29272), .Z(n29275) );
  XNOR U28635 ( .A(n29270), .B(n29269), .Z(n29272) );
  XNOR U28636 ( .A(n29267), .B(n29266), .Z(n29269) );
  XNOR U28637 ( .A(n29264), .B(n29263), .Z(n29266) );
  XNOR U28638 ( .A(n29261), .B(n29260), .Z(n29263) );
  XNOR U28639 ( .A(n29258), .B(n29257), .Z(n29260) );
  XNOR U28640 ( .A(n29255), .B(n29254), .Z(n29257) );
  XNOR U28641 ( .A(n29252), .B(n29251), .Z(n29254) );
  XNOR U28642 ( .A(n29249), .B(n29248), .Z(n29251) );
  XNOR U28643 ( .A(n29246), .B(n29245), .Z(n29248) );
  XNOR U28644 ( .A(n29243), .B(n29242), .Z(n29245) );
  XNOR U28645 ( .A(n29240), .B(n29239), .Z(n29242) );
  XNOR U28646 ( .A(n29237), .B(n29236), .Z(n29239) );
  XNOR U28647 ( .A(n29234), .B(n29233), .Z(n29236) );
  XNOR U28648 ( .A(n29231), .B(n29230), .Z(n29233) );
  XNOR U28649 ( .A(n29228), .B(n29227), .Z(n29230) );
  XNOR U28650 ( .A(n29225), .B(n29224), .Z(n29227) );
  XNOR U28651 ( .A(n29222), .B(n29221), .Z(n29224) );
  XNOR U28652 ( .A(n29219), .B(n29218), .Z(n29221) );
  XNOR U28653 ( .A(n29216), .B(n29215), .Z(n29218) );
  XNOR U28654 ( .A(n29213), .B(n29212), .Z(n29215) );
  XNOR U28655 ( .A(n29210), .B(n29209), .Z(n29212) );
  XNOR U28656 ( .A(n29207), .B(n29206), .Z(n29209) );
  XNOR U28657 ( .A(n29204), .B(n29203), .Z(n29206) );
  XNOR U28658 ( .A(n29201), .B(n29200), .Z(n29203) );
  XNOR U28659 ( .A(n29198), .B(n29197), .Z(n29200) );
  XNOR U28660 ( .A(n29195), .B(n29194), .Z(n29197) );
  XNOR U28661 ( .A(n29192), .B(n29191), .Z(n29194) );
  XNOR U28662 ( .A(n29189), .B(n29188), .Z(n29191) );
  XNOR U28663 ( .A(n29186), .B(n29185), .Z(n29188) );
  XNOR U28664 ( .A(n29183), .B(n29182), .Z(n29185) );
  XNOR U28665 ( .A(n29180), .B(n29179), .Z(n29182) );
  XNOR U28666 ( .A(n29177), .B(n29176), .Z(n29179) );
  XNOR U28667 ( .A(n29174), .B(n29173), .Z(n29176) );
  XNOR U28668 ( .A(n29171), .B(n29170), .Z(n29173) );
  XNOR U28669 ( .A(n29168), .B(n29167), .Z(n29170) );
  XNOR U28670 ( .A(n29165), .B(n29164), .Z(n29167) );
  XNOR U28671 ( .A(n29162), .B(n29161), .Z(n29164) );
  XNOR U28672 ( .A(n29159), .B(n29158), .Z(n29161) );
  XNOR U28673 ( .A(n29156), .B(n29155), .Z(n29158) );
  XNOR U28674 ( .A(n29153), .B(n29152), .Z(n29155) );
  XNOR U28675 ( .A(n29150), .B(n29149), .Z(n29152) );
  XNOR U28676 ( .A(n29147), .B(n29146), .Z(n29149) );
  XNOR U28677 ( .A(n29144), .B(n29143), .Z(n29146) );
  XNOR U28678 ( .A(n29141), .B(n29140), .Z(n29143) );
  XNOR U28679 ( .A(n29138), .B(n29137), .Z(n29140) );
  XNOR U28680 ( .A(n29135), .B(n29134), .Z(n29137) );
  XNOR U28681 ( .A(n29132), .B(n29131), .Z(n29134) );
  XNOR U28682 ( .A(n29129), .B(n29128), .Z(n29131) );
  XNOR U28683 ( .A(n29126), .B(n29125), .Z(n29128) );
  XNOR U28684 ( .A(n29123), .B(n29122), .Z(n29125) );
  XNOR U28685 ( .A(n29120), .B(n29119), .Z(n29122) );
  XNOR U28686 ( .A(n29117), .B(n29116), .Z(n29119) );
  XNOR U28687 ( .A(n29114), .B(n29113), .Z(n29116) );
  XNOR U28688 ( .A(n29111), .B(n29110), .Z(n29113) );
  XNOR U28689 ( .A(n29108), .B(n29107), .Z(n29110) );
  XNOR U28690 ( .A(n29105), .B(n29104), .Z(n29107) );
  XNOR U28691 ( .A(n29102), .B(n29101), .Z(n29104) );
  XNOR U28692 ( .A(n29099), .B(n29098), .Z(n29101) );
  XNOR U28693 ( .A(n29096), .B(n29095), .Z(n29098) );
  XNOR U28694 ( .A(n29093), .B(n29092), .Z(n29095) );
  XNOR U28695 ( .A(n29090), .B(n29089), .Z(n29092) );
  XNOR U28696 ( .A(n29087), .B(n29086), .Z(n29089) );
  XNOR U28697 ( .A(n29084), .B(n29083), .Z(n29086) );
  XNOR U28698 ( .A(n29081), .B(n29080), .Z(n29083) );
  XNOR U28699 ( .A(n29078), .B(n29077), .Z(n29080) );
  XNOR U28700 ( .A(n29075), .B(n29074), .Z(n29077) );
  XNOR U28701 ( .A(n29072), .B(n29071), .Z(n29074) );
  XNOR U28702 ( .A(n29069), .B(n29068), .Z(n29071) );
  XNOR U28703 ( .A(n29066), .B(n29065), .Z(n29068) );
  XNOR U28704 ( .A(n29063), .B(n29062), .Z(n29065) );
  XNOR U28705 ( .A(n29060), .B(n29059), .Z(n29062) );
  XNOR U28706 ( .A(n29057), .B(n29056), .Z(n29059) );
  XNOR U28707 ( .A(n29054), .B(n29053), .Z(n29056) );
  XNOR U28708 ( .A(n29051), .B(n29050), .Z(n29053) );
  XNOR U28709 ( .A(n29048), .B(n29047), .Z(n29050) );
  XNOR U28710 ( .A(n29045), .B(n29044), .Z(n29047) );
  XNOR U28711 ( .A(n29042), .B(n29041), .Z(n29044) );
  XNOR U28712 ( .A(n29039), .B(n29038), .Z(n29041) );
  XNOR U28713 ( .A(n29036), .B(n29035), .Z(n29038) );
  XNOR U28714 ( .A(n29033), .B(n29032), .Z(n29035) );
  XNOR U28715 ( .A(n29030), .B(n29029), .Z(n29032) );
  XNOR U28716 ( .A(n29027), .B(n29026), .Z(n29029) );
  XNOR U28717 ( .A(n29024), .B(n29023), .Z(n29026) );
  XNOR U28718 ( .A(n29021), .B(n29020), .Z(n29023) );
  XNOR U28719 ( .A(n29018), .B(n29017), .Z(n29020) );
  XNOR U28720 ( .A(n29015), .B(n29014), .Z(n29017) );
  XNOR U28721 ( .A(n29012), .B(n29011), .Z(n29014) );
  XNOR U28722 ( .A(n29009), .B(n29008), .Z(n29011) );
  XNOR U28723 ( .A(n29006), .B(n29005), .Z(n29008) );
  XNOR U28724 ( .A(n29003), .B(n29002), .Z(n29005) );
  XNOR U28725 ( .A(n29000), .B(n28999), .Z(n29002) );
  XNOR U28726 ( .A(n28997), .B(n28996), .Z(n28999) );
  XNOR U28727 ( .A(n28994), .B(n28993), .Z(n28996) );
  XNOR U28728 ( .A(n28991), .B(n28990), .Z(n28993) );
  XNOR U28729 ( .A(n28988), .B(n28987), .Z(n28990) );
  XNOR U28730 ( .A(n28985), .B(n28984), .Z(n28987) );
  XNOR U28731 ( .A(n28982), .B(n28981), .Z(n28984) );
  XNOR U28732 ( .A(n28979), .B(n28978), .Z(n28981) );
  XNOR U28733 ( .A(n28976), .B(n28975), .Z(n28978) );
  XNOR U28734 ( .A(n28973), .B(n28972), .Z(n28975) );
  XNOR U28735 ( .A(n28970), .B(n28969), .Z(n28972) );
  XNOR U28736 ( .A(n28967), .B(n28966), .Z(n28969) );
  XNOR U28737 ( .A(n28964), .B(n28963), .Z(n28966) );
  XNOR U28738 ( .A(n28961), .B(n28960), .Z(n28963) );
  XNOR U28739 ( .A(n28958), .B(n28957), .Z(n28960) );
  XNOR U28740 ( .A(n28955), .B(n28954), .Z(n28957) );
  XNOR U28741 ( .A(n28952), .B(n28951), .Z(n28954) );
  XNOR U28742 ( .A(n28949), .B(n28948), .Z(n28951) );
  XNOR U28743 ( .A(n28946), .B(n28945), .Z(n28948) );
  XNOR U28744 ( .A(n28943), .B(n28942), .Z(n28945) );
  XNOR U28745 ( .A(n28940), .B(n28939), .Z(n28942) );
  XNOR U28746 ( .A(n28937), .B(n28936), .Z(n28939) );
  XNOR U28747 ( .A(n28934), .B(n28933), .Z(n28936) );
  XNOR U28748 ( .A(n28931), .B(n28930), .Z(n28933) );
  XNOR U28749 ( .A(n28928), .B(n28927), .Z(n28930) );
  XNOR U28750 ( .A(n28925), .B(n28924), .Z(n28927) );
  XNOR U28751 ( .A(n28922), .B(n28921), .Z(n28924) );
  XNOR U28752 ( .A(n28919), .B(n28918), .Z(n28921) );
  XNOR U28753 ( .A(n28916), .B(n28915), .Z(n28918) );
  XNOR U28754 ( .A(n28913), .B(n28912), .Z(n28915) );
  XNOR U28755 ( .A(n28910), .B(n28909), .Z(n28912) );
  XNOR U28756 ( .A(n28907), .B(n28906), .Z(n28909) );
  XNOR U28757 ( .A(n28904), .B(n28903), .Z(n28906) );
  XNOR U28758 ( .A(n28901), .B(n28900), .Z(n28903) );
  XNOR U28759 ( .A(n28898), .B(n28897), .Z(n28900) );
  XNOR U28760 ( .A(n28895), .B(n28894), .Z(n28897) );
  XNOR U28761 ( .A(n28892), .B(n28891), .Z(n28894) );
  XNOR U28762 ( .A(n28889), .B(n28888), .Z(n28891) );
  XNOR U28763 ( .A(n28886), .B(n28885), .Z(n28888) );
  XNOR U28764 ( .A(n28883), .B(n28882), .Z(n28885) );
  XNOR U28765 ( .A(n28880), .B(n28879), .Z(n28882) );
  XNOR U28766 ( .A(n28877), .B(n28876), .Z(n28879) );
  XNOR U28767 ( .A(n28874), .B(n28873), .Z(n28876) );
  XNOR U28768 ( .A(n28871), .B(n28870), .Z(n28873) );
  XNOR U28769 ( .A(n28868), .B(n28867), .Z(n28870) );
  XNOR U28770 ( .A(n28865), .B(n28864), .Z(n28867) );
  XNOR U28771 ( .A(n28862), .B(n28861), .Z(n28864) );
  XNOR U28772 ( .A(n28859), .B(n28858), .Z(n28861) );
  XNOR U28773 ( .A(n28856), .B(n28855), .Z(n28858) );
  XNOR U28774 ( .A(n28853), .B(n28852), .Z(n28855) );
  XNOR U28775 ( .A(n28850), .B(n28849), .Z(n28852) );
  XNOR U28776 ( .A(n28847), .B(n28846), .Z(n28849) );
  XNOR U28777 ( .A(n28844), .B(n28843), .Z(n28846) );
  XNOR U28778 ( .A(n28841), .B(n28840), .Z(n28843) );
  XNOR U28779 ( .A(n28838), .B(n28837), .Z(n28840) );
  XNOR U28780 ( .A(n28835), .B(n28834), .Z(n28837) );
  XNOR U28781 ( .A(n28832), .B(n28831), .Z(n28834) );
  XNOR U28782 ( .A(n28829), .B(n28828), .Z(n28831) );
  XNOR U28783 ( .A(n28826), .B(n28825), .Z(n28828) );
  XNOR U28784 ( .A(n28823), .B(n28822), .Z(n28825) );
  XNOR U28785 ( .A(n28820), .B(n28819), .Z(n28822) );
  XNOR U28786 ( .A(n28817), .B(n28816), .Z(n28819) );
  XNOR U28787 ( .A(n28814), .B(n28813), .Z(n28816) );
  XNOR U28788 ( .A(n28811), .B(n28810), .Z(n28813) );
  XNOR U28789 ( .A(n28808), .B(n28807), .Z(n28810) );
  XNOR U28790 ( .A(n28805), .B(n28804), .Z(n28807) );
  XNOR U28791 ( .A(n28802), .B(n28801), .Z(n28804) );
  XNOR U28792 ( .A(n28799), .B(n28798), .Z(n28801) );
  XNOR U28793 ( .A(n28796), .B(n28795), .Z(n28798) );
  XNOR U28794 ( .A(n28793), .B(n28792), .Z(n28795) );
  XNOR U28795 ( .A(n28790), .B(n28789), .Z(n28792) );
  XNOR U28796 ( .A(n28787), .B(n28786), .Z(n28789) );
  XNOR U28797 ( .A(n28784), .B(n28783), .Z(n28786) );
  XNOR U28798 ( .A(n28781), .B(n28780), .Z(n28783) );
  XNOR U28799 ( .A(n28778), .B(n28777), .Z(n28780) );
  XNOR U28800 ( .A(n28775), .B(n28774), .Z(n28777) );
  XNOR U28801 ( .A(n28772), .B(n28771), .Z(n28774) );
  XNOR U28802 ( .A(n28769), .B(n28768), .Z(n28771) );
  XNOR U28803 ( .A(n28766), .B(n28765), .Z(n28768) );
  XNOR U28804 ( .A(n28763), .B(n28762), .Z(n28765) );
  XNOR U28805 ( .A(n28760), .B(n28759), .Z(n28762) );
  XNOR U28806 ( .A(n28757), .B(n28756), .Z(n28759) );
  XNOR U28807 ( .A(n28754), .B(n28753), .Z(n28756) );
  XNOR U28808 ( .A(n28751), .B(n28750), .Z(n28753) );
  XNOR U28809 ( .A(n28748), .B(n28747), .Z(n28750) );
  XNOR U28810 ( .A(n28745), .B(n28744), .Z(n28747) );
  XNOR U28811 ( .A(n28742), .B(n28741), .Z(n28744) );
  XNOR U28812 ( .A(n28739), .B(n28738), .Z(n28741) );
  XNOR U28813 ( .A(n28736), .B(n28735), .Z(n28738) );
  XNOR U28814 ( .A(n28733), .B(n28732), .Z(n28735) );
  XNOR U28815 ( .A(n28730), .B(n28729), .Z(n28732) );
  XNOR U28816 ( .A(n28727), .B(n28726), .Z(n28729) );
  XNOR U28817 ( .A(n28724), .B(n28723), .Z(n28726) );
  XNOR U28818 ( .A(n28721), .B(n28720), .Z(n28723) );
  XNOR U28819 ( .A(n28718), .B(n28717), .Z(n28720) );
  XNOR U28820 ( .A(n28715), .B(n28714), .Z(n28717) );
  XNOR U28821 ( .A(n28712), .B(n28711), .Z(n28714) );
  XNOR U28822 ( .A(n28709), .B(n28708), .Z(n28711) );
  XNOR U28823 ( .A(n28706), .B(n28705), .Z(n28708) );
  XNOR U28824 ( .A(n28703), .B(n28702), .Z(n28705) );
  XNOR U28825 ( .A(n28700), .B(n28699), .Z(n28702) );
  XNOR U28826 ( .A(n28697), .B(n28696), .Z(n28699) );
  XNOR U28827 ( .A(n28694), .B(n28693), .Z(n28696) );
  XNOR U28828 ( .A(n28691), .B(n28690), .Z(n28693) );
  XNOR U28829 ( .A(n28688), .B(n28687), .Z(n28690) );
  XNOR U28830 ( .A(n28685), .B(n28684), .Z(n28687) );
  XNOR U28831 ( .A(n28682), .B(n28681), .Z(n28684) );
  XNOR U28832 ( .A(n28679), .B(n28678), .Z(n28681) );
  XNOR U28833 ( .A(n28676), .B(n28675), .Z(n28678) );
  XNOR U28834 ( .A(n28673), .B(n28672), .Z(n28675) );
  XNOR U28835 ( .A(n28670), .B(n28669), .Z(n28672) );
  XNOR U28836 ( .A(n28667), .B(n28666), .Z(n28669) );
  XOR U28837 ( .A(n28664), .B(n28381), .Z(n28666) );
  XNOR U28838 ( .A(n28382), .B(n28379), .Z(n28381) );
  XNOR U28839 ( .A(n28380), .B(n28375), .Z(n28379) );
  XOR U28840 ( .A(n28376), .B(n28396), .Z(n28375) );
  XOR U28841 ( .A(n31274), .B(n28394), .Z(n28396) );
  XNOR U28842 ( .A(n28395), .B(n28662), .Z(n28394) );
  XNOR U28843 ( .A(n28663), .B(n28661), .Z(n28662) );
  XNOR U28844 ( .A(n28391), .B(n28658), .Z(n28661) );
  XNOR U28845 ( .A(n28390), .B(n28413), .Z(n28658) );
  XNOR U28846 ( .A(n28408), .B(n28657), .Z(n28413) );
  XNOR U28847 ( .A(n28407), .B(n28652), .Z(n28657) );
  XOR U28848 ( .A(n28409), .B(n28651), .Z(n28652) );
  XOR U28849 ( .A(n28412), .B(n28648), .Z(n28651) );
  XOR U28850 ( .A(n28418), .B(n28646), .Z(n28648) );
  XOR U28851 ( .A(n28647), .B(n28643), .Z(n28646) );
  XOR U28852 ( .A(n28638), .B(n28637), .Z(n28643) );
  XOR U28853 ( .A(n28434), .B(n28636), .Z(n28637) );
  AND U28854 ( .A(n31275), .B(n31276), .Z(n28636) );
  XOR U28855 ( .A(n28635), .B(n28428), .Z(n28434) );
  AND U28856 ( .A(n31277), .B(n31278), .Z(n28428) );
  XOR U28857 ( .A(n28632), .B(n28433), .Z(n28635) );
  AND U28858 ( .A(n31279), .B(n31280), .Z(n28433) );
  XOR U28859 ( .A(n28631), .B(n28431), .Z(n28632) );
  AND U28860 ( .A(n31281), .B(n31282), .Z(n28431) );
  XNOR U28861 ( .A(n28625), .B(n28430), .Z(n28631) );
  AND U28862 ( .A(n31283), .B(n31284), .Z(n28430) );
  XNOR U28863 ( .A(n28616), .B(n28626), .Z(n28625) );
  AND U28864 ( .A(n31285), .B(n31286), .Z(n28626) );
  XOR U28865 ( .A(n28614), .B(n28615), .Z(n28616) );
  AND U28866 ( .A(n31287), .B(n31288), .Z(n28615) );
  XOR U28867 ( .A(n28621), .B(n28613), .Z(n28614) );
  AND U28868 ( .A(n31289), .B(n31290), .Z(n28613) );
  XNOR U28869 ( .A(n28588), .B(n28620), .Z(n28621) );
  AND U28870 ( .A(n31291), .B(n31292), .Z(n28620) );
  XNOR U28871 ( .A(n28610), .B(n28589), .Z(n28588) );
  AND U28872 ( .A(n31293), .B(n31294), .Z(n28589) );
  XOR U28873 ( .A(n28609), .B(n28586), .Z(n28610) );
  AND U28874 ( .A(n31295), .B(n31296), .Z(n28586) );
  XOR U28875 ( .A(n28619), .B(n28585), .Z(n28609) );
  AND U28876 ( .A(n31297), .B(n31298), .Z(n28585) );
  XNOR U28877 ( .A(n28597), .B(n28584), .Z(n28619) );
  AND U28878 ( .A(n31299), .B(n31300), .Z(n28584) );
  XNOR U28879 ( .A(n28602), .B(n28598), .Z(n28597) );
  AND U28880 ( .A(n31301), .B(n31302), .Z(n28598) );
  XOR U28881 ( .A(n28601), .B(n28595), .Z(n28602) );
  AND U28882 ( .A(n31303), .B(n31304), .Z(n28595) );
  XOR U28883 ( .A(n28581), .B(n28594), .Z(n28601) );
  AND U28884 ( .A(n31305), .B(n31306), .Z(n28594) );
  XNOR U28885 ( .A(n28552), .B(n28580), .Z(n28581) );
  AND U28886 ( .A(n31307), .B(n31308), .Z(n28580) );
  XNOR U28887 ( .A(n28575), .B(n28553), .Z(n28552) );
  AND U28888 ( .A(n31309), .B(n31310), .Z(n28553) );
  XOR U28889 ( .A(n28574), .B(n28550), .Z(n28575) );
  AND U28890 ( .A(n31311), .B(n31312), .Z(n28550) );
  XOR U28891 ( .A(n28579), .B(n28549), .Z(n28574) );
  AND U28892 ( .A(n31313), .B(n31314), .Z(n28549) );
  XNOR U28893 ( .A(n28562), .B(n28548), .Z(n28579) );
  AND U28894 ( .A(n31315), .B(n31316), .Z(n28548) );
  XNOR U28895 ( .A(n28567), .B(n28563), .Z(n28562) );
  AND U28896 ( .A(n31317), .B(n31318), .Z(n28563) );
  XOR U28897 ( .A(n28566), .B(n28560), .Z(n28567) );
  AND U28898 ( .A(n31319), .B(n31320), .Z(n28560) );
  XOR U28899 ( .A(n28576), .B(n28559), .Z(n28566) );
  AND U28900 ( .A(n31321), .B(n31322), .Z(n28559) );
  XNOR U28901 ( .A(n28459), .B(n28558), .Z(n28576) );
  AND U28902 ( .A(n31323), .B(n31324), .Z(n28558) );
  XNOR U28903 ( .A(n28541), .B(n28460), .Z(n28459) );
  AND U28904 ( .A(n31325), .B(n31326), .Z(n28460) );
  XOR U28905 ( .A(n28540), .B(n28457), .Z(n28541) );
  AND U28906 ( .A(n31327), .B(n31328), .Z(n28457) );
  XOR U28907 ( .A(n28545), .B(n28456), .Z(n28540) );
  AND U28908 ( .A(n31329), .B(n31330), .Z(n28456) );
  XNOR U28909 ( .A(n28467), .B(n28455), .Z(n28545) );
  AND U28910 ( .A(n31331), .B(n31332), .Z(n28455) );
  XNOR U28911 ( .A(n28537), .B(n28468), .Z(n28467) );
  AND U28912 ( .A(n31333), .B(n31334), .Z(n28468) );
  XOR U28913 ( .A(n28536), .B(n28465), .Z(n28537) );
  AND U28914 ( .A(n31335), .B(n31336), .Z(n28465) );
  XOR U28915 ( .A(n28544), .B(n28464), .Z(n28536) );
  AND U28916 ( .A(n31337), .B(n31338), .Z(n28464) );
  XNOR U28917 ( .A(n28477), .B(n28463), .Z(n28544) );
  AND U28918 ( .A(n31339), .B(n31340), .Z(n28463) );
  XNOR U28919 ( .A(n28484), .B(n28478), .Z(n28477) );
  AND U28920 ( .A(n31341), .B(n31342), .Z(n28478) );
  XOR U28921 ( .A(n28483), .B(n28475), .Z(n28484) );
  AND U28922 ( .A(n31343), .B(n31344), .Z(n28475) );
  XOR U28923 ( .A(n28529), .B(n28474), .Z(n28483) );
  AND U28924 ( .A(n31345), .B(n31346), .Z(n28474) );
  XNOR U28925 ( .A(n28495), .B(n28473), .Z(n28529) );
  AND U28926 ( .A(n31347), .B(n31348), .Z(n28473) );
  XNOR U28927 ( .A(n28502), .B(n28496), .Z(n28495) );
  AND U28928 ( .A(n31349), .B(n31350), .Z(n28496) );
  XOR U28929 ( .A(n28501), .B(n28493), .Z(n28502) );
  AND U28930 ( .A(n31351), .B(n31352), .Z(n28493) );
  XOR U28931 ( .A(n28528), .B(n28492), .Z(n28501) );
  AND U28932 ( .A(n31353), .B(n31354), .Z(n28492) );
  XNOR U28933 ( .A(n28513), .B(n28491), .Z(n28528) );
  AND U28934 ( .A(n31355), .B(n31356), .Z(n28491) );
  XOR U28935 ( .A(n31357), .B(n28514), .Z(n28513) );
  AND U28936 ( .A(n31358), .B(n31359), .Z(n28514) );
  XOR U28937 ( .A(n31360), .B(n31361), .Z(n31357) );
  XOR U28938 ( .A(n31362), .B(n31363), .Z(n31361) );
  XOR U28939 ( .A(n28526), .B(n28527), .Z(n31363) );
  AND U28940 ( .A(n31364), .B(n31365), .Z(n28527) );
  AND U28941 ( .A(n31366), .B(n31367), .Z(n28526) );
  XNOR U28942 ( .A(n28524), .B(n28523), .Z(n31362) );
  IV U28943 ( .A(n31368), .Z(n28523) );
  AND U28944 ( .A(n31369), .B(n31370), .Z(n31368) );
  AND U28945 ( .A(n31371), .B(n31372), .Z(n28524) );
  XOR U28946 ( .A(n31373), .B(n31374), .Z(n31360) );
  XNOR U28947 ( .A(n28509), .B(n28518), .Z(n31374) );
  IV U28948 ( .A(n28510), .Z(n28518) );
  AND U28949 ( .A(n31375), .B(n31376), .Z(n28510) );
  AND U28950 ( .A(n31377), .B(n31378), .Z(n28509) );
  XOR U28951 ( .A(n28525), .B(n28511), .Z(n31373) );
  AND U28952 ( .A(n31379), .B(n31380), .Z(n28511) );
  XNOR U28953 ( .A(n31381), .B(n31382), .Z(n28525) );
  AND U28954 ( .A(n31383), .B(n31384), .Z(n31382) );
  NOR U28955 ( .A(n31385), .B(n31386), .Z(n31384) );
  NOR U28956 ( .A(n31387), .B(n31388), .Z(n31383) );
  AND U28957 ( .A(n31389), .B(n31390), .Z(n31388) );
  AND U28958 ( .A(n31391), .B(n31392), .Z(n31381) );
  NOR U28959 ( .A(n31393), .B(n31394), .Z(n31392) );
  AND U28960 ( .A(n31386), .B(n31395), .Z(n31394) );
  AND U28961 ( .A(n31387), .B(n31396), .Z(n31393) );
  NOR U28962 ( .A(n31397), .B(n31398), .Z(n31391) );
  XOR U28963 ( .A(n31399), .B(n31400), .Z(n31398) );
  AND U28964 ( .A(n31401), .B(n31402), .Z(n31400) );
  NOR U28965 ( .A(n31403), .B(n31404), .Z(n31402) );
  NOR U28966 ( .A(n31405), .B(n31406), .Z(n31401) );
  AND U28967 ( .A(n31407), .B(n31408), .Z(n31406) );
  AND U28968 ( .A(n31409), .B(n31410), .Z(n31399) );
  NOR U28969 ( .A(n31411), .B(n31412), .Z(n31410) );
  AND U28970 ( .A(n31404), .B(n31413), .Z(n31412) );
  AND U28971 ( .A(n31405), .B(n31414), .Z(n31411) );
  NOR U28972 ( .A(n31415), .B(n31416), .Z(n31409) );
  XOR U28973 ( .A(n31417), .B(n31418), .Z(n31416) );
  AND U28974 ( .A(n31419), .B(n31420), .Z(n31418) );
  NOR U28975 ( .A(n31421), .B(n31422), .Z(n31420) );
  NOR U28976 ( .A(n31423), .B(n31424), .Z(n31419) );
  AND U28977 ( .A(n31425), .B(n31426), .Z(n31424) );
  AND U28978 ( .A(n31427), .B(n31428), .Z(n31417) );
  NOR U28979 ( .A(n31429), .B(n31430), .Z(n31428) );
  AND U28980 ( .A(n31422), .B(n31431), .Z(n31430) );
  AND U28981 ( .A(n31423), .B(n31432), .Z(n31429) );
  NOR U28982 ( .A(n31433), .B(n31434), .Z(n31427) );
  XOR U28983 ( .A(n31435), .B(n31436), .Z(n31434) );
  AND U28984 ( .A(n31437), .B(n31438), .Z(n31436) );
  NOR U28985 ( .A(n31439), .B(n31440), .Z(n31438) );
  NOR U28986 ( .A(n31441), .B(n31442), .Z(n31437) );
  AND U28987 ( .A(n31443), .B(n31444), .Z(n31442) );
  AND U28988 ( .A(n31445), .B(n31446), .Z(n31435) );
  NOR U28989 ( .A(n31447), .B(n31448), .Z(n31446) );
  AND U28990 ( .A(n31440), .B(n31449), .Z(n31448) );
  AND U28991 ( .A(n31441), .B(n31450), .Z(n31447) );
  NOR U28992 ( .A(n31451), .B(n31452), .Z(n31445) );
  AND U28993 ( .A(n31453), .B(n31454), .Z(n31452) );
  AND U28994 ( .A(n31455), .B(n31456), .Z(n31454) );
  AND U28995 ( .A(n31457), .B(n31458), .Z(n31456) );
  AND U28996 ( .A(n31459), .B(n31460), .Z(n31458) );
  NOR U28997 ( .A(n31461), .B(n31462), .Z(n31459) );
  NOR U28998 ( .A(n31463), .B(n31464), .Z(n31457) );
  AND U28999 ( .A(n31465), .B(n31466), .Z(n31455) );
  NOR U29000 ( .A(n31467), .B(n31468), .Z(n31466) );
  NOR U29001 ( .A(n31469), .B(n31470), .Z(n31465) );
  AND U29002 ( .A(n31471), .B(n31472), .Z(n31453) );
  AND U29003 ( .A(n31473), .B(n31474), .Z(n31472) );
  NOR U29004 ( .A(n31475), .B(n31476), .Z(n31474) );
  NOR U29005 ( .A(n31477), .B(n31478), .Z(n31473) );
  AND U29006 ( .A(n31479), .B(n31480), .Z(n31471) );
  NOR U29007 ( .A(n31481), .B(n31482), .Z(n31480) );
  NOR U29008 ( .A(n31483), .B(n31484), .Z(n31479) );
  AND U29009 ( .A(n31439), .B(n31485), .Z(n31451) );
  AND U29010 ( .A(n31421), .B(n31486), .Z(n31433) );
  AND U29011 ( .A(n31403), .B(n31487), .Z(n31415) );
  AND U29012 ( .A(n31385), .B(n31488), .Z(n31397) );
  XOR U29013 ( .A(n31489), .B(n31490), .Z(n28638) );
  AND U29014 ( .A(n31489), .B(n31491), .Z(n31490) );
  IV U29015 ( .A(n28639), .Z(n28647) );
  XNOR U29016 ( .A(n31492), .B(n31493), .Z(n28639) );
  AND U29017 ( .A(n31492), .B(n31494), .Z(n31493) );
  XOR U29018 ( .A(n31495), .B(n31496), .Z(n28418) );
  AND U29019 ( .A(n31495), .B(n31497), .Z(n31496) );
  XOR U29020 ( .A(n31498), .B(n31499), .Z(n28412) );
  AND U29021 ( .A(n31498), .B(n31500), .Z(n31499) );
  XNOR U29022 ( .A(n31501), .B(n31502), .Z(n28409) );
  AND U29023 ( .A(n31501), .B(n31503), .Z(n31502) );
  XNOR U29024 ( .A(n31504), .B(n31505), .Z(n28407) );
  AND U29025 ( .A(n31506), .B(n31504), .Z(n31505) );
  XOR U29026 ( .A(n31507), .B(n31508), .Z(n28408) );
  NOR U29027 ( .A(n31509), .B(n31507), .Z(n31508) );
  XOR U29028 ( .A(n31510), .B(n31511), .Z(n28390) );
  NOR U29029 ( .A(n31512), .B(n31510), .Z(n31511) );
  XOR U29030 ( .A(n31513), .B(n31514), .Z(n28391) );
  NOR U29031 ( .A(n31515), .B(n31513), .Z(n31514) );
  XOR U29032 ( .A(n31516), .B(n31517), .Z(n28663) );
  NOR U29033 ( .A(n31518), .B(n31516), .Z(n31517) );
  XOR U29034 ( .A(n31519), .B(n31520), .Z(n28395) );
  NOR U29035 ( .A(n31521), .B(n31519), .Z(n31520) );
  IV U29036 ( .A(n28374), .Z(n31274) );
  XNOR U29037 ( .A(n31522), .B(n31523), .Z(n28374) );
  NOR U29038 ( .A(n31524), .B(n31522), .Z(n31523) );
  XOR U29039 ( .A(n31525), .B(n31526), .Z(n28376) );
  NOR U29040 ( .A(n31527), .B(n31525), .Z(n31526) );
  XOR U29041 ( .A(n31528), .B(n31529), .Z(n28380) );
  NOR U29042 ( .A(n31530), .B(n31528), .Z(n31529) );
  XNOR U29043 ( .A(n31531), .B(n31532), .Z(n28382) );
  NOR U29044 ( .A(n31533), .B(n31531), .Z(n31532) );
  XOR U29045 ( .A(n31534), .B(n31535), .Z(n28664) );
  NOR U29046 ( .A(n31536), .B(n31534), .Z(n31535) );
  XOR U29047 ( .A(n31537), .B(n31538), .Z(n28667) );
  NOR U29048 ( .A(n31539), .B(n31537), .Z(n31538) );
  XOR U29049 ( .A(n31540), .B(n31541), .Z(n28670) );
  NOR U29050 ( .A(n31542), .B(n31540), .Z(n31541) );
  XOR U29051 ( .A(n31543), .B(n31544), .Z(n28673) );
  NOR U29052 ( .A(n31545), .B(n31543), .Z(n31544) );
  XOR U29053 ( .A(n31546), .B(n31547), .Z(n28676) );
  NOR U29054 ( .A(n31548), .B(n31546), .Z(n31547) );
  XOR U29055 ( .A(n31549), .B(n31550), .Z(n28679) );
  NOR U29056 ( .A(n31551), .B(n31549), .Z(n31550) );
  XOR U29057 ( .A(n31552), .B(n31553), .Z(n28682) );
  NOR U29058 ( .A(n31554), .B(n31552), .Z(n31553) );
  XOR U29059 ( .A(n31555), .B(n31556), .Z(n28685) );
  NOR U29060 ( .A(n31557), .B(n31555), .Z(n31556) );
  XOR U29061 ( .A(n31558), .B(n31559), .Z(n28688) );
  NOR U29062 ( .A(n31560), .B(n31558), .Z(n31559) );
  XOR U29063 ( .A(n31561), .B(n31562), .Z(n28691) );
  NOR U29064 ( .A(n31563), .B(n31561), .Z(n31562) );
  XOR U29065 ( .A(n31564), .B(n31565), .Z(n28694) );
  NOR U29066 ( .A(n31566), .B(n31564), .Z(n31565) );
  XOR U29067 ( .A(n31567), .B(n31568), .Z(n28697) );
  NOR U29068 ( .A(n31569), .B(n31567), .Z(n31568) );
  XOR U29069 ( .A(n31570), .B(n31571), .Z(n28700) );
  NOR U29070 ( .A(n31572), .B(n31570), .Z(n31571) );
  XOR U29071 ( .A(n31573), .B(n31574), .Z(n28703) );
  NOR U29072 ( .A(n31575), .B(n31573), .Z(n31574) );
  XOR U29073 ( .A(n31576), .B(n31577), .Z(n28706) );
  NOR U29074 ( .A(n31578), .B(n31576), .Z(n31577) );
  XOR U29075 ( .A(n31579), .B(n31580), .Z(n28709) );
  NOR U29076 ( .A(n31581), .B(n31579), .Z(n31580) );
  XOR U29077 ( .A(n31582), .B(n31583), .Z(n28712) );
  NOR U29078 ( .A(n31584), .B(n31582), .Z(n31583) );
  XOR U29079 ( .A(n31585), .B(n31586), .Z(n28715) );
  NOR U29080 ( .A(n31587), .B(n31585), .Z(n31586) );
  XOR U29081 ( .A(n31588), .B(n31589), .Z(n28718) );
  NOR U29082 ( .A(n31590), .B(n31588), .Z(n31589) );
  XOR U29083 ( .A(n31591), .B(n31592), .Z(n28721) );
  NOR U29084 ( .A(n31593), .B(n31591), .Z(n31592) );
  XOR U29085 ( .A(n31594), .B(n31595), .Z(n28724) );
  NOR U29086 ( .A(n31596), .B(n31594), .Z(n31595) );
  XOR U29087 ( .A(n31597), .B(n31598), .Z(n28727) );
  NOR U29088 ( .A(n31599), .B(n31597), .Z(n31598) );
  XOR U29089 ( .A(n31600), .B(n31601), .Z(n28730) );
  NOR U29090 ( .A(n31602), .B(n31600), .Z(n31601) );
  XOR U29091 ( .A(n31603), .B(n31604), .Z(n28733) );
  NOR U29092 ( .A(n31605), .B(n31603), .Z(n31604) );
  XOR U29093 ( .A(n31606), .B(n31607), .Z(n28736) );
  NOR U29094 ( .A(n31608), .B(n31606), .Z(n31607) );
  XOR U29095 ( .A(n31609), .B(n31610), .Z(n28739) );
  NOR U29096 ( .A(n31611), .B(n31609), .Z(n31610) );
  XOR U29097 ( .A(n31612), .B(n31613), .Z(n28742) );
  NOR U29098 ( .A(n31614), .B(n31612), .Z(n31613) );
  XOR U29099 ( .A(n31615), .B(n31616), .Z(n28745) );
  NOR U29100 ( .A(n31617), .B(n31615), .Z(n31616) );
  XOR U29101 ( .A(n31618), .B(n31619), .Z(n28748) );
  NOR U29102 ( .A(n31620), .B(n31618), .Z(n31619) );
  XOR U29103 ( .A(n31621), .B(n31622), .Z(n28751) );
  NOR U29104 ( .A(n31623), .B(n31621), .Z(n31622) );
  XOR U29105 ( .A(n31624), .B(n31625), .Z(n28754) );
  NOR U29106 ( .A(n31626), .B(n31624), .Z(n31625) );
  XOR U29107 ( .A(n31627), .B(n31628), .Z(n28757) );
  NOR U29108 ( .A(n31629), .B(n31627), .Z(n31628) );
  XOR U29109 ( .A(n31630), .B(n31631), .Z(n28760) );
  NOR U29110 ( .A(n31632), .B(n31630), .Z(n31631) );
  XOR U29111 ( .A(n31633), .B(n31634), .Z(n28763) );
  NOR U29112 ( .A(n31635), .B(n31633), .Z(n31634) );
  XOR U29113 ( .A(n31636), .B(n31637), .Z(n28766) );
  NOR U29114 ( .A(n31638), .B(n31636), .Z(n31637) );
  XOR U29115 ( .A(n31639), .B(n31640), .Z(n28769) );
  NOR U29116 ( .A(n31641), .B(n31639), .Z(n31640) );
  XOR U29117 ( .A(n31642), .B(n31643), .Z(n28772) );
  NOR U29118 ( .A(n31644), .B(n31642), .Z(n31643) );
  XOR U29119 ( .A(n31645), .B(n31646), .Z(n28775) );
  NOR U29120 ( .A(n31647), .B(n31645), .Z(n31646) );
  XOR U29121 ( .A(n31648), .B(n31649), .Z(n28778) );
  NOR U29122 ( .A(n31650), .B(n31648), .Z(n31649) );
  XOR U29123 ( .A(n31651), .B(n31652), .Z(n28781) );
  NOR U29124 ( .A(n31653), .B(n31651), .Z(n31652) );
  XOR U29125 ( .A(n31654), .B(n31655), .Z(n28784) );
  NOR U29126 ( .A(n31656), .B(n31654), .Z(n31655) );
  XOR U29127 ( .A(n31657), .B(n31658), .Z(n28787) );
  NOR U29128 ( .A(n31659), .B(n31657), .Z(n31658) );
  XOR U29129 ( .A(n31660), .B(n31661), .Z(n28790) );
  NOR U29130 ( .A(n31662), .B(n31660), .Z(n31661) );
  XOR U29131 ( .A(n31663), .B(n31664), .Z(n28793) );
  NOR U29132 ( .A(n31665), .B(n31663), .Z(n31664) );
  XOR U29133 ( .A(n31666), .B(n31667), .Z(n28796) );
  NOR U29134 ( .A(n31668), .B(n31666), .Z(n31667) );
  XOR U29135 ( .A(n31669), .B(n31670), .Z(n28799) );
  NOR U29136 ( .A(n31671), .B(n31669), .Z(n31670) );
  XOR U29137 ( .A(n31672), .B(n31673), .Z(n28802) );
  NOR U29138 ( .A(n31674), .B(n31672), .Z(n31673) );
  XOR U29139 ( .A(n31675), .B(n31676), .Z(n28805) );
  NOR U29140 ( .A(n31677), .B(n31675), .Z(n31676) );
  XOR U29141 ( .A(n31678), .B(n31679), .Z(n28808) );
  NOR U29142 ( .A(n31680), .B(n31678), .Z(n31679) );
  XOR U29143 ( .A(n31681), .B(n31682), .Z(n28811) );
  NOR U29144 ( .A(n31683), .B(n31681), .Z(n31682) );
  XOR U29145 ( .A(n31684), .B(n31685), .Z(n28814) );
  NOR U29146 ( .A(n31686), .B(n31684), .Z(n31685) );
  XOR U29147 ( .A(n31687), .B(n31688), .Z(n28817) );
  NOR U29148 ( .A(n31689), .B(n31687), .Z(n31688) );
  XOR U29149 ( .A(n31690), .B(n31691), .Z(n28820) );
  NOR U29150 ( .A(n31692), .B(n31690), .Z(n31691) );
  XOR U29151 ( .A(n31693), .B(n31694), .Z(n28823) );
  NOR U29152 ( .A(n31695), .B(n31693), .Z(n31694) );
  XOR U29153 ( .A(n31696), .B(n31697), .Z(n28826) );
  NOR U29154 ( .A(n31698), .B(n31696), .Z(n31697) );
  XOR U29155 ( .A(n31699), .B(n31700), .Z(n28829) );
  NOR U29156 ( .A(n31701), .B(n31699), .Z(n31700) );
  XOR U29157 ( .A(n31702), .B(n31703), .Z(n28832) );
  NOR U29158 ( .A(n31704), .B(n31702), .Z(n31703) );
  XOR U29159 ( .A(n31705), .B(n31706), .Z(n28835) );
  NOR U29160 ( .A(n31707), .B(n31705), .Z(n31706) );
  XOR U29161 ( .A(n31708), .B(n31709), .Z(n28838) );
  NOR U29162 ( .A(n31710), .B(n31708), .Z(n31709) );
  XOR U29163 ( .A(n31711), .B(n31712), .Z(n28841) );
  NOR U29164 ( .A(n31713), .B(n31711), .Z(n31712) );
  XOR U29165 ( .A(n31714), .B(n31715), .Z(n28844) );
  NOR U29166 ( .A(n31716), .B(n31714), .Z(n31715) );
  XOR U29167 ( .A(n31717), .B(n31718), .Z(n28847) );
  NOR U29168 ( .A(n31719), .B(n31717), .Z(n31718) );
  XOR U29169 ( .A(n31720), .B(n31721), .Z(n28850) );
  NOR U29170 ( .A(n31722), .B(n31720), .Z(n31721) );
  XOR U29171 ( .A(n31723), .B(n31724), .Z(n28853) );
  NOR U29172 ( .A(n31725), .B(n31723), .Z(n31724) );
  XOR U29173 ( .A(n31726), .B(n31727), .Z(n28856) );
  NOR U29174 ( .A(n31728), .B(n31726), .Z(n31727) );
  XOR U29175 ( .A(n31729), .B(n31730), .Z(n28859) );
  NOR U29176 ( .A(n31731), .B(n31729), .Z(n31730) );
  XOR U29177 ( .A(n31732), .B(n31733), .Z(n28862) );
  NOR U29178 ( .A(n31734), .B(n31732), .Z(n31733) );
  XOR U29179 ( .A(n31735), .B(n31736), .Z(n28865) );
  NOR U29180 ( .A(n31737), .B(n31735), .Z(n31736) );
  XOR U29181 ( .A(n31738), .B(n31739), .Z(n28868) );
  NOR U29182 ( .A(n31740), .B(n31738), .Z(n31739) );
  XOR U29183 ( .A(n31741), .B(n31742), .Z(n28871) );
  NOR U29184 ( .A(n31743), .B(n31741), .Z(n31742) );
  XOR U29185 ( .A(n31744), .B(n31745), .Z(n28874) );
  NOR U29186 ( .A(n31746), .B(n31744), .Z(n31745) );
  XOR U29187 ( .A(n31747), .B(n31748), .Z(n28877) );
  NOR U29188 ( .A(n31749), .B(n31747), .Z(n31748) );
  XOR U29189 ( .A(n31750), .B(n31751), .Z(n28880) );
  NOR U29190 ( .A(n31752), .B(n31750), .Z(n31751) );
  XOR U29191 ( .A(n31753), .B(n31754), .Z(n28883) );
  NOR U29192 ( .A(n31755), .B(n31753), .Z(n31754) );
  XOR U29193 ( .A(n31756), .B(n31757), .Z(n28886) );
  NOR U29194 ( .A(n31758), .B(n31756), .Z(n31757) );
  XOR U29195 ( .A(n31759), .B(n31760), .Z(n28889) );
  NOR U29196 ( .A(n31761), .B(n31759), .Z(n31760) );
  XOR U29197 ( .A(n31762), .B(n31763), .Z(n28892) );
  NOR U29198 ( .A(n31764), .B(n31762), .Z(n31763) );
  XOR U29199 ( .A(n31765), .B(n31766), .Z(n28895) );
  NOR U29200 ( .A(n31767), .B(n31765), .Z(n31766) );
  XOR U29201 ( .A(n31768), .B(n31769), .Z(n28898) );
  NOR U29202 ( .A(n31770), .B(n31768), .Z(n31769) );
  XOR U29203 ( .A(n31771), .B(n31772), .Z(n28901) );
  NOR U29204 ( .A(n31773), .B(n31771), .Z(n31772) );
  XOR U29205 ( .A(n31774), .B(n31775), .Z(n28904) );
  NOR U29206 ( .A(n31776), .B(n31774), .Z(n31775) );
  XOR U29207 ( .A(n31777), .B(n31778), .Z(n28907) );
  NOR U29208 ( .A(n31779), .B(n31777), .Z(n31778) );
  XOR U29209 ( .A(n31780), .B(n31781), .Z(n28910) );
  NOR U29210 ( .A(n31782), .B(n31780), .Z(n31781) );
  XOR U29211 ( .A(n31783), .B(n31784), .Z(n28913) );
  NOR U29212 ( .A(n31785), .B(n31783), .Z(n31784) );
  XOR U29213 ( .A(n31786), .B(n31787), .Z(n28916) );
  NOR U29214 ( .A(n31788), .B(n31786), .Z(n31787) );
  XOR U29215 ( .A(n31789), .B(n31790), .Z(n28919) );
  NOR U29216 ( .A(n31791), .B(n31789), .Z(n31790) );
  XOR U29217 ( .A(n31792), .B(n31793), .Z(n28922) );
  NOR U29218 ( .A(n31794), .B(n31792), .Z(n31793) );
  XOR U29219 ( .A(n31795), .B(n31796), .Z(n28925) );
  NOR U29220 ( .A(n31797), .B(n31795), .Z(n31796) );
  XOR U29221 ( .A(n31798), .B(n31799), .Z(n28928) );
  NOR U29222 ( .A(n31800), .B(n31798), .Z(n31799) );
  XOR U29223 ( .A(n31801), .B(n31802), .Z(n28931) );
  NOR U29224 ( .A(n31803), .B(n31801), .Z(n31802) );
  XOR U29225 ( .A(n31804), .B(n31805), .Z(n28934) );
  NOR U29226 ( .A(n31806), .B(n31804), .Z(n31805) );
  XOR U29227 ( .A(n31807), .B(n31808), .Z(n28937) );
  NOR U29228 ( .A(n31809), .B(n31807), .Z(n31808) );
  XOR U29229 ( .A(n31810), .B(n31811), .Z(n28940) );
  NOR U29230 ( .A(n31812), .B(n31810), .Z(n31811) );
  XOR U29231 ( .A(n31813), .B(n31814), .Z(n28943) );
  NOR U29232 ( .A(n31815), .B(n31813), .Z(n31814) );
  XOR U29233 ( .A(n31816), .B(n31817), .Z(n28946) );
  NOR U29234 ( .A(n31818), .B(n31816), .Z(n31817) );
  XOR U29235 ( .A(n31819), .B(n31820), .Z(n28949) );
  NOR U29236 ( .A(n31821), .B(n31819), .Z(n31820) );
  XOR U29237 ( .A(n31822), .B(n31823), .Z(n28952) );
  NOR U29238 ( .A(n31824), .B(n31822), .Z(n31823) );
  XOR U29239 ( .A(n31825), .B(n31826), .Z(n28955) );
  NOR U29240 ( .A(n31827), .B(n31825), .Z(n31826) );
  XOR U29241 ( .A(n31828), .B(n31829), .Z(n28958) );
  NOR U29242 ( .A(n31830), .B(n31828), .Z(n31829) );
  XOR U29243 ( .A(n31831), .B(n31832), .Z(n28961) );
  NOR U29244 ( .A(n31833), .B(n31831), .Z(n31832) );
  XOR U29245 ( .A(n31834), .B(n31835), .Z(n28964) );
  NOR U29246 ( .A(n31836), .B(n31834), .Z(n31835) );
  XOR U29247 ( .A(n31837), .B(n31838), .Z(n28967) );
  NOR U29248 ( .A(n31839), .B(n31837), .Z(n31838) );
  XOR U29249 ( .A(n31840), .B(n31841), .Z(n28970) );
  NOR U29250 ( .A(n31842), .B(n31840), .Z(n31841) );
  XOR U29251 ( .A(n31843), .B(n31844), .Z(n28973) );
  NOR U29252 ( .A(n31845), .B(n31843), .Z(n31844) );
  XOR U29253 ( .A(n31846), .B(n31847), .Z(n28976) );
  NOR U29254 ( .A(n31848), .B(n31846), .Z(n31847) );
  XOR U29255 ( .A(n31849), .B(n31850), .Z(n28979) );
  NOR U29256 ( .A(n31851), .B(n31849), .Z(n31850) );
  XOR U29257 ( .A(n31852), .B(n31853), .Z(n28982) );
  NOR U29258 ( .A(n31854), .B(n31852), .Z(n31853) );
  XOR U29259 ( .A(n31855), .B(n31856), .Z(n28985) );
  NOR U29260 ( .A(n31857), .B(n31855), .Z(n31856) );
  XOR U29261 ( .A(n31858), .B(n31859), .Z(n28988) );
  NOR U29262 ( .A(n31860), .B(n31858), .Z(n31859) );
  XOR U29263 ( .A(n31861), .B(n31862), .Z(n28991) );
  NOR U29264 ( .A(n31863), .B(n31861), .Z(n31862) );
  XOR U29265 ( .A(n31864), .B(n31865), .Z(n28994) );
  NOR U29266 ( .A(n31866), .B(n31864), .Z(n31865) );
  XOR U29267 ( .A(n31867), .B(n31868), .Z(n28997) );
  NOR U29268 ( .A(n31869), .B(n31867), .Z(n31868) );
  XOR U29269 ( .A(n31870), .B(n31871), .Z(n29000) );
  NOR U29270 ( .A(n31872), .B(n31870), .Z(n31871) );
  XOR U29271 ( .A(n31873), .B(n31874), .Z(n29003) );
  NOR U29272 ( .A(n31875), .B(n31873), .Z(n31874) );
  XOR U29273 ( .A(n31876), .B(n31877), .Z(n29006) );
  NOR U29274 ( .A(n31878), .B(n31876), .Z(n31877) );
  XOR U29275 ( .A(n31879), .B(n31880), .Z(n29009) );
  NOR U29276 ( .A(n31881), .B(n31879), .Z(n31880) );
  XOR U29277 ( .A(n31882), .B(n31883), .Z(n29012) );
  NOR U29278 ( .A(n31884), .B(n31882), .Z(n31883) );
  XOR U29279 ( .A(n31885), .B(n31886), .Z(n29015) );
  NOR U29280 ( .A(n31887), .B(n31885), .Z(n31886) );
  XOR U29281 ( .A(n31888), .B(n31889), .Z(n29018) );
  NOR U29282 ( .A(n31890), .B(n31888), .Z(n31889) );
  XOR U29283 ( .A(n31891), .B(n31892), .Z(n29021) );
  NOR U29284 ( .A(n31893), .B(n31891), .Z(n31892) );
  XOR U29285 ( .A(n31894), .B(n31895), .Z(n29024) );
  NOR U29286 ( .A(n31896), .B(n31894), .Z(n31895) );
  XOR U29287 ( .A(n31897), .B(n31898), .Z(n29027) );
  NOR U29288 ( .A(n31899), .B(n31897), .Z(n31898) );
  XOR U29289 ( .A(n31900), .B(n31901), .Z(n29030) );
  NOR U29290 ( .A(n31902), .B(n31900), .Z(n31901) );
  XOR U29291 ( .A(n31903), .B(n31904), .Z(n29033) );
  NOR U29292 ( .A(n31905), .B(n31903), .Z(n31904) );
  XOR U29293 ( .A(n31906), .B(n31907), .Z(n29036) );
  NOR U29294 ( .A(n31908), .B(n31906), .Z(n31907) );
  XOR U29295 ( .A(n31909), .B(n31910), .Z(n29039) );
  NOR U29296 ( .A(n31911), .B(n31909), .Z(n31910) );
  XOR U29297 ( .A(n31912), .B(n31913), .Z(n29042) );
  NOR U29298 ( .A(n31914), .B(n31912), .Z(n31913) );
  XOR U29299 ( .A(n31915), .B(n31916), .Z(n29045) );
  NOR U29300 ( .A(n31917), .B(n31915), .Z(n31916) );
  XOR U29301 ( .A(n31918), .B(n31919), .Z(n29048) );
  NOR U29302 ( .A(n31920), .B(n31918), .Z(n31919) );
  XOR U29303 ( .A(n31921), .B(n31922), .Z(n29051) );
  NOR U29304 ( .A(n31923), .B(n31921), .Z(n31922) );
  XOR U29305 ( .A(n31924), .B(n31925), .Z(n29054) );
  NOR U29306 ( .A(n31926), .B(n31924), .Z(n31925) );
  XOR U29307 ( .A(n31927), .B(n31928), .Z(n29057) );
  NOR U29308 ( .A(n31929), .B(n31927), .Z(n31928) );
  XOR U29309 ( .A(n31930), .B(n31931), .Z(n29060) );
  NOR U29310 ( .A(n31932), .B(n31930), .Z(n31931) );
  XOR U29311 ( .A(n31933), .B(n31934), .Z(n29063) );
  NOR U29312 ( .A(n31935), .B(n31933), .Z(n31934) );
  XOR U29313 ( .A(n31936), .B(n31937), .Z(n29066) );
  NOR U29314 ( .A(n31938), .B(n31936), .Z(n31937) );
  XOR U29315 ( .A(n31939), .B(n31940), .Z(n29069) );
  NOR U29316 ( .A(n31941), .B(n31939), .Z(n31940) );
  XOR U29317 ( .A(n31942), .B(n31943), .Z(n29072) );
  NOR U29318 ( .A(n31944), .B(n31942), .Z(n31943) );
  XOR U29319 ( .A(n31945), .B(n31946), .Z(n29075) );
  NOR U29320 ( .A(n31947), .B(n31945), .Z(n31946) );
  XOR U29321 ( .A(n31948), .B(n31949), .Z(n29078) );
  NOR U29322 ( .A(n31950), .B(n31948), .Z(n31949) );
  XOR U29323 ( .A(n31951), .B(n31952), .Z(n29081) );
  NOR U29324 ( .A(n31953), .B(n31951), .Z(n31952) );
  XOR U29325 ( .A(n31954), .B(n31955), .Z(n29084) );
  NOR U29326 ( .A(n31956), .B(n31954), .Z(n31955) );
  XOR U29327 ( .A(n31957), .B(n31958), .Z(n29087) );
  NOR U29328 ( .A(n31959), .B(n31957), .Z(n31958) );
  XOR U29329 ( .A(n31960), .B(n31961), .Z(n29090) );
  NOR U29330 ( .A(n31962), .B(n31960), .Z(n31961) );
  XOR U29331 ( .A(n31963), .B(n31964), .Z(n29093) );
  NOR U29332 ( .A(n31965), .B(n31963), .Z(n31964) );
  XOR U29333 ( .A(n31966), .B(n31967), .Z(n29096) );
  NOR U29334 ( .A(n31968), .B(n31966), .Z(n31967) );
  XOR U29335 ( .A(n31969), .B(n31970), .Z(n29099) );
  NOR U29336 ( .A(n31971), .B(n31969), .Z(n31970) );
  XOR U29337 ( .A(n31972), .B(n31973), .Z(n29102) );
  NOR U29338 ( .A(n31974), .B(n31972), .Z(n31973) );
  XOR U29339 ( .A(n31975), .B(n31976), .Z(n29105) );
  NOR U29340 ( .A(n31977), .B(n31975), .Z(n31976) );
  XOR U29341 ( .A(n31978), .B(n31979), .Z(n29108) );
  NOR U29342 ( .A(n31980), .B(n31978), .Z(n31979) );
  XOR U29343 ( .A(n31981), .B(n31982), .Z(n29111) );
  NOR U29344 ( .A(n31983), .B(n31981), .Z(n31982) );
  XOR U29345 ( .A(n31984), .B(n31985), .Z(n29114) );
  NOR U29346 ( .A(n31986), .B(n31984), .Z(n31985) );
  XOR U29347 ( .A(n31987), .B(n31988), .Z(n29117) );
  NOR U29348 ( .A(n31989), .B(n31987), .Z(n31988) );
  XOR U29349 ( .A(n31990), .B(n31991), .Z(n29120) );
  NOR U29350 ( .A(n31992), .B(n31990), .Z(n31991) );
  XOR U29351 ( .A(n31993), .B(n31994), .Z(n29123) );
  NOR U29352 ( .A(n31995), .B(n31993), .Z(n31994) );
  XOR U29353 ( .A(n31996), .B(n31997), .Z(n29126) );
  NOR U29354 ( .A(n31998), .B(n31996), .Z(n31997) );
  XOR U29355 ( .A(n31999), .B(n32000), .Z(n29129) );
  NOR U29356 ( .A(n32001), .B(n31999), .Z(n32000) );
  XOR U29357 ( .A(n32002), .B(n32003), .Z(n29132) );
  NOR U29358 ( .A(n32004), .B(n32002), .Z(n32003) );
  XOR U29359 ( .A(n32005), .B(n32006), .Z(n29135) );
  NOR U29360 ( .A(n32007), .B(n32005), .Z(n32006) );
  XOR U29361 ( .A(n32008), .B(n32009), .Z(n29138) );
  NOR U29362 ( .A(n32010), .B(n32008), .Z(n32009) );
  XOR U29363 ( .A(n32011), .B(n32012), .Z(n29141) );
  NOR U29364 ( .A(n32013), .B(n32011), .Z(n32012) );
  XOR U29365 ( .A(n32014), .B(n32015), .Z(n29144) );
  NOR U29366 ( .A(n32016), .B(n32014), .Z(n32015) );
  XOR U29367 ( .A(n32017), .B(n32018), .Z(n29147) );
  NOR U29368 ( .A(n32019), .B(n32017), .Z(n32018) );
  XOR U29369 ( .A(n32020), .B(n32021), .Z(n29150) );
  NOR U29370 ( .A(n32022), .B(n32020), .Z(n32021) );
  XOR U29371 ( .A(n32023), .B(n32024), .Z(n29153) );
  NOR U29372 ( .A(n32025), .B(n32023), .Z(n32024) );
  XOR U29373 ( .A(n32026), .B(n32027), .Z(n29156) );
  NOR U29374 ( .A(n32028), .B(n32026), .Z(n32027) );
  XOR U29375 ( .A(n32029), .B(n32030), .Z(n29159) );
  NOR U29376 ( .A(n32031), .B(n32029), .Z(n32030) );
  XOR U29377 ( .A(n32032), .B(n32033), .Z(n29162) );
  NOR U29378 ( .A(n32034), .B(n32032), .Z(n32033) );
  XOR U29379 ( .A(n32035), .B(n32036), .Z(n29165) );
  NOR U29380 ( .A(n32037), .B(n32035), .Z(n32036) );
  XOR U29381 ( .A(n32038), .B(n32039), .Z(n29168) );
  NOR U29382 ( .A(n32040), .B(n32038), .Z(n32039) );
  XOR U29383 ( .A(n32041), .B(n32042), .Z(n29171) );
  NOR U29384 ( .A(n32043), .B(n32041), .Z(n32042) );
  XOR U29385 ( .A(n32044), .B(n32045), .Z(n29174) );
  NOR U29386 ( .A(n32046), .B(n32044), .Z(n32045) );
  XOR U29387 ( .A(n32047), .B(n32048), .Z(n29177) );
  NOR U29388 ( .A(n32049), .B(n32047), .Z(n32048) );
  XOR U29389 ( .A(n32050), .B(n32051), .Z(n29180) );
  NOR U29390 ( .A(n32052), .B(n32050), .Z(n32051) );
  XOR U29391 ( .A(n32053), .B(n32054), .Z(n29183) );
  NOR U29392 ( .A(n32055), .B(n32053), .Z(n32054) );
  XOR U29393 ( .A(n32056), .B(n32057), .Z(n29186) );
  NOR U29394 ( .A(n32058), .B(n32056), .Z(n32057) );
  XOR U29395 ( .A(n32059), .B(n32060), .Z(n29189) );
  NOR U29396 ( .A(n32061), .B(n32059), .Z(n32060) );
  XOR U29397 ( .A(n32062), .B(n32063), .Z(n29192) );
  NOR U29398 ( .A(n32064), .B(n32062), .Z(n32063) );
  XOR U29399 ( .A(n32065), .B(n32066), .Z(n29195) );
  NOR U29400 ( .A(n32067), .B(n32065), .Z(n32066) );
  XOR U29401 ( .A(n32068), .B(n32069), .Z(n29198) );
  NOR U29402 ( .A(n32070), .B(n32068), .Z(n32069) );
  XOR U29403 ( .A(n32071), .B(n32072), .Z(n29201) );
  NOR U29404 ( .A(n32073), .B(n32071), .Z(n32072) );
  XOR U29405 ( .A(n32074), .B(n32075), .Z(n29204) );
  NOR U29406 ( .A(n32076), .B(n32074), .Z(n32075) );
  XOR U29407 ( .A(n32077), .B(n32078), .Z(n29207) );
  NOR U29408 ( .A(n32079), .B(n32077), .Z(n32078) );
  XOR U29409 ( .A(n32080), .B(n32081), .Z(n29210) );
  NOR U29410 ( .A(n32082), .B(n32080), .Z(n32081) );
  XOR U29411 ( .A(n32083), .B(n32084), .Z(n29213) );
  NOR U29412 ( .A(n32085), .B(n32083), .Z(n32084) );
  XOR U29413 ( .A(n32086), .B(n32087), .Z(n29216) );
  NOR U29414 ( .A(n32088), .B(n32086), .Z(n32087) );
  XOR U29415 ( .A(n32089), .B(n32090), .Z(n29219) );
  NOR U29416 ( .A(n32091), .B(n32089), .Z(n32090) );
  XOR U29417 ( .A(n32092), .B(n32093), .Z(n29222) );
  NOR U29418 ( .A(n32094), .B(n32092), .Z(n32093) );
  XOR U29419 ( .A(n32095), .B(n32096), .Z(n29225) );
  NOR U29420 ( .A(n32097), .B(n32095), .Z(n32096) );
  XOR U29421 ( .A(n32098), .B(n32099), .Z(n29228) );
  NOR U29422 ( .A(n32100), .B(n32098), .Z(n32099) );
  XOR U29423 ( .A(n32101), .B(n32102), .Z(n29231) );
  NOR U29424 ( .A(n32103), .B(n32101), .Z(n32102) );
  XOR U29425 ( .A(n32104), .B(n32105), .Z(n29234) );
  NOR U29426 ( .A(n32106), .B(n32104), .Z(n32105) );
  XOR U29427 ( .A(n32107), .B(n32108), .Z(n29237) );
  NOR U29428 ( .A(n32109), .B(n32107), .Z(n32108) );
  XOR U29429 ( .A(n32110), .B(n32111), .Z(n29240) );
  NOR U29430 ( .A(n32112), .B(n32110), .Z(n32111) );
  XOR U29431 ( .A(n32113), .B(n32114), .Z(n29243) );
  NOR U29432 ( .A(n32115), .B(n32113), .Z(n32114) );
  XOR U29433 ( .A(n32116), .B(n32117), .Z(n29246) );
  NOR U29434 ( .A(n32118), .B(n32116), .Z(n32117) );
  XOR U29435 ( .A(n32119), .B(n32120), .Z(n29249) );
  NOR U29436 ( .A(n32121), .B(n32119), .Z(n32120) );
  XOR U29437 ( .A(n32122), .B(n32123), .Z(n29252) );
  NOR U29438 ( .A(n32124), .B(n32122), .Z(n32123) );
  XOR U29439 ( .A(n32125), .B(n32126), .Z(n29255) );
  NOR U29440 ( .A(n32127), .B(n32125), .Z(n32126) );
  XOR U29441 ( .A(n32128), .B(n32129), .Z(n29258) );
  NOR U29442 ( .A(n32130), .B(n32128), .Z(n32129) );
  XOR U29443 ( .A(n32131), .B(n32132), .Z(n29261) );
  NOR U29444 ( .A(n32133), .B(n32131), .Z(n32132) );
  XOR U29445 ( .A(n32134), .B(n32135), .Z(n29264) );
  NOR U29446 ( .A(n32136), .B(n32134), .Z(n32135) );
  XOR U29447 ( .A(n32137), .B(n32138), .Z(n29267) );
  NOR U29448 ( .A(n32139), .B(n32137), .Z(n32138) );
  XOR U29449 ( .A(n32140), .B(n32141), .Z(n29270) );
  NOR U29450 ( .A(n32142), .B(n32140), .Z(n32141) );
  XOR U29451 ( .A(n32143), .B(n32144), .Z(n29273) );
  NOR U29452 ( .A(n32145), .B(n32143), .Z(n32144) );
  XOR U29453 ( .A(n32146), .B(n32147), .Z(n29276) );
  NOR U29454 ( .A(n32148), .B(n32146), .Z(n32147) );
  XOR U29455 ( .A(n32149), .B(n32150), .Z(n29279) );
  NOR U29456 ( .A(n32151), .B(n32149), .Z(n32150) );
  XOR U29457 ( .A(n32152), .B(n32153), .Z(n29282) );
  NOR U29458 ( .A(n32154), .B(n32152), .Z(n32153) );
  XOR U29459 ( .A(n32155), .B(n32156), .Z(n29285) );
  NOR U29460 ( .A(n32157), .B(n32155), .Z(n32156) );
  XOR U29461 ( .A(n32158), .B(n32159), .Z(n29288) );
  NOR U29462 ( .A(n32160), .B(n32158), .Z(n32159) );
  XOR U29463 ( .A(n32161), .B(n32162), .Z(n29291) );
  NOR U29464 ( .A(n32163), .B(n32161), .Z(n32162) );
  XOR U29465 ( .A(n32164), .B(n32165), .Z(n29294) );
  NOR U29466 ( .A(n32166), .B(n32164), .Z(n32165) );
  XOR U29467 ( .A(n32167), .B(n32168), .Z(n29297) );
  NOR U29468 ( .A(n32169), .B(n32167), .Z(n32168) );
  XOR U29469 ( .A(n32170), .B(n32171), .Z(n29300) );
  NOR U29470 ( .A(n32172), .B(n32170), .Z(n32171) );
  XOR U29471 ( .A(n32173), .B(n32174), .Z(n29303) );
  NOR U29472 ( .A(n32175), .B(n32173), .Z(n32174) );
  XOR U29473 ( .A(n32176), .B(n32177), .Z(n29306) );
  NOR U29474 ( .A(n32178), .B(n32176), .Z(n32177) );
  XOR U29475 ( .A(n32179), .B(n32180), .Z(n29309) );
  NOR U29476 ( .A(n32181), .B(n32179), .Z(n32180) );
  XOR U29477 ( .A(n32182), .B(n32183), .Z(n29312) );
  NOR U29478 ( .A(n32184), .B(n32182), .Z(n32183) );
  XOR U29479 ( .A(n32185), .B(n32186), .Z(n29315) );
  NOR U29480 ( .A(n32187), .B(n32185), .Z(n32186) );
  XOR U29481 ( .A(n32188), .B(n32189), .Z(n29318) );
  NOR U29482 ( .A(n32190), .B(n32188), .Z(n32189) );
  XOR U29483 ( .A(n32191), .B(n32192), .Z(n29321) );
  NOR U29484 ( .A(n32193), .B(n32191), .Z(n32192) );
  XOR U29485 ( .A(n32194), .B(n32195), .Z(n29324) );
  NOR U29486 ( .A(n32196), .B(n32194), .Z(n32195) );
  XOR U29487 ( .A(n32197), .B(n32198), .Z(n29327) );
  NOR U29488 ( .A(n32199), .B(n32197), .Z(n32198) );
  XOR U29489 ( .A(n32200), .B(n32201), .Z(n29330) );
  NOR U29490 ( .A(n32202), .B(n32200), .Z(n32201) );
  XOR U29491 ( .A(n32203), .B(n32204), .Z(n29333) );
  NOR U29492 ( .A(n32205), .B(n32203), .Z(n32204) );
  XOR U29493 ( .A(n32206), .B(n32207), .Z(n29336) );
  NOR U29494 ( .A(n32208), .B(n32206), .Z(n32207) );
  XOR U29495 ( .A(n32209), .B(n32210), .Z(n29339) );
  NOR U29496 ( .A(n32211), .B(n32209), .Z(n32210) );
  XOR U29497 ( .A(n32212), .B(n32213), .Z(n29342) );
  NOR U29498 ( .A(n32214), .B(n32212), .Z(n32213) );
  XOR U29499 ( .A(n32215), .B(n32216), .Z(n29345) );
  NOR U29500 ( .A(n32217), .B(n32215), .Z(n32216) );
  XOR U29501 ( .A(n32218), .B(n32219), .Z(n29348) );
  NOR U29502 ( .A(n32220), .B(n32218), .Z(n32219) );
  XOR U29503 ( .A(n32221), .B(n32222), .Z(n29351) );
  NOR U29504 ( .A(n32223), .B(n32221), .Z(n32222) );
  XOR U29505 ( .A(n32224), .B(n32225), .Z(n29354) );
  NOR U29506 ( .A(n32226), .B(n32224), .Z(n32225) );
  XOR U29507 ( .A(n32227), .B(n32228), .Z(n29357) );
  NOR U29508 ( .A(n32229), .B(n32227), .Z(n32228) );
  XOR U29509 ( .A(n32230), .B(n32231), .Z(n29360) );
  NOR U29510 ( .A(n32232), .B(n32230), .Z(n32231) );
  XOR U29511 ( .A(n32233), .B(n32234), .Z(n29363) );
  NOR U29512 ( .A(n32235), .B(n32233), .Z(n32234) );
  XOR U29513 ( .A(n32236), .B(n32237), .Z(n29366) );
  NOR U29514 ( .A(n32238), .B(n32236), .Z(n32237) );
  XOR U29515 ( .A(n32239), .B(n32240), .Z(n29369) );
  NOR U29516 ( .A(n32241), .B(n32239), .Z(n32240) );
  XOR U29517 ( .A(n32242), .B(n32243), .Z(n29372) );
  NOR U29518 ( .A(n32244), .B(n32242), .Z(n32243) );
  XOR U29519 ( .A(n32245), .B(n32246), .Z(n29375) );
  NOR U29520 ( .A(n32247), .B(n32245), .Z(n32246) );
  XOR U29521 ( .A(n32248), .B(n32249), .Z(n29378) );
  NOR U29522 ( .A(n32250), .B(n32248), .Z(n32249) );
  XOR U29523 ( .A(n32251), .B(n32252), .Z(n29381) );
  NOR U29524 ( .A(n32253), .B(n32251), .Z(n32252) );
  XOR U29525 ( .A(n32254), .B(n32255), .Z(n29384) );
  NOR U29526 ( .A(n32256), .B(n32254), .Z(n32255) );
  XOR U29527 ( .A(n32257), .B(n32258), .Z(n29387) );
  NOR U29528 ( .A(n32259), .B(n32257), .Z(n32258) );
  XOR U29529 ( .A(n32260), .B(n32261), .Z(n29390) );
  NOR U29530 ( .A(n32262), .B(n32260), .Z(n32261) );
  XOR U29531 ( .A(n32263), .B(n32264), .Z(n29393) );
  NOR U29532 ( .A(n32265), .B(n32263), .Z(n32264) );
  XOR U29533 ( .A(n32266), .B(n32267), .Z(n29396) );
  NOR U29534 ( .A(n32268), .B(n32266), .Z(n32267) );
  XOR U29535 ( .A(n32269), .B(n32270), .Z(n29399) );
  NOR U29536 ( .A(n32271), .B(n32269), .Z(n32270) );
  XOR U29537 ( .A(n32272), .B(n32273), .Z(n29402) );
  NOR U29538 ( .A(n32274), .B(n32272), .Z(n32273) );
  XOR U29539 ( .A(n32275), .B(n32276), .Z(n29405) );
  NOR U29540 ( .A(n32277), .B(n32275), .Z(n32276) );
  XOR U29541 ( .A(n32278), .B(n32279), .Z(n29408) );
  NOR U29542 ( .A(n32280), .B(n32278), .Z(n32279) );
  XOR U29543 ( .A(n32281), .B(n32282), .Z(n29411) );
  NOR U29544 ( .A(n32283), .B(n32281), .Z(n32282) );
  XOR U29545 ( .A(n32284), .B(n32285), .Z(n29414) );
  NOR U29546 ( .A(n32286), .B(n32284), .Z(n32285) );
  XOR U29547 ( .A(n32287), .B(n32288), .Z(n29417) );
  NOR U29548 ( .A(n32289), .B(n32287), .Z(n32288) );
  XOR U29549 ( .A(n32290), .B(n32291), .Z(n29420) );
  NOR U29550 ( .A(n32292), .B(n32290), .Z(n32291) );
  XOR U29551 ( .A(n32293), .B(n32294), .Z(n29423) );
  NOR U29552 ( .A(n32295), .B(n32293), .Z(n32294) );
  XOR U29553 ( .A(n32296), .B(n32297), .Z(n29426) );
  NOR U29554 ( .A(n32298), .B(n32296), .Z(n32297) );
  XOR U29555 ( .A(n32299), .B(n32300), .Z(n29429) );
  NOR U29556 ( .A(n32301), .B(n32299), .Z(n32300) );
  XOR U29557 ( .A(n32302), .B(n32303), .Z(n29432) );
  NOR U29558 ( .A(n32304), .B(n32302), .Z(n32303) );
  XOR U29559 ( .A(n32305), .B(n32306), .Z(n29435) );
  NOR U29560 ( .A(n32307), .B(n32305), .Z(n32306) );
  XOR U29561 ( .A(n32308), .B(n32309), .Z(n29438) );
  NOR U29562 ( .A(n32310), .B(n32308), .Z(n32309) );
  XOR U29563 ( .A(n32311), .B(n32312), .Z(n29441) );
  NOR U29564 ( .A(n32313), .B(n32311), .Z(n32312) );
  XOR U29565 ( .A(n32314), .B(n32315), .Z(n29444) );
  NOR U29566 ( .A(n32316), .B(n32314), .Z(n32315) );
  XOR U29567 ( .A(n32317), .B(n32318), .Z(n29447) );
  NOR U29568 ( .A(n32319), .B(n32317), .Z(n32318) );
  XOR U29569 ( .A(n32320), .B(n32321), .Z(n29450) );
  NOR U29570 ( .A(n32322), .B(n32320), .Z(n32321) );
  XOR U29571 ( .A(n32323), .B(n32324), .Z(n29453) );
  NOR U29572 ( .A(n32325), .B(n32323), .Z(n32324) );
  XOR U29573 ( .A(n32326), .B(n32327), .Z(n29456) );
  NOR U29574 ( .A(n32328), .B(n32326), .Z(n32327) );
  XOR U29575 ( .A(n32329), .B(n32330), .Z(n29459) );
  NOR U29576 ( .A(n32331), .B(n32329), .Z(n32330) );
  XOR U29577 ( .A(n32332), .B(n32333), .Z(n29462) );
  NOR U29578 ( .A(n32334), .B(n32332), .Z(n32333) );
  XOR U29579 ( .A(n32335), .B(n32336), .Z(n29465) );
  NOR U29580 ( .A(n32337), .B(n32335), .Z(n32336) );
  XOR U29581 ( .A(n32338), .B(n32339), .Z(n29468) );
  NOR U29582 ( .A(n32340), .B(n32338), .Z(n32339) );
  XOR U29583 ( .A(n32341), .B(n32342), .Z(n29471) );
  NOR U29584 ( .A(n32343), .B(n32341), .Z(n32342) );
  XOR U29585 ( .A(n32344), .B(n32345), .Z(n29474) );
  NOR U29586 ( .A(n32346), .B(n32344), .Z(n32345) );
  XOR U29587 ( .A(n32347), .B(n32348), .Z(n29477) );
  NOR U29588 ( .A(n32349), .B(n32347), .Z(n32348) );
  XOR U29589 ( .A(n32350), .B(n32351), .Z(n29480) );
  NOR U29590 ( .A(n32352), .B(n32350), .Z(n32351) );
  XOR U29591 ( .A(n32353), .B(n32354), .Z(n29483) );
  NOR U29592 ( .A(n32355), .B(n32353), .Z(n32354) );
  XOR U29593 ( .A(n32356), .B(n32357), .Z(n29486) );
  NOR U29594 ( .A(n32358), .B(n32356), .Z(n32357) );
  XOR U29595 ( .A(n32359), .B(n32360), .Z(n29489) );
  NOR U29596 ( .A(n32361), .B(n32359), .Z(n32360) );
  XOR U29597 ( .A(n32362), .B(n32363), .Z(n29492) );
  NOR U29598 ( .A(n32364), .B(n32362), .Z(n32363) );
  XOR U29599 ( .A(n32365), .B(n32366), .Z(n29495) );
  NOR U29600 ( .A(n32367), .B(n32365), .Z(n32366) );
  XOR U29601 ( .A(n32368), .B(n32369), .Z(n29498) );
  NOR U29602 ( .A(n32370), .B(n32368), .Z(n32369) );
  XOR U29603 ( .A(n32371), .B(n32372), .Z(n29501) );
  NOR U29604 ( .A(n32373), .B(n32371), .Z(n32372) );
  XOR U29605 ( .A(n32374), .B(n32375), .Z(n29504) );
  NOR U29606 ( .A(n32376), .B(n32374), .Z(n32375) );
  XOR U29607 ( .A(n32377), .B(n32378), .Z(n29507) );
  NOR U29608 ( .A(n32379), .B(n32377), .Z(n32378) );
  XOR U29609 ( .A(n32380), .B(n32381), .Z(n29510) );
  NOR U29610 ( .A(n32382), .B(n32380), .Z(n32381) );
  XOR U29611 ( .A(n32383), .B(n32384), .Z(n29513) );
  NOR U29612 ( .A(n32385), .B(n32383), .Z(n32384) );
  XOR U29613 ( .A(n32386), .B(n32387), .Z(n29516) );
  NOR U29614 ( .A(n32388), .B(n32386), .Z(n32387) );
  XOR U29615 ( .A(n32389), .B(n32390), .Z(n29519) );
  NOR U29616 ( .A(n32391), .B(n32389), .Z(n32390) );
  XOR U29617 ( .A(n32392), .B(n32393), .Z(n29522) );
  NOR U29618 ( .A(n32394), .B(n32392), .Z(n32393) );
  XOR U29619 ( .A(n32395), .B(n32396), .Z(n29525) );
  NOR U29620 ( .A(n32397), .B(n32395), .Z(n32396) );
  XOR U29621 ( .A(n32398), .B(n32399), .Z(n29528) );
  NOR U29622 ( .A(n32400), .B(n32398), .Z(n32399) );
  XOR U29623 ( .A(n32401), .B(n32402), .Z(n29531) );
  NOR U29624 ( .A(n32403), .B(n32401), .Z(n32402) );
  XOR U29625 ( .A(n32404), .B(n32405), .Z(n29534) );
  NOR U29626 ( .A(n32406), .B(n32404), .Z(n32405) );
  XOR U29627 ( .A(n32407), .B(n32408), .Z(n29537) );
  NOR U29628 ( .A(n32409), .B(n32407), .Z(n32408) );
  XOR U29629 ( .A(n32410), .B(n32411), .Z(n29540) );
  NOR U29630 ( .A(n32412), .B(n32410), .Z(n32411) );
  XOR U29631 ( .A(n32413), .B(n32414), .Z(n29543) );
  NOR U29632 ( .A(n32415), .B(n32413), .Z(n32414) );
  XOR U29633 ( .A(n32416), .B(n32417), .Z(n29546) );
  NOR U29634 ( .A(n32418), .B(n32416), .Z(n32417) );
  XOR U29635 ( .A(n32419), .B(n32420), .Z(n29549) );
  NOR U29636 ( .A(n32421), .B(n32419), .Z(n32420) );
  XOR U29637 ( .A(n32422), .B(n32423), .Z(n29552) );
  NOR U29638 ( .A(n32424), .B(n32422), .Z(n32423) );
  XOR U29639 ( .A(n32425), .B(n32426), .Z(n29555) );
  NOR U29640 ( .A(n32427), .B(n32425), .Z(n32426) );
  XOR U29641 ( .A(n32428), .B(n32429), .Z(n29558) );
  NOR U29642 ( .A(n32430), .B(n32428), .Z(n32429) );
  XOR U29643 ( .A(n32431), .B(n32432), .Z(n29561) );
  NOR U29644 ( .A(n32433), .B(n32431), .Z(n32432) );
  XOR U29645 ( .A(n32434), .B(n32435), .Z(n29564) );
  NOR U29646 ( .A(n32436), .B(n32434), .Z(n32435) );
  XOR U29647 ( .A(n32437), .B(n32438), .Z(n29567) );
  NOR U29648 ( .A(n32439), .B(n32437), .Z(n32438) );
  XOR U29649 ( .A(n32440), .B(n32441), .Z(n29570) );
  NOR U29650 ( .A(n32442), .B(n32440), .Z(n32441) );
  XOR U29651 ( .A(n32443), .B(n32444), .Z(n29573) );
  NOR U29652 ( .A(n32445), .B(n32443), .Z(n32444) );
  XOR U29653 ( .A(n32446), .B(n32447), .Z(n29576) );
  NOR U29654 ( .A(n32448), .B(n32446), .Z(n32447) );
  XOR U29655 ( .A(n32449), .B(n32450), .Z(n29579) );
  NOR U29656 ( .A(n32451), .B(n32449), .Z(n32450) );
  XOR U29657 ( .A(n32452), .B(n32453), .Z(n29582) );
  NOR U29658 ( .A(n32454), .B(n32452), .Z(n32453) );
  XOR U29659 ( .A(n32455), .B(n32456), .Z(n29585) );
  NOR U29660 ( .A(n32457), .B(n32455), .Z(n32456) );
  XOR U29661 ( .A(n32458), .B(n32459), .Z(n29588) );
  NOR U29662 ( .A(n32460), .B(n32458), .Z(n32459) );
  XOR U29663 ( .A(n32461), .B(n32462), .Z(n29591) );
  NOR U29664 ( .A(n32463), .B(n32461), .Z(n32462) );
  XOR U29665 ( .A(n32464), .B(n32465), .Z(n29594) );
  NOR U29666 ( .A(n32466), .B(n32464), .Z(n32465) );
  XOR U29667 ( .A(n32467), .B(n32468), .Z(n29597) );
  NOR U29668 ( .A(n32469), .B(n32467), .Z(n32468) );
  XOR U29669 ( .A(n32470), .B(n32471), .Z(n29600) );
  NOR U29670 ( .A(n32472), .B(n32470), .Z(n32471) );
  XOR U29671 ( .A(n32473), .B(n32474), .Z(n29603) );
  NOR U29672 ( .A(n32475), .B(n32473), .Z(n32474) );
  XOR U29673 ( .A(n32476), .B(n32477), .Z(n29606) );
  NOR U29674 ( .A(n32478), .B(n32476), .Z(n32477) );
  XOR U29675 ( .A(n32479), .B(n32480), .Z(n29609) );
  NOR U29676 ( .A(n32481), .B(n32479), .Z(n32480) );
  XOR U29677 ( .A(n32482), .B(n32483), .Z(n29612) );
  NOR U29678 ( .A(n32484), .B(n32482), .Z(n32483) );
  XOR U29679 ( .A(n32485), .B(n32486), .Z(n29615) );
  NOR U29680 ( .A(n32487), .B(n32485), .Z(n32486) );
  XOR U29681 ( .A(n32488), .B(n32489), .Z(n29618) );
  NOR U29682 ( .A(n32490), .B(n32488), .Z(n32489) );
  XOR U29683 ( .A(n32491), .B(n32492), .Z(n29621) );
  NOR U29684 ( .A(n32493), .B(n32491), .Z(n32492) );
  XOR U29685 ( .A(n32494), .B(n32495), .Z(n29624) );
  NOR U29686 ( .A(n32496), .B(n32494), .Z(n32495) );
  XOR U29687 ( .A(n32497), .B(n32498), .Z(n29627) );
  NOR U29688 ( .A(n32499), .B(n32497), .Z(n32498) );
  XOR U29689 ( .A(n32500), .B(n32501), .Z(n29630) );
  NOR U29690 ( .A(n32502), .B(n32500), .Z(n32501) );
  XOR U29691 ( .A(n32503), .B(n32504), .Z(n29633) );
  NOR U29692 ( .A(n32505), .B(n32503), .Z(n32504) );
  XOR U29693 ( .A(n32506), .B(n32507), .Z(n29636) );
  NOR U29694 ( .A(n32508), .B(n32506), .Z(n32507) );
  XOR U29695 ( .A(n32509), .B(n32510), .Z(n29639) );
  NOR U29696 ( .A(n32511), .B(n32509), .Z(n32510) );
  XOR U29697 ( .A(n32512), .B(n32513), .Z(n29642) );
  NOR U29698 ( .A(n32514), .B(n32512), .Z(n32513) );
  XOR U29699 ( .A(n32515), .B(n32516), .Z(n29645) );
  NOR U29700 ( .A(n32517), .B(n32515), .Z(n32516) );
  XOR U29701 ( .A(n32518), .B(n32519), .Z(n29648) );
  NOR U29702 ( .A(n32520), .B(n32518), .Z(n32519) );
  XOR U29703 ( .A(n32521), .B(n32522), .Z(n29651) );
  NOR U29704 ( .A(n32523), .B(n32521), .Z(n32522) );
  XOR U29705 ( .A(n32524), .B(n32525), .Z(n29654) );
  NOR U29706 ( .A(n32526), .B(n32524), .Z(n32525) );
  XOR U29707 ( .A(n32527), .B(n32528), .Z(n29657) );
  NOR U29708 ( .A(n32529), .B(n32527), .Z(n32528) );
  XOR U29709 ( .A(n32530), .B(n32531), .Z(n29660) );
  NOR U29710 ( .A(n32532), .B(n32530), .Z(n32531) );
  XOR U29711 ( .A(n32533), .B(n32534), .Z(n29663) );
  NOR U29712 ( .A(n32535), .B(n32533), .Z(n32534) );
  XOR U29713 ( .A(n32536), .B(n32537), .Z(n29666) );
  NOR U29714 ( .A(n32538), .B(n32536), .Z(n32537) );
  XOR U29715 ( .A(n32539), .B(n32540), .Z(n29669) );
  NOR U29716 ( .A(n32541), .B(n32539), .Z(n32540) );
  XOR U29717 ( .A(n32542), .B(n32543), .Z(n29672) );
  NOR U29718 ( .A(n32544), .B(n32542), .Z(n32543) );
  XOR U29719 ( .A(n32545), .B(n32546), .Z(n29675) );
  NOR U29720 ( .A(n32547), .B(n32545), .Z(n32546) );
  XOR U29721 ( .A(n32548), .B(n32549), .Z(n29678) );
  NOR U29722 ( .A(n32550), .B(n32548), .Z(n32549) );
  XOR U29723 ( .A(n32551), .B(n32552), .Z(n29681) );
  NOR U29724 ( .A(n32553), .B(n32551), .Z(n32552) );
  XOR U29725 ( .A(n32554), .B(n32555), .Z(n29684) );
  NOR U29726 ( .A(n32556), .B(n32554), .Z(n32555) );
  XOR U29727 ( .A(n32557), .B(n32558), .Z(n29687) );
  NOR U29728 ( .A(n32559), .B(n32557), .Z(n32558) );
  XOR U29729 ( .A(n32560), .B(n32561), .Z(n29690) );
  NOR U29730 ( .A(n32562), .B(n32560), .Z(n32561) );
  XOR U29731 ( .A(n32563), .B(n32564), .Z(n29693) );
  NOR U29732 ( .A(n32565), .B(n32563), .Z(n32564) );
  XOR U29733 ( .A(n32566), .B(n32567), .Z(n29696) );
  NOR U29734 ( .A(n32568), .B(n32566), .Z(n32567) );
  XOR U29735 ( .A(n32569), .B(n32570), .Z(n29699) );
  NOR U29736 ( .A(n32571), .B(n32569), .Z(n32570) );
  XOR U29737 ( .A(n32572), .B(n32573), .Z(n29702) );
  NOR U29738 ( .A(n32574), .B(n32572), .Z(n32573) );
  XOR U29739 ( .A(n32575), .B(n32576), .Z(n29705) );
  NOR U29740 ( .A(n32577), .B(n32575), .Z(n32576) );
  XOR U29741 ( .A(n32578), .B(n32579), .Z(n29708) );
  NOR U29742 ( .A(n32580), .B(n32578), .Z(n32579) );
  XOR U29743 ( .A(n32581), .B(n32582), .Z(n29711) );
  NOR U29744 ( .A(n32583), .B(n32581), .Z(n32582) );
  XOR U29745 ( .A(n32584), .B(n32585), .Z(n29714) );
  NOR U29746 ( .A(n32586), .B(n32584), .Z(n32585) );
  XOR U29747 ( .A(n32587), .B(n32588), .Z(n29717) );
  NOR U29748 ( .A(n32589), .B(n32587), .Z(n32588) );
  XOR U29749 ( .A(n32590), .B(n32591), .Z(n29720) );
  NOR U29750 ( .A(n32592), .B(n32590), .Z(n32591) );
  XOR U29751 ( .A(n32593), .B(n32594), .Z(n29723) );
  NOR U29752 ( .A(n32595), .B(n32593), .Z(n32594) );
  XOR U29753 ( .A(n32596), .B(n32597), .Z(n29726) );
  NOR U29754 ( .A(n32598), .B(n32596), .Z(n32597) );
  XOR U29755 ( .A(n32599), .B(n32600), .Z(n29729) );
  NOR U29756 ( .A(n32601), .B(n32599), .Z(n32600) );
  XOR U29757 ( .A(n32602), .B(n32603), .Z(n29732) );
  NOR U29758 ( .A(n32604), .B(n32602), .Z(n32603) );
  XOR U29759 ( .A(n32605), .B(n32606), .Z(n29735) );
  NOR U29760 ( .A(n32607), .B(n32605), .Z(n32606) );
  XOR U29761 ( .A(n32608), .B(n32609), .Z(n29738) );
  NOR U29762 ( .A(n32610), .B(n32608), .Z(n32609) );
  XOR U29763 ( .A(n32611), .B(n32612), .Z(n29741) );
  NOR U29764 ( .A(n32613), .B(n32611), .Z(n32612) );
  XOR U29765 ( .A(n32614), .B(n32615), .Z(n29744) );
  NOR U29766 ( .A(n32616), .B(n32614), .Z(n32615) );
  XOR U29767 ( .A(n32617), .B(n32618), .Z(n29747) );
  NOR U29768 ( .A(n32619), .B(n32617), .Z(n32618) );
  XOR U29769 ( .A(n32620), .B(n32621), .Z(n29750) );
  NOR U29770 ( .A(n32622), .B(n32620), .Z(n32621) );
  XOR U29771 ( .A(n32623), .B(n32624), .Z(n29753) );
  NOR U29772 ( .A(n32625), .B(n32623), .Z(n32624) );
  XOR U29773 ( .A(n32626), .B(n32627), .Z(n29756) );
  NOR U29774 ( .A(n32628), .B(n32626), .Z(n32627) );
  XOR U29775 ( .A(n32629), .B(n32630), .Z(n29759) );
  NOR U29776 ( .A(n32631), .B(n32629), .Z(n32630) );
  XOR U29777 ( .A(n32632), .B(n32633), .Z(n29762) );
  NOR U29778 ( .A(n32634), .B(n32632), .Z(n32633) );
  XOR U29779 ( .A(n32635), .B(n32636), .Z(n29765) );
  NOR U29780 ( .A(n32637), .B(n32635), .Z(n32636) );
  XOR U29781 ( .A(n32638), .B(n32639), .Z(n29768) );
  NOR U29782 ( .A(n32640), .B(n32638), .Z(n32639) );
  XOR U29783 ( .A(n32641), .B(n32642), .Z(n29771) );
  NOR U29784 ( .A(n32643), .B(n32641), .Z(n32642) );
  XOR U29785 ( .A(n32644), .B(n32645), .Z(n29774) );
  NOR U29786 ( .A(n32646), .B(n32644), .Z(n32645) );
  XOR U29787 ( .A(n32647), .B(n32648), .Z(n29777) );
  NOR U29788 ( .A(n32649), .B(n32647), .Z(n32648) );
  XOR U29789 ( .A(n32650), .B(n32651), .Z(n29780) );
  NOR U29790 ( .A(n32652), .B(n32650), .Z(n32651) );
  XOR U29791 ( .A(n32653), .B(n32654), .Z(n29783) );
  NOR U29792 ( .A(n32655), .B(n32653), .Z(n32654) );
  XOR U29793 ( .A(n32656), .B(n32657), .Z(n29786) );
  NOR U29794 ( .A(n32658), .B(n32656), .Z(n32657) );
  XOR U29795 ( .A(n32659), .B(n32660), .Z(n29789) );
  NOR U29796 ( .A(n32661), .B(n32659), .Z(n32660) );
  XOR U29797 ( .A(n32662), .B(n32663), .Z(n29792) );
  NOR U29798 ( .A(n32664), .B(n32662), .Z(n32663) );
  XOR U29799 ( .A(n32665), .B(n32666), .Z(n29795) );
  NOR U29800 ( .A(n32667), .B(n32665), .Z(n32666) );
  XOR U29801 ( .A(n32668), .B(n32669), .Z(n29798) );
  NOR U29802 ( .A(n32670), .B(n32668), .Z(n32669) );
  XOR U29803 ( .A(n32671), .B(n32672), .Z(n29801) );
  NOR U29804 ( .A(n32673), .B(n32671), .Z(n32672) );
  XOR U29805 ( .A(n32674), .B(n32675), .Z(n29804) );
  NOR U29806 ( .A(n32676), .B(n32674), .Z(n32675) );
  XOR U29807 ( .A(n32677), .B(n32678), .Z(n29807) );
  NOR U29808 ( .A(n32679), .B(n32677), .Z(n32678) );
  XOR U29809 ( .A(n32680), .B(n32681), .Z(n29810) );
  NOR U29810 ( .A(n32682), .B(n32680), .Z(n32681) );
  XOR U29811 ( .A(n32683), .B(n32684), .Z(n29813) );
  AND U29812 ( .A(n32685), .B(n32683), .Z(n32684) );
  XOR U29813 ( .A(n32686), .B(n32687), .Z(n29816) );
  AND U29814 ( .A(n94), .B(n32686), .Z(n32687) );
  XOR U29815 ( .A(n76), .B(n31270), .Z(n31272) );
  XOR U29816 ( .A(n31267), .B(n31266), .Z(n76) );
  XNOR U29817 ( .A(n31264), .B(n31263), .Z(n31266) );
  XNOR U29818 ( .A(n31261), .B(n31260), .Z(n31263) );
  XNOR U29819 ( .A(n31258), .B(n31257), .Z(n31260) );
  XNOR U29820 ( .A(n31255), .B(n31254), .Z(n31257) );
  XNOR U29821 ( .A(n31252), .B(n31251), .Z(n31254) );
  XNOR U29822 ( .A(n31249), .B(n31248), .Z(n31251) );
  XNOR U29823 ( .A(n31246), .B(n31245), .Z(n31248) );
  XNOR U29824 ( .A(n31243), .B(n31242), .Z(n31245) );
  XNOR U29825 ( .A(n31240), .B(n31239), .Z(n31242) );
  XNOR U29826 ( .A(n31237), .B(n31236), .Z(n31239) );
  XNOR U29827 ( .A(n31234), .B(n31233), .Z(n31236) );
  XNOR U29828 ( .A(n31231), .B(n31230), .Z(n31233) );
  XNOR U29829 ( .A(n31228), .B(n31227), .Z(n31230) );
  XNOR U29830 ( .A(n31225), .B(n31224), .Z(n31227) );
  XNOR U29831 ( .A(n31222), .B(n31221), .Z(n31224) );
  XNOR U29832 ( .A(n31219), .B(n31218), .Z(n31221) );
  XNOR U29833 ( .A(n31216), .B(n31215), .Z(n31218) );
  XNOR U29834 ( .A(n31213), .B(n31212), .Z(n31215) );
  XNOR U29835 ( .A(n31210), .B(n31209), .Z(n31212) );
  XNOR U29836 ( .A(n31207), .B(n31206), .Z(n31209) );
  XNOR U29837 ( .A(n31204), .B(n31203), .Z(n31206) );
  XNOR U29838 ( .A(n31201), .B(n31200), .Z(n31203) );
  XNOR U29839 ( .A(n31198), .B(n31197), .Z(n31200) );
  XNOR U29840 ( .A(n31195), .B(n31194), .Z(n31197) );
  XNOR U29841 ( .A(n31192), .B(n31191), .Z(n31194) );
  XNOR U29842 ( .A(n31189), .B(n31188), .Z(n31191) );
  XNOR U29843 ( .A(n31186), .B(n31185), .Z(n31188) );
  XNOR U29844 ( .A(n31183), .B(n31182), .Z(n31185) );
  XNOR U29845 ( .A(n31180), .B(n31179), .Z(n31182) );
  XNOR U29846 ( .A(n31177), .B(n31176), .Z(n31179) );
  XNOR U29847 ( .A(n31174), .B(n31173), .Z(n31176) );
  XNOR U29848 ( .A(n31171), .B(n31170), .Z(n31173) );
  XNOR U29849 ( .A(n31168), .B(n31167), .Z(n31170) );
  XNOR U29850 ( .A(n31165), .B(n31164), .Z(n31167) );
  XNOR U29851 ( .A(n31162), .B(n31161), .Z(n31164) );
  XNOR U29852 ( .A(n31159), .B(n31158), .Z(n31161) );
  XNOR U29853 ( .A(n31156), .B(n31155), .Z(n31158) );
  XNOR U29854 ( .A(n31153), .B(n31152), .Z(n31155) );
  XNOR U29855 ( .A(n31150), .B(n31149), .Z(n31152) );
  XNOR U29856 ( .A(n31147), .B(n31146), .Z(n31149) );
  XNOR U29857 ( .A(n31144), .B(n31143), .Z(n31146) );
  XNOR U29858 ( .A(n31141), .B(n31140), .Z(n31143) );
  XNOR U29859 ( .A(n31138), .B(n31137), .Z(n31140) );
  XNOR U29860 ( .A(n31135), .B(n31134), .Z(n31137) );
  XNOR U29861 ( .A(n31132), .B(n31131), .Z(n31134) );
  XNOR U29862 ( .A(n31129), .B(n31128), .Z(n31131) );
  XNOR U29863 ( .A(n31126), .B(n31125), .Z(n31128) );
  XNOR U29864 ( .A(n31123), .B(n31122), .Z(n31125) );
  XNOR U29865 ( .A(n31120), .B(n31119), .Z(n31122) );
  XNOR U29866 ( .A(n31117), .B(n31116), .Z(n31119) );
  XNOR U29867 ( .A(n31114), .B(n31113), .Z(n31116) );
  XNOR U29868 ( .A(n31111), .B(n31110), .Z(n31113) );
  XNOR U29869 ( .A(n31108), .B(n31107), .Z(n31110) );
  XNOR U29870 ( .A(n31105), .B(n31104), .Z(n31107) );
  XNOR U29871 ( .A(n31102), .B(n31101), .Z(n31104) );
  XNOR U29872 ( .A(n31099), .B(n31098), .Z(n31101) );
  XNOR U29873 ( .A(n31096), .B(n31095), .Z(n31098) );
  XNOR U29874 ( .A(n31093), .B(n31092), .Z(n31095) );
  XNOR U29875 ( .A(n31090), .B(n31089), .Z(n31092) );
  XNOR U29876 ( .A(n31087), .B(n31086), .Z(n31089) );
  XNOR U29877 ( .A(n31084), .B(n31083), .Z(n31086) );
  XNOR U29878 ( .A(n31081), .B(n31080), .Z(n31083) );
  XNOR U29879 ( .A(n31078), .B(n31077), .Z(n31080) );
  XNOR U29880 ( .A(n31075), .B(n31074), .Z(n31077) );
  XNOR U29881 ( .A(n31072), .B(n31071), .Z(n31074) );
  XNOR U29882 ( .A(n31069), .B(n31068), .Z(n31071) );
  XNOR U29883 ( .A(n31066), .B(n31065), .Z(n31068) );
  XNOR U29884 ( .A(n31063), .B(n31062), .Z(n31065) );
  XNOR U29885 ( .A(n31060), .B(n31059), .Z(n31062) );
  XNOR U29886 ( .A(n31057), .B(n31056), .Z(n31059) );
  XNOR U29887 ( .A(n31054), .B(n31053), .Z(n31056) );
  XNOR U29888 ( .A(n31051), .B(n31050), .Z(n31053) );
  XNOR U29889 ( .A(n31048), .B(n31047), .Z(n31050) );
  XNOR U29890 ( .A(n31045), .B(n31044), .Z(n31047) );
  XNOR U29891 ( .A(n31042), .B(n31041), .Z(n31044) );
  XNOR U29892 ( .A(n31039), .B(n31038), .Z(n31041) );
  XNOR U29893 ( .A(n31036), .B(n31035), .Z(n31038) );
  XNOR U29894 ( .A(n31033), .B(n31032), .Z(n31035) );
  XNOR U29895 ( .A(n31030), .B(n31029), .Z(n31032) );
  XNOR U29896 ( .A(n31027), .B(n31026), .Z(n31029) );
  XNOR U29897 ( .A(n31024), .B(n31023), .Z(n31026) );
  XNOR U29898 ( .A(n31021), .B(n31020), .Z(n31023) );
  XNOR U29899 ( .A(n31018), .B(n31017), .Z(n31020) );
  XNOR U29900 ( .A(n31015), .B(n31014), .Z(n31017) );
  XNOR U29901 ( .A(n31012), .B(n31011), .Z(n31014) );
  XNOR U29902 ( .A(n31009), .B(n31008), .Z(n31011) );
  XNOR U29903 ( .A(n31006), .B(n31005), .Z(n31008) );
  XNOR U29904 ( .A(n31003), .B(n31002), .Z(n31005) );
  XNOR U29905 ( .A(n31000), .B(n30999), .Z(n31002) );
  XNOR U29906 ( .A(n30997), .B(n30996), .Z(n30999) );
  XNOR U29907 ( .A(n30994), .B(n30993), .Z(n30996) );
  XNOR U29908 ( .A(n30991), .B(n30990), .Z(n30993) );
  XNOR U29909 ( .A(n30988), .B(n30987), .Z(n30990) );
  XNOR U29910 ( .A(n30985), .B(n30984), .Z(n30987) );
  XNOR U29911 ( .A(n30982), .B(n30981), .Z(n30984) );
  XNOR U29912 ( .A(n30979), .B(n30978), .Z(n30981) );
  XNOR U29913 ( .A(n30976), .B(n30975), .Z(n30978) );
  XNOR U29914 ( .A(n30973), .B(n30972), .Z(n30975) );
  XNOR U29915 ( .A(n30970), .B(n30969), .Z(n30972) );
  XNOR U29916 ( .A(n30967), .B(n30966), .Z(n30969) );
  XNOR U29917 ( .A(n30964), .B(n30963), .Z(n30966) );
  XNOR U29918 ( .A(n30961), .B(n30960), .Z(n30963) );
  XNOR U29919 ( .A(n30958), .B(n30957), .Z(n30960) );
  XNOR U29920 ( .A(n30955), .B(n30954), .Z(n30957) );
  XNOR U29921 ( .A(n30952), .B(n30951), .Z(n30954) );
  XNOR U29922 ( .A(n30949), .B(n30948), .Z(n30951) );
  XNOR U29923 ( .A(n30946), .B(n30945), .Z(n30948) );
  XNOR U29924 ( .A(n30943), .B(n30942), .Z(n30945) );
  XNOR U29925 ( .A(n30940), .B(n30939), .Z(n30942) );
  XNOR U29926 ( .A(n30937), .B(n30936), .Z(n30939) );
  XNOR U29927 ( .A(n30934), .B(n30933), .Z(n30936) );
  XNOR U29928 ( .A(n30931), .B(n30930), .Z(n30933) );
  XNOR U29929 ( .A(n30928), .B(n30927), .Z(n30930) );
  XNOR U29930 ( .A(n30925), .B(n30924), .Z(n30927) );
  XNOR U29931 ( .A(n30922), .B(n30921), .Z(n30924) );
  XNOR U29932 ( .A(n30919), .B(n30918), .Z(n30921) );
  XNOR U29933 ( .A(n30916), .B(n30915), .Z(n30918) );
  XNOR U29934 ( .A(n30913), .B(n30912), .Z(n30915) );
  XNOR U29935 ( .A(n30910), .B(n30909), .Z(n30912) );
  XNOR U29936 ( .A(n30907), .B(n30906), .Z(n30909) );
  XNOR U29937 ( .A(n30904), .B(n30903), .Z(n30906) );
  XNOR U29938 ( .A(n30901), .B(n30900), .Z(n30903) );
  XNOR U29939 ( .A(n30898), .B(n30897), .Z(n30900) );
  XNOR U29940 ( .A(n30895), .B(n30894), .Z(n30897) );
  XNOR U29941 ( .A(n30892), .B(n30891), .Z(n30894) );
  XNOR U29942 ( .A(n30889), .B(n30888), .Z(n30891) );
  XNOR U29943 ( .A(n30886), .B(n30885), .Z(n30888) );
  XNOR U29944 ( .A(n30883), .B(n30882), .Z(n30885) );
  XNOR U29945 ( .A(n30880), .B(n30879), .Z(n30882) );
  XNOR U29946 ( .A(n30877), .B(n30876), .Z(n30879) );
  XNOR U29947 ( .A(n30874), .B(n30873), .Z(n30876) );
  XNOR U29948 ( .A(n30871), .B(n30870), .Z(n30873) );
  XNOR U29949 ( .A(n30868), .B(n30867), .Z(n30870) );
  XNOR U29950 ( .A(n30865), .B(n30864), .Z(n30867) );
  XNOR U29951 ( .A(n30862), .B(n30861), .Z(n30864) );
  XNOR U29952 ( .A(n30859), .B(n30858), .Z(n30861) );
  XNOR U29953 ( .A(n30856), .B(n30855), .Z(n30858) );
  XNOR U29954 ( .A(n30853), .B(n30852), .Z(n30855) );
  XNOR U29955 ( .A(n30850), .B(n30849), .Z(n30852) );
  XNOR U29956 ( .A(n30847), .B(n30846), .Z(n30849) );
  XNOR U29957 ( .A(n30844), .B(n30843), .Z(n30846) );
  XNOR U29958 ( .A(n30841), .B(n30840), .Z(n30843) );
  XNOR U29959 ( .A(n30838), .B(n30837), .Z(n30840) );
  XNOR U29960 ( .A(n30835), .B(n30834), .Z(n30837) );
  XNOR U29961 ( .A(n30832), .B(n30831), .Z(n30834) );
  XNOR U29962 ( .A(n30829), .B(n30828), .Z(n30831) );
  XNOR U29963 ( .A(n30826), .B(n30825), .Z(n30828) );
  XNOR U29964 ( .A(n30823), .B(n30822), .Z(n30825) );
  XNOR U29965 ( .A(n30820), .B(n30819), .Z(n30822) );
  XNOR U29966 ( .A(n30817), .B(n30816), .Z(n30819) );
  XNOR U29967 ( .A(n30814), .B(n30813), .Z(n30816) );
  XNOR U29968 ( .A(n30811), .B(n30810), .Z(n30813) );
  XNOR U29969 ( .A(n30808), .B(n30807), .Z(n30810) );
  XNOR U29970 ( .A(n30805), .B(n30804), .Z(n30807) );
  XNOR U29971 ( .A(n30802), .B(n30801), .Z(n30804) );
  XNOR U29972 ( .A(n30799), .B(n30798), .Z(n30801) );
  XNOR U29973 ( .A(n30796), .B(n30795), .Z(n30798) );
  XNOR U29974 ( .A(n30793), .B(n30792), .Z(n30795) );
  XNOR U29975 ( .A(n30790), .B(n30789), .Z(n30792) );
  XNOR U29976 ( .A(n30787), .B(n30786), .Z(n30789) );
  XNOR U29977 ( .A(n30784), .B(n30783), .Z(n30786) );
  XNOR U29978 ( .A(n30781), .B(n30780), .Z(n30783) );
  XNOR U29979 ( .A(n30778), .B(n30777), .Z(n30780) );
  XNOR U29980 ( .A(n30775), .B(n30774), .Z(n30777) );
  XNOR U29981 ( .A(n30772), .B(n30771), .Z(n30774) );
  XNOR U29982 ( .A(n30769), .B(n30768), .Z(n30771) );
  XNOR U29983 ( .A(n30766), .B(n30765), .Z(n30768) );
  XNOR U29984 ( .A(n30763), .B(n30762), .Z(n30765) );
  XNOR U29985 ( .A(n30760), .B(n30759), .Z(n30762) );
  XNOR U29986 ( .A(n30757), .B(n30756), .Z(n30759) );
  XNOR U29987 ( .A(n30754), .B(n30753), .Z(n30756) );
  XNOR U29988 ( .A(n30751), .B(n30750), .Z(n30753) );
  XNOR U29989 ( .A(n30748), .B(n30747), .Z(n30750) );
  XNOR U29990 ( .A(n30745), .B(n30744), .Z(n30747) );
  XNOR U29991 ( .A(n30742), .B(n30741), .Z(n30744) );
  XNOR U29992 ( .A(n30739), .B(n30738), .Z(n30741) );
  XNOR U29993 ( .A(n30736), .B(n30735), .Z(n30738) );
  XNOR U29994 ( .A(n30733), .B(n30732), .Z(n30735) );
  XNOR U29995 ( .A(n30730), .B(n30729), .Z(n30732) );
  XNOR U29996 ( .A(n30727), .B(n30726), .Z(n30729) );
  XNOR U29997 ( .A(n30724), .B(n30723), .Z(n30726) );
  XNOR U29998 ( .A(n30721), .B(n30720), .Z(n30723) );
  XNOR U29999 ( .A(n30718), .B(n30717), .Z(n30720) );
  XNOR U30000 ( .A(n30715), .B(n30714), .Z(n30717) );
  XNOR U30001 ( .A(n30712), .B(n30711), .Z(n30714) );
  XNOR U30002 ( .A(n30709), .B(n30708), .Z(n30711) );
  XNOR U30003 ( .A(n30706), .B(n30705), .Z(n30708) );
  XNOR U30004 ( .A(n30703), .B(n30702), .Z(n30705) );
  XNOR U30005 ( .A(n30700), .B(n30699), .Z(n30702) );
  XNOR U30006 ( .A(n30697), .B(n30696), .Z(n30699) );
  XNOR U30007 ( .A(n30694), .B(n30693), .Z(n30696) );
  XNOR U30008 ( .A(n30691), .B(n30690), .Z(n30693) );
  XNOR U30009 ( .A(n30688), .B(n30687), .Z(n30690) );
  XNOR U30010 ( .A(n30685), .B(n30684), .Z(n30687) );
  XNOR U30011 ( .A(n30682), .B(n30681), .Z(n30684) );
  XNOR U30012 ( .A(n30679), .B(n30678), .Z(n30681) );
  XNOR U30013 ( .A(n30676), .B(n30675), .Z(n30678) );
  XNOR U30014 ( .A(n30673), .B(n30672), .Z(n30675) );
  XNOR U30015 ( .A(n30670), .B(n30669), .Z(n30672) );
  XNOR U30016 ( .A(n30667), .B(n30666), .Z(n30669) );
  XNOR U30017 ( .A(n30664), .B(n30663), .Z(n30666) );
  XNOR U30018 ( .A(n30661), .B(n30660), .Z(n30663) );
  XNOR U30019 ( .A(n30658), .B(n30657), .Z(n30660) );
  XNOR U30020 ( .A(n30655), .B(n30654), .Z(n30657) );
  XNOR U30021 ( .A(n30652), .B(n30651), .Z(n30654) );
  XNOR U30022 ( .A(n30649), .B(n30648), .Z(n30651) );
  XNOR U30023 ( .A(n30646), .B(n30645), .Z(n30648) );
  XNOR U30024 ( .A(n30643), .B(n30642), .Z(n30645) );
  XNOR U30025 ( .A(n30640), .B(n30639), .Z(n30642) );
  XNOR U30026 ( .A(n30637), .B(n30636), .Z(n30639) );
  XNOR U30027 ( .A(n30634), .B(n30633), .Z(n30636) );
  XNOR U30028 ( .A(n30631), .B(n30630), .Z(n30633) );
  XNOR U30029 ( .A(n30628), .B(n30627), .Z(n30630) );
  XNOR U30030 ( .A(n30625), .B(n30624), .Z(n30627) );
  XNOR U30031 ( .A(n30622), .B(n30621), .Z(n30624) );
  XNOR U30032 ( .A(n30619), .B(n30618), .Z(n30621) );
  XNOR U30033 ( .A(n30616), .B(n30615), .Z(n30618) );
  XNOR U30034 ( .A(n30613), .B(n30612), .Z(n30615) );
  XNOR U30035 ( .A(n30610), .B(n30609), .Z(n30612) );
  XNOR U30036 ( .A(n30607), .B(n30606), .Z(n30609) );
  XNOR U30037 ( .A(n30604), .B(n30603), .Z(n30606) );
  XNOR U30038 ( .A(n30601), .B(n30600), .Z(n30603) );
  XNOR U30039 ( .A(n30598), .B(n30597), .Z(n30600) );
  XNOR U30040 ( .A(n30595), .B(n30594), .Z(n30597) );
  XNOR U30041 ( .A(n30592), .B(n30591), .Z(n30594) );
  XNOR U30042 ( .A(n30589), .B(n30588), .Z(n30591) );
  XNOR U30043 ( .A(n30586), .B(n30585), .Z(n30588) );
  XNOR U30044 ( .A(n30583), .B(n30582), .Z(n30585) );
  XNOR U30045 ( .A(n30580), .B(n30579), .Z(n30582) );
  XNOR U30046 ( .A(n30577), .B(n30576), .Z(n30579) );
  XNOR U30047 ( .A(n30574), .B(n30573), .Z(n30576) );
  XNOR U30048 ( .A(n30571), .B(n30570), .Z(n30573) );
  XNOR U30049 ( .A(n30568), .B(n30567), .Z(n30570) );
  XNOR U30050 ( .A(n30565), .B(n30564), .Z(n30567) );
  XNOR U30051 ( .A(n30562), .B(n30561), .Z(n30564) );
  XNOR U30052 ( .A(n30559), .B(n30558), .Z(n30561) );
  XNOR U30053 ( .A(n30556), .B(n30555), .Z(n30558) );
  XNOR U30054 ( .A(n30553), .B(n30552), .Z(n30555) );
  XNOR U30055 ( .A(n30550), .B(n30549), .Z(n30552) );
  XNOR U30056 ( .A(n30547), .B(n30546), .Z(n30549) );
  XNOR U30057 ( .A(n30544), .B(n30543), .Z(n30546) );
  XNOR U30058 ( .A(n30541), .B(n30540), .Z(n30543) );
  XNOR U30059 ( .A(n30538), .B(n30537), .Z(n30540) );
  XNOR U30060 ( .A(n30535), .B(n30534), .Z(n30537) );
  XNOR U30061 ( .A(n30532), .B(n30531), .Z(n30534) );
  XNOR U30062 ( .A(n30529), .B(n30528), .Z(n30531) );
  XNOR U30063 ( .A(n30526), .B(n30525), .Z(n30528) );
  XNOR U30064 ( .A(n30523), .B(n30522), .Z(n30525) );
  XNOR U30065 ( .A(n30520), .B(n30519), .Z(n30522) );
  XNOR U30066 ( .A(n30517), .B(n30516), .Z(n30519) );
  XNOR U30067 ( .A(n30514), .B(n30513), .Z(n30516) );
  XNOR U30068 ( .A(n30511), .B(n30510), .Z(n30513) );
  XNOR U30069 ( .A(n30508), .B(n30507), .Z(n30510) );
  XNOR U30070 ( .A(n30505), .B(n30504), .Z(n30507) );
  XNOR U30071 ( .A(n30502), .B(n30501), .Z(n30504) );
  XNOR U30072 ( .A(n30499), .B(n30498), .Z(n30501) );
  XNOR U30073 ( .A(n30496), .B(n30495), .Z(n30498) );
  XNOR U30074 ( .A(n30493), .B(n30492), .Z(n30495) );
  XNOR U30075 ( .A(n30490), .B(n30489), .Z(n30492) );
  XNOR U30076 ( .A(n30487), .B(n30486), .Z(n30489) );
  XNOR U30077 ( .A(n30484), .B(n30483), .Z(n30486) );
  XNOR U30078 ( .A(n30481), .B(n30480), .Z(n30483) );
  XNOR U30079 ( .A(n30478), .B(n30477), .Z(n30480) );
  XNOR U30080 ( .A(n30475), .B(n30474), .Z(n30477) );
  XNOR U30081 ( .A(n30472), .B(n30471), .Z(n30474) );
  XNOR U30082 ( .A(n30469), .B(n30468), .Z(n30471) );
  XNOR U30083 ( .A(n30466), .B(n30465), .Z(n30468) );
  XNOR U30084 ( .A(n30463), .B(n30462), .Z(n30465) );
  XNOR U30085 ( .A(n30460), .B(n30459), .Z(n30462) );
  XNOR U30086 ( .A(n30457), .B(n30456), .Z(n30459) );
  XNOR U30087 ( .A(n30454), .B(n30453), .Z(n30456) );
  XNOR U30088 ( .A(n30451), .B(n30450), .Z(n30453) );
  XNOR U30089 ( .A(n30448), .B(n30447), .Z(n30450) );
  XNOR U30090 ( .A(n30445), .B(n30444), .Z(n30447) );
  XNOR U30091 ( .A(n30442), .B(n30441), .Z(n30444) );
  XNOR U30092 ( .A(n30439), .B(n30438), .Z(n30441) );
  XNOR U30093 ( .A(n30436), .B(n30435), .Z(n30438) );
  XNOR U30094 ( .A(n30433), .B(n30432), .Z(n30435) );
  XNOR U30095 ( .A(n30430), .B(n30429), .Z(n30432) );
  XNOR U30096 ( .A(n30427), .B(n30426), .Z(n30429) );
  XNOR U30097 ( .A(n30424), .B(n30423), .Z(n30426) );
  XNOR U30098 ( .A(n30421), .B(n30420), .Z(n30423) );
  XNOR U30099 ( .A(n30418), .B(n30417), .Z(n30420) );
  XNOR U30100 ( .A(n30415), .B(n30414), .Z(n30417) );
  XNOR U30101 ( .A(n30412), .B(n30411), .Z(n30414) );
  XNOR U30102 ( .A(n30409), .B(n30408), .Z(n30411) );
  XNOR U30103 ( .A(n30406), .B(n30405), .Z(n30408) );
  XNOR U30104 ( .A(n30403), .B(n30402), .Z(n30405) );
  XNOR U30105 ( .A(n30400), .B(n30399), .Z(n30402) );
  XNOR U30106 ( .A(n30397), .B(n30396), .Z(n30399) );
  XNOR U30107 ( .A(n30394), .B(n30393), .Z(n30396) );
  XNOR U30108 ( .A(n30391), .B(n30390), .Z(n30393) );
  XNOR U30109 ( .A(n30388), .B(n30387), .Z(n30390) );
  XNOR U30110 ( .A(n30385), .B(n30384), .Z(n30387) );
  XNOR U30111 ( .A(n30382), .B(n30381), .Z(n30384) );
  XNOR U30112 ( .A(n30379), .B(n30378), .Z(n30381) );
  XNOR U30113 ( .A(n30376), .B(n30375), .Z(n30378) );
  XNOR U30114 ( .A(n30373), .B(n30372), .Z(n30375) );
  XNOR U30115 ( .A(n30370), .B(n30369), .Z(n30372) );
  XNOR U30116 ( .A(n30367), .B(n30366), .Z(n30369) );
  XNOR U30117 ( .A(n30364), .B(n30363), .Z(n30366) );
  XNOR U30118 ( .A(n30361), .B(n30360), .Z(n30363) );
  XNOR U30119 ( .A(n30358), .B(n30357), .Z(n30360) );
  XNOR U30120 ( .A(n30355), .B(n30354), .Z(n30357) );
  XNOR U30121 ( .A(n30352), .B(n30351), .Z(n30354) );
  XNOR U30122 ( .A(n30349), .B(n30348), .Z(n30351) );
  XNOR U30123 ( .A(n30346), .B(n30345), .Z(n30348) );
  XNOR U30124 ( .A(n30343), .B(n30342), .Z(n30345) );
  XNOR U30125 ( .A(n30340), .B(n30339), .Z(n30342) );
  XNOR U30126 ( .A(n30337), .B(n30336), .Z(n30339) );
  XNOR U30127 ( .A(n30334), .B(n30333), .Z(n30336) );
  XNOR U30128 ( .A(n30331), .B(n30330), .Z(n30333) );
  XNOR U30129 ( .A(n30328), .B(n30327), .Z(n30330) );
  XNOR U30130 ( .A(n30325), .B(n30324), .Z(n30327) );
  XNOR U30131 ( .A(n30322), .B(n30321), .Z(n30324) );
  XNOR U30132 ( .A(n30319), .B(n30318), .Z(n30321) );
  XNOR U30133 ( .A(n30316), .B(n30315), .Z(n30318) );
  XNOR U30134 ( .A(n30313), .B(n30312), .Z(n30315) );
  XNOR U30135 ( .A(n30310), .B(n30309), .Z(n30312) );
  XNOR U30136 ( .A(n30307), .B(n30306), .Z(n30309) );
  XNOR U30137 ( .A(n30304), .B(n30303), .Z(n30306) );
  XNOR U30138 ( .A(n30301), .B(n30300), .Z(n30303) );
  XNOR U30139 ( .A(n30298), .B(n30297), .Z(n30300) );
  XNOR U30140 ( .A(n30295), .B(n30294), .Z(n30297) );
  XNOR U30141 ( .A(n30292), .B(n30291), .Z(n30294) );
  XNOR U30142 ( .A(n30289), .B(n30288), .Z(n30291) );
  XNOR U30143 ( .A(n30286), .B(n30285), .Z(n30288) );
  XNOR U30144 ( .A(n30283), .B(n30282), .Z(n30285) );
  XNOR U30145 ( .A(n30280), .B(n30279), .Z(n30282) );
  XNOR U30146 ( .A(n30277), .B(n30276), .Z(n30279) );
  XNOR U30147 ( .A(n30274), .B(n30273), .Z(n30276) );
  XNOR U30148 ( .A(n30271), .B(n30270), .Z(n30273) );
  XNOR U30149 ( .A(n30268), .B(n30267), .Z(n30270) );
  XNOR U30150 ( .A(n30265), .B(n30264), .Z(n30267) );
  XNOR U30151 ( .A(n30262), .B(n30261), .Z(n30264) );
  XNOR U30152 ( .A(n30259), .B(n30258), .Z(n30261) );
  XNOR U30153 ( .A(n30256), .B(n30255), .Z(n30258) );
  XNOR U30154 ( .A(n30253), .B(n30252), .Z(n30255) );
  XNOR U30155 ( .A(n30250), .B(n30249), .Z(n30252) );
  XNOR U30156 ( .A(n30247), .B(n30246), .Z(n30249) );
  XNOR U30157 ( .A(n30244), .B(n30243), .Z(n30246) );
  XNOR U30158 ( .A(n30241), .B(n30240), .Z(n30243) );
  XNOR U30159 ( .A(n30238), .B(n30237), .Z(n30240) );
  XNOR U30160 ( .A(n30235), .B(n30234), .Z(n30237) );
  XNOR U30161 ( .A(n30232), .B(n30231), .Z(n30234) );
  XNOR U30162 ( .A(n30229), .B(n30228), .Z(n30231) );
  XNOR U30163 ( .A(n30226), .B(n30225), .Z(n30228) );
  XNOR U30164 ( .A(n30223), .B(n30222), .Z(n30225) );
  XNOR U30165 ( .A(n30220), .B(n30219), .Z(n30222) );
  XNOR U30166 ( .A(n30217), .B(n30216), .Z(n30219) );
  XNOR U30167 ( .A(n30214), .B(n30213), .Z(n30216) );
  XNOR U30168 ( .A(n30211), .B(n30210), .Z(n30213) );
  XNOR U30169 ( .A(n30208), .B(n30207), .Z(n30210) );
  XNOR U30170 ( .A(n30205), .B(n30204), .Z(n30207) );
  XNOR U30171 ( .A(n30202), .B(n30201), .Z(n30204) );
  XNOR U30172 ( .A(n30199), .B(n30198), .Z(n30201) );
  XNOR U30173 ( .A(n30196), .B(n30195), .Z(n30198) );
  XNOR U30174 ( .A(n30193), .B(n30192), .Z(n30195) );
  XNOR U30175 ( .A(n30190), .B(n30189), .Z(n30192) );
  XNOR U30176 ( .A(n30187), .B(n30186), .Z(n30189) );
  XNOR U30177 ( .A(n30184), .B(n30183), .Z(n30186) );
  XNOR U30178 ( .A(n30181), .B(n30180), .Z(n30183) );
  XNOR U30179 ( .A(n30178), .B(n30177), .Z(n30180) );
  XNOR U30180 ( .A(n30175), .B(n30174), .Z(n30177) );
  XNOR U30181 ( .A(n30172), .B(n30171), .Z(n30174) );
  XNOR U30182 ( .A(n30169), .B(n30168), .Z(n30171) );
  XNOR U30183 ( .A(n30166), .B(n30165), .Z(n30168) );
  XNOR U30184 ( .A(n30163), .B(n30162), .Z(n30165) );
  XNOR U30185 ( .A(n30160), .B(n30159), .Z(n30162) );
  XNOR U30186 ( .A(n30157), .B(n30156), .Z(n30159) );
  XNOR U30187 ( .A(n30154), .B(n30153), .Z(n30156) );
  XNOR U30188 ( .A(n30151), .B(n30150), .Z(n30153) );
  XNOR U30189 ( .A(n30148), .B(n30147), .Z(n30150) );
  XNOR U30190 ( .A(n30145), .B(n30144), .Z(n30147) );
  XNOR U30191 ( .A(n30142), .B(n30141), .Z(n30144) );
  XNOR U30192 ( .A(n30139), .B(n30138), .Z(n30141) );
  XNOR U30193 ( .A(n30136), .B(n30135), .Z(n30138) );
  XNOR U30194 ( .A(n30133), .B(n30132), .Z(n30135) );
  XNOR U30195 ( .A(n30130), .B(n30129), .Z(n30132) );
  XNOR U30196 ( .A(n30127), .B(n30126), .Z(n30129) );
  XNOR U30197 ( .A(n30124), .B(n30123), .Z(n30126) );
  XNOR U30198 ( .A(n30121), .B(n30120), .Z(n30123) );
  XNOR U30199 ( .A(n30118), .B(n30117), .Z(n30120) );
  XOR U30200 ( .A(n30115), .B(n29842), .Z(n30117) );
  XOR U30201 ( .A(n32688), .B(n29830), .Z(n29842) );
  XNOR U30202 ( .A(n29831), .B(n29828), .Z(n29830) );
  XNOR U30203 ( .A(n29829), .B(n29825), .Z(n29828) );
  XNOR U30204 ( .A(n29824), .B(n29851), .Z(n29825) );
  XNOR U30205 ( .A(n29850), .B(n30114), .Z(n29851) );
  XNOR U30206 ( .A(n30105), .B(n30113), .Z(n30114) );
  XNOR U30207 ( .A(n30104), .B(n30110), .Z(n30113) );
  XNOR U30208 ( .A(n30109), .B(n30092), .Z(n30110) );
  XNOR U30209 ( .A(n29857), .B(n30103), .Z(n30092) );
  XNOR U30210 ( .A(n30094), .B(n30102), .Z(n30103) );
  XOR U30211 ( .A(n30093), .B(n30099), .Z(n30102) );
  XOR U30212 ( .A(n30098), .B(n30082), .Z(n30099) );
  XOR U30213 ( .A(n29860), .B(n30091), .Z(n30082) );
  XOR U30214 ( .A(n30078), .B(n30088), .Z(n30091) );
  XOR U30215 ( .A(n30081), .B(n30087), .Z(n30088) );
  XOR U30216 ( .A(n30077), .B(n29856), .Z(n30087) );
  AND U30217 ( .A(n32689), .B(n32690), .Z(n29856) );
  XOR U30218 ( .A(n30076), .B(n30072), .Z(n30077) );
  AND U30219 ( .A(n32691), .B(n32692), .Z(n30072) );
  XOR U30220 ( .A(n30073), .B(n30066), .Z(n30076) );
  AND U30221 ( .A(n32693), .B(n32694), .Z(n30066) );
  XNOR U30222 ( .A(n30067), .B(n30065), .Z(n30073) );
  AND U30223 ( .A(n32695), .B(n32696), .Z(n30065) );
  XOR U30224 ( .A(n30018), .B(n30068), .Z(n30067) );
  AND U30225 ( .A(n32697), .B(n32698), .Z(n30068) );
  XNOR U30226 ( .A(n30062), .B(n30019), .Z(n30018) );
  AND U30227 ( .A(n32699), .B(n32700), .Z(n30019) );
  XOR U30228 ( .A(n30061), .B(n30053), .Z(n30062) );
  AND U30229 ( .A(n32701), .B(n32702), .Z(n30053) );
  XNOR U30230 ( .A(n30056), .B(n30052), .Z(n30061) );
  AND U30231 ( .A(n32703), .B(n32704), .Z(n30052) );
  XOR U30232 ( .A(n30022), .B(n30057), .Z(n30056) );
  AND U30233 ( .A(n32705), .B(n32706), .Z(n30057) );
  XNOR U30234 ( .A(n30051), .B(n30023), .Z(n30022) );
  AND U30235 ( .A(n32707), .B(n32708), .Z(n30023) );
  XOR U30236 ( .A(n30050), .B(n30040), .Z(n30051) );
  AND U30237 ( .A(n32709), .B(n32710), .Z(n30040) );
  XNOR U30238 ( .A(n30045), .B(n30039), .Z(n30050) );
  AND U30239 ( .A(n32711), .B(n32712), .Z(n30039) );
  XOR U30240 ( .A(n29982), .B(n30046), .Z(n30045) );
  AND U30241 ( .A(n32713), .B(n32714), .Z(n30046) );
  XNOR U30242 ( .A(n30038), .B(n29983), .Z(n29982) );
  AND U30243 ( .A(n32715), .B(n32716), .Z(n29983) );
  XOR U30244 ( .A(n30037), .B(n30025), .Z(n30038) );
  AND U30245 ( .A(n32717), .B(n32718), .Z(n30025) );
  XNOR U30246 ( .A(n30032), .B(n30024), .Z(n30037) );
  AND U30247 ( .A(n32719), .B(n32720), .Z(n30024) );
  XOR U30248 ( .A(n29986), .B(n30033), .Z(n30032) );
  AND U30249 ( .A(n32721), .B(n32722), .Z(n30033) );
  XNOR U30250 ( .A(n30017), .B(n29987), .Z(n29986) );
  AND U30251 ( .A(n32723), .B(n32724), .Z(n29987) );
  XOR U30252 ( .A(n30016), .B(n30008), .Z(n30017) );
  AND U30253 ( .A(n32725), .B(n32726), .Z(n30008) );
  XNOR U30254 ( .A(n30011), .B(n30007), .Z(n30016) );
  AND U30255 ( .A(n32727), .B(n32728), .Z(n30007) );
  XOR U30256 ( .A(n29988), .B(n30012), .Z(n30011) );
  AND U30257 ( .A(n32729), .B(n32730), .Z(n30012) );
  XNOR U30258 ( .A(n30004), .B(n29989), .Z(n29988) );
  AND U30259 ( .A(n32731), .B(n32732), .Z(n29989) );
  XOR U30260 ( .A(n30003), .B(n29995), .Z(n30004) );
  AND U30261 ( .A(n32733), .B(n32734), .Z(n29995) );
  XNOR U30262 ( .A(n29998), .B(n29994), .Z(n30003) );
  AND U30263 ( .A(n32735), .B(n32736), .Z(n29994) );
  XOR U30264 ( .A(n29939), .B(n29999), .Z(n29998) );
  AND U30265 ( .A(n32737), .B(n32738), .Z(n29999) );
  XNOR U30266 ( .A(n29981), .B(n29940), .Z(n29939) );
  AND U30267 ( .A(n32739), .B(n32740), .Z(n29940) );
  XOR U30268 ( .A(n29980), .B(n29972), .Z(n29981) );
  AND U30269 ( .A(n32741), .B(n32742), .Z(n29972) );
  XNOR U30270 ( .A(n29975), .B(n29971), .Z(n29980) );
  AND U30271 ( .A(n32743), .B(n32744), .Z(n29971) );
  XOR U30272 ( .A(n29943), .B(n29976), .Z(n29975) );
  AND U30273 ( .A(n32745), .B(n32746), .Z(n29976) );
  XNOR U30274 ( .A(n29968), .B(n29944), .Z(n29943) );
  AND U30275 ( .A(n32747), .B(n32748), .Z(n29944) );
  XOR U30276 ( .A(n29967), .B(n29959), .Z(n29968) );
  AND U30277 ( .A(n32749), .B(n32750), .Z(n29959) );
  XNOR U30278 ( .A(n29962), .B(n29958), .Z(n29967) );
  AND U30279 ( .A(n32751), .B(n32752), .Z(n29958) );
  XOR U30280 ( .A(n29892), .B(n29963), .Z(n29962) );
  AND U30281 ( .A(n32753), .B(n32754), .Z(n29963) );
  XNOR U30282 ( .A(n29953), .B(n29893), .Z(n29892) );
  AND U30283 ( .A(n32755), .B(n32756), .Z(n29893) );
  XOR U30284 ( .A(n29952), .B(n29938), .Z(n29953) );
  AND U30285 ( .A(n32757), .B(n32758), .Z(n29938) );
  XNOR U30286 ( .A(n29947), .B(n29937), .Z(n29952) );
  AND U30287 ( .A(n32759), .B(n32760), .Z(n29937) );
  XOR U30288 ( .A(n29894), .B(n29948), .Z(n29947) );
  AND U30289 ( .A(n32761), .B(n32762), .Z(n29948) );
  XNOR U30290 ( .A(n29936), .B(n29895), .Z(n29894) );
  AND U30291 ( .A(n32763), .B(n32764), .Z(n29895) );
  XOR U30292 ( .A(n29935), .B(n29925), .Z(n29936) );
  AND U30293 ( .A(n32765), .B(n32766), .Z(n29925) );
  XNOR U30294 ( .A(n29930), .B(n29924), .Z(n29935) );
  AND U30295 ( .A(n32767), .B(n32768), .Z(n29924) );
  XOR U30296 ( .A(n32769), .B(n29923), .Z(n29930) );
  XOR U30297 ( .A(n29922), .B(n29910), .Z(n29923) );
  AND U30298 ( .A(n32770), .B(n32771), .Z(n29910) );
  XNOR U30299 ( .A(n29917), .B(n29909), .Z(n29922) );
  AND U30300 ( .A(n32772), .B(n32773), .Z(n29909) );
  XOR U30301 ( .A(n32774), .B(n32775), .Z(n29917) );
  XOR U30302 ( .A(n29907), .B(n32776), .Z(n32775) );
  XOR U30303 ( .A(n29903), .B(n29901), .Z(n32776) );
  AND U30304 ( .A(n32777), .B(n32778), .Z(n29901) );
  AND U30305 ( .A(n32779), .B(n32780), .Z(n29903) );
  AND U30306 ( .A(n32781), .B(n32782), .Z(n29907) );
  XNOR U30307 ( .A(n32783), .B(n29904), .Z(n32774) );
  XOR U30308 ( .A(n32784), .B(n32785), .Z(n29904) );
  XOR U30309 ( .A(n32786), .B(n32787), .Z(n32785) );
  XOR U30310 ( .A(n32788), .B(n32789), .Z(n32787) );
  NOR U30311 ( .A(n32790), .B(n32791), .Z(n32789) );
  NOR U30312 ( .A(n32792), .B(n32793), .Z(n32788) );
  AND U30313 ( .A(n32794), .B(n32795), .Z(n32793) );
  IV U30314 ( .A(n32796), .Z(n32792) );
  NOR U30315 ( .A(n32797), .B(n32798), .Z(n32796) );
  AND U30316 ( .A(n32790), .B(n32799), .Z(n32798) );
  AND U30317 ( .A(n32791), .B(n32800), .Z(n32797) );
  NOR U30318 ( .A(n32801), .B(n32802), .Z(n32786) );
  AND U30319 ( .A(n32803), .B(n32804), .Z(n32802) );
  IV U30320 ( .A(n32805), .Z(n32801) );
  NOR U30321 ( .A(n32806), .B(n32807), .Z(n32805) );
  AND U30322 ( .A(n32808), .B(n32809), .Z(n32807) );
  AND U30323 ( .A(n32810), .B(n32811), .Z(n32806) );
  XOR U30324 ( .A(n32812), .B(n32813), .Z(n32784) );
  XOR U30325 ( .A(n32814), .B(n32815), .Z(n32813) );
  XOR U30326 ( .A(n32816), .B(n32817), .Z(n32815) );
  XOR U30327 ( .A(n32818), .B(n32819), .Z(n32817) );
  AND U30328 ( .A(n32820), .B(n32821), .Z(n32819) );
  AND U30329 ( .A(n32822), .B(n32823), .Z(n32818) );
  XOR U30330 ( .A(n32824), .B(n32825), .Z(n32816) );
  AND U30331 ( .A(n32826), .B(n32827), .Z(n32825) );
  AND U30332 ( .A(n32828), .B(n32829), .Z(n32824) );
  AND U30333 ( .A(n32830), .B(n32831), .Z(n32829) );
  AND U30334 ( .A(n32832), .B(n32833), .Z(n32831) );
  NOR U30335 ( .A(n32834), .B(n32835), .Z(n32833) );
  IV U30336 ( .A(n32836), .Z(n32834) );
  NOR U30337 ( .A(n32837), .B(n32838), .Z(n32836) );
  NOR U30338 ( .A(n32839), .B(n32840), .Z(n32832) );
  AND U30339 ( .A(n32841), .B(n32842), .Z(n32830) );
  NOR U30340 ( .A(n32843), .B(n32844), .Z(n32842) );
  NOR U30341 ( .A(n32845), .B(n32846), .Z(n32841) );
  AND U30342 ( .A(n32847), .B(n32848), .Z(n32828) );
  AND U30343 ( .A(n32849), .B(n32850), .Z(n32848) );
  NOR U30344 ( .A(n32851), .B(n32852), .Z(n32850) );
  NOR U30345 ( .A(n32853), .B(n32854), .Z(n32849) );
  AND U30346 ( .A(n32855), .B(n32856), .Z(n32847) );
  NOR U30347 ( .A(n32857), .B(n32858), .Z(n32856) );
  NOR U30348 ( .A(n32859), .B(n32860), .Z(n32855) );
  XOR U30349 ( .A(n32861), .B(n32862), .Z(n32814) );
  XOR U30350 ( .A(n32863), .B(n32864), .Z(n32862) );
  NOR U30351 ( .A(n32865), .B(n32866), .Z(n32864) );
  NOR U30352 ( .A(n32867), .B(n32868), .Z(n32863) );
  AND U30353 ( .A(n32869), .B(n32870), .Z(n32868) );
  IV U30354 ( .A(n32871), .Z(n32867) );
  NOR U30355 ( .A(n32872), .B(n32873), .Z(n32871) );
  AND U30356 ( .A(n32865), .B(n32874), .Z(n32873) );
  AND U30357 ( .A(n32866), .B(n32875), .Z(n32872) );
  XOR U30358 ( .A(n32876), .B(n32877), .Z(n32861) );
  NOR U30359 ( .A(n32878), .B(n32879), .Z(n32877) );
  NOR U30360 ( .A(n32880), .B(n32881), .Z(n32876) );
  AND U30361 ( .A(n32882), .B(n32883), .Z(n32881) );
  IV U30362 ( .A(n32884), .Z(n32880) );
  NOR U30363 ( .A(n32885), .B(n32886), .Z(n32884) );
  AND U30364 ( .A(n32878), .B(n32887), .Z(n32886) );
  AND U30365 ( .A(n32879), .B(n32888), .Z(n32885) );
  XNOR U30366 ( .A(n32889), .B(n32890), .Z(n32812) );
  AND U30367 ( .A(n32891), .B(n32892), .Z(n32890) );
  NOR U30368 ( .A(n32808), .B(n32810), .Z(n32889) );
  XNOR U30369 ( .A(n29908), .B(n29918), .Z(n32783) );
  AND U30370 ( .A(n32893), .B(n32894), .Z(n29918) );
  AND U30371 ( .A(n32895), .B(n32896), .Z(n29908) );
  XOR U30372 ( .A(n29906), .B(n29931), .Z(n32769) );
  AND U30373 ( .A(n32897), .B(n32898), .Z(n29931) );
  IV U30374 ( .A(n32899), .Z(n29906) );
  AND U30375 ( .A(n32900), .B(n32901), .Z(n32899) );
  XOR U30376 ( .A(n32902), .B(n32903), .Z(n30081) );
  AND U30377 ( .A(n32902), .B(n32904), .Z(n32903) );
  XOR U30378 ( .A(n32905), .B(n32906), .Z(n30078) );
  AND U30379 ( .A(n32905), .B(n32907), .Z(n32906) );
  XOR U30380 ( .A(n32908), .B(n32909), .Z(n29860) );
  AND U30381 ( .A(n32908), .B(n32910), .Z(n32909) );
  XOR U30382 ( .A(n32911), .B(n32912), .Z(n30098) );
  AND U30383 ( .A(n32911), .B(n32913), .Z(n32912) );
  XNOR U30384 ( .A(n32914), .B(n32915), .Z(n30093) );
  AND U30385 ( .A(n32914), .B(n32916), .Z(n32915) );
  XNOR U30386 ( .A(n32917), .B(n32918), .Z(n30094) );
  AND U30387 ( .A(n32919), .B(n32917), .Z(n32918) );
  XOR U30388 ( .A(n32920), .B(n32921), .Z(n29857) );
  NOR U30389 ( .A(n32922), .B(n32920), .Z(n32921) );
  XOR U30390 ( .A(n32923), .B(n32924), .Z(n30109) );
  NOR U30391 ( .A(n32925), .B(n32923), .Z(n32924) );
  XOR U30392 ( .A(n32926), .B(n32927), .Z(n30104) );
  NOR U30393 ( .A(n32928), .B(n32926), .Z(n32927) );
  XOR U30394 ( .A(n32929), .B(n32930), .Z(n30105) );
  NOR U30395 ( .A(n32931), .B(n32929), .Z(n32930) );
  XOR U30396 ( .A(n32932), .B(n32933), .Z(n29850) );
  NOR U30397 ( .A(n32934), .B(n32932), .Z(n32933) );
  XOR U30398 ( .A(n32935), .B(n32936), .Z(n29824) );
  NOR U30399 ( .A(n32937), .B(n32935), .Z(n32936) );
  XOR U30400 ( .A(n32938), .B(n32939), .Z(n29829) );
  NOR U30401 ( .A(n32940), .B(n32938), .Z(n32939) );
  XOR U30402 ( .A(n32941), .B(n32942), .Z(n29831) );
  NOR U30403 ( .A(n32943), .B(n32941), .Z(n32942) );
  IV U30404 ( .A(n29841), .Z(n32688) );
  XNOR U30405 ( .A(n32944), .B(n32945), .Z(n29841) );
  NOR U30406 ( .A(n32946), .B(n32944), .Z(n32945) );
  XOR U30407 ( .A(n32947), .B(n32948), .Z(n30115) );
  NOR U30408 ( .A(n32949), .B(n32947), .Z(n32948) );
  XOR U30409 ( .A(n32950), .B(n32951), .Z(n30118) );
  NOR U30410 ( .A(n32952), .B(n32950), .Z(n32951) );
  XOR U30411 ( .A(n32953), .B(n32954), .Z(n30121) );
  NOR U30412 ( .A(n32955), .B(n32953), .Z(n32954) );
  XOR U30413 ( .A(n32956), .B(n32957), .Z(n30124) );
  NOR U30414 ( .A(n32958), .B(n32956), .Z(n32957) );
  XOR U30415 ( .A(n32959), .B(n32960), .Z(n30127) );
  NOR U30416 ( .A(n32961), .B(n32959), .Z(n32960) );
  XOR U30417 ( .A(n32962), .B(n32963), .Z(n30130) );
  NOR U30418 ( .A(n32964), .B(n32962), .Z(n32963) );
  XOR U30419 ( .A(n32965), .B(n32966), .Z(n30133) );
  NOR U30420 ( .A(n32967), .B(n32965), .Z(n32966) );
  XOR U30421 ( .A(n32968), .B(n32969), .Z(n30136) );
  NOR U30422 ( .A(n32970), .B(n32968), .Z(n32969) );
  XOR U30423 ( .A(n32971), .B(n32972), .Z(n30139) );
  NOR U30424 ( .A(n32973), .B(n32971), .Z(n32972) );
  XOR U30425 ( .A(n32974), .B(n32975), .Z(n30142) );
  NOR U30426 ( .A(n32976), .B(n32974), .Z(n32975) );
  XOR U30427 ( .A(n32977), .B(n32978), .Z(n30145) );
  NOR U30428 ( .A(n32979), .B(n32977), .Z(n32978) );
  XOR U30429 ( .A(n32980), .B(n32981), .Z(n30148) );
  NOR U30430 ( .A(n32982), .B(n32980), .Z(n32981) );
  XOR U30431 ( .A(n32983), .B(n32984), .Z(n30151) );
  NOR U30432 ( .A(n32985), .B(n32983), .Z(n32984) );
  XOR U30433 ( .A(n32986), .B(n32987), .Z(n30154) );
  NOR U30434 ( .A(n32988), .B(n32986), .Z(n32987) );
  XOR U30435 ( .A(n32989), .B(n32990), .Z(n30157) );
  NOR U30436 ( .A(n32991), .B(n32989), .Z(n32990) );
  XOR U30437 ( .A(n32992), .B(n32993), .Z(n30160) );
  NOR U30438 ( .A(n32994), .B(n32992), .Z(n32993) );
  XOR U30439 ( .A(n32995), .B(n32996), .Z(n30163) );
  NOR U30440 ( .A(n32997), .B(n32995), .Z(n32996) );
  XOR U30441 ( .A(n32998), .B(n32999), .Z(n30166) );
  NOR U30442 ( .A(n33000), .B(n32998), .Z(n32999) );
  XOR U30443 ( .A(n33001), .B(n33002), .Z(n30169) );
  NOR U30444 ( .A(n33003), .B(n33001), .Z(n33002) );
  XOR U30445 ( .A(n33004), .B(n33005), .Z(n30172) );
  NOR U30446 ( .A(n33006), .B(n33004), .Z(n33005) );
  XOR U30447 ( .A(n33007), .B(n33008), .Z(n30175) );
  NOR U30448 ( .A(n33009), .B(n33007), .Z(n33008) );
  XOR U30449 ( .A(n33010), .B(n33011), .Z(n30178) );
  NOR U30450 ( .A(n33012), .B(n33010), .Z(n33011) );
  XOR U30451 ( .A(n33013), .B(n33014), .Z(n30181) );
  NOR U30452 ( .A(n33015), .B(n33013), .Z(n33014) );
  XOR U30453 ( .A(n33016), .B(n33017), .Z(n30184) );
  NOR U30454 ( .A(n33018), .B(n33016), .Z(n33017) );
  XOR U30455 ( .A(n33019), .B(n33020), .Z(n30187) );
  NOR U30456 ( .A(n33021), .B(n33019), .Z(n33020) );
  XOR U30457 ( .A(n33022), .B(n33023), .Z(n30190) );
  NOR U30458 ( .A(n33024), .B(n33022), .Z(n33023) );
  XOR U30459 ( .A(n33025), .B(n33026), .Z(n30193) );
  NOR U30460 ( .A(n33027), .B(n33025), .Z(n33026) );
  XOR U30461 ( .A(n33028), .B(n33029), .Z(n30196) );
  NOR U30462 ( .A(n33030), .B(n33028), .Z(n33029) );
  XOR U30463 ( .A(n33031), .B(n33032), .Z(n30199) );
  NOR U30464 ( .A(n33033), .B(n33031), .Z(n33032) );
  XOR U30465 ( .A(n33034), .B(n33035), .Z(n30202) );
  NOR U30466 ( .A(n33036), .B(n33034), .Z(n33035) );
  XOR U30467 ( .A(n33037), .B(n33038), .Z(n30205) );
  NOR U30468 ( .A(n33039), .B(n33037), .Z(n33038) );
  XOR U30469 ( .A(n33040), .B(n33041), .Z(n30208) );
  NOR U30470 ( .A(n33042), .B(n33040), .Z(n33041) );
  XOR U30471 ( .A(n33043), .B(n33044), .Z(n30211) );
  NOR U30472 ( .A(n33045), .B(n33043), .Z(n33044) );
  XOR U30473 ( .A(n33046), .B(n33047), .Z(n30214) );
  NOR U30474 ( .A(n33048), .B(n33046), .Z(n33047) );
  XOR U30475 ( .A(n33049), .B(n33050), .Z(n30217) );
  NOR U30476 ( .A(n33051), .B(n33049), .Z(n33050) );
  XOR U30477 ( .A(n33052), .B(n33053), .Z(n30220) );
  NOR U30478 ( .A(n33054), .B(n33052), .Z(n33053) );
  XOR U30479 ( .A(n33055), .B(n33056), .Z(n30223) );
  NOR U30480 ( .A(n33057), .B(n33055), .Z(n33056) );
  XOR U30481 ( .A(n33058), .B(n33059), .Z(n30226) );
  NOR U30482 ( .A(n33060), .B(n33058), .Z(n33059) );
  XOR U30483 ( .A(n33061), .B(n33062), .Z(n30229) );
  NOR U30484 ( .A(n33063), .B(n33061), .Z(n33062) );
  XOR U30485 ( .A(n33064), .B(n33065), .Z(n30232) );
  NOR U30486 ( .A(n33066), .B(n33064), .Z(n33065) );
  XOR U30487 ( .A(n33067), .B(n33068), .Z(n30235) );
  NOR U30488 ( .A(n33069), .B(n33067), .Z(n33068) );
  XOR U30489 ( .A(n33070), .B(n33071), .Z(n30238) );
  NOR U30490 ( .A(n33072), .B(n33070), .Z(n33071) );
  XOR U30491 ( .A(n33073), .B(n33074), .Z(n30241) );
  NOR U30492 ( .A(n33075), .B(n33073), .Z(n33074) );
  XOR U30493 ( .A(n33076), .B(n33077), .Z(n30244) );
  NOR U30494 ( .A(n33078), .B(n33076), .Z(n33077) );
  XOR U30495 ( .A(n33079), .B(n33080), .Z(n30247) );
  NOR U30496 ( .A(n33081), .B(n33079), .Z(n33080) );
  XOR U30497 ( .A(n33082), .B(n33083), .Z(n30250) );
  NOR U30498 ( .A(n33084), .B(n33082), .Z(n33083) );
  XOR U30499 ( .A(n33085), .B(n33086), .Z(n30253) );
  NOR U30500 ( .A(n33087), .B(n33085), .Z(n33086) );
  XOR U30501 ( .A(n33088), .B(n33089), .Z(n30256) );
  NOR U30502 ( .A(n33090), .B(n33088), .Z(n33089) );
  XOR U30503 ( .A(n33091), .B(n33092), .Z(n30259) );
  NOR U30504 ( .A(n33093), .B(n33091), .Z(n33092) );
  XOR U30505 ( .A(n33094), .B(n33095), .Z(n30262) );
  NOR U30506 ( .A(n33096), .B(n33094), .Z(n33095) );
  XOR U30507 ( .A(n33097), .B(n33098), .Z(n30265) );
  NOR U30508 ( .A(n33099), .B(n33097), .Z(n33098) );
  XOR U30509 ( .A(n33100), .B(n33101), .Z(n30268) );
  NOR U30510 ( .A(n33102), .B(n33100), .Z(n33101) );
  XOR U30511 ( .A(n33103), .B(n33104), .Z(n30271) );
  NOR U30512 ( .A(n33105), .B(n33103), .Z(n33104) );
  XOR U30513 ( .A(n33106), .B(n33107), .Z(n30274) );
  NOR U30514 ( .A(n33108), .B(n33106), .Z(n33107) );
  XOR U30515 ( .A(n33109), .B(n33110), .Z(n30277) );
  NOR U30516 ( .A(n33111), .B(n33109), .Z(n33110) );
  XOR U30517 ( .A(n33112), .B(n33113), .Z(n30280) );
  NOR U30518 ( .A(n33114), .B(n33112), .Z(n33113) );
  XOR U30519 ( .A(n33115), .B(n33116), .Z(n30283) );
  NOR U30520 ( .A(n33117), .B(n33115), .Z(n33116) );
  XOR U30521 ( .A(n33118), .B(n33119), .Z(n30286) );
  NOR U30522 ( .A(n33120), .B(n33118), .Z(n33119) );
  XOR U30523 ( .A(n33121), .B(n33122), .Z(n30289) );
  NOR U30524 ( .A(n33123), .B(n33121), .Z(n33122) );
  XOR U30525 ( .A(n33124), .B(n33125), .Z(n30292) );
  NOR U30526 ( .A(n33126), .B(n33124), .Z(n33125) );
  XOR U30527 ( .A(n33127), .B(n33128), .Z(n30295) );
  NOR U30528 ( .A(n33129), .B(n33127), .Z(n33128) );
  XOR U30529 ( .A(n33130), .B(n33131), .Z(n30298) );
  NOR U30530 ( .A(n33132), .B(n33130), .Z(n33131) );
  XOR U30531 ( .A(n33133), .B(n33134), .Z(n30301) );
  NOR U30532 ( .A(n33135), .B(n33133), .Z(n33134) );
  XOR U30533 ( .A(n33136), .B(n33137), .Z(n30304) );
  NOR U30534 ( .A(n33138), .B(n33136), .Z(n33137) );
  XOR U30535 ( .A(n33139), .B(n33140), .Z(n30307) );
  NOR U30536 ( .A(n33141), .B(n33139), .Z(n33140) );
  XOR U30537 ( .A(n33142), .B(n33143), .Z(n30310) );
  NOR U30538 ( .A(n33144), .B(n33142), .Z(n33143) );
  XOR U30539 ( .A(n33145), .B(n33146), .Z(n30313) );
  NOR U30540 ( .A(n33147), .B(n33145), .Z(n33146) );
  XOR U30541 ( .A(n33148), .B(n33149), .Z(n30316) );
  NOR U30542 ( .A(n33150), .B(n33148), .Z(n33149) );
  XOR U30543 ( .A(n33151), .B(n33152), .Z(n30319) );
  NOR U30544 ( .A(n33153), .B(n33151), .Z(n33152) );
  XOR U30545 ( .A(n33154), .B(n33155), .Z(n30322) );
  NOR U30546 ( .A(n33156), .B(n33154), .Z(n33155) );
  XOR U30547 ( .A(n33157), .B(n33158), .Z(n30325) );
  NOR U30548 ( .A(n33159), .B(n33157), .Z(n33158) );
  XOR U30549 ( .A(n33160), .B(n33161), .Z(n30328) );
  NOR U30550 ( .A(n33162), .B(n33160), .Z(n33161) );
  XOR U30551 ( .A(n33163), .B(n33164), .Z(n30331) );
  NOR U30552 ( .A(n33165), .B(n33163), .Z(n33164) );
  XOR U30553 ( .A(n33166), .B(n33167), .Z(n30334) );
  NOR U30554 ( .A(n33168), .B(n33166), .Z(n33167) );
  XOR U30555 ( .A(n33169), .B(n33170), .Z(n30337) );
  NOR U30556 ( .A(n33171), .B(n33169), .Z(n33170) );
  XOR U30557 ( .A(n33172), .B(n33173), .Z(n30340) );
  NOR U30558 ( .A(n33174), .B(n33172), .Z(n33173) );
  XOR U30559 ( .A(n33175), .B(n33176), .Z(n30343) );
  NOR U30560 ( .A(n33177), .B(n33175), .Z(n33176) );
  XOR U30561 ( .A(n33178), .B(n33179), .Z(n30346) );
  NOR U30562 ( .A(n33180), .B(n33178), .Z(n33179) );
  XOR U30563 ( .A(n33181), .B(n33182), .Z(n30349) );
  NOR U30564 ( .A(n33183), .B(n33181), .Z(n33182) );
  XOR U30565 ( .A(n33184), .B(n33185), .Z(n30352) );
  NOR U30566 ( .A(n33186), .B(n33184), .Z(n33185) );
  XOR U30567 ( .A(n33187), .B(n33188), .Z(n30355) );
  NOR U30568 ( .A(n33189), .B(n33187), .Z(n33188) );
  XOR U30569 ( .A(n33190), .B(n33191), .Z(n30358) );
  NOR U30570 ( .A(n33192), .B(n33190), .Z(n33191) );
  XOR U30571 ( .A(n33193), .B(n33194), .Z(n30361) );
  NOR U30572 ( .A(n33195), .B(n33193), .Z(n33194) );
  XOR U30573 ( .A(n33196), .B(n33197), .Z(n30364) );
  NOR U30574 ( .A(n33198), .B(n33196), .Z(n33197) );
  XOR U30575 ( .A(n33199), .B(n33200), .Z(n30367) );
  NOR U30576 ( .A(n33201), .B(n33199), .Z(n33200) );
  XOR U30577 ( .A(n33202), .B(n33203), .Z(n30370) );
  NOR U30578 ( .A(n33204), .B(n33202), .Z(n33203) );
  XOR U30579 ( .A(n33205), .B(n33206), .Z(n30373) );
  NOR U30580 ( .A(n33207), .B(n33205), .Z(n33206) );
  XOR U30581 ( .A(n33208), .B(n33209), .Z(n30376) );
  NOR U30582 ( .A(n33210), .B(n33208), .Z(n33209) );
  XOR U30583 ( .A(n33211), .B(n33212), .Z(n30379) );
  NOR U30584 ( .A(n33213), .B(n33211), .Z(n33212) );
  XOR U30585 ( .A(n33214), .B(n33215), .Z(n30382) );
  NOR U30586 ( .A(n33216), .B(n33214), .Z(n33215) );
  XOR U30587 ( .A(n33217), .B(n33218), .Z(n30385) );
  NOR U30588 ( .A(n33219), .B(n33217), .Z(n33218) );
  XOR U30589 ( .A(n33220), .B(n33221), .Z(n30388) );
  NOR U30590 ( .A(n33222), .B(n33220), .Z(n33221) );
  XOR U30591 ( .A(n33223), .B(n33224), .Z(n30391) );
  NOR U30592 ( .A(n33225), .B(n33223), .Z(n33224) );
  XOR U30593 ( .A(n33226), .B(n33227), .Z(n30394) );
  NOR U30594 ( .A(n33228), .B(n33226), .Z(n33227) );
  XOR U30595 ( .A(n33229), .B(n33230), .Z(n30397) );
  NOR U30596 ( .A(n33231), .B(n33229), .Z(n33230) );
  XOR U30597 ( .A(n33232), .B(n33233), .Z(n30400) );
  NOR U30598 ( .A(n33234), .B(n33232), .Z(n33233) );
  XOR U30599 ( .A(n33235), .B(n33236), .Z(n30403) );
  NOR U30600 ( .A(n33237), .B(n33235), .Z(n33236) );
  XOR U30601 ( .A(n33238), .B(n33239), .Z(n30406) );
  NOR U30602 ( .A(n33240), .B(n33238), .Z(n33239) );
  XOR U30603 ( .A(n33241), .B(n33242), .Z(n30409) );
  NOR U30604 ( .A(n33243), .B(n33241), .Z(n33242) );
  XOR U30605 ( .A(n33244), .B(n33245), .Z(n30412) );
  NOR U30606 ( .A(n33246), .B(n33244), .Z(n33245) );
  XOR U30607 ( .A(n33247), .B(n33248), .Z(n30415) );
  NOR U30608 ( .A(n33249), .B(n33247), .Z(n33248) );
  XOR U30609 ( .A(n33250), .B(n33251), .Z(n30418) );
  NOR U30610 ( .A(n33252), .B(n33250), .Z(n33251) );
  XOR U30611 ( .A(n33253), .B(n33254), .Z(n30421) );
  NOR U30612 ( .A(n33255), .B(n33253), .Z(n33254) );
  XOR U30613 ( .A(n33256), .B(n33257), .Z(n30424) );
  NOR U30614 ( .A(n33258), .B(n33256), .Z(n33257) );
  XOR U30615 ( .A(n33259), .B(n33260), .Z(n30427) );
  NOR U30616 ( .A(n33261), .B(n33259), .Z(n33260) );
  XOR U30617 ( .A(n33262), .B(n33263), .Z(n30430) );
  NOR U30618 ( .A(n33264), .B(n33262), .Z(n33263) );
  XOR U30619 ( .A(n33265), .B(n33266), .Z(n30433) );
  NOR U30620 ( .A(n33267), .B(n33265), .Z(n33266) );
  XOR U30621 ( .A(n33268), .B(n33269), .Z(n30436) );
  NOR U30622 ( .A(n33270), .B(n33268), .Z(n33269) );
  XOR U30623 ( .A(n33271), .B(n33272), .Z(n30439) );
  NOR U30624 ( .A(n33273), .B(n33271), .Z(n33272) );
  XOR U30625 ( .A(n33274), .B(n33275), .Z(n30442) );
  NOR U30626 ( .A(n33276), .B(n33274), .Z(n33275) );
  XOR U30627 ( .A(n33277), .B(n33278), .Z(n30445) );
  NOR U30628 ( .A(n33279), .B(n33277), .Z(n33278) );
  XOR U30629 ( .A(n33280), .B(n33281), .Z(n30448) );
  NOR U30630 ( .A(n33282), .B(n33280), .Z(n33281) );
  XOR U30631 ( .A(n33283), .B(n33284), .Z(n30451) );
  NOR U30632 ( .A(n33285), .B(n33283), .Z(n33284) );
  XOR U30633 ( .A(n33286), .B(n33287), .Z(n30454) );
  NOR U30634 ( .A(n33288), .B(n33286), .Z(n33287) );
  XOR U30635 ( .A(n33289), .B(n33290), .Z(n30457) );
  NOR U30636 ( .A(n33291), .B(n33289), .Z(n33290) );
  XOR U30637 ( .A(n33292), .B(n33293), .Z(n30460) );
  NOR U30638 ( .A(n33294), .B(n33292), .Z(n33293) );
  XOR U30639 ( .A(n33295), .B(n33296), .Z(n30463) );
  NOR U30640 ( .A(n33297), .B(n33295), .Z(n33296) );
  XOR U30641 ( .A(n33298), .B(n33299), .Z(n30466) );
  NOR U30642 ( .A(n33300), .B(n33298), .Z(n33299) );
  XOR U30643 ( .A(n33301), .B(n33302), .Z(n30469) );
  NOR U30644 ( .A(n33303), .B(n33301), .Z(n33302) );
  XOR U30645 ( .A(n33304), .B(n33305), .Z(n30472) );
  NOR U30646 ( .A(n33306), .B(n33304), .Z(n33305) );
  XOR U30647 ( .A(n33307), .B(n33308), .Z(n30475) );
  NOR U30648 ( .A(n33309), .B(n33307), .Z(n33308) );
  XOR U30649 ( .A(n33310), .B(n33311), .Z(n30478) );
  NOR U30650 ( .A(n33312), .B(n33310), .Z(n33311) );
  XOR U30651 ( .A(n33313), .B(n33314), .Z(n30481) );
  NOR U30652 ( .A(n33315), .B(n33313), .Z(n33314) );
  XOR U30653 ( .A(n33316), .B(n33317), .Z(n30484) );
  NOR U30654 ( .A(n33318), .B(n33316), .Z(n33317) );
  XOR U30655 ( .A(n33319), .B(n33320), .Z(n30487) );
  NOR U30656 ( .A(n33321), .B(n33319), .Z(n33320) );
  XOR U30657 ( .A(n33322), .B(n33323), .Z(n30490) );
  NOR U30658 ( .A(n33324), .B(n33322), .Z(n33323) );
  XOR U30659 ( .A(n33325), .B(n33326), .Z(n30493) );
  NOR U30660 ( .A(n33327), .B(n33325), .Z(n33326) );
  XOR U30661 ( .A(n33328), .B(n33329), .Z(n30496) );
  NOR U30662 ( .A(n33330), .B(n33328), .Z(n33329) );
  XOR U30663 ( .A(n33331), .B(n33332), .Z(n30499) );
  NOR U30664 ( .A(n33333), .B(n33331), .Z(n33332) );
  XOR U30665 ( .A(n33334), .B(n33335), .Z(n30502) );
  NOR U30666 ( .A(n33336), .B(n33334), .Z(n33335) );
  XOR U30667 ( .A(n33337), .B(n33338), .Z(n30505) );
  NOR U30668 ( .A(n33339), .B(n33337), .Z(n33338) );
  XOR U30669 ( .A(n33340), .B(n33341), .Z(n30508) );
  NOR U30670 ( .A(n33342), .B(n33340), .Z(n33341) );
  XOR U30671 ( .A(n33343), .B(n33344), .Z(n30511) );
  NOR U30672 ( .A(n33345), .B(n33343), .Z(n33344) );
  XOR U30673 ( .A(n33346), .B(n33347), .Z(n30514) );
  NOR U30674 ( .A(n33348), .B(n33346), .Z(n33347) );
  XOR U30675 ( .A(n33349), .B(n33350), .Z(n30517) );
  NOR U30676 ( .A(n33351), .B(n33349), .Z(n33350) );
  XOR U30677 ( .A(n33352), .B(n33353), .Z(n30520) );
  NOR U30678 ( .A(n33354), .B(n33352), .Z(n33353) );
  XOR U30679 ( .A(n33355), .B(n33356), .Z(n30523) );
  NOR U30680 ( .A(n33357), .B(n33355), .Z(n33356) );
  XOR U30681 ( .A(n33358), .B(n33359), .Z(n30526) );
  NOR U30682 ( .A(n33360), .B(n33358), .Z(n33359) );
  XOR U30683 ( .A(n33361), .B(n33362), .Z(n30529) );
  NOR U30684 ( .A(n33363), .B(n33361), .Z(n33362) );
  XOR U30685 ( .A(n33364), .B(n33365), .Z(n30532) );
  NOR U30686 ( .A(n33366), .B(n33364), .Z(n33365) );
  XOR U30687 ( .A(n33367), .B(n33368), .Z(n30535) );
  NOR U30688 ( .A(n33369), .B(n33367), .Z(n33368) );
  XOR U30689 ( .A(n33370), .B(n33371), .Z(n30538) );
  NOR U30690 ( .A(n33372), .B(n33370), .Z(n33371) );
  XOR U30691 ( .A(n33373), .B(n33374), .Z(n30541) );
  NOR U30692 ( .A(n33375), .B(n33373), .Z(n33374) );
  XOR U30693 ( .A(n33376), .B(n33377), .Z(n30544) );
  NOR U30694 ( .A(n33378), .B(n33376), .Z(n33377) );
  XOR U30695 ( .A(n33379), .B(n33380), .Z(n30547) );
  NOR U30696 ( .A(n33381), .B(n33379), .Z(n33380) );
  XOR U30697 ( .A(n33382), .B(n33383), .Z(n30550) );
  NOR U30698 ( .A(n33384), .B(n33382), .Z(n33383) );
  XOR U30699 ( .A(n33385), .B(n33386), .Z(n30553) );
  NOR U30700 ( .A(n33387), .B(n33385), .Z(n33386) );
  XOR U30701 ( .A(n33388), .B(n33389), .Z(n30556) );
  NOR U30702 ( .A(n33390), .B(n33388), .Z(n33389) );
  XOR U30703 ( .A(n33391), .B(n33392), .Z(n30559) );
  NOR U30704 ( .A(n33393), .B(n33391), .Z(n33392) );
  XOR U30705 ( .A(n33394), .B(n33395), .Z(n30562) );
  NOR U30706 ( .A(n33396), .B(n33394), .Z(n33395) );
  XOR U30707 ( .A(n33397), .B(n33398), .Z(n30565) );
  NOR U30708 ( .A(n33399), .B(n33397), .Z(n33398) );
  XOR U30709 ( .A(n33400), .B(n33401), .Z(n30568) );
  NOR U30710 ( .A(n33402), .B(n33400), .Z(n33401) );
  XOR U30711 ( .A(n33403), .B(n33404), .Z(n30571) );
  NOR U30712 ( .A(n33405), .B(n33403), .Z(n33404) );
  XOR U30713 ( .A(n33406), .B(n33407), .Z(n30574) );
  NOR U30714 ( .A(n33408), .B(n33406), .Z(n33407) );
  XOR U30715 ( .A(n33409), .B(n33410), .Z(n30577) );
  NOR U30716 ( .A(n33411), .B(n33409), .Z(n33410) );
  XOR U30717 ( .A(n33412), .B(n33413), .Z(n30580) );
  NOR U30718 ( .A(n33414), .B(n33412), .Z(n33413) );
  XOR U30719 ( .A(n33415), .B(n33416), .Z(n30583) );
  NOR U30720 ( .A(n33417), .B(n33415), .Z(n33416) );
  XOR U30721 ( .A(n33418), .B(n33419), .Z(n30586) );
  NOR U30722 ( .A(n33420), .B(n33418), .Z(n33419) );
  XOR U30723 ( .A(n33421), .B(n33422), .Z(n30589) );
  NOR U30724 ( .A(n33423), .B(n33421), .Z(n33422) );
  XOR U30725 ( .A(n33424), .B(n33425), .Z(n30592) );
  NOR U30726 ( .A(n33426), .B(n33424), .Z(n33425) );
  XOR U30727 ( .A(n33427), .B(n33428), .Z(n30595) );
  NOR U30728 ( .A(n33429), .B(n33427), .Z(n33428) );
  XOR U30729 ( .A(n33430), .B(n33431), .Z(n30598) );
  NOR U30730 ( .A(n33432), .B(n33430), .Z(n33431) );
  XOR U30731 ( .A(n33433), .B(n33434), .Z(n30601) );
  NOR U30732 ( .A(n33435), .B(n33433), .Z(n33434) );
  XOR U30733 ( .A(n33436), .B(n33437), .Z(n30604) );
  NOR U30734 ( .A(n33438), .B(n33436), .Z(n33437) );
  XOR U30735 ( .A(n33439), .B(n33440), .Z(n30607) );
  NOR U30736 ( .A(n33441), .B(n33439), .Z(n33440) );
  XOR U30737 ( .A(n33442), .B(n33443), .Z(n30610) );
  NOR U30738 ( .A(n33444), .B(n33442), .Z(n33443) );
  XOR U30739 ( .A(n33445), .B(n33446), .Z(n30613) );
  NOR U30740 ( .A(n33447), .B(n33445), .Z(n33446) );
  XOR U30741 ( .A(n33448), .B(n33449), .Z(n30616) );
  NOR U30742 ( .A(n33450), .B(n33448), .Z(n33449) );
  XOR U30743 ( .A(n33451), .B(n33452), .Z(n30619) );
  NOR U30744 ( .A(n33453), .B(n33451), .Z(n33452) );
  XOR U30745 ( .A(n33454), .B(n33455), .Z(n30622) );
  NOR U30746 ( .A(n33456), .B(n33454), .Z(n33455) );
  XOR U30747 ( .A(n33457), .B(n33458), .Z(n30625) );
  NOR U30748 ( .A(n33459), .B(n33457), .Z(n33458) );
  XOR U30749 ( .A(n33460), .B(n33461), .Z(n30628) );
  NOR U30750 ( .A(n33462), .B(n33460), .Z(n33461) );
  XOR U30751 ( .A(n33463), .B(n33464), .Z(n30631) );
  NOR U30752 ( .A(n33465), .B(n33463), .Z(n33464) );
  XOR U30753 ( .A(n33466), .B(n33467), .Z(n30634) );
  NOR U30754 ( .A(n33468), .B(n33466), .Z(n33467) );
  XOR U30755 ( .A(n33469), .B(n33470), .Z(n30637) );
  NOR U30756 ( .A(n33471), .B(n33469), .Z(n33470) );
  XOR U30757 ( .A(n33472), .B(n33473), .Z(n30640) );
  NOR U30758 ( .A(n33474), .B(n33472), .Z(n33473) );
  XOR U30759 ( .A(n33475), .B(n33476), .Z(n30643) );
  NOR U30760 ( .A(n33477), .B(n33475), .Z(n33476) );
  XOR U30761 ( .A(n33478), .B(n33479), .Z(n30646) );
  NOR U30762 ( .A(n33480), .B(n33478), .Z(n33479) );
  XOR U30763 ( .A(n33481), .B(n33482), .Z(n30649) );
  NOR U30764 ( .A(n33483), .B(n33481), .Z(n33482) );
  XOR U30765 ( .A(n33484), .B(n33485), .Z(n30652) );
  NOR U30766 ( .A(n33486), .B(n33484), .Z(n33485) );
  XOR U30767 ( .A(n33487), .B(n33488), .Z(n30655) );
  NOR U30768 ( .A(n33489), .B(n33487), .Z(n33488) );
  XOR U30769 ( .A(n33490), .B(n33491), .Z(n30658) );
  NOR U30770 ( .A(n33492), .B(n33490), .Z(n33491) );
  XOR U30771 ( .A(n33493), .B(n33494), .Z(n30661) );
  NOR U30772 ( .A(n33495), .B(n33493), .Z(n33494) );
  XOR U30773 ( .A(n33496), .B(n33497), .Z(n30664) );
  NOR U30774 ( .A(n33498), .B(n33496), .Z(n33497) );
  XOR U30775 ( .A(n33499), .B(n33500), .Z(n30667) );
  NOR U30776 ( .A(n33501), .B(n33499), .Z(n33500) );
  XOR U30777 ( .A(n33502), .B(n33503), .Z(n30670) );
  NOR U30778 ( .A(n33504), .B(n33502), .Z(n33503) );
  XOR U30779 ( .A(n33505), .B(n33506), .Z(n30673) );
  NOR U30780 ( .A(n33507), .B(n33505), .Z(n33506) );
  XOR U30781 ( .A(n33508), .B(n33509), .Z(n30676) );
  NOR U30782 ( .A(n33510), .B(n33508), .Z(n33509) );
  XOR U30783 ( .A(n33511), .B(n33512), .Z(n30679) );
  NOR U30784 ( .A(n33513), .B(n33511), .Z(n33512) );
  XOR U30785 ( .A(n33514), .B(n33515), .Z(n30682) );
  NOR U30786 ( .A(n33516), .B(n33514), .Z(n33515) );
  XOR U30787 ( .A(n33517), .B(n33518), .Z(n30685) );
  NOR U30788 ( .A(n33519), .B(n33517), .Z(n33518) );
  XOR U30789 ( .A(n33520), .B(n33521), .Z(n30688) );
  NOR U30790 ( .A(n33522), .B(n33520), .Z(n33521) );
  XOR U30791 ( .A(n33523), .B(n33524), .Z(n30691) );
  NOR U30792 ( .A(n33525), .B(n33523), .Z(n33524) );
  XOR U30793 ( .A(n33526), .B(n33527), .Z(n30694) );
  NOR U30794 ( .A(n33528), .B(n33526), .Z(n33527) );
  XOR U30795 ( .A(n33529), .B(n33530), .Z(n30697) );
  NOR U30796 ( .A(n33531), .B(n33529), .Z(n33530) );
  XOR U30797 ( .A(n33532), .B(n33533), .Z(n30700) );
  NOR U30798 ( .A(n33534), .B(n33532), .Z(n33533) );
  XOR U30799 ( .A(n33535), .B(n33536), .Z(n30703) );
  NOR U30800 ( .A(n33537), .B(n33535), .Z(n33536) );
  XOR U30801 ( .A(n33538), .B(n33539), .Z(n30706) );
  NOR U30802 ( .A(n33540), .B(n33538), .Z(n33539) );
  XOR U30803 ( .A(n33541), .B(n33542), .Z(n30709) );
  NOR U30804 ( .A(n33543), .B(n33541), .Z(n33542) );
  XOR U30805 ( .A(n33544), .B(n33545), .Z(n30712) );
  NOR U30806 ( .A(n33546), .B(n33544), .Z(n33545) );
  XOR U30807 ( .A(n33547), .B(n33548), .Z(n30715) );
  NOR U30808 ( .A(n33549), .B(n33547), .Z(n33548) );
  XOR U30809 ( .A(n33550), .B(n33551), .Z(n30718) );
  NOR U30810 ( .A(n33552), .B(n33550), .Z(n33551) );
  XOR U30811 ( .A(n33553), .B(n33554), .Z(n30721) );
  NOR U30812 ( .A(n33555), .B(n33553), .Z(n33554) );
  XOR U30813 ( .A(n33556), .B(n33557), .Z(n30724) );
  NOR U30814 ( .A(n33558), .B(n33556), .Z(n33557) );
  XOR U30815 ( .A(n33559), .B(n33560), .Z(n30727) );
  NOR U30816 ( .A(n33561), .B(n33559), .Z(n33560) );
  XOR U30817 ( .A(n33562), .B(n33563), .Z(n30730) );
  NOR U30818 ( .A(n33564), .B(n33562), .Z(n33563) );
  XOR U30819 ( .A(n33565), .B(n33566), .Z(n30733) );
  NOR U30820 ( .A(n33567), .B(n33565), .Z(n33566) );
  XOR U30821 ( .A(n33568), .B(n33569), .Z(n30736) );
  NOR U30822 ( .A(n33570), .B(n33568), .Z(n33569) );
  XOR U30823 ( .A(n33571), .B(n33572), .Z(n30739) );
  NOR U30824 ( .A(n33573), .B(n33571), .Z(n33572) );
  XOR U30825 ( .A(n33574), .B(n33575), .Z(n30742) );
  NOR U30826 ( .A(n33576), .B(n33574), .Z(n33575) );
  XOR U30827 ( .A(n33577), .B(n33578), .Z(n30745) );
  NOR U30828 ( .A(n33579), .B(n33577), .Z(n33578) );
  XOR U30829 ( .A(n33580), .B(n33581), .Z(n30748) );
  NOR U30830 ( .A(n33582), .B(n33580), .Z(n33581) );
  XOR U30831 ( .A(n33583), .B(n33584), .Z(n30751) );
  NOR U30832 ( .A(n33585), .B(n33583), .Z(n33584) );
  XOR U30833 ( .A(n33586), .B(n33587), .Z(n30754) );
  NOR U30834 ( .A(n33588), .B(n33586), .Z(n33587) );
  XOR U30835 ( .A(n33589), .B(n33590), .Z(n30757) );
  NOR U30836 ( .A(n33591), .B(n33589), .Z(n33590) );
  XOR U30837 ( .A(n33592), .B(n33593), .Z(n30760) );
  NOR U30838 ( .A(n33594), .B(n33592), .Z(n33593) );
  XOR U30839 ( .A(n33595), .B(n33596), .Z(n30763) );
  NOR U30840 ( .A(n33597), .B(n33595), .Z(n33596) );
  XOR U30841 ( .A(n33598), .B(n33599), .Z(n30766) );
  NOR U30842 ( .A(n33600), .B(n33598), .Z(n33599) );
  XOR U30843 ( .A(n33601), .B(n33602), .Z(n30769) );
  NOR U30844 ( .A(n33603), .B(n33601), .Z(n33602) );
  XOR U30845 ( .A(n33604), .B(n33605), .Z(n30772) );
  NOR U30846 ( .A(n33606), .B(n33604), .Z(n33605) );
  XOR U30847 ( .A(n33607), .B(n33608), .Z(n30775) );
  NOR U30848 ( .A(n33609), .B(n33607), .Z(n33608) );
  XOR U30849 ( .A(n33610), .B(n33611), .Z(n30778) );
  NOR U30850 ( .A(n33612), .B(n33610), .Z(n33611) );
  XOR U30851 ( .A(n33613), .B(n33614), .Z(n30781) );
  NOR U30852 ( .A(n33615), .B(n33613), .Z(n33614) );
  XOR U30853 ( .A(n33616), .B(n33617), .Z(n30784) );
  NOR U30854 ( .A(n33618), .B(n33616), .Z(n33617) );
  XOR U30855 ( .A(n33619), .B(n33620), .Z(n30787) );
  NOR U30856 ( .A(n33621), .B(n33619), .Z(n33620) );
  XOR U30857 ( .A(n33622), .B(n33623), .Z(n30790) );
  NOR U30858 ( .A(n33624), .B(n33622), .Z(n33623) );
  XOR U30859 ( .A(n33625), .B(n33626), .Z(n30793) );
  NOR U30860 ( .A(n33627), .B(n33625), .Z(n33626) );
  XOR U30861 ( .A(n33628), .B(n33629), .Z(n30796) );
  NOR U30862 ( .A(n33630), .B(n33628), .Z(n33629) );
  XOR U30863 ( .A(n33631), .B(n33632), .Z(n30799) );
  NOR U30864 ( .A(n33633), .B(n33631), .Z(n33632) );
  XOR U30865 ( .A(n33634), .B(n33635), .Z(n30802) );
  NOR U30866 ( .A(n33636), .B(n33634), .Z(n33635) );
  XOR U30867 ( .A(n33637), .B(n33638), .Z(n30805) );
  NOR U30868 ( .A(n33639), .B(n33637), .Z(n33638) );
  XOR U30869 ( .A(n33640), .B(n33641), .Z(n30808) );
  NOR U30870 ( .A(n33642), .B(n33640), .Z(n33641) );
  XOR U30871 ( .A(n33643), .B(n33644), .Z(n30811) );
  NOR U30872 ( .A(n33645), .B(n33643), .Z(n33644) );
  XOR U30873 ( .A(n33646), .B(n33647), .Z(n30814) );
  NOR U30874 ( .A(n33648), .B(n33646), .Z(n33647) );
  XOR U30875 ( .A(n33649), .B(n33650), .Z(n30817) );
  NOR U30876 ( .A(n33651), .B(n33649), .Z(n33650) );
  XOR U30877 ( .A(n33652), .B(n33653), .Z(n30820) );
  NOR U30878 ( .A(n33654), .B(n33652), .Z(n33653) );
  XOR U30879 ( .A(n33655), .B(n33656), .Z(n30823) );
  NOR U30880 ( .A(n33657), .B(n33655), .Z(n33656) );
  XOR U30881 ( .A(n33658), .B(n33659), .Z(n30826) );
  NOR U30882 ( .A(n33660), .B(n33658), .Z(n33659) );
  XOR U30883 ( .A(n33661), .B(n33662), .Z(n30829) );
  NOR U30884 ( .A(n33663), .B(n33661), .Z(n33662) );
  XOR U30885 ( .A(n33664), .B(n33665), .Z(n30832) );
  NOR U30886 ( .A(n33666), .B(n33664), .Z(n33665) );
  XOR U30887 ( .A(n33667), .B(n33668), .Z(n30835) );
  NOR U30888 ( .A(n33669), .B(n33667), .Z(n33668) );
  XOR U30889 ( .A(n33670), .B(n33671), .Z(n30838) );
  NOR U30890 ( .A(n33672), .B(n33670), .Z(n33671) );
  XOR U30891 ( .A(n33673), .B(n33674), .Z(n30841) );
  NOR U30892 ( .A(n33675), .B(n33673), .Z(n33674) );
  XOR U30893 ( .A(n33676), .B(n33677), .Z(n30844) );
  NOR U30894 ( .A(n33678), .B(n33676), .Z(n33677) );
  XOR U30895 ( .A(n33679), .B(n33680), .Z(n30847) );
  NOR U30896 ( .A(n33681), .B(n33679), .Z(n33680) );
  XOR U30897 ( .A(n33682), .B(n33683), .Z(n30850) );
  NOR U30898 ( .A(n33684), .B(n33682), .Z(n33683) );
  XOR U30899 ( .A(n33685), .B(n33686), .Z(n30853) );
  NOR U30900 ( .A(n33687), .B(n33685), .Z(n33686) );
  XOR U30901 ( .A(n33688), .B(n33689), .Z(n30856) );
  NOR U30902 ( .A(n33690), .B(n33688), .Z(n33689) );
  XOR U30903 ( .A(n33691), .B(n33692), .Z(n30859) );
  NOR U30904 ( .A(n33693), .B(n33691), .Z(n33692) );
  XOR U30905 ( .A(n33694), .B(n33695), .Z(n30862) );
  NOR U30906 ( .A(n33696), .B(n33694), .Z(n33695) );
  XOR U30907 ( .A(n33697), .B(n33698), .Z(n30865) );
  NOR U30908 ( .A(n33699), .B(n33697), .Z(n33698) );
  XOR U30909 ( .A(n33700), .B(n33701), .Z(n30868) );
  NOR U30910 ( .A(n33702), .B(n33700), .Z(n33701) );
  XOR U30911 ( .A(n33703), .B(n33704), .Z(n30871) );
  NOR U30912 ( .A(n33705), .B(n33703), .Z(n33704) );
  XOR U30913 ( .A(n33706), .B(n33707), .Z(n30874) );
  NOR U30914 ( .A(n33708), .B(n33706), .Z(n33707) );
  XOR U30915 ( .A(n33709), .B(n33710), .Z(n30877) );
  NOR U30916 ( .A(n33711), .B(n33709), .Z(n33710) );
  XOR U30917 ( .A(n33712), .B(n33713), .Z(n30880) );
  NOR U30918 ( .A(n33714), .B(n33712), .Z(n33713) );
  XOR U30919 ( .A(n33715), .B(n33716), .Z(n30883) );
  NOR U30920 ( .A(n33717), .B(n33715), .Z(n33716) );
  XOR U30921 ( .A(n33718), .B(n33719), .Z(n30886) );
  NOR U30922 ( .A(n33720), .B(n33718), .Z(n33719) );
  XOR U30923 ( .A(n33721), .B(n33722), .Z(n30889) );
  NOR U30924 ( .A(n33723), .B(n33721), .Z(n33722) );
  XOR U30925 ( .A(n33724), .B(n33725), .Z(n30892) );
  NOR U30926 ( .A(n33726), .B(n33724), .Z(n33725) );
  XOR U30927 ( .A(n33727), .B(n33728), .Z(n30895) );
  NOR U30928 ( .A(n33729), .B(n33727), .Z(n33728) );
  XOR U30929 ( .A(n33730), .B(n33731), .Z(n30898) );
  NOR U30930 ( .A(n33732), .B(n33730), .Z(n33731) );
  XOR U30931 ( .A(n33733), .B(n33734), .Z(n30901) );
  NOR U30932 ( .A(n33735), .B(n33733), .Z(n33734) );
  XOR U30933 ( .A(n33736), .B(n33737), .Z(n30904) );
  NOR U30934 ( .A(n33738), .B(n33736), .Z(n33737) );
  XOR U30935 ( .A(n33739), .B(n33740), .Z(n30907) );
  NOR U30936 ( .A(n33741), .B(n33739), .Z(n33740) );
  XOR U30937 ( .A(n33742), .B(n33743), .Z(n30910) );
  NOR U30938 ( .A(n33744), .B(n33742), .Z(n33743) );
  XOR U30939 ( .A(n33745), .B(n33746), .Z(n30913) );
  NOR U30940 ( .A(n33747), .B(n33745), .Z(n33746) );
  XOR U30941 ( .A(n33748), .B(n33749), .Z(n30916) );
  NOR U30942 ( .A(n33750), .B(n33748), .Z(n33749) );
  XOR U30943 ( .A(n33751), .B(n33752), .Z(n30919) );
  NOR U30944 ( .A(n33753), .B(n33751), .Z(n33752) );
  XOR U30945 ( .A(n33754), .B(n33755), .Z(n30922) );
  NOR U30946 ( .A(n33756), .B(n33754), .Z(n33755) );
  XOR U30947 ( .A(n33757), .B(n33758), .Z(n30925) );
  NOR U30948 ( .A(n33759), .B(n33757), .Z(n33758) );
  XOR U30949 ( .A(n33760), .B(n33761), .Z(n30928) );
  NOR U30950 ( .A(n33762), .B(n33760), .Z(n33761) );
  XOR U30951 ( .A(n33763), .B(n33764), .Z(n30931) );
  NOR U30952 ( .A(n33765), .B(n33763), .Z(n33764) );
  XOR U30953 ( .A(n33766), .B(n33767), .Z(n30934) );
  NOR U30954 ( .A(n33768), .B(n33766), .Z(n33767) );
  XOR U30955 ( .A(n33769), .B(n33770), .Z(n30937) );
  NOR U30956 ( .A(n33771), .B(n33769), .Z(n33770) );
  XOR U30957 ( .A(n33772), .B(n33773), .Z(n30940) );
  NOR U30958 ( .A(n33774), .B(n33772), .Z(n33773) );
  XOR U30959 ( .A(n33775), .B(n33776), .Z(n30943) );
  NOR U30960 ( .A(n33777), .B(n33775), .Z(n33776) );
  XOR U30961 ( .A(n33778), .B(n33779), .Z(n30946) );
  NOR U30962 ( .A(n33780), .B(n33778), .Z(n33779) );
  XOR U30963 ( .A(n33781), .B(n33782), .Z(n30949) );
  NOR U30964 ( .A(n33783), .B(n33781), .Z(n33782) );
  XOR U30965 ( .A(n33784), .B(n33785), .Z(n30952) );
  NOR U30966 ( .A(n33786), .B(n33784), .Z(n33785) );
  XOR U30967 ( .A(n33787), .B(n33788), .Z(n30955) );
  NOR U30968 ( .A(n33789), .B(n33787), .Z(n33788) );
  XOR U30969 ( .A(n33790), .B(n33791), .Z(n30958) );
  NOR U30970 ( .A(n33792), .B(n33790), .Z(n33791) );
  XOR U30971 ( .A(n33793), .B(n33794), .Z(n30961) );
  NOR U30972 ( .A(n33795), .B(n33793), .Z(n33794) );
  XOR U30973 ( .A(n33796), .B(n33797), .Z(n30964) );
  NOR U30974 ( .A(n33798), .B(n33796), .Z(n33797) );
  XOR U30975 ( .A(n33799), .B(n33800), .Z(n30967) );
  NOR U30976 ( .A(n33801), .B(n33799), .Z(n33800) );
  XOR U30977 ( .A(n33802), .B(n33803), .Z(n30970) );
  NOR U30978 ( .A(n33804), .B(n33802), .Z(n33803) );
  XOR U30979 ( .A(n33805), .B(n33806), .Z(n30973) );
  NOR U30980 ( .A(n33807), .B(n33805), .Z(n33806) );
  XOR U30981 ( .A(n33808), .B(n33809), .Z(n30976) );
  NOR U30982 ( .A(n33810), .B(n33808), .Z(n33809) );
  XOR U30983 ( .A(n33811), .B(n33812), .Z(n30979) );
  NOR U30984 ( .A(n33813), .B(n33811), .Z(n33812) );
  XOR U30985 ( .A(n33814), .B(n33815), .Z(n30982) );
  NOR U30986 ( .A(n33816), .B(n33814), .Z(n33815) );
  XOR U30987 ( .A(n33817), .B(n33818), .Z(n30985) );
  NOR U30988 ( .A(n33819), .B(n33817), .Z(n33818) );
  XOR U30989 ( .A(n33820), .B(n33821), .Z(n30988) );
  NOR U30990 ( .A(n33822), .B(n33820), .Z(n33821) );
  XOR U30991 ( .A(n33823), .B(n33824), .Z(n30991) );
  NOR U30992 ( .A(n33825), .B(n33823), .Z(n33824) );
  XOR U30993 ( .A(n33826), .B(n33827), .Z(n30994) );
  NOR U30994 ( .A(n33828), .B(n33826), .Z(n33827) );
  XOR U30995 ( .A(n33829), .B(n33830), .Z(n30997) );
  NOR U30996 ( .A(n33831), .B(n33829), .Z(n33830) );
  XOR U30997 ( .A(n33832), .B(n33833), .Z(n31000) );
  NOR U30998 ( .A(n33834), .B(n33832), .Z(n33833) );
  XOR U30999 ( .A(n33835), .B(n33836), .Z(n31003) );
  NOR U31000 ( .A(n33837), .B(n33835), .Z(n33836) );
  XOR U31001 ( .A(n33838), .B(n33839), .Z(n31006) );
  NOR U31002 ( .A(n33840), .B(n33838), .Z(n33839) );
  XOR U31003 ( .A(n33841), .B(n33842), .Z(n31009) );
  NOR U31004 ( .A(n33843), .B(n33841), .Z(n33842) );
  XOR U31005 ( .A(n33844), .B(n33845), .Z(n31012) );
  NOR U31006 ( .A(n33846), .B(n33844), .Z(n33845) );
  XOR U31007 ( .A(n33847), .B(n33848), .Z(n31015) );
  NOR U31008 ( .A(n33849), .B(n33847), .Z(n33848) );
  XOR U31009 ( .A(n33850), .B(n33851), .Z(n31018) );
  NOR U31010 ( .A(n33852), .B(n33850), .Z(n33851) );
  XOR U31011 ( .A(n33853), .B(n33854), .Z(n31021) );
  NOR U31012 ( .A(n33855), .B(n33853), .Z(n33854) );
  XOR U31013 ( .A(n33856), .B(n33857), .Z(n31024) );
  NOR U31014 ( .A(n33858), .B(n33856), .Z(n33857) );
  XOR U31015 ( .A(n33859), .B(n33860), .Z(n31027) );
  NOR U31016 ( .A(n33861), .B(n33859), .Z(n33860) );
  XOR U31017 ( .A(n33862), .B(n33863), .Z(n31030) );
  NOR U31018 ( .A(n33864), .B(n33862), .Z(n33863) );
  XOR U31019 ( .A(n33865), .B(n33866), .Z(n31033) );
  NOR U31020 ( .A(n33867), .B(n33865), .Z(n33866) );
  XOR U31021 ( .A(n33868), .B(n33869), .Z(n31036) );
  NOR U31022 ( .A(n33870), .B(n33868), .Z(n33869) );
  XOR U31023 ( .A(n33871), .B(n33872), .Z(n31039) );
  NOR U31024 ( .A(n33873), .B(n33871), .Z(n33872) );
  XOR U31025 ( .A(n33874), .B(n33875), .Z(n31042) );
  NOR U31026 ( .A(n33876), .B(n33874), .Z(n33875) );
  XOR U31027 ( .A(n33877), .B(n33878), .Z(n31045) );
  NOR U31028 ( .A(n33879), .B(n33877), .Z(n33878) );
  XOR U31029 ( .A(n33880), .B(n33881), .Z(n31048) );
  NOR U31030 ( .A(n33882), .B(n33880), .Z(n33881) );
  XOR U31031 ( .A(n33883), .B(n33884), .Z(n31051) );
  NOR U31032 ( .A(n33885), .B(n33883), .Z(n33884) );
  XOR U31033 ( .A(n33886), .B(n33887), .Z(n31054) );
  NOR U31034 ( .A(n33888), .B(n33886), .Z(n33887) );
  XOR U31035 ( .A(n33889), .B(n33890), .Z(n31057) );
  NOR U31036 ( .A(n33891), .B(n33889), .Z(n33890) );
  XOR U31037 ( .A(n33892), .B(n33893), .Z(n31060) );
  NOR U31038 ( .A(n33894), .B(n33892), .Z(n33893) );
  XOR U31039 ( .A(n33895), .B(n33896), .Z(n31063) );
  NOR U31040 ( .A(n33897), .B(n33895), .Z(n33896) );
  XOR U31041 ( .A(n33898), .B(n33899), .Z(n31066) );
  NOR U31042 ( .A(n33900), .B(n33898), .Z(n33899) );
  XOR U31043 ( .A(n33901), .B(n33902), .Z(n31069) );
  NOR U31044 ( .A(n33903), .B(n33901), .Z(n33902) );
  XOR U31045 ( .A(n33904), .B(n33905), .Z(n31072) );
  NOR U31046 ( .A(n33906), .B(n33904), .Z(n33905) );
  XOR U31047 ( .A(n33907), .B(n33908), .Z(n31075) );
  NOR U31048 ( .A(n33909), .B(n33907), .Z(n33908) );
  XOR U31049 ( .A(n33910), .B(n33911), .Z(n31078) );
  NOR U31050 ( .A(n33912), .B(n33910), .Z(n33911) );
  XOR U31051 ( .A(n33913), .B(n33914), .Z(n31081) );
  NOR U31052 ( .A(n33915), .B(n33913), .Z(n33914) );
  XOR U31053 ( .A(n33916), .B(n33917), .Z(n31084) );
  NOR U31054 ( .A(n33918), .B(n33916), .Z(n33917) );
  XOR U31055 ( .A(n33919), .B(n33920), .Z(n31087) );
  NOR U31056 ( .A(n33921), .B(n33919), .Z(n33920) );
  XOR U31057 ( .A(n33922), .B(n33923), .Z(n31090) );
  NOR U31058 ( .A(n33924), .B(n33922), .Z(n33923) );
  XOR U31059 ( .A(n33925), .B(n33926), .Z(n31093) );
  NOR U31060 ( .A(n33927), .B(n33925), .Z(n33926) );
  XOR U31061 ( .A(n33928), .B(n33929), .Z(n31096) );
  NOR U31062 ( .A(n33930), .B(n33928), .Z(n33929) );
  XOR U31063 ( .A(n33931), .B(n33932), .Z(n31099) );
  NOR U31064 ( .A(n33933), .B(n33931), .Z(n33932) );
  XOR U31065 ( .A(n33934), .B(n33935), .Z(n31102) );
  NOR U31066 ( .A(n33936), .B(n33934), .Z(n33935) );
  XOR U31067 ( .A(n33937), .B(n33938), .Z(n31105) );
  NOR U31068 ( .A(n33939), .B(n33937), .Z(n33938) );
  XOR U31069 ( .A(n33940), .B(n33941), .Z(n31108) );
  NOR U31070 ( .A(n33942), .B(n33940), .Z(n33941) );
  XOR U31071 ( .A(n33943), .B(n33944), .Z(n31111) );
  NOR U31072 ( .A(n33945), .B(n33943), .Z(n33944) );
  XOR U31073 ( .A(n33946), .B(n33947), .Z(n31114) );
  NOR U31074 ( .A(n33948), .B(n33946), .Z(n33947) );
  XOR U31075 ( .A(n33949), .B(n33950), .Z(n31117) );
  NOR U31076 ( .A(n33951), .B(n33949), .Z(n33950) );
  XOR U31077 ( .A(n33952), .B(n33953), .Z(n31120) );
  NOR U31078 ( .A(n33954), .B(n33952), .Z(n33953) );
  XOR U31079 ( .A(n33955), .B(n33956), .Z(n31123) );
  NOR U31080 ( .A(n33957), .B(n33955), .Z(n33956) );
  XOR U31081 ( .A(n33958), .B(n33959), .Z(n31126) );
  NOR U31082 ( .A(n33960), .B(n33958), .Z(n33959) );
  XOR U31083 ( .A(n33961), .B(n33962), .Z(n31129) );
  NOR U31084 ( .A(n33963), .B(n33961), .Z(n33962) );
  XOR U31085 ( .A(n33964), .B(n33965), .Z(n31132) );
  NOR U31086 ( .A(n33966), .B(n33964), .Z(n33965) );
  XOR U31087 ( .A(n33967), .B(n33968), .Z(n31135) );
  NOR U31088 ( .A(n33969), .B(n33967), .Z(n33968) );
  XOR U31089 ( .A(n33970), .B(n33971), .Z(n31138) );
  NOR U31090 ( .A(n33972), .B(n33970), .Z(n33971) );
  XOR U31091 ( .A(n33973), .B(n33974), .Z(n31141) );
  NOR U31092 ( .A(n33975), .B(n33973), .Z(n33974) );
  XOR U31093 ( .A(n33976), .B(n33977), .Z(n31144) );
  NOR U31094 ( .A(n33978), .B(n33976), .Z(n33977) );
  XOR U31095 ( .A(n33979), .B(n33980), .Z(n31147) );
  NOR U31096 ( .A(n33981), .B(n33979), .Z(n33980) );
  XOR U31097 ( .A(n33982), .B(n33983), .Z(n31150) );
  NOR U31098 ( .A(n33984), .B(n33982), .Z(n33983) );
  XOR U31099 ( .A(n33985), .B(n33986), .Z(n31153) );
  NOR U31100 ( .A(n33987), .B(n33985), .Z(n33986) );
  XOR U31101 ( .A(n33988), .B(n33989), .Z(n31156) );
  NOR U31102 ( .A(n33990), .B(n33988), .Z(n33989) );
  XOR U31103 ( .A(n33991), .B(n33992), .Z(n31159) );
  NOR U31104 ( .A(n33993), .B(n33991), .Z(n33992) );
  XOR U31105 ( .A(n33994), .B(n33995), .Z(n31162) );
  NOR U31106 ( .A(n33996), .B(n33994), .Z(n33995) );
  XOR U31107 ( .A(n33997), .B(n33998), .Z(n31165) );
  NOR U31108 ( .A(n33999), .B(n33997), .Z(n33998) );
  XOR U31109 ( .A(n34000), .B(n34001), .Z(n31168) );
  NOR U31110 ( .A(n34002), .B(n34000), .Z(n34001) );
  XOR U31111 ( .A(n34003), .B(n34004), .Z(n31171) );
  NOR U31112 ( .A(n34005), .B(n34003), .Z(n34004) );
  XOR U31113 ( .A(n34006), .B(n34007), .Z(n31174) );
  NOR U31114 ( .A(n34008), .B(n34006), .Z(n34007) );
  XOR U31115 ( .A(n34009), .B(n34010), .Z(n31177) );
  NOR U31116 ( .A(n34011), .B(n34009), .Z(n34010) );
  XOR U31117 ( .A(n34012), .B(n34013), .Z(n31180) );
  NOR U31118 ( .A(n34014), .B(n34012), .Z(n34013) );
  XOR U31119 ( .A(n34015), .B(n34016), .Z(n31183) );
  NOR U31120 ( .A(n34017), .B(n34015), .Z(n34016) );
  XOR U31121 ( .A(n34018), .B(n34019), .Z(n31186) );
  NOR U31122 ( .A(n34020), .B(n34018), .Z(n34019) );
  XOR U31123 ( .A(n34021), .B(n34022), .Z(n31189) );
  NOR U31124 ( .A(n34023), .B(n34021), .Z(n34022) );
  XOR U31125 ( .A(n34024), .B(n34025), .Z(n31192) );
  NOR U31126 ( .A(n34026), .B(n34024), .Z(n34025) );
  XOR U31127 ( .A(n34027), .B(n34028), .Z(n31195) );
  NOR U31128 ( .A(n34029), .B(n34027), .Z(n34028) );
  XOR U31129 ( .A(n34030), .B(n34031), .Z(n31198) );
  NOR U31130 ( .A(n34032), .B(n34030), .Z(n34031) );
  XOR U31131 ( .A(n34033), .B(n34034), .Z(n31201) );
  NOR U31132 ( .A(n34035), .B(n34033), .Z(n34034) );
  XOR U31133 ( .A(n34036), .B(n34037), .Z(n31204) );
  NOR U31134 ( .A(n34038), .B(n34036), .Z(n34037) );
  XOR U31135 ( .A(n34039), .B(n34040), .Z(n31207) );
  NOR U31136 ( .A(n34041), .B(n34039), .Z(n34040) );
  XOR U31137 ( .A(n34042), .B(n34043), .Z(n31210) );
  NOR U31138 ( .A(n34044), .B(n34042), .Z(n34043) );
  XOR U31139 ( .A(n34045), .B(n34046), .Z(n31213) );
  NOR U31140 ( .A(n34047), .B(n34045), .Z(n34046) );
  XOR U31141 ( .A(n34048), .B(n34049), .Z(n31216) );
  NOR U31142 ( .A(n34050), .B(n34048), .Z(n34049) );
  XOR U31143 ( .A(n34051), .B(n34052), .Z(n31219) );
  NOR U31144 ( .A(n34053), .B(n34051), .Z(n34052) );
  XOR U31145 ( .A(n34054), .B(n34055), .Z(n31222) );
  NOR U31146 ( .A(n34056), .B(n34054), .Z(n34055) );
  XOR U31147 ( .A(n34057), .B(n34058), .Z(n31225) );
  NOR U31148 ( .A(n34059), .B(n34057), .Z(n34058) );
  XOR U31149 ( .A(n34060), .B(n34061), .Z(n31228) );
  NOR U31150 ( .A(n34062), .B(n34060), .Z(n34061) );
  XOR U31151 ( .A(n34063), .B(n34064), .Z(n31231) );
  NOR U31152 ( .A(n34065), .B(n34063), .Z(n34064) );
  XOR U31153 ( .A(n34066), .B(n34067), .Z(n31234) );
  NOR U31154 ( .A(n34068), .B(n34066), .Z(n34067) );
  XOR U31155 ( .A(n34069), .B(n34070), .Z(n31237) );
  NOR U31156 ( .A(n34071), .B(n34069), .Z(n34070) );
  XOR U31157 ( .A(n34072), .B(n34073), .Z(n31240) );
  NOR U31158 ( .A(n34074), .B(n34072), .Z(n34073) );
  XOR U31159 ( .A(n34075), .B(n34076), .Z(n31243) );
  NOR U31160 ( .A(n34077), .B(n34075), .Z(n34076) );
  XOR U31161 ( .A(n34078), .B(n34079), .Z(n31246) );
  NOR U31162 ( .A(n34080), .B(n34078), .Z(n34079) );
  XOR U31163 ( .A(n34081), .B(n34082), .Z(n31249) );
  NOR U31164 ( .A(n34083), .B(n34081), .Z(n34082) );
  XOR U31165 ( .A(n34084), .B(n34085), .Z(n31252) );
  NOR U31166 ( .A(n34086), .B(n34084), .Z(n34085) );
  XOR U31167 ( .A(n34087), .B(n34088), .Z(n31255) );
  NOR U31168 ( .A(n34089), .B(n34087), .Z(n34088) );
  XOR U31169 ( .A(n34090), .B(n34091), .Z(n31258) );
  NOR U31170 ( .A(n34092), .B(n34090), .Z(n34091) );
  XOR U31171 ( .A(n34093), .B(n34094), .Z(n31261) );
  NOR U31172 ( .A(n34095), .B(n34093), .Z(n34094) );
  XOR U31173 ( .A(n34096), .B(n34097), .Z(n31264) );
  NOR U31174 ( .A(n34098), .B(n34096), .Z(n34097) );
  XOR U31175 ( .A(n34099), .B(n34100), .Z(n31267) );
  NOR U31176 ( .A(n91), .B(n34101), .Z(n34100) );
  IV U31177 ( .A(n34099), .Z(n34101) );
  XOR U31178 ( .A(n34102), .B(n34103), .Z(n31270) );
  AND U31179 ( .A(n34104), .B(n34105), .Z(n34103) );
  XOR U31180 ( .A(n34102), .B(n94), .Z(n34105) );
  XOR U31181 ( .A(n32686), .B(n32685), .Z(n94) );
  XNOR U31182 ( .A(n32683), .B(n32682), .Z(n32685) );
  XNOR U31183 ( .A(n32680), .B(n32679), .Z(n32682) );
  XNOR U31184 ( .A(n32677), .B(n32676), .Z(n32679) );
  XNOR U31185 ( .A(n32674), .B(n32673), .Z(n32676) );
  XNOR U31186 ( .A(n32671), .B(n32670), .Z(n32673) );
  XNOR U31187 ( .A(n32668), .B(n32667), .Z(n32670) );
  XNOR U31188 ( .A(n32665), .B(n32664), .Z(n32667) );
  XNOR U31189 ( .A(n32662), .B(n32661), .Z(n32664) );
  XNOR U31190 ( .A(n32659), .B(n32658), .Z(n32661) );
  XNOR U31191 ( .A(n32656), .B(n32655), .Z(n32658) );
  XNOR U31192 ( .A(n32653), .B(n32652), .Z(n32655) );
  XNOR U31193 ( .A(n32650), .B(n32649), .Z(n32652) );
  XNOR U31194 ( .A(n32647), .B(n32646), .Z(n32649) );
  XNOR U31195 ( .A(n32644), .B(n32643), .Z(n32646) );
  XNOR U31196 ( .A(n32641), .B(n32640), .Z(n32643) );
  XNOR U31197 ( .A(n32638), .B(n32637), .Z(n32640) );
  XNOR U31198 ( .A(n32635), .B(n32634), .Z(n32637) );
  XNOR U31199 ( .A(n32632), .B(n32631), .Z(n32634) );
  XNOR U31200 ( .A(n32629), .B(n32628), .Z(n32631) );
  XNOR U31201 ( .A(n32626), .B(n32625), .Z(n32628) );
  XNOR U31202 ( .A(n32623), .B(n32622), .Z(n32625) );
  XNOR U31203 ( .A(n32620), .B(n32619), .Z(n32622) );
  XNOR U31204 ( .A(n32617), .B(n32616), .Z(n32619) );
  XNOR U31205 ( .A(n32614), .B(n32613), .Z(n32616) );
  XNOR U31206 ( .A(n32611), .B(n32610), .Z(n32613) );
  XNOR U31207 ( .A(n32608), .B(n32607), .Z(n32610) );
  XNOR U31208 ( .A(n32605), .B(n32604), .Z(n32607) );
  XNOR U31209 ( .A(n32602), .B(n32601), .Z(n32604) );
  XNOR U31210 ( .A(n32599), .B(n32598), .Z(n32601) );
  XNOR U31211 ( .A(n32596), .B(n32595), .Z(n32598) );
  XNOR U31212 ( .A(n32593), .B(n32592), .Z(n32595) );
  XNOR U31213 ( .A(n32590), .B(n32589), .Z(n32592) );
  XNOR U31214 ( .A(n32587), .B(n32586), .Z(n32589) );
  XNOR U31215 ( .A(n32584), .B(n32583), .Z(n32586) );
  XNOR U31216 ( .A(n32581), .B(n32580), .Z(n32583) );
  XNOR U31217 ( .A(n32578), .B(n32577), .Z(n32580) );
  XNOR U31218 ( .A(n32575), .B(n32574), .Z(n32577) );
  XNOR U31219 ( .A(n32572), .B(n32571), .Z(n32574) );
  XNOR U31220 ( .A(n32569), .B(n32568), .Z(n32571) );
  XNOR U31221 ( .A(n32566), .B(n32565), .Z(n32568) );
  XNOR U31222 ( .A(n32563), .B(n32562), .Z(n32565) );
  XNOR U31223 ( .A(n32560), .B(n32559), .Z(n32562) );
  XNOR U31224 ( .A(n32557), .B(n32556), .Z(n32559) );
  XNOR U31225 ( .A(n32554), .B(n32553), .Z(n32556) );
  XNOR U31226 ( .A(n32551), .B(n32550), .Z(n32553) );
  XNOR U31227 ( .A(n32548), .B(n32547), .Z(n32550) );
  XNOR U31228 ( .A(n32545), .B(n32544), .Z(n32547) );
  XNOR U31229 ( .A(n32542), .B(n32541), .Z(n32544) );
  XNOR U31230 ( .A(n32539), .B(n32538), .Z(n32541) );
  XNOR U31231 ( .A(n32536), .B(n32535), .Z(n32538) );
  XNOR U31232 ( .A(n32533), .B(n32532), .Z(n32535) );
  XNOR U31233 ( .A(n32530), .B(n32529), .Z(n32532) );
  XNOR U31234 ( .A(n32527), .B(n32526), .Z(n32529) );
  XNOR U31235 ( .A(n32524), .B(n32523), .Z(n32526) );
  XNOR U31236 ( .A(n32521), .B(n32520), .Z(n32523) );
  XNOR U31237 ( .A(n32518), .B(n32517), .Z(n32520) );
  XNOR U31238 ( .A(n32515), .B(n32514), .Z(n32517) );
  XNOR U31239 ( .A(n32512), .B(n32511), .Z(n32514) );
  XNOR U31240 ( .A(n32509), .B(n32508), .Z(n32511) );
  XNOR U31241 ( .A(n32506), .B(n32505), .Z(n32508) );
  XNOR U31242 ( .A(n32503), .B(n32502), .Z(n32505) );
  XNOR U31243 ( .A(n32500), .B(n32499), .Z(n32502) );
  XNOR U31244 ( .A(n32497), .B(n32496), .Z(n32499) );
  XNOR U31245 ( .A(n32494), .B(n32493), .Z(n32496) );
  XNOR U31246 ( .A(n32491), .B(n32490), .Z(n32493) );
  XNOR U31247 ( .A(n32488), .B(n32487), .Z(n32490) );
  XNOR U31248 ( .A(n32485), .B(n32484), .Z(n32487) );
  XNOR U31249 ( .A(n32482), .B(n32481), .Z(n32484) );
  XNOR U31250 ( .A(n32479), .B(n32478), .Z(n32481) );
  XNOR U31251 ( .A(n32476), .B(n32475), .Z(n32478) );
  XNOR U31252 ( .A(n32473), .B(n32472), .Z(n32475) );
  XNOR U31253 ( .A(n32470), .B(n32469), .Z(n32472) );
  XNOR U31254 ( .A(n32467), .B(n32466), .Z(n32469) );
  XNOR U31255 ( .A(n32464), .B(n32463), .Z(n32466) );
  XNOR U31256 ( .A(n32461), .B(n32460), .Z(n32463) );
  XNOR U31257 ( .A(n32458), .B(n32457), .Z(n32460) );
  XNOR U31258 ( .A(n32455), .B(n32454), .Z(n32457) );
  XNOR U31259 ( .A(n32452), .B(n32451), .Z(n32454) );
  XNOR U31260 ( .A(n32449), .B(n32448), .Z(n32451) );
  XNOR U31261 ( .A(n32446), .B(n32445), .Z(n32448) );
  XNOR U31262 ( .A(n32443), .B(n32442), .Z(n32445) );
  XNOR U31263 ( .A(n32440), .B(n32439), .Z(n32442) );
  XNOR U31264 ( .A(n32437), .B(n32436), .Z(n32439) );
  XNOR U31265 ( .A(n32434), .B(n32433), .Z(n32436) );
  XNOR U31266 ( .A(n32431), .B(n32430), .Z(n32433) );
  XNOR U31267 ( .A(n32428), .B(n32427), .Z(n32430) );
  XNOR U31268 ( .A(n32425), .B(n32424), .Z(n32427) );
  XNOR U31269 ( .A(n32422), .B(n32421), .Z(n32424) );
  XNOR U31270 ( .A(n32419), .B(n32418), .Z(n32421) );
  XNOR U31271 ( .A(n32416), .B(n32415), .Z(n32418) );
  XNOR U31272 ( .A(n32413), .B(n32412), .Z(n32415) );
  XNOR U31273 ( .A(n32410), .B(n32409), .Z(n32412) );
  XNOR U31274 ( .A(n32407), .B(n32406), .Z(n32409) );
  XNOR U31275 ( .A(n32404), .B(n32403), .Z(n32406) );
  XNOR U31276 ( .A(n32401), .B(n32400), .Z(n32403) );
  XNOR U31277 ( .A(n32398), .B(n32397), .Z(n32400) );
  XNOR U31278 ( .A(n32395), .B(n32394), .Z(n32397) );
  XNOR U31279 ( .A(n32392), .B(n32391), .Z(n32394) );
  XNOR U31280 ( .A(n32389), .B(n32388), .Z(n32391) );
  XNOR U31281 ( .A(n32386), .B(n32385), .Z(n32388) );
  XNOR U31282 ( .A(n32383), .B(n32382), .Z(n32385) );
  XNOR U31283 ( .A(n32380), .B(n32379), .Z(n32382) );
  XNOR U31284 ( .A(n32377), .B(n32376), .Z(n32379) );
  XNOR U31285 ( .A(n32374), .B(n32373), .Z(n32376) );
  XNOR U31286 ( .A(n32371), .B(n32370), .Z(n32373) );
  XNOR U31287 ( .A(n32368), .B(n32367), .Z(n32370) );
  XNOR U31288 ( .A(n32365), .B(n32364), .Z(n32367) );
  XNOR U31289 ( .A(n32362), .B(n32361), .Z(n32364) );
  XNOR U31290 ( .A(n32359), .B(n32358), .Z(n32361) );
  XNOR U31291 ( .A(n32356), .B(n32355), .Z(n32358) );
  XNOR U31292 ( .A(n32353), .B(n32352), .Z(n32355) );
  XNOR U31293 ( .A(n32350), .B(n32349), .Z(n32352) );
  XNOR U31294 ( .A(n32347), .B(n32346), .Z(n32349) );
  XNOR U31295 ( .A(n32344), .B(n32343), .Z(n32346) );
  XNOR U31296 ( .A(n32341), .B(n32340), .Z(n32343) );
  XNOR U31297 ( .A(n32338), .B(n32337), .Z(n32340) );
  XNOR U31298 ( .A(n32335), .B(n32334), .Z(n32337) );
  XNOR U31299 ( .A(n32332), .B(n32331), .Z(n32334) );
  XNOR U31300 ( .A(n32329), .B(n32328), .Z(n32331) );
  XNOR U31301 ( .A(n32326), .B(n32325), .Z(n32328) );
  XNOR U31302 ( .A(n32323), .B(n32322), .Z(n32325) );
  XNOR U31303 ( .A(n32320), .B(n32319), .Z(n32322) );
  XNOR U31304 ( .A(n32317), .B(n32316), .Z(n32319) );
  XNOR U31305 ( .A(n32314), .B(n32313), .Z(n32316) );
  XNOR U31306 ( .A(n32311), .B(n32310), .Z(n32313) );
  XNOR U31307 ( .A(n32308), .B(n32307), .Z(n32310) );
  XNOR U31308 ( .A(n32305), .B(n32304), .Z(n32307) );
  XNOR U31309 ( .A(n32302), .B(n32301), .Z(n32304) );
  XNOR U31310 ( .A(n32299), .B(n32298), .Z(n32301) );
  XNOR U31311 ( .A(n32296), .B(n32295), .Z(n32298) );
  XNOR U31312 ( .A(n32293), .B(n32292), .Z(n32295) );
  XNOR U31313 ( .A(n32290), .B(n32289), .Z(n32292) );
  XNOR U31314 ( .A(n32287), .B(n32286), .Z(n32289) );
  XNOR U31315 ( .A(n32284), .B(n32283), .Z(n32286) );
  XNOR U31316 ( .A(n32281), .B(n32280), .Z(n32283) );
  XNOR U31317 ( .A(n32278), .B(n32277), .Z(n32280) );
  XNOR U31318 ( .A(n32275), .B(n32274), .Z(n32277) );
  XNOR U31319 ( .A(n32272), .B(n32271), .Z(n32274) );
  XNOR U31320 ( .A(n32269), .B(n32268), .Z(n32271) );
  XNOR U31321 ( .A(n32266), .B(n32265), .Z(n32268) );
  XNOR U31322 ( .A(n32263), .B(n32262), .Z(n32265) );
  XNOR U31323 ( .A(n32260), .B(n32259), .Z(n32262) );
  XNOR U31324 ( .A(n32257), .B(n32256), .Z(n32259) );
  XNOR U31325 ( .A(n32254), .B(n32253), .Z(n32256) );
  XNOR U31326 ( .A(n32251), .B(n32250), .Z(n32253) );
  XNOR U31327 ( .A(n32248), .B(n32247), .Z(n32250) );
  XNOR U31328 ( .A(n32245), .B(n32244), .Z(n32247) );
  XNOR U31329 ( .A(n32242), .B(n32241), .Z(n32244) );
  XNOR U31330 ( .A(n32239), .B(n32238), .Z(n32241) );
  XNOR U31331 ( .A(n32236), .B(n32235), .Z(n32238) );
  XNOR U31332 ( .A(n32233), .B(n32232), .Z(n32235) );
  XNOR U31333 ( .A(n32230), .B(n32229), .Z(n32232) );
  XNOR U31334 ( .A(n32227), .B(n32226), .Z(n32229) );
  XNOR U31335 ( .A(n32224), .B(n32223), .Z(n32226) );
  XNOR U31336 ( .A(n32221), .B(n32220), .Z(n32223) );
  XNOR U31337 ( .A(n32218), .B(n32217), .Z(n32220) );
  XNOR U31338 ( .A(n32215), .B(n32214), .Z(n32217) );
  XNOR U31339 ( .A(n32212), .B(n32211), .Z(n32214) );
  XNOR U31340 ( .A(n32209), .B(n32208), .Z(n32211) );
  XNOR U31341 ( .A(n32206), .B(n32205), .Z(n32208) );
  XNOR U31342 ( .A(n32203), .B(n32202), .Z(n32205) );
  XNOR U31343 ( .A(n32200), .B(n32199), .Z(n32202) );
  XNOR U31344 ( .A(n32197), .B(n32196), .Z(n32199) );
  XNOR U31345 ( .A(n32194), .B(n32193), .Z(n32196) );
  XNOR U31346 ( .A(n32191), .B(n32190), .Z(n32193) );
  XNOR U31347 ( .A(n32188), .B(n32187), .Z(n32190) );
  XNOR U31348 ( .A(n32185), .B(n32184), .Z(n32187) );
  XNOR U31349 ( .A(n32182), .B(n32181), .Z(n32184) );
  XNOR U31350 ( .A(n32179), .B(n32178), .Z(n32181) );
  XNOR U31351 ( .A(n32176), .B(n32175), .Z(n32178) );
  XNOR U31352 ( .A(n32173), .B(n32172), .Z(n32175) );
  XNOR U31353 ( .A(n32170), .B(n32169), .Z(n32172) );
  XNOR U31354 ( .A(n32167), .B(n32166), .Z(n32169) );
  XNOR U31355 ( .A(n32164), .B(n32163), .Z(n32166) );
  XNOR U31356 ( .A(n32161), .B(n32160), .Z(n32163) );
  XNOR U31357 ( .A(n32158), .B(n32157), .Z(n32160) );
  XNOR U31358 ( .A(n32155), .B(n32154), .Z(n32157) );
  XNOR U31359 ( .A(n32152), .B(n32151), .Z(n32154) );
  XNOR U31360 ( .A(n32149), .B(n32148), .Z(n32151) );
  XNOR U31361 ( .A(n32146), .B(n32145), .Z(n32148) );
  XNOR U31362 ( .A(n32143), .B(n32142), .Z(n32145) );
  XNOR U31363 ( .A(n32140), .B(n32139), .Z(n32142) );
  XNOR U31364 ( .A(n32137), .B(n32136), .Z(n32139) );
  XNOR U31365 ( .A(n32134), .B(n32133), .Z(n32136) );
  XNOR U31366 ( .A(n32131), .B(n32130), .Z(n32133) );
  XNOR U31367 ( .A(n32128), .B(n32127), .Z(n32130) );
  XNOR U31368 ( .A(n32125), .B(n32124), .Z(n32127) );
  XNOR U31369 ( .A(n32122), .B(n32121), .Z(n32124) );
  XNOR U31370 ( .A(n32119), .B(n32118), .Z(n32121) );
  XNOR U31371 ( .A(n32116), .B(n32115), .Z(n32118) );
  XNOR U31372 ( .A(n32113), .B(n32112), .Z(n32115) );
  XNOR U31373 ( .A(n32110), .B(n32109), .Z(n32112) );
  XNOR U31374 ( .A(n32107), .B(n32106), .Z(n32109) );
  XNOR U31375 ( .A(n32104), .B(n32103), .Z(n32106) );
  XNOR U31376 ( .A(n32101), .B(n32100), .Z(n32103) );
  XNOR U31377 ( .A(n32098), .B(n32097), .Z(n32100) );
  XNOR U31378 ( .A(n32095), .B(n32094), .Z(n32097) );
  XNOR U31379 ( .A(n32092), .B(n32091), .Z(n32094) );
  XNOR U31380 ( .A(n32089), .B(n32088), .Z(n32091) );
  XNOR U31381 ( .A(n32086), .B(n32085), .Z(n32088) );
  XNOR U31382 ( .A(n32083), .B(n32082), .Z(n32085) );
  XNOR U31383 ( .A(n32080), .B(n32079), .Z(n32082) );
  XNOR U31384 ( .A(n32077), .B(n32076), .Z(n32079) );
  XNOR U31385 ( .A(n32074), .B(n32073), .Z(n32076) );
  XNOR U31386 ( .A(n32071), .B(n32070), .Z(n32073) );
  XNOR U31387 ( .A(n32068), .B(n32067), .Z(n32070) );
  XNOR U31388 ( .A(n32065), .B(n32064), .Z(n32067) );
  XNOR U31389 ( .A(n32062), .B(n32061), .Z(n32064) );
  XNOR U31390 ( .A(n32059), .B(n32058), .Z(n32061) );
  XNOR U31391 ( .A(n32056), .B(n32055), .Z(n32058) );
  XNOR U31392 ( .A(n32053), .B(n32052), .Z(n32055) );
  XNOR U31393 ( .A(n32050), .B(n32049), .Z(n32052) );
  XNOR U31394 ( .A(n32047), .B(n32046), .Z(n32049) );
  XNOR U31395 ( .A(n32044), .B(n32043), .Z(n32046) );
  XNOR U31396 ( .A(n32041), .B(n32040), .Z(n32043) );
  XNOR U31397 ( .A(n32038), .B(n32037), .Z(n32040) );
  XNOR U31398 ( .A(n32035), .B(n32034), .Z(n32037) );
  XNOR U31399 ( .A(n32032), .B(n32031), .Z(n32034) );
  XNOR U31400 ( .A(n32029), .B(n32028), .Z(n32031) );
  XNOR U31401 ( .A(n32026), .B(n32025), .Z(n32028) );
  XNOR U31402 ( .A(n32023), .B(n32022), .Z(n32025) );
  XNOR U31403 ( .A(n32020), .B(n32019), .Z(n32022) );
  XNOR U31404 ( .A(n32017), .B(n32016), .Z(n32019) );
  XNOR U31405 ( .A(n32014), .B(n32013), .Z(n32016) );
  XNOR U31406 ( .A(n32011), .B(n32010), .Z(n32013) );
  XNOR U31407 ( .A(n32008), .B(n32007), .Z(n32010) );
  XNOR U31408 ( .A(n32005), .B(n32004), .Z(n32007) );
  XNOR U31409 ( .A(n32002), .B(n32001), .Z(n32004) );
  XNOR U31410 ( .A(n31999), .B(n31998), .Z(n32001) );
  XNOR U31411 ( .A(n31996), .B(n31995), .Z(n31998) );
  XNOR U31412 ( .A(n31993), .B(n31992), .Z(n31995) );
  XNOR U31413 ( .A(n31990), .B(n31989), .Z(n31992) );
  XNOR U31414 ( .A(n31987), .B(n31986), .Z(n31989) );
  XNOR U31415 ( .A(n31984), .B(n31983), .Z(n31986) );
  XNOR U31416 ( .A(n31981), .B(n31980), .Z(n31983) );
  XNOR U31417 ( .A(n31978), .B(n31977), .Z(n31980) );
  XNOR U31418 ( .A(n31975), .B(n31974), .Z(n31977) );
  XNOR U31419 ( .A(n31972), .B(n31971), .Z(n31974) );
  XNOR U31420 ( .A(n31969), .B(n31968), .Z(n31971) );
  XNOR U31421 ( .A(n31966), .B(n31965), .Z(n31968) );
  XNOR U31422 ( .A(n31963), .B(n31962), .Z(n31965) );
  XNOR U31423 ( .A(n31960), .B(n31959), .Z(n31962) );
  XNOR U31424 ( .A(n31957), .B(n31956), .Z(n31959) );
  XNOR U31425 ( .A(n31954), .B(n31953), .Z(n31956) );
  XNOR U31426 ( .A(n31951), .B(n31950), .Z(n31953) );
  XNOR U31427 ( .A(n31948), .B(n31947), .Z(n31950) );
  XNOR U31428 ( .A(n31945), .B(n31944), .Z(n31947) );
  XNOR U31429 ( .A(n31942), .B(n31941), .Z(n31944) );
  XNOR U31430 ( .A(n31939), .B(n31938), .Z(n31941) );
  XNOR U31431 ( .A(n31936), .B(n31935), .Z(n31938) );
  XNOR U31432 ( .A(n31933), .B(n31932), .Z(n31935) );
  XNOR U31433 ( .A(n31930), .B(n31929), .Z(n31932) );
  XNOR U31434 ( .A(n31927), .B(n31926), .Z(n31929) );
  XNOR U31435 ( .A(n31924), .B(n31923), .Z(n31926) );
  XNOR U31436 ( .A(n31921), .B(n31920), .Z(n31923) );
  XNOR U31437 ( .A(n31918), .B(n31917), .Z(n31920) );
  XNOR U31438 ( .A(n31915), .B(n31914), .Z(n31917) );
  XNOR U31439 ( .A(n31912), .B(n31911), .Z(n31914) );
  XNOR U31440 ( .A(n31909), .B(n31908), .Z(n31911) );
  XNOR U31441 ( .A(n31906), .B(n31905), .Z(n31908) );
  XNOR U31442 ( .A(n31903), .B(n31902), .Z(n31905) );
  XNOR U31443 ( .A(n31900), .B(n31899), .Z(n31902) );
  XNOR U31444 ( .A(n31897), .B(n31896), .Z(n31899) );
  XNOR U31445 ( .A(n31894), .B(n31893), .Z(n31896) );
  XNOR U31446 ( .A(n31891), .B(n31890), .Z(n31893) );
  XNOR U31447 ( .A(n31888), .B(n31887), .Z(n31890) );
  XNOR U31448 ( .A(n31885), .B(n31884), .Z(n31887) );
  XNOR U31449 ( .A(n31882), .B(n31881), .Z(n31884) );
  XNOR U31450 ( .A(n31879), .B(n31878), .Z(n31881) );
  XNOR U31451 ( .A(n31876), .B(n31875), .Z(n31878) );
  XNOR U31452 ( .A(n31873), .B(n31872), .Z(n31875) );
  XNOR U31453 ( .A(n31870), .B(n31869), .Z(n31872) );
  XNOR U31454 ( .A(n31867), .B(n31866), .Z(n31869) );
  XNOR U31455 ( .A(n31864), .B(n31863), .Z(n31866) );
  XNOR U31456 ( .A(n31861), .B(n31860), .Z(n31863) );
  XNOR U31457 ( .A(n31858), .B(n31857), .Z(n31860) );
  XNOR U31458 ( .A(n31855), .B(n31854), .Z(n31857) );
  XNOR U31459 ( .A(n31852), .B(n31851), .Z(n31854) );
  XNOR U31460 ( .A(n31849), .B(n31848), .Z(n31851) );
  XNOR U31461 ( .A(n31846), .B(n31845), .Z(n31848) );
  XNOR U31462 ( .A(n31843), .B(n31842), .Z(n31845) );
  XNOR U31463 ( .A(n31840), .B(n31839), .Z(n31842) );
  XNOR U31464 ( .A(n31837), .B(n31836), .Z(n31839) );
  XNOR U31465 ( .A(n31834), .B(n31833), .Z(n31836) );
  XNOR U31466 ( .A(n31831), .B(n31830), .Z(n31833) );
  XNOR U31467 ( .A(n31828), .B(n31827), .Z(n31830) );
  XNOR U31468 ( .A(n31825), .B(n31824), .Z(n31827) );
  XNOR U31469 ( .A(n31822), .B(n31821), .Z(n31824) );
  XNOR U31470 ( .A(n31819), .B(n31818), .Z(n31821) );
  XNOR U31471 ( .A(n31816), .B(n31815), .Z(n31818) );
  XNOR U31472 ( .A(n31813), .B(n31812), .Z(n31815) );
  XNOR U31473 ( .A(n31810), .B(n31809), .Z(n31812) );
  XNOR U31474 ( .A(n31807), .B(n31806), .Z(n31809) );
  XNOR U31475 ( .A(n31804), .B(n31803), .Z(n31806) );
  XNOR U31476 ( .A(n31801), .B(n31800), .Z(n31803) );
  XNOR U31477 ( .A(n31798), .B(n31797), .Z(n31800) );
  XNOR U31478 ( .A(n31795), .B(n31794), .Z(n31797) );
  XNOR U31479 ( .A(n31792), .B(n31791), .Z(n31794) );
  XNOR U31480 ( .A(n31789), .B(n31788), .Z(n31791) );
  XNOR U31481 ( .A(n31786), .B(n31785), .Z(n31788) );
  XNOR U31482 ( .A(n31783), .B(n31782), .Z(n31785) );
  XNOR U31483 ( .A(n31780), .B(n31779), .Z(n31782) );
  XNOR U31484 ( .A(n31777), .B(n31776), .Z(n31779) );
  XNOR U31485 ( .A(n31774), .B(n31773), .Z(n31776) );
  XNOR U31486 ( .A(n31771), .B(n31770), .Z(n31773) );
  XNOR U31487 ( .A(n31768), .B(n31767), .Z(n31770) );
  XNOR U31488 ( .A(n31765), .B(n31764), .Z(n31767) );
  XNOR U31489 ( .A(n31762), .B(n31761), .Z(n31764) );
  XNOR U31490 ( .A(n31759), .B(n31758), .Z(n31761) );
  XNOR U31491 ( .A(n31756), .B(n31755), .Z(n31758) );
  XNOR U31492 ( .A(n31753), .B(n31752), .Z(n31755) );
  XNOR U31493 ( .A(n31750), .B(n31749), .Z(n31752) );
  XNOR U31494 ( .A(n31747), .B(n31746), .Z(n31749) );
  XNOR U31495 ( .A(n31744), .B(n31743), .Z(n31746) );
  XNOR U31496 ( .A(n31741), .B(n31740), .Z(n31743) );
  XNOR U31497 ( .A(n31738), .B(n31737), .Z(n31740) );
  XNOR U31498 ( .A(n31735), .B(n31734), .Z(n31737) );
  XNOR U31499 ( .A(n31732), .B(n31731), .Z(n31734) );
  XNOR U31500 ( .A(n31729), .B(n31728), .Z(n31731) );
  XNOR U31501 ( .A(n31726), .B(n31725), .Z(n31728) );
  XNOR U31502 ( .A(n31723), .B(n31722), .Z(n31725) );
  XNOR U31503 ( .A(n31720), .B(n31719), .Z(n31722) );
  XNOR U31504 ( .A(n31717), .B(n31716), .Z(n31719) );
  XNOR U31505 ( .A(n31714), .B(n31713), .Z(n31716) );
  XNOR U31506 ( .A(n31711), .B(n31710), .Z(n31713) );
  XNOR U31507 ( .A(n31708), .B(n31707), .Z(n31710) );
  XNOR U31508 ( .A(n31705), .B(n31704), .Z(n31707) );
  XNOR U31509 ( .A(n31702), .B(n31701), .Z(n31704) );
  XNOR U31510 ( .A(n31699), .B(n31698), .Z(n31701) );
  XNOR U31511 ( .A(n31696), .B(n31695), .Z(n31698) );
  XNOR U31512 ( .A(n31693), .B(n31692), .Z(n31695) );
  XNOR U31513 ( .A(n31690), .B(n31689), .Z(n31692) );
  XNOR U31514 ( .A(n31687), .B(n31686), .Z(n31689) );
  XNOR U31515 ( .A(n31684), .B(n31683), .Z(n31686) );
  XNOR U31516 ( .A(n31681), .B(n31680), .Z(n31683) );
  XNOR U31517 ( .A(n31678), .B(n31677), .Z(n31680) );
  XNOR U31518 ( .A(n31675), .B(n31674), .Z(n31677) );
  XNOR U31519 ( .A(n31672), .B(n31671), .Z(n31674) );
  XNOR U31520 ( .A(n31669), .B(n31668), .Z(n31671) );
  XNOR U31521 ( .A(n31666), .B(n31665), .Z(n31668) );
  XNOR U31522 ( .A(n31663), .B(n31662), .Z(n31665) );
  XNOR U31523 ( .A(n31660), .B(n31659), .Z(n31662) );
  XNOR U31524 ( .A(n31657), .B(n31656), .Z(n31659) );
  XNOR U31525 ( .A(n31654), .B(n31653), .Z(n31656) );
  XNOR U31526 ( .A(n31651), .B(n31650), .Z(n31653) );
  XNOR U31527 ( .A(n31648), .B(n31647), .Z(n31650) );
  XNOR U31528 ( .A(n31645), .B(n31644), .Z(n31647) );
  XNOR U31529 ( .A(n31642), .B(n31641), .Z(n31644) );
  XNOR U31530 ( .A(n31639), .B(n31638), .Z(n31641) );
  XNOR U31531 ( .A(n31636), .B(n31635), .Z(n31638) );
  XNOR U31532 ( .A(n31633), .B(n31632), .Z(n31635) );
  XNOR U31533 ( .A(n31630), .B(n31629), .Z(n31632) );
  XNOR U31534 ( .A(n31627), .B(n31626), .Z(n31629) );
  XNOR U31535 ( .A(n31624), .B(n31623), .Z(n31626) );
  XNOR U31536 ( .A(n31621), .B(n31620), .Z(n31623) );
  XNOR U31537 ( .A(n31618), .B(n31617), .Z(n31620) );
  XNOR U31538 ( .A(n31615), .B(n31614), .Z(n31617) );
  XNOR U31539 ( .A(n31612), .B(n31611), .Z(n31614) );
  XNOR U31540 ( .A(n31609), .B(n31608), .Z(n31611) );
  XNOR U31541 ( .A(n31606), .B(n31605), .Z(n31608) );
  XNOR U31542 ( .A(n31603), .B(n31602), .Z(n31605) );
  XNOR U31543 ( .A(n31600), .B(n31599), .Z(n31602) );
  XNOR U31544 ( .A(n31597), .B(n31596), .Z(n31599) );
  XNOR U31545 ( .A(n31594), .B(n31593), .Z(n31596) );
  XNOR U31546 ( .A(n31591), .B(n31590), .Z(n31593) );
  XNOR U31547 ( .A(n31588), .B(n31587), .Z(n31590) );
  XNOR U31548 ( .A(n31585), .B(n31584), .Z(n31587) );
  XNOR U31549 ( .A(n31582), .B(n31581), .Z(n31584) );
  XNOR U31550 ( .A(n31579), .B(n31578), .Z(n31581) );
  XNOR U31551 ( .A(n31576), .B(n31575), .Z(n31578) );
  XNOR U31552 ( .A(n31573), .B(n31572), .Z(n31575) );
  XNOR U31553 ( .A(n31570), .B(n31569), .Z(n31572) );
  XNOR U31554 ( .A(n31567), .B(n31566), .Z(n31569) );
  XNOR U31555 ( .A(n31564), .B(n31563), .Z(n31566) );
  XNOR U31556 ( .A(n31561), .B(n31560), .Z(n31563) );
  XNOR U31557 ( .A(n31558), .B(n31557), .Z(n31560) );
  XNOR U31558 ( .A(n31555), .B(n31554), .Z(n31557) );
  XNOR U31559 ( .A(n31552), .B(n31551), .Z(n31554) );
  XNOR U31560 ( .A(n31549), .B(n31548), .Z(n31551) );
  XNOR U31561 ( .A(n31546), .B(n31545), .Z(n31548) );
  XNOR U31562 ( .A(n31543), .B(n31542), .Z(n31545) );
  XNOR U31563 ( .A(n31540), .B(n31539), .Z(n31542) );
  XNOR U31564 ( .A(n31537), .B(n31536), .Z(n31539) );
  XNOR U31565 ( .A(n31534), .B(n31533), .Z(n31536) );
  XNOR U31566 ( .A(n31531), .B(n31530), .Z(n31533) );
  XNOR U31567 ( .A(n31528), .B(n31527), .Z(n31530) );
  XNOR U31568 ( .A(n31525), .B(n31524), .Z(n31527) );
  XNOR U31569 ( .A(n31522), .B(n31521), .Z(n31524) );
  XNOR U31570 ( .A(n31519), .B(n31518), .Z(n31521) );
  XNOR U31571 ( .A(n31516), .B(n31515), .Z(n31518) );
  XNOR U31572 ( .A(n31513), .B(n31512), .Z(n31515) );
  XOR U31573 ( .A(n34106), .B(n31509), .Z(n31512) );
  XOR U31574 ( .A(n31507), .B(n31506), .Z(n31509) );
  XOR U31575 ( .A(n31504), .B(n31503), .Z(n31506) );
  XOR U31576 ( .A(n31500), .B(n31501), .Z(n31503) );
  AND U31577 ( .A(n34107), .B(n34108), .Z(n31501) );
  XOR U31578 ( .A(n31497), .B(n31498), .Z(n31500) );
  AND U31579 ( .A(n34109), .B(n34110), .Z(n31498) );
  XOR U31580 ( .A(n31494), .B(n31495), .Z(n31497) );
  AND U31581 ( .A(n34111), .B(n34112), .Z(n31495) );
  XOR U31582 ( .A(n31491), .B(n31492), .Z(n31494) );
  AND U31583 ( .A(n34113), .B(n34114), .Z(n31492) );
  XNOR U31584 ( .A(n31275), .B(n31489), .Z(n31491) );
  AND U31585 ( .A(n34115), .B(n34116), .Z(n31489) );
  XOR U31586 ( .A(n31277), .B(n31276), .Z(n31275) );
  AND U31587 ( .A(n34117), .B(n34118), .Z(n31276) );
  XOR U31588 ( .A(n31279), .B(n31278), .Z(n31277) );
  AND U31589 ( .A(n34119), .B(n34120), .Z(n31278) );
  XOR U31590 ( .A(n31281), .B(n31280), .Z(n31279) );
  AND U31591 ( .A(n34121), .B(n34122), .Z(n31280) );
  XOR U31592 ( .A(n31283), .B(n31282), .Z(n31281) );
  AND U31593 ( .A(n34123), .B(n34124), .Z(n31282) );
  XOR U31594 ( .A(n31285), .B(n31284), .Z(n31283) );
  AND U31595 ( .A(n34125), .B(n34126), .Z(n31284) );
  XOR U31596 ( .A(n31287), .B(n31286), .Z(n31285) );
  AND U31597 ( .A(n34127), .B(n34128), .Z(n31286) );
  XOR U31598 ( .A(n31289), .B(n31288), .Z(n31287) );
  AND U31599 ( .A(n34129), .B(n34130), .Z(n31288) );
  XOR U31600 ( .A(n31291), .B(n31290), .Z(n31289) );
  AND U31601 ( .A(n34131), .B(n34132), .Z(n31290) );
  XOR U31602 ( .A(n31293), .B(n31292), .Z(n31291) );
  AND U31603 ( .A(n34133), .B(n34134), .Z(n31292) );
  XOR U31604 ( .A(n31295), .B(n31294), .Z(n31293) );
  AND U31605 ( .A(n34135), .B(n34136), .Z(n31294) );
  XOR U31606 ( .A(n31297), .B(n31296), .Z(n31295) );
  AND U31607 ( .A(n34137), .B(n34138), .Z(n31296) );
  XOR U31608 ( .A(n31299), .B(n31298), .Z(n31297) );
  AND U31609 ( .A(n34139), .B(n34140), .Z(n31298) );
  XOR U31610 ( .A(n31301), .B(n31300), .Z(n31299) );
  AND U31611 ( .A(n34141), .B(n34142), .Z(n31300) );
  XOR U31612 ( .A(n31303), .B(n31302), .Z(n31301) );
  AND U31613 ( .A(n34143), .B(n34144), .Z(n31302) );
  XOR U31614 ( .A(n31305), .B(n31304), .Z(n31303) );
  AND U31615 ( .A(n34145), .B(n34146), .Z(n31304) );
  XOR U31616 ( .A(n31307), .B(n31306), .Z(n31305) );
  AND U31617 ( .A(n34147), .B(n34148), .Z(n31306) );
  XOR U31618 ( .A(n31309), .B(n31308), .Z(n31307) );
  AND U31619 ( .A(n34149), .B(n34150), .Z(n31308) );
  XOR U31620 ( .A(n31311), .B(n31310), .Z(n31309) );
  AND U31621 ( .A(n34151), .B(n34152), .Z(n31310) );
  XOR U31622 ( .A(n31313), .B(n31312), .Z(n31311) );
  AND U31623 ( .A(n34153), .B(n34154), .Z(n31312) );
  XOR U31624 ( .A(n31315), .B(n31314), .Z(n31313) );
  AND U31625 ( .A(n34155), .B(n34156), .Z(n31314) );
  XOR U31626 ( .A(n31317), .B(n31316), .Z(n31315) );
  AND U31627 ( .A(n34157), .B(n34158), .Z(n31316) );
  XOR U31628 ( .A(n31319), .B(n31318), .Z(n31317) );
  AND U31629 ( .A(n34159), .B(n34160), .Z(n31318) );
  XOR U31630 ( .A(n31321), .B(n31320), .Z(n31319) );
  AND U31631 ( .A(n34161), .B(n34162), .Z(n31320) );
  XOR U31632 ( .A(n31323), .B(n31322), .Z(n31321) );
  AND U31633 ( .A(n34163), .B(n34164), .Z(n31322) );
  XOR U31634 ( .A(n31325), .B(n31324), .Z(n31323) );
  AND U31635 ( .A(n34165), .B(n34166), .Z(n31324) );
  XOR U31636 ( .A(n31327), .B(n31326), .Z(n31325) );
  AND U31637 ( .A(n34167), .B(n34168), .Z(n31326) );
  XOR U31638 ( .A(n31329), .B(n31328), .Z(n31327) );
  AND U31639 ( .A(n34169), .B(n34170), .Z(n31328) );
  XOR U31640 ( .A(n31331), .B(n31330), .Z(n31329) );
  AND U31641 ( .A(n34171), .B(n34172), .Z(n31330) );
  XOR U31642 ( .A(n31333), .B(n31332), .Z(n31331) );
  AND U31643 ( .A(n34173), .B(n34174), .Z(n31332) );
  XOR U31644 ( .A(n31335), .B(n31334), .Z(n31333) );
  AND U31645 ( .A(n34175), .B(n34176), .Z(n31334) );
  XOR U31646 ( .A(n31337), .B(n31336), .Z(n31335) );
  AND U31647 ( .A(n34177), .B(n34178), .Z(n31336) );
  XOR U31648 ( .A(n31339), .B(n31338), .Z(n31337) );
  AND U31649 ( .A(n34179), .B(n34180), .Z(n31338) );
  XOR U31650 ( .A(n31341), .B(n31340), .Z(n31339) );
  AND U31651 ( .A(n34181), .B(n34182), .Z(n31340) );
  XOR U31652 ( .A(n31343), .B(n31342), .Z(n31341) );
  AND U31653 ( .A(n34183), .B(n34184), .Z(n31342) );
  XOR U31654 ( .A(n31345), .B(n31344), .Z(n31343) );
  AND U31655 ( .A(n34185), .B(n34186), .Z(n31344) );
  XOR U31656 ( .A(n31347), .B(n31346), .Z(n31345) );
  AND U31657 ( .A(n34187), .B(n34188), .Z(n31346) );
  XOR U31658 ( .A(n31349), .B(n31348), .Z(n31347) );
  AND U31659 ( .A(n34189), .B(n34190), .Z(n31348) );
  XOR U31660 ( .A(n31351), .B(n31350), .Z(n31349) );
  AND U31661 ( .A(n34191), .B(n34192), .Z(n31350) );
  XOR U31662 ( .A(n31353), .B(n31352), .Z(n31351) );
  AND U31663 ( .A(n34193), .B(n34194), .Z(n31352) );
  XOR U31664 ( .A(n31355), .B(n31354), .Z(n31353) );
  AND U31665 ( .A(n34195), .B(n34196), .Z(n31354) );
  XOR U31666 ( .A(n31358), .B(n31356), .Z(n31355) );
  AND U31667 ( .A(n34197), .B(n34198), .Z(n31356) );
  XOR U31668 ( .A(n31379), .B(n31359), .Z(n31358) );
  AND U31669 ( .A(n34199), .B(n34200), .Z(n31359) );
  XOR U31670 ( .A(n31375), .B(n31380), .Z(n31379) );
  AND U31671 ( .A(n34201), .B(n34202), .Z(n31380) );
  XOR U31672 ( .A(n31377), .B(n31376), .Z(n31375) );
  AND U31673 ( .A(n34203), .B(n34204), .Z(n31376) );
  XOR U31674 ( .A(n31364), .B(n31378), .Z(n31377) );
  AND U31675 ( .A(n34205), .B(n34206), .Z(n31378) );
  XOR U31676 ( .A(n31366), .B(n31365), .Z(n31364) );
  AND U31677 ( .A(n34207), .B(n34208), .Z(n31365) );
  XOR U31678 ( .A(n31369), .B(n31367), .Z(n31366) );
  AND U31679 ( .A(n34209), .B(n34210), .Z(n31367) );
  XOR U31680 ( .A(n31371), .B(n31370), .Z(n31369) );
  AND U31681 ( .A(n34211), .B(n34212), .Z(n31370) );
  XOR U31682 ( .A(n31389), .B(n31372), .Z(n31371) );
  AND U31683 ( .A(n34213), .B(n34214), .Z(n31372) );
  XNOR U31684 ( .A(n31396), .B(n31390), .Z(n31389) );
  AND U31685 ( .A(n34215), .B(n34216), .Z(n31390) );
  XOR U31686 ( .A(n31395), .B(n31387), .Z(n31396) );
  AND U31687 ( .A(n34217), .B(n34218), .Z(n31387) );
  XOR U31688 ( .A(n31488), .B(n31386), .Z(n31395) );
  AND U31689 ( .A(n34219), .B(n34220), .Z(n31386) );
  XNOR U31690 ( .A(n31407), .B(n31385), .Z(n31488) );
  AND U31691 ( .A(n34221), .B(n34222), .Z(n31385) );
  XNOR U31692 ( .A(n31414), .B(n31408), .Z(n31407) );
  AND U31693 ( .A(n34223), .B(n34224), .Z(n31408) );
  XOR U31694 ( .A(n31413), .B(n31405), .Z(n31414) );
  AND U31695 ( .A(n34225), .B(n34226), .Z(n31405) );
  XOR U31696 ( .A(n31487), .B(n31404), .Z(n31413) );
  AND U31697 ( .A(n34227), .B(n34228), .Z(n31404) );
  XNOR U31698 ( .A(n31425), .B(n31403), .Z(n31487) );
  AND U31699 ( .A(n34229), .B(n34230), .Z(n31403) );
  XNOR U31700 ( .A(n31432), .B(n31426), .Z(n31425) );
  AND U31701 ( .A(n34231), .B(n34232), .Z(n31426) );
  XOR U31702 ( .A(n31431), .B(n31423), .Z(n31432) );
  AND U31703 ( .A(n34233), .B(n34234), .Z(n31423) );
  XOR U31704 ( .A(n31486), .B(n31422), .Z(n31431) );
  AND U31705 ( .A(n34235), .B(n34236), .Z(n31422) );
  XNOR U31706 ( .A(n31443), .B(n31421), .Z(n31486) );
  AND U31707 ( .A(n34237), .B(n34238), .Z(n31421) );
  XNOR U31708 ( .A(n31450), .B(n31444), .Z(n31443) );
  AND U31709 ( .A(n34239), .B(n34240), .Z(n31444) );
  XOR U31710 ( .A(n31449), .B(n31441), .Z(n31450) );
  AND U31711 ( .A(n34241), .B(n34242), .Z(n31441) );
  XOR U31712 ( .A(n31485), .B(n31440), .Z(n31449) );
  AND U31713 ( .A(n34243), .B(n34244), .Z(n31440) );
  XNOR U31714 ( .A(n34245), .B(n34246), .Z(n31485) );
  XOR U31715 ( .A(n31483), .B(n31484), .Z(n34246) );
  AND U31716 ( .A(n34247), .B(n34248), .Z(n31484) );
  AND U31717 ( .A(n34249), .B(n34250), .Z(n31483) );
  XOR U31718 ( .A(n34251), .B(n31439), .Z(n34245) );
  AND U31719 ( .A(n34252), .B(n34253), .Z(n31439) );
  XOR U31720 ( .A(n34254), .B(n34255), .Z(n34251) );
  XOR U31721 ( .A(n34256), .B(n34257), .Z(n34255) );
  XOR U31722 ( .A(n31476), .B(n31477), .Z(n34257) );
  AND U31723 ( .A(n34258), .B(n34259), .Z(n31477) );
  AND U31724 ( .A(n34260), .B(n34261), .Z(n31476) );
  XOR U31725 ( .A(n31470), .B(n31475), .Z(n34256) );
  AND U31726 ( .A(n34262), .B(n34263), .Z(n31475) );
  AND U31727 ( .A(n34264), .B(n34265), .Z(n31470) );
  XOR U31728 ( .A(n34266), .B(n34267), .Z(n34254) );
  XOR U31729 ( .A(n31478), .B(n31481), .Z(n34267) );
  AND U31730 ( .A(n34268), .B(n34269), .Z(n31481) );
  AND U31731 ( .A(n34270), .B(n34271), .Z(n31478) );
  XOR U31732 ( .A(n34272), .B(n31482), .Z(n34266) );
  AND U31733 ( .A(n34273), .B(n34274), .Z(n31482) );
  XOR U31734 ( .A(n34275), .B(n34276), .Z(n34272) );
  XOR U31735 ( .A(n34277), .B(n34278), .Z(n34276) );
  XOR U31736 ( .A(n31463), .B(n31464), .Z(n34278) );
  AND U31737 ( .A(n34279), .B(n34280), .Z(n31464) );
  AND U31738 ( .A(n34281), .B(n34282), .Z(n31463) );
  XNOR U31739 ( .A(n31461), .B(n31460), .Z(n34277) );
  IV U31740 ( .A(n34283), .Z(n31460) );
  AND U31741 ( .A(n34284), .B(n34285), .Z(n34283) );
  AND U31742 ( .A(n34286), .B(n34287), .Z(n31461) );
  XOR U31743 ( .A(n34288), .B(n34289), .Z(n34275) );
  XOR U31744 ( .A(n31467), .B(n31468), .Z(n34289) );
  AND U31745 ( .A(n34290), .B(n34291), .Z(n31468) );
  AND U31746 ( .A(n34292), .B(n34293), .Z(n31467) );
  XOR U31747 ( .A(n31462), .B(n31469), .Z(n34288) );
  AND U31748 ( .A(n34294), .B(n34295), .Z(n31469) );
  XNOR U31749 ( .A(n34296), .B(n34297), .Z(n31462) );
  AND U31750 ( .A(n34298), .B(n34299), .Z(n34297) );
  NOR U31751 ( .A(n34300), .B(n34301), .Z(n34299) );
  NOR U31752 ( .A(n34302), .B(n34303), .Z(n34298) );
  AND U31753 ( .A(n34304), .B(n34305), .Z(n34303) );
  AND U31754 ( .A(n34306), .B(n34307), .Z(n34296) );
  NOR U31755 ( .A(n34308), .B(n34309), .Z(n34307) );
  AND U31756 ( .A(n34301), .B(n34310), .Z(n34309) );
  AND U31757 ( .A(n34302), .B(n34311), .Z(n34308) );
  NOR U31758 ( .A(n34312), .B(n34313), .Z(n34306) );
  XOR U31759 ( .A(n34314), .B(n34315), .Z(n34313) );
  AND U31760 ( .A(n34316), .B(n34317), .Z(n34315) );
  NOR U31761 ( .A(n34318), .B(n34319), .Z(n34317) );
  NOR U31762 ( .A(n34320), .B(n34321), .Z(n34316) );
  AND U31763 ( .A(n34322), .B(n34323), .Z(n34321) );
  AND U31764 ( .A(n34324), .B(n34325), .Z(n34314) );
  NOR U31765 ( .A(n34326), .B(n34327), .Z(n34325) );
  AND U31766 ( .A(n34319), .B(n34328), .Z(n34327) );
  AND U31767 ( .A(n34320), .B(n34329), .Z(n34326) );
  NOR U31768 ( .A(n34330), .B(n34331), .Z(n34324) );
  AND U31769 ( .A(n34332), .B(n34333), .Z(n34331) );
  AND U31770 ( .A(n34334), .B(n34335), .Z(n34333) );
  AND U31771 ( .A(n34336), .B(n34337), .Z(n34335) );
  NOR U31772 ( .A(n34338), .B(n34339), .Z(n34336) );
  NOR U31773 ( .A(n34340), .B(n34341), .Z(n34334) );
  AND U31774 ( .A(n34342), .B(n34343), .Z(n34332) );
  NOR U31775 ( .A(n34344), .B(n34345), .Z(n34343) );
  NOR U31776 ( .A(n34346), .B(n34347), .Z(n34342) );
  AND U31777 ( .A(n34318), .B(n34348), .Z(n34330) );
  AND U31778 ( .A(n34300), .B(n34349), .Z(n34312) );
  XOR U31779 ( .A(n34350), .B(n34351), .Z(n31504) );
  AND U31780 ( .A(n34350), .B(n34352), .Z(n34351) );
  XNOR U31781 ( .A(n34353), .B(n34354), .Z(n31507) );
  AND U31782 ( .A(n34353), .B(n34355), .Z(n34354) );
  IV U31783 ( .A(n31510), .Z(n34106) );
  XNOR U31784 ( .A(n34356), .B(n34357), .Z(n31510) );
  AND U31785 ( .A(n34356), .B(n34358), .Z(n34357) );
  XNOR U31786 ( .A(n34359), .B(n34360), .Z(n31513) );
  AND U31787 ( .A(n34359), .B(n34361), .Z(n34360) );
  XNOR U31788 ( .A(n34362), .B(n34363), .Z(n31516) );
  AND U31789 ( .A(n34364), .B(n34362), .Z(n34363) );
  XOR U31790 ( .A(n34365), .B(n34366), .Z(n31519) );
  NOR U31791 ( .A(n34367), .B(n34365), .Z(n34366) );
  XOR U31792 ( .A(n34368), .B(n34369), .Z(n31522) );
  NOR U31793 ( .A(n34370), .B(n34368), .Z(n34369) );
  XOR U31794 ( .A(n34371), .B(n34372), .Z(n31525) );
  NOR U31795 ( .A(n34373), .B(n34371), .Z(n34372) );
  XOR U31796 ( .A(n34374), .B(n34375), .Z(n31528) );
  NOR U31797 ( .A(n34376), .B(n34374), .Z(n34375) );
  XOR U31798 ( .A(n34377), .B(n34378), .Z(n31531) );
  NOR U31799 ( .A(n34379), .B(n34377), .Z(n34378) );
  XOR U31800 ( .A(n34380), .B(n34381), .Z(n31534) );
  NOR U31801 ( .A(n34382), .B(n34380), .Z(n34381) );
  XOR U31802 ( .A(n34383), .B(n34384), .Z(n31537) );
  NOR U31803 ( .A(n34385), .B(n34383), .Z(n34384) );
  XOR U31804 ( .A(n34386), .B(n34387), .Z(n31540) );
  NOR U31805 ( .A(n34388), .B(n34386), .Z(n34387) );
  XOR U31806 ( .A(n34389), .B(n34390), .Z(n31543) );
  NOR U31807 ( .A(n34391), .B(n34389), .Z(n34390) );
  XOR U31808 ( .A(n34392), .B(n34393), .Z(n31546) );
  NOR U31809 ( .A(n34394), .B(n34392), .Z(n34393) );
  XOR U31810 ( .A(n34395), .B(n34396), .Z(n31549) );
  NOR U31811 ( .A(n34397), .B(n34395), .Z(n34396) );
  XOR U31812 ( .A(n34398), .B(n34399), .Z(n31552) );
  NOR U31813 ( .A(n34400), .B(n34398), .Z(n34399) );
  XOR U31814 ( .A(n34401), .B(n34402), .Z(n31555) );
  NOR U31815 ( .A(n34403), .B(n34401), .Z(n34402) );
  XOR U31816 ( .A(n34404), .B(n34405), .Z(n31558) );
  NOR U31817 ( .A(n34406), .B(n34404), .Z(n34405) );
  XOR U31818 ( .A(n34407), .B(n34408), .Z(n31561) );
  NOR U31819 ( .A(n34409), .B(n34407), .Z(n34408) );
  XOR U31820 ( .A(n34410), .B(n34411), .Z(n31564) );
  NOR U31821 ( .A(n34412), .B(n34410), .Z(n34411) );
  XOR U31822 ( .A(n34413), .B(n34414), .Z(n31567) );
  NOR U31823 ( .A(n34415), .B(n34413), .Z(n34414) );
  XOR U31824 ( .A(n34416), .B(n34417), .Z(n31570) );
  NOR U31825 ( .A(n34418), .B(n34416), .Z(n34417) );
  XOR U31826 ( .A(n34419), .B(n34420), .Z(n31573) );
  NOR U31827 ( .A(n34421), .B(n34419), .Z(n34420) );
  XOR U31828 ( .A(n34422), .B(n34423), .Z(n31576) );
  NOR U31829 ( .A(n34424), .B(n34422), .Z(n34423) );
  XOR U31830 ( .A(n34425), .B(n34426), .Z(n31579) );
  NOR U31831 ( .A(n34427), .B(n34425), .Z(n34426) );
  XOR U31832 ( .A(n34428), .B(n34429), .Z(n31582) );
  NOR U31833 ( .A(n34430), .B(n34428), .Z(n34429) );
  XOR U31834 ( .A(n34431), .B(n34432), .Z(n31585) );
  NOR U31835 ( .A(n34433), .B(n34431), .Z(n34432) );
  XOR U31836 ( .A(n34434), .B(n34435), .Z(n31588) );
  NOR U31837 ( .A(n34436), .B(n34434), .Z(n34435) );
  XOR U31838 ( .A(n34437), .B(n34438), .Z(n31591) );
  NOR U31839 ( .A(n34439), .B(n34437), .Z(n34438) );
  XOR U31840 ( .A(n34440), .B(n34441), .Z(n31594) );
  NOR U31841 ( .A(n34442), .B(n34440), .Z(n34441) );
  XOR U31842 ( .A(n34443), .B(n34444), .Z(n31597) );
  NOR U31843 ( .A(n34445), .B(n34443), .Z(n34444) );
  XOR U31844 ( .A(n34446), .B(n34447), .Z(n31600) );
  NOR U31845 ( .A(n34448), .B(n34446), .Z(n34447) );
  XOR U31846 ( .A(n34449), .B(n34450), .Z(n31603) );
  NOR U31847 ( .A(n34451), .B(n34449), .Z(n34450) );
  XOR U31848 ( .A(n34452), .B(n34453), .Z(n31606) );
  NOR U31849 ( .A(n34454), .B(n34452), .Z(n34453) );
  XOR U31850 ( .A(n34455), .B(n34456), .Z(n31609) );
  NOR U31851 ( .A(n34457), .B(n34455), .Z(n34456) );
  XOR U31852 ( .A(n34458), .B(n34459), .Z(n31612) );
  NOR U31853 ( .A(n34460), .B(n34458), .Z(n34459) );
  XOR U31854 ( .A(n34461), .B(n34462), .Z(n31615) );
  NOR U31855 ( .A(n34463), .B(n34461), .Z(n34462) );
  XOR U31856 ( .A(n34464), .B(n34465), .Z(n31618) );
  NOR U31857 ( .A(n34466), .B(n34464), .Z(n34465) );
  XOR U31858 ( .A(n34467), .B(n34468), .Z(n31621) );
  NOR U31859 ( .A(n34469), .B(n34467), .Z(n34468) );
  XOR U31860 ( .A(n34470), .B(n34471), .Z(n31624) );
  NOR U31861 ( .A(n34472), .B(n34470), .Z(n34471) );
  XOR U31862 ( .A(n34473), .B(n34474), .Z(n31627) );
  NOR U31863 ( .A(n34475), .B(n34473), .Z(n34474) );
  XOR U31864 ( .A(n34476), .B(n34477), .Z(n31630) );
  NOR U31865 ( .A(n34478), .B(n34476), .Z(n34477) );
  XOR U31866 ( .A(n34479), .B(n34480), .Z(n31633) );
  NOR U31867 ( .A(n34481), .B(n34479), .Z(n34480) );
  XOR U31868 ( .A(n34482), .B(n34483), .Z(n31636) );
  NOR U31869 ( .A(n34484), .B(n34482), .Z(n34483) );
  XOR U31870 ( .A(n34485), .B(n34486), .Z(n31639) );
  NOR U31871 ( .A(n34487), .B(n34485), .Z(n34486) );
  XOR U31872 ( .A(n34488), .B(n34489), .Z(n31642) );
  NOR U31873 ( .A(n34490), .B(n34488), .Z(n34489) );
  XOR U31874 ( .A(n34491), .B(n34492), .Z(n31645) );
  NOR U31875 ( .A(n34493), .B(n34491), .Z(n34492) );
  XOR U31876 ( .A(n34494), .B(n34495), .Z(n31648) );
  NOR U31877 ( .A(n34496), .B(n34494), .Z(n34495) );
  XOR U31878 ( .A(n34497), .B(n34498), .Z(n31651) );
  NOR U31879 ( .A(n34499), .B(n34497), .Z(n34498) );
  XOR U31880 ( .A(n34500), .B(n34501), .Z(n31654) );
  NOR U31881 ( .A(n34502), .B(n34500), .Z(n34501) );
  XOR U31882 ( .A(n34503), .B(n34504), .Z(n31657) );
  NOR U31883 ( .A(n34505), .B(n34503), .Z(n34504) );
  XOR U31884 ( .A(n34506), .B(n34507), .Z(n31660) );
  NOR U31885 ( .A(n34508), .B(n34506), .Z(n34507) );
  XOR U31886 ( .A(n34509), .B(n34510), .Z(n31663) );
  NOR U31887 ( .A(n34511), .B(n34509), .Z(n34510) );
  XOR U31888 ( .A(n34512), .B(n34513), .Z(n31666) );
  NOR U31889 ( .A(n34514), .B(n34512), .Z(n34513) );
  XOR U31890 ( .A(n34515), .B(n34516), .Z(n31669) );
  NOR U31891 ( .A(n34517), .B(n34515), .Z(n34516) );
  XOR U31892 ( .A(n34518), .B(n34519), .Z(n31672) );
  NOR U31893 ( .A(n34520), .B(n34518), .Z(n34519) );
  XOR U31894 ( .A(n34521), .B(n34522), .Z(n31675) );
  NOR U31895 ( .A(n34523), .B(n34521), .Z(n34522) );
  XOR U31896 ( .A(n34524), .B(n34525), .Z(n31678) );
  NOR U31897 ( .A(n34526), .B(n34524), .Z(n34525) );
  XOR U31898 ( .A(n34527), .B(n34528), .Z(n31681) );
  NOR U31899 ( .A(n34529), .B(n34527), .Z(n34528) );
  XOR U31900 ( .A(n34530), .B(n34531), .Z(n31684) );
  NOR U31901 ( .A(n34532), .B(n34530), .Z(n34531) );
  XOR U31902 ( .A(n34533), .B(n34534), .Z(n31687) );
  NOR U31903 ( .A(n34535), .B(n34533), .Z(n34534) );
  XOR U31904 ( .A(n34536), .B(n34537), .Z(n31690) );
  NOR U31905 ( .A(n34538), .B(n34536), .Z(n34537) );
  XOR U31906 ( .A(n34539), .B(n34540), .Z(n31693) );
  NOR U31907 ( .A(n34541), .B(n34539), .Z(n34540) );
  XOR U31908 ( .A(n34542), .B(n34543), .Z(n31696) );
  NOR U31909 ( .A(n34544), .B(n34542), .Z(n34543) );
  XOR U31910 ( .A(n34545), .B(n34546), .Z(n31699) );
  NOR U31911 ( .A(n34547), .B(n34545), .Z(n34546) );
  XOR U31912 ( .A(n34548), .B(n34549), .Z(n31702) );
  NOR U31913 ( .A(n34550), .B(n34548), .Z(n34549) );
  XOR U31914 ( .A(n34551), .B(n34552), .Z(n31705) );
  NOR U31915 ( .A(n34553), .B(n34551), .Z(n34552) );
  XOR U31916 ( .A(n34554), .B(n34555), .Z(n31708) );
  NOR U31917 ( .A(n34556), .B(n34554), .Z(n34555) );
  XOR U31918 ( .A(n34557), .B(n34558), .Z(n31711) );
  NOR U31919 ( .A(n34559), .B(n34557), .Z(n34558) );
  XOR U31920 ( .A(n34560), .B(n34561), .Z(n31714) );
  NOR U31921 ( .A(n34562), .B(n34560), .Z(n34561) );
  XOR U31922 ( .A(n34563), .B(n34564), .Z(n31717) );
  NOR U31923 ( .A(n34565), .B(n34563), .Z(n34564) );
  XOR U31924 ( .A(n34566), .B(n34567), .Z(n31720) );
  NOR U31925 ( .A(n34568), .B(n34566), .Z(n34567) );
  XOR U31926 ( .A(n34569), .B(n34570), .Z(n31723) );
  NOR U31927 ( .A(n34571), .B(n34569), .Z(n34570) );
  XOR U31928 ( .A(n34572), .B(n34573), .Z(n31726) );
  NOR U31929 ( .A(n34574), .B(n34572), .Z(n34573) );
  XOR U31930 ( .A(n34575), .B(n34576), .Z(n31729) );
  NOR U31931 ( .A(n34577), .B(n34575), .Z(n34576) );
  XOR U31932 ( .A(n34578), .B(n34579), .Z(n31732) );
  NOR U31933 ( .A(n34580), .B(n34578), .Z(n34579) );
  XOR U31934 ( .A(n34581), .B(n34582), .Z(n31735) );
  NOR U31935 ( .A(n34583), .B(n34581), .Z(n34582) );
  XOR U31936 ( .A(n34584), .B(n34585), .Z(n31738) );
  NOR U31937 ( .A(n34586), .B(n34584), .Z(n34585) );
  XOR U31938 ( .A(n34587), .B(n34588), .Z(n31741) );
  NOR U31939 ( .A(n34589), .B(n34587), .Z(n34588) );
  XOR U31940 ( .A(n34590), .B(n34591), .Z(n31744) );
  NOR U31941 ( .A(n34592), .B(n34590), .Z(n34591) );
  XOR U31942 ( .A(n34593), .B(n34594), .Z(n31747) );
  NOR U31943 ( .A(n34595), .B(n34593), .Z(n34594) );
  XOR U31944 ( .A(n34596), .B(n34597), .Z(n31750) );
  NOR U31945 ( .A(n34598), .B(n34596), .Z(n34597) );
  XOR U31946 ( .A(n34599), .B(n34600), .Z(n31753) );
  NOR U31947 ( .A(n34601), .B(n34599), .Z(n34600) );
  XOR U31948 ( .A(n34602), .B(n34603), .Z(n31756) );
  NOR U31949 ( .A(n34604), .B(n34602), .Z(n34603) );
  XOR U31950 ( .A(n34605), .B(n34606), .Z(n31759) );
  NOR U31951 ( .A(n34607), .B(n34605), .Z(n34606) );
  XOR U31952 ( .A(n34608), .B(n34609), .Z(n31762) );
  NOR U31953 ( .A(n34610), .B(n34608), .Z(n34609) );
  XOR U31954 ( .A(n34611), .B(n34612), .Z(n31765) );
  NOR U31955 ( .A(n34613), .B(n34611), .Z(n34612) );
  XOR U31956 ( .A(n34614), .B(n34615), .Z(n31768) );
  NOR U31957 ( .A(n34616), .B(n34614), .Z(n34615) );
  XOR U31958 ( .A(n34617), .B(n34618), .Z(n31771) );
  NOR U31959 ( .A(n34619), .B(n34617), .Z(n34618) );
  XOR U31960 ( .A(n34620), .B(n34621), .Z(n31774) );
  NOR U31961 ( .A(n34622), .B(n34620), .Z(n34621) );
  XOR U31962 ( .A(n34623), .B(n34624), .Z(n31777) );
  NOR U31963 ( .A(n34625), .B(n34623), .Z(n34624) );
  XOR U31964 ( .A(n34626), .B(n34627), .Z(n31780) );
  NOR U31965 ( .A(n34628), .B(n34626), .Z(n34627) );
  XOR U31966 ( .A(n34629), .B(n34630), .Z(n31783) );
  NOR U31967 ( .A(n34631), .B(n34629), .Z(n34630) );
  XOR U31968 ( .A(n34632), .B(n34633), .Z(n31786) );
  NOR U31969 ( .A(n34634), .B(n34632), .Z(n34633) );
  XOR U31970 ( .A(n34635), .B(n34636), .Z(n31789) );
  NOR U31971 ( .A(n34637), .B(n34635), .Z(n34636) );
  XOR U31972 ( .A(n34638), .B(n34639), .Z(n31792) );
  NOR U31973 ( .A(n34640), .B(n34638), .Z(n34639) );
  XOR U31974 ( .A(n34641), .B(n34642), .Z(n31795) );
  NOR U31975 ( .A(n34643), .B(n34641), .Z(n34642) );
  XOR U31976 ( .A(n34644), .B(n34645), .Z(n31798) );
  NOR U31977 ( .A(n34646), .B(n34644), .Z(n34645) );
  XOR U31978 ( .A(n34647), .B(n34648), .Z(n31801) );
  NOR U31979 ( .A(n34649), .B(n34647), .Z(n34648) );
  XOR U31980 ( .A(n34650), .B(n34651), .Z(n31804) );
  NOR U31981 ( .A(n34652), .B(n34650), .Z(n34651) );
  XOR U31982 ( .A(n34653), .B(n34654), .Z(n31807) );
  NOR U31983 ( .A(n34655), .B(n34653), .Z(n34654) );
  XOR U31984 ( .A(n34656), .B(n34657), .Z(n31810) );
  NOR U31985 ( .A(n34658), .B(n34656), .Z(n34657) );
  XOR U31986 ( .A(n34659), .B(n34660), .Z(n31813) );
  NOR U31987 ( .A(n34661), .B(n34659), .Z(n34660) );
  XOR U31988 ( .A(n34662), .B(n34663), .Z(n31816) );
  NOR U31989 ( .A(n34664), .B(n34662), .Z(n34663) );
  XOR U31990 ( .A(n34665), .B(n34666), .Z(n31819) );
  NOR U31991 ( .A(n34667), .B(n34665), .Z(n34666) );
  XOR U31992 ( .A(n34668), .B(n34669), .Z(n31822) );
  NOR U31993 ( .A(n34670), .B(n34668), .Z(n34669) );
  XOR U31994 ( .A(n34671), .B(n34672), .Z(n31825) );
  NOR U31995 ( .A(n34673), .B(n34671), .Z(n34672) );
  XOR U31996 ( .A(n34674), .B(n34675), .Z(n31828) );
  NOR U31997 ( .A(n34676), .B(n34674), .Z(n34675) );
  XOR U31998 ( .A(n34677), .B(n34678), .Z(n31831) );
  NOR U31999 ( .A(n34679), .B(n34677), .Z(n34678) );
  XOR U32000 ( .A(n34680), .B(n34681), .Z(n31834) );
  NOR U32001 ( .A(n34682), .B(n34680), .Z(n34681) );
  XOR U32002 ( .A(n34683), .B(n34684), .Z(n31837) );
  NOR U32003 ( .A(n34685), .B(n34683), .Z(n34684) );
  XOR U32004 ( .A(n34686), .B(n34687), .Z(n31840) );
  NOR U32005 ( .A(n34688), .B(n34686), .Z(n34687) );
  XOR U32006 ( .A(n34689), .B(n34690), .Z(n31843) );
  NOR U32007 ( .A(n34691), .B(n34689), .Z(n34690) );
  XOR U32008 ( .A(n34692), .B(n34693), .Z(n31846) );
  NOR U32009 ( .A(n34694), .B(n34692), .Z(n34693) );
  XOR U32010 ( .A(n34695), .B(n34696), .Z(n31849) );
  NOR U32011 ( .A(n34697), .B(n34695), .Z(n34696) );
  XOR U32012 ( .A(n34698), .B(n34699), .Z(n31852) );
  NOR U32013 ( .A(n34700), .B(n34698), .Z(n34699) );
  XOR U32014 ( .A(n34701), .B(n34702), .Z(n31855) );
  NOR U32015 ( .A(n34703), .B(n34701), .Z(n34702) );
  XOR U32016 ( .A(n34704), .B(n34705), .Z(n31858) );
  NOR U32017 ( .A(n34706), .B(n34704), .Z(n34705) );
  XOR U32018 ( .A(n34707), .B(n34708), .Z(n31861) );
  NOR U32019 ( .A(n34709), .B(n34707), .Z(n34708) );
  XOR U32020 ( .A(n34710), .B(n34711), .Z(n31864) );
  NOR U32021 ( .A(n34712), .B(n34710), .Z(n34711) );
  XOR U32022 ( .A(n34713), .B(n34714), .Z(n31867) );
  NOR U32023 ( .A(n34715), .B(n34713), .Z(n34714) );
  XOR U32024 ( .A(n34716), .B(n34717), .Z(n31870) );
  NOR U32025 ( .A(n34718), .B(n34716), .Z(n34717) );
  XOR U32026 ( .A(n34719), .B(n34720), .Z(n31873) );
  NOR U32027 ( .A(n34721), .B(n34719), .Z(n34720) );
  XOR U32028 ( .A(n34722), .B(n34723), .Z(n31876) );
  NOR U32029 ( .A(n34724), .B(n34722), .Z(n34723) );
  XOR U32030 ( .A(n34725), .B(n34726), .Z(n31879) );
  NOR U32031 ( .A(n34727), .B(n34725), .Z(n34726) );
  XOR U32032 ( .A(n34728), .B(n34729), .Z(n31882) );
  NOR U32033 ( .A(n34730), .B(n34728), .Z(n34729) );
  XOR U32034 ( .A(n34731), .B(n34732), .Z(n31885) );
  NOR U32035 ( .A(n34733), .B(n34731), .Z(n34732) );
  XOR U32036 ( .A(n34734), .B(n34735), .Z(n31888) );
  NOR U32037 ( .A(n34736), .B(n34734), .Z(n34735) );
  XOR U32038 ( .A(n34737), .B(n34738), .Z(n31891) );
  NOR U32039 ( .A(n34739), .B(n34737), .Z(n34738) );
  XOR U32040 ( .A(n34740), .B(n34741), .Z(n31894) );
  NOR U32041 ( .A(n34742), .B(n34740), .Z(n34741) );
  XOR U32042 ( .A(n34743), .B(n34744), .Z(n31897) );
  NOR U32043 ( .A(n34745), .B(n34743), .Z(n34744) );
  XOR U32044 ( .A(n34746), .B(n34747), .Z(n31900) );
  NOR U32045 ( .A(n34748), .B(n34746), .Z(n34747) );
  XOR U32046 ( .A(n34749), .B(n34750), .Z(n31903) );
  NOR U32047 ( .A(n34751), .B(n34749), .Z(n34750) );
  XOR U32048 ( .A(n34752), .B(n34753), .Z(n31906) );
  NOR U32049 ( .A(n34754), .B(n34752), .Z(n34753) );
  XOR U32050 ( .A(n34755), .B(n34756), .Z(n31909) );
  NOR U32051 ( .A(n34757), .B(n34755), .Z(n34756) );
  XOR U32052 ( .A(n34758), .B(n34759), .Z(n31912) );
  NOR U32053 ( .A(n34760), .B(n34758), .Z(n34759) );
  XOR U32054 ( .A(n34761), .B(n34762), .Z(n31915) );
  NOR U32055 ( .A(n34763), .B(n34761), .Z(n34762) );
  XOR U32056 ( .A(n34764), .B(n34765), .Z(n31918) );
  NOR U32057 ( .A(n34766), .B(n34764), .Z(n34765) );
  XOR U32058 ( .A(n34767), .B(n34768), .Z(n31921) );
  NOR U32059 ( .A(n34769), .B(n34767), .Z(n34768) );
  XOR U32060 ( .A(n34770), .B(n34771), .Z(n31924) );
  NOR U32061 ( .A(n34772), .B(n34770), .Z(n34771) );
  XOR U32062 ( .A(n34773), .B(n34774), .Z(n31927) );
  NOR U32063 ( .A(n34775), .B(n34773), .Z(n34774) );
  XOR U32064 ( .A(n34776), .B(n34777), .Z(n31930) );
  NOR U32065 ( .A(n34778), .B(n34776), .Z(n34777) );
  XOR U32066 ( .A(n34779), .B(n34780), .Z(n31933) );
  NOR U32067 ( .A(n34781), .B(n34779), .Z(n34780) );
  XOR U32068 ( .A(n34782), .B(n34783), .Z(n31936) );
  NOR U32069 ( .A(n34784), .B(n34782), .Z(n34783) );
  XOR U32070 ( .A(n34785), .B(n34786), .Z(n31939) );
  NOR U32071 ( .A(n34787), .B(n34785), .Z(n34786) );
  XOR U32072 ( .A(n34788), .B(n34789), .Z(n31942) );
  NOR U32073 ( .A(n34790), .B(n34788), .Z(n34789) );
  XOR U32074 ( .A(n34791), .B(n34792), .Z(n31945) );
  NOR U32075 ( .A(n34793), .B(n34791), .Z(n34792) );
  XOR U32076 ( .A(n34794), .B(n34795), .Z(n31948) );
  NOR U32077 ( .A(n34796), .B(n34794), .Z(n34795) );
  XOR U32078 ( .A(n34797), .B(n34798), .Z(n31951) );
  NOR U32079 ( .A(n34799), .B(n34797), .Z(n34798) );
  XOR U32080 ( .A(n34800), .B(n34801), .Z(n31954) );
  NOR U32081 ( .A(n34802), .B(n34800), .Z(n34801) );
  XOR U32082 ( .A(n34803), .B(n34804), .Z(n31957) );
  NOR U32083 ( .A(n34805), .B(n34803), .Z(n34804) );
  XOR U32084 ( .A(n34806), .B(n34807), .Z(n31960) );
  NOR U32085 ( .A(n34808), .B(n34806), .Z(n34807) );
  XOR U32086 ( .A(n34809), .B(n34810), .Z(n31963) );
  NOR U32087 ( .A(n34811), .B(n34809), .Z(n34810) );
  XOR U32088 ( .A(n34812), .B(n34813), .Z(n31966) );
  NOR U32089 ( .A(n34814), .B(n34812), .Z(n34813) );
  XOR U32090 ( .A(n34815), .B(n34816), .Z(n31969) );
  NOR U32091 ( .A(n34817), .B(n34815), .Z(n34816) );
  XOR U32092 ( .A(n34818), .B(n34819), .Z(n31972) );
  NOR U32093 ( .A(n34820), .B(n34818), .Z(n34819) );
  XOR U32094 ( .A(n34821), .B(n34822), .Z(n31975) );
  NOR U32095 ( .A(n34823), .B(n34821), .Z(n34822) );
  XOR U32096 ( .A(n34824), .B(n34825), .Z(n31978) );
  NOR U32097 ( .A(n34826), .B(n34824), .Z(n34825) );
  XOR U32098 ( .A(n34827), .B(n34828), .Z(n31981) );
  NOR U32099 ( .A(n34829), .B(n34827), .Z(n34828) );
  XOR U32100 ( .A(n34830), .B(n34831), .Z(n31984) );
  NOR U32101 ( .A(n34832), .B(n34830), .Z(n34831) );
  XOR U32102 ( .A(n34833), .B(n34834), .Z(n31987) );
  NOR U32103 ( .A(n34835), .B(n34833), .Z(n34834) );
  XOR U32104 ( .A(n34836), .B(n34837), .Z(n31990) );
  NOR U32105 ( .A(n34838), .B(n34836), .Z(n34837) );
  XOR U32106 ( .A(n34839), .B(n34840), .Z(n31993) );
  NOR U32107 ( .A(n34841), .B(n34839), .Z(n34840) );
  XOR U32108 ( .A(n34842), .B(n34843), .Z(n31996) );
  NOR U32109 ( .A(n34844), .B(n34842), .Z(n34843) );
  XOR U32110 ( .A(n34845), .B(n34846), .Z(n31999) );
  NOR U32111 ( .A(n34847), .B(n34845), .Z(n34846) );
  XOR U32112 ( .A(n34848), .B(n34849), .Z(n32002) );
  NOR U32113 ( .A(n34850), .B(n34848), .Z(n34849) );
  XOR U32114 ( .A(n34851), .B(n34852), .Z(n32005) );
  NOR U32115 ( .A(n34853), .B(n34851), .Z(n34852) );
  XOR U32116 ( .A(n34854), .B(n34855), .Z(n32008) );
  NOR U32117 ( .A(n34856), .B(n34854), .Z(n34855) );
  XOR U32118 ( .A(n34857), .B(n34858), .Z(n32011) );
  NOR U32119 ( .A(n34859), .B(n34857), .Z(n34858) );
  XOR U32120 ( .A(n34860), .B(n34861), .Z(n32014) );
  NOR U32121 ( .A(n34862), .B(n34860), .Z(n34861) );
  XOR U32122 ( .A(n34863), .B(n34864), .Z(n32017) );
  NOR U32123 ( .A(n34865), .B(n34863), .Z(n34864) );
  XOR U32124 ( .A(n34866), .B(n34867), .Z(n32020) );
  NOR U32125 ( .A(n34868), .B(n34866), .Z(n34867) );
  XOR U32126 ( .A(n34869), .B(n34870), .Z(n32023) );
  NOR U32127 ( .A(n34871), .B(n34869), .Z(n34870) );
  XOR U32128 ( .A(n34872), .B(n34873), .Z(n32026) );
  NOR U32129 ( .A(n34874), .B(n34872), .Z(n34873) );
  XOR U32130 ( .A(n34875), .B(n34876), .Z(n32029) );
  NOR U32131 ( .A(n34877), .B(n34875), .Z(n34876) );
  XOR U32132 ( .A(n34878), .B(n34879), .Z(n32032) );
  NOR U32133 ( .A(n34880), .B(n34878), .Z(n34879) );
  XOR U32134 ( .A(n34881), .B(n34882), .Z(n32035) );
  NOR U32135 ( .A(n34883), .B(n34881), .Z(n34882) );
  XOR U32136 ( .A(n34884), .B(n34885), .Z(n32038) );
  NOR U32137 ( .A(n34886), .B(n34884), .Z(n34885) );
  XOR U32138 ( .A(n34887), .B(n34888), .Z(n32041) );
  NOR U32139 ( .A(n34889), .B(n34887), .Z(n34888) );
  XOR U32140 ( .A(n34890), .B(n34891), .Z(n32044) );
  NOR U32141 ( .A(n34892), .B(n34890), .Z(n34891) );
  XOR U32142 ( .A(n34893), .B(n34894), .Z(n32047) );
  NOR U32143 ( .A(n34895), .B(n34893), .Z(n34894) );
  XOR U32144 ( .A(n34896), .B(n34897), .Z(n32050) );
  NOR U32145 ( .A(n34898), .B(n34896), .Z(n34897) );
  XOR U32146 ( .A(n34899), .B(n34900), .Z(n32053) );
  NOR U32147 ( .A(n34901), .B(n34899), .Z(n34900) );
  XOR U32148 ( .A(n34902), .B(n34903), .Z(n32056) );
  NOR U32149 ( .A(n34904), .B(n34902), .Z(n34903) );
  XOR U32150 ( .A(n34905), .B(n34906), .Z(n32059) );
  NOR U32151 ( .A(n34907), .B(n34905), .Z(n34906) );
  XOR U32152 ( .A(n34908), .B(n34909), .Z(n32062) );
  NOR U32153 ( .A(n34910), .B(n34908), .Z(n34909) );
  XOR U32154 ( .A(n34911), .B(n34912), .Z(n32065) );
  NOR U32155 ( .A(n34913), .B(n34911), .Z(n34912) );
  XOR U32156 ( .A(n34914), .B(n34915), .Z(n32068) );
  NOR U32157 ( .A(n34916), .B(n34914), .Z(n34915) );
  XOR U32158 ( .A(n34917), .B(n34918), .Z(n32071) );
  NOR U32159 ( .A(n34919), .B(n34917), .Z(n34918) );
  XOR U32160 ( .A(n34920), .B(n34921), .Z(n32074) );
  NOR U32161 ( .A(n34922), .B(n34920), .Z(n34921) );
  XOR U32162 ( .A(n34923), .B(n34924), .Z(n32077) );
  NOR U32163 ( .A(n34925), .B(n34923), .Z(n34924) );
  XOR U32164 ( .A(n34926), .B(n34927), .Z(n32080) );
  NOR U32165 ( .A(n34928), .B(n34926), .Z(n34927) );
  XOR U32166 ( .A(n34929), .B(n34930), .Z(n32083) );
  NOR U32167 ( .A(n34931), .B(n34929), .Z(n34930) );
  XOR U32168 ( .A(n34932), .B(n34933), .Z(n32086) );
  NOR U32169 ( .A(n34934), .B(n34932), .Z(n34933) );
  XOR U32170 ( .A(n34935), .B(n34936), .Z(n32089) );
  NOR U32171 ( .A(n34937), .B(n34935), .Z(n34936) );
  XOR U32172 ( .A(n34938), .B(n34939), .Z(n32092) );
  NOR U32173 ( .A(n34940), .B(n34938), .Z(n34939) );
  XOR U32174 ( .A(n34941), .B(n34942), .Z(n32095) );
  NOR U32175 ( .A(n34943), .B(n34941), .Z(n34942) );
  XOR U32176 ( .A(n34944), .B(n34945), .Z(n32098) );
  NOR U32177 ( .A(n34946), .B(n34944), .Z(n34945) );
  XOR U32178 ( .A(n34947), .B(n34948), .Z(n32101) );
  NOR U32179 ( .A(n34949), .B(n34947), .Z(n34948) );
  XOR U32180 ( .A(n34950), .B(n34951), .Z(n32104) );
  NOR U32181 ( .A(n34952), .B(n34950), .Z(n34951) );
  XOR U32182 ( .A(n34953), .B(n34954), .Z(n32107) );
  NOR U32183 ( .A(n34955), .B(n34953), .Z(n34954) );
  XOR U32184 ( .A(n34956), .B(n34957), .Z(n32110) );
  NOR U32185 ( .A(n34958), .B(n34956), .Z(n34957) );
  XOR U32186 ( .A(n34959), .B(n34960), .Z(n32113) );
  NOR U32187 ( .A(n34961), .B(n34959), .Z(n34960) );
  XOR U32188 ( .A(n34962), .B(n34963), .Z(n32116) );
  NOR U32189 ( .A(n34964), .B(n34962), .Z(n34963) );
  XOR U32190 ( .A(n34965), .B(n34966), .Z(n32119) );
  NOR U32191 ( .A(n34967), .B(n34965), .Z(n34966) );
  XOR U32192 ( .A(n34968), .B(n34969), .Z(n32122) );
  NOR U32193 ( .A(n34970), .B(n34968), .Z(n34969) );
  XOR U32194 ( .A(n34971), .B(n34972), .Z(n32125) );
  NOR U32195 ( .A(n34973), .B(n34971), .Z(n34972) );
  XOR U32196 ( .A(n34974), .B(n34975), .Z(n32128) );
  NOR U32197 ( .A(n34976), .B(n34974), .Z(n34975) );
  XOR U32198 ( .A(n34977), .B(n34978), .Z(n32131) );
  NOR U32199 ( .A(n34979), .B(n34977), .Z(n34978) );
  XOR U32200 ( .A(n34980), .B(n34981), .Z(n32134) );
  NOR U32201 ( .A(n34982), .B(n34980), .Z(n34981) );
  XOR U32202 ( .A(n34983), .B(n34984), .Z(n32137) );
  NOR U32203 ( .A(n34985), .B(n34983), .Z(n34984) );
  XOR U32204 ( .A(n34986), .B(n34987), .Z(n32140) );
  NOR U32205 ( .A(n34988), .B(n34986), .Z(n34987) );
  XOR U32206 ( .A(n34989), .B(n34990), .Z(n32143) );
  NOR U32207 ( .A(n34991), .B(n34989), .Z(n34990) );
  XOR U32208 ( .A(n34992), .B(n34993), .Z(n32146) );
  NOR U32209 ( .A(n34994), .B(n34992), .Z(n34993) );
  XOR U32210 ( .A(n34995), .B(n34996), .Z(n32149) );
  NOR U32211 ( .A(n34997), .B(n34995), .Z(n34996) );
  XOR U32212 ( .A(n34998), .B(n34999), .Z(n32152) );
  NOR U32213 ( .A(n35000), .B(n34998), .Z(n34999) );
  XOR U32214 ( .A(n35001), .B(n35002), .Z(n32155) );
  NOR U32215 ( .A(n35003), .B(n35001), .Z(n35002) );
  XOR U32216 ( .A(n35004), .B(n35005), .Z(n32158) );
  NOR U32217 ( .A(n35006), .B(n35004), .Z(n35005) );
  XOR U32218 ( .A(n35007), .B(n35008), .Z(n32161) );
  NOR U32219 ( .A(n35009), .B(n35007), .Z(n35008) );
  XOR U32220 ( .A(n35010), .B(n35011), .Z(n32164) );
  NOR U32221 ( .A(n35012), .B(n35010), .Z(n35011) );
  XOR U32222 ( .A(n35013), .B(n35014), .Z(n32167) );
  NOR U32223 ( .A(n35015), .B(n35013), .Z(n35014) );
  XOR U32224 ( .A(n35016), .B(n35017), .Z(n32170) );
  NOR U32225 ( .A(n35018), .B(n35016), .Z(n35017) );
  XOR U32226 ( .A(n35019), .B(n35020), .Z(n32173) );
  NOR U32227 ( .A(n35021), .B(n35019), .Z(n35020) );
  XOR U32228 ( .A(n35022), .B(n35023), .Z(n32176) );
  NOR U32229 ( .A(n35024), .B(n35022), .Z(n35023) );
  XOR U32230 ( .A(n35025), .B(n35026), .Z(n32179) );
  NOR U32231 ( .A(n35027), .B(n35025), .Z(n35026) );
  XOR U32232 ( .A(n35028), .B(n35029), .Z(n32182) );
  NOR U32233 ( .A(n35030), .B(n35028), .Z(n35029) );
  XOR U32234 ( .A(n35031), .B(n35032), .Z(n32185) );
  NOR U32235 ( .A(n35033), .B(n35031), .Z(n35032) );
  XOR U32236 ( .A(n35034), .B(n35035), .Z(n32188) );
  NOR U32237 ( .A(n35036), .B(n35034), .Z(n35035) );
  XOR U32238 ( .A(n35037), .B(n35038), .Z(n32191) );
  NOR U32239 ( .A(n35039), .B(n35037), .Z(n35038) );
  XOR U32240 ( .A(n35040), .B(n35041), .Z(n32194) );
  NOR U32241 ( .A(n35042), .B(n35040), .Z(n35041) );
  XOR U32242 ( .A(n35043), .B(n35044), .Z(n32197) );
  NOR U32243 ( .A(n35045), .B(n35043), .Z(n35044) );
  XOR U32244 ( .A(n35046), .B(n35047), .Z(n32200) );
  NOR U32245 ( .A(n35048), .B(n35046), .Z(n35047) );
  XOR U32246 ( .A(n35049), .B(n35050), .Z(n32203) );
  NOR U32247 ( .A(n35051), .B(n35049), .Z(n35050) );
  XOR U32248 ( .A(n35052), .B(n35053), .Z(n32206) );
  NOR U32249 ( .A(n35054), .B(n35052), .Z(n35053) );
  XOR U32250 ( .A(n35055), .B(n35056), .Z(n32209) );
  NOR U32251 ( .A(n35057), .B(n35055), .Z(n35056) );
  XOR U32252 ( .A(n35058), .B(n35059), .Z(n32212) );
  NOR U32253 ( .A(n35060), .B(n35058), .Z(n35059) );
  XOR U32254 ( .A(n35061), .B(n35062), .Z(n32215) );
  NOR U32255 ( .A(n35063), .B(n35061), .Z(n35062) );
  XOR U32256 ( .A(n35064), .B(n35065), .Z(n32218) );
  NOR U32257 ( .A(n35066), .B(n35064), .Z(n35065) );
  XOR U32258 ( .A(n35067), .B(n35068), .Z(n32221) );
  NOR U32259 ( .A(n35069), .B(n35067), .Z(n35068) );
  XOR U32260 ( .A(n35070), .B(n35071), .Z(n32224) );
  NOR U32261 ( .A(n35072), .B(n35070), .Z(n35071) );
  XOR U32262 ( .A(n35073), .B(n35074), .Z(n32227) );
  NOR U32263 ( .A(n35075), .B(n35073), .Z(n35074) );
  XOR U32264 ( .A(n35076), .B(n35077), .Z(n32230) );
  NOR U32265 ( .A(n35078), .B(n35076), .Z(n35077) );
  XOR U32266 ( .A(n35079), .B(n35080), .Z(n32233) );
  NOR U32267 ( .A(n35081), .B(n35079), .Z(n35080) );
  XOR U32268 ( .A(n35082), .B(n35083), .Z(n32236) );
  NOR U32269 ( .A(n35084), .B(n35082), .Z(n35083) );
  XOR U32270 ( .A(n35085), .B(n35086), .Z(n32239) );
  NOR U32271 ( .A(n35087), .B(n35085), .Z(n35086) );
  XOR U32272 ( .A(n35088), .B(n35089), .Z(n32242) );
  NOR U32273 ( .A(n35090), .B(n35088), .Z(n35089) );
  XOR U32274 ( .A(n35091), .B(n35092), .Z(n32245) );
  NOR U32275 ( .A(n35093), .B(n35091), .Z(n35092) );
  XOR U32276 ( .A(n35094), .B(n35095), .Z(n32248) );
  NOR U32277 ( .A(n35096), .B(n35094), .Z(n35095) );
  XOR U32278 ( .A(n35097), .B(n35098), .Z(n32251) );
  NOR U32279 ( .A(n35099), .B(n35097), .Z(n35098) );
  XOR U32280 ( .A(n35100), .B(n35101), .Z(n32254) );
  NOR U32281 ( .A(n35102), .B(n35100), .Z(n35101) );
  XOR U32282 ( .A(n35103), .B(n35104), .Z(n32257) );
  NOR U32283 ( .A(n35105), .B(n35103), .Z(n35104) );
  XOR U32284 ( .A(n35106), .B(n35107), .Z(n32260) );
  NOR U32285 ( .A(n35108), .B(n35106), .Z(n35107) );
  XOR U32286 ( .A(n35109), .B(n35110), .Z(n32263) );
  NOR U32287 ( .A(n35111), .B(n35109), .Z(n35110) );
  XOR U32288 ( .A(n35112), .B(n35113), .Z(n32266) );
  NOR U32289 ( .A(n35114), .B(n35112), .Z(n35113) );
  XOR U32290 ( .A(n35115), .B(n35116), .Z(n32269) );
  NOR U32291 ( .A(n35117), .B(n35115), .Z(n35116) );
  XOR U32292 ( .A(n35118), .B(n35119), .Z(n32272) );
  NOR U32293 ( .A(n35120), .B(n35118), .Z(n35119) );
  XOR U32294 ( .A(n35121), .B(n35122), .Z(n32275) );
  NOR U32295 ( .A(n35123), .B(n35121), .Z(n35122) );
  XOR U32296 ( .A(n35124), .B(n35125), .Z(n32278) );
  NOR U32297 ( .A(n35126), .B(n35124), .Z(n35125) );
  XOR U32298 ( .A(n35127), .B(n35128), .Z(n32281) );
  NOR U32299 ( .A(n35129), .B(n35127), .Z(n35128) );
  XOR U32300 ( .A(n35130), .B(n35131), .Z(n32284) );
  NOR U32301 ( .A(n35132), .B(n35130), .Z(n35131) );
  XOR U32302 ( .A(n35133), .B(n35134), .Z(n32287) );
  NOR U32303 ( .A(n35135), .B(n35133), .Z(n35134) );
  XOR U32304 ( .A(n35136), .B(n35137), .Z(n32290) );
  NOR U32305 ( .A(n35138), .B(n35136), .Z(n35137) );
  XOR U32306 ( .A(n35139), .B(n35140), .Z(n32293) );
  NOR U32307 ( .A(n35141), .B(n35139), .Z(n35140) );
  XOR U32308 ( .A(n35142), .B(n35143), .Z(n32296) );
  NOR U32309 ( .A(n35144), .B(n35142), .Z(n35143) );
  XOR U32310 ( .A(n35145), .B(n35146), .Z(n32299) );
  NOR U32311 ( .A(n35147), .B(n35145), .Z(n35146) );
  XOR U32312 ( .A(n35148), .B(n35149), .Z(n32302) );
  NOR U32313 ( .A(n35150), .B(n35148), .Z(n35149) );
  XOR U32314 ( .A(n35151), .B(n35152), .Z(n32305) );
  NOR U32315 ( .A(n35153), .B(n35151), .Z(n35152) );
  XOR U32316 ( .A(n35154), .B(n35155), .Z(n32308) );
  NOR U32317 ( .A(n35156), .B(n35154), .Z(n35155) );
  XOR U32318 ( .A(n35157), .B(n35158), .Z(n32311) );
  NOR U32319 ( .A(n35159), .B(n35157), .Z(n35158) );
  XOR U32320 ( .A(n35160), .B(n35161), .Z(n32314) );
  NOR U32321 ( .A(n35162), .B(n35160), .Z(n35161) );
  XOR U32322 ( .A(n35163), .B(n35164), .Z(n32317) );
  NOR U32323 ( .A(n35165), .B(n35163), .Z(n35164) );
  XOR U32324 ( .A(n35166), .B(n35167), .Z(n32320) );
  NOR U32325 ( .A(n35168), .B(n35166), .Z(n35167) );
  XOR U32326 ( .A(n35169), .B(n35170), .Z(n32323) );
  NOR U32327 ( .A(n35171), .B(n35169), .Z(n35170) );
  XOR U32328 ( .A(n35172), .B(n35173), .Z(n32326) );
  NOR U32329 ( .A(n35174), .B(n35172), .Z(n35173) );
  XOR U32330 ( .A(n35175), .B(n35176), .Z(n32329) );
  NOR U32331 ( .A(n35177), .B(n35175), .Z(n35176) );
  XOR U32332 ( .A(n35178), .B(n35179), .Z(n32332) );
  NOR U32333 ( .A(n35180), .B(n35178), .Z(n35179) );
  XOR U32334 ( .A(n35181), .B(n35182), .Z(n32335) );
  NOR U32335 ( .A(n35183), .B(n35181), .Z(n35182) );
  XOR U32336 ( .A(n35184), .B(n35185), .Z(n32338) );
  NOR U32337 ( .A(n35186), .B(n35184), .Z(n35185) );
  XOR U32338 ( .A(n35187), .B(n35188), .Z(n32341) );
  NOR U32339 ( .A(n35189), .B(n35187), .Z(n35188) );
  XOR U32340 ( .A(n35190), .B(n35191), .Z(n32344) );
  NOR U32341 ( .A(n35192), .B(n35190), .Z(n35191) );
  XOR U32342 ( .A(n35193), .B(n35194), .Z(n32347) );
  NOR U32343 ( .A(n35195), .B(n35193), .Z(n35194) );
  XOR U32344 ( .A(n35196), .B(n35197), .Z(n32350) );
  NOR U32345 ( .A(n35198), .B(n35196), .Z(n35197) );
  XOR U32346 ( .A(n35199), .B(n35200), .Z(n32353) );
  NOR U32347 ( .A(n35201), .B(n35199), .Z(n35200) );
  XOR U32348 ( .A(n35202), .B(n35203), .Z(n32356) );
  NOR U32349 ( .A(n35204), .B(n35202), .Z(n35203) );
  XOR U32350 ( .A(n35205), .B(n35206), .Z(n32359) );
  NOR U32351 ( .A(n35207), .B(n35205), .Z(n35206) );
  XOR U32352 ( .A(n35208), .B(n35209), .Z(n32362) );
  NOR U32353 ( .A(n35210), .B(n35208), .Z(n35209) );
  XOR U32354 ( .A(n35211), .B(n35212), .Z(n32365) );
  NOR U32355 ( .A(n35213), .B(n35211), .Z(n35212) );
  XOR U32356 ( .A(n35214), .B(n35215), .Z(n32368) );
  NOR U32357 ( .A(n35216), .B(n35214), .Z(n35215) );
  XOR U32358 ( .A(n35217), .B(n35218), .Z(n32371) );
  NOR U32359 ( .A(n35219), .B(n35217), .Z(n35218) );
  XOR U32360 ( .A(n35220), .B(n35221), .Z(n32374) );
  NOR U32361 ( .A(n35222), .B(n35220), .Z(n35221) );
  XOR U32362 ( .A(n35223), .B(n35224), .Z(n32377) );
  NOR U32363 ( .A(n35225), .B(n35223), .Z(n35224) );
  XOR U32364 ( .A(n35226), .B(n35227), .Z(n32380) );
  NOR U32365 ( .A(n35228), .B(n35226), .Z(n35227) );
  XOR U32366 ( .A(n35229), .B(n35230), .Z(n32383) );
  NOR U32367 ( .A(n35231), .B(n35229), .Z(n35230) );
  XOR U32368 ( .A(n35232), .B(n35233), .Z(n32386) );
  NOR U32369 ( .A(n35234), .B(n35232), .Z(n35233) );
  XOR U32370 ( .A(n35235), .B(n35236), .Z(n32389) );
  NOR U32371 ( .A(n35237), .B(n35235), .Z(n35236) );
  XOR U32372 ( .A(n35238), .B(n35239), .Z(n32392) );
  NOR U32373 ( .A(n35240), .B(n35238), .Z(n35239) );
  XOR U32374 ( .A(n35241), .B(n35242), .Z(n32395) );
  NOR U32375 ( .A(n35243), .B(n35241), .Z(n35242) );
  XOR U32376 ( .A(n35244), .B(n35245), .Z(n32398) );
  NOR U32377 ( .A(n35246), .B(n35244), .Z(n35245) );
  XOR U32378 ( .A(n35247), .B(n35248), .Z(n32401) );
  NOR U32379 ( .A(n35249), .B(n35247), .Z(n35248) );
  XOR U32380 ( .A(n35250), .B(n35251), .Z(n32404) );
  NOR U32381 ( .A(n35252), .B(n35250), .Z(n35251) );
  XOR U32382 ( .A(n35253), .B(n35254), .Z(n32407) );
  NOR U32383 ( .A(n35255), .B(n35253), .Z(n35254) );
  XOR U32384 ( .A(n35256), .B(n35257), .Z(n32410) );
  NOR U32385 ( .A(n35258), .B(n35256), .Z(n35257) );
  XOR U32386 ( .A(n35259), .B(n35260), .Z(n32413) );
  NOR U32387 ( .A(n35261), .B(n35259), .Z(n35260) );
  XOR U32388 ( .A(n35262), .B(n35263), .Z(n32416) );
  NOR U32389 ( .A(n35264), .B(n35262), .Z(n35263) );
  XOR U32390 ( .A(n35265), .B(n35266), .Z(n32419) );
  NOR U32391 ( .A(n35267), .B(n35265), .Z(n35266) );
  XOR U32392 ( .A(n35268), .B(n35269), .Z(n32422) );
  NOR U32393 ( .A(n35270), .B(n35268), .Z(n35269) );
  XOR U32394 ( .A(n35271), .B(n35272), .Z(n32425) );
  NOR U32395 ( .A(n35273), .B(n35271), .Z(n35272) );
  XOR U32396 ( .A(n35274), .B(n35275), .Z(n32428) );
  NOR U32397 ( .A(n35276), .B(n35274), .Z(n35275) );
  XOR U32398 ( .A(n35277), .B(n35278), .Z(n32431) );
  NOR U32399 ( .A(n35279), .B(n35277), .Z(n35278) );
  XOR U32400 ( .A(n35280), .B(n35281), .Z(n32434) );
  NOR U32401 ( .A(n35282), .B(n35280), .Z(n35281) );
  XOR U32402 ( .A(n35283), .B(n35284), .Z(n32437) );
  NOR U32403 ( .A(n35285), .B(n35283), .Z(n35284) );
  XOR U32404 ( .A(n35286), .B(n35287), .Z(n32440) );
  NOR U32405 ( .A(n35288), .B(n35286), .Z(n35287) );
  XOR U32406 ( .A(n35289), .B(n35290), .Z(n32443) );
  NOR U32407 ( .A(n35291), .B(n35289), .Z(n35290) );
  XOR U32408 ( .A(n35292), .B(n35293), .Z(n32446) );
  NOR U32409 ( .A(n35294), .B(n35292), .Z(n35293) );
  XOR U32410 ( .A(n35295), .B(n35296), .Z(n32449) );
  NOR U32411 ( .A(n35297), .B(n35295), .Z(n35296) );
  XOR U32412 ( .A(n35298), .B(n35299), .Z(n32452) );
  NOR U32413 ( .A(n35300), .B(n35298), .Z(n35299) );
  XOR U32414 ( .A(n35301), .B(n35302), .Z(n32455) );
  NOR U32415 ( .A(n35303), .B(n35301), .Z(n35302) );
  XOR U32416 ( .A(n35304), .B(n35305), .Z(n32458) );
  NOR U32417 ( .A(n35306), .B(n35304), .Z(n35305) );
  XOR U32418 ( .A(n35307), .B(n35308), .Z(n32461) );
  NOR U32419 ( .A(n35309), .B(n35307), .Z(n35308) );
  XOR U32420 ( .A(n35310), .B(n35311), .Z(n32464) );
  NOR U32421 ( .A(n35312), .B(n35310), .Z(n35311) );
  XOR U32422 ( .A(n35313), .B(n35314), .Z(n32467) );
  NOR U32423 ( .A(n35315), .B(n35313), .Z(n35314) );
  XOR U32424 ( .A(n35316), .B(n35317), .Z(n32470) );
  NOR U32425 ( .A(n35318), .B(n35316), .Z(n35317) );
  XOR U32426 ( .A(n35319), .B(n35320), .Z(n32473) );
  NOR U32427 ( .A(n35321), .B(n35319), .Z(n35320) );
  XOR U32428 ( .A(n35322), .B(n35323), .Z(n32476) );
  NOR U32429 ( .A(n35324), .B(n35322), .Z(n35323) );
  XOR U32430 ( .A(n35325), .B(n35326), .Z(n32479) );
  NOR U32431 ( .A(n35327), .B(n35325), .Z(n35326) );
  XOR U32432 ( .A(n35328), .B(n35329), .Z(n32482) );
  NOR U32433 ( .A(n35330), .B(n35328), .Z(n35329) );
  XOR U32434 ( .A(n35331), .B(n35332), .Z(n32485) );
  NOR U32435 ( .A(n35333), .B(n35331), .Z(n35332) );
  XOR U32436 ( .A(n35334), .B(n35335), .Z(n32488) );
  NOR U32437 ( .A(n35336), .B(n35334), .Z(n35335) );
  XOR U32438 ( .A(n35337), .B(n35338), .Z(n32491) );
  NOR U32439 ( .A(n35339), .B(n35337), .Z(n35338) );
  XOR U32440 ( .A(n35340), .B(n35341), .Z(n32494) );
  NOR U32441 ( .A(n35342), .B(n35340), .Z(n35341) );
  XOR U32442 ( .A(n35343), .B(n35344), .Z(n32497) );
  NOR U32443 ( .A(n35345), .B(n35343), .Z(n35344) );
  XOR U32444 ( .A(n35346), .B(n35347), .Z(n32500) );
  NOR U32445 ( .A(n35348), .B(n35346), .Z(n35347) );
  XOR U32446 ( .A(n35349), .B(n35350), .Z(n32503) );
  NOR U32447 ( .A(n35351), .B(n35349), .Z(n35350) );
  XOR U32448 ( .A(n35352), .B(n35353), .Z(n32506) );
  NOR U32449 ( .A(n35354), .B(n35352), .Z(n35353) );
  XOR U32450 ( .A(n35355), .B(n35356), .Z(n32509) );
  NOR U32451 ( .A(n35357), .B(n35355), .Z(n35356) );
  XOR U32452 ( .A(n35358), .B(n35359), .Z(n32512) );
  NOR U32453 ( .A(n35360), .B(n35358), .Z(n35359) );
  XOR U32454 ( .A(n35361), .B(n35362), .Z(n32515) );
  NOR U32455 ( .A(n35363), .B(n35361), .Z(n35362) );
  XOR U32456 ( .A(n35364), .B(n35365), .Z(n32518) );
  NOR U32457 ( .A(n35366), .B(n35364), .Z(n35365) );
  XOR U32458 ( .A(n35367), .B(n35368), .Z(n32521) );
  NOR U32459 ( .A(n35369), .B(n35367), .Z(n35368) );
  XOR U32460 ( .A(n35370), .B(n35371), .Z(n32524) );
  NOR U32461 ( .A(n35372), .B(n35370), .Z(n35371) );
  XOR U32462 ( .A(n35373), .B(n35374), .Z(n32527) );
  NOR U32463 ( .A(n35375), .B(n35373), .Z(n35374) );
  XOR U32464 ( .A(n35376), .B(n35377), .Z(n32530) );
  NOR U32465 ( .A(n35378), .B(n35376), .Z(n35377) );
  XOR U32466 ( .A(n35379), .B(n35380), .Z(n32533) );
  NOR U32467 ( .A(n35381), .B(n35379), .Z(n35380) );
  XOR U32468 ( .A(n35382), .B(n35383), .Z(n32536) );
  NOR U32469 ( .A(n35384), .B(n35382), .Z(n35383) );
  XOR U32470 ( .A(n35385), .B(n35386), .Z(n32539) );
  NOR U32471 ( .A(n35387), .B(n35385), .Z(n35386) );
  XOR U32472 ( .A(n35388), .B(n35389), .Z(n32542) );
  NOR U32473 ( .A(n35390), .B(n35388), .Z(n35389) );
  XOR U32474 ( .A(n35391), .B(n35392), .Z(n32545) );
  NOR U32475 ( .A(n35393), .B(n35391), .Z(n35392) );
  XOR U32476 ( .A(n35394), .B(n35395), .Z(n32548) );
  NOR U32477 ( .A(n35396), .B(n35394), .Z(n35395) );
  XOR U32478 ( .A(n35397), .B(n35398), .Z(n32551) );
  NOR U32479 ( .A(n35399), .B(n35397), .Z(n35398) );
  XOR U32480 ( .A(n35400), .B(n35401), .Z(n32554) );
  NOR U32481 ( .A(n35402), .B(n35400), .Z(n35401) );
  XOR U32482 ( .A(n35403), .B(n35404), .Z(n32557) );
  NOR U32483 ( .A(n35405), .B(n35403), .Z(n35404) );
  XOR U32484 ( .A(n35406), .B(n35407), .Z(n32560) );
  NOR U32485 ( .A(n35408), .B(n35406), .Z(n35407) );
  XOR U32486 ( .A(n35409), .B(n35410), .Z(n32563) );
  NOR U32487 ( .A(n35411), .B(n35409), .Z(n35410) );
  XOR U32488 ( .A(n35412), .B(n35413), .Z(n32566) );
  NOR U32489 ( .A(n35414), .B(n35412), .Z(n35413) );
  XOR U32490 ( .A(n35415), .B(n35416), .Z(n32569) );
  NOR U32491 ( .A(n35417), .B(n35415), .Z(n35416) );
  XOR U32492 ( .A(n35418), .B(n35419), .Z(n32572) );
  NOR U32493 ( .A(n35420), .B(n35418), .Z(n35419) );
  XOR U32494 ( .A(n35421), .B(n35422), .Z(n32575) );
  NOR U32495 ( .A(n35423), .B(n35421), .Z(n35422) );
  XOR U32496 ( .A(n35424), .B(n35425), .Z(n32578) );
  NOR U32497 ( .A(n35426), .B(n35424), .Z(n35425) );
  XOR U32498 ( .A(n35427), .B(n35428), .Z(n32581) );
  NOR U32499 ( .A(n35429), .B(n35427), .Z(n35428) );
  XOR U32500 ( .A(n35430), .B(n35431), .Z(n32584) );
  NOR U32501 ( .A(n35432), .B(n35430), .Z(n35431) );
  XOR U32502 ( .A(n35433), .B(n35434), .Z(n32587) );
  NOR U32503 ( .A(n35435), .B(n35433), .Z(n35434) );
  XOR U32504 ( .A(n35436), .B(n35437), .Z(n32590) );
  NOR U32505 ( .A(n35438), .B(n35436), .Z(n35437) );
  XOR U32506 ( .A(n35439), .B(n35440), .Z(n32593) );
  NOR U32507 ( .A(n35441), .B(n35439), .Z(n35440) );
  XOR U32508 ( .A(n35442), .B(n35443), .Z(n32596) );
  NOR U32509 ( .A(n35444), .B(n35442), .Z(n35443) );
  XOR U32510 ( .A(n35445), .B(n35446), .Z(n32599) );
  NOR U32511 ( .A(n35447), .B(n35445), .Z(n35446) );
  XOR U32512 ( .A(n35448), .B(n35449), .Z(n32602) );
  NOR U32513 ( .A(n35450), .B(n35448), .Z(n35449) );
  XOR U32514 ( .A(n35451), .B(n35452), .Z(n32605) );
  NOR U32515 ( .A(n35453), .B(n35451), .Z(n35452) );
  XOR U32516 ( .A(n35454), .B(n35455), .Z(n32608) );
  NOR U32517 ( .A(n35456), .B(n35454), .Z(n35455) );
  XOR U32518 ( .A(n35457), .B(n35458), .Z(n32611) );
  NOR U32519 ( .A(n35459), .B(n35457), .Z(n35458) );
  XOR U32520 ( .A(n35460), .B(n35461), .Z(n32614) );
  NOR U32521 ( .A(n35462), .B(n35460), .Z(n35461) );
  XOR U32522 ( .A(n35463), .B(n35464), .Z(n32617) );
  NOR U32523 ( .A(n35465), .B(n35463), .Z(n35464) );
  XOR U32524 ( .A(n35466), .B(n35467), .Z(n32620) );
  NOR U32525 ( .A(n35468), .B(n35466), .Z(n35467) );
  XOR U32526 ( .A(n35469), .B(n35470), .Z(n32623) );
  NOR U32527 ( .A(n35471), .B(n35469), .Z(n35470) );
  XOR U32528 ( .A(n35472), .B(n35473), .Z(n32626) );
  NOR U32529 ( .A(n35474), .B(n35472), .Z(n35473) );
  XOR U32530 ( .A(n35475), .B(n35476), .Z(n32629) );
  NOR U32531 ( .A(n35477), .B(n35475), .Z(n35476) );
  XOR U32532 ( .A(n35478), .B(n35479), .Z(n32632) );
  NOR U32533 ( .A(n35480), .B(n35478), .Z(n35479) );
  XOR U32534 ( .A(n35481), .B(n35482), .Z(n32635) );
  NOR U32535 ( .A(n35483), .B(n35481), .Z(n35482) );
  XOR U32536 ( .A(n35484), .B(n35485), .Z(n32638) );
  NOR U32537 ( .A(n35486), .B(n35484), .Z(n35485) );
  XOR U32538 ( .A(n35487), .B(n35488), .Z(n32641) );
  NOR U32539 ( .A(n35489), .B(n35487), .Z(n35488) );
  XOR U32540 ( .A(n35490), .B(n35491), .Z(n32644) );
  NOR U32541 ( .A(n35492), .B(n35490), .Z(n35491) );
  XOR U32542 ( .A(n35493), .B(n35494), .Z(n32647) );
  NOR U32543 ( .A(n35495), .B(n35493), .Z(n35494) );
  XOR U32544 ( .A(n35496), .B(n35497), .Z(n32650) );
  NOR U32545 ( .A(n35498), .B(n35496), .Z(n35497) );
  XOR U32546 ( .A(n35499), .B(n35500), .Z(n32653) );
  NOR U32547 ( .A(n35501), .B(n35499), .Z(n35500) );
  XOR U32548 ( .A(n35502), .B(n35503), .Z(n32656) );
  NOR U32549 ( .A(n35504), .B(n35502), .Z(n35503) );
  XOR U32550 ( .A(n35505), .B(n35506), .Z(n32659) );
  NOR U32551 ( .A(n35507), .B(n35505), .Z(n35506) );
  XOR U32552 ( .A(n35508), .B(n35509), .Z(n32662) );
  NOR U32553 ( .A(n35510), .B(n35508), .Z(n35509) );
  XOR U32554 ( .A(n35511), .B(n35512), .Z(n32665) );
  NOR U32555 ( .A(n35513), .B(n35511), .Z(n35512) );
  XOR U32556 ( .A(n35514), .B(n35515), .Z(n32668) );
  NOR U32557 ( .A(n35516), .B(n35514), .Z(n35515) );
  XOR U32558 ( .A(n35517), .B(n35518), .Z(n32671) );
  NOR U32559 ( .A(n35519), .B(n35517), .Z(n35518) );
  XOR U32560 ( .A(n35520), .B(n35521), .Z(n32674) );
  NOR U32561 ( .A(n35522), .B(n35520), .Z(n35521) );
  XOR U32562 ( .A(n35523), .B(n35524), .Z(n32677) );
  NOR U32563 ( .A(n35525), .B(n35523), .Z(n35524) );
  XOR U32564 ( .A(n35526), .B(n35527), .Z(n32680) );
  NOR U32565 ( .A(n35528), .B(n35526), .Z(n35527) );
  XOR U32566 ( .A(n35529), .B(n35530), .Z(n32683) );
  AND U32567 ( .A(n35531), .B(n35529), .Z(n35530) );
  XOR U32568 ( .A(n35532), .B(n35533), .Z(n32686) );
  AND U32569 ( .A(n109), .B(n35532), .Z(n35533) );
  XOR U32570 ( .A(n91), .B(n34102), .Z(n34104) );
  XOR U32571 ( .A(n34099), .B(n34098), .Z(n91) );
  XNOR U32572 ( .A(n34096), .B(n34095), .Z(n34098) );
  XNOR U32573 ( .A(n34093), .B(n34092), .Z(n34095) );
  XNOR U32574 ( .A(n34090), .B(n34089), .Z(n34092) );
  XNOR U32575 ( .A(n34087), .B(n34086), .Z(n34089) );
  XNOR U32576 ( .A(n34084), .B(n34083), .Z(n34086) );
  XNOR U32577 ( .A(n34081), .B(n34080), .Z(n34083) );
  XNOR U32578 ( .A(n34078), .B(n34077), .Z(n34080) );
  XNOR U32579 ( .A(n34075), .B(n34074), .Z(n34077) );
  XNOR U32580 ( .A(n34072), .B(n34071), .Z(n34074) );
  XNOR U32581 ( .A(n34069), .B(n34068), .Z(n34071) );
  XNOR U32582 ( .A(n34066), .B(n34065), .Z(n34068) );
  XNOR U32583 ( .A(n34063), .B(n34062), .Z(n34065) );
  XNOR U32584 ( .A(n34060), .B(n34059), .Z(n34062) );
  XNOR U32585 ( .A(n34057), .B(n34056), .Z(n34059) );
  XNOR U32586 ( .A(n34054), .B(n34053), .Z(n34056) );
  XNOR U32587 ( .A(n34051), .B(n34050), .Z(n34053) );
  XNOR U32588 ( .A(n34048), .B(n34047), .Z(n34050) );
  XNOR U32589 ( .A(n34045), .B(n34044), .Z(n34047) );
  XNOR U32590 ( .A(n34042), .B(n34041), .Z(n34044) );
  XNOR U32591 ( .A(n34039), .B(n34038), .Z(n34041) );
  XNOR U32592 ( .A(n34036), .B(n34035), .Z(n34038) );
  XNOR U32593 ( .A(n34033), .B(n34032), .Z(n34035) );
  XNOR U32594 ( .A(n34030), .B(n34029), .Z(n34032) );
  XNOR U32595 ( .A(n34027), .B(n34026), .Z(n34029) );
  XNOR U32596 ( .A(n34024), .B(n34023), .Z(n34026) );
  XNOR U32597 ( .A(n34021), .B(n34020), .Z(n34023) );
  XNOR U32598 ( .A(n34018), .B(n34017), .Z(n34020) );
  XNOR U32599 ( .A(n34015), .B(n34014), .Z(n34017) );
  XNOR U32600 ( .A(n34012), .B(n34011), .Z(n34014) );
  XNOR U32601 ( .A(n34009), .B(n34008), .Z(n34011) );
  XNOR U32602 ( .A(n34006), .B(n34005), .Z(n34008) );
  XNOR U32603 ( .A(n34003), .B(n34002), .Z(n34005) );
  XNOR U32604 ( .A(n34000), .B(n33999), .Z(n34002) );
  XNOR U32605 ( .A(n33997), .B(n33996), .Z(n33999) );
  XNOR U32606 ( .A(n33994), .B(n33993), .Z(n33996) );
  XNOR U32607 ( .A(n33991), .B(n33990), .Z(n33993) );
  XNOR U32608 ( .A(n33988), .B(n33987), .Z(n33990) );
  XNOR U32609 ( .A(n33985), .B(n33984), .Z(n33987) );
  XNOR U32610 ( .A(n33982), .B(n33981), .Z(n33984) );
  XNOR U32611 ( .A(n33979), .B(n33978), .Z(n33981) );
  XNOR U32612 ( .A(n33976), .B(n33975), .Z(n33978) );
  XNOR U32613 ( .A(n33973), .B(n33972), .Z(n33975) );
  XNOR U32614 ( .A(n33970), .B(n33969), .Z(n33972) );
  XNOR U32615 ( .A(n33967), .B(n33966), .Z(n33969) );
  XNOR U32616 ( .A(n33964), .B(n33963), .Z(n33966) );
  XNOR U32617 ( .A(n33961), .B(n33960), .Z(n33963) );
  XNOR U32618 ( .A(n33958), .B(n33957), .Z(n33960) );
  XNOR U32619 ( .A(n33955), .B(n33954), .Z(n33957) );
  XNOR U32620 ( .A(n33952), .B(n33951), .Z(n33954) );
  XNOR U32621 ( .A(n33949), .B(n33948), .Z(n33951) );
  XNOR U32622 ( .A(n33946), .B(n33945), .Z(n33948) );
  XNOR U32623 ( .A(n33943), .B(n33942), .Z(n33945) );
  XNOR U32624 ( .A(n33940), .B(n33939), .Z(n33942) );
  XNOR U32625 ( .A(n33937), .B(n33936), .Z(n33939) );
  XNOR U32626 ( .A(n33934), .B(n33933), .Z(n33936) );
  XNOR U32627 ( .A(n33931), .B(n33930), .Z(n33933) );
  XNOR U32628 ( .A(n33928), .B(n33927), .Z(n33930) );
  XNOR U32629 ( .A(n33925), .B(n33924), .Z(n33927) );
  XNOR U32630 ( .A(n33922), .B(n33921), .Z(n33924) );
  XNOR U32631 ( .A(n33919), .B(n33918), .Z(n33921) );
  XNOR U32632 ( .A(n33916), .B(n33915), .Z(n33918) );
  XNOR U32633 ( .A(n33913), .B(n33912), .Z(n33915) );
  XNOR U32634 ( .A(n33910), .B(n33909), .Z(n33912) );
  XNOR U32635 ( .A(n33907), .B(n33906), .Z(n33909) );
  XNOR U32636 ( .A(n33904), .B(n33903), .Z(n33906) );
  XNOR U32637 ( .A(n33901), .B(n33900), .Z(n33903) );
  XNOR U32638 ( .A(n33898), .B(n33897), .Z(n33900) );
  XNOR U32639 ( .A(n33895), .B(n33894), .Z(n33897) );
  XNOR U32640 ( .A(n33892), .B(n33891), .Z(n33894) );
  XNOR U32641 ( .A(n33889), .B(n33888), .Z(n33891) );
  XNOR U32642 ( .A(n33886), .B(n33885), .Z(n33888) );
  XNOR U32643 ( .A(n33883), .B(n33882), .Z(n33885) );
  XNOR U32644 ( .A(n33880), .B(n33879), .Z(n33882) );
  XNOR U32645 ( .A(n33877), .B(n33876), .Z(n33879) );
  XNOR U32646 ( .A(n33874), .B(n33873), .Z(n33876) );
  XNOR U32647 ( .A(n33871), .B(n33870), .Z(n33873) );
  XNOR U32648 ( .A(n33868), .B(n33867), .Z(n33870) );
  XNOR U32649 ( .A(n33865), .B(n33864), .Z(n33867) );
  XNOR U32650 ( .A(n33862), .B(n33861), .Z(n33864) );
  XNOR U32651 ( .A(n33859), .B(n33858), .Z(n33861) );
  XNOR U32652 ( .A(n33856), .B(n33855), .Z(n33858) );
  XNOR U32653 ( .A(n33853), .B(n33852), .Z(n33855) );
  XNOR U32654 ( .A(n33850), .B(n33849), .Z(n33852) );
  XNOR U32655 ( .A(n33847), .B(n33846), .Z(n33849) );
  XNOR U32656 ( .A(n33844), .B(n33843), .Z(n33846) );
  XNOR U32657 ( .A(n33841), .B(n33840), .Z(n33843) );
  XNOR U32658 ( .A(n33838), .B(n33837), .Z(n33840) );
  XNOR U32659 ( .A(n33835), .B(n33834), .Z(n33837) );
  XNOR U32660 ( .A(n33832), .B(n33831), .Z(n33834) );
  XNOR U32661 ( .A(n33829), .B(n33828), .Z(n33831) );
  XNOR U32662 ( .A(n33826), .B(n33825), .Z(n33828) );
  XNOR U32663 ( .A(n33823), .B(n33822), .Z(n33825) );
  XNOR U32664 ( .A(n33820), .B(n33819), .Z(n33822) );
  XNOR U32665 ( .A(n33817), .B(n33816), .Z(n33819) );
  XNOR U32666 ( .A(n33814), .B(n33813), .Z(n33816) );
  XNOR U32667 ( .A(n33811), .B(n33810), .Z(n33813) );
  XNOR U32668 ( .A(n33808), .B(n33807), .Z(n33810) );
  XNOR U32669 ( .A(n33805), .B(n33804), .Z(n33807) );
  XNOR U32670 ( .A(n33802), .B(n33801), .Z(n33804) );
  XNOR U32671 ( .A(n33799), .B(n33798), .Z(n33801) );
  XNOR U32672 ( .A(n33796), .B(n33795), .Z(n33798) );
  XNOR U32673 ( .A(n33793), .B(n33792), .Z(n33795) );
  XNOR U32674 ( .A(n33790), .B(n33789), .Z(n33792) );
  XNOR U32675 ( .A(n33787), .B(n33786), .Z(n33789) );
  XNOR U32676 ( .A(n33784), .B(n33783), .Z(n33786) );
  XNOR U32677 ( .A(n33781), .B(n33780), .Z(n33783) );
  XNOR U32678 ( .A(n33778), .B(n33777), .Z(n33780) );
  XNOR U32679 ( .A(n33775), .B(n33774), .Z(n33777) );
  XNOR U32680 ( .A(n33772), .B(n33771), .Z(n33774) );
  XNOR U32681 ( .A(n33769), .B(n33768), .Z(n33771) );
  XNOR U32682 ( .A(n33766), .B(n33765), .Z(n33768) );
  XNOR U32683 ( .A(n33763), .B(n33762), .Z(n33765) );
  XNOR U32684 ( .A(n33760), .B(n33759), .Z(n33762) );
  XNOR U32685 ( .A(n33757), .B(n33756), .Z(n33759) );
  XNOR U32686 ( .A(n33754), .B(n33753), .Z(n33756) );
  XNOR U32687 ( .A(n33751), .B(n33750), .Z(n33753) );
  XNOR U32688 ( .A(n33748), .B(n33747), .Z(n33750) );
  XNOR U32689 ( .A(n33745), .B(n33744), .Z(n33747) );
  XNOR U32690 ( .A(n33742), .B(n33741), .Z(n33744) );
  XNOR U32691 ( .A(n33739), .B(n33738), .Z(n33741) );
  XNOR U32692 ( .A(n33736), .B(n33735), .Z(n33738) );
  XNOR U32693 ( .A(n33733), .B(n33732), .Z(n33735) );
  XNOR U32694 ( .A(n33730), .B(n33729), .Z(n33732) );
  XNOR U32695 ( .A(n33727), .B(n33726), .Z(n33729) );
  XNOR U32696 ( .A(n33724), .B(n33723), .Z(n33726) );
  XNOR U32697 ( .A(n33721), .B(n33720), .Z(n33723) );
  XNOR U32698 ( .A(n33718), .B(n33717), .Z(n33720) );
  XNOR U32699 ( .A(n33715), .B(n33714), .Z(n33717) );
  XNOR U32700 ( .A(n33712), .B(n33711), .Z(n33714) );
  XNOR U32701 ( .A(n33709), .B(n33708), .Z(n33711) );
  XNOR U32702 ( .A(n33706), .B(n33705), .Z(n33708) );
  XNOR U32703 ( .A(n33703), .B(n33702), .Z(n33705) );
  XNOR U32704 ( .A(n33700), .B(n33699), .Z(n33702) );
  XNOR U32705 ( .A(n33697), .B(n33696), .Z(n33699) );
  XNOR U32706 ( .A(n33694), .B(n33693), .Z(n33696) );
  XNOR U32707 ( .A(n33691), .B(n33690), .Z(n33693) );
  XNOR U32708 ( .A(n33688), .B(n33687), .Z(n33690) );
  XNOR U32709 ( .A(n33685), .B(n33684), .Z(n33687) );
  XNOR U32710 ( .A(n33682), .B(n33681), .Z(n33684) );
  XNOR U32711 ( .A(n33679), .B(n33678), .Z(n33681) );
  XNOR U32712 ( .A(n33676), .B(n33675), .Z(n33678) );
  XNOR U32713 ( .A(n33673), .B(n33672), .Z(n33675) );
  XNOR U32714 ( .A(n33670), .B(n33669), .Z(n33672) );
  XNOR U32715 ( .A(n33667), .B(n33666), .Z(n33669) );
  XNOR U32716 ( .A(n33664), .B(n33663), .Z(n33666) );
  XNOR U32717 ( .A(n33661), .B(n33660), .Z(n33663) );
  XNOR U32718 ( .A(n33658), .B(n33657), .Z(n33660) );
  XNOR U32719 ( .A(n33655), .B(n33654), .Z(n33657) );
  XNOR U32720 ( .A(n33652), .B(n33651), .Z(n33654) );
  XNOR U32721 ( .A(n33649), .B(n33648), .Z(n33651) );
  XNOR U32722 ( .A(n33646), .B(n33645), .Z(n33648) );
  XNOR U32723 ( .A(n33643), .B(n33642), .Z(n33645) );
  XNOR U32724 ( .A(n33640), .B(n33639), .Z(n33642) );
  XNOR U32725 ( .A(n33637), .B(n33636), .Z(n33639) );
  XNOR U32726 ( .A(n33634), .B(n33633), .Z(n33636) );
  XNOR U32727 ( .A(n33631), .B(n33630), .Z(n33633) );
  XNOR U32728 ( .A(n33628), .B(n33627), .Z(n33630) );
  XNOR U32729 ( .A(n33625), .B(n33624), .Z(n33627) );
  XNOR U32730 ( .A(n33622), .B(n33621), .Z(n33624) );
  XNOR U32731 ( .A(n33619), .B(n33618), .Z(n33621) );
  XNOR U32732 ( .A(n33616), .B(n33615), .Z(n33618) );
  XNOR U32733 ( .A(n33613), .B(n33612), .Z(n33615) );
  XNOR U32734 ( .A(n33610), .B(n33609), .Z(n33612) );
  XNOR U32735 ( .A(n33607), .B(n33606), .Z(n33609) );
  XNOR U32736 ( .A(n33604), .B(n33603), .Z(n33606) );
  XNOR U32737 ( .A(n33601), .B(n33600), .Z(n33603) );
  XNOR U32738 ( .A(n33598), .B(n33597), .Z(n33600) );
  XNOR U32739 ( .A(n33595), .B(n33594), .Z(n33597) );
  XNOR U32740 ( .A(n33592), .B(n33591), .Z(n33594) );
  XNOR U32741 ( .A(n33589), .B(n33588), .Z(n33591) );
  XNOR U32742 ( .A(n33586), .B(n33585), .Z(n33588) );
  XNOR U32743 ( .A(n33583), .B(n33582), .Z(n33585) );
  XNOR U32744 ( .A(n33580), .B(n33579), .Z(n33582) );
  XNOR U32745 ( .A(n33577), .B(n33576), .Z(n33579) );
  XNOR U32746 ( .A(n33574), .B(n33573), .Z(n33576) );
  XNOR U32747 ( .A(n33571), .B(n33570), .Z(n33573) );
  XNOR U32748 ( .A(n33568), .B(n33567), .Z(n33570) );
  XNOR U32749 ( .A(n33565), .B(n33564), .Z(n33567) );
  XNOR U32750 ( .A(n33562), .B(n33561), .Z(n33564) );
  XNOR U32751 ( .A(n33559), .B(n33558), .Z(n33561) );
  XNOR U32752 ( .A(n33556), .B(n33555), .Z(n33558) );
  XNOR U32753 ( .A(n33553), .B(n33552), .Z(n33555) );
  XNOR U32754 ( .A(n33550), .B(n33549), .Z(n33552) );
  XNOR U32755 ( .A(n33547), .B(n33546), .Z(n33549) );
  XNOR U32756 ( .A(n33544), .B(n33543), .Z(n33546) );
  XNOR U32757 ( .A(n33541), .B(n33540), .Z(n33543) );
  XNOR U32758 ( .A(n33538), .B(n33537), .Z(n33540) );
  XNOR U32759 ( .A(n33535), .B(n33534), .Z(n33537) );
  XNOR U32760 ( .A(n33532), .B(n33531), .Z(n33534) );
  XNOR U32761 ( .A(n33529), .B(n33528), .Z(n33531) );
  XNOR U32762 ( .A(n33526), .B(n33525), .Z(n33528) );
  XNOR U32763 ( .A(n33523), .B(n33522), .Z(n33525) );
  XNOR U32764 ( .A(n33520), .B(n33519), .Z(n33522) );
  XNOR U32765 ( .A(n33517), .B(n33516), .Z(n33519) );
  XNOR U32766 ( .A(n33514), .B(n33513), .Z(n33516) );
  XNOR U32767 ( .A(n33511), .B(n33510), .Z(n33513) );
  XNOR U32768 ( .A(n33508), .B(n33507), .Z(n33510) );
  XNOR U32769 ( .A(n33505), .B(n33504), .Z(n33507) );
  XNOR U32770 ( .A(n33502), .B(n33501), .Z(n33504) );
  XNOR U32771 ( .A(n33499), .B(n33498), .Z(n33501) );
  XNOR U32772 ( .A(n33496), .B(n33495), .Z(n33498) );
  XNOR U32773 ( .A(n33493), .B(n33492), .Z(n33495) );
  XNOR U32774 ( .A(n33490), .B(n33489), .Z(n33492) );
  XNOR U32775 ( .A(n33487), .B(n33486), .Z(n33489) );
  XNOR U32776 ( .A(n33484), .B(n33483), .Z(n33486) );
  XNOR U32777 ( .A(n33481), .B(n33480), .Z(n33483) );
  XNOR U32778 ( .A(n33478), .B(n33477), .Z(n33480) );
  XNOR U32779 ( .A(n33475), .B(n33474), .Z(n33477) );
  XNOR U32780 ( .A(n33472), .B(n33471), .Z(n33474) );
  XNOR U32781 ( .A(n33469), .B(n33468), .Z(n33471) );
  XNOR U32782 ( .A(n33466), .B(n33465), .Z(n33468) );
  XNOR U32783 ( .A(n33463), .B(n33462), .Z(n33465) );
  XNOR U32784 ( .A(n33460), .B(n33459), .Z(n33462) );
  XNOR U32785 ( .A(n33457), .B(n33456), .Z(n33459) );
  XNOR U32786 ( .A(n33454), .B(n33453), .Z(n33456) );
  XNOR U32787 ( .A(n33451), .B(n33450), .Z(n33453) );
  XNOR U32788 ( .A(n33448), .B(n33447), .Z(n33450) );
  XNOR U32789 ( .A(n33445), .B(n33444), .Z(n33447) );
  XNOR U32790 ( .A(n33442), .B(n33441), .Z(n33444) );
  XNOR U32791 ( .A(n33439), .B(n33438), .Z(n33441) );
  XNOR U32792 ( .A(n33436), .B(n33435), .Z(n33438) );
  XNOR U32793 ( .A(n33433), .B(n33432), .Z(n33435) );
  XNOR U32794 ( .A(n33430), .B(n33429), .Z(n33432) );
  XNOR U32795 ( .A(n33427), .B(n33426), .Z(n33429) );
  XNOR U32796 ( .A(n33424), .B(n33423), .Z(n33426) );
  XNOR U32797 ( .A(n33421), .B(n33420), .Z(n33423) );
  XNOR U32798 ( .A(n33418), .B(n33417), .Z(n33420) );
  XNOR U32799 ( .A(n33415), .B(n33414), .Z(n33417) );
  XNOR U32800 ( .A(n33412), .B(n33411), .Z(n33414) );
  XNOR U32801 ( .A(n33409), .B(n33408), .Z(n33411) );
  XNOR U32802 ( .A(n33406), .B(n33405), .Z(n33408) );
  XNOR U32803 ( .A(n33403), .B(n33402), .Z(n33405) );
  XNOR U32804 ( .A(n33400), .B(n33399), .Z(n33402) );
  XNOR U32805 ( .A(n33397), .B(n33396), .Z(n33399) );
  XNOR U32806 ( .A(n33394), .B(n33393), .Z(n33396) );
  XNOR U32807 ( .A(n33391), .B(n33390), .Z(n33393) );
  XNOR U32808 ( .A(n33388), .B(n33387), .Z(n33390) );
  XNOR U32809 ( .A(n33385), .B(n33384), .Z(n33387) );
  XNOR U32810 ( .A(n33382), .B(n33381), .Z(n33384) );
  XNOR U32811 ( .A(n33379), .B(n33378), .Z(n33381) );
  XNOR U32812 ( .A(n33376), .B(n33375), .Z(n33378) );
  XNOR U32813 ( .A(n33373), .B(n33372), .Z(n33375) );
  XNOR U32814 ( .A(n33370), .B(n33369), .Z(n33372) );
  XNOR U32815 ( .A(n33367), .B(n33366), .Z(n33369) );
  XNOR U32816 ( .A(n33364), .B(n33363), .Z(n33366) );
  XNOR U32817 ( .A(n33361), .B(n33360), .Z(n33363) );
  XNOR U32818 ( .A(n33358), .B(n33357), .Z(n33360) );
  XNOR U32819 ( .A(n33355), .B(n33354), .Z(n33357) );
  XNOR U32820 ( .A(n33352), .B(n33351), .Z(n33354) );
  XNOR U32821 ( .A(n33349), .B(n33348), .Z(n33351) );
  XNOR U32822 ( .A(n33346), .B(n33345), .Z(n33348) );
  XNOR U32823 ( .A(n33343), .B(n33342), .Z(n33345) );
  XNOR U32824 ( .A(n33340), .B(n33339), .Z(n33342) );
  XNOR U32825 ( .A(n33337), .B(n33336), .Z(n33339) );
  XNOR U32826 ( .A(n33334), .B(n33333), .Z(n33336) );
  XNOR U32827 ( .A(n33331), .B(n33330), .Z(n33333) );
  XNOR U32828 ( .A(n33328), .B(n33327), .Z(n33330) );
  XNOR U32829 ( .A(n33325), .B(n33324), .Z(n33327) );
  XNOR U32830 ( .A(n33322), .B(n33321), .Z(n33324) );
  XNOR U32831 ( .A(n33319), .B(n33318), .Z(n33321) );
  XNOR U32832 ( .A(n33316), .B(n33315), .Z(n33318) );
  XNOR U32833 ( .A(n33313), .B(n33312), .Z(n33315) );
  XNOR U32834 ( .A(n33310), .B(n33309), .Z(n33312) );
  XNOR U32835 ( .A(n33307), .B(n33306), .Z(n33309) );
  XNOR U32836 ( .A(n33304), .B(n33303), .Z(n33306) );
  XNOR U32837 ( .A(n33301), .B(n33300), .Z(n33303) );
  XNOR U32838 ( .A(n33298), .B(n33297), .Z(n33300) );
  XNOR U32839 ( .A(n33295), .B(n33294), .Z(n33297) );
  XNOR U32840 ( .A(n33292), .B(n33291), .Z(n33294) );
  XNOR U32841 ( .A(n33289), .B(n33288), .Z(n33291) );
  XNOR U32842 ( .A(n33286), .B(n33285), .Z(n33288) );
  XNOR U32843 ( .A(n33283), .B(n33282), .Z(n33285) );
  XNOR U32844 ( .A(n33280), .B(n33279), .Z(n33282) );
  XNOR U32845 ( .A(n33277), .B(n33276), .Z(n33279) );
  XNOR U32846 ( .A(n33274), .B(n33273), .Z(n33276) );
  XNOR U32847 ( .A(n33271), .B(n33270), .Z(n33273) );
  XNOR U32848 ( .A(n33268), .B(n33267), .Z(n33270) );
  XNOR U32849 ( .A(n33265), .B(n33264), .Z(n33267) );
  XNOR U32850 ( .A(n33262), .B(n33261), .Z(n33264) );
  XNOR U32851 ( .A(n33259), .B(n33258), .Z(n33261) );
  XNOR U32852 ( .A(n33256), .B(n33255), .Z(n33258) );
  XNOR U32853 ( .A(n33253), .B(n33252), .Z(n33255) );
  XNOR U32854 ( .A(n33250), .B(n33249), .Z(n33252) );
  XNOR U32855 ( .A(n33247), .B(n33246), .Z(n33249) );
  XNOR U32856 ( .A(n33244), .B(n33243), .Z(n33246) );
  XNOR U32857 ( .A(n33241), .B(n33240), .Z(n33243) );
  XNOR U32858 ( .A(n33238), .B(n33237), .Z(n33240) );
  XNOR U32859 ( .A(n33235), .B(n33234), .Z(n33237) );
  XNOR U32860 ( .A(n33232), .B(n33231), .Z(n33234) );
  XNOR U32861 ( .A(n33229), .B(n33228), .Z(n33231) );
  XNOR U32862 ( .A(n33226), .B(n33225), .Z(n33228) );
  XNOR U32863 ( .A(n33223), .B(n33222), .Z(n33225) );
  XNOR U32864 ( .A(n33220), .B(n33219), .Z(n33222) );
  XNOR U32865 ( .A(n33217), .B(n33216), .Z(n33219) );
  XNOR U32866 ( .A(n33214), .B(n33213), .Z(n33216) );
  XNOR U32867 ( .A(n33211), .B(n33210), .Z(n33213) );
  XNOR U32868 ( .A(n33208), .B(n33207), .Z(n33210) );
  XNOR U32869 ( .A(n33205), .B(n33204), .Z(n33207) );
  XNOR U32870 ( .A(n33202), .B(n33201), .Z(n33204) );
  XNOR U32871 ( .A(n33199), .B(n33198), .Z(n33201) );
  XNOR U32872 ( .A(n33196), .B(n33195), .Z(n33198) );
  XNOR U32873 ( .A(n33193), .B(n33192), .Z(n33195) );
  XNOR U32874 ( .A(n33190), .B(n33189), .Z(n33192) );
  XNOR U32875 ( .A(n33187), .B(n33186), .Z(n33189) );
  XNOR U32876 ( .A(n33184), .B(n33183), .Z(n33186) );
  XNOR U32877 ( .A(n33181), .B(n33180), .Z(n33183) );
  XNOR U32878 ( .A(n33178), .B(n33177), .Z(n33180) );
  XNOR U32879 ( .A(n33175), .B(n33174), .Z(n33177) );
  XNOR U32880 ( .A(n33172), .B(n33171), .Z(n33174) );
  XNOR U32881 ( .A(n33169), .B(n33168), .Z(n33171) );
  XNOR U32882 ( .A(n33166), .B(n33165), .Z(n33168) );
  XNOR U32883 ( .A(n33163), .B(n33162), .Z(n33165) );
  XNOR U32884 ( .A(n33160), .B(n33159), .Z(n33162) );
  XNOR U32885 ( .A(n33157), .B(n33156), .Z(n33159) );
  XNOR U32886 ( .A(n33154), .B(n33153), .Z(n33156) );
  XNOR U32887 ( .A(n33151), .B(n33150), .Z(n33153) );
  XNOR U32888 ( .A(n33148), .B(n33147), .Z(n33150) );
  XNOR U32889 ( .A(n33145), .B(n33144), .Z(n33147) );
  XNOR U32890 ( .A(n33142), .B(n33141), .Z(n33144) );
  XNOR U32891 ( .A(n33139), .B(n33138), .Z(n33141) );
  XNOR U32892 ( .A(n33136), .B(n33135), .Z(n33138) );
  XNOR U32893 ( .A(n33133), .B(n33132), .Z(n33135) );
  XNOR U32894 ( .A(n33130), .B(n33129), .Z(n33132) );
  XNOR U32895 ( .A(n33127), .B(n33126), .Z(n33129) );
  XNOR U32896 ( .A(n33124), .B(n33123), .Z(n33126) );
  XNOR U32897 ( .A(n33121), .B(n33120), .Z(n33123) );
  XNOR U32898 ( .A(n33118), .B(n33117), .Z(n33120) );
  XNOR U32899 ( .A(n33115), .B(n33114), .Z(n33117) );
  XNOR U32900 ( .A(n33112), .B(n33111), .Z(n33114) );
  XNOR U32901 ( .A(n33109), .B(n33108), .Z(n33111) );
  XNOR U32902 ( .A(n33106), .B(n33105), .Z(n33108) );
  XNOR U32903 ( .A(n33103), .B(n33102), .Z(n33105) );
  XNOR U32904 ( .A(n33100), .B(n33099), .Z(n33102) );
  XNOR U32905 ( .A(n33097), .B(n33096), .Z(n33099) );
  XNOR U32906 ( .A(n33094), .B(n33093), .Z(n33096) );
  XNOR U32907 ( .A(n33091), .B(n33090), .Z(n33093) );
  XNOR U32908 ( .A(n33088), .B(n33087), .Z(n33090) );
  XNOR U32909 ( .A(n33085), .B(n33084), .Z(n33087) );
  XNOR U32910 ( .A(n33082), .B(n33081), .Z(n33084) );
  XNOR U32911 ( .A(n33079), .B(n33078), .Z(n33081) );
  XNOR U32912 ( .A(n33076), .B(n33075), .Z(n33078) );
  XNOR U32913 ( .A(n33073), .B(n33072), .Z(n33075) );
  XNOR U32914 ( .A(n33070), .B(n33069), .Z(n33072) );
  XNOR U32915 ( .A(n33067), .B(n33066), .Z(n33069) );
  XNOR U32916 ( .A(n33064), .B(n33063), .Z(n33066) );
  XNOR U32917 ( .A(n33061), .B(n33060), .Z(n33063) );
  XNOR U32918 ( .A(n33058), .B(n33057), .Z(n33060) );
  XNOR U32919 ( .A(n33055), .B(n33054), .Z(n33057) );
  XNOR U32920 ( .A(n33052), .B(n33051), .Z(n33054) );
  XNOR U32921 ( .A(n33049), .B(n33048), .Z(n33051) );
  XNOR U32922 ( .A(n33046), .B(n33045), .Z(n33048) );
  XNOR U32923 ( .A(n33043), .B(n33042), .Z(n33045) );
  XNOR U32924 ( .A(n33040), .B(n33039), .Z(n33042) );
  XNOR U32925 ( .A(n33037), .B(n33036), .Z(n33039) );
  XNOR U32926 ( .A(n33034), .B(n33033), .Z(n33036) );
  XNOR U32927 ( .A(n33031), .B(n33030), .Z(n33033) );
  XNOR U32928 ( .A(n33028), .B(n33027), .Z(n33030) );
  XNOR U32929 ( .A(n33025), .B(n33024), .Z(n33027) );
  XNOR U32930 ( .A(n33022), .B(n33021), .Z(n33024) );
  XNOR U32931 ( .A(n33019), .B(n33018), .Z(n33021) );
  XNOR U32932 ( .A(n33016), .B(n33015), .Z(n33018) );
  XNOR U32933 ( .A(n33013), .B(n33012), .Z(n33015) );
  XNOR U32934 ( .A(n33010), .B(n33009), .Z(n33012) );
  XNOR U32935 ( .A(n33007), .B(n33006), .Z(n33009) );
  XNOR U32936 ( .A(n33004), .B(n33003), .Z(n33006) );
  XNOR U32937 ( .A(n33001), .B(n33000), .Z(n33003) );
  XNOR U32938 ( .A(n32998), .B(n32997), .Z(n33000) );
  XNOR U32939 ( .A(n32995), .B(n32994), .Z(n32997) );
  XNOR U32940 ( .A(n32992), .B(n32991), .Z(n32994) );
  XNOR U32941 ( .A(n32989), .B(n32988), .Z(n32991) );
  XNOR U32942 ( .A(n32986), .B(n32985), .Z(n32988) );
  XNOR U32943 ( .A(n32983), .B(n32982), .Z(n32985) );
  XNOR U32944 ( .A(n32980), .B(n32979), .Z(n32982) );
  XNOR U32945 ( .A(n32977), .B(n32976), .Z(n32979) );
  XNOR U32946 ( .A(n32974), .B(n32973), .Z(n32976) );
  XNOR U32947 ( .A(n32971), .B(n32970), .Z(n32973) );
  XNOR U32948 ( .A(n32968), .B(n32967), .Z(n32970) );
  XNOR U32949 ( .A(n32965), .B(n32964), .Z(n32967) );
  XNOR U32950 ( .A(n32962), .B(n32961), .Z(n32964) );
  XNOR U32951 ( .A(n32959), .B(n32958), .Z(n32961) );
  XNOR U32952 ( .A(n32956), .B(n32955), .Z(n32958) );
  XNOR U32953 ( .A(n32953), .B(n32952), .Z(n32955) );
  XNOR U32954 ( .A(n32950), .B(n32949), .Z(n32952) );
  XNOR U32955 ( .A(n32947), .B(n32946), .Z(n32949) );
  XNOR U32956 ( .A(n32944), .B(n32943), .Z(n32946) );
  XNOR U32957 ( .A(n32941), .B(n32940), .Z(n32943) );
  XNOR U32958 ( .A(n32938), .B(n32937), .Z(n32940) );
  XNOR U32959 ( .A(n32935), .B(n32934), .Z(n32937) );
  XNOR U32960 ( .A(n32932), .B(n32931), .Z(n32934) );
  XNOR U32961 ( .A(n32929), .B(n32928), .Z(n32931) );
  XNOR U32962 ( .A(n32926), .B(n32925), .Z(n32928) );
  XOR U32963 ( .A(n35534), .B(n32922), .Z(n32925) );
  XOR U32964 ( .A(n32920), .B(n32919), .Z(n32922) );
  XOR U32965 ( .A(n32917), .B(n32916), .Z(n32919) );
  XOR U32966 ( .A(n32913), .B(n32914), .Z(n32916) );
  AND U32967 ( .A(n35535), .B(n35536), .Z(n32914) );
  XOR U32968 ( .A(n32910), .B(n32911), .Z(n32913) );
  AND U32969 ( .A(n35537), .B(n35538), .Z(n32911) );
  XOR U32970 ( .A(n32907), .B(n32908), .Z(n32910) );
  AND U32971 ( .A(n35539), .B(n35540), .Z(n32908) );
  XOR U32972 ( .A(n32904), .B(n32905), .Z(n32907) );
  AND U32973 ( .A(n35541), .B(n35542), .Z(n32905) );
  XNOR U32974 ( .A(n32689), .B(n32902), .Z(n32904) );
  AND U32975 ( .A(n35543), .B(n35544), .Z(n32902) );
  XOR U32976 ( .A(n32691), .B(n32690), .Z(n32689) );
  AND U32977 ( .A(n35545), .B(n35546), .Z(n32690) );
  XOR U32978 ( .A(n32693), .B(n32692), .Z(n32691) );
  AND U32979 ( .A(n35547), .B(n35548), .Z(n32692) );
  XOR U32980 ( .A(n32695), .B(n32694), .Z(n32693) );
  AND U32981 ( .A(n35549), .B(n35550), .Z(n32694) );
  XOR U32982 ( .A(n32697), .B(n32696), .Z(n32695) );
  AND U32983 ( .A(n35551), .B(n35552), .Z(n32696) );
  XOR U32984 ( .A(n32699), .B(n32698), .Z(n32697) );
  AND U32985 ( .A(n35553), .B(n35554), .Z(n32698) );
  XOR U32986 ( .A(n32701), .B(n32700), .Z(n32699) );
  AND U32987 ( .A(n35555), .B(n35556), .Z(n32700) );
  XOR U32988 ( .A(n32703), .B(n32702), .Z(n32701) );
  AND U32989 ( .A(n35557), .B(n35558), .Z(n32702) );
  XOR U32990 ( .A(n32705), .B(n32704), .Z(n32703) );
  AND U32991 ( .A(n35559), .B(n35560), .Z(n32704) );
  XOR U32992 ( .A(n32707), .B(n32706), .Z(n32705) );
  AND U32993 ( .A(n35561), .B(n35562), .Z(n32706) );
  XOR U32994 ( .A(n32709), .B(n32708), .Z(n32707) );
  AND U32995 ( .A(n35563), .B(n35564), .Z(n32708) );
  XOR U32996 ( .A(n32711), .B(n32710), .Z(n32709) );
  AND U32997 ( .A(n35565), .B(n35566), .Z(n32710) );
  XOR U32998 ( .A(n32713), .B(n32712), .Z(n32711) );
  AND U32999 ( .A(n35567), .B(n35568), .Z(n32712) );
  XOR U33000 ( .A(n32715), .B(n32714), .Z(n32713) );
  AND U33001 ( .A(n35569), .B(n35570), .Z(n32714) );
  XOR U33002 ( .A(n32717), .B(n32716), .Z(n32715) );
  AND U33003 ( .A(n35571), .B(n35572), .Z(n32716) );
  XOR U33004 ( .A(n32719), .B(n32718), .Z(n32717) );
  AND U33005 ( .A(n35573), .B(n35574), .Z(n32718) );
  XOR U33006 ( .A(n32721), .B(n32720), .Z(n32719) );
  AND U33007 ( .A(n35575), .B(n35576), .Z(n32720) );
  XOR U33008 ( .A(n32723), .B(n32722), .Z(n32721) );
  AND U33009 ( .A(n35577), .B(n35578), .Z(n32722) );
  XOR U33010 ( .A(n32725), .B(n32724), .Z(n32723) );
  AND U33011 ( .A(n35579), .B(n35580), .Z(n32724) );
  XOR U33012 ( .A(n32727), .B(n32726), .Z(n32725) );
  AND U33013 ( .A(n35581), .B(n35582), .Z(n32726) );
  XOR U33014 ( .A(n32729), .B(n32728), .Z(n32727) );
  AND U33015 ( .A(n35583), .B(n35584), .Z(n32728) );
  XOR U33016 ( .A(n32731), .B(n32730), .Z(n32729) );
  AND U33017 ( .A(n35585), .B(n35586), .Z(n32730) );
  XOR U33018 ( .A(n32733), .B(n32732), .Z(n32731) );
  AND U33019 ( .A(n35587), .B(n35588), .Z(n32732) );
  XOR U33020 ( .A(n32735), .B(n32734), .Z(n32733) );
  AND U33021 ( .A(n35589), .B(n35590), .Z(n32734) );
  XOR U33022 ( .A(n32737), .B(n32736), .Z(n32735) );
  AND U33023 ( .A(n35591), .B(n35592), .Z(n32736) );
  XOR U33024 ( .A(n32739), .B(n32738), .Z(n32737) );
  AND U33025 ( .A(n35593), .B(n35594), .Z(n32738) );
  XOR U33026 ( .A(n32741), .B(n32740), .Z(n32739) );
  AND U33027 ( .A(n35595), .B(n35596), .Z(n32740) );
  XOR U33028 ( .A(n32743), .B(n32742), .Z(n32741) );
  AND U33029 ( .A(n35597), .B(n35598), .Z(n32742) );
  XOR U33030 ( .A(n32745), .B(n32744), .Z(n32743) );
  AND U33031 ( .A(n35599), .B(n35600), .Z(n32744) );
  XOR U33032 ( .A(n32747), .B(n32746), .Z(n32745) );
  AND U33033 ( .A(n35601), .B(n35602), .Z(n32746) );
  XOR U33034 ( .A(n32749), .B(n32748), .Z(n32747) );
  AND U33035 ( .A(n35603), .B(n35604), .Z(n32748) );
  XOR U33036 ( .A(n32751), .B(n32750), .Z(n32749) );
  AND U33037 ( .A(n35605), .B(n35606), .Z(n32750) );
  XOR U33038 ( .A(n32753), .B(n32752), .Z(n32751) );
  AND U33039 ( .A(n35607), .B(n35608), .Z(n32752) );
  XOR U33040 ( .A(n32755), .B(n32754), .Z(n32753) );
  AND U33041 ( .A(n35609), .B(n35610), .Z(n32754) );
  XOR U33042 ( .A(n32757), .B(n32756), .Z(n32755) );
  AND U33043 ( .A(n35611), .B(n35612), .Z(n32756) );
  XOR U33044 ( .A(n32759), .B(n32758), .Z(n32757) );
  AND U33045 ( .A(n35613), .B(n35614), .Z(n32758) );
  XOR U33046 ( .A(n32761), .B(n32760), .Z(n32759) );
  AND U33047 ( .A(n35615), .B(n35616), .Z(n32760) );
  XOR U33048 ( .A(n32763), .B(n32762), .Z(n32761) );
  AND U33049 ( .A(n35617), .B(n35618), .Z(n32762) );
  XOR U33050 ( .A(n32765), .B(n32764), .Z(n32763) );
  AND U33051 ( .A(n35619), .B(n35620), .Z(n32764) );
  XOR U33052 ( .A(n32767), .B(n32766), .Z(n32765) );
  AND U33053 ( .A(n35621), .B(n35622), .Z(n32766) );
  XOR U33054 ( .A(n32897), .B(n32768), .Z(n32767) );
  AND U33055 ( .A(n35623), .B(n35624), .Z(n32768) );
  XOR U33056 ( .A(n32900), .B(n32898), .Z(n32897) );
  AND U33057 ( .A(n35625), .B(n35626), .Z(n32898) );
  XOR U33058 ( .A(n32770), .B(n32901), .Z(n32900) );
  AND U33059 ( .A(n35627), .B(n35628), .Z(n32901) );
  XOR U33060 ( .A(n32772), .B(n32771), .Z(n32770) );
  AND U33061 ( .A(n35629), .B(n35630), .Z(n32771) );
  XOR U33062 ( .A(n32893), .B(n32773), .Z(n32772) );
  AND U33063 ( .A(n35631), .B(n35632), .Z(n32773) );
  XOR U33064 ( .A(n32895), .B(n32894), .Z(n32893) );
  AND U33065 ( .A(n35633), .B(n35634), .Z(n32894) );
  XOR U33066 ( .A(n32781), .B(n32896), .Z(n32895) );
  AND U33067 ( .A(n35635), .B(n35636), .Z(n32896) );
  XOR U33068 ( .A(n32777), .B(n32782), .Z(n32781) );
  AND U33069 ( .A(n35637), .B(n35638), .Z(n32782) );
  XOR U33070 ( .A(n32779), .B(n32778), .Z(n32777) );
  AND U33071 ( .A(n35639), .B(n35640), .Z(n32778) );
  XOR U33072 ( .A(n32891), .B(n32780), .Z(n32779) );
  AND U33073 ( .A(n35641), .B(n35642), .Z(n32780) );
  XNOR U33074 ( .A(n32800), .B(n32892), .Z(n32891) );
  AND U33075 ( .A(n35643), .B(n35644), .Z(n32892) );
  XOR U33076 ( .A(n32799), .B(n32791), .Z(n32800) );
  AND U33077 ( .A(n35645), .B(n35646), .Z(n32791) );
  XNOR U33078 ( .A(n32794), .B(n32790), .Z(n32799) );
  AND U33079 ( .A(n35647), .B(n35648), .Z(n32790) );
  XOR U33080 ( .A(n32820), .B(n32795), .Z(n32794) );
  AND U33081 ( .A(n35649), .B(n35650), .Z(n32795) );
  XNOR U33082 ( .A(n32811), .B(n32821), .Z(n32820) );
  AND U33083 ( .A(n35651), .B(n35652), .Z(n32821) );
  XOR U33084 ( .A(n32809), .B(n32810), .Z(n32811) );
  AND U33085 ( .A(n35653), .B(n35654), .Z(n32810) );
  XNOR U33086 ( .A(n32803), .B(n32808), .Z(n32809) );
  AND U33087 ( .A(n35655), .B(n35656), .Z(n32808) );
  XOR U33088 ( .A(n32822), .B(n32804), .Z(n32803) );
  AND U33089 ( .A(n35657), .B(n35658), .Z(n32804) );
  XNOR U33090 ( .A(n32888), .B(n32823), .Z(n32822) );
  AND U33091 ( .A(n35659), .B(n35660), .Z(n32823) );
  XOR U33092 ( .A(n32887), .B(n32879), .Z(n32888) );
  AND U33093 ( .A(n35661), .B(n35662), .Z(n32879) );
  XNOR U33094 ( .A(n32882), .B(n32878), .Z(n32887) );
  AND U33095 ( .A(n35663), .B(n35664), .Z(n32878) );
  XOR U33096 ( .A(n32826), .B(n32883), .Z(n32882) );
  AND U33097 ( .A(n35665), .B(n35666), .Z(n32883) );
  XNOR U33098 ( .A(n32875), .B(n32827), .Z(n32826) );
  AND U33099 ( .A(n35667), .B(n35668), .Z(n32827) );
  XOR U33100 ( .A(n32874), .B(n32866), .Z(n32875) );
  AND U33101 ( .A(n35669), .B(n35670), .Z(n32866) );
  XNOR U33102 ( .A(n32869), .B(n32865), .Z(n32874) );
  AND U33103 ( .A(n35671), .B(n35672), .Z(n32865) );
  XOR U33104 ( .A(n35673), .B(n35674), .Z(n32869) );
  XOR U33105 ( .A(n32859), .B(n32860), .Z(n35674) );
  AND U33106 ( .A(n35675), .B(n35676), .Z(n32860) );
  AND U33107 ( .A(n35677), .B(n35678), .Z(n32859) );
  XOR U33108 ( .A(n35679), .B(n32870), .Z(n35673) );
  AND U33109 ( .A(n35680), .B(n35681), .Z(n32870) );
  XOR U33110 ( .A(n35682), .B(n35683), .Z(n35679) );
  XOR U33111 ( .A(n35684), .B(n35685), .Z(n35683) );
  XOR U33112 ( .A(n32852), .B(n32853), .Z(n35685) );
  AND U33113 ( .A(n35686), .B(n35687), .Z(n32853) );
  AND U33114 ( .A(n35688), .B(n35689), .Z(n32852) );
  XOR U33115 ( .A(n32846), .B(n32851), .Z(n35684) );
  AND U33116 ( .A(n35690), .B(n35691), .Z(n32851) );
  AND U33117 ( .A(n35692), .B(n35693), .Z(n32846) );
  XOR U33118 ( .A(n35694), .B(n35695), .Z(n35682) );
  XOR U33119 ( .A(n32854), .B(n32857), .Z(n35695) );
  AND U33120 ( .A(n35696), .B(n35697), .Z(n32857) );
  AND U33121 ( .A(n35698), .B(n35699), .Z(n32854) );
  XOR U33122 ( .A(n35700), .B(n32858), .Z(n35694) );
  AND U33123 ( .A(n35701), .B(n35702), .Z(n32858) );
  XOR U33124 ( .A(n35703), .B(n35704), .Z(n35700) );
  XOR U33125 ( .A(n35705), .B(n35706), .Z(n35704) );
  XOR U33126 ( .A(n32839), .B(n32840), .Z(n35706) );
  AND U33127 ( .A(n35707), .B(n35708), .Z(n32840) );
  AND U33128 ( .A(n35709), .B(n35710), .Z(n32839) );
  XOR U33129 ( .A(n32837), .B(n32835), .Z(n35705) );
  AND U33130 ( .A(n35711), .B(n35712), .Z(n32835) );
  AND U33131 ( .A(n35713), .B(n35714), .Z(n32837) );
  XOR U33132 ( .A(n35715), .B(n35716), .Z(n35703) );
  XOR U33133 ( .A(n32843), .B(n32844), .Z(n35716) );
  AND U33134 ( .A(n35717), .B(n35718), .Z(n32844) );
  AND U33135 ( .A(n35719), .B(n35720), .Z(n32843) );
  XOR U33136 ( .A(n32838), .B(n32845), .Z(n35715) );
  AND U33137 ( .A(n35721), .B(n35722), .Z(n32845) );
  XOR U33138 ( .A(n35723), .B(n35724), .Z(n32838) );
  XOR U33139 ( .A(n35725), .B(n35726), .Z(n35724) );
  XOR U33140 ( .A(n35727), .B(n35728), .Z(n35726) );
  NOR U33141 ( .A(n35729), .B(n35730), .Z(n35728) );
  NOR U33142 ( .A(n35731), .B(n35732), .Z(n35727) );
  AND U33143 ( .A(n35733), .B(n35734), .Z(n35732) );
  IV U33144 ( .A(n35735), .Z(n35731) );
  NOR U33145 ( .A(n35736), .B(n35737), .Z(n35735) );
  AND U33146 ( .A(n35729), .B(n35738), .Z(n35737) );
  AND U33147 ( .A(n35730), .B(n35739), .Z(n35736) );
  XOR U33148 ( .A(n35740), .B(n35741), .Z(n35725) );
  NOR U33149 ( .A(n35742), .B(n35743), .Z(n35741) );
  NOR U33150 ( .A(n35744), .B(n35745), .Z(n35740) );
  AND U33151 ( .A(n35746), .B(n35747), .Z(n35745) );
  IV U33152 ( .A(n35748), .Z(n35744) );
  NOR U33153 ( .A(n35749), .B(n35750), .Z(n35748) );
  AND U33154 ( .A(n35742), .B(n35751), .Z(n35750) );
  AND U33155 ( .A(n35743), .B(n35752), .Z(n35749) );
  XOR U33156 ( .A(n35753), .B(n35754), .Z(n35723) );
  AND U33157 ( .A(n35755), .B(n35756), .Z(n35754) );
  XNOR U33158 ( .A(n35757), .B(n35758), .Z(n35753) );
  AND U33159 ( .A(n35759), .B(n35760), .Z(n35758) );
  AND U33160 ( .A(n35761), .B(n35762), .Z(n35757) );
  AND U33161 ( .A(n35763), .B(n35764), .Z(n35762) );
  NOR U33162 ( .A(n35765), .B(n35766), .Z(n35764) );
  IV U33163 ( .A(n35767), .Z(n35765) );
  NOR U33164 ( .A(n35768), .B(n35769), .Z(n35767) );
  NOR U33165 ( .A(n35770), .B(n35771), .Z(n35763) );
  AND U33166 ( .A(n35772), .B(n35773), .Z(n35761) );
  NOR U33167 ( .A(n35774), .B(n35775), .Z(n35773) );
  NOR U33168 ( .A(n35776), .B(n35777), .Z(n35772) );
  XOR U33169 ( .A(n35778), .B(n35779), .Z(n32917) );
  AND U33170 ( .A(n35778), .B(n35780), .Z(n35779) );
  XNOR U33171 ( .A(n35781), .B(n35782), .Z(n32920) );
  AND U33172 ( .A(n35781), .B(n35783), .Z(n35782) );
  IV U33173 ( .A(n32923), .Z(n35534) );
  XNOR U33174 ( .A(n35784), .B(n35785), .Z(n32923) );
  AND U33175 ( .A(n35784), .B(n35786), .Z(n35785) );
  XNOR U33176 ( .A(n35787), .B(n35788), .Z(n32926) );
  AND U33177 ( .A(n35787), .B(n35789), .Z(n35788) );
  XNOR U33178 ( .A(n35790), .B(n35791), .Z(n32929) );
  AND U33179 ( .A(n35792), .B(n35790), .Z(n35791) );
  XOR U33180 ( .A(n35793), .B(n35794), .Z(n32932) );
  NOR U33181 ( .A(n35795), .B(n35793), .Z(n35794) );
  XOR U33182 ( .A(n35796), .B(n35797), .Z(n32935) );
  NOR U33183 ( .A(n35798), .B(n35796), .Z(n35797) );
  XOR U33184 ( .A(n35799), .B(n35800), .Z(n32938) );
  NOR U33185 ( .A(n35801), .B(n35799), .Z(n35800) );
  XOR U33186 ( .A(n35802), .B(n35803), .Z(n32941) );
  NOR U33187 ( .A(n35804), .B(n35802), .Z(n35803) );
  XOR U33188 ( .A(n35805), .B(n35806), .Z(n32944) );
  NOR U33189 ( .A(n35807), .B(n35805), .Z(n35806) );
  XOR U33190 ( .A(n35808), .B(n35809), .Z(n32947) );
  NOR U33191 ( .A(n35810), .B(n35808), .Z(n35809) );
  XOR U33192 ( .A(n35811), .B(n35812), .Z(n32950) );
  NOR U33193 ( .A(n35813), .B(n35811), .Z(n35812) );
  XOR U33194 ( .A(n35814), .B(n35815), .Z(n32953) );
  NOR U33195 ( .A(n35816), .B(n35814), .Z(n35815) );
  XOR U33196 ( .A(n35817), .B(n35818), .Z(n32956) );
  NOR U33197 ( .A(n35819), .B(n35817), .Z(n35818) );
  XOR U33198 ( .A(n35820), .B(n35821), .Z(n32959) );
  NOR U33199 ( .A(n35822), .B(n35820), .Z(n35821) );
  XOR U33200 ( .A(n35823), .B(n35824), .Z(n32962) );
  NOR U33201 ( .A(n35825), .B(n35823), .Z(n35824) );
  XOR U33202 ( .A(n35826), .B(n35827), .Z(n32965) );
  NOR U33203 ( .A(n35828), .B(n35826), .Z(n35827) );
  XOR U33204 ( .A(n35829), .B(n35830), .Z(n32968) );
  NOR U33205 ( .A(n35831), .B(n35829), .Z(n35830) );
  XOR U33206 ( .A(n35832), .B(n35833), .Z(n32971) );
  NOR U33207 ( .A(n35834), .B(n35832), .Z(n35833) );
  XOR U33208 ( .A(n35835), .B(n35836), .Z(n32974) );
  NOR U33209 ( .A(n35837), .B(n35835), .Z(n35836) );
  XOR U33210 ( .A(n35838), .B(n35839), .Z(n32977) );
  NOR U33211 ( .A(n35840), .B(n35838), .Z(n35839) );
  XOR U33212 ( .A(n35841), .B(n35842), .Z(n32980) );
  NOR U33213 ( .A(n35843), .B(n35841), .Z(n35842) );
  XOR U33214 ( .A(n35844), .B(n35845), .Z(n32983) );
  NOR U33215 ( .A(n35846), .B(n35844), .Z(n35845) );
  XOR U33216 ( .A(n35847), .B(n35848), .Z(n32986) );
  NOR U33217 ( .A(n35849), .B(n35847), .Z(n35848) );
  XOR U33218 ( .A(n35850), .B(n35851), .Z(n32989) );
  NOR U33219 ( .A(n35852), .B(n35850), .Z(n35851) );
  XOR U33220 ( .A(n35853), .B(n35854), .Z(n32992) );
  NOR U33221 ( .A(n35855), .B(n35853), .Z(n35854) );
  XOR U33222 ( .A(n35856), .B(n35857), .Z(n32995) );
  NOR U33223 ( .A(n35858), .B(n35856), .Z(n35857) );
  XOR U33224 ( .A(n35859), .B(n35860), .Z(n32998) );
  NOR U33225 ( .A(n35861), .B(n35859), .Z(n35860) );
  XOR U33226 ( .A(n35862), .B(n35863), .Z(n33001) );
  NOR U33227 ( .A(n35864), .B(n35862), .Z(n35863) );
  XOR U33228 ( .A(n35865), .B(n35866), .Z(n33004) );
  NOR U33229 ( .A(n35867), .B(n35865), .Z(n35866) );
  XOR U33230 ( .A(n35868), .B(n35869), .Z(n33007) );
  NOR U33231 ( .A(n35870), .B(n35868), .Z(n35869) );
  XOR U33232 ( .A(n35871), .B(n35872), .Z(n33010) );
  NOR U33233 ( .A(n35873), .B(n35871), .Z(n35872) );
  XOR U33234 ( .A(n35874), .B(n35875), .Z(n33013) );
  NOR U33235 ( .A(n35876), .B(n35874), .Z(n35875) );
  XOR U33236 ( .A(n35877), .B(n35878), .Z(n33016) );
  NOR U33237 ( .A(n35879), .B(n35877), .Z(n35878) );
  XOR U33238 ( .A(n35880), .B(n35881), .Z(n33019) );
  NOR U33239 ( .A(n35882), .B(n35880), .Z(n35881) );
  XOR U33240 ( .A(n35883), .B(n35884), .Z(n33022) );
  NOR U33241 ( .A(n35885), .B(n35883), .Z(n35884) );
  XOR U33242 ( .A(n35886), .B(n35887), .Z(n33025) );
  NOR U33243 ( .A(n35888), .B(n35886), .Z(n35887) );
  XOR U33244 ( .A(n35889), .B(n35890), .Z(n33028) );
  NOR U33245 ( .A(n35891), .B(n35889), .Z(n35890) );
  XOR U33246 ( .A(n35892), .B(n35893), .Z(n33031) );
  NOR U33247 ( .A(n35894), .B(n35892), .Z(n35893) );
  XOR U33248 ( .A(n35895), .B(n35896), .Z(n33034) );
  NOR U33249 ( .A(n35897), .B(n35895), .Z(n35896) );
  XOR U33250 ( .A(n35898), .B(n35899), .Z(n33037) );
  NOR U33251 ( .A(n35900), .B(n35898), .Z(n35899) );
  XOR U33252 ( .A(n35901), .B(n35902), .Z(n33040) );
  NOR U33253 ( .A(n35903), .B(n35901), .Z(n35902) );
  XOR U33254 ( .A(n35904), .B(n35905), .Z(n33043) );
  NOR U33255 ( .A(n35906), .B(n35904), .Z(n35905) );
  XOR U33256 ( .A(n35907), .B(n35908), .Z(n33046) );
  NOR U33257 ( .A(n35909), .B(n35907), .Z(n35908) );
  XOR U33258 ( .A(n35910), .B(n35911), .Z(n33049) );
  NOR U33259 ( .A(n35912), .B(n35910), .Z(n35911) );
  XOR U33260 ( .A(n35913), .B(n35914), .Z(n33052) );
  NOR U33261 ( .A(n35915), .B(n35913), .Z(n35914) );
  XOR U33262 ( .A(n35916), .B(n35917), .Z(n33055) );
  NOR U33263 ( .A(n35918), .B(n35916), .Z(n35917) );
  XOR U33264 ( .A(n35919), .B(n35920), .Z(n33058) );
  NOR U33265 ( .A(n35921), .B(n35919), .Z(n35920) );
  XOR U33266 ( .A(n35922), .B(n35923), .Z(n33061) );
  NOR U33267 ( .A(n35924), .B(n35922), .Z(n35923) );
  XOR U33268 ( .A(n35925), .B(n35926), .Z(n33064) );
  NOR U33269 ( .A(n35927), .B(n35925), .Z(n35926) );
  XOR U33270 ( .A(n35928), .B(n35929), .Z(n33067) );
  NOR U33271 ( .A(n35930), .B(n35928), .Z(n35929) );
  XOR U33272 ( .A(n35931), .B(n35932), .Z(n33070) );
  NOR U33273 ( .A(n35933), .B(n35931), .Z(n35932) );
  XOR U33274 ( .A(n35934), .B(n35935), .Z(n33073) );
  NOR U33275 ( .A(n35936), .B(n35934), .Z(n35935) );
  XOR U33276 ( .A(n35937), .B(n35938), .Z(n33076) );
  NOR U33277 ( .A(n35939), .B(n35937), .Z(n35938) );
  XOR U33278 ( .A(n35940), .B(n35941), .Z(n33079) );
  NOR U33279 ( .A(n35942), .B(n35940), .Z(n35941) );
  XOR U33280 ( .A(n35943), .B(n35944), .Z(n33082) );
  NOR U33281 ( .A(n35945), .B(n35943), .Z(n35944) );
  XOR U33282 ( .A(n35946), .B(n35947), .Z(n33085) );
  NOR U33283 ( .A(n35948), .B(n35946), .Z(n35947) );
  XOR U33284 ( .A(n35949), .B(n35950), .Z(n33088) );
  NOR U33285 ( .A(n35951), .B(n35949), .Z(n35950) );
  XOR U33286 ( .A(n35952), .B(n35953), .Z(n33091) );
  NOR U33287 ( .A(n35954), .B(n35952), .Z(n35953) );
  XOR U33288 ( .A(n35955), .B(n35956), .Z(n33094) );
  NOR U33289 ( .A(n35957), .B(n35955), .Z(n35956) );
  XOR U33290 ( .A(n35958), .B(n35959), .Z(n33097) );
  NOR U33291 ( .A(n35960), .B(n35958), .Z(n35959) );
  XOR U33292 ( .A(n35961), .B(n35962), .Z(n33100) );
  NOR U33293 ( .A(n35963), .B(n35961), .Z(n35962) );
  XOR U33294 ( .A(n35964), .B(n35965), .Z(n33103) );
  NOR U33295 ( .A(n35966), .B(n35964), .Z(n35965) );
  XOR U33296 ( .A(n35967), .B(n35968), .Z(n33106) );
  NOR U33297 ( .A(n35969), .B(n35967), .Z(n35968) );
  XOR U33298 ( .A(n35970), .B(n35971), .Z(n33109) );
  NOR U33299 ( .A(n35972), .B(n35970), .Z(n35971) );
  XOR U33300 ( .A(n35973), .B(n35974), .Z(n33112) );
  NOR U33301 ( .A(n35975), .B(n35973), .Z(n35974) );
  XOR U33302 ( .A(n35976), .B(n35977), .Z(n33115) );
  NOR U33303 ( .A(n35978), .B(n35976), .Z(n35977) );
  XOR U33304 ( .A(n35979), .B(n35980), .Z(n33118) );
  NOR U33305 ( .A(n35981), .B(n35979), .Z(n35980) );
  XOR U33306 ( .A(n35982), .B(n35983), .Z(n33121) );
  NOR U33307 ( .A(n35984), .B(n35982), .Z(n35983) );
  XOR U33308 ( .A(n35985), .B(n35986), .Z(n33124) );
  NOR U33309 ( .A(n35987), .B(n35985), .Z(n35986) );
  XOR U33310 ( .A(n35988), .B(n35989), .Z(n33127) );
  NOR U33311 ( .A(n35990), .B(n35988), .Z(n35989) );
  XOR U33312 ( .A(n35991), .B(n35992), .Z(n33130) );
  NOR U33313 ( .A(n35993), .B(n35991), .Z(n35992) );
  XOR U33314 ( .A(n35994), .B(n35995), .Z(n33133) );
  NOR U33315 ( .A(n35996), .B(n35994), .Z(n35995) );
  XOR U33316 ( .A(n35997), .B(n35998), .Z(n33136) );
  NOR U33317 ( .A(n35999), .B(n35997), .Z(n35998) );
  XOR U33318 ( .A(n36000), .B(n36001), .Z(n33139) );
  NOR U33319 ( .A(n36002), .B(n36000), .Z(n36001) );
  XOR U33320 ( .A(n36003), .B(n36004), .Z(n33142) );
  NOR U33321 ( .A(n36005), .B(n36003), .Z(n36004) );
  XOR U33322 ( .A(n36006), .B(n36007), .Z(n33145) );
  NOR U33323 ( .A(n36008), .B(n36006), .Z(n36007) );
  XOR U33324 ( .A(n36009), .B(n36010), .Z(n33148) );
  NOR U33325 ( .A(n36011), .B(n36009), .Z(n36010) );
  XOR U33326 ( .A(n36012), .B(n36013), .Z(n33151) );
  NOR U33327 ( .A(n36014), .B(n36012), .Z(n36013) );
  XOR U33328 ( .A(n36015), .B(n36016), .Z(n33154) );
  NOR U33329 ( .A(n36017), .B(n36015), .Z(n36016) );
  XOR U33330 ( .A(n36018), .B(n36019), .Z(n33157) );
  NOR U33331 ( .A(n36020), .B(n36018), .Z(n36019) );
  XOR U33332 ( .A(n36021), .B(n36022), .Z(n33160) );
  NOR U33333 ( .A(n36023), .B(n36021), .Z(n36022) );
  XOR U33334 ( .A(n36024), .B(n36025), .Z(n33163) );
  NOR U33335 ( .A(n36026), .B(n36024), .Z(n36025) );
  XOR U33336 ( .A(n36027), .B(n36028), .Z(n33166) );
  NOR U33337 ( .A(n36029), .B(n36027), .Z(n36028) );
  XOR U33338 ( .A(n36030), .B(n36031), .Z(n33169) );
  NOR U33339 ( .A(n36032), .B(n36030), .Z(n36031) );
  XOR U33340 ( .A(n36033), .B(n36034), .Z(n33172) );
  NOR U33341 ( .A(n36035), .B(n36033), .Z(n36034) );
  XOR U33342 ( .A(n36036), .B(n36037), .Z(n33175) );
  NOR U33343 ( .A(n36038), .B(n36036), .Z(n36037) );
  XOR U33344 ( .A(n36039), .B(n36040), .Z(n33178) );
  NOR U33345 ( .A(n36041), .B(n36039), .Z(n36040) );
  XOR U33346 ( .A(n36042), .B(n36043), .Z(n33181) );
  NOR U33347 ( .A(n36044), .B(n36042), .Z(n36043) );
  XOR U33348 ( .A(n36045), .B(n36046), .Z(n33184) );
  NOR U33349 ( .A(n36047), .B(n36045), .Z(n36046) );
  XOR U33350 ( .A(n36048), .B(n36049), .Z(n33187) );
  NOR U33351 ( .A(n36050), .B(n36048), .Z(n36049) );
  XOR U33352 ( .A(n36051), .B(n36052), .Z(n33190) );
  NOR U33353 ( .A(n36053), .B(n36051), .Z(n36052) );
  XOR U33354 ( .A(n36054), .B(n36055), .Z(n33193) );
  NOR U33355 ( .A(n36056), .B(n36054), .Z(n36055) );
  XOR U33356 ( .A(n36057), .B(n36058), .Z(n33196) );
  NOR U33357 ( .A(n36059), .B(n36057), .Z(n36058) );
  XOR U33358 ( .A(n36060), .B(n36061), .Z(n33199) );
  NOR U33359 ( .A(n36062), .B(n36060), .Z(n36061) );
  XOR U33360 ( .A(n36063), .B(n36064), .Z(n33202) );
  NOR U33361 ( .A(n36065), .B(n36063), .Z(n36064) );
  XOR U33362 ( .A(n36066), .B(n36067), .Z(n33205) );
  NOR U33363 ( .A(n36068), .B(n36066), .Z(n36067) );
  XOR U33364 ( .A(n36069), .B(n36070), .Z(n33208) );
  NOR U33365 ( .A(n36071), .B(n36069), .Z(n36070) );
  XOR U33366 ( .A(n36072), .B(n36073), .Z(n33211) );
  NOR U33367 ( .A(n36074), .B(n36072), .Z(n36073) );
  XOR U33368 ( .A(n36075), .B(n36076), .Z(n33214) );
  NOR U33369 ( .A(n36077), .B(n36075), .Z(n36076) );
  XOR U33370 ( .A(n36078), .B(n36079), .Z(n33217) );
  NOR U33371 ( .A(n36080), .B(n36078), .Z(n36079) );
  XOR U33372 ( .A(n36081), .B(n36082), .Z(n33220) );
  NOR U33373 ( .A(n36083), .B(n36081), .Z(n36082) );
  XOR U33374 ( .A(n36084), .B(n36085), .Z(n33223) );
  NOR U33375 ( .A(n36086), .B(n36084), .Z(n36085) );
  XOR U33376 ( .A(n36087), .B(n36088), .Z(n33226) );
  NOR U33377 ( .A(n36089), .B(n36087), .Z(n36088) );
  XOR U33378 ( .A(n36090), .B(n36091), .Z(n33229) );
  NOR U33379 ( .A(n36092), .B(n36090), .Z(n36091) );
  XOR U33380 ( .A(n36093), .B(n36094), .Z(n33232) );
  NOR U33381 ( .A(n36095), .B(n36093), .Z(n36094) );
  XOR U33382 ( .A(n36096), .B(n36097), .Z(n33235) );
  NOR U33383 ( .A(n36098), .B(n36096), .Z(n36097) );
  XOR U33384 ( .A(n36099), .B(n36100), .Z(n33238) );
  NOR U33385 ( .A(n36101), .B(n36099), .Z(n36100) );
  XOR U33386 ( .A(n36102), .B(n36103), .Z(n33241) );
  NOR U33387 ( .A(n36104), .B(n36102), .Z(n36103) );
  XOR U33388 ( .A(n36105), .B(n36106), .Z(n33244) );
  NOR U33389 ( .A(n36107), .B(n36105), .Z(n36106) );
  XOR U33390 ( .A(n36108), .B(n36109), .Z(n33247) );
  NOR U33391 ( .A(n36110), .B(n36108), .Z(n36109) );
  XOR U33392 ( .A(n36111), .B(n36112), .Z(n33250) );
  NOR U33393 ( .A(n36113), .B(n36111), .Z(n36112) );
  XOR U33394 ( .A(n36114), .B(n36115), .Z(n33253) );
  NOR U33395 ( .A(n36116), .B(n36114), .Z(n36115) );
  XOR U33396 ( .A(n36117), .B(n36118), .Z(n33256) );
  NOR U33397 ( .A(n36119), .B(n36117), .Z(n36118) );
  XOR U33398 ( .A(n36120), .B(n36121), .Z(n33259) );
  NOR U33399 ( .A(n36122), .B(n36120), .Z(n36121) );
  XOR U33400 ( .A(n36123), .B(n36124), .Z(n33262) );
  NOR U33401 ( .A(n36125), .B(n36123), .Z(n36124) );
  XOR U33402 ( .A(n36126), .B(n36127), .Z(n33265) );
  NOR U33403 ( .A(n36128), .B(n36126), .Z(n36127) );
  XOR U33404 ( .A(n36129), .B(n36130), .Z(n33268) );
  NOR U33405 ( .A(n36131), .B(n36129), .Z(n36130) );
  XOR U33406 ( .A(n36132), .B(n36133), .Z(n33271) );
  NOR U33407 ( .A(n36134), .B(n36132), .Z(n36133) );
  XOR U33408 ( .A(n36135), .B(n36136), .Z(n33274) );
  NOR U33409 ( .A(n36137), .B(n36135), .Z(n36136) );
  XOR U33410 ( .A(n36138), .B(n36139), .Z(n33277) );
  NOR U33411 ( .A(n36140), .B(n36138), .Z(n36139) );
  XOR U33412 ( .A(n36141), .B(n36142), .Z(n33280) );
  NOR U33413 ( .A(n36143), .B(n36141), .Z(n36142) );
  XOR U33414 ( .A(n36144), .B(n36145), .Z(n33283) );
  NOR U33415 ( .A(n36146), .B(n36144), .Z(n36145) );
  XOR U33416 ( .A(n36147), .B(n36148), .Z(n33286) );
  NOR U33417 ( .A(n36149), .B(n36147), .Z(n36148) );
  XOR U33418 ( .A(n36150), .B(n36151), .Z(n33289) );
  NOR U33419 ( .A(n36152), .B(n36150), .Z(n36151) );
  XOR U33420 ( .A(n36153), .B(n36154), .Z(n33292) );
  NOR U33421 ( .A(n36155), .B(n36153), .Z(n36154) );
  XOR U33422 ( .A(n36156), .B(n36157), .Z(n33295) );
  NOR U33423 ( .A(n36158), .B(n36156), .Z(n36157) );
  XOR U33424 ( .A(n36159), .B(n36160), .Z(n33298) );
  NOR U33425 ( .A(n36161), .B(n36159), .Z(n36160) );
  XOR U33426 ( .A(n36162), .B(n36163), .Z(n33301) );
  NOR U33427 ( .A(n36164), .B(n36162), .Z(n36163) );
  XOR U33428 ( .A(n36165), .B(n36166), .Z(n33304) );
  NOR U33429 ( .A(n36167), .B(n36165), .Z(n36166) );
  XOR U33430 ( .A(n36168), .B(n36169), .Z(n33307) );
  NOR U33431 ( .A(n36170), .B(n36168), .Z(n36169) );
  XOR U33432 ( .A(n36171), .B(n36172), .Z(n33310) );
  NOR U33433 ( .A(n36173), .B(n36171), .Z(n36172) );
  XOR U33434 ( .A(n36174), .B(n36175), .Z(n33313) );
  NOR U33435 ( .A(n36176), .B(n36174), .Z(n36175) );
  XOR U33436 ( .A(n36177), .B(n36178), .Z(n33316) );
  NOR U33437 ( .A(n36179), .B(n36177), .Z(n36178) );
  XOR U33438 ( .A(n36180), .B(n36181), .Z(n33319) );
  NOR U33439 ( .A(n36182), .B(n36180), .Z(n36181) );
  XOR U33440 ( .A(n36183), .B(n36184), .Z(n33322) );
  NOR U33441 ( .A(n36185), .B(n36183), .Z(n36184) );
  XOR U33442 ( .A(n36186), .B(n36187), .Z(n33325) );
  NOR U33443 ( .A(n36188), .B(n36186), .Z(n36187) );
  XOR U33444 ( .A(n36189), .B(n36190), .Z(n33328) );
  NOR U33445 ( .A(n36191), .B(n36189), .Z(n36190) );
  XOR U33446 ( .A(n36192), .B(n36193), .Z(n33331) );
  NOR U33447 ( .A(n36194), .B(n36192), .Z(n36193) );
  XOR U33448 ( .A(n36195), .B(n36196), .Z(n33334) );
  NOR U33449 ( .A(n36197), .B(n36195), .Z(n36196) );
  XOR U33450 ( .A(n36198), .B(n36199), .Z(n33337) );
  NOR U33451 ( .A(n36200), .B(n36198), .Z(n36199) );
  XOR U33452 ( .A(n36201), .B(n36202), .Z(n33340) );
  NOR U33453 ( .A(n36203), .B(n36201), .Z(n36202) );
  XOR U33454 ( .A(n36204), .B(n36205), .Z(n33343) );
  NOR U33455 ( .A(n36206), .B(n36204), .Z(n36205) );
  XOR U33456 ( .A(n36207), .B(n36208), .Z(n33346) );
  NOR U33457 ( .A(n36209), .B(n36207), .Z(n36208) );
  XOR U33458 ( .A(n36210), .B(n36211), .Z(n33349) );
  NOR U33459 ( .A(n36212), .B(n36210), .Z(n36211) );
  XOR U33460 ( .A(n36213), .B(n36214), .Z(n33352) );
  NOR U33461 ( .A(n36215), .B(n36213), .Z(n36214) );
  XOR U33462 ( .A(n36216), .B(n36217), .Z(n33355) );
  NOR U33463 ( .A(n36218), .B(n36216), .Z(n36217) );
  XOR U33464 ( .A(n36219), .B(n36220), .Z(n33358) );
  NOR U33465 ( .A(n36221), .B(n36219), .Z(n36220) );
  XOR U33466 ( .A(n36222), .B(n36223), .Z(n33361) );
  NOR U33467 ( .A(n36224), .B(n36222), .Z(n36223) );
  XOR U33468 ( .A(n36225), .B(n36226), .Z(n33364) );
  NOR U33469 ( .A(n36227), .B(n36225), .Z(n36226) );
  XOR U33470 ( .A(n36228), .B(n36229), .Z(n33367) );
  NOR U33471 ( .A(n36230), .B(n36228), .Z(n36229) );
  XOR U33472 ( .A(n36231), .B(n36232), .Z(n33370) );
  NOR U33473 ( .A(n36233), .B(n36231), .Z(n36232) );
  XOR U33474 ( .A(n36234), .B(n36235), .Z(n33373) );
  NOR U33475 ( .A(n36236), .B(n36234), .Z(n36235) );
  XOR U33476 ( .A(n36237), .B(n36238), .Z(n33376) );
  NOR U33477 ( .A(n36239), .B(n36237), .Z(n36238) );
  XOR U33478 ( .A(n36240), .B(n36241), .Z(n33379) );
  NOR U33479 ( .A(n36242), .B(n36240), .Z(n36241) );
  XOR U33480 ( .A(n36243), .B(n36244), .Z(n33382) );
  NOR U33481 ( .A(n36245), .B(n36243), .Z(n36244) );
  XOR U33482 ( .A(n36246), .B(n36247), .Z(n33385) );
  NOR U33483 ( .A(n36248), .B(n36246), .Z(n36247) );
  XOR U33484 ( .A(n36249), .B(n36250), .Z(n33388) );
  NOR U33485 ( .A(n36251), .B(n36249), .Z(n36250) );
  XOR U33486 ( .A(n36252), .B(n36253), .Z(n33391) );
  NOR U33487 ( .A(n36254), .B(n36252), .Z(n36253) );
  XOR U33488 ( .A(n36255), .B(n36256), .Z(n33394) );
  NOR U33489 ( .A(n36257), .B(n36255), .Z(n36256) );
  XOR U33490 ( .A(n36258), .B(n36259), .Z(n33397) );
  NOR U33491 ( .A(n36260), .B(n36258), .Z(n36259) );
  XOR U33492 ( .A(n36261), .B(n36262), .Z(n33400) );
  NOR U33493 ( .A(n36263), .B(n36261), .Z(n36262) );
  XOR U33494 ( .A(n36264), .B(n36265), .Z(n33403) );
  NOR U33495 ( .A(n36266), .B(n36264), .Z(n36265) );
  XOR U33496 ( .A(n36267), .B(n36268), .Z(n33406) );
  NOR U33497 ( .A(n36269), .B(n36267), .Z(n36268) );
  XOR U33498 ( .A(n36270), .B(n36271), .Z(n33409) );
  NOR U33499 ( .A(n36272), .B(n36270), .Z(n36271) );
  XOR U33500 ( .A(n36273), .B(n36274), .Z(n33412) );
  NOR U33501 ( .A(n36275), .B(n36273), .Z(n36274) );
  XOR U33502 ( .A(n36276), .B(n36277), .Z(n33415) );
  NOR U33503 ( .A(n36278), .B(n36276), .Z(n36277) );
  XOR U33504 ( .A(n36279), .B(n36280), .Z(n33418) );
  NOR U33505 ( .A(n36281), .B(n36279), .Z(n36280) );
  XOR U33506 ( .A(n36282), .B(n36283), .Z(n33421) );
  NOR U33507 ( .A(n36284), .B(n36282), .Z(n36283) );
  XOR U33508 ( .A(n36285), .B(n36286), .Z(n33424) );
  NOR U33509 ( .A(n36287), .B(n36285), .Z(n36286) );
  XOR U33510 ( .A(n36288), .B(n36289), .Z(n33427) );
  NOR U33511 ( .A(n36290), .B(n36288), .Z(n36289) );
  XOR U33512 ( .A(n36291), .B(n36292), .Z(n33430) );
  NOR U33513 ( .A(n36293), .B(n36291), .Z(n36292) );
  XOR U33514 ( .A(n36294), .B(n36295), .Z(n33433) );
  NOR U33515 ( .A(n36296), .B(n36294), .Z(n36295) );
  XOR U33516 ( .A(n36297), .B(n36298), .Z(n33436) );
  NOR U33517 ( .A(n36299), .B(n36297), .Z(n36298) );
  XOR U33518 ( .A(n36300), .B(n36301), .Z(n33439) );
  NOR U33519 ( .A(n36302), .B(n36300), .Z(n36301) );
  XOR U33520 ( .A(n36303), .B(n36304), .Z(n33442) );
  NOR U33521 ( .A(n36305), .B(n36303), .Z(n36304) );
  XOR U33522 ( .A(n36306), .B(n36307), .Z(n33445) );
  NOR U33523 ( .A(n36308), .B(n36306), .Z(n36307) );
  XOR U33524 ( .A(n36309), .B(n36310), .Z(n33448) );
  NOR U33525 ( .A(n36311), .B(n36309), .Z(n36310) );
  XOR U33526 ( .A(n36312), .B(n36313), .Z(n33451) );
  NOR U33527 ( .A(n36314), .B(n36312), .Z(n36313) );
  XOR U33528 ( .A(n36315), .B(n36316), .Z(n33454) );
  NOR U33529 ( .A(n36317), .B(n36315), .Z(n36316) );
  XOR U33530 ( .A(n36318), .B(n36319), .Z(n33457) );
  NOR U33531 ( .A(n36320), .B(n36318), .Z(n36319) );
  XOR U33532 ( .A(n36321), .B(n36322), .Z(n33460) );
  NOR U33533 ( .A(n36323), .B(n36321), .Z(n36322) );
  XOR U33534 ( .A(n36324), .B(n36325), .Z(n33463) );
  NOR U33535 ( .A(n36326), .B(n36324), .Z(n36325) );
  XOR U33536 ( .A(n36327), .B(n36328), .Z(n33466) );
  NOR U33537 ( .A(n36329), .B(n36327), .Z(n36328) );
  XOR U33538 ( .A(n36330), .B(n36331), .Z(n33469) );
  NOR U33539 ( .A(n36332), .B(n36330), .Z(n36331) );
  XOR U33540 ( .A(n36333), .B(n36334), .Z(n33472) );
  NOR U33541 ( .A(n36335), .B(n36333), .Z(n36334) );
  XOR U33542 ( .A(n36336), .B(n36337), .Z(n33475) );
  NOR U33543 ( .A(n36338), .B(n36336), .Z(n36337) );
  XOR U33544 ( .A(n36339), .B(n36340), .Z(n33478) );
  NOR U33545 ( .A(n36341), .B(n36339), .Z(n36340) );
  XOR U33546 ( .A(n36342), .B(n36343), .Z(n33481) );
  NOR U33547 ( .A(n36344), .B(n36342), .Z(n36343) );
  XOR U33548 ( .A(n36345), .B(n36346), .Z(n33484) );
  NOR U33549 ( .A(n36347), .B(n36345), .Z(n36346) );
  XOR U33550 ( .A(n36348), .B(n36349), .Z(n33487) );
  NOR U33551 ( .A(n36350), .B(n36348), .Z(n36349) );
  XOR U33552 ( .A(n36351), .B(n36352), .Z(n33490) );
  NOR U33553 ( .A(n36353), .B(n36351), .Z(n36352) );
  XOR U33554 ( .A(n36354), .B(n36355), .Z(n33493) );
  NOR U33555 ( .A(n36356), .B(n36354), .Z(n36355) );
  XOR U33556 ( .A(n36357), .B(n36358), .Z(n33496) );
  NOR U33557 ( .A(n36359), .B(n36357), .Z(n36358) );
  XOR U33558 ( .A(n36360), .B(n36361), .Z(n33499) );
  NOR U33559 ( .A(n36362), .B(n36360), .Z(n36361) );
  XOR U33560 ( .A(n36363), .B(n36364), .Z(n33502) );
  NOR U33561 ( .A(n36365), .B(n36363), .Z(n36364) );
  XOR U33562 ( .A(n36366), .B(n36367), .Z(n33505) );
  NOR U33563 ( .A(n36368), .B(n36366), .Z(n36367) );
  XOR U33564 ( .A(n36369), .B(n36370), .Z(n33508) );
  NOR U33565 ( .A(n36371), .B(n36369), .Z(n36370) );
  XOR U33566 ( .A(n36372), .B(n36373), .Z(n33511) );
  NOR U33567 ( .A(n36374), .B(n36372), .Z(n36373) );
  XOR U33568 ( .A(n36375), .B(n36376), .Z(n33514) );
  NOR U33569 ( .A(n36377), .B(n36375), .Z(n36376) );
  XOR U33570 ( .A(n36378), .B(n36379), .Z(n33517) );
  NOR U33571 ( .A(n36380), .B(n36378), .Z(n36379) );
  XOR U33572 ( .A(n36381), .B(n36382), .Z(n33520) );
  NOR U33573 ( .A(n36383), .B(n36381), .Z(n36382) );
  XOR U33574 ( .A(n36384), .B(n36385), .Z(n33523) );
  NOR U33575 ( .A(n36386), .B(n36384), .Z(n36385) );
  XOR U33576 ( .A(n36387), .B(n36388), .Z(n33526) );
  NOR U33577 ( .A(n36389), .B(n36387), .Z(n36388) );
  XOR U33578 ( .A(n36390), .B(n36391), .Z(n33529) );
  NOR U33579 ( .A(n36392), .B(n36390), .Z(n36391) );
  XOR U33580 ( .A(n36393), .B(n36394), .Z(n33532) );
  NOR U33581 ( .A(n36395), .B(n36393), .Z(n36394) );
  XOR U33582 ( .A(n36396), .B(n36397), .Z(n33535) );
  NOR U33583 ( .A(n36398), .B(n36396), .Z(n36397) );
  XOR U33584 ( .A(n36399), .B(n36400), .Z(n33538) );
  NOR U33585 ( .A(n36401), .B(n36399), .Z(n36400) );
  XOR U33586 ( .A(n36402), .B(n36403), .Z(n33541) );
  NOR U33587 ( .A(n36404), .B(n36402), .Z(n36403) );
  XOR U33588 ( .A(n36405), .B(n36406), .Z(n33544) );
  NOR U33589 ( .A(n36407), .B(n36405), .Z(n36406) );
  XOR U33590 ( .A(n36408), .B(n36409), .Z(n33547) );
  NOR U33591 ( .A(n36410), .B(n36408), .Z(n36409) );
  XOR U33592 ( .A(n36411), .B(n36412), .Z(n33550) );
  NOR U33593 ( .A(n36413), .B(n36411), .Z(n36412) );
  XOR U33594 ( .A(n36414), .B(n36415), .Z(n33553) );
  NOR U33595 ( .A(n36416), .B(n36414), .Z(n36415) );
  XOR U33596 ( .A(n36417), .B(n36418), .Z(n33556) );
  NOR U33597 ( .A(n36419), .B(n36417), .Z(n36418) );
  XOR U33598 ( .A(n36420), .B(n36421), .Z(n33559) );
  NOR U33599 ( .A(n36422), .B(n36420), .Z(n36421) );
  XOR U33600 ( .A(n36423), .B(n36424), .Z(n33562) );
  NOR U33601 ( .A(n36425), .B(n36423), .Z(n36424) );
  XOR U33602 ( .A(n36426), .B(n36427), .Z(n33565) );
  NOR U33603 ( .A(n36428), .B(n36426), .Z(n36427) );
  XOR U33604 ( .A(n36429), .B(n36430), .Z(n33568) );
  NOR U33605 ( .A(n36431), .B(n36429), .Z(n36430) );
  XOR U33606 ( .A(n36432), .B(n36433), .Z(n33571) );
  NOR U33607 ( .A(n36434), .B(n36432), .Z(n36433) );
  XOR U33608 ( .A(n36435), .B(n36436), .Z(n33574) );
  NOR U33609 ( .A(n36437), .B(n36435), .Z(n36436) );
  XOR U33610 ( .A(n36438), .B(n36439), .Z(n33577) );
  NOR U33611 ( .A(n36440), .B(n36438), .Z(n36439) );
  XOR U33612 ( .A(n36441), .B(n36442), .Z(n33580) );
  NOR U33613 ( .A(n36443), .B(n36441), .Z(n36442) );
  XOR U33614 ( .A(n36444), .B(n36445), .Z(n33583) );
  NOR U33615 ( .A(n36446), .B(n36444), .Z(n36445) );
  XOR U33616 ( .A(n36447), .B(n36448), .Z(n33586) );
  NOR U33617 ( .A(n36449), .B(n36447), .Z(n36448) );
  XOR U33618 ( .A(n36450), .B(n36451), .Z(n33589) );
  NOR U33619 ( .A(n36452), .B(n36450), .Z(n36451) );
  XOR U33620 ( .A(n36453), .B(n36454), .Z(n33592) );
  NOR U33621 ( .A(n36455), .B(n36453), .Z(n36454) );
  XOR U33622 ( .A(n36456), .B(n36457), .Z(n33595) );
  NOR U33623 ( .A(n36458), .B(n36456), .Z(n36457) );
  XOR U33624 ( .A(n36459), .B(n36460), .Z(n33598) );
  NOR U33625 ( .A(n36461), .B(n36459), .Z(n36460) );
  XOR U33626 ( .A(n36462), .B(n36463), .Z(n33601) );
  NOR U33627 ( .A(n36464), .B(n36462), .Z(n36463) );
  XOR U33628 ( .A(n36465), .B(n36466), .Z(n33604) );
  NOR U33629 ( .A(n36467), .B(n36465), .Z(n36466) );
  XOR U33630 ( .A(n36468), .B(n36469), .Z(n33607) );
  NOR U33631 ( .A(n36470), .B(n36468), .Z(n36469) );
  XOR U33632 ( .A(n36471), .B(n36472), .Z(n33610) );
  NOR U33633 ( .A(n36473), .B(n36471), .Z(n36472) );
  XOR U33634 ( .A(n36474), .B(n36475), .Z(n33613) );
  NOR U33635 ( .A(n36476), .B(n36474), .Z(n36475) );
  XOR U33636 ( .A(n36477), .B(n36478), .Z(n33616) );
  NOR U33637 ( .A(n36479), .B(n36477), .Z(n36478) );
  XOR U33638 ( .A(n36480), .B(n36481), .Z(n33619) );
  NOR U33639 ( .A(n36482), .B(n36480), .Z(n36481) );
  XOR U33640 ( .A(n36483), .B(n36484), .Z(n33622) );
  NOR U33641 ( .A(n36485), .B(n36483), .Z(n36484) );
  XOR U33642 ( .A(n36486), .B(n36487), .Z(n33625) );
  NOR U33643 ( .A(n36488), .B(n36486), .Z(n36487) );
  XOR U33644 ( .A(n36489), .B(n36490), .Z(n33628) );
  NOR U33645 ( .A(n36491), .B(n36489), .Z(n36490) );
  XOR U33646 ( .A(n36492), .B(n36493), .Z(n33631) );
  NOR U33647 ( .A(n36494), .B(n36492), .Z(n36493) );
  XOR U33648 ( .A(n36495), .B(n36496), .Z(n33634) );
  NOR U33649 ( .A(n36497), .B(n36495), .Z(n36496) );
  XOR U33650 ( .A(n36498), .B(n36499), .Z(n33637) );
  NOR U33651 ( .A(n36500), .B(n36498), .Z(n36499) );
  XOR U33652 ( .A(n36501), .B(n36502), .Z(n33640) );
  NOR U33653 ( .A(n36503), .B(n36501), .Z(n36502) );
  XOR U33654 ( .A(n36504), .B(n36505), .Z(n33643) );
  NOR U33655 ( .A(n36506), .B(n36504), .Z(n36505) );
  XOR U33656 ( .A(n36507), .B(n36508), .Z(n33646) );
  NOR U33657 ( .A(n36509), .B(n36507), .Z(n36508) );
  XOR U33658 ( .A(n36510), .B(n36511), .Z(n33649) );
  NOR U33659 ( .A(n36512), .B(n36510), .Z(n36511) );
  XOR U33660 ( .A(n36513), .B(n36514), .Z(n33652) );
  NOR U33661 ( .A(n36515), .B(n36513), .Z(n36514) );
  XOR U33662 ( .A(n36516), .B(n36517), .Z(n33655) );
  NOR U33663 ( .A(n36518), .B(n36516), .Z(n36517) );
  XOR U33664 ( .A(n36519), .B(n36520), .Z(n33658) );
  NOR U33665 ( .A(n36521), .B(n36519), .Z(n36520) );
  XOR U33666 ( .A(n36522), .B(n36523), .Z(n33661) );
  NOR U33667 ( .A(n36524), .B(n36522), .Z(n36523) );
  XOR U33668 ( .A(n36525), .B(n36526), .Z(n33664) );
  NOR U33669 ( .A(n36527), .B(n36525), .Z(n36526) );
  XOR U33670 ( .A(n36528), .B(n36529), .Z(n33667) );
  NOR U33671 ( .A(n36530), .B(n36528), .Z(n36529) );
  XOR U33672 ( .A(n36531), .B(n36532), .Z(n33670) );
  NOR U33673 ( .A(n36533), .B(n36531), .Z(n36532) );
  XOR U33674 ( .A(n36534), .B(n36535), .Z(n33673) );
  NOR U33675 ( .A(n36536), .B(n36534), .Z(n36535) );
  XOR U33676 ( .A(n36537), .B(n36538), .Z(n33676) );
  NOR U33677 ( .A(n36539), .B(n36537), .Z(n36538) );
  XOR U33678 ( .A(n36540), .B(n36541), .Z(n33679) );
  NOR U33679 ( .A(n36542), .B(n36540), .Z(n36541) );
  XOR U33680 ( .A(n36543), .B(n36544), .Z(n33682) );
  NOR U33681 ( .A(n36545), .B(n36543), .Z(n36544) );
  XOR U33682 ( .A(n36546), .B(n36547), .Z(n33685) );
  NOR U33683 ( .A(n36548), .B(n36546), .Z(n36547) );
  XOR U33684 ( .A(n36549), .B(n36550), .Z(n33688) );
  NOR U33685 ( .A(n36551), .B(n36549), .Z(n36550) );
  XOR U33686 ( .A(n36552), .B(n36553), .Z(n33691) );
  NOR U33687 ( .A(n36554), .B(n36552), .Z(n36553) );
  XOR U33688 ( .A(n36555), .B(n36556), .Z(n33694) );
  NOR U33689 ( .A(n36557), .B(n36555), .Z(n36556) );
  XOR U33690 ( .A(n36558), .B(n36559), .Z(n33697) );
  NOR U33691 ( .A(n36560), .B(n36558), .Z(n36559) );
  XOR U33692 ( .A(n36561), .B(n36562), .Z(n33700) );
  NOR U33693 ( .A(n36563), .B(n36561), .Z(n36562) );
  XOR U33694 ( .A(n36564), .B(n36565), .Z(n33703) );
  NOR U33695 ( .A(n36566), .B(n36564), .Z(n36565) );
  XOR U33696 ( .A(n36567), .B(n36568), .Z(n33706) );
  NOR U33697 ( .A(n36569), .B(n36567), .Z(n36568) );
  XOR U33698 ( .A(n36570), .B(n36571), .Z(n33709) );
  NOR U33699 ( .A(n36572), .B(n36570), .Z(n36571) );
  XOR U33700 ( .A(n36573), .B(n36574), .Z(n33712) );
  NOR U33701 ( .A(n36575), .B(n36573), .Z(n36574) );
  XOR U33702 ( .A(n36576), .B(n36577), .Z(n33715) );
  NOR U33703 ( .A(n36578), .B(n36576), .Z(n36577) );
  XOR U33704 ( .A(n36579), .B(n36580), .Z(n33718) );
  NOR U33705 ( .A(n36581), .B(n36579), .Z(n36580) );
  XOR U33706 ( .A(n36582), .B(n36583), .Z(n33721) );
  NOR U33707 ( .A(n36584), .B(n36582), .Z(n36583) );
  XOR U33708 ( .A(n36585), .B(n36586), .Z(n33724) );
  NOR U33709 ( .A(n36587), .B(n36585), .Z(n36586) );
  XOR U33710 ( .A(n36588), .B(n36589), .Z(n33727) );
  NOR U33711 ( .A(n36590), .B(n36588), .Z(n36589) );
  XOR U33712 ( .A(n36591), .B(n36592), .Z(n33730) );
  NOR U33713 ( .A(n36593), .B(n36591), .Z(n36592) );
  XOR U33714 ( .A(n36594), .B(n36595), .Z(n33733) );
  NOR U33715 ( .A(n36596), .B(n36594), .Z(n36595) );
  XOR U33716 ( .A(n36597), .B(n36598), .Z(n33736) );
  NOR U33717 ( .A(n36599), .B(n36597), .Z(n36598) );
  XOR U33718 ( .A(n36600), .B(n36601), .Z(n33739) );
  NOR U33719 ( .A(n36602), .B(n36600), .Z(n36601) );
  XOR U33720 ( .A(n36603), .B(n36604), .Z(n33742) );
  NOR U33721 ( .A(n36605), .B(n36603), .Z(n36604) );
  XOR U33722 ( .A(n36606), .B(n36607), .Z(n33745) );
  NOR U33723 ( .A(n36608), .B(n36606), .Z(n36607) );
  XOR U33724 ( .A(n36609), .B(n36610), .Z(n33748) );
  NOR U33725 ( .A(n36611), .B(n36609), .Z(n36610) );
  XOR U33726 ( .A(n36612), .B(n36613), .Z(n33751) );
  NOR U33727 ( .A(n36614), .B(n36612), .Z(n36613) );
  XOR U33728 ( .A(n36615), .B(n36616), .Z(n33754) );
  NOR U33729 ( .A(n36617), .B(n36615), .Z(n36616) );
  XOR U33730 ( .A(n36618), .B(n36619), .Z(n33757) );
  NOR U33731 ( .A(n36620), .B(n36618), .Z(n36619) );
  XOR U33732 ( .A(n36621), .B(n36622), .Z(n33760) );
  NOR U33733 ( .A(n36623), .B(n36621), .Z(n36622) );
  XOR U33734 ( .A(n36624), .B(n36625), .Z(n33763) );
  NOR U33735 ( .A(n36626), .B(n36624), .Z(n36625) );
  XOR U33736 ( .A(n36627), .B(n36628), .Z(n33766) );
  NOR U33737 ( .A(n36629), .B(n36627), .Z(n36628) );
  XOR U33738 ( .A(n36630), .B(n36631), .Z(n33769) );
  NOR U33739 ( .A(n36632), .B(n36630), .Z(n36631) );
  XOR U33740 ( .A(n36633), .B(n36634), .Z(n33772) );
  NOR U33741 ( .A(n36635), .B(n36633), .Z(n36634) );
  XOR U33742 ( .A(n36636), .B(n36637), .Z(n33775) );
  NOR U33743 ( .A(n36638), .B(n36636), .Z(n36637) );
  XOR U33744 ( .A(n36639), .B(n36640), .Z(n33778) );
  NOR U33745 ( .A(n36641), .B(n36639), .Z(n36640) );
  XOR U33746 ( .A(n36642), .B(n36643), .Z(n33781) );
  NOR U33747 ( .A(n36644), .B(n36642), .Z(n36643) );
  XOR U33748 ( .A(n36645), .B(n36646), .Z(n33784) );
  NOR U33749 ( .A(n36647), .B(n36645), .Z(n36646) );
  XOR U33750 ( .A(n36648), .B(n36649), .Z(n33787) );
  NOR U33751 ( .A(n36650), .B(n36648), .Z(n36649) );
  XOR U33752 ( .A(n36651), .B(n36652), .Z(n33790) );
  NOR U33753 ( .A(n36653), .B(n36651), .Z(n36652) );
  XOR U33754 ( .A(n36654), .B(n36655), .Z(n33793) );
  NOR U33755 ( .A(n36656), .B(n36654), .Z(n36655) );
  XOR U33756 ( .A(n36657), .B(n36658), .Z(n33796) );
  NOR U33757 ( .A(n36659), .B(n36657), .Z(n36658) );
  XOR U33758 ( .A(n36660), .B(n36661), .Z(n33799) );
  NOR U33759 ( .A(n36662), .B(n36660), .Z(n36661) );
  XOR U33760 ( .A(n36663), .B(n36664), .Z(n33802) );
  NOR U33761 ( .A(n36665), .B(n36663), .Z(n36664) );
  XOR U33762 ( .A(n36666), .B(n36667), .Z(n33805) );
  NOR U33763 ( .A(n36668), .B(n36666), .Z(n36667) );
  XOR U33764 ( .A(n36669), .B(n36670), .Z(n33808) );
  NOR U33765 ( .A(n36671), .B(n36669), .Z(n36670) );
  XOR U33766 ( .A(n36672), .B(n36673), .Z(n33811) );
  NOR U33767 ( .A(n36674), .B(n36672), .Z(n36673) );
  XOR U33768 ( .A(n36675), .B(n36676), .Z(n33814) );
  NOR U33769 ( .A(n36677), .B(n36675), .Z(n36676) );
  XOR U33770 ( .A(n36678), .B(n36679), .Z(n33817) );
  NOR U33771 ( .A(n36680), .B(n36678), .Z(n36679) );
  XOR U33772 ( .A(n36681), .B(n36682), .Z(n33820) );
  NOR U33773 ( .A(n36683), .B(n36681), .Z(n36682) );
  XOR U33774 ( .A(n36684), .B(n36685), .Z(n33823) );
  NOR U33775 ( .A(n36686), .B(n36684), .Z(n36685) );
  XOR U33776 ( .A(n36687), .B(n36688), .Z(n33826) );
  NOR U33777 ( .A(n36689), .B(n36687), .Z(n36688) );
  XOR U33778 ( .A(n36690), .B(n36691), .Z(n33829) );
  NOR U33779 ( .A(n36692), .B(n36690), .Z(n36691) );
  XOR U33780 ( .A(n36693), .B(n36694), .Z(n33832) );
  NOR U33781 ( .A(n36695), .B(n36693), .Z(n36694) );
  XOR U33782 ( .A(n36696), .B(n36697), .Z(n33835) );
  NOR U33783 ( .A(n36698), .B(n36696), .Z(n36697) );
  XOR U33784 ( .A(n36699), .B(n36700), .Z(n33838) );
  NOR U33785 ( .A(n36701), .B(n36699), .Z(n36700) );
  XOR U33786 ( .A(n36702), .B(n36703), .Z(n33841) );
  NOR U33787 ( .A(n36704), .B(n36702), .Z(n36703) );
  XOR U33788 ( .A(n36705), .B(n36706), .Z(n33844) );
  NOR U33789 ( .A(n36707), .B(n36705), .Z(n36706) );
  XOR U33790 ( .A(n36708), .B(n36709), .Z(n33847) );
  NOR U33791 ( .A(n36710), .B(n36708), .Z(n36709) );
  XOR U33792 ( .A(n36711), .B(n36712), .Z(n33850) );
  NOR U33793 ( .A(n36713), .B(n36711), .Z(n36712) );
  XOR U33794 ( .A(n36714), .B(n36715), .Z(n33853) );
  NOR U33795 ( .A(n36716), .B(n36714), .Z(n36715) );
  XOR U33796 ( .A(n36717), .B(n36718), .Z(n33856) );
  NOR U33797 ( .A(n36719), .B(n36717), .Z(n36718) );
  XOR U33798 ( .A(n36720), .B(n36721), .Z(n33859) );
  NOR U33799 ( .A(n36722), .B(n36720), .Z(n36721) );
  XOR U33800 ( .A(n36723), .B(n36724), .Z(n33862) );
  NOR U33801 ( .A(n36725), .B(n36723), .Z(n36724) );
  XOR U33802 ( .A(n36726), .B(n36727), .Z(n33865) );
  NOR U33803 ( .A(n36728), .B(n36726), .Z(n36727) );
  XOR U33804 ( .A(n36729), .B(n36730), .Z(n33868) );
  NOR U33805 ( .A(n36731), .B(n36729), .Z(n36730) );
  XOR U33806 ( .A(n36732), .B(n36733), .Z(n33871) );
  NOR U33807 ( .A(n36734), .B(n36732), .Z(n36733) );
  XOR U33808 ( .A(n36735), .B(n36736), .Z(n33874) );
  NOR U33809 ( .A(n36737), .B(n36735), .Z(n36736) );
  XOR U33810 ( .A(n36738), .B(n36739), .Z(n33877) );
  NOR U33811 ( .A(n36740), .B(n36738), .Z(n36739) );
  XOR U33812 ( .A(n36741), .B(n36742), .Z(n33880) );
  NOR U33813 ( .A(n36743), .B(n36741), .Z(n36742) );
  XOR U33814 ( .A(n36744), .B(n36745), .Z(n33883) );
  NOR U33815 ( .A(n36746), .B(n36744), .Z(n36745) );
  XOR U33816 ( .A(n36747), .B(n36748), .Z(n33886) );
  NOR U33817 ( .A(n36749), .B(n36747), .Z(n36748) );
  XOR U33818 ( .A(n36750), .B(n36751), .Z(n33889) );
  NOR U33819 ( .A(n36752), .B(n36750), .Z(n36751) );
  XOR U33820 ( .A(n36753), .B(n36754), .Z(n33892) );
  NOR U33821 ( .A(n36755), .B(n36753), .Z(n36754) );
  XOR U33822 ( .A(n36756), .B(n36757), .Z(n33895) );
  NOR U33823 ( .A(n36758), .B(n36756), .Z(n36757) );
  XOR U33824 ( .A(n36759), .B(n36760), .Z(n33898) );
  NOR U33825 ( .A(n36761), .B(n36759), .Z(n36760) );
  XOR U33826 ( .A(n36762), .B(n36763), .Z(n33901) );
  NOR U33827 ( .A(n36764), .B(n36762), .Z(n36763) );
  XOR U33828 ( .A(n36765), .B(n36766), .Z(n33904) );
  NOR U33829 ( .A(n36767), .B(n36765), .Z(n36766) );
  XOR U33830 ( .A(n36768), .B(n36769), .Z(n33907) );
  NOR U33831 ( .A(n36770), .B(n36768), .Z(n36769) );
  XOR U33832 ( .A(n36771), .B(n36772), .Z(n33910) );
  NOR U33833 ( .A(n36773), .B(n36771), .Z(n36772) );
  XOR U33834 ( .A(n36774), .B(n36775), .Z(n33913) );
  NOR U33835 ( .A(n36776), .B(n36774), .Z(n36775) );
  XOR U33836 ( .A(n36777), .B(n36778), .Z(n33916) );
  NOR U33837 ( .A(n36779), .B(n36777), .Z(n36778) );
  XOR U33838 ( .A(n36780), .B(n36781), .Z(n33919) );
  NOR U33839 ( .A(n36782), .B(n36780), .Z(n36781) );
  XOR U33840 ( .A(n36783), .B(n36784), .Z(n33922) );
  NOR U33841 ( .A(n36785), .B(n36783), .Z(n36784) );
  XOR U33842 ( .A(n36786), .B(n36787), .Z(n33925) );
  NOR U33843 ( .A(n36788), .B(n36786), .Z(n36787) );
  XOR U33844 ( .A(n36789), .B(n36790), .Z(n33928) );
  NOR U33845 ( .A(n36791), .B(n36789), .Z(n36790) );
  XOR U33846 ( .A(n36792), .B(n36793), .Z(n33931) );
  NOR U33847 ( .A(n36794), .B(n36792), .Z(n36793) );
  XOR U33848 ( .A(n36795), .B(n36796), .Z(n33934) );
  NOR U33849 ( .A(n36797), .B(n36795), .Z(n36796) );
  XOR U33850 ( .A(n36798), .B(n36799), .Z(n33937) );
  NOR U33851 ( .A(n36800), .B(n36798), .Z(n36799) );
  XOR U33852 ( .A(n36801), .B(n36802), .Z(n33940) );
  NOR U33853 ( .A(n36803), .B(n36801), .Z(n36802) );
  XOR U33854 ( .A(n36804), .B(n36805), .Z(n33943) );
  NOR U33855 ( .A(n36806), .B(n36804), .Z(n36805) );
  XOR U33856 ( .A(n36807), .B(n36808), .Z(n33946) );
  NOR U33857 ( .A(n36809), .B(n36807), .Z(n36808) );
  XOR U33858 ( .A(n36810), .B(n36811), .Z(n33949) );
  NOR U33859 ( .A(n36812), .B(n36810), .Z(n36811) );
  XOR U33860 ( .A(n36813), .B(n36814), .Z(n33952) );
  NOR U33861 ( .A(n36815), .B(n36813), .Z(n36814) );
  XOR U33862 ( .A(n36816), .B(n36817), .Z(n33955) );
  NOR U33863 ( .A(n36818), .B(n36816), .Z(n36817) );
  XOR U33864 ( .A(n36819), .B(n36820), .Z(n33958) );
  NOR U33865 ( .A(n36821), .B(n36819), .Z(n36820) );
  XOR U33866 ( .A(n36822), .B(n36823), .Z(n33961) );
  NOR U33867 ( .A(n36824), .B(n36822), .Z(n36823) );
  XOR U33868 ( .A(n36825), .B(n36826), .Z(n33964) );
  NOR U33869 ( .A(n36827), .B(n36825), .Z(n36826) );
  XOR U33870 ( .A(n36828), .B(n36829), .Z(n33967) );
  NOR U33871 ( .A(n36830), .B(n36828), .Z(n36829) );
  XOR U33872 ( .A(n36831), .B(n36832), .Z(n33970) );
  NOR U33873 ( .A(n36833), .B(n36831), .Z(n36832) );
  XOR U33874 ( .A(n36834), .B(n36835), .Z(n33973) );
  NOR U33875 ( .A(n36836), .B(n36834), .Z(n36835) );
  XOR U33876 ( .A(n36837), .B(n36838), .Z(n33976) );
  NOR U33877 ( .A(n36839), .B(n36837), .Z(n36838) );
  XOR U33878 ( .A(n36840), .B(n36841), .Z(n33979) );
  NOR U33879 ( .A(n36842), .B(n36840), .Z(n36841) );
  XOR U33880 ( .A(n36843), .B(n36844), .Z(n33982) );
  NOR U33881 ( .A(n36845), .B(n36843), .Z(n36844) );
  XOR U33882 ( .A(n36846), .B(n36847), .Z(n33985) );
  NOR U33883 ( .A(n36848), .B(n36846), .Z(n36847) );
  XOR U33884 ( .A(n36849), .B(n36850), .Z(n33988) );
  NOR U33885 ( .A(n36851), .B(n36849), .Z(n36850) );
  XOR U33886 ( .A(n36852), .B(n36853), .Z(n33991) );
  NOR U33887 ( .A(n36854), .B(n36852), .Z(n36853) );
  XOR U33888 ( .A(n36855), .B(n36856), .Z(n33994) );
  NOR U33889 ( .A(n36857), .B(n36855), .Z(n36856) );
  XOR U33890 ( .A(n36858), .B(n36859), .Z(n33997) );
  NOR U33891 ( .A(n36860), .B(n36858), .Z(n36859) );
  XOR U33892 ( .A(n36861), .B(n36862), .Z(n34000) );
  NOR U33893 ( .A(n36863), .B(n36861), .Z(n36862) );
  XOR U33894 ( .A(n36864), .B(n36865), .Z(n34003) );
  NOR U33895 ( .A(n36866), .B(n36864), .Z(n36865) );
  XOR U33896 ( .A(n36867), .B(n36868), .Z(n34006) );
  NOR U33897 ( .A(n36869), .B(n36867), .Z(n36868) );
  XOR U33898 ( .A(n36870), .B(n36871), .Z(n34009) );
  NOR U33899 ( .A(n36872), .B(n36870), .Z(n36871) );
  XOR U33900 ( .A(n36873), .B(n36874), .Z(n34012) );
  NOR U33901 ( .A(n36875), .B(n36873), .Z(n36874) );
  XOR U33902 ( .A(n36876), .B(n36877), .Z(n34015) );
  NOR U33903 ( .A(n36878), .B(n36876), .Z(n36877) );
  XOR U33904 ( .A(n36879), .B(n36880), .Z(n34018) );
  NOR U33905 ( .A(n36881), .B(n36879), .Z(n36880) );
  XOR U33906 ( .A(n36882), .B(n36883), .Z(n34021) );
  NOR U33907 ( .A(n36884), .B(n36882), .Z(n36883) );
  XOR U33908 ( .A(n36885), .B(n36886), .Z(n34024) );
  NOR U33909 ( .A(n36887), .B(n36885), .Z(n36886) );
  XOR U33910 ( .A(n36888), .B(n36889), .Z(n34027) );
  NOR U33911 ( .A(n36890), .B(n36888), .Z(n36889) );
  XOR U33912 ( .A(n36891), .B(n36892), .Z(n34030) );
  NOR U33913 ( .A(n36893), .B(n36891), .Z(n36892) );
  XOR U33914 ( .A(n36894), .B(n36895), .Z(n34033) );
  NOR U33915 ( .A(n36896), .B(n36894), .Z(n36895) );
  XOR U33916 ( .A(n36897), .B(n36898), .Z(n34036) );
  NOR U33917 ( .A(n36899), .B(n36897), .Z(n36898) );
  XOR U33918 ( .A(n36900), .B(n36901), .Z(n34039) );
  NOR U33919 ( .A(n36902), .B(n36900), .Z(n36901) );
  XOR U33920 ( .A(n36903), .B(n36904), .Z(n34042) );
  NOR U33921 ( .A(n36905), .B(n36903), .Z(n36904) );
  XOR U33922 ( .A(n36906), .B(n36907), .Z(n34045) );
  NOR U33923 ( .A(n36908), .B(n36906), .Z(n36907) );
  XOR U33924 ( .A(n36909), .B(n36910), .Z(n34048) );
  NOR U33925 ( .A(n36911), .B(n36909), .Z(n36910) );
  XOR U33926 ( .A(n36912), .B(n36913), .Z(n34051) );
  NOR U33927 ( .A(n36914), .B(n36912), .Z(n36913) );
  XOR U33928 ( .A(n36915), .B(n36916), .Z(n34054) );
  NOR U33929 ( .A(n36917), .B(n36915), .Z(n36916) );
  XOR U33930 ( .A(n36918), .B(n36919), .Z(n34057) );
  NOR U33931 ( .A(n36920), .B(n36918), .Z(n36919) );
  XOR U33932 ( .A(n36921), .B(n36922), .Z(n34060) );
  NOR U33933 ( .A(n36923), .B(n36921), .Z(n36922) );
  XOR U33934 ( .A(n36924), .B(n36925), .Z(n34063) );
  NOR U33935 ( .A(n36926), .B(n36924), .Z(n36925) );
  XOR U33936 ( .A(n36927), .B(n36928), .Z(n34066) );
  NOR U33937 ( .A(n36929), .B(n36927), .Z(n36928) );
  XOR U33938 ( .A(n36930), .B(n36931), .Z(n34069) );
  NOR U33939 ( .A(n36932), .B(n36930), .Z(n36931) );
  XOR U33940 ( .A(n36933), .B(n36934), .Z(n34072) );
  NOR U33941 ( .A(n36935), .B(n36933), .Z(n36934) );
  XOR U33942 ( .A(n36936), .B(n36937), .Z(n34075) );
  NOR U33943 ( .A(n36938), .B(n36936), .Z(n36937) );
  XOR U33944 ( .A(n36939), .B(n36940), .Z(n34078) );
  NOR U33945 ( .A(n36941), .B(n36939), .Z(n36940) );
  XOR U33946 ( .A(n36942), .B(n36943), .Z(n34081) );
  NOR U33947 ( .A(n36944), .B(n36942), .Z(n36943) );
  XOR U33948 ( .A(n36945), .B(n36946), .Z(n34084) );
  NOR U33949 ( .A(n36947), .B(n36945), .Z(n36946) );
  XOR U33950 ( .A(n36948), .B(n36949), .Z(n34087) );
  NOR U33951 ( .A(n36950), .B(n36948), .Z(n36949) );
  XOR U33952 ( .A(n36951), .B(n36952), .Z(n34090) );
  NOR U33953 ( .A(n36953), .B(n36951), .Z(n36952) );
  XOR U33954 ( .A(n36954), .B(n36955), .Z(n34093) );
  NOR U33955 ( .A(n36956), .B(n36954), .Z(n36955) );
  XOR U33956 ( .A(n36957), .B(n36958), .Z(n34096) );
  NOR U33957 ( .A(n36959), .B(n36957), .Z(n36958) );
  XOR U33958 ( .A(n36960), .B(n36961), .Z(n34099) );
  NOR U33959 ( .A(n106), .B(n36962), .Z(n36961) );
  IV U33960 ( .A(n36960), .Z(n36962) );
  XOR U33961 ( .A(n36963), .B(n36964), .Z(n34102) );
  AND U33962 ( .A(n36965), .B(n36966), .Z(n36964) );
  XOR U33963 ( .A(n36963), .B(n109), .Z(n36966) );
  XOR U33964 ( .A(n35532), .B(n35531), .Z(n109) );
  XNOR U33965 ( .A(n35529), .B(n35528), .Z(n35531) );
  XNOR U33966 ( .A(n35526), .B(n35525), .Z(n35528) );
  XNOR U33967 ( .A(n35523), .B(n35522), .Z(n35525) );
  XNOR U33968 ( .A(n35520), .B(n35519), .Z(n35522) );
  XNOR U33969 ( .A(n35517), .B(n35516), .Z(n35519) );
  XNOR U33970 ( .A(n35514), .B(n35513), .Z(n35516) );
  XNOR U33971 ( .A(n35511), .B(n35510), .Z(n35513) );
  XNOR U33972 ( .A(n35508), .B(n35507), .Z(n35510) );
  XNOR U33973 ( .A(n35505), .B(n35504), .Z(n35507) );
  XNOR U33974 ( .A(n35502), .B(n35501), .Z(n35504) );
  XNOR U33975 ( .A(n35499), .B(n35498), .Z(n35501) );
  XNOR U33976 ( .A(n35496), .B(n35495), .Z(n35498) );
  XNOR U33977 ( .A(n35493), .B(n35492), .Z(n35495) );
  XNOR U33978 ( .A(n35490), .B(n35489), .Z(n35492) );
  XNOR U33979 ( .A(n35487), .B(n35486), .Z(n35489) );
  XNOR U33980 ( .A(n35484), .B(n35483), .Z(n35486) );
  XNOR U33981 ( .A(n35481), .B(n35480), .Z(n35483) );
  XNOR U33982 ( .A(n35478), .B(n35477), .Z(n35480) );
  XNOR U33983 ( .A(n35475), .B(n35474), .Z(n35477) );
  XNOR U33984 ( .A(n35472), .B(n35471), .Z(n35474) );
  XNOR U33985 ( .A(n35469), .B(n35468), .Z(n35471) );
  XNOR U33986 ( .A(n35466), .B(n35465), .Z(n35468) );
  XNOR U33987 ( .A(n35463), .B(n35462), .Z(n35465) );
  XNOR U33988 ( .A(n35460), .B(n35459), .Z(n35462) );
  XNOR U33989 ( .A(n35457), .B(n35456), .Z(n35459) );
  XNOR U33990 ( .A(n35454), .B(n35453), .Z(n35456) );
  XNOR U33991 ( .A(n35451), .B(n35450), .Z(n35453) );
  XNOR U33992 ( .A(n35448), .B(n35447), .Z(n35450) );
  XNOR U33993 ( .A(n35445), .B(n35444), .Z(n35447) );
  XNOR U33994 ( .A(n35442), .B(n35441), .Z(n35444) );
  XNOR U33995 ( .A(n35439), .B(n35438), .Z(n35441) );
  XNOR U33996 ( .A(n35436), .B(n35435), .Z(n35438) );
  XNOR U33997 ( .A(n35433), .B(n35432), .Z(n35435) );
  XNOR U33998 ( .A(n35430), .B(n35429), .Z(n35432) );
  XNOR U33999 ( .A(n35427), .B(n35426), .Z(n35429) );
  XNOR U34000 ( .A(n35424), .B(n35423), .Z(n35426) );
  XNOR U34001 ( .A(n35421), .B(n35420), .Z(n35423) );
  XNOR U34002 ( .A(n35418), .B(n35417), .Z(n35420) );
  XNOR U34003 ( .A(n35415), .B(n35414), .Z(n35417) );
  XNOR U34004 ( .A(n35412), .B(n35411), .Z(n35414) );
  XNOR U34005 ( .A(n35409), .B(n35408), .Z(n35411) );
  XNOR U34006 ( .A(n35406), .B(n35405), .Z(n35408) );
  XNOR U34007 ( .A(n35403), .B(n35402), .Z(n35405) );
  XNOR U34008 ( .A(n35400), .B(n35399), .Z(n35402) );
  XNOR U34009 ( .A(n35397), .B(n35396), .Z(n35399) );
  XNOR U34010 ( .A(n35394), .B(n35393), .Z(n35396) );
  XNOR U34011 ( .A(n35391), .B(n35390), .Z(n35393) );
  XNOR U34012 ( .A(n35388), .B(n35387), .Z(n35390) );
  XNOR U34013 ( .A(n35385), .B(n35384), .Z(n35387) );
  XNOR U34014 ( .A(n35382), .B(n35381), .Z(n35384) );
  XNOR U34015 ( .A(n35379), .B(n35378), .Z(n35381) );
  XNOR U34016 ( .A(n35376), .B(n35375), .Z(n35378) );
  XNOR U34017 ( .A(n35373), .B(n35372), .Z(n35375) );
  XNOR U34018 ( .A(n35370), .B(n35369), .Z(n35372) );
  XNOR U34019 ( .A(n35367), .B(n35366), .Z(n35369) );
  XNOR U34020 ( .A(n35364), .B(n35363), .Z(n35366) );
  XNOR U34021 ( .A(n35361), .B(n35360), .Z(n35363) );
  XNOR U34022 ( .A(n35358), .B(n35357), .Z(n35360) );
  XNOR U34023 ( .A(n35355), .B(n35354), .Z(n35357) );
  XNOR U34024 ( .A(n35352), .B(n35351), .Z(n35354) );
  XNOR U34025 ( .A(n35349), .B(n35348), .Z(n35351) );
  XNOR U34026 ( .A(n35346), .B(n35345), .Z(n35348) );
  XNOR U34027 ( .A(n35343), .B(n35342), .Z(n35345) );
  XNOR U34028 ( .A(n35340), .B(n35339), .Z(n35342) );
  XNOR U34029 ( .A(n35337), .B(n35336), .Z(n35339) );
  XNOR U34030 ( .A(n35334), .B(n35333), .Z(n35336) );
  XNOR U34031 ( .A(n35331), .B(n35330), .Z(n35333) );
  XNOR U34032 ( .A(n35328), .B(n35327), .Z(n35330) );
  XNOR U34033 ( .A(n35325), .B(n35324), .Z(n35327) );
  XNOR U34034 ( .A(n35322), .B(n35321), .Z(n35324) );
  XNOR U34035 ( .A(n35319), .B(n35318), .Z(n35321) );
  XNOR U34036 ( .A(n35316), .B(n35315), .Z(n35318) );
  XNOR U34037 ( .A(n35313), .B(n35312), .Z(n35315) );
  XNOR U34038 ( .A(n35310), .B(n35309), .Z(n35312) );
  XNOR U34039 ( .A(n35307), .B(n35306), .Z(n35309) );
  XNOR U34040 ( .A(n35304), .B(n35303), .Z(n35306) );
  XNOR U34041 ( .A(n35301), .B(n35300), .Z(n35303) );
  XNOR U34042 ( .A(n35298), .B(n35297), .Z(n35300) );
  XNOR U34043 ( .A(n35295), .B(n35294), .Z(n35297) );
  XNOR U34044 ( .A(n35292), .B(n35291), .Z(n35294) );
  XNOR U34045 ( .A(n35289), .B(n35288), .Z(n35291) );
  XNOR U34046 ( .A(n35286), .B(n35285), .Z(n35288) );
  XNOR U34047 ( .A(n35283), .B(n35282), .Z(n35285) );
  XNOR U34048 ( .A(n35280), .B(n35279), .Z(n35282) );
  XNOR U34049 ( .A(n35277), .B(n35276), .Z(n35279) );
  XNOR U34050 ( .A(n35274), .B(n35273), .Z(n35276) );
  XNOR U34051 ( .A(n35271), .B(n35270), .Z(n35273) );
  XNOR U34052 ( .A(n35268), .B(n35267), .Z(n35270) );
  XNOR U34053 ( .A(n35265), .B(n35264), .Z(n35267) );
  XNOR U34054 ( .A(n35262), .B(n35261), .Z(n35264) );
  XNOR U34055 ( .A(n35259), .B(n35258), .Z(n35261) );
  XNOR U34056 ( .A(n35256), .B(n35255), .Z(n35258) );
  XNOR U34057 ( .A(n35253), .B(n35252), .Z(n35255) );
  XNOR U34058 ( .A(n35250), .B(n35249), .Z(n35252) );
  XNOR U34059 ( .A(n35247), .B(n35246), .Z(n35249) );
  XNOR U34060 ( .A(n35244), .B(n35243), .Z(n35246) );
  XNOR U34061 ( .A(n35241), .B(n35240), .Z(n35243) );
  XNOR U34062 ( .A(n35238), .B(n35237), .Z(n35240) );
  XNOR U34063 ( .A(n35235), .B(n35234), .Z(n35237) );
  XNOR U34064 ( .A(n35232), .B(n35231), .Z(n35234) );
  XNOR U34065 ( .A(n35229), .B(n35228), .Z(n35231) );
  XNOR U34066 ( .A(n35226), .B(n35225), .Z(n35228) );
  XNOR U34067 ( .A(n35223), .B(n35222), .Z(n35225) );
  XNOR U34068 ( .A(n35220), .B(n35219), .Z(n35222) );
  XNOR U34069 ( .A(n35217), .B(n35216), .Z(n35219) );
  XNOR U34070 ( .A(n35214), .B(n35213), .Z(n35216) );
  XNOR U34071 ( .A(n35211), .B(n35210), .Z(n35213) );
  XNOR U34072 ( .A(n35208), .B(n35207), .Z(n35210) );
  XNOR U34073 ( .A(n35205), .B(n35204), .Z(n35207) );
  XNOR U34074 ( .A(n35202), .B(n35201), .Z(n35204) );
  XNOR U34075 ( .A(n35199), .B(n35198), .Z(n35201) );
  XNOR U34076 ( .A(n35196), .B(n35195), .Z(n35198) );
  XNOR U34077 ( .A(n35193), .B(n35192), .Z(n35195) );
  XNOR U34078 ( .A(n35190), .B(n35189), .Z(n35192) );
  XNOR U34079 ( .A(n35187), .B(n35186), .Z(n35189) );
  XNOR U34080 ( .A(n35184), .B(n35183), .Z(n35186) );
  XNOR U34081 ( .A(n35181), .B(n35180), .Z(n35183) );
  XNOR U34082 ( .A(n35178), .B(n35177), .Z(n35180) );
  XNOR U34083 ( .A(n35175), .B(n35174), .Z(n35177) );
  XNOR U34084 ( .A(n35172), .B(n35171), .Z(n35174) );
  XNOR U34085 ( .A(n35169), .B(n35168), .Z(n35171) );
  XNOR U34086 ( .A(n35166), .B(n35165), .Z(n35168) );
  XNOR U34087 ( .A(n35163), .B(n35162), .Z(n35165) );
  XNOR U34088 ( .A(n35160), .B(n35159), .Z(n35162) );
  XNOR U34089 ( .A(n35157), .B(n35156), .Z(n35159) );
  XNOR U34090 ( .A(n35154), .B(n35153), .Z(n35156) );
  XNOR U34091 ( .A(n35151), .B(n35150), .Z(n35153) );
  XNOR U34092 ( .A(n35148), .B(n35147), .Z(n35150) );
  XNOR U34093 ( .A(n35145), .B(n35144), .Z(n35147) );
  XNOR U34094 ( .A(n35142), .B(n35141), .Z(n35144) );
  XNOR U34095 ( .A(n35139), .B(n35138), .Z(n35141) );
  XNOR U34096 ( .A(n35136), .B(n35135), .Z(n35138) );
  XNOR U34097 ( .A(n35133), .B(n35132), .Z(n35135) );
  XNOR U34098 ( .A(n35130), .B(n35129), .Z(n35132) );
  XNOR U34099 ( .A(n35127), .B(n35126), .Z(n35129) );
  XNOR U34100 ( .A(n35124), .B(n35123), .Z(n35126) );
  XNOR U34101 ( .A(n35121), .B(n35120), .Z(n35123) );
  XNOR U34102 ( .A(n35118), .B(n35117), .Z(n35120) );
  XNOR U34103 ( .A(n35115), .B(n35114), .Z(n35117) );
  XNOR U34104 ( .A(n35112), .B(n35111), .Z(n35114) );
  XNOR U34105 ( .A(n35109), .B(n35108), .Z(n35111) );
  XNOR U34106 ( .A(n35106), .B(n35105), .Z(n35108) );
  XNOR U34107 ( .A(n35103), .B(n35102), .Z(n35105) );
  XNOR U34108 ( .A(n35100), .B(n35099), .Z(n35102) );
  XNOR U34109 ( .A(n35097), .B(n35096), .Z(n35099) );
  XNOR U34110 ( .A(n35094), .B(n35093), .Z(n35096) );
  XNOR U34111 ( .A(n35091), .B(n35090), .Z(n35093) );
  XNOR U34112 ( .A(n35088), .B(n35087), .Z(n35090) );
  XNOR U34113 ( .A(n35085), .B(n35084), .Z(n35087) );
  XNOR U34114 ( .A(n35082), .B(n35081), .Z(n35084) );
  XNOR U34115 ( .A(n35079), .B(n35078), .Z(n35081) );
  XNOR U34116 ( .A(n35076), .B(n35075), .Z(n35078) );
  XNOR U34117 ( .A(n35073), .B(n35072), .Z(n35075) );
  XNOR U34118 ( .A(n35070), .B(n35069), .Z(n35072) );
  XNOR U34119 ( .A(n35067), .B(n35066), .Z(n35069) );
  XNOR U34120 ( .A(n35064), .B(n35063), .Z(n35066) );
  XNOR U34121 ( .A(n35061), .B(n35060), .Z(n35063) );
  XNOR U34122 ( .A(n35058), .B(n35057), .Z(n35060) );
  XNOR U34123 ( .A(n35055), .B(n35054), .Z(n35057) );
  XNOR U34124 ( .A(n35052), .B(n35051), .Z(n35054) );
  XNOR U34125 ( .A(n35049), .B(n35048), .Z(n35051) );
  XNOR U34126 ( .A(n35046), .B(n35045), .Z(n35048) );
  XNOR U34127 ( .A(n35043), .B(n35042), .Z(n35045) );
  XNOR U34128 ( .A(n35040), .B(n35039), .Z(n35042) );
  XNOR U34129 ( .A(n35037), .B(n35036), .Z(n35039) );
  XNOR U34130 ( .A(n35034), .B(n35033), .Z(n35036) );
  XNOR U34131 ( .A(n35031), .B(n35030), .Z(n35033) );
  XNOR U34132 ( .A(n35028), .B(n35027), .Z(n35030) );
  XNOR U34133 ( .A(n35025), .B(n35024), .Z(n35027) );
  XNOR U34134 ( .A(n35022), .B(n35021), .Z(n35024) );
  XNOR U34135 ( .A(n35019), .B(n35018), .Z(n35021) );
  XNOR U34136 ( .A(n35016), .B(n35015), .Z(n35018) );
  XNOR U34137 ( .A(n35013), .B(n35012), .Z(n35015) );
  XNOR U34138 ( .A(n35010), .B(n35009), .Z(n35012) );
  XNOR U34139 ( .A(n35007), .B(n35006), .Z(n35009) );
  XNOR U34140 ( .A(n35004), .B(n35003), .Z(n35006) );
  XNOR U34141 ( .A(n35001), .B(n35000), .Z(n35003) );
  XNOR U34142 ( .A(n34998), .B(n34997), .Z(n35000) );
  XNOR U34143 ( .A(n34995), .B(n34994), .Z(n34997) );
  XNOR U34144 ( .A(n34992), .B(n34991), .Z(n34994) );
  XNOR U34145 ( .A(n34989), .B(n34988), .Z(n34991) );
  XNOR U34146 ( .A(n34986), .B(n34985), .Z(n34988) );
  XNOR U34147 ( .A(n34983), .B(n34982), .Z(n34985) );
  XNOR U34148 ( .A(n34980), .B(n34979), .Z(n34982) );
  XNOR U34149 ( .A(n34977), .B(n34976), .Z(n34979) );
  XNOR U34150 ( .A(n34974), .B(n34973), .Z(n34976) );
  XNOR U34151 ( .A(n34971), .B(n34970), .Z(n34973) );
  XNOR U34152 ( .A(n34968), .B(n34967), .Z(n34970) );
  XNOR U34153 ( .A(n34965), .B(n34964), .Z(n34967) );
  XNOR U34154 ( .A(n34962), .B(n34961), .Z(n34964) );
  XNOR U34155 ( .A(n34959), .B(n34958), .Z(n34961) );
  XNOR U34156 ( .A(n34956), .B(n34955), .Z(n34958) );
  XNOR U34157 ( .A(n34953), .B(n34952), .Z(n34955) );
  XNOR U34158 ( .A(n34950), .B(n34949), .Z(n34952) );
  XNOR U34159 ( .A(n34947), .B(n34946), .Z(n34949) );
  XNOR U34160 ( .A(n34944), .B(n34943), .Z(n34946) );
  XNOR U34161 ( .A(n34941), .B(n34940), .Z(n34943) );
  XNOR U34162 ( .A(n34938), .B(n34937), .Z(n34940) );
  XNOR U34163 ( .A(n34935), .B(n34934), .Z(n34937) );
  XNOR U34164 ( .A(n34932), .B(n34931), .Z(n34934) );
  XNOR U34165 ( .A(n34929), .B(n34928), .Z(n34931) );
  XNOR U34166 ( .A(n34926), .B(n34925), .Z(n34928) );
  XNOR U34167 ( .A(n34923), .B(n34922), .Z(n34925) );
  XNOR U34168 ( .A(n34920), .B(n34919), .Z(n34922) );
  XNOR U34169 ( .A(n34917), .B(n34916), .Z(n34919) );
  XNOR U34170 ( .A(n34914), .B(n34913), .Z(n34916) );
  XNOR U34171 ( .A(n34911), .B(n34910), .Z(n34913) );
  XNOR U34172 ( .A(n34908), .B(n34907), .Z(n34910) );
  XNOR U34173 ( .A(n34905), .B(n34904), .Z(n34907) );
  XNOR U34174 ( .A(n34902), .B(n34901), .Z(n34904) );
  XNOR U34175 ( .A(n34899), .B(n34898), .Z(n34901) );
  XNOR U34176 ( .A(n34896), .B(n34895), .Z(n34898) );
  XNOR U34177 ( .A(n34893), .B(n34892), .Z(n34895) );
  XNOR U34178 ( .A(n34890), .B(n34889), .Z(n34892) );
  XNOR U34179 ( .A(n34887), .B(n34886), .Z(n34889) );
  XNOR U34180 ( .A(n34884), .B(n34883), .Z(n34886) );
  XNOR U34181 ( .A(n34881), .B(n34880), .Z(n34883) );
  XNOR U34182 ( .A(n34878), .B(n34877), .Z(n34880) );
  XNOR U34183 ( .A(n34875), .B(n34874), .Z(n34877) );
  XNOR U34184 ( .A(n34872), .B(n34871), .Z(n34874) );
  XNOR U34185 ( .A(n34869), .B(n34868), .Z(n34871) );
  XNOR U34186 ( .A(n34866), .B(n34865), .Z(n34868) );
  XNOR U34187 ( .A(n34863), .B(n34862), .Z(n34865) );
  XNOR U34188 ( .A(n34860), .B(n34859), .Z(n34862) );
  XNOR U34189 ( .A(n34857), .B(n34856), .Z(n34859) );
  XNOR U34190 ( .A(n34854), .B(n34853), .Z(n34856) );
  XNOR U34191 ( .A(n34851), .B(n34850), .Z(n34853) );
  XNOR U34192 ( .A(n34848), .B(n34847), .Z(n34850) );
  XNOR U34193 ( .A(n34845), .B(n34844), .Z(n34847) );
  XNOR U34194 ( .A(n34842), .B(n34841), .Z(n34844) );
  XNOR U34195 ( .A(n34839), .B(n34838), .Z(n34841) );
  XNOR U34196 ( .A(n34836), .B(n34835), .Z(n34838) );
  XNOR U34197 ( .A(n34833), .B(n34832), .Z(n34835) );
  XNOR U34198 ( .A(n34830), .B(n34829), .Z(n34832) );
  XNOR U34199 ( .A(n34827), .B(n34826), .Z(n34829) );
  XNOR U34200 ( .A(n34824), .B(n34823), .Z(n34826) );
  XNOR U34201 ( .A(n34821), .B(n34820), .Z(n34823) );
  XNOR U34202 ( .A(n34818), .B(n34817), .Z(n34820) );
  XNOR U34203 ( .A(n34815), .B(n34814), .Z(n34817) );
  XNOR U34204 ( .A(n34812), .B(n34811), .Z(n34814) );
  XNOR U34205 ( .A(n34809), .B(n34808), .Z(n34811) );
  XNOR U34206 ( .A(n34806), .B(n34805), .Z(n34808) );
  XNOR U34207 ( .A(n34803), .B(n34802), .Z(n34805) );
  XNOR U34208 ( .A(n34800), .B(n34799), .Z(n34802) );
  XNOR U34209 ( .A(n34797), .B(n34796), .Z(n34799) );
  XNOR U34210 ( .A(n34794), .B(n34793), .Z(n34796) );
  XNOR U34211 ( .A(n34791), .B(n34790), .Z(n34793) );
  XNOR U34212 ( .A(n34788), .B(n34787), .Z(n34790) );
  XNOR U34213 ( .A(n34785), .B(n34784), .Z(n34787) );
  XNOR U34214 ( .A(n34782), .B(n34781), .Z(n34784) );
  XNOR U34215 ( .A(n34779), .B(n34778), .Z(n34781) );
  XNOR U34216 ( .A(n34776), .B(n34775), .Z(n34778) );
  XNOR U34217 ( .A(n34773), .B(n34772), .Z(n34775) );
  XNOR U34218 ( .A(n34770), .B(n34769), .Z(n34772) );
  XNOR U34219 ( .A(n34767), .B(n34766), .Z(n34769) );
  XNOR U34220 ( .A(n34764), .B(n34763), .Z(n34766) );
  XNOR U34221 ( .A(n34761), .B(n34760), .Z(n34763) );
  XNOR U34222 ( .A(n34758), .B(n34757), .Z(n34760) );
  XNOR U34223 ( .A(n34755), .B(n34754), .Z(n34757) );
  XNOR U34224 ( .A(n34752), .B(n34751), .Z(n34754) );
  XNOR U34225 ( .A(n34749), .B(n34748), .Z(n34751) );
  XNOR U34226 ( .A(n34746), .B(n34745), .Z(n34748) );
  XNOR U34227 ( .A(n34743), .B(n34742), .Z(n34745) );
  XNOR U34228 ( .A(n34740), .B(n34739), .Z(n34742) );
  XNOR U34229 ( .A(n34737), .B(n34736), .Z(n34739) );
  XNOR U34230 ( .A(n34734), .B(n34733), .Z(n34736) );
  XNOR U34231 ( .A(n34731), .B(n34730), .Z(n34733) );
  XNOR U34232 ( .A(n34728), .B(n34727), .Z(n34730) );
  XNOR U34233 ( .A(n34725), .B(n34724), .Z(n34727) );
  XNOR U34234 ( .A(n34722), .B(n34721), .Z(n34724) );
  XNOR U34235 ( .A(n34719), .B(n34718), .Z(n34721) );
  XNOR U34236 ( .A(n34716), .B(n34715), .Z(n34718) );
  XNOR U34237 ( .A(n34713), .B(n34712), .Z(n34715) );
  XNOR U34238 ( .A(n34710), .B(n34709), .Z(n34712) );
  XNOR U34239 ( .A(n34707), .B(n34706), .Z(n34709) );
  XNOR U34240 ( .A(n34704), .B(n34703), .Z(n34706) );
  XNOR U34241 ( .A(n34701), .B(n34700), .Z(n34703) );
  XNOR U34242 ( .A(n34698), .B(n34697), .Z(n34700) );
  XNOR U34243 ( .A(n34695), .B(n34694), .Z(n34697) );
  XNOR U34244 ( .A(n34692), .B(n34691), .Z(n34694) );
  XNOR U34245 ( .A(n34689), .B(n34688), .Z(n34691) );
  XNOR U34246 ( .A(n34686), .B(n34685), .Z(n34688) );
  XNOR U34247 ( .A(n34683), .B(n34682), .Z(n34685) );
  XNOR U34248 ( .A(n34680), .B(n34679), .Z(n34682) );
  XNOR U34249 ( .A(n34677), .B(n34676), .Z(n34679) );
  XNOR U34250 ( .A(n34674), .B(n34673), .Z(n34676) );
  XNOR U34251 ( .A(n34671), .B(n34670), .Z(n34673) );
  XNOR U34252 ( .A(n34668), .B(n34667), .Z(n34670) );
  XNOR U34253 ( .A(n34665), .B(n34664), .Z(n34667) );
  XNOR U34254 ( .A(n34662), .B(n34661), .Z(n34664) );
  XNOR U34255 ( .A(n34659), .B(n34658), .Z(n34661) );
  XNOR U34256 ( .A(n34656), .B(n34655), .Z(n34658) );
  XNOR U34257 ( .A(n34653), .B(n34652), .Z(n34655) );
  XNOR U34258 ( .A(n34650), .B(n34649), .Z(n34652) );
  XNOR U34259 ( .A(n34647), .B(n34646), .Z(n34649) );
  XNOR U34260 ( .A(n34644), .B(n34643), .Z(n34646) );
  XNOR U34261 ( .A(n34641), .B(n34640), .Z(n34643) );
  XNOR U34262 ( .A(n34638), .B(n34637), .Z(n34640) );
  XNOR U34263 ( .A(n34635), .B(n34634), .Z(n34637) );
  XNOR U34264 ( .A(n34632), .B(n34631), .Z(n34634) );
  XNOR U34265 ( .A(n34629), .B(n34628), .Z(n34631) );
  XNOR U34266 ( .A(n34626), .B(n34625), .Z(n34628) );
  XNOR U34267 ( .A(n34623), .B(n34622), .Z(n34625) );
  XNOR U34268 ( .A(n34620), .B(n34619), .Z(n34622) );
  XNOR U34269 ( .A(n34617), .B(n34616), .Z(n34619) );
  XNOR U34270 ( .A(n34614), .B(n34613), .Z(n34616) );
  XNOR U34271 ( .A(n34611), .B(n34610), .Z(n34613) );
  XNOR U34272 ( .A(n34608), .B(n34607), .Z(n34610) );
  XNOR U34273 ( .A(n34605), .B(n34604), .Z(n34607) );
  XNOR U34274 ( .A(n34602), .B(n34601), .Z(n34604) );
  XNOR U34275 ( .A(n34599), .B(n34598), .Z(n34601) );
  XNOR U34276 ( .A(n34596), .B(n34595), .Z(n34598) );
  XNOR U34277 ( .A(n34593), .B(n34592), .Z(n34595) );
  XNOR U34278 ( .A(n34590), .B(n34589), .Z(n34592) );
  XNOR U34279 ( .A(n34587), .B(n34586), .Z(n34589) );
  XNOR U34280 ( .A(n34584), .B(n34583), .Z(n34586) );
  XNOR U34281 ( .A(n34581), .B(n34580), .Z(n34583) );
  XNOR U34282 ( .A(n34578), .B(n34577), .Z(n34580) );
  XNOR U34283 ( .A(n34575), .B(n34574), .Z(n34577) );
  XNOR U34284 ( .A(n34572), .B(n34571), .Z(n34574) );
  XNOR U34285 ( .A(n34569), .B(n34568), .Z(n34571) );
  XNOR U34286 ( .A(n34566), .B(n34565), .Z(n34568) );
  XNOR U34287 ( .A(n34563), .B(n34562), .Z(n34565) );
  XNOR U34288 ( .A(n34560), .B(n34559), .Z(n34562) );
  XNOR U34289 ( .A(n34557), .B(n34556), .Z(n34559) );
  XNOR U34290 ( .A(n34554), .B(n34553), .Z(n34556) );
  XNOR U34291 ( .A(n34551), .B(n34550), .Z(n34553) );
  XNOR U34292 ( .A(n34548), .B(n34547), .Z(n34550) );
  XNOR U34293 ( .A(n34545), .B(n34544), .Z(n34547) );
  XNOR U34294 ( .A(n34542), .B(n34541), .Z(n34544) );
  XNOR U34295 ( .A(n34539), .B(n34538), .Z(n34541) );
  XNOR U34296 ( .A(n34536), .B(n34535), .Z(n34538) );
  XNOR U34297 ( .A(n34533), .B(n34532), .Z(n34535) );
  XNOR U34298 ( .A(n34530), .B(n34529), .Z(n34532) );
  XNOR U34299 ( .A(n34527), .B(n34526), .Z(n34529) );
  XNOR U34300 ( .A(n34524), .B(n34523), .Z(n34526) );
  XNOR U34301 ( .A(n34521), .B(n34520), .Z(n34523) );
  XNOR U34302 ( .A(n34518), .B(n34517), .Z(n34520) );
  XNOR U34303 ( .A(n34515), .B(n34514), .Z(n34517) );
  XNOR U34304 ( .A(n34512), .B(n34511), .Z(n34514) );
  XNOR U34305 ( .A(n34509), .B(n34508), .Z(n34511) );
  XNOR U34306 ( .A(n34506), .B(n34505), .Z(n34508) );
  XNOR U34307 ( .A(n34503), .B(n34502), .Z(n34505) );
  XNOR U34308 ( .A(n34500), .B(n34499), .Z(n34502) );
  XNOR U34309 ( .A(n34497), .B(n34496), .Z(n34499) );
  XNOR U34310 ( .A(n34494), .B(n34493), .Z(n34496) );
  XNOR U34311 ( .A(n34491), .B(n34490), .Z(n34493) );
  XNOR U34312 ( .A(n34488), .B(n34487), .Z(n34490) );
  XNOR U34313 ( .A(n34485), .B(n34484), .Z(n34487) );
  XNOR U34314 ( .A(n34482), .B(n34481), .Z(n34484) );
  XNOR U34315 ( .A(n34479), .B(n34478), .Z(n34481) );
  XNOR U34316 ( .A(n34476), .B(n34475), .Z(n34478) );
  XNOR U34317 ( .A(n34473), .B(n34472), .Z(n34475) );
  XNOR U34318 ( .A(n34470), .B(n34469), .Z(n34472) );
  XNOR U34319 ( .A(n34467), .B(n34466), .Z(n34469) );
  XNOR U34320 ( .A(n34464), .B(n34463), .Z(n34466) );
  XNOR U34321 ( .A(n34461), .B(n34460), .Z(n34463) );
  XNOR U34322 ( .A(n34458), .B(n34457), .Z(n34460) );
  XNOR U34323 ( .A(n34455), .B(n34454), .Z(n34457) );
  XNOR U34324 ( .A(n34452), .B(n34451), .Z(n34454) );
  XNOR U34325 ( .A(n34449), .B(n34448), .Z(n34451) );
  XNOR U34326 ( .A(n34446), .B(n34445), .Z(n34448) );
  XNOR U34327 ( .A(n34443), .B(n34442), .Z(n34445) );
  XNOR U34328 ( .A(n34440), .B(n34439), .Z(n34442) );
  XNOR U34329 ( .A(n34437), .B(n34436), .Z(n34439) );
  XNOR U34330 ( .A(n34434), .B(n34433), .Z(n34436) );
  XNOR U34331 ( .A(n34431), .B(n34430), .Z(n34433) );
  XNOR U34332 ( .A(n34428), .B(n34427), .Z(n34430) );
  XNOR U34333 ( .A(n34425), .B(n34424), .Z(n34427) );
  XNOR U34334 ( .A(n34422), .B(n34421), .Z(n34424) );
  XNOR U34335 ( .A(n34419), .B(n34418), .Z(n34421) );
  XNOR U34336 ( .A(n34416), .B(n34415), .Z(n34418) );
  XNOR U34337 ( .A(n34413), .B(n34412), .Z(n34415) );
  XNOR U34338 ( .A(n34410), .B(n34409), .Z(n34412) );
  XNOR U34339 ( .A(n34407), .B(n34406), .Z(n34409) );
  XNOR U34340 ( .A(n34404), .B(n34403), .Z(n34406) );
  XNOR U34341 ( .A(n34401), .B(n34400), .Z(n34403) );
  XNOR U34342 ( .A(n34398), .B(n34397), .Z(n34400) );
  XNOR U34343 ( .A(n34395), .B(n34394), .Z(n34397) );
  XNOR U34344 ( .A(n34392), .B(n34391), .Z(n34394) );
  XNOR U34345 ( .A(n34389), .B(n34388), .Z(n34391) );
  XNOR U34346 ( .A(n34386), .B(n34385), .Z(n34388) );
  XNOR U34347 ( .A(n34383), .B(n34382), .Z(n34385) );
  XNOR U34348 ( .A(n34380), .B(n34379), .Z(n34382) );
  XNOR U34349 ( .A(n34377), .B(n34376), .Z(n34379) );
  XNOR U34350 ( .A(n34374), .B(n34373), .Z(n34376) );
  XNOR U34351 ( .A(n34371), .B(n34370), .Z(n34373) );
  XNOR U34352 ( .A(n34368), .B(n34367), .Z(n34370) );
  XOR U34353 ( .A(n34365), .B(n34364), .Z(n34367) );
  XOR U34354 ( .A(n34362), .B(n34361), .Z(n34364) );
  XOR U34355 ( .A(n34358), .B(n34359), .Z(n34361) );
  AND U34356 ( .A(n36967), .B(n36968), .Z(n34359) );
  XOR U34357 ( .A(n34355), .B(n34356), .Z(n34358) );
  AND U34358 ( .A(n36969), .B(n36970), .Z(n34356) );
  XOR U34359 ( .A(n34352), .B(n34353), .Z(n34355) );
  AND U34360 ( .A(n36971), .B(n36972), .Z(n34353) );
  XNOR U34361 ( .A(n34107), .B(n34350), .Z(n34352) );
  AND U34362 ( .A(n36973), .B(n36974), .Z(n34350) );
  XOR U34363 ( .A(n34109), .B(n34108), .Z(n34107) );
  AND U34364 ( .A(n36975), .B(n36976), .Z(n34108) );
  XOR U34365 ( .A(n34111), .B(n34110), .Z(n34109) );
  AND U34366 ( .A(n36977), .B(n36978), .Z(n34110) );
  XOR U34367 ( .A(n34113), .B(n34112), .Z(n34111) );
  AND U34368 ( .A(n36979), .B(n36980), .Z(n34112) );
  XOR U34369 ( .A(n34115), .B(n34114), .Z(n34113) );
  AND U34370 ( .A(n36981), .B(n36982), .Z(n34114) );
  XOR U34371 ( .A(n34117), .B(n34116), .Z(n34115) );
  AND U34372 ( .A(n36983), .B(n36984), .Z(n34116) );
  XOR U34373 ( .A(n34119), .B(n34118), .Z(n34117) );
  AND U34374 ( .A(n36985), .B(n36986), .Z(n34118) );
  XOR U34375 ( .A(n34121), .B(n34120), .Z(n34119) );
  AND U34376 ( .A(n36987), .B(n36988), .Z(n34120) );
  XOR U34377 ( .A(n34123), .B(n34122), .Z(n34121) );
  AND U34378 ( .A(n36989), .B(n36990), .Z(n34122) );
  XOR U34379 ( .A(n34125), .B(n34124), .Z(n34123) );
  AND U34380 ( .A(n36991), .B(n36992), .Z(n34124) );
  XOR U34381 ( .A(n34127), .B(n34126), .Z(n34125) );
  AND U34382 ( .A(n36993), .B(n36994), .Z(n34126) );
  XOR U34383 ( .A(n34129), .B(n34128), .Z(n34127) );
  AND U34384 ( .A(n36995), .B(n36996), .Z(n34128) );
  XOR U34385 ( .A(n34131), .B(n34130), .Z(n34129) );
  AND U34386 ( .A(n36997), .B(n36998), .Z(n34130) );
  XOR U34387 ( .A(n34133), .B(n34132), .Z(n34131) );
  AND U34388 ( .A(n36999), .B(n37000), .Z(n34132) );
  XOR U34389 ( .A(n34135), .B(n34134), .Z(n34133) );
  AND U34390 ( .A(n37001), .B(n37002), .Z(n34134) );
  XOR U34391 ( .A(n34137), .B(n34136), .Z(n34135) );
  AND U34392 ( .A(n37003), .B(n37004), .Z(n34136) );
  XOR U34393 ( .A(n34139), .B(n34138), .Z(n34137) );
  AND U34394 ( .A(n37005), .B(n37006), .Z(n34138) );
  XOR U34395 ( .A(n34141), .B(n34140), .Z(n34139) );
  AND U34396 ( .A(n37007), .B(n37008), .Z(n34140) );
  XOR U34397 ( .A(n34143), .B(n34142), .Z(n34141) );
  AND U34398 ( .A(n37009), .B(n37010), .Z(n34142) );
  XOR U34399 ( .A(n34145), .B(n34144), .Z(n34143) );
  AND U34400 ( .A(n37011), .B(n37012), .Z(n34144) );
  XOR U34401 ( .A(n34147), .B(n34146), .Z(n34145) );
  AND U34402 ( .A(n37013), .B(n37014), .Z(n34146) );
  XOR U34403 ( .A(n34149), .B(n34148), .Z(n34147) );
  AND U34404 ( .A(n37015), .B(n37016), .Z(n34148) );
  XOR U34405 ( .A(n34151), .B(n34150), .Z(n34149) );
  AND U34406 ( .A(n37017), .B(n37018), .Z(n34150) );
  XOR U34407 ( .A(n34153), .B(n34152), .Z(n34151) );
  AND U34408 ( .A(n37019), .B(n37020), .Z(n34152) );
  XOR U34409 ( .A(n34155), .B(n34154), .Z(n34153) );
  AND U34410 ( .A(n37021), .B(n37022), .Z(n34154) );
  XOR U34411 ( .A(n34157), .B(n34156), .Z(n34155) );
  AND U34412 ( .A(n37023), .B(n37024), .Z(n34156) );
  XOR U34413 ( .A(n34159), .B(n34158), .Z(n34157) );
  AND U34414 ( .A(n37025), .B(n37026), .Z(n34158) );
  XOR U34415 ( .A(n34161), .B(n34160), .Z(n34159) );
  AND U34416 ( .A(n37027), .B(n37028), .Z(n34160) );
  XOR U34417 ( .A(n34163), .B(n34162), .Z(n34161) );
  AND U34418 ( .A(n37029), .B(n37030), .Z(n34162) );
  XOR U34419 ( .A(n34165), .B(n34164), .Z(n34163) );
  AND U34420 ( .A(n37031), .B(n37032), .Z(n34164) );
  XOR U34421 ( .A(n34167), .B(n34166), .Z(n34165) );
  AND U34422 ( .A(n37033), .B(n37034), .Z(n34166) );
  XOR U34423 ( .A(n34169), .B(n34168), .Z(n34167) );
  AND U34424 ( .A(n37035), .B(n37036), .Z(n34168) );
  XOR U34425 ( .A(n34171), .B(n34170), .Z(n34169) );
  AND U34426 ( .A(n37037), .B(n37038), .Z(n34170) );
  XOR U34427 ( .A(n34173), .B(n34172), .Z(n34171) );
  AND U34428 ( .A(n37039), .B(n37040), .Z(n34172) );
  XOR U34429 ( .A(n34175), .B(n34174), .Z(n34173) );
  AND U34430 ( .A(n37041), .B(n37042), .Z(n34174) );
  XOR U34431 ( .A(n34177), .B(n34176), .Z(n34175) );
  AND U34432 ( .A(n37043), .B(n37044), .Z(n34176) );
  XOR U34433 ( .A(n34179), .B(n34178), .Z(n34177) );
  AND U34434 ( .A(n37045), .B(n37046), .Z(n34178) );
  XOR U34435 ( .A(n34181), .B(n34180), .Z(n34179) );
  AND U34436 ( .A(n37047), .B(n37048), .Z(n34180) );
  XOR U34437 ( .A(n34183), .B(n34182), .Z(n34181) );
  AND U34438 ( .A(n37049), .B(n37050), .Z(n34182) );
  XOR U34439 ( .A(n34185), .B(n34184), .Z(n34183) );
  AND U34440 ( .A(n37051), .B(n37052), .Z(n34184) );
  XOR U34441 ( .A(n34187), .B(n34186), .Z(n34185) );
  AND U34442 ( .A(n37053), .B(n37054), .Z(n34186) );
  XOR U34443 ( .A(n34189), .B(n34188), .Z(n34187) );
  AND U34444 ( .A(n37055), .B(n37056), .Z(n34188) );
  XOR U34445 ( .A(n34191), .B(n34190), .Z(n34189) );
  AND U34446 ( .A(n37057), .B(n37058), .Z(n34190) );
  XOR U34447 ( .A(n34193), .B(n34192), .Z(n34191) );
  AND U34448 ( .A(n37059), .B(n37060), .Z(n34192) );
  XOR U34449 ( .A(n34195), .B(n34194), .Z(n34193) );
  AND U34450 ( .A(n37061), .B(n37062), .Z(n34194) );
  XOR U34451 ( .A(n34197), .B(n34196), .Z(n34195) );
  AND U34452 ( .A(n37063), .B(n37064), .Z(n34196) );
  XOR U34453 ( .A(n34199), .B(n34198), .Z(n34197) );
  AND U34454 ( .A(n37065), .B(n37066), .Z(n34198) );
  XOR U34455 ( .A(n34201), .B(n34200), .Z(n34199) );
  AND U34456 ( .A(n37067), .B(n37068), .Z(n34200) );
  XOR U34457 ( .A(n34203), .B(n34202), .Z(n34201) );
  AND U34458 ( .A(n37069), .B(n37070), .Z(n34202) );
  XOR U34459 ( .A(n34205), .B(n34204), .Z(n34203) );
  AND U34460 ( .A(n37071), .B(n37072), .Z(n34204) );
  XOR U34461 ( .A(n34207), .B(n34206), .Z(n34205) );
  AND U34462 ( .A(n37073), .B(n37074), .Z(n34206) );
  XOR U34463 ( .A(n34209), .B(n34208), .Z(n34207) );
  AND U34464 ( .A(n37075), .B(n37076), .Z(n34208) );
  XOR U34465 ( .A(n34211), .B(n34210), .Z(n34209) );
  AND U34466 ( .A(n37077), .B(n37078), .Z(n34210) );
  XOR U34467 ( .A(n34213), .B(n34212), .Z(n34211) );
  AND U34468 ( .A(n37079), .B(n37080), .Z(n34212) );
  XOR U34469 ( .A(n34215), .B(n34214), .Z(n34213) );
  AND U34470 ( .A(n37081), .B(n37082), .Z(n34214) );
  XOR U34471 ( .A(n34217), .B(n34216), .Z(n34215) );
  AND U34472 ( .A(n37083), .B(n37084), .Z(n34216) );
  XOR U34473 ( .A(n34219), .B(n34218), .Z(n34217) );
  AND U34474 ( .A(n37085), .B(n37086), .Z(n34218) );
  XOR U34475 ( .A(n34221), .B(n34220), .Z(n34219) );
  AND U34476 ( .A(n37087), .B(n37088), .Z(n34220) );
  XOR U34477 ( .A(n34223), .B(n34222), .Z(n34221) );
  AND U34478 ( .A(n37089), .B(n37090), .Z(n34222) );
  XOR U34479 ( .A(n34225), .B(n34224), .Z(n34223) );
  AND U34480 ( .A(n37091), .B(n37092), .Z(n34224) );
  XOR U34481 ( .A(n34227), .B(n34226), .Z(n34225) );
  AND U34482 ( .A(n37093), .B(n37094), .Z(n34226) );
  XOR U34483 ( .A(n34229), .B(n34228), .Z(n34227) );
  AND U34484 ( .A(n37095), .B(n37096), .Z(n34228) );
  XOR U34485 ( .A(n34231), .B(n34230), .Z(n34229) );
  AND U34486 ( .A(n37097), .B(n37098), .Z(n34230) );
  XOR U34487 ( .A(n34233), .B(n34232), .Z(n34231) );
  AND U34488 ( .A(n37099), .B(n37100), .Z(n34232) );
  XOR U34489 ( .A(n34235), .B(n34234), .Z(n34233) );
  AND U34490 ( .A(n37101), .B(n37102), .Z(n34234) );
  XOR U34491 ( .A(n34237), .B(n34236), .Z(n34235) );
  AND U34492 ( .A(n37103), .B(n37104), .Z(n34236) );
  XOR U34493 ( .A(n34239), .B(n34238), .Z(n34237) );
  AND U34494 ( .A(n37105), .B(n37106), .Z(n34238) );
  XOR U34495 ( .A(n34241), .B(n34240), .Z(n34239) );
  AND U34496 ( .A(n37107), .B(n37108), .Z(n34240) );
  XOR U34497 ( .A(n34243), .B(n34242), .Z(n34241) );
  AND U34498 ( .A(n37109), .B(n37110), .Z(n34242) );
  XOR U34499 ( .A(n34252), .B(n34244), .Z(n34243) );
  AND U34500 ( .A(n37111), .B(n37112), .Z(n34244) );
  XOR U34501 ( .A(n34247), .B(n34253), .Z(n34252) );
  AND U34502 ( .A(n37113), .B(n37114), .Z(n34253) );
  XOR U34503 ( .A(n34249), .B(n34248), .Z(n34247) );
  AND U34504 ( .A(n37115), .B(n37116), .Z(n34248) );
  XOR U34505 ( .A(n34273), .B(n34250), .Z(n34249) );
  AND U34506 ( .A(n37117), .B(n37118), .Z(n34250) );
  XOR U34507 ( .A(n34268), .B(n34274), .Z(n34273) );
  AND U34508 ( .A(n37119), .B(n37120), .Z(n34274) );
  XOR U34509 ( .A(n34270), .B(n34269), .Z(n34268) );
  AND U34510 ( .A(n37121), .B(n37122), .Z(n34269) );
  XOR U34511 ( .A(n34258), .B(n34271), .Z(n34270) );
  AND U34512 ( .A(n37123), .B(n37124), .Z(n34271) );
  XOR U34513 ( .A(n34260), .B(n34259), .Z(n34258) );
  AND U34514 ( .A(n37125), .B(n37126), .Z(n34259) );
  XOR U34515 ( .A(n34262), .B(n34261), .Z(n34260) );
  AND U34516 ( .A(n37127), .B(n37128), .Z(n34261) );
  XOR U34517 ( .A(n34264), .B(n34263), .Z(n34262) );
  AND U34518 ( .A(n37129), .B(n37130), .Z(n34263) );
  XOR U34519 ( .A(n34294), .B(n34265), .Z(n34264) );
  AND U34520 ( .A(n37131), .B(n37132), .Z(n34265) );
  XOR U34521 ( .A(n34290), .B(n34295), .Z(n34294) );
  AND U34522 ( .A(n37133), .B(n37134), .Z(n34295) );
  XOR U34523 ( .A(n34292), .B(n34291), .Z(n34290) );
  AND U34524 ( .A(n37135), .B(n37136), .Z(n34291) );
  XOR U34525 ( .A(n34279), .B(n34293), .Z(n34292) );
  AND U34526 ( .A(n37137), .B(n37138), .Z(n34293) );
  XOR U34527 ( .A(n34281), .B(n34280), .Z(n34279) );
  AND U34528 ( .A(n37139), .B(n37140), .Z(n34280) );
  XOR U34529 ( .A(n34284), .B(n34282), .Z(n34281) );
  AND U34530 ( .A(n37141), .B(n37142), .Z(n34282) );
  XOR U34531 ( .A(n34286), .B(n34285), .Z(n34284) );
  AND U34532 ( .A(n37143), .B(n37144), .Z(n34285) );
  XOR U34533 ( .A(n34304), .B(n34287), .Z(n34286) );
  AND U34534 ( .A(n37145), .B(n37146), .Z(n34287) );
  XNOR U34535 ( .A(n34311), .B(n34305), .Z(n34304) );
  AND U34536 ( .A(n37147), .B(n37148), .Z(n34305) );
  XOR U34537 ( .A(n34310), .B(n34302), .Z(n34311) );
  AND U34538 ( .A(n37149), .B(n37150), .Z(n34302) );
  XOR U34539 ( .A(n34349), .B(n34301), .Z(n34310) );
  AND U34540 ( .A(n37151), .B(n37152), .Z(n34301) );
  XNOR U34541 ( .A(n34322), .B(n34300), .Z(n34349) );
  AND U34542 ( .A(n37153), .B(n37154), .Z(n34300) );
  XNOR U34543 ( .A(n34329), .B(n34323), .Z(n34322) );
  AND U34544 ( .A(n37155), .B(n37156), .Z(n34323) );
  XOR U34545 ( .A(n34328), .B(n34320), .Z(n34329) );
  AND U34546 ( .A(n37157), .B(n37158), .Z(n34320) );
  XOR U34547 ( .A(n34348), .B(n34319), .Z(n34328) );
  AND U34548 ( .A(n37159), .B(n37160), .Z(n34319) );
  XNOR U34549 ( .A(n37161), .B(n37162), .Z(n34348) );
  XOR U34550 ( .A(n37163), .B(n37164), .Z(n37162) );
  XOR U34551 ( .A(n37165), .B(n37166), .Z(n37164) );
  XNOR U34552 ( .A(n34346), .B(n34339), .Z(n37166) );
  XNOR U34553 ( .A(n37167), .B(n37168), .Z(n34339) );
  AND U34554 ( .A(n37169), .B(n37170), .Z(n37168) );
  NOR U34555 ( .A(n37171), .B(n37172), .Z(n37170) );
  NOR U34556 ( .A(n37173), .B(n37174), .Z(n37169) );
  AND U34557 ( .A(n37175), .B(n37176), .Z(n37174) );
  AND U34558 ( .A(n37177), .B(n37178), .Z(n37167) );
  NOR U34559 ( .A(n37179), .B(n37180), .Z(n37178) );
  AND U34560 ( .A(n37172), .B(n37181), .Z(n37180) );
  AND U34561 ( .A(n37173), .B(n37182), .Z(n37179) );
  NOR U34562 ( .A(n37183), .B(n37184), .Z(n37177) );
  AND U34563 ( .A(n37185), .B(n37186), .Z(n37184) );
  NOR U34564 ( .A(n37187), .B(n37188), .Z(n37186) );
  IV U34565 ( .A(n37189), .Z(n37187) );
  NOR U34566 ( .A(n37190), .B(n37191), .Z(n37189) );
  NOR U34567 ( .A(n37192), .B(n37193), .Z(n37185) );
  AND U34568 ( .A(n37171), .B(n37194), .Z(n37183) );
  AND U34569 ( .A(n37195), .B(n37196), .Z(n34346) );
  XOR U34570 ( .A(n34344), .B(n34345), .Z(n37165) );
  AND U34571 ( .A(n37197), .B(n37198), .Z(n34345) );
  AND U34572 ( .A(n37199), .B(n37200), .Z(n34344) );
  XOR U34573 ( .A(n37201), .B(n37202), .Z(n37163) );
  XOR U34574 ( .A(n34340), .B(n34341), .Z(n37202) );
  AND U34575 ( .A(n37203), .B(n37204), .Z(n34341) );
  AND U34576 ( .A(n37205), .B(n37206), .Z(n34340) );
  XNOR U34577 ( .A(n34338), .B(n34337), .Z(n37201) );
  IV U34578 ( .A(n37207), .Z(n34337) );
  AND U34579 ( .A(n37208), .B(n37209), .Z(n37207) );
  AND U34580 ( .A(n37210), .B(n37211), .Z(n34338) );
  XNOR U34581 ( .A(n34347), .B(n34318), .Z(n37161) );
  AND U34582 ( .A(n37212), .B(n37213), .Z(n34318) );
  AND U34583 ( .A(n37214), .B(n37215), .Z(n34347) );
  XOR U34584 ( .A(n37216), .B(n37217), .Z(n34362) );
  AND U34585 ( .A(n37216), .B(n37218), .Z(n37217) );
  XNOR U34586 ( .A(n37219), .B(n37220), .Z(n34365) );
  AND U34587 ( .A(n37219), .B(n37221), .Z(n37220) );
  XNOR U34588 ( .A(n37222), .B(n37223), .Z(n34368) );
  AND U34589 ( .A(n37222), .B(n37224), .Z(n37223) );
  XNOR U34590 ( .A(n37225), .B(n37226), .Z(n34371) );
  AND U34591 ( .A(n37225), .B(n37227), .Z(n37226) );
  XNOR U34592 ( .A(n37228), .B(n37229), .Z(n34374) );
  AND U34593 ( .A(n37230), .B(n37228), .Z(n37229) );
  XOR U34594 ( .A(n37231), .B(n37232), .Z(n34377) );
  NOR U34595 ( .A(n37233), .B(n37231), .Z(n37232) );
  XOR U34596 ( .A(n37234), .B(n37235), .Z(n34380) );
  NOR U34597 ( .A(n37236), .B(n37234), .Z(n37235) );
  XOR U34598 ( .A(n37237), .B(n37238), .Z(n34383) );
  NOR U34599 ( .A(n37239), .B(n37237), .Z(n37238) );
  XOR U34600 ( .A(n37240), .B(n37241), .Z(n34386) );
  NOR U34601 ( .A(n37242), .B(n37240), .Z(n37241) );
  XOR U34602 ( .A(n37243), .B(n37244), .Z(n34389) );
  NOR U34603 ( .A(n37245), .B(n37243), .Z(n37244) );
  XOR U34604 ( .A(n37246), .B(n37247), .Z(n34392) );
  NOR U34605 ( .A(n37248), .B(n37246), .Z(n37247) );
  XOR U34606 ( .A(n37249), .B(n37250), .Z(n34395) );
  NOR U34607 ( .A(n37251), .B(n37249), .Z(n37250) );
  XOR U34608 ( .A(n37252), .B(n37253), .Z(n34398) );
  NOR U34609 ( .A(n37254), .B(n37252), .Z(n37253) );
  XOR U34610 ( .A(n37255), .B(n37256), .Z(n34401) );
  NOR U34611 ( .A(n37257), .B(n37255), .Z(n37256) );
  XOR U34612 ( .A(n37258), .B(n37259), .Z(n34404) );
  NOR U34613 ( .A(n37260), .B(n37258), .Z(n37259) );
  XOR U34614 ( .A(n37261), .B(n37262), .Z(n34407) );
  NOR U34615 ( .A(n37263), .B(n37261), .Z(n37262) );
  XOR U34616 ( .A(n37264), .B(n37265), .Z(n34410) );
  NOR U34617 ( .A(n37266), .B(n37264), .Z(n37265) );
  XOR U34618 ( .A(n37267), .B(n37268), .Z(n34413) );
  NOR U34619 ( .A(n37269), .B(n37267), .Z(n37268) );
  XOR U34620 ( .A(n37270), .B(n37271), .Z(n34416) );
  NOR U34621 ( .A(n37272), .B(n37270), .Z(n37271) );
  XOR U34622 ( .A(n37273), .B(n37274), .Z(n34419) );
  NOR U34623 ( .A(n37275), .B(n37273), .Z(n37274) );
  XOR U34624 ( .A(n37276), .B(n37277), .Z(n34422) );
  NOR U34625 ( .A(n37278), .B(n37276), .Z(n37277) );
  XOR U34626 ( .A(n37279), .B(n37280), .Z(n34425) );
  NOR U34627 ( .A(n37281), .B(n37279), .Z(n37280) );
  XOR U34628 ( .A(n37282), .B(n37283), .Z(n34428) );
  NOR U34629 ( .A(n37284), .B(n37282), .Z(n37283) );
  XOR U34630 ( .A(n37285), .B(n37286), .Z(n34431) );
  NOR U34631 ( .A(n37287), .B(n37285), .Z(n37286) );
  XOR U34632 ( .A(n37288), .B(n37289), .Z(n34434) );
  NOR U34633 ( .A(n37290), .B(n37288), .Z(n37289) );
  XOR U34634 ( .A(n37291), .B(n37292), .Z(n34437) );
  NOR U34635 ( .A(n37293), .B(n37291), .Z(n37292) );
  XOR U34636 ( .A(n37294), .B(n37295), .Z(n34440) );
  NOR U34637 ( .A(n37296), .B(n37294), .Z(n37295) );
  XOR U34638 ( .A(n37297), .B(n37298), .Z(n34443) );
  NOR U34639 ( .A(n37299), .B(n37297), .Z(n37298) );
  XOR U34640 ( .A(n37300), .B(n37301), .Z(n34446) );
  NOR U34641 ( .A(n37302), .B(n37300), .Z(n37301) );
  XOR U34642 ( .A(n37303), .B(n37304), .Z(n34449) );
  NOR U34643 ( .A(n37305), .B(n37303), .Z(n37304) );
  XOR U34644 ( .A(n37306), .B(n37307), .Z(n34452) );
  NOR U34645 ( .A(n37308), .B(n37306), .Z(n37307) );
  XOR U34646 ( .A(n37309), .B(n37310), .Z(n34455) );
  NOR U34647 ( .A(n37311), .B(n37309), .Z(n37310) );
  XOR U34648 ( .A(n37312), .B(n37313), .Z(n34458) );
  NOR U34649 ( .A(n37314), .B(n37312), .Z(n37313) );
  XOR U34650 ( .A(n37315), .B(n37316), .Z(n34461) );
  NOR U34651 ( .A(n37317), .B(n37315), .Z(n37316) );
  XOR U34652 ( .A(n37318), .B(n37319), .Z(n34464) );
  NOR U34653 ( .A(n37320), .B(n37318), .Z(n37319) );
  XOR U34654 ( .A(n37321), .B(n37322), .Z(n34467) );
  NOR U34655 ( .A(n37323), .B(n37321), .Z(n37322) );
  XOR U34656 ( .A(n37324), .B(n37325), .Z(n34470) );
  NOR U34657 ( .A(n37326), .B(n37324), .Z(n37325) );
  XOR U34658 ( .A(n37327), .B(n37328), .Z(n34473) );
  NOR U34659 ( .A(n37329), .B(n37327), .Z(n37328) );
  XOR U34660 ( .A(n37330), .B(n37331), .Z(n34476) );
  NOR U34661 ( .A(n37332), .B(n37330), .Z(n37331) );
  XOR U34662 ( .A(n37333), .B(n37334), .Z(n34479) );
  NOR U34663 ( .A(n37335), .B(n37333), .Z(n37334) );
  XOR U34664 ( .A(n37336), .B(n37337), .Z(n34482) );
  NOR U34665 ( .A(n37338), .B(n37336), .Z(n37337) );
  XOR U34666 ( .A(n37339), .B(n37340), .Z(n34485) );
  NOR U34667 ( .A(n37341), .B(n37339), .Z(n37340) );
  XOR U34668 ( .A(n37342), .B(n37343), .Z(n34488) );
  NOR U34669 ( .A(n37344), .B(n37342), .Z(n37343) );
  XOR U34670 ( .A(n37345), .B(n37346), .Z(n34491) );
  NOR U34671 ( .A(n37347), .B(n37345), .Z(n37346) );
  XOR U34672 ( .A(n37348), .B(n37349), .Z(n34494) );
  NOR U34673 ( .A(n37350), .B(n37348), .Z(n37349) );
  XOR U34674 ( .A(n37351), .B(n37352), .Z(n34497) );
  NOR U34675 ( .A(n37353), .B(n37351), .Z(n37352) );
  XOR U34676 ( .A(n37354), .B(n37355), .Z(n34500) );
  NOR U34677 ( .A(n37356), .B(n37354), .Z(n37355) );
  XOR U34678 ( .A(n37357), .B(n37358), .Z(n34503) );
  NOR U34679 ( .A(n37359), .B(n37357), .Z(n37358) );
  XOR U34680 ( .A(n37360), .B(n37361), .Z(n34506) );
  NOR U34681 ( .A(n37362), .B(n37360), .Z(n37361) );
  XOR U34682 ( .A(n37363), .B(n37364), .Z(n34509) );
  NOR U34683 ( .A(n37365), .B(n37363), .Z(n37364) );
  XOR U34684 ( .A(n37366), .B(n37367), .Z(n34512) );
  NOR U34685 ( .A(n37368), .B(n37366), .Z(n37367) );
  XOR U34686 ( .A(n37369), .B(n37370), .Z(n34515) );
  NOR U34687 ( .A(n37371), .B(n37369), .Z(n37370) );
  XOR U34688 ( .A(n37372), .B(n37373), .Z(n34518) );
  NOR U34689 ( .A(n37374), .B(n37372), .Z(n37373) );
  XOR U34690 ( .A(n37375), .B(n37376), .Z(n34521) );
  NOR U34691 ( .A(n37377), .B(n37375), .Z(n37376) );
  XOR U34692 ( .A(n37378), .B(n37379), .Z(n34524) );
  NOR U34693 ( .A(n37380), .B(n37378), .Z(n37379) );
  XOR U34694 ( .A(n37381), .B(n37382), .Z(n34527) );
  NOR U34695 ( .A(n37383), .B(n37381), .Z(n37382) );
  XOR U34696 ( .A(n37384), .B(n37385), .Z(n34530) );
  NOR U34697 ( .A(n37386), .B(n37384), .Z(n37385) );
  XOR U34698 ( .A(n37387), .B(n37388), .Z(n34533) );
  NOR U34699 ( .A(n37389), .B(n37387), .Z(n37388) );
  XOR U34700 ( .A(n37390), .B(n37391), .Z(n34536) );
  NOR U34701 ( .A(n37392), .B(n37390), .Z(n37391) );
  XOR U34702 ( .A(n37393), .B(n37394), .Z(n34539) );
  NOR U34703 ( .A(n37395), .B(n37393), .Z(n37394) );
  XOR U34704 ( .A(n37396), .B(n37397), .Z(n34542) );
  NOR U34705 ( .A(n37398), .B(n37396), .Z(n37397) );
  XOR U34706 ( .A(n37399), .B(n37400), .Z(n34545) );
  NOR U34707 ( .A(n37401), .B(n37399), .Z(n37400) );
  XOR U34708 ( .A(n37402), .B(n37403), .Z(n34548) );
  NOR U34709 ( .A(n37404), .B(n37402), .Z(n37403) );
  XOR U34710 ( .A(n37405), .B(n37406), .Z(n34551) );
  NOR U34711 ( .A(n37407), .B(n37405), .Z(n37406) );
  XOR U34712 ( .A(n37408), .B(n37409), .Z(n34554) );
  NOR U34713 ( .A(n37410), .B(n37408), .Z(n37409) );
  XOR U34714 ( .A(n37411), .B(n37412), .Z(n34557) );
  NOR U34715 ( .A(n37413), .B(n37411), .Z(n37412) );
  XOR U34716 ( .A(n37414), .B(n37415), .Z(n34560) );
  NOR U34717 ( .A(n37416), .B(n37414), .Z(n37415) );
  XOR U34718 ( .A(n37417), .B(n37418), .Z(n34563) );
  NOR U34719 ( .A(n37419), .B(n37417), .Z(n37418) );
  XOR U34720 ( .A(n37420), .B(n37421), .Z(n34566) );
  NOR U34721 ( .A(n37422), .B(n37420), .Z(n37421) );
  XOR U34722 ( .A(n37423), .B(n37424), .Z(n34569) );
  NOR U34723 ( .A(n37425), .B(n37423), .Z(n37424) );
  XOR U34724 ( .A(n37426), .B(n37427), .Z(n34572) );
  NOR U34725 ( .A(n37428), .B(n37426), .Z(n37427) );
  XOR U34726 ( .A(n37429), .B(n37430), .Z(n34575) );
  NOR U34727 ( .A(n37431), .B(n37429), .Z(n37430) );
  XOR U34728 ( .A(n37432), .B(n37433), .Z(n34578) );
  NOR U34729 ( .A(n37434), .B(n37432), .Z(n37433) );
  XOR U34730 ( .A(n37435), .B(n37436), .Z(n34581) );
  NOR U34731 ( .A(n37437), .B(n37435), .Z(n37436) );
  XOR U34732 ( .A(n37438), .B(n37439), .Z(n34584) );
  NOR U34733 ( .A(n37440), .B(n37438), .Z(n37439) );
  XOR U34734 ( .A(n37441), .B(n37442), .Z(n34587) );
  NOR U34735 ( .A(n37443), .B(n37441), .Z(n37442) );
  XOR U34736 ( .A(n37444), .B(n37445), .Z(n34590) );
  NOR U34737 ( .A(n37446), .B(n37444), .Z(n37445) );
  XOR U34738 ( .A(n37447), .B(n37448), .Z(n34593) );
  NOR U34739 ( .A(n37449), .B(n37447), .Z(n37448) );
  XOR U34740 ( .A(n37450), .B(n37451), .Z(n34596) );
  NOR U34741 ( .A(n37452), .B(n37450), .Z(n37451) );
  XOR U34742 ( .A(n37453), .B(n37454), .Z(n34599) );
  NOR U34743 ( .A(n37455), .B(n37453), .Z(n37454) );
  XOR U34744 ( .A(n37456), .B(n37457), .Z(n34602) );
  NOR U34745 ( .A(n37458), .B(n37456), .Z(n37457) );
  XOR U34746 ( .A(n37459), .B(n37460), .Z(n34605) );
  NOR U34747 ( .A(n37461), .B(n37459), .Z(n37460) );
  XOR U34748 ( .A(n37462), .B(n37463), .Z(n34608) );
  NOR U34749 ( .A(n37464), .B(n37462), .Z(n37463) );
  XOR U34750 ( .A(n37465), .B(n37466), .Z(n34611) );
  NOR U34751 ( .A(n37467), .B(n37465), .Z(n37466) );
  XOR U34752 ( .A(n37468), .B(n37469), .Z(n34614) );
  NOR U34753 ( .A(n37470), .B(n37468), .Z(n37469) );
  XOR U34754 ( .A(n37471), .B(n37472), .Z(n34617) );
  NOR U34755 ( .A(n37473), .B(n37471), .Z(n37472) );
  XOR U34756 ( .A(n37474), .B(n37475), .Z(n34620) );
  NOR U34757 ( .A(n37476), .B(n37474), .Z(n37475) );
  XOR U34758 ( .A(n37477), .B(n37478), .Z(n34623) );
  NOR U34759 ( .A(n37479), .B(n37477), .Z(n37478) );
  XOR U34760 ( .A(n37480), .B(n37481), .Z(n34626) );
  NOR U34761 ( .A(n37482), .B(n37480), .Z(n37481) );
  XOR U34762 ( .A(n37483), .B(n37484), .Z(n34629) );
  NOR U34763 ( .A(n37485), .B(n37483), .Z(n37484) );
  XOR U34764 ( .A(n37486), .B(n37487), .Z(n34632) );
  NOR U34765 ( .A(n37488), .B(n37486), .Z(n37487) );
  XOR U34766 ( .A(n37489), .B(n37490), .Z(n34635) );
  NOR U34767 ( .A(n37491), .B(n37489), .Z(n37490) );
  XOR U34768 ( .A(n37492), .B(n37493), .Z(n34638) );
  NOR U34769 ( .A(n37494), .B(n37492), .Z(n37493) );
  XOR U34770 ( .A(n37495), .B(n37496), .Z(n34641) );
  NOR U34771 ( .A(n37497), .B(n37495), .Z(n37496) );
  XOR U34772 ( .A(n37498), .B(n37499), .Z(n34644) );
  NOR U34773 ( .A(n37500), .B(n37498), .Z(n37499) );
  XOR U34774 ( .A(n37501), .B(n37502), .Z(n34647) );
  NOR U34775 ( .A(n37503), .B(n37501), .Z(n37502) );
  XOR U34776 ( .A(n37504), .B(n37505), .Z(n34650) );
  NOR U34777 ( .A(n37506), .B(n37504), .Z(n37505) );
  XOR U34778 ( .A(n37507), .B(n37508), .Z(n34653) );
  NOR U34779 ( .A(n37509), .B(n37507), .Z(n37508) );
  XOR U34780 ( .A(n37510), .B(n37511), .Z(n34656) );
  NOR U34781 ( .A(n37512), .B(n37510), .Z(n37511) );
  XOR U34782 ( .A(n37513), .B(n37514), .Z(n34659) );
  NOR U34783 ( .A(n37515), .B(n37513), .Z(n37514) );
  XOR U34784 ( .A(n37516), .B(n37517), .Z(n34662) );
  NOR U34785 ( .A(n37518), .B(n37516), .Z(n37517) );
  XOR U34786 ( .A(n37519), .B(n37520), .Z(n34665) );
  NOR U34787 ( .A(n37521), .B(n37519), .Z(n37520) );
  XOR U34788 ( .A(n37522), .B(n37523), .Z(n34668) );
  NOR U34789 ( .A(n37524), .B(n37522), .Z(n37523) );
  XOR U34790 ( .A(n37525), .B(n37526), .Z(n34671) );
  NOR U34791 ( .A(n37527), .B(n37525), .Z(n37526) );
  XOR U34792 ( .A(n37528), .B(n37529), .Z(n34674) );
  NOR U34793 ( .A(n37530), .B(n37528), .Z(n37529) );
  XOR U34794 ( .A(n37531), .B(n37532), .Z(n34677) );
  NOR U34795 ( .A(n37533), .B(n37531), .Z(n37532) );
  XOR U34796 ( .A(n37534), .B(n37535), .Z(n34680) );
  NOR U34797 ( .A(n37536), .B(n37534), .Z(n37535) );
  XOR U34798 ( .A(n37537), .B(n37538), .Z(n34683) );
  NOR U34799 ( .A(n37539), .B(n37537), .Z(n37538) );
  XOR U34800 ( .A(n37540), .B(n37541), .Z(n34686) );
  NOR U34801 ( .A(n37542), .B(n37540), .Z(n37541) );
  XOR U34802 ( .A(n37543), .B(n37544), .Z(n34689) );
  NOR U34803 ( .A(n37545), .B(n37543), .Z(n37544) );
  XOR U34804 ( .A(n37546), .B(n37547), .Z(n34692) );
  NOR U34805 ( .A(n37548), .B(n37546), .Z(n37547) );
  XOR U34806 ( .A(n37549), .B(n37550), .Z(n34695) );
  NOR U34807 ( .A(n37551), .B(n37549), .Z(n37550) );
  XOR U34808 ( .A(n37552), .B(n37553), .Z(n34698) );
  NOR U34809 ( .A(n37554), .B(n37552), .Z(n37553) );
  XOR U34810 ( .A(n37555), .B(n37556), .Z(n34701) );
  NOR U34811 ( .A(n37557), .B(n37555), .Z(n37556) );
  XOR U34812 ( .A(n37558), .B(n37559), .Z(n34704) );
  NOR U34813 ( .A(n37560), .B(n37558), .Z(n37559) );
  XOR U34814 ( .A(n37561), .B(n37562), .Z(n34707) );
  NOR U34815 ( .A(n37563), .B(n37561), .Z(n37562) );
  XOR U34816 ( .A(n37564), .B(n37565), .Z(n34710) );
  NOR U34817 ( .A(n37566), .B(n37564), .Z(n37565) );
  XOR U34818 ( .A(n37567), .B(n37568), .Z(n34713) );
  NOR U34819 ( .A(n37569), .B(n37567), .Z(n37568) );
  XOR U34820 ( .A(n37570), .B(n37571), .Z(n34716) );
  NOR U34821 ( .A(n37572), .B(n37570), .Z(n37571) );
  XOR U34822 ( .A(n37573), .B(n37574), .Z(n34719) );
  NOR U34823 ( .A(n37575), .B(n37573), .Z(n37574) );
  XOR U34824 ( .A(n37576), .B(n37577), .Z(n34722) );
  NOR U34825 ( .A(n37578), .B(n37576), .Z(n37577) );
  XOR U34826 ( .A(n37579), .B(n37580), .Z(n34725) );
  NOR U34827 ( .A(n37581), .B(n37579), .Z(n37580) );
  XOR U34828 ( .A(n37582), .B(n37583), .Z(n34728) );
  NOR U34829 ( .A(n37584), .B(n37582), .Z(n37583) );
  XOR U34830 ( .A(n37585), .B(n37586), .Z(n34731) );
  NOR U34831 ( .A(n37587), .B(n37585), .Z(n37586) );
  XOR U34832 ( .A(n37588), .B(n37589), .Z(n34734) );
  NOR U34833 ( .A(n37590), .B(n37588), .Z(n37589) );
  XOR U34834 ( .A(n37591), .B(n37592), .Z(n34737) );
  NOR U34835 ( .A(n37593), .B(n37591), .Z(n37592) );
  XOR U34836 ( .A(n37594), .B(n37595), .Z(n34740) );
  NOR U34837 ( .A(n37596), .B(n37594), .Z(n37595) );
  XOR U34838 ( .A(n37597), .B(n37598), .Z(n34743) );
  NOR U34839 ( .A(n37599), .B(n37597), .Z(n37598) );
  XOR U34840 ( .A(n37600), .B(n37601), .Z(n34746) );
  NOR U34841 ( .A(n37602), .B(n37600), .Z(n37601) );
  XOR U34842 ( .A(n37603), .B(n37604), .Z(n34749) );
  NOR U34843 ( .A(n37605), .B(n37603), .Z(n37604) );
  XOR U34844 ( .A(n37606), .B(n37607), .Z(n34752) );
  NOR U34845 ( .A(n37608), .B(n37606), .Z(n37607) );
  XOR U34846 ( .A(n37609), .B(n37610), .Z(n34755) );
  NOR U34847 ( .A(n37611), .B(n37609), .Z(n37610) );
  XOR U34848 ( .A(n37612), .B(n37613), .Z(n34758) );
  NOR U34849 ( .A(n37614), .B(n37612), .Z(n37613) );
  XOR U34850 ( .A(n37615), .B(n37616), .Z(n34761) );
  NOR U34851 ( .A(n37617), .B(n37615), .Z(n37616) );
  XOR U34852 ( .A(n37618), .B(n37619), .Z(n34764) );
  NOR U34853 ( .A(n37620), .B(n37618), .Z(n37619) );
  XOR U34854 ( .A(n37621), .B(n37622), .Z(n34767) );
  NOR U34855 ( .A(n37623), .B(n37621), .Z(n37622) );
  XOR U34856 ( .A(n37624), .B(n37625), .Z(n34770) );
  NOR U34857 ( .A(n37626), .B(n37624), .Z(n37625) );
  XOR U34858 ( .A(n37627), .B(n37628), .Z(n34773) );
  NOR U34859 ( .A(n37629), .B(n37627), .Z(n37628) );
  XOR U34860 ( .A(n37630), .B(n37631), .Z(n34776) );
  NOR U34861 ( .A(n37632), .B(n37630), .Z(n37631) );
  XOR U34862 ( .A(n37633), .B(n37634), .Z(n34779) );
  NOR U34863 ( .A(n37635), .B(n37633), .Z(n37634) );
  XOR U34864 ( .A(n37636), .B(n37637), .Z(n34782) );
  NOR U34865 ( .A(n37638), .B(n37636), .Z(n37637) );
  XOR U34866 ( .A(n37639), .B(n37640), .Z(n34785) );
  NOR U34867 ( .A(n37641), .B(n37639), .Z(n37640) );
  XOR U34868 ( .A(n37642), .B(n37643), .Z(n34788) );
  NOR U34869 ( .A(n37644), .B(n37642), .Z(n37643) );
  XOR U34870 ( .A(n37645), .B(n37646), .Z(n34791) );
  NOR U34871 ( .A(n37647), .B(n37645), .Z(n37646) );
  XOR U34872 ( .A(n37648), .B(n37649), .Z(n34794) );
  NOR U34873 ( .A(n37650), .B(n37648), .Z(n37649) );
  XOR U34874 ( .A(n37651), .B(n37652), .Z(n34797) );
  NOR U34875 ( .A(n37653), .B(n37651), .Z(n37652) );
  XOR U34876 ( .A(n37654), .B(n37655), .Z(n34800) );
  NOR U34877 ( .A(n37656), .B(n37654), .Z(n37655) );
  XOR U34878 ( .A(n37657), .B(n37658), .Z(n34803) );
  NOR U34879 ( .A(n37659), .B(n37657), .Z(n37658) );
  XOR U34880 ( .A(n37660), .B(n37661), .Z(n34806) );
  NOR U34881 ( .A(n37662), .B(n37660), .Z(n37661) );
  XOR U34882 ( .A(n37663), .B(n37664), .Z(n34809) );
  NOR U34883 ( .A(n37665), .B(n37663), .Z(n37664) );
  XOR U34884 ( .A(n37666), .B(n37667), .Z(n34812) );
  NOR U34885 ( .A(n37668), .B(n37666), .Z(n37667) );
  XOR U34886 ( .A(n37669), .B(n37670), .Z(n34815) );
  NOR U34887 ( .A(n37671), .B(n37669), .Z(n37670) );
  XOR U34888 ( .A(n37672), .B(n37673), .Z(n34818) );
  NOR U34889 ( .A(n37674), .B(n37672), .Z(n37673) );
  XOR U34890 ( .A(n37675), .B(n37676), .Z(n34821) );
  NOR U34891 ( .A(n37677), .B(n37675), .Z(n37676) );
  XOR U34892 ( .A(n37678), .B(n37679), .Z(n34824) );
  NOR U34893 ( .A(n37680), .B(n37678), .Z(n37679) );
  XOR U34894 ( .A(n37681), .B(n37682), .Z(n34827) );
  NOR U34895 ( .A(n37683), .B(n37681), .Z(n37682) );
  XOR U34896 ( .A(n37684), .B(n37685), .Z(n34830) );
  NOR U34897 ( .A(n37686), .B(n37684), .Z(n37685) );
  XOR U34898 ( .A(n37687), .B(n37688), .Z(n34833) );
  NOR U34899 ( .A(n37689), .B(n37687), .Z(n37688) );
  XOR U34900 ( .A(n37690), .B(n37691), .Z(n34836) );
  NOR U34901 ( .A(n37692), .B(n37690), .Z(n37691) );
  XOR U34902 ( .A(n37693), .B(n37694), .Z(n34839) );
  NOR U34903 ( .A(n37695), .B(n37693), .Z(n37694) );
  XOR U34904 ( .A(n37696), .B(n37697), .Z(n34842) );
  NOR U34905 ( .A(n37698), .B(n37696), .Z(n37697) );
  XOR U34906 ( .A(n37699), .B(n37700), .Z(n34845) );
  NOR U34907 ( .A(n37701), .B(n37699), .Z(n37700) );
  XOR U34908 ( .A(n37702), .B(n37703), .Z(n34848) );
  NOR U34909 ( .A(n37704), .B(n37702), .Z(n37703) );
  XOR U34910 ( .A(n37705), .B(n37706), .Z(n34851) );
  NOR U34911 ( .A(n37707), .B(n37705), .Z(n37706) );
  XOR U34912 ( .A(n37708), .B(n37709), .Z(n34854) );
  NOR U34913 ( .A(n37710), .B(n37708), .Z(n37709) );
  XOR U34914 ( .A(n37711), .B(n37712), .Z(n34857) );
  NOR U34915 ( .A(n37713), .B(n37711), .Z(n37712) );
  XOR U34916 ( .A(n37714), .B(n37715), .Z(n34860) );
  NOR U34917 ( .A(n37716), .B(n37714), .Z(n37715) );
  XOR U34918 ( .A(n37717), .B(n37718), .Z(n34863) );
  NOR U34919 ( .A(n37719), .B(n37717), .Z(n37718) );
  XOR U34920 ( .A(n37720), .B(n37721), .Z(n34866) );
  NOR U34921 ( .A(n37722), .B(n37720), .Z(n37721) );
  XOR U34922 ( .A(n37723), .B(n37724), .Z(n34869) );
  NOR U34923 ( .A(n37725), .B(n37723), .Z(n37724) );
  XOR U34924 ( .A(n37726), .B(n37727), .Z(n34872) );
  NOR U34925 ( .A(n37728), .B(n37726), .Z(n37727) );
  XOR U34926 ( .A(n37729), .B(n37730), .Z(n34875) );
  NOR U34927 ( .A(n37731), .B(n37729), .Z(n37730) );
  XOR U34928 ( .A(n37732), .B(n37733), .Z(n34878) );
  NOR U34929 ( .A(n37734), .B(n37732), .Z(n37733) );
  XOR U34930 ( .A(n37735), .B(n37736), .Z(n34881) );
  NOR U34931 ( .A(n37737), .B(n37735), .Z(n37736) );
  XOR U34932 ( .A(n37738), .B(n37739), .Z(n34884) );
  NOR U34933 ( .A(n37740), .B(n37738), .Z(n37739) );
  XOR U34934 ( .A(n37741), .B(n37742), .Z(n34887) );
  NOR U34935 ( .A(n37743), .B(n37741), .Z(n37742) );
  XOR U34936 ( .A(n37744), .B(n37745), .Z(n34890) );
  NOR U34937 ( .A(n37746), .B(n37744), .Z(n37745) );
  XOR U34938 ( .A(n37747), .B(n37748), .Z(n34893) );
  NOR U34939 ( .A(n37749), .B(n37747), .Z(n37748) );
  XOR U34940 ( .A(n37750), .B(n37751), .Z(n34896) );
  NOR U34941 ( .A(n37752), .B(n37750), .Z(n37751) );
  XOR U34942 ( .A(n37753), .B(n37754), .Z(n34899) );
  NOR U34943 ( .A(n37755), .B(n37753), .Z(n37754) );
  XOR U34944 ( .A(n37756), .B(n37757), .Z(n34902) );
  NOR U34945 ( .A(n37758), .B(n37756), .Z(n37757) );
  XOR U34946 ( .A(n37759), .B(n37760), .Z(n34905) );
  NOR U34947 ( .A(n37761), .B(n37759), .Z(n37760) );
  XOR U34948 ( .A(n37762), .B(n37763), .Z(n34908) );
  NOR U34949 ( .A(n37764), .B(n37762), .Z(n37763) );
  XOR U34950 ( .A(n37765), .B(n37766), .Z(n34911) );
  NOR U34951 ( .A(n37767), .B(n37765), .Z(n37766) );
  XOR U34952 ( .A(n37768), .B(n37769), .Z(n34914) );
  NOR U34953 ( .A(n37770), .B(n37768), .Z(n37769) );
  XOR U34954 ( .A(n37771), .B(n37772), .Z(n34917) );
  NOR U34955 ( .A(n37773), .B(n37771), .Z(n37772) );
  XOR U34956 ( .A(n37774), .B(n37775), .Z(n34920) );
  NOR U34957 ( .A(n37776), .B(n37774), .Z(n37775) );
  XOR U34958 ( .A(n37777), .B(n37778), .Z(n34923) );
  NOR U34959 ( .A(n37779), .B(n37777), .Z(n37778) );
  XOR U34960 ( .A(n37780), .B(n37781), .Z(n34926) );
  NOR U34961 ( .A(n37782), .B(n37780), .Z(n37781) );
  XOR U34962 ( .A(n37783), .B(n37784), .Z(n34929) );
  NOR U34963 ( .A(n37785), .B(n37783), .Z(n37784) );
  XOR U34964 ( .A(n37786), .B(n37787), .Z(n34932) );
  NOR U34965 ( .A(n37788), .B(n37786), .Z(n37787) );
  XOR U34966 ( .A(n37789), .B(n37790), .Z(n34935) );
  NOR U34967 ( .A(n37791), .B(n37789), .Z(n37790) );
  XOR U34968 ( .A(n37792), .B(n37793), .Z(n34938) );
  NOR U34969 ( .A(n37794), .B(n37792), .Z(n37793) );
  XOR U34970 ( .A(n37795), .B(n37796), .Z(n34941) );
  NOR U34971 ( .A(n37797), .B(n37795), .Z(n37796) );
  XOR U34972 ( .A(n37798), .B(n37799), .Z(n34944) );
  NOR U34973 ( .A(n37800), .B(n37798), .Z(n37799) );
  XOR U34974 ( .A(n37801), .B(n37802), .Z(n34947) );
  NOR U34975 ( .A(n37803), .B(n37801), .Z(n37802) );
  XOR U34976 ( .A(n37804), .B(n37805), .Z(n34950) );
  NOR U34977 ( .A(n37806), .B(n37804), .Z(n37805) );
  XOR U34978 ( .A(n37807), .B(n37808), .Z(n34953) );
  NOR U34979 ( .A(n37809), .B(n37807), .Z(n37808) );
  XOR U34980 ( .A(n37810), .B(n37811), .Z(n34956) );
  NOR U34981 ( .A(n37812), .B(n37810), .Z(n37811) );
  XOR U34982 ( .A(n37813), .B(n37814), .Z(n34959) );
  NOR U34983 ( .A(n37815), .B(n37813), .Z(n37814) );
  XOR U34984 ( .A(n37816), .B(n37817), .Z(n34962) );
  NOR U34985 ( .A(n37818), .B(n37816), .Z(n37817) );
  XOR U34986 ( .A(n37819), .B(n37820), .Z(n34965) );
  NOR U34987 ( .A(n37821), .B(n37819), .Z(n37820) );
  XOR U34988 ( .A(n37822), .B(n37823), .Z(n34968) );
  NOR U34989 ( .A(n37824), .B(n37822), .Z(n37823) );
  XOR U34990 ( .A(n37825), .B(n37826), .Z(n34971) );
  NOR U34991 ( .A(n37827), .B(n37825), .Z(n37826) );
  XOR U34992 ( .A(n37828), .B(n37829), .Z(n34974) );
  NOR U34993 ( .A(n37830), .B(n37828), .Z(n37829) );
  XOR U34994 ( .A(n37831), .B(n37832), .Z(n34977) );
  NOR U34995 ( .A(n37833), .B(n37831), .Z(n37832) );
  XOR U34996 ( .A(n37834), .B(n37835), .Z(n34980) );
  NOR U34997 ( .A(n37836), .B(n37834), .Z(n37835) );
  XOR U34998 ( .A(n37837), .B(n37838), .Z(n34983) );
  NOR U34999 ( .A(n37839), .B(n37837), .Z(n37838) );
  XOR U35000 ( .A(n37840), .B(n37841), .Z(n34986) );
  NOR U35001 ( .A(n37842), .B(n37840), .Z(n37841) );
  XOR U35002 ( .A(n37843), .B(n37844), .Z(n34989) );
  NOR U35003 ( .A(n37845), .B(n37843), .Z(n37844) );
  XOR U35004 ( .A(n37846), .B(n37847), .Z(n34992) );
  NOR U35005 ( .A(n37848), .B(n37846), .Z(n37847) );
  XOR U35006 ( .A(n37849), .B(n37850), .Z(n34995) );
  NOR U35007 ( .A(n37851), .B(n37849), .Z(n37850) );
  XOR U35008 ( .A(n37852), .B(n37853), .Z(n34998) );
  NOR U35009 ( .A(n37854), .B(n37852), .Z(n37853) );
  XOR U35010 ( .A(n37855), .B(n37856), .Z(n35001) );
  NOR U35011 ( .A(n37857), .B(n37855), .Z(n37856) );
  XOR U35012 ( .A(n37858), .B(n37859), .Z(n35004) );
  NOR U35013 ( .A(n37860), .B(n37858), .Z(n37859) );
  XOR U35014 ( .A(n37861), .B(n37862), .Z(n35007) );
  NOR U35015 ( .A(n37863), .B(n37861), .Z(n37862) );
  XOR U35016 ( .A(n37864), .B(n37865), .Z(n35010) );
  NOR U35017 ( .A(n37866), .B(n37864), .Z(n37865) );
  XOR U35018 ( .A(n37867), .B(n37868), .Z(n35013) );
  NOR U35019 ( .A(n37869), .B(n37867), .Z(n37868) );
  XOR U35020 ( .A(n37870), .B(n37871), .Z(n35016) );
  NOR U35021 ( .A(n37872), .B(n37870), .Z(n37871) );
  XOR U35022 ( .A(n37873), .B(n37874), .Z(n35019) );
  NOR U35023 ( .A(n37875), .B(n37873), .Z(n37874) );
  XOR U35024 ( .A(n37876), .B(n37877), .Z(n35022) );
  NOR U35025 ( .A(n37878), .B(n37876), .Z(n37877) );
  XOR U35026 ( .A(n37879), .B(n37880), .Z(n35025) );
  NOR U35027 ( .A(n37881), .B(n37879), .Z(n37880) );
  XOR U35028 ( .A(n37882), .B(n37883), .Z(n35028) );
  NOR U35029 ( .A(n37884), .B(n37882), .Z(n37883) );
  XOR U35030 ( .A(n37885), .B(n37886), .Z(n35031) );
  NOR U35031 ( .A(n37887), .B(n37885), .Z(n37886) );
  XOR U35032 ( .A(n37888), .B(n37889), .Z(n35034) );
  NOR U35033 ( .A(n37890), .B(n37888), .Z(n37889) );
  XOR U35034 ( .A(n37891), .B(n37892), .Z(n35037) );
  NOR U35035 ( .A(n37893), .B(n37891), .Z(n37892) );
  XOR U35036 ( .A(n37894), .B(n37895), .Z(n35040) );
  NOR U35037 ( .A(n37896), .B(n37894), .Z(n37895) );
  XOR U35038 ( .A(n37897), .B(n37898), .Z(n35043) );
  NOR U35039 ( .A(n37899), .B(n37897), .Z(n37898) );
  XOR U35040 ( .A(n37900), .B(n37901), .Z(n35046) );
  NOR U35041 ( .A(n37902), .B(n37900), .Z(n37901) );
  XOR U35042 ( .A(n37903), .B(n37904), .Z(n35049) );
  NOR U35043 ( .A(n37905), .B(n37903), .Z(n37904) );
  XOR U35044 ( .A(n37906), .B(n37907), .Z(n35052) );
  NOR U35045 ( .A(n37908), .B(n37906), .Z(n37907) );
  XOR U35046 ( .A(n37909), .B(n37910), .Z(n35055) );
  NOR U35047 ( .A(n37911), .B(n37909), .Z(n37910) );
  XOR U35048 ( .A(n37912), .B(n37913), .Z(n35058) );
  NOR U35049 ( .A(n37914), .B(n37912), .Z(n37913) );
  XOR U35050 ( .A(n37915), .B(n37916), .Z(n35061) );
  NOR U35051 ( .A(n37917), .B(n37915), .Z(n37916) );
  XOR U35052 ( .A(n37918), .B(n37919), .Z(n35064) );
  NOR U35053 ( .A(n37920), .B(n37918), .Z(n37919) );
  XOR U35054 ( .A(n37921), .B(n37922), .Z(n35067) );
  NOR U35055 ( .A(n37923), .B(n37921), .Z(n37922) );
  XOR U35056 ( .A(n37924), .B(n37925), .Z(n35070) );
  NOR U35057 ( .A(n37926), .B(n37924), .Z(n37925) );
  XOR U35058 ( .A(n37927), .B(n37928), .Z(n35073) );
  NOR U35059 ( .A(n37929), .B(n37927), .Z(n37928) );
  XOR U35060 ( .A(n37930), .B(n37931), .Z(n35076) );
  NOR U35061 ( .A(n37932), .B(n37930), .Z(n37931) );
  XOR U35062 ( .A(n37933), .B(n37934), .Z(n35079) );
  NOR U35063 ( .A(n37935), .B(n37933), .Z(n37934) );
  XOR U35064 ( .A(n37936), .B(n37937), .Z(n35082) );
  NOR U35065 ( .A(n37938), .B(n37936), .Z(n37937) );
  XOR U35066 ( .A(n37939), .B(n37940), .Z(n35085) );
  NOR U35067 ( .A(n37941), .B(n37939), .Z(n37940) );
  XOR U35068 ( .A(n37942), .B(n37943), .Z(n35088) );
  NOR U35069 ( .A(n37944), .B(n37942), .Z(n37943) );
  XOR U35070 ( .A(n37945), .B(n37946), .Z(n35091) );
  NOR U35071 ( .A(n37947), .B(n37945), .Z(n37946) );
  XOR U35072 ( .A(n37948), .B(n37949), .Z(n35094) );
  NOR U35073 ( .A(n37950), .B(n37948), .Z(n37949) );
  XOR U35074 ( .A(n37951), .B(n37952), .Z(n35097) );
  NOR U35075 ( .A(n37953), .B(n37951), .Z(n37952) );
  XOR U35076 ( .A(n37954), .B(n37955), .Z(n35100) );
  NOR U35077 ( .A(n37956), .B(n37954), .Z(n37955) );
  XOR U35078 ( .A(n37957), .B(n37958), .Z(n35103) );
  NOR U35079 ( .A(n37959), .B(n37957), .Z(n37958) );
  XOR U35080 ( .A(n37960), .B(n37961), .Z(n35106) );
  NOR U35081 ( .A(n37962), .B(n37960), .Z(n37961) );
  XOR U35082 ( .A(n37963), .B(n37964), .Z(n35109) );
  NOR U35083 ( .A(n37965), .B(n37963), .Z(n37964) );
  XOR U35084 ( .A(n37966), .B(n37967), .Z(n35112) );
  NOR U35085 ( .A(n37968), .B(n37966), .Z(n37967) );
  XOR U35086 ( .A(n37969), .B(n37970), .Z(n35115) );
  NOR U35087 ( .A(n37971), .B(n37969), .Z(n37970) );
  XOR U35088 ( .A(n37972), .B(n37973), .Z(n35118) );
  NOR U35089 ( .A(n37974), .B(n37972), .Z(n37973) );
  XOR U35090 ( .A(n37975), .B(n37976), .Z(n35121) );
  NOR U35091 ( .A(n37977), .B(n37975), .Z(n37976) );
  XOR U35092 ( .A(n37978), .B(n37979), .Z(n35124) );
  NOR U35093 ( .A(n37980), .B(n37978), .Z(n37979) );
  XOR U35094 ( .A(n37981), .B(n37982), .Z(n35127) );
  NOR U35095 ( .A(n37983), .B(n37981), .Z(n37982) );
  XOR U35096 ( .A(n37984), .B(n37985), .Z(n35130) );
  NOR U35097 ( .A(n37986), .B(n37984), .Z(n37985) );
  XOR U35098 ( .A(n37987), .B(n37988), .Z(n35133) );
  NOR U35099 ( .A(n37989), .B(n37987), .Z(n37988) );
  XOR U35100 ( .A(n37990), .B(n37991), .Z(n35136) );
  NOR U35101 ( .A(n37992), .B(n37990), .Z(n37991) );
  XOR U35102 ( .A(n37993), .B(n37994), .Z(n35139) );
  NOR U35103 ( .A(n37995), .B(n37993), .Z(n37994) );
  XOR U35104 ( .A(n37996), .B(n37997), .Z(n35142) );
  NOR U35105 ( .A(n37998), .B(n37996), .Z(n37997) );
  XOR U35106 ( .A(n37999), .B(n38000), .Z(n35145) );
  NOR U35107 ( .A(n38001), .B(n37999), .Z(n38000) );
  XOR U35108 ( .A(n38002), .B(n38003), .Z(n35148) );
  NOR U35109 ( .A(n38004), .B(n38002), .Z(n38003) );
  XOR U35110 ( .A(n38005), .B(n38006), .Z(n35151) );
  NOR U35111 ( .A(n38007), .B(n38005), .Z(n38006) );
  XOR U35112 ( .A(n38008), .B(n38009), .Z(n35154) );
  NOR U35113 ( .A(n38010), .B(n38008), .Z(n38009) );
  XOR U35114 ( .A(n38011), .B(n38012), .Z(n35157) );
  NOR U35115 ( .A(n38013), .B(n38011), .Z(n38012) );
  XOR U35116 ( .A(n38014), .B(n38015), .Z(n35160) );
  NOR U35117 ( .A(n38016), .B(n38014), .Z(n38015) );
  XOR U35118 ( .A(n38017), .B(n38018), .Z(n35163) );
  NOR U35119 ( .A(n38019), .B(n38017), .Z(n38018) );
  XOR U35120 ( .A(n38020), .B(n38021), .Z(n35166) );
  NOR U35121 ( .A(n38022), .B(n38020), .Z(n38021) );
  XOR U35122 ( .A(n38023), .B(n38024), .Z(n35169) );
  NOR U35123 ( .A(n38025), .B(n38023), .Z(n38024) );
  XOR U35124 ( .A(n38026), .B(n38027), .Z(n35172) );
  NOR U35125 ( .A(n38028), .B(n38026), .Z(n38027) );
  XOR U35126 ( .A(n38029), .B(n38030), .Z(n35175) );
  NOR U35127 ( .A(n38031), .B(n38029), .Z(n38030) );
  XOR U35128 ( .A(n38032), .B(n38033), .Z(n35178) );
  NOR U35129 ( .A(n38034), .B(n38032), .Z(n38033) );
  XOR U35130 ( .A(n38035), .B(n38036), .Z(n35181) );
  NOR U35131 ( .A(n38037), .B(n38035), .Z(n38036) );
  XOR U35132 ( .A(n38038), .B(n38039), .Z(n35184) );
  NOR U35133 ( .A(n38040), .B(n38038), .Z(n38039) );
  XOR U35134 ( .A(n38041), .B(n38042), .Z(n35187) );
  NOR U35135 ( .A(n38043), .B(n38041), .Z(n38042) );
  XOR U35136 ( .A(n38044), .B(n38045), .Z(n35190) );
  NOR U35137 ( .A(n38046), .B(n38044), .Z(n38045) );
  XOR U35138 ( .A(n38047), .B(n38048), .Z(n35193) );
  NOR U35139 ( .A(n38049), .B(n38047), .Z(n38048) );
  XOR U35140 ( .A(n38050), .B(n38051), .Z(n35196) );
  NOR U35141 ( .A(n38052), .B(n38050), .Z(n38051) );
  XOR U35142 ( .A(n38053), .B(n38054), .Z(n35199) );
  NOR U35143 ( .A(n38055), .B(n38053), .Z(n38054) );
  XOR U35144 ( .A(n38056), .B(n38057), .Z(n35202) );
  NOR U35145 ( .A(n38058), .B(n38056), .Z(n38057) );
  XOR U35146 ( .A(n38059), .B(n38060), .Z(n35205) );
  NOR U35147 ( .A(n38061), .B(n38059), .Z(n38060) );
  XOR U35148 ( .A(n38062), .B(n38063), .Z(n35208) );
  NOR U35149 ( .A(n38064), .B(n38062), .Z(n38063) );
  XOR U35150 ( .A(n38065), .B(n38066), .Z(n35211) );
  NOR U35151 ( .A(n38067), .B(n38065), .Z(n38066) );
  XOR U35152 ( .A(n38068), .B(n38069), .Z(n35214) );
  NOR U35153 ( .A(n38070), .B(n38068), .Z(n38069) );
  XOR U35154 ( .A(n38071), .B(n38072), .Z(n35217) );
  NOR U35155 ( .A(n38073), .B(n38071), .Z(n38072) );
  XOR U35156 ( .A(n38074), .B(n38075), .Z(n35220) );
  NOR U35157 ( .A(n38076), .B(n38074), .Z(n38075) );
  XOR U35158 ( .A(n38077), .B(n38078), .Z(n35223) );
  NOR U35159 ( .A(n38079), .B(n38077), .Z(n38078) );
  XOR U35160 ( .A(n38080), .B(n38081), .Z(n35226) );
  NOR U35161 ( .A(n38082), .B(n38080), .Z(n38081) );
  XOR U35162 ( .A(n38083), .B(n38084), .Z(n35229) );
  NOR U35163 ( .A(n38085), .B(n38083), .Z(n38084) );
  XOR U35164 ( .A(n38086), .B(n38087), .Z(n35232) );
  NOR U35165 ( .A(n38088), .B(n38086), .Z(n38087) );
  XOR U35166 ( .A(n38089), .B(n38090), .Z(n35235) );
  NOR U35167 ( .A(n38091), .B(n38089), .Z(n38090) );
  XOR U35168 ( .A(n38092), .B(n38093), .Z(n35238) );
  NOR U35169 ( .A(n38094), .B(n38092), .Z(n38093) );
  XOR U35170 ( .A(n38095), .B(n38096), .Z(n35241) );
  NOR U35171 ( .A(n38097), .B(n38095), .Z(n38096) );
  XOR U35172 ( .A(n38098), .B(n38099), .Z(n35244) );
  NOR U35173 ( .A(n38100), .B(n38098), .Z(n38099) );
  XOR U35174 ( .A(n38101), .B(n38102), .Z(n35247) );
  NOR U35175 ( .A(n38103), .B(n38101), .Z(n38102) );
  XOR U35176 ( .A(n38104), .B(n38105), .Z(n35250) );
  NOR U35177 ( .A(n38106), .B(n38104), .Z(n38105) );
  XOR U35178 ( .A(n38107), .B(n38108), .Z(n35253) );
  NOR U35179 ( .A(n38109), .B(n38107), .Z(n38108) );
  XOR U35180 ( .A(n38110), .B(n38111), .Z(n35256) );
  NOR U35181 ( .A(n38112), .B(n38110), .Z(n38111) );
  XOR U35182 ( .A(n38113), .B(n38114), .Z(n35259) );
  NOR U35183 ( .A(n38115), .B(n38113), .Z(n38114) );
  XOR U35184 ( .A(n38116), .B(n38117), .Z(n35262) );
  NOR U35185 ( .A(n38118), .B(n38116), .Z(n38117) );
  XOR U35186 ( .A(n38119), .B(n38120), .Z(n35265) );
  NOR U35187 ( .A(n38121), .B(n38119), .Z(n38120) );
  XOR U35188 ( .A(n38122), .B(n38123), .Z(n35268) );
  NOR U35189 ( .A(n38124), .B(n38122), .Z(n38123) );
  XOR U35190 ( .A(n38125), .B(n38126), .Z(n35271) );
  NOR U35191 ( .A(n38127), .B(n38125), .Z(n38126) );
  XOR U35192 ( .A(n38128), .B(n38129), .Z(n35274) );
  NOR U35193 ( .A(n38130), .B(n38128), .Z(n38129) );
  XOR U35194 ( .A(n38131), .B(n38132), .Z(n35277) );
  NOR U35195 ( .A(n38133), .B(n38131), .Z(n38132) );
  XOR U35196 ( .A(n38134), .B(n38135), .Z(n35280) );
  NOR U35197 ( .A(n38136), .B(n38134), .Z(n38135) );
  XOR U35198 ( .A(n38137), .B(n38138), .Z(n35283) );
  NOR U35199 ( .A(n38139), .B(n38137), .Z(n38138) );
  XOR U35200 ( .A(n38140), .B(n38141), .Z(n35286) );
  NOR U35201 ( .A(n38142), .B(n38140), .Z(n38141) );
  XOR U35202 ( .A(n38143), .B(n38144), .Z(n35289) );
  NOR U35203 ( .A(n38145), .B(n38143), .Z(n38144) );
  XOR U35204 ( .A(n38146), .B(n38147), .Z(n35292) );
  NOR U35205 ( .A(n38148), .B(n38146), .Z(n38147) );
  XOR U35206 ( .A(n38149), .B(n38150), .Z(n35295) );
  NOR U35207 ( .A(n38151), .B(n38149), .Z(n38150) );
  XOR U35208 ( .A(n38152), .B(n38153), .Z(n35298) );
  NOR U35209 ( .A(n38154), .B(n38152), .Z(n38153) );
  XOR U35210 ( .A(n38155), .B(n38156), .Z(n35301) );
  NOR U35211 ( .A(n38157), .B(n38155), .Z(n38156) );
  XOR U35212 ( .A(n38158), .B(n38159), .Z(n35304) );
  NOR U35213 ( .A(n38160), .B(n38158), .Z(n38159) );
  XOR U35214 ( .A(n38161), .B(n38162), .Z(n35307) );
  NOR U35215 ( .A(n38163), .B(n38161), .Z(n38162) );
  XOR U35216 ( .A(n38164), .B(n38165), .Z(n35310) );
  NOR U35217 ( .A(n38166), .B(n38164), .Z(n38165) );
  XOR U35218 ( .A(n38167), .B(n38168), .Z(n35313) );
  NOR U35219 ( .A(n38169), .B(n38167), .Z(n38168) );
  XOR U35220 ( .A(n38170), .B(n38171), .Z(n35316) );
  NOR U35221 ( .A(n38172), .B(n38170), .Z(n38171) );
  XOR U35222 ( .A(n38173), .B(n38174), .Z(n35319) );
  NOR U35223 ( .A(n38175), .B(n38173), .Z(n38174) );
  XOR U35224 ( .A(n38176), .B(n38177), .Z(n35322) );
  NOR U35225 ( .A(n38178), .B(n38176), .Z(n38177) );
  XOR U35226 ( .A(n38179), .B(n38180), .Z(n35325) );
  NOR U35227 ( .A(n38181), .B(n38179), .Z(n38180) );
  XOR U35228 ( .A(n38182), .B(n38183), .Z(n35328) );
  NOR U35229 ( .A(n38184), .B(n38182), .Z(n38183) );
  XOR U35230 ( .A(n38185), .B(n38186), .Z(n35331) );
  NOR U35231 ( .A(n38187), .B(n38185), .Z(n38186) );
  XOR U35232 ( .A(n38188), .B(n38189), .Z(n35334) );
  NOR U35233 ( .A(n38190), .B(n38188), .Z(n38189) );
  XOR U35234 ( .A(n38191), .B(n38192), .Z(n35337) );
  NOR U35235 ( .A(n38193), .B(n38191), .Z(n38192) );
  XOR U35236 ( .A(n38194), .B(n38195), .Z(n35340) );
  NOR U35237 ( .A(n38196), .B(n38194), .Z(n38195) );
  XOR U35238 ( .A(n38197), .B(n38198), .Z(n35343) );
  NOR U35239 ( .A(n38199), .B(n38197), .Z(n38198) );
  XOR U35240 ( .A(n38200), .B(n38201), .Z(n35346) );
  NOR U35241 ( .A(n38202), .B(n38200), .Z(n38201) );
  XOR U35242 ( .A(n38203), .B(n38204), .Z(n35349) );
  NOR U35243 ( .A(n38205), .B(n38203), .Z(n38204) );
  XOR U35244 ( .A(n38206), .B(n38207), .Z(n35352) );
  NOR U35245 ( .A(n38208), .B(n38206), .Z(n38207) );
  XOR U35246 ( .A(n38209), .B(n38210), .Z(n35355) );
  NOR U35247 ( .A(n38211), .B(n38209), .Z(n38210) );
  XOR U35248 ( .A(n38212), .B(n38213), .Z(n35358) );
  NOR U35249 ( .A(n38214), .B(n38212), .Z(n38213) );
  XOR U35250 ( .A(n38215), .B(n38216), .Z(n35361) );
  NOR U35251 ( .A(n38217), .B(n38215), .Z(n38216) );
  XOR U35252 ( .A(n38218), .B(n38219), .Z(n35364) );
  NOR U35253 ( .A(n38220), .B(n38218), .Z(n38219) );
  XOR U35254 ( .A(n38221), .B(n38222), .Z(n35367) );
  NOR U35255 ( .A(n38223), .B(n38221), .Z(n38222) );
  XOR U35256 ( .A(n38224), .B(n38225), .Z(n35370) );
  NOR U35257 ( .A(n38226), .B(n38224), .Z(n38225) );
  XOR U35258 ( .A(n38227), .B(n38228), .Z(n35373) );
  NOR U35259 ( .A(n38229), .B(n38227), .Z(n38228) );
  XOR U35260 ( .A(n38230), .B(n38231), .Z(n35376) );
  NOR U35261 ( .A(n38232), .B(n38230), .Z(n38231) );
  XOR U35262 ( .A(n38233), .B(n38234), .Z(n35379) );
  NOR U35263 ( .A(n38235), .B(n38233), .Z(n38234) );
  XOR U35264 ( .A(n38236), .B(n38237), .Z(n35382) );
  NOR U35265 ( .A(n38238), .B(n38236), .Z(n38237) );
  XOR U35266 ( .A(n38239), .B(n38240), .Z(n35385) );
  NOR U35267 ( .A(n38241), .B(n38239), .Z(n38240) );
  XOR U35268 ( .A(n38242), .B(n38243), .Z(n35388) );
  NOR U35269 ( .A(n38244), .B(n38242), .Z(n38243) );
  XOR U35270 ( .A(n38245), .B(n38246), .Z(n35391) );
  NOR U35271 ( .A(n38247), .B(n38245), .Z(n38246) );
  XOR U35272 ( .A(n38248), .B(n38249), .Z(n35394) );
  NOR U35273 ( .A(n38250), .B(n38248), .Z(n38249) );
  XOR U35274 ( .A(n38251), .B(n38252), .Z(n35397) );
  NOR U35275 ( .A(n38253), .B(n38251), .Z(n38252) );
  XOR U35276 ( .A(n38254), .B(n38255), .Z(n35400) );
  NOR U35277 ( .A(n38256), .B(n38254), .Z(n38255) );
  XOR U35278 ( .A(n38257), .B(n38258), .Z(n35403) );
  NOR U35279 ( .A(n38259), .B(n38257), .Z(n38258) );
  XOR U35280 ( .A(n38260), .B(n38261), .Z(n35406) );
  NOR U35281 ( .A(n38262), .B(n38260), .Z(n38261) );
  XOR U35282 ( .A(n38263), .B(n38264), .Z(n35409) );
  NOR U35283 ( .A(n38265), .B(n38263), .Z(n38264) );
  XOR U35284 ( .A(n38266), .B(n38267), .Z(n35412) );
  NOR U35285 ( .A(n38268), .B(n38266), .Z(n38267) );
  XOR U35286 ( .A(n38269), .B(n38270), .Z(n35415) );
  NOR U35287 ( .A(n38271), .B(n38269), .Z(n38270) );
  XOR U35288 ( .A(n38272), .B(n38273), .Z(n35418) );
  NOR U35289 ( .A(n38274), .B(n38272), .Z(n38273) );
  XOR U35290 ( .A(n38275), .B(n38276), .Z(n35421) );
  NOR U35291 ( .A(n38277), .B(n38275), .Z(n38276) );
  XOR U35292 ( .A(n38278), .B(n38279), .Z(n35424) );
  NOR U35293 ( .A(n38280), .B(n38278), .Z(n38279) );
  XOR U35294 ( .A(n38281), .B(n38282), .Z(n35427) );
  NOR U35295 ( .A(n38283), .B(n38281), .Z(n38282) );
  XOR U35296 ( .A(n38284), .B(n38285), .Z(n35430) );
  NOR U35297 ( .A(n38286), .B(n38284), .Z(n38285) );
  XOR U35298 ( .A(n38287), .B(n38288), .Z(n35433) );
  NOR U35299 ( .A(n38289), .B(n38287), .Z(n38288) );
  XOR U35300 ( .A(n38290), .B(n38291), .Z(n35436) );
  NOR U35301 ( .A(n38292), .B(n38290), .Z(n38291) );
  XOR U35302 ( .A(n38293), .B(n38294), .Z(n35439) );
  NOR U35303 ( .A(n38295), .B(n38293), .Z(n38294) );
  XOR U35304 ( .A(n38296), .B(n38297), .Z(n35442) );
  NOR U35305 ( .A(n38298), .B(n38296), .Z(n38297) );
  XOR U35306 ( .A(n38299), .B(n38300), .Z(n35445) );
  NOR U35307 ( .A(n38301), .B(n38299), .Z(n38300) );
  XOR U35308 ( .A(n38302), .B(n38303), .Z(n35448) );
  NOR U35309 ( .A(n38304), .B(n38302), .Z(n38303) );
  XOR U35310 ( .A(n38305), .B(n38306), .Z(n35451) );
  NOR U35311 ( .A(n38307), .B(n38305), .Z(n38306) );
  XOR U35312 ( .A(n38308), .B(n38309), .Z(n35454) );
  NOR U35313 ( .A(n38310), .B(n38308), .Z(n38309) );
  XOR U35314 ( .A(n38311), .B(n38312), .Z(n35457) );
  NOR U35315 ( .A(n38313), .B(n38311), .Z(n38312) );
  XOR U35316 ( .A(n38314), .B(n38315), .Z(n35460) );
  NOR U35317 ( .A(n38316), .B(n38314), .Z(n38315) );
  XOR U35318 ( .A(n38317), .B(n38318), .Z(n35463) );
  NOR U35319 ( .A(n38319), .B(n38317), .Z(n38318) );
  XOR U35320 ( .A(n38320), .B(n38321), .Z(n35466) );
  NOR U35321 ( .A(n38322), .B(n38320), .Z(n38321) );
  XOR U35322 ( .A(n38323), .B(n38324), .Z(n35469) );
  NOR U35323 ( .A(n38325), .B(n38323), .Z(n38324) );
  XOR U35324 ( .A(n38326), .B(n38327), .Z(n35472) );
  NOR U35325 ( .A(n38328), .B(n38326), .Z(n38327) );
  XOR U35326 ( .A(n38329), .B(n38330), .Z(n35475) );
  NOR U35327 ( .A(n38331), .B(n38329), .Z(n38330) );
  XOR U35328 ( .A(n38332), .B(n38333), .Z(n35478) );
  NOR U35329 ( .A(n38334), .B(n38332), .Z(n38333) );
  XOR U35330 ( .A(n38335), .B(n38336), .Z(n35481) );
  NOR U35331 ( .A(n38337), .B(n38335), .Z(n38336) );
  XOR U35332 ( .A(n38338), .B(n38339), .Z(n35484) );
  NOR U35333 ( .A(n38340), .B(n38338), .Z(n38339) );
  XOR U35334 ( .A(n38341), .B(n38342), .Z(n35487) );
  NOR U35335 ( .A(n38343), .B(n38341), .Z(n38342) );
  XOR U35336 ( .A(n38344), .B(n38345), .Z(n35490) );
  NOR U35337 ( .A(n38346), .B(n38344), .Z(n38345) );
  XOR U35338 ( .A(n38347), .B(n38348), .Z(n35493) );
  NOR U35339 ( .A(n38349), .B(n38347), .Z(n38348) );
  XOR U35340 ( .A(n38350), .B(n38351), .Z(n35496) );
  NOR U35341 ( .A(n38352), .B(n38350), .Z(n38351) );
  XOR U35342 ( .A(n38353), .B(n38354), .Z(n35499) );
  NOR U35343 ( .A(n38355), .B(n38353), .Z(n38354) );
  XOR U35344 ( .A(n38356), .B(n38357), .Z(n35502) );
  NOR U35345 ( .A(n38358), .B(n38356), .Z(n38357) );
  XOR U35346 ( .A(n38359), .B(n38360), .Z(n35505) );
  NOR U35347 ( .A(n38361), .B(n38359), .Z(n38360) );
  XOR U35348 ( .A(n38362), .B(n38363), .Z(n35508) );
  NOR U35349 ( .A(n38364), .B(n38362), .Z(n38363) );
  XOR U35350 ( .A(n38365), .B(n38366), .Z(n35511) );
  NOR U35351 ( .A(n38367), .B(n38365), .Z(n38366) );
  XOR U35352 ( .A(n38368), .B(n38369), .Z(n35514) );
  NOR U35353 ( .A(n38370), .B(n38368), .Z(n38369) );
  XOR U35354 ( .A(n38371), .B(n38372), .Z(n35517) );
  NOR U35355 ( .A(n38373), .B(n38371), .Z(n38372) );
  XOR U35356 ( .A(n38374), .B(n38375), .Z(n35520) );
  NOR U35357 ( .A(n38376), .B(n38374), .Z(n38375) );
  XOR U35358 ( .A(n38377), .B(n38378), .Z(n35523) );
  NOR U35359 ( .A(n38379), .B(n38377), .Z(n38378) );
  XOR U35360 ( .A(n38380), .B(n38381), .Z(n35526) );
  NOR U35361 ( .A(n38382), .B(n38380), .Z(n38381) );
  XNOR U35362 ( .A(n38383), .B(n38384), .Z(n35529) );
  NOR U35363 ( .A(n38385), .B(n38383), .Z(n38384) );
  XOR U35364 ( .A(n38386), .B(n38387), .Z(n35532) );
  AND U35365 ( .A(n124), .B(n38386), .Z(n38387) );
  XOR U35366 ( .A(n106), .B(n36963), .Z(n36965) );
  XOR U35367 ( .A(n36960), .B(n36959), .Z(n106) );
  XNOR U35368 ( .A(n36957), .B(n36956), .Z(n36959) );
  XNOR U35369 ( .A(n36954), .B(n36953), .Z(n36956) );
  XNOR U35370 ( .A(n36951), .B(n36950), .Z(n36953) );
  XNOR U35371 ( .A(n36948), .B(n36947), .Z(n36950) );
  XNOR U35372 ( .A(n36945), .B(n36944), .Z(n36947) );
  XNOR U35373 ( .A(n36942), .B(n36941), .Z(n36944) );
  XNOR U35374 ( .A(n36939), .B(n36938), .Z(n36941) );
  XNOR U35375 ( .A(n36936), .B(n36935), .Z(n36938) );
  XNOR U35376 ( .A(n36933), .B(n36932), .Z(n36935) );
  XNOR U35377 ( .A(n36930), .B(n36929), .Z(n36932) );
  XNOR U35378 ( .A(n36927), .B(n36926), .Z(n36929) );
  XNOR U35379 ( .A(n36924), .B(n36923), .Z(n36926) );
  XNOR U35380 ( .A(n36921), .B(n36920), .Z(n36923) );
  XNOR U35381 ( .A(n36918), .B(n36917), .Z(n36920) );
  XNOR U35382 ( .A(n36915), .B(n36914), .Z(n36917) );
  XNOR U35383 ( .A(n36912), .B(n36911), .Z(n36914) );
  XNOR U35384 ( .A(n36909), .B(n36908), .Z(n36911) );
  XNOR U35385 ( .A(n36906), .B(n36905), .Z(n36908) );
  XNOR U35386 ( .A(n36903), .B(n36902), .Z(n36905) );
  XNOR U35387 ( .A(n36900), .B(n36899), .Z(n36902) );
  XNOR U35388 ( .A(n36897), .B(n36896), .Z(n36899) );
  XNOR U35389 ( .A(n36894), .B(n36893), .Z(n36896) );
  XNOR U35390 ( .A(n36891), .B(n36890), .Z(n36893) );
  XNOR U35391 ( .A(n36888), .B(n36887), .Z(n36890) );
  XNOR U35392 ( .A(n36885), .B(n36884), .Z(n36887) );
  XNOR U35393 ( .A(n36882), .B(n36881), .Z(n36884) );
  XNOR U35394 ( .A(n36879), .B(n36878), .Z(n36881) );
  XNOR U35395 ( .A(n36876), .B(n36875), .Z(n36878) );
  XNOR U35396 ( .A(n36873), .B(n36872), .Z(n36875) );
  XNOR U35397 ( .A(n36870), .B(n36869), .Z(n36872) );
  XNOR U35398 ( .A(n36867), .B(n36866), .Z(n36869) );
  XNOR U35399 ( .A(n36864), .B(n36863), .Z(n36866) );
  XNOR U35400 ( .A(n36861), .B(n36860), .Z(n36863) );
  XNOR U35401 ( .A(n36858), .B(n36857), .Z(n36860) );
  XNOR U35402 ( .A(n36855), .B(n36854), .Z(n36857) );
  XNOR U35403 ( .A(n36852), .B(n36851), .Z(n36854) );
  XNOR U35404 ( .A(n36849), .B(n36848), .Z(n36851) );
  XNOR U35405 ( .A(n36846), .B(n36845), .Z(n36848) );
  XNOR U35406 ( .A(n36843), .B(n36842), .Z(n36845) );
  XNOR U35407 ( .A(n36840), .B(n36839), .Z(n36842) );
  XNOR U35408 ( .A(n36837), .B(n36836), .Z(n36839) );
  XNOR U35409 ( .A(n36834), .B(n36833), .Z(n36836) );
  XNOR U35410 ( .A(n36831), .B(n36830), .Z(n36833) );
  XNOR U35411 ( .A(n36828), .B(n36827), .Z(n36830) );
  XNOR U35412 ( .A(n36825), .B(n36824), .Z(n36827) );
  XNOR U35413 ( .A(n36822), .B(n36821), .Z(n36824) );
  XNOR U35414 ( .A(n36819), .B(n36818), .Z(n36821) );
  XNOR U35415 ( .A(n36816), .B(n36815), .Z(n36818) );
  XNOR U35416 ( .A(n36813), .B(n36812), .Z(n36815) );
  XNOR U35417 ( .A(n36810), .B(n36809), .Z(n36812) );
  XNOR U35418 ( .A(n36807), .B(n36806), .Z(n36809) );
  XNOR U35419 ( .A(n36804), .B(n36803), .Z(n36806) );
  XNOR U35420 ( .A(n36801), .B(n36800), .Z(n36803) );
  XNOR U35421 ( .A(n36798), .B(n36797), .Z(n36800) );
  XNOR U35422 ( .A(n36795), .B(n36794), .Z(n36797) );
  XNOR U35423 ( .A(n36792), .B(n36791), .Z(n36794) );
  XNOR U35424 ( .A(n36789), .B(n36788), .Z(n36791) );
  XNOR U35425 ( .A(n36786), .B(n36785), .Z(n36788) );
  XNOR U35426 ( .A(n36783), .B(n36782), .Z(n36785) );
  XNOR U35427 ( .A(n36780), .B(n36779), .Z(n36782) );
  XNOR U35428 ( .A(n36777), .B(n36776), .Z(n36779) );
  XNOR U35429 ( .A(n36774), .B(n36773), .Z(n36776) );
  XNOR U35430 ( .A(n36771), .B(n36770), .Z(n36773) );
  XNOR U35431 ( .A(n36768), .B(n36767), .Z(n36770) );
  XNOR U35432 ( .A(n36765), .B(n36764), .Z(n36767) );
  XNOR U35433 ( .A(n36762), .B(n36761), .Z(n36764) );
  XNOR U35434 ( .A(n36759), .B(n36758), .Z(n36761) );
  XNOR U35435 ( .A(n36756), .B(n36755), .Z(n36758) );
  XNOR U35436 ( .A(n36753), .B(n36752), .Z(n36755) );
  XNOR U35437 ( .A(n36750), .B(n36749), .Z(n36752) );
  XNOR U35438 ( .A(n36747), .B(n36746), .Z(n36749) );
  XNOR U35439 ( .A(n36744), .B(n36743), .Z(n36746) );
  XNOR U35440 ( .A(n36741), .B(n36740), .Z(n36743) );
  XNOR U35441 ( .A(n36738), .B(n36737), .Z(n36740) );
  XNOR U35442 ( .A(n36735), .B(n36734), .Z(n36737) );
  XNOR U35443 ( .A(n36732), .B(n36731), .Z(n36734) );
  XNOR U35444 ( .A(n36729), .B(n36728), .Z(n36731) );
  XNOR U35445 ( .A(n36726), .B(n36725), .Z(n36728) );
  XNOR U35446 ( .A(n36723), .B(n36722), .Z(n36725) );
  XNOR U35447 ( .A(n36720), .B(n36719), .Z(n36722) );
  XNOR U35448 ( .A(n36717), .B(n36716), .Z(n36719) );
  XNOR U35449 ( .A(n36714), .B(n36713), .Z(n36716) );
  XNOR U35450 ( .A(n36711), .B(n36710), .Z(n36713) );
  XNOR U35451 ( .A(n36708), .B(n36707), .Z(n36710) );
  XNOR U35452 ( .A(n36705), .B(n36704), .Z(n36707) );
  XNOR U35453 ( .A(n36702), .B(n36701), .Z(n36704) );
  XNOR U35454 ( .A(n36699), .B(n36698), .Z(n36701) );
  XNOR U35455 ( .A(n36696), .B(n36695), .Z(n36698) );
  XNOR U35456 ( .A(n36693), .B(n36692), .Z(n36695) );
  XNOR U35457 ( .A(n36690), .B(n36689), .Z(n36692) );
  XNOR U35458 ( .A(n36687), .B(n36686), .Z(n36689) );
  XNOR U35459 ( .A(n36684), .B(n36683), .Z(n36686) );
  XNOR U35460 ( .A(n36681), .B(n36680), .Z(n36683) );
  XNOR U35461 ( .A(n36678), .B(n36677), .Z(n36680) );
  XNOR U35462 ( .A(n36675), .B(n36674), .Z(n36677) );
  XNOR U35463 ( .A(n36672), .B(n36671), .Z(n36674) );
  XNOR U35464 ( .A(n36669), .B(n36668), .Z(n36671) );
  XNOR U35465 ( .A(n36666), .B(n36665), .Z(n36668) );
  XNOR U35466 ( .A(n36663), .B(n36662), .Z(n36665) );
  XNOR U35467 ( .A(n36660), .B(n36659), .Z(n36662) );
  XNOR U35468 ( .A(n36657), .B(n36656), .Z(n36659) );
  XNOR U35469 ( .A(n36654), .B(n36653), .Z(n36656) );
  XNOR U35470 ( .A(n36651), .B(n36650), .Z(n36653) );
  XNOR U35471 ( .A(n36648), .B(n36647), .Z(n36650) );
  XNOR U35472 ( .A(n36645), .B(n36644), .Z(n36647) );
  XNOR U35473 ( .A(n36642), .B(n36641), .Z(n36644) );
  XNOR U35474 ( .A(n36639), .B(n36638), .Z(n36641) );
  XNOR U35475 ( .A(n36636), .B(n36635), .Z(n36638) );
  XNOR U35476 ( .A(n36633), .B(n36632), .Z(n36635) );
  XNOR U35477 ( .A(n36630), .B(n36629), .Z(n36632) );
  XNOR U35478 ( .A(n36627), .B(n36626), .Z(n36629) );
  XNOR U35479 ( .A(n36624), .B(n36623), .Z(n36626) );
  XNOR U35480 ( .A(n36621), .B(n36620), .Z(n36623) );
  XNOR U35481 ( .A(n36618), .B(n36617), .Z(n36620) );
  XNOR U35482 ( .A(n36615), .B(n36614), .Z(n36617) );
  XNOR U35483 ( .A(n36612), .B(n36611), .Z(n36614) );
  XNOR U35484 ( .A(n36609), .B(n36608), .Z(n36611) );
  XNOR U35485 ( .A(n36606), .B(n36605), .Z(n36608) );
  XNOR U35486 ( .A(n36603), .B(n36602), .Z(n36605) );
  XNOR U35487 ( .A(n36600), .B(n36599), .Z(n36602) );
  XNOR U35488 ( .A(n36597), .B(n36596), .Z(n36599) );
  XNOR U35489 ( .A(n36594), .B(n36593), .Z(n36596) );
  XNOR U35490 ( .A(n36591), .B(n36590), .Z(n36593) );
  XNOR U35491 ( .A(n36588), .B(n36587), .Z(n36590) );
  XNOR U35492 ( .A(n36585), .B(n36584), .Z(n36587) );
  XNOR U35493 ( .A(n36582), .B(n36581), .Z(n36584) );
  XNOR U35494 ( .A(n36579), .B(n36578), .Z(n36581) );
  XNOR U35495 ( .A(n36576), .B(n36575), .Z(n36578) );
  XNOR U35496 ( .A(n36573), .B(n36572), .Z(n36575) );
  XNOR U35497 ( .A(n36570), .B(n36569), .Z(n36572) );
  XNOR U35498 ( .A(n36567), .B(n36566), .Z(n36569) );
  XNOR U35499 ( .A(n36564), .B(n36563), .Z(n36566) );
  XNOR U35500 ( .A(n36561), .B(n36560), .Z(n36563) );
  XNOR U35501 ( .A(n36558), .B(n36557), .Z(n36560) );
  XNOR U35502 ( .A(n36555), .B(n36554), .Z(n36557) );
  XNOR U35503 ( .A(n36552), .B(n36551), .Z(n36554) );
  XNOR U35504 ( .A(n36549), .B(n36548), .Z(n36551) );
  XNOR U35505 ( .A(n36546), .B(n36545), .Z(n36548) );
  XNOR U35506 ( .A(n36543), .B(n36542), .Z(n36545) );
  XNOR U35507 ( .A(n36540), .B(n36539), .Z(n36542) );
  XNOR U35508 ( .A(n36537), .B(n36536), .Z(n36539) );
  XNOR U35509 ( .A(n36534), .B(n36533), .Z(n36536) );
  XNOR U35510 ( .A(n36531), .B(n36530), .Z(n36533) );
  XNOR U35511 ( .A(n36528), .B(n36527), .Z(n36530) );
  XNOR U35512 ( .A(n36525), .B(n36524), .Z(n36527) );
  XNOR U35513 ( .A(n36522), .B(n36521), .Z(n36524) );
  XNOR U35514 ( .A(n36519), .B(n36518), .Z(n36521) );
  XNOR U35515 ( .A(n36516), .B(n36515), .Z(n36518) );
  XNOR U35516 ( .A(n36513), .B(n36512), .Z(n36515) );
  XNOR U35517 ( .A(n36510), .B(n36509), .Z(n36512) );
  XNOR U35518 ( .A(n36507), .B(n36506), .Z(n36509) );
  XNOR U35519 ( .A(n36504), .B(n36503), .Z(n36506) );
  XNOR U35520 ( .A(n36501), .B(n36500), .Z(n36503) );
  XNOR U35521 ( .A(n36498), .B(n36497), .Z(n36500) );
  XNOR U35522 ( .A(n36495), .B(n36494), .Z(n36497) );
  XNOR U35523 ( .A(n36492), .B(n36491), .Z(n36494) );
  XNOR U35524 ( .A(n36489), .B(n36488), .Z(n36491) );
  XNOR U35525 ( .A(n36486), .B(n36485), .Z(n36488) );
  XNOR U35526 ( .A(n36483), .B(n36482), .Z(n36485) );
  XNOR U35527 ( .A(n36480), .B(n36479), .Z(n36482) );
  XNOR U35528 ( .A(n36477), .B(n36476), .Z(n36479) );
  XNOR U35529 ( .A(n36474), .B(n36473), .Z(n36476) );
  XNOR U35530 ( .A(n36471), .B(n36470), .Z(n36473) );
  XNOR U35531 ( .A(n36468), .B(n36467), .Z(n36470) );
  XNOR U35532 ( .A(n36465), .B(n36464), .Z(n36467) );
  XNOR U35533 ( .A(n36462), .B(n36461), .Z(n36464) );
  XNOR U35534 ( .A(n36459), .B(n36458), .Z(n36461) );
  XNOR U35535 ( .A(n36456), .B(n36455), .Z(n36458) );
  XNOR U35536 ( .A(n36453), .B(n36452), .Z(n36455) );
  XNOR U35537 ( .A(n36450), .B(n36449), .Z(n36452) );
  XNOR U35538 ( .A(n36447), .B(n36446), .Z(n36449) );
  XNOR U35539 ( .A(n36444), .B(n36443), .Z(n36446) );
  XNOR U35540 ( .A(n36441), .B(n36440), .Z(n36443) );
  XNOR U35541 ( .A(n36438), .B(n36437), .Z(n36440) );
  XNOR U35542 ( .A(n36435), .B(n36434), .Z(n36437) );
  XNOR U35543 ( .A(n36432), .B(n36431), .Z(n36434) );
  XNOR U35544 ( .A(n36429), .B(n36428), .Z(n36431) );
  XNOR U35545 ( .A(n36426), .B(n36425), .Z(n36428) );
  XNOR U35546 ( .A(n36423), .B(n36422), .Z(n36425) );
  XNOR U35547 ( .A(n36420), .B(n36419), .Z(n36422) );
  XNOR U35548 ( .A(n36417), .B(n36416), .Z(n36419) );
  XNOR U35549 ( .A(n36414), .B(n36413), .Z(n36416) );
  XNOR U35550 ( .A(n36411), .B(n36410), .Z(n36413) );
  XNOR U35551 ( .A(n36408), .B(n36407), .Z(n36410) );
  XNOR U35552 ( .A(n36405), .B(n36404), .Z(n36407) );
  XNOR U35553 ( .A(n36402), .B(n36401), .Z(n36404) );
  XNOR U35554 ( .A(n36399), .B(n36398), .Z(n36401) );
  XNOR U35555 ( .A(n36396), .B(n36395), .Z(n36398) );
  XNOR U35556 ( .A(n36393), .B(n36392), .Z(n36395) );
  XNOR U35557 ( .A(n36390), .B(n36389), .Z(n36392) );
  XNOR U35558 ( .A(n36387), .B(n36386), .Z(n36389) );
  XNOR U35559 ( .A(n36384), .B(n36383), .Z(n36386) );
  XNOR U35560 ( .A(n36381), .B(n36380), .Z(n36383) );
  XNOR U35561 ( .A(n36378), .B(n36377), .Z(n36380) );
  XNOR U35562 ( .A(n36375), .B(n36374), .Z(n36377) );
  XNOR U35563 ( .A(n36372), .B(n36371), .Z(n36374) );
  XNOR U35564 ( .A(n36369), .B(n36368), .Z(n36371) );
  XNOR U35565 ( .A(n36366), .B(n36365), .Z(n36368) );
  XNOR U35566 ( .A(n36363), .B(n36362), .Z(n36365) );
  XNOR U35567 ( .A(n36360), .B(n36359), .Z(n36362) );
  XNOR U35568 ( .A(n36357), .B(n36356), .Z(n36359) );
  XNOR U35569 ( .A(n36354), .B(n36353), .Z(n36356) );
  XNOR U35570 ( .A(n36351), .B(n36350), .Z(n36353) );
  XNOR U35571 ( .A(n36348), .B(n36347), .Z(n36350) );
  XNOR U35572 ( .A(n36345), .B(n36344), .Z(n36347) );
  XNOR U35573 ( .A(n36342), .B(n36341), .Z(n36344) );
  XNOR U35574 ( .A(n36339), .B(n36338), .Z(n36341) );
  XNOR U35575 ( .A(n36336), .B(n36335), .Z(n36338) );
  XNOR U35576 ( .A(n36333), .B(n36332), .Z(n36335) );
  XNOR U35577 ( .A(n36330), .B(n36329), .Z(n36332) );
  XNOR U35578 ( .A(n36327), .B(n36326), .Z(n36329) );
  XNOR U35579 ( .A(n36324), .B(n36323), .Z(n36326) );
  XNOR U35580 ( .A(n36321), .B(n36320), .Z(n36323) );
  XNOR U35581 ( .A(n36318), .B(n36317), .Z(n36320) );
  XNOR U35582 ( .A(n36315), .B(n36314), .Z(n36317) );
  XNOR U35583 ( .A(n36312), .B(n36311), .Z(n36314) );
  XNOR U35584 ( .A(n36309), .B(n36308), .Z(n36311) );
  XNOR U35585 ( .A(n36306), .B(n36305), .Z(n36308) );
  XNOR U35586 ( .A(n36303), .B(n36302), .Z(n36305) );
  XNOR U35587 ( .A(n36300), .B(n36299), .Z(n36302) );
  XNOR U35588 ( .A(n36297), .B(n36296), .Z(n36299) );
  XNOR U35589 ( .A(n36294), .B(n36293), .Z(n36296) );
  XNOR U35590 ( .A(n36291), .B(n36290), .Z(n36293) );
  XNOR U35591 ( .A(n36288), .B(n36287), .Z(n36290) );
  XNOR U35592 ( .A(n36285), .B(n36284), .Z(n36287) );
  XNOR U35593 ( .A(n36282), .B(n36281), .Z(n36284) );
  XNOR U35594 ( .A(n36279), .B(n36278), .Z(n36281) );
  XNOR U35595 ( .A(n36276), .B(n36275), .Z(n36278) );
  XNOR U35596 ( .A(n36273), .B(n36272), .Z(n36275) );
  XNOR U35597 ( .A(n36270), .B(n36269), .Z(n36272) );
  XNOR U35598 ( .A(n36267), .B(n36266), .Z(n36269) );
  XNOR U35599 ( .A(n36264), .B(n36263), .Z(n36266) );
  XNOR U35600 ( .A(n36261), .B(n36260), .Z(n36263) );
  XNOR U35601 ( .A(n36258), .B(n36257), .Z(n36260) );
  XNOR U35602 ( .A(n36255), .B(n36254), .Z(n36257) );
  XNOR U35603 ( .A(n36252), .B(n36251), .Z(n36254) );
  XNOR U35604 ( .A(n36249), .B(n36248), .Z(n36251) );
  XNOR U35605 ( .A(n36246), .B(n36245), .Z(n36248) );
  XNOR U35606 ( .A(n36243), .B(n36242), .Z(n36245) );
  XNOR U35607 ( .A(n36240), .B(n36239), .Z(n36242) );
  XNOR U35608 ( .A(n36237), .B(n36236), .Z(n36239) );
  XNOR U35609 ( .A(n36234), .B(n36233), .Z(n36236) );
  XNOR U35610 ( .A(n36231), .B(n36230), .Z(n36233) );
  XNOR U35611 ( .A(n36228), .B(n36227), .Z(n36230) );
  XNOR U35612 ( .A(n36225), .B(n36224), .Z(n36227) );
  XNOR U35613 ( .A(n36222), .B(n36221), .Z(n36224) );
  XNOR U35614 ( .A(n36219), .B(n36218), .Z(n36221) );
  XNOR U35615 ( .A(n36216), .B(n36215), .Z(n36218) );
  XNOR U35616 ( .A(n36213), .B(n36212), .Z(n36215) );
  XNOR U35617 ( .A(n36210), .B(n36209), .Z(n36212) );
  XNOR U35618 ( .A(n36207), .B(n36206), .Z(n36209) );
  XNOR U35619 ( .A(n36204), .B(n36203), .Z(n36206) );
  XNOR U35620 ( .A(n36201), .B(n36200), .Z(n36203) );
  XNOR U35621 ( .A(n36198), .B(n36197), .Z(n36200) );
  XNOR U35622 ( .A(n36195), .B(n36194), .Z(n36197) );
  XNOR U35623 ( .A(n36192), .B(n36191), .Z(n36194) );
  XNOR U35624 ( .A(n36189), .B(n36188), .Z(n36191) );
  XNOR U35625 ( .A(n36186), .B(n36185), .Z(n36188) );
  XNOR U35626 ( .A(n36183), .B(n36182), .Z(n36185) );
  XNOR U35627 ( .A(n36180), .B(n36179), .Z(n36182) );
  XNOR U35628 ( .A(n36177), .B(n36176), .Z(n36179) );
  XNOR U35629 ( .A(n36174), .B(n36173), .Z(n36176) );
  XNOR U35630 ( .A(n36171), .B(n36170), .Z(n36173) );
  XNOR U35631 ( .A(n36168), .B(n36167), .Z(n36170) );
  XNOR U35632 ( .A(n36165), .B(n36164), .Z(n36167) );
  XNOR U35633 ( .A(n36162), .B(n36161), .Z(n36164) );
  XNOR U35634 ( .A(n36159), .B(n36158), .Z(n36161) );
  XNOR U35635 ( .A(n36156), .B(n36155), .Z(n36158) );
  XNOR U35636 ( .A(n36153), .B(n36152), .Z(n36155) );
  XNOR U35637 ( .A(n36150), .B(n36149), .Z(n36152) );
  XNOR U35638 ( .A(n36147), .B(n36146), .Z(n36149) );
  XNOR U35639 ( .A(n36144), .B(n36143), .Z(n36146) );
  XNOR U35640 ( .A(n36141), .B(n36140), .Z(n36143) );
  XNOR U35641 ( .A(n36138), .B(n36137), .Z(n36140) );
  XNOR U35642 ( .A(n36135), .B(n36134), .Z(n36137) );
  XNOR U35643 ( .A(n36132), .B(n36131), .Z(n36134) );
  XNOR U35644 ( .A(n36129), .B(n36128), .Z(n36131) );
  XNOR U35645 ( .A(n36126), .B(n36125), .Z(n36128) );
  XNOR U35646 ( .A(n36123), .B(n36122), .Z(n36125) );
  XNOR U35647 ( .A(n36120), .B(n36119), .Z(n36122) );
  XNOR U35648 ( .A(n36117), .B(n36116), .Z(n36119) );
  XNOR U35649 ( .A(n36114), .B(n36113), .Z(n36116) );
  XNOR U35650 ( .A(n36111), .B(n36110), .Z(n36113) );
  XNOR U35651 ( .A(n36108), .B(n36107), .Z(n36110) );
  XNOR U35652 ( .A(n36105), .B(n36104), .Z(n36107) );
  XNOR U35653 ( .A(n36102), .B(n36101), .Z(n36104) );
  XNOR U35654 ( .A(n36099), .B(n36098), .Z(n36101) );
  XNOR U35655 ( .A(n36096), .B(n36095), .Z(n36098) );
  XNOR U35656 ( .A(n36093), .B(n36092), .Z(n36095) );
  XNOR U35657 ( .A(n36090), .B(n36089), .Z(n36092) );
  XNOR U35658 ( .A(n36087), .B(n36086), .Z(n36089) );
  XNOR U35659 ( .A(n36084), .B(n36083), .Z(n36086) );
  XNOR U35660 ( .A(n36081), .B(n36080), .Z(n36083) );
  XNOR U35661 ( .A(n36078), .B(n36077), .Z(n36080) );
  XNOR U35662 ( .A(n36075), .B(n36074), .Z(n36077) );
  XNOR U35663 ( .A(n36072), .B(n36071), .Z(n36074) );
  XNOR U35664 ( .A(n36069), .B(n36068), .Z(n36071) );
  XNOR U35665 ( .A(n36066), .B(n36065), .Z(n36068) );
  XNOR U35666 ( .A(n36063), .B(n36062), .Z(n36065) );
  XNOR U35667 ( .A(n36060), .B(n36059), .Z(n36062) );
  XNOR U35668 ( .A(n36057), .B(n36056), .Z(n36059) );
  XNOR U35669 ( .A(n36054), .B(n36053), .Z(n36056) );
  XNOR U35670 ( .A(n36051), .B(n36050), .Z(n36053) );
  XNOR U35671 ( .A(n36048), .B(n36047), .Z(n36050) );
  XNOR U35672 ( .A(n36045), .B(n36044), .Z(n36047) );
  XNOR U35673 ( .A(n36042), .B(n36041), .Z(n36044) );
  XNOR U35674 ( .A(n36039), .B(n36038), .Z(n36041) );
  XNOR U35675 ( .A(n36036), .B(n36035), .Z(n36038) );
  XNOR U35676 ( .A(n36033), .B(n36032), .Z(n36035) );
  XNOR U35677 ( .A(n36030), .B(n36029), .Z(n36032) );
  XNOR U35678 ( .A(n36027), .B(n36026), .Z(n36029) );
  XNOR U35679 ( .A(n36024), .B(n36023), .Z(n36026) );
  XNOR U35680 ( .A(n36021), .B(n36020), .Z(n36023) );
  XNOR U35681 ( .A(n36018), .B(n36017), .Z(n36020) );
  XNOR U35682 ( .A(n36015), .B(n36014), .Z(n36017) );
  XNOR U35683 ( .A(n36012), .B(n36011), .Z(n36014) );
  XNOR U35684 ( .A(n36009), .B(n36008), .Z(n36011) );
  XNOR U35685 ( .A(n36006), .B(n36005), .Z(n36008) );
  XNOR U35686 ( .A(n36003), .B(n36002), .Z(n36005) );
  XNOR U35687 ( .A(n36000), .B(n35999), .Z(n36002) );
  XNOR U35688 ( .A(n35997), .B(n35996), .Z(n35999) );
  XNOR U35689 ( .A(n35994), .B(n35993), .Z(n35996) );
  XNOR U35690 ( .A(n35991), .B(n35990), .Z(n35993) );
  XNOR U35691 ( .A(n35988), .B(n35987), .Z(n35990) );
  XNOR U35692 ( .A(n35985), .B(n35984), .Z(n35987) );
  XNOR U35693 ( .A(n35982), .B(n35981), .Z(n35984) );
  XNOR U35694 ( .A(n35979), .B(n35978), .Z(n35981) );
  XNOR U35695 ( .A(n35976), .B(n35975), .Z(n35978) );
  XNOR U35696 ( .A(n35973), .B(n35972), .Z(n35975) );
  XNOR U35697 ( .A(n35970), .B(n35969), .Z(n35972) );
  XNOR U35698 ( .A(n35967), .B(n35966), .Z(n35969) );
  XNOR U35699 ( .A(n35964), .B(n35963), .Z(n35966) );
  XNOR U35700 ( .A(n35961), .B(n35960), .Z(n35963) );
  XNOR U35701 ( .A(n35958), .B(n35957), .Z(n35960) );
  XNOR U35702 ( .A(n35955), .B(n35954), .Z(n35957) );
  XNOR U35703 ( .A(n35952), .B(n35951), .Z(n35954) );
  XNOR U35704 ( .A(n35949), .B(n35948), .Z(n35951) );
  XNOR U35705 ( .A(n35946), .B(n35945), .Z(n35948) );
  XNOR U35706 ( .A(n35943), .B(n35942), .Z(n35945) );
  XNOR U35707 ( .A(n35940), .B(n35939), .Z(n35942) );
  XNOR U35708 ( .A(n35937), .B(n35936), .Z(n35939) );
  XNOR U35709 ( .A(n35934), .B(n35933), .Z(n35936) );
  XNOR U35710 ( .A(n35931), .B(n35930), .Z(n35933) );
  XNOR U35711 ( .A(n35928), .B(n35927), .Z(n35930) );
  XNOR U35712 ( .A(n35925), .B(n35924), .Z(n35927) );
  XNOR U35713 ( .A(n35922), .B(n35921), .Z(n35924) );
  XNOR U35714 ( .A(n35919), .B(n35918), .Z(n35921) );
  XNOR U35715 ( .A(n35916), .B(n35915), .Z(n35918) );
  XNOR U35716 ( .A(n35913), .B(n35912), .Z(n35915) );
  XNOR U35717 ( .A(n35910), .B(n35909), .Z(n35912) );
  XNOR U35718 ( .A(n35907), .B(n35906), .Z(n35909) );
  XNOR U35719 ( .A(n35904), .B(n35903), .Z(n35906) );
  XNOR U35720 ( .A(n35901), .B(n35900), .Z(n35903) );
  XNOR U35721 ( .A(n35898), .B(n35897), .Z(n35900) );
  XNOR U35722 ( .A(n35895), .B(n35894), .Z(n35897) );
  XNOR U35723 ( .A(n35892), .B(n35891), .Z(n35894) );
  XNOR U35724 ( .A(n35889), .B(n35888), .Z(n35891) );
  XNOR U35725 ( .A(n35886), .B(n35885), .Z(n35888) );
  XNOR U35726 ( .A(n35883), .B(n35882), .Z(n35885) );
  XNOR U35727 ( .A(n35880), .B(n35879), .Z(n35882) );
  XNOR U35728 ( .A(n35877), .B(n35876), .Z(n35879) );
  XNOR U35729 ( .A(n35874), .B(n35873), .Z(n35876) );
  XNOR U35730 ( .A(n35871), .B(n35870), .Z(n35873) );
  XNOR U35731 ( .A(n35868), .B(n35867), .Z(n35870) );
  XNOR U35732 ( .A(n35865), .B(n35864), .Z(n35867) );
  XNOR U35733 ( .A(n35862), .B(n35861), .Z(n35864) );
  XNOR U35734 ( .A(n35859), .B(n35858), .Z(n35861) );
  XNOR U35735 ( .A(n35856), .B(n35855), .Z(n35858) );
  XNOR U35736 ( .A(n35853), .B(n35852), .Z(n35855) );
  XNOR U35737 ( .A(n35850), .B(n35849), .Z(n35852) );
  XNOR U35738 ( .A(n35847), .B(n35846), .Z(n35849) );
  XNOR U35739 ( .A(n35844), .B(n35843), .Z(n35846) );
  XNOR U35740 ( .A(n35841), .B(n35840), .Z(n35843) );
  XNOR U35741 ( .A(n35838), .B(n35837), .Z(n35840) );
  XNOR U35742 ( .A(n35835), .B(n35834), .Z(n35837) );
  XNOR U35743 ( .A(n35832), .B(n35831), .Z(n35834) );
  XNOR U35744 ( .A(n35829), .B(n35828), .Z(n35831) );
  XNOR U35745 ( .A(n35826), .B(n35825), .Z(n35828) );
  XNOR U35746 ( .A(n35823), .B(n35822), .Z(n35825) );
  XNOR U35747 ( .A(n35820), .B(n35819), .Z(n35822) );
  XNOR U35748 ( .A(n35817), .B(n35816), .Z(n35819) );
  XNOR U35749 ( .A(n35814), .B(n35813), .Z(n35816) );
  XNOR U35750 ( .A(n35811), .B(n35810), .Z(n35813) );
  XNOR U35751 ( .A(n35808), .B(n35807), .Z(n35810) );
  XNOR U35752 ( .A(n35805), .B(n35804), .Z(n35807) );
  XNOR U35753 ( .A(n35802), .B(n35801), .Z(n35804) );
  XNOR U35754 ( .A(n35799), .B(n35798), .Z(n35801) );
  XNOR U35755 ( .A(n35796), .B(n35795), .Z(n35798) );
  XOR U35756 ( .A(n35793), .B(n35792), .Z(n35795) );
  XOR U35757 ( .A(n35790), .B(n35789), .Z(n35792) );
  XOR U35758 ( .A(n35786), .B(n35787), .Z(n35789) );
  AND U35759 ( .A(n38388), .B(n38389), .Z(n35787) );
  XOR U35760 ( .A(n35783), .B(n35784), .Z(n35786) );
  AND U35761 ( .A(n38390), .B(n38391), .Z(n35784) );
  XOR U35762 ( .A(n35780), .B(n35781), .Z(n35783) );
  AND U35763 ( .A(n38392), .B(n38393), .Z(n35781) );
  XNOR U35764 ( .A(n35535), .B(n35778), .Z(n35780) );
  AND U35765 ( .A(n38394), .B(n38395), .Z(n35778) );
  XOR U35766 ( .A(n35537), .B(n35536), .Z(n35535) );
  AND U35767 ( .A(n38396), .B(n38397), .Z(n35536) );
  XOR U35768 ( .A(n35539), .B(n35538), .Z(n35537) );
  AND U35769 ( .A(n38398), .B(n38399), .Z(n35538) );
  XOR U35770 ( .A(n35541), .B(n35540), .Z(n35539) );
  AND U35771 ( .A(n38400), .B(n38401), .Z(n35540) );
  XOR U35772 ( .A(n35543), .B(n35542), .Z(n35541) );
  AND U35773 ( .A(n38402), .B(n38403), .Z(n35542) );
  XOR U35774 ( .A(n35545), .B(n35544), .Z(n35543) );
  AND U35775 ( .A(n38404), .B(n38405), .Z(n35544) );
  XOR U35776 ( .A(n35547), .B(n35546), .Z(n35545) );
  AND U35777 ( .A(n38406), .B(n38407), .Z(n35546) );
  XOR U35778 ( .A(n35549), .B(n35548), .Z(n35547) );
  AND U35779 ( .A(n38408), .B(n38409), .Z(n35548) );
  XOR U35780 ( .A(n35551), .B(n35550), .Z(n35549) );
  AND U35781 ( .A(n38410), .B(n38411), .Z(n35550) );
  XOR U35782 ( .A(n35553), .B(n35552), .Z(n35551) );
  AND U35783 ( .A(n38412), .B(n38413), .Z(n35552) );
  XOR U35784 ( .A(n35555), .B(n35554), .Z(n35553) );
  AND U35785 ( .A(n38414), .B(n38415), .Z(n35554) );
  XOR U35786 ( .A(n35557), .B(n35556), .Z(n35555) );
  AND U35787 ( .A(n38416), .B(n38417), .Z(n35556) );
  XOR U35788 ( .A(n35559), .B(n35558), .Z(n35557) );
  AND U35789 ( .A(n38418), .B(n38419), .Z(n35558) );
  XOR U35790 ( .A(n35561), .B(n35560), .Z(n35559) );
  AND U35791 ( .A(n38420), .B(n38421), .Z(n35560) );
  XOR U35792 ( .A(n35563), .B(n35562), .Z(n35561) );
  AND U35793 ( .A(n38422), .B(n38423), .Z(n35562) );
  XOR U35794 ( .A(n35565), .B(n35564), .Z(n35563) );
  AND U35795 ( .A(n38424), .B(n38425), .Z(n35564) );
  XOR U35796 ( .A(n35567), .B(n35566), .Z(n35565) );
  AND U35797 ( .A(n38426), .B(n38427), .Z(n35566) );
  XOR U35798 ( .A(n35569), .B(n35568), .Z(n35567) );
  AND U35799 ( .A(n38428), .B(n38429), .Z(n35568) );
  XOR U35800 ( .A(n35571), .B(n35570), .Z(n35569) );
  AND U35801 ( .A(n38430), .B(n38431), .Z(n35570) );
  XOR U35802 ( .A(n35573), .B(n35572), .Z(n35571) );
  AND U35803 ( .A(n38432), .B(n38433), .Z(n35572) );
  XOR U35804 ( .A(n35575), .B(n35574), .Z(n35573) );
  AND U35805 ( .A(n38434), .B(n38435), .Z(n35574) );
  XOR U35806 ( .A(n35577), .B(n35576), .Z(n35575) );
  AND U35807 ( .A(n38436), .B(n38437), .Z(n35576) );
  XOR U35808 ( .A(n35579), .B(n35578), .Z(n35577) );
  AND U35809 ( .A(n38438), .B(n38439), .Z(n35578) );
  XOR U35810 ( .A(n35581), .B(n35580), .Z(n35579) );
  AND U35811 ( .A(n38440), .B(n38441), .Z(n35580) );
  XOR U35812 ( .A(n35583), .B(n35582), .Z(n35581) );
  AND U35813 ( .A(n38442), .B(n38443), .Z(n35582) );
  XOR U35814 ( .A(n35585), .B(n35584), .Z(n35583) );
  AND U35815 ( .A(n38444), .B(n38445), .Z(n35584) );
  XOR U35816 ( .A(n35587), .B(n35586), .Z(n35585) );
  AND U35817 ( .A(n38446), .B(n38447), .Z(n35586) );
  XOR U35818 ( .A(n35589), .B(n35588), .Z(n35587) );
  AND U35819 ( .A(n38448), .B(n38449), .Z(n35588) );
  XOR U35820 ( .A(n35591), .B(n35590), .Z(n35589) );
  AND U35821 ( .A(n38450), .B(n38451), .Z(n35590) );
  XOR U35822 ( .A(n35593), .B(n35592), .Z(n35591) );
  AND U35823 ( .A(n38452), .B(n38453), .Z(n35592) );
  XOR U35824 ( .A(n35595), .B(n35594), .Z(n35593) );
  AND U35825 ( .A(n38454), .B(n38455), .Z(n35594) );
  XOR U35826 ( .A(n35597), .B(n35596), .Z(n35595) );
  AND U35827 ( .A(n38456), .B(n38457), .Z(n35596) );
  XOR U35828 ( .A(n35599), .B(n35598), .Z(n35597) );
  AND U35829 ( .A(n38458), .B(n38459), .Z(n35598) );
  XOR U35830 ( .A(n35601), .B(n35600), .Z(n35599) );
  AND U35831 ( .A(n38460), .B(n38461), .Z(n35600) );
  XOR U35832 ( .A(n35603), .B(n35602), .Z(n35601) );
  AND U35833 ( .A(n38462), .B(n38463), .Z(n35602) );
  XOR U35834 ( .A(n35605), .B(n35604), .Z(n35603) );
  AND U35835 ( .A(n38464), .B(n38465), .Z(n35604) );
  XOR U35836 ( .A(n35607), .B(n35606), .Z(n35605) );
  AND U35837 ( .A(n38466), .B(n38467), .Z(n35606) );
  XOR U35838 ( .A(n35609), .B(n35608), .Z(n35607) );
  AND U35839 ( .A(n38468), .B(n38469), .Z(n35608) );
  XOR U35840 ( .A(n35611), .B(n35610), .Z(n35609) );
  AND U35841 ( .A(n38470), .B(n38471), .Z(n35610) );
  XOR U35842 ( .A(n35613), .B(n35612), .Z(n35611) );
  AND U35843 ( .A(n38472), .B(n38473), .Z(n35612) );
  XOR U35844 ( .A(n35615), .B(n35614), .Z(n35613) );
  AND U35845 ( .A(n38474), .B(n38475), .Z(n35614) );
  XOR U35846 ( .A(n35617), .B(n35616), .Z(n35615) );
  AND U35847 ( .A(n38476), .B(n38477), .Z(n35616) );
  XOR U35848 ( .A(n35619), .B(n35618), .Z(n35617) );
  AND U35849 ( .A(n38478), .B(n38479), .Z(n35618) );
  XOR U35850 ( .A(n35621), .B(n35620), .Z(n35619) );
  AND U35851 ( .A(n38480), .B(n38481), .Z(n35620) );
  XOR U35852 ( .A(n35623), .B(n35622), .Z(n35621) );
  AND U35853 ( .A(n38482), .B(n38483), .Z(n35622) );
  XOR U35854 ( .A(n35625), .B(n35624), .Z(n35623) );
  AND U35855 ( .A(n38484), .B(n38485), .Z(n35624) );
  XOR U35856 ( .A(n35627), .B(n35626), .Z(n35625) );
  AND U35857 ( .A(n38486), .B(n38487), .Z(n35626) );
  XOR U35858 ( .A(n35629), .B(n35628), .Z(n35627) );
  AND U35859 ( .A(n38488), .B(n38489), .Z(n35628) );
  XOR U35860 ( .A(n35631), .B(n35630), .Z(n35629) );
  AND U35861 ( .A(n38490), .B(n38491), .Z(n35630) );
  XOR U35862 ( .A(n35633), .B(n35632), .Z(n35631) );
  AND U35863 ( .A(n38492), .B(n38493), .Z(n35632) );
  XOR U35864 ( .A(n35635), .B(n35634), .Z(n35633) );
  AND U35865 ( .A(n38494), .B(n38495), .Z(n35634) );
  XOR U35866 ( .A(n35637), .B(n35636), .Z(n35635) );
  AND U35867 ( .A(n38496), .B(n38497), .Z(n35636) );
  XOR U35868 ( .A(n35639), .B(n35638), .Z(n35637) );
  AND U35869 ( .A(n38498), .B(n38499), .Z(n35638) );
  XOR U35870 ( .A(n35641), .B(n35640), .Z(n35639) );
  AND U35871 ( .A(n38500), .B(n38501), .Z(n35640) );
  XOR U35872 ( .A(n35643), .B(n35642), .Z(n35641) );
  AND U35873 ( .A(n38502), .B(n38503), .Z(n35642) );
  XOR U35874 ( .A(n35645), .B(n35644), .Z(n35643) );
  AND U35875 ( .A(n38504), .B(n38505), .Z(n35644) );
  XOR U35876 ( .A(n35647), .B(n35646), .Z(n35645) );
  AND U35877 ( .A(n38506), .B(n38507), .Z(n35646) );
  XOR U35878 ( .A(n35649), .B(n35648), .Z(n35647) );
  AND U35879 ( .A(n38508), .B(n38509), .Z(n35648) );
  XOR U35880 ( .A(n35651), .B(n35650), .Z(n35649) );
  AND U35881 ( .A(n38510), .B(n38511), .Z(n35650) );
  XOR U35882 ( .A(n35653), .B(n35652), .Z(n35651) );
  AND U35883 ( .A(n38512), .B(n38513), .Z(n35652) );
  XOR U35884 ( .A(n35655), .B(n35654), .Z(n35653) );
  AND U35885 ( .A(n38514), .B(n38515), .Z(n35654) );
  XOR U35886 ( .A(n35657), .B(n35656), .Z(n35655) );
  AND U35887 ( .A(n38516), .B(n38517), .Z(n35656) );
  XOR U35888 ( .A(n35659), .B(n35658), .Z(n35657) );
  AND U35889 ( .A(n38518), .B(n38519), .Z(n35658) );
  XOR U35890 ( .A(n35661), .B(n35660), .Z(n35659) );
  AND U35891 ( .A(n38520), .B(n38521), .Z(n35660) );
  XOR U35892 ( .A(n35663), .B(n35662), .Z(n35661) );
  AND U35893 ( .A(n38522), .B(n38523), .Z(n35662) );
  XOR U35894 ( .A(n35665), .B(n35664), .Z(n35663) );
  AND U35895 ( .A(n38524), .B(n38525), .Z(n35664) );
  XOR U35896 ( .A(n35667), .B(n35666), .Z(n35665) );
  AND U35897 ( .A(n38526), .B(n38527), .Z(n35666) );
  XOR U35898 ( .A(n35669), .B(n35668), .Z(n35667) );
  AND U35899 ( .A(n38528), .B(n38529), .Z(n35668) );
  XOR U35900 ( .A(n35671), .B(n35670), .Z(n35669) );
  AND U35901 ( .A(n38530), .B(n38531), .Z(n35670) );
  XOR U35902 ( .A(n35680), .B(n35672), .Z(n35671) );
  AND U35903 ( .A(n38532), .B(n38533), .Z(n35672) );
  XOR U35904 ( .A(n35675), .B(n35681), .Z(n35680) );
  AND U35905 ( .A(n38534), .B(n38535), .Z(n35681) );
  XOR U35906 ( .A(n35677), .B(n35676), .Z(n35675) );
  AND U35907 ( .A(n38536), .B(n38537), .Z(n35676) );
  XOR U35908 ( .A(n35701), .B(n35678), .Z(n35677) );
  AND U35909 ( .A(n38538), .B(n38539), .Z(n35678) );
  XOR U35910 ( .A(n35696), .B(n35702), .Z(n35701) );
  AND U35911 ( .A(n38540), .B(n38541), .Z(n35702) );
  XOR U35912 ( .A(n35698), .B(n35697), .Z(n35696) );
  AND U35913 ( .A(n38542), .B(n38543), .Z(n35697) );
  XOR U35914 ( .A(n35686), .B(n35699), .Z(n35698) );
  AND U35915 ( .A(n38544), .B(n38545), .Z(n35699) );
  XOR U35916 ( .A(n35688), .B(n35687), .Z(n35686) );
  AND U35917 ( .A(n38546), .B(n38547), .Z(n35687) );
  XOR U35918 ( .A(n35690), .B(n35689), .Z(n35688) );
  AND U35919 ( .A(n38548), .B(n38549), .Z(n35689) );
  XOR U35920 ( .A(n35692), .B(n35691), .Z(n35690) );
  AND U35921 ( .A(n38550), .B(n38551), .Z(n35691) );
  XOR U35922 ( .A(n35721), .B(n35693), .Z(n35692) );
  AND U35923 ( .A(n38552), .B(n38553), .Z(n35693) );
  XOR U35924 ( .A(n35717), .B(n35722), .Z(n35721) );
  AND U35925 ( .A(n38554), .B(n38555), .Z(n35722) );
  XOR U35926 ( .A(n35719), .B(n35718), .Z(n35717) );
  AND U35927 ( .A(n38556), .B(n38557), .Z(n35718) );
  XOR U35928 ( .A(n35707), .B(n35720), .Z(n35719) );
  AND U35929 ( .A(n38558), .B(n38559), .Z(n35720) );
  XOR U35930 ( .A(n35709), .B(n35708), .Z(n35707) );
  AND U35931 ( .A(n38560), .B(n38561), .Z(n35708) );
  XOR U35932 ( .A(n35711), .B(n35710), .Z(n35709) );
  AND U35933 ( .A(n38562), .B(n38563), .Z(n35710) );
  XOR U35934 ( .A(n35713), .B(n35712), .Z(n35711) );
  AND U35935 ( .A(n38564), .B(n38565), .Z(n35712) );
  XOR U35936 ( .A(n35755), .B(n35714), .Z(n35713) );
  AND U35937 ( .A(n38566), .B(n38567), .Z(n35714) );
  XNOR U35938 ( .A(n35752), .B(n35756), .Z(n35755) );
  AND U35939 ( .A(n38568), .B(n38569), .Z(n35756) );
  XOR U35940 ( .A(n35751), .B(n35743), .Z(n35752) );
  AND U35941 ( .A(n38570), .B(n38571), .Z(n35743) );
  XNOR U35942 ( .A(n35746), .B(n35742), .Z(n35751) );
  AND U35943 ( .A(n38572), .B(n38573), .Z(n35742) );
  XOR U35944 ( .A(n35759), .B(n35747), .Z(n35746) );
  AND U35945 ( .A(n38574), .B(n38575), .Z(n35747) );
  XNOR U35946 ( .A(n35739), .B(n35760), .Z(n35759) );
  AND U35947 ( .A(n38576), .B(n38577), .Z(n35760) );
  XOR U35948 ( .A(n35738), .B(n35730), .Z(n35739) );
  AND U35949 ( .A(n38578), .B(n38579), .Z(n35730) );
  XNOR U35950 ( .A(n35733), .B(n35729), .Z(n35738) );
  AND U35951 ( .A(n38580), .B(n38581), .Z(n35729) );
  XOR U35952 ( .A(n38582), .B(n38583), .Z(n35733) );
  XOR U35953 ( .A(n38584), .B(n38585), .Z(n38583) );
  XOR U35954 ( .A(n38586), .B(n38587), .Z(n38585) );
  XNOR U35955 ( .A(n35776), .B(n35769), .Z(n38587) );
  XOR U35956 ( .A(n38588), .B(n38589), .Z(n35769) );
  XOR U35957 ( .A(n38590), .B(n38591), .Z(n38589) );
  NOR U35958 ( .A(n38592), .B(n38593), .Z(n38591) );
  NOR U35959 ( .A(n38594), .B(n38595), .Z(n38590) );
  AND U35960 ( .A(n38596), .B(n38597), .Z(n38595) );
  IV U35961 ( .A(n38598), .Z(n38594) );
  NOR U35962 ( .A(n38599), .B(n38600), .Z(n38598) );
  AND U35963 ( .A(n38592), .B(n38601), .Z(n38600) );
  AND U35964 ( .A(n38593), .B(n38602), .Z(n38599) );
  XNOR U35965 ( .A(n38603), .B(n38604), .Z(n38588) );
  AND U35966 ( .A(n38605), .B(n38606), .Z(n38604) );
  AND U35967 ( .A(n38607), .B(n38608), .Z(n38603) );
  NOR U35968 ( .A(n38609), .B(n38610), .Z(n38608) );
  IV U35969 ( .A(n38611), .Z(n38609) );
  NOR U35970 ( .A(n38612), .B(n38613), .Z(n38611) );
  NOR U35971 ( .A(n38614), .B(n38615), .Z(n38607) );
  AND U35972 ( .A(n38616), .B(n38617), .Z(n35776) );
  XOR U35973 ( .A(n35774), .B(n35775), .Z(n38586) );
  AND U35974 ( .A(n38618), .B(n38619), .Z(n35775) );
  AND U35975 ( .A(n38620), .B(n38621), .Z(n35774) );
  XOR U35976 ( .A(n38622), .B(n38623), .Z(n38584) );
  XOR U35977 ( .A(n35770), .B(n35771), .Z(n38623) );
  AND U35978 ( .A(n38624), .B(n38625), .Z(n35771) );
  AND U35979 ( .A(n38626), .B(n38627), .Z(n35770) );
  XOR U35980 ( .A(n35768), .B(n35766), .Z(n38622) );
  AND U35981 ( .A(n38628), .B(n38629), .Z(n35766) );
  AND U35982 ( .A(n38630), .B(n38631), .Z(n35768) );
  XNOR U35983 ( .A(n35777), .B(n35734), .Z(n38582) );
  AND U35984 ( .A(n38632), .B(n38633), .Z(n35734) );
  AND U35985 ( .A(n38634), .B(n38635), .Z(n35777) );
  XOR U35986 ( .A(n38636), .B(n38637), .Z(n35790) );
  AND U35987 ( .A(n38636), .B(n38638), .Z(n38637) );
  XNOR U35988 ( .A(n38639), .B(n38640), .Z(n35793) );
  AND U35989 ( .A(n38639), .B(n38641), .Z(n38640) );
  XNOR U35990 ( .A(n38642), .B(n38643), .Z(n35796) );
  AND U35991 ( .A(n38642), .B(n38644), .Z(n38643) );
  XNOR U35992 ( .A(n38645), .B(n38646), .Z(n35799) );
  AND U35993 ( .A(n38645), .B(n38647), .Z(n38646) );
  XNOR U35994 ( .A(n38648), .B(n38649), .Z(n35802) );
  AND U35995 ( .A(n38650), .B(n38648), .Z(n38649) );
  XOR U35996 ( .A(n38651), .B(n38652), .Z(n35805) );
  NOR U35997 ( .A(n38653), .B(n38651), .Z(n38652) );
  XOR U35998 ( .A(n38654), .B(n38655), .Z(n35808) );
  NOR U35999 ( .A(n38656), .B(n38654), .Z(n38655) );
  XOR U36000 ( .A(n38657), .B(n38658), .Z(n35811) );
  NOR U36001 ( .A(n38659), .B(n38657), .Z(n38658) );
  XOR U36002 ( .A(n38660), .B(n38661), .Z(n35814) );
  NOR U36003 ( .A(n38662), .B(n38660), .Z(n38661) );
  XOR U36004 ( .A(n38663), .B(n38664), .Z(n35817) );
  NOR U36005 ( .A(n38665), .B(n38663), .Z(n38664) );
  XOR U36006 ( .A(n38666), .B(n38667), .Z(n35820) );
  NOR U36007 ( .A(n38668), .B(n38666), .Z(n38667) );
  XOR U36008 ( .A(n38669), .B(n38670), .Z(n35823) );
  NOR U36009 ( .A(n38671), .B(n38669), .Z(n38670) );
  XOR U36010 ( .A(n38672), .B(n38673), .Z(n35826) );
  NOR U36011 ( .A(n38674), .B(n38672), .Z(n38673) );
  XOR U36012 ( .A(n38675), .B(n38676), .Z(n35829) );
  NOR U36013 ( .A(n38677), .B(n38675), .Z(n38676) );
  XOR U36014 ( .A(n38678), .B(n38679), .Z(n35832) );
  NOR U36015 ( .A(n38680), .B(n38678), .Z(n38679) );
  XOR U36016 ( .A(n38681), .B(n38682), .Z(n35835) );
  NOR U36017 ( .A(n38683), .B(n38681), .Z(n38682) );
  XOR U36018 ( .A(n38684), .B(n38685), .Z(n35838) );
  NOR U36019 ( .A(n38686), .B(n38684), .Z(n38685) );
  XOR U36020 ( .A(n38687), .B(n38688), .Z(n35841) );
  NOR U36021 ( .A(n38689), .B(n38687), .Z(n38688) );
  XOR U36022 ( .A(n38690), .B(n38691), .Z(n35844) );
  NOR U36023 ( .A(n38692), .B(n38690), .Z(n38691) );
  XOR U36024 ( .A(n38693), .B(n38694), .Z(n35847) );
  NOR U36025 ( .A(n38695), .B(n38693), .Z(n38694) );
  XOR U36026 ( .A(n38696), .B(n38697), .Z(n35850) );
  NOR U36027 ( .A(n38698), .B(n38696), .Z(n38697) );
  XOR U36028 ( .A(n38699), .B(n38700), .Z(n35853) );
  NOR U36029 ( .A(n38701), .B(n38699), .Z(n38700) );
  XOR U36030 ( .A(n38702), .B(n38703), .Z(n35856) );
  NOR U36031 ( .A(n38704), .B(n38702), .Z(n38703) );
  XOR U36032 ( .A(n38705), .B(n38706), .Z(n35859) );
  NOR U36033 ( .A(n38707), .B(n38705), .Z(n38706) );
  XOR U36034 ( .A(n38708), .B(n38709), .Z(n35862) );
  NOR U36035 ( .A(n38710), .B(n38708), .Z(n38709) );
  XOR U36036 ( .A(n38711), .B(n38712), .Z(n35865) );
  NOR U36037 ( .A(n38713), .B(n38711), .Z(n38712) );
  XOR U36038 ( .A(n38714), .B(n38715), .Z(n35868) );
  NOR U36039 ( .A(n38716), .B(n38714), .Z(n38715) );
  XOR U36040 ( .A(n38717), .B(n38718), .Z(n35871) );
  NOR U36041 ( .A(n38719), .B(n38717), .Z(n38718) );
  XOR U36042 ( .A(n38720), .B(n38721), .Z(n35874) );
  NOR U36043 ( .A(n38722), .B(n38720), .Z(n38721) );
  XOR U36044 ( .A(n38723), .B(n38724), .Z(n35877) );
  NOR U36045 ( .A(n38725), .B(n38723), .Z(n38724) );
  XOR U36046 ( .A(n38726), .B(n38727), .Z(n35880) );
  NOR U36047 ( .A(n38728), .B(n38726), .Z(n38727) );
  XOR U36048 ( .A(n38729), .B(n38730), .Z(n35883) );
  NOR U36049 ( .A(n38731), .B(n38729), .Z(n38730) );
  XOR U36050 ( .A(n38732), .B(n38733), .Z(n35886) );
  NOR U36051 ( .A(n38734), .B(n38732), .Z(n38733) );
  XOR U36052 ( .A(n38735), .B(n38736), .Z(n35889) );
  NOR U36053 ( .A(n38737), .B(n38735), .Z(n38736) );
  XOR U36054 ( .A(n38738), .B(n38739), .Z(n35892) );
  NOR U36055 ( .A(n38740), .B(n38738), .Z(n38739) );
  XOR U36056 ( .A(n38741), .B(n38742), .Z(n35895) );
  NOR U36057 ( .A(n38743), .B(n38741), .Z(n38742) );
  XOR U36058 ( .A(n38744), .B(n38745), .Z(n35898) );
  NOR U36059 ( .A(n38746), .B(n38744), .Z(n38745) );
  XOR U36060 ( .A(n38747), .B(n38748), .Z(n35901) );
  NOR U36061 ( .A(n38749), .B(n38747), .Z(n38748) );
  XOR U36062 ( .A(n38750), .B(n38751), .Z(n35904) );
  NOR U36063 ( .A(n38752), .B(n38750), .Z(n38751) );
  XOR U36064 ( .A(n38753), .B(n38754), .Z(n35907) );
  NOR U36065 ( .A(n38755), .B(n38753), .Z(n38754) );
  XOR U36066 ( .A(n38756), .B(n38757), .Z(n35910) );
  NOR U36067 ( .A(n38758), .B(n38756), .Z(n38757) );
  XOR U36068 ( .A(n38759), .B(n38760), .Z(n35913) );
  NOR U36069 ( .A(n38761), .B(n38759), .Z(n38760) );
  XOR U36070 ( .A(n38762), .B(n38763), .Z(n35916) );
  NOR U36071 ( .A(n38764), .B(n38762), .Z(n38763) );
  XOR U36072 ( .A(n38765), .B(n38766), .Z(n35919) );
  NOR U36073 ( .A(n38767), .B(n38765), .Z(n38766) );
  XOR U36074 ( .A(n38768), .B(n38769), .Z(n35922) );
  NOR U36075 ( .A(n38770), .B(n38768), .Z(n38769) );
  XOR U36076 ( .A(n38771), .B(n38772), .Z(n35925) );
  NOR U36077 ( .A(n38773), .B(n38771), .Z(n38772) );
  XOR U36078 ( .A(n38774), .B(n38775), .Z(n35928) );
  NOR U36079 ( .A(n38776), .B(n38774), .Z(n38775) );
  XOR U36080 ( .A(n38777), .B(n38778), .Z(n35931) );
  NOR U36081 ( .A(n38779), .B(n38777), .Z(n38778) );
  XOR U36082 ( .A(n38780), .B(n38781), .Z(n35934) );
  NOR U36083 ( .A(n38782), .B(n38780), .Z(n38781) );
  XOR U36084 ( .A(n38783), .B(n38784), .Z(n35937) );
  NOR U36085 ( .A(n38785), .B(n38783), .Z(n38784) );
  XOR U36086 ( .A(n38786), .B(n38787), .Z(n35940) );
  NOR U36087 ( .A(n38788), .B(n38786), .Z(n38787) );
  XOR U36088 ( .A(n38789), .B(n38790), .Z(n35943) );
  NOR U36089 ( .A(n38791), .B(n38789), .Z(n38790) );
  XOR U36090 ( .A(n38792), .B(n38793), .Z(n35946) );
  NOR U36091 ( .A(n38794), .B(n38792), .Z(n38793) );
  XOR U36092 ( .A(n38795), .B(n38796), .Z(n35949) );
  NOR U36093 ( .A(n38797), .B(n38795), .Z(n38796) );
  XOR U36094 ( .A(n38798), .B(n38799), .Z(n35952) );
  NOR U36095 ( .A(n38800), .B(n38798), .Z(n38799) );
  XOR U36096 ( .A(n38801), .B(n38802), .Z(n35955) );
  NOR U36097 ( .A(n38803), .B(n38801), .Z(n38802) );
  XOR U36098 ( .A(n38804), .B(n38805), .Z(n35958) );
  NOR U36099 ( .A(n38806), .B(n38804), .Z(n38805) );
  XOR U36100 ( .A(n38807), .B(n38808), .Z(n35961) );
  NOR U36101 ( .A(n38809), .B(n38807), .Z(n38808) );
  XOR U36102 ( .A(n38810), .B(n38811), .Z(n35964) );
  NOR U36103 ( .A(n38812), .B(n38810), .Z(n38811) );
  XOR U36104 ( .A(n38813), .B(n38814), .Z(n35967) );
  NOR U36105 ( .A(n38815), .B(n38813), .Z(n38814) );
  XOR U36106 ( .A(n38816), .B(n38817), .Z(n35970) );
  NOR U36107 ( .A(n38818), .B(n38816), .Z(n38817) );
  XOR U36108 ( .A(n38819), .B(n38820), .Z(n35973) );
  NOR U36109 ( .A(n38821), .B(n38819), .Z(n38820) );
  XOR U36110 ( .A(n38822), .B(n38823), .Z(n35976) );
  NOR U36111 ( .A(n38824), .B(n38822), .Z(n38823) );
  XOR U36112 ( .A(n38825), .B(n38826), .Z(n35979) );
  NOR U36113 ( .A(n38827), .B(n38825), .Z(n38826) );
  XOR U36114 ( .A(n38828), .B(n38829), .Z(n35982) );
  NOR U36115 ( .A(n38830), .B(n38828), .Z(n38829) );
  XOR U36116 ( .A(n38831), .B(n38832), .Z(n35985) );
  NOR U36117 ( .A(n38833), .B(n38831), .Z(n38832) );
  XOR U36118 ( .A(n38834), .B(n38835), .Z(n35988) );
  NOR U36119 ( .A(n38836), .B(n38834), .Z(n38835) );
  XOR U36120 ( .A(n38837), .B(n38838), .Z(n35991) );
  NOR U36121 ( .A(n38839), .B(n38837), .Z(n38838) );
  XOR U36122 ( .A(n38840), .B(n38841), .Z(n35994) );
  NOR U36123 ( .A(n38842), .B(n38840), .Z(n38841) );
  XOR U36124 ( .A(n38843), .B(n38844), .Z(n35997) );
  NOR U36125 ( .A(n38845), .B(n38843), .Z(n38844) );
  XOR U36126 ( .A(n38846), .B(n38847), .Z(n36000) );
  NOR U36127 ( .A(n38848), .B(n38846), .Z(n38847) );
  XOR U36128 ( .A(n38849), .B(n38850), .Z(n36003) );
  NOR U36129 ( .A(n38851), .B(n38849), .Z(n38850) );
  XOR U36130 ( .A(n38852), .B(n38853), .Z(n36006) );
  NOR U36131 ( .A(n38854), .B(n38852), .Z(n38853) );
  XOR U36132 ( .A(n38855), .B(n38856), .Z(n36009) );
  NOR U36133 ( .A(n38857), .B(n38855), .Z(n38856) );
  XOR U36134 ( .A(n38858), .B(n38859), .Z(n36012) );
  NOR U36135 ( .A(n38860), .B(n38858), .Z(n38859) );
  XOR U36136 ( .A(n38861), .B(n38862), .Z(n36015) );
  NOR U36137 ( .A(n38863), .B(n38861), .Z(n38862) );
  XOR U36138 ( .A(n38864), .B(n38865), .Z(n36018) );
  NOR U36139 ( .A(n38866), .B(n38864), .Z(n38865) );
  XOR U36140 ( .A(n38867), .B(n38868), .Z(n36021) );
  NOR U36141 ( .A(n38869), .B(n38867), .Z(n38868) );
  XOR U36142 ( .A(n38870), .B(n38871), .Z(n36024) );
  NOR U36143 ( .A(n38872), .B(n38870), .Z(n38871) );
  XOR U36144 ( .A(n38873), .B(n38874), .Z(n36027) );
  NOR U36145 ( .A(n38875), .B(n38873), .Z(n38874) );
  XOR U36146 ( .A(n38876), .B(n38877), .Z(n36030) );
  NOR U36147 ( .A(n38878), .B(n38876), .Z(n38877) );
  XOR U36148 ( .A(n38879), .B(n38880), .Z(n36033) );
  NOR U36149 ( .A(n38881), .B(n38879), .Z(n38880) );
  XOR U36150 ( .A(n38882), .B(n38883), .Z(n36036) );
  NOR U36151 ( .A(n38884), .B(n38882), .Z(n38883) );
  XOR U36152 ( .A(n38885), .B(n38886), .Z(n36039) );
  NOR U36153 ( .A(n38887), .B(n38885), .Z(n38886) );
  XOR U36154 ( .A(n38888), .B(n38889), .Z(n36042) );
  NOR U36155 ( .A(n38890), .B(n38888), .Z(n38889) );
  XOR U36156 ( .A(n38891), .B(n38892), .Z(n36045) );
  NOR U36157 ( .A(n38893), .B(n38891), .Z(n38892) );
  XOR U36158 ( .A(n38894), .B(n38895), .Z(n36048) );
  NOR U36159 ( .A(n38896), .B(n38894), .Z(n38895) );
  XOR U36160 ( .A(n38897), .B(n38898), .Z(n36051) );
  NOR U36161 ( .A(n38899), .B(n38897), .Z(n38898) );
  XOR U36162 ( .A(n38900), .B(n38901), .Z(n36054) );
  NOR U36163 ( .A(n38902), .B(n38900), .Z(n38901) );
  XOR U36164 ( .A(n38903), .B(n38904), .Z(n36057) );
  NOR U36165 ( .A(n38905), .B(n38903), .Z(n38904) );
  XOR U36166 ( .A(n38906), .B(n38907), .Z(n36060) );
  NOR U36167 ( .A(n38908), .B(n38906), .Z(n38907) );
  XOR U36168 ( .A(n38909), .B(n38910), .Z(n36063) );
  NOR U36169 ( .A(n38911), .B(n38909), .Z(n38910) );
  XOR U36170 ( .A(n38912), .B(n38913), .Z(n36066) );
  NOR U36171 ( .A(n38914), .B(n38912), .Z(n38913) );
  XOR U36172 ( .A(n38915), .B(n38916), .Z(n36069) );
  NOR U36173 ( .A(n38917), .B(n38915), .Z(n38916) );
  XOR U36174 ( .A(n38918), .B(n38919), .Z(n36072) );
  NOR U36175 ( .A(n38920), .B(n38918), .Z(n38919) );
  XOR U36176 ( .A(n38921), .B(n38922), .Z(n36075) );
  NOR U36177 ( .A(n38923), .B(n38921), .Z(n38922) );
  XOR U36178 ( .A(n38924), .B(n38925), .Z(n36078) );
  NOR U36179 ( .A(n38926), .B(n38924), .Z(n38925) );
  XOR U36180 ( .A(n38927), .B(n38928), .Z(n36081) );
  NOR U36181 ( .A(n38929), .B(n38927), .Z(n38928) );
  XOR U36182 ( .A(n38930), .B(n38931), .Z(n36084) );
  NOR U36183 ( .A(n38932), .B(n38930), .Z(n38931) );
  XOR U36184 ( .A(n38933), .B(n38934), .Z(n36087) );
  NOR U36185 ( .A(n38935), .B(n38933), .Z(n38934) );
  XOR U36186 ( .A(n38936), .B(n38937), .Z(n36090) );
  NOR U36187 ( .A(n38938), .B(n38936), .Z(n38937) );
  XOR U36188 ( .A(n38939), .B(n38940), .Z(n36093) );
  NOR U36189 ( .A(n38941), .B(n38939), .Z(n38940) );
  XOR U36190 ( .A(n38942), .B(n38943), .Z(n36096) );
  NOR U36191 ( .A(n38944), .B(n38942), .Z(n38943) );
  XOR U36192 ( .A(n38945), .B(n38946), .Z(n36099) );
  NOR U36193 ( .A(n38947), .B(n38945), .Z(n38946) );
  XOR U36194 ( .A(n38948), .B(n38949), .Z(n36102) );
  NOR U36195 ( .A(n38950), .B(n38948), .Z(n38949) );
  XOR U36196 ( .A(n38951), .B(n38952), .Z(n36105) );
  NOR U36197 ( .A(n38953), .B(n38951), .Z(n38952) );
  XOR U36198 ( .A(n38954), .B(n38955), .Z(n36108) );
  NOR U36199 ( .A(n38956), .B(n38954), .Z(n38955) );
  XOR U36200 ( .A(n38957), .B(n38958), .Z(n36111) );
  NOR U36201 ( .A(n38959), .B(n38957), .Z(n38958) );
  XOR U36202 ( .A(n38960), .B(n38961), .Z(n36114) );
  NOR U36203 ( .A(n38962), .B(n38960), .Z(n38961) );
  XOR U36204 ( .A(n38963), .B(n38964), .Z(n36117) );
  NOR U36205 ( .A(n38965), .B(n38963), .Z(n38964) );
  XOR U36206 ( .A(n38966), .B(n38967), .Z(n36120) );
  NOR U36207 ( .A(n38968), .B(n38966), .Z(n38967) );
  XOR U36208 ( .A(n38969), .B(n38970), .Z(n36123) );
  NOR U36209 ( .A(n38971), .B(n38969), .Z(n38970) );
  XOR U36210 ( .A(n38972), .B(n38973), .Z(n36126) );
  NOR U36211 ( .A(n38974), .B(n38972), .Z(n38973) );
  XOR U36212 ( .A(n38975), .B(n38976), .Z(n36129) );
  NOR U36213 ( .A(n38977), .B(n38975), .Z(n38976) );
  XOR U36214 ( .A(n38978), .B(n38979), .Z(n36132) );
  NOR U36215 ( .A(n38980), .B(n38978), .Z(n38979) );
  XOR U36216 ( .A(n38981), .B(n38982), .Z(n36135) );
  NOR U36217 ( .A(n38983), .B(n38981), .Z(n38982) );
  XOR U36218 ( .A(n38984), .B(n38985), .Z(n36138) );
  NOR U36219 ( .A(n38986), .B(n38984), .Z(n38985) );
  XOR U36220 ( .A(n38987), .B(n38988), .Z(n36141) );
  NOR U36221 ( .A(n38989), .B(n38987), .Z(n38988) );
  XOR U36222 ( .A(n38990), .B(n38991), .Z(n36144) );
  NOR U36223 ( .A(n38992), .B(n38990), .Z(n38991) );
  XOR U36224 ( .A(n38993), .B(n38994), .Z(n36147) );
  NOR U36225 ( .A(n38995), .B(n38993), .Z(n38994) );
  XOR U36226 ( .A(n38996), .B(n38997), .Z(n36150) );
  NOR U36227 ( .A(n38998), .B(n38996), .Z(n38997) );
  XOR U36228 ( .A(n38999), .B(n39000), .Z(n36153) );
  NOR U36229 ( .A(n39001), .B(n38999), .Z(n39000) );
  XOR U36230 ( .A(n39002), .B(n39003), .Z(n36156) );
  NOR U36231 ( .A(n39004), .B(n39002), .Z(n39003) );
  XOR U36232 ( .A(n39005), .B(n39006), .Z(n36159) );
  NOR U36233 ( .A(n39007), .B(n39005), .Z(n39006) );
  XOR U36234 ( .A(n39008), .B(n39009), .Z(n36162) );
  NOR U36235 ( .A(n39010), .B(n39008), .Z(n39009) );
  XOR U36236 ( .A(n39011), .B(n39012), .Z(n36165) );
  NOR U36237 ( .A(n39013), .B(n39011), .Z(n39012) );
  XOR U36238 ( .A(n39014), .B(n39015), .Z(n36168) );
  NOR U36239 ( .A(n39016), .B(n39014), .Z(n39015) );
  XOR U36240 ( .A(n39017), .B(n39018), .Z(n36171) );
  NOR U36241 ( .A(n39019), .B(n39017), .Z(n39018) );
  XOR U36242 ( .A(n39020), .B(n39021), .Z(n36174) );
  NOR U36243 ( .A(n39022), .B(n39020), .Z(n39021) );
  XOR U36244 ( .A(n39023), .B(n39024), .Z(n36177) );
  NOR U36245 ( .A(n39025), .B(n39023), .Z(n39024) );
  XOR U36246 ( .A(n39026), .B(n39027), .Z(n36180) );
  NOR U36247 ( .A(n39028), .B(n39026), .Z(n39027) );
  XOR U36248 ( .A(n39029), .B(n39030), .Z(n36183) );
  NOR U36249 ( .A(n39031), .B(n39029), .Z(n39030) );
  XOR U36250 ( .A(n39032), .B(n39033), .Z(n36186) );
  NOR U36251 ( .A(n39034), .B(n39032), .Z(n39033) );
  XOR U36252 ( .A(n39035), .B(n39036), .Z(n36189) );
  NOR U36253 ( .A(n39037), .B(n39035), .Z(n39036) );
  XOR U36254 ( .A(n39038), .B(n39039), .Z(n36192) );
  NOR U36255 ( .A(n39040), .B(n39038), .Z(n39039) );
  XOR U36256 ( .A(n39041), .B(n39042), .Z(n36195) );
  NOR U36257 ( .A(n39043), .B(n39041), .Z(n39042) );
  XOR U36258 ( .A(n39044), .B(n39045), .Z(n36198) );
  NOR U36259 ( .A(n39046), .B(n39044), .Z(n39045) );
  XOR U36260 ( .A(n39047), .B(n39048), .Z(n36201) );
  NOR U36261 ( .A(n39049), .B(n39047), .Z(n39048) );
  XOR U36262 ( .A(n39050), .B(n39051), .Z(n36204) );
  NOR U36263 ( .A(n39052), .B(n39050), .Z(n39051) );
  XOR U36264 ( .A(n39053), .B(n39054), .Z(n36207) );
  NOR U36265 ( .A(n39055), .B(n39053), .Z(n39054) );
  XOR U36266 ( .A(n39056), .B(n39057), .Z(n36210) );
  NOR U36267 ( .A(n39058), .B(n39056), .Z(n39057) );
  XOR U36268 ( .A(n39059), .B(n39060), .Z(n36213) );
  NOR U36269 ( .A(n39061), .B(n39059), .Z(n39060) );
  XOR U36270 ( .A(n39062), .B(n39063), .Z(n36216) );
  NOR U36271 ( .A(n39064), .B(n39062), .Z(n39063) );
  XOR U36272 ( .A(n39065), .B(n39066), .Z(n36219) );
  NOR U36273 ( .A(n39067), .B(n39065), .Z(n39066) );
  XOR U36274 ( .A(n39068), .B(n39069), .Z(n36222) );
  NOR U36275 ( .A(n39070), .B(n39068), .Z(n39069) );
  XOR U36276 ( .A(n39071), .B(n39072), .Z(n36225) );
  NOR U36277 ( .A(n39073), .B(n39071), .Z(n39072) );
  XOR U36278 ( .A(n39074), .B(n39075), .Z(n36228) );
  NOR U36279 ( .A(n39076), .B(n39074), .Z(n39075) );
  XOR U36280 ( .A(n39077), .B(n39078), .Z(n36231) );
  NOR U36281 ( .A(n39079), .B(n39077), .Z(n39078) );
  XOR U36282 ( .A(n39080), .B(n39081), .Z(n36234) );
  NOR U36283 ( .A(n39082), .B(n39080), .Z(n39081) );
  XOR U36284 ( .A(n39083), .B(n39084), .Z(n36237) );
  NOR U36285 ( .A(n39085), .B(n39083), .Z(n39084) );
  XOR U36286 ( .A(n39086), .B(n39087), .Z(n36240) );
  NOR U36287 ( .A(n39088), .B(n39086), .Z(n39087) );
  XOR U36288 ( .A(n39089), .B(n39090), .Z(n36243) );
  NOR U36289 ( .A(n39091), .B(n39089), .Z(n39090) );
  XOR U36290 ( .A(n39092), .B(n39093), .Z(n36246) );
  NOR U36291 ( .A(n39094), .B(n39092), .Z(n39093) );
  XOR U36292 ( .A(n39095), .B(n39096), .Z(n36249) );
  NOR U36293 ( .A(n39097), .B(n39095), .Z(n39096) );
  XOR U36294 ( .A(n39098), .B(n39099), .Z(n36252) );
  NOR U36295 ( .A(n39100), .B(n39098), .Z(n39099) );
  XOR U36296 ( .A(n39101), .B(n39102), .Z(n36255) );
  NOR U36297 ( .A(n39103), .B(n39101), .Z(n39102) );
  XOR U36298 ( .A(n39104), .B(n39105), .Z(n36258) );
  NOR U36299 ( .A(n39106), .B(n39104), .Z(n39105) );
  XOR U36300 ( .A(n39107), .B(n39108), .Z(n36261) );
  NOR U36301 ( .A(n39109), .B(n39107), .Z(n39108) );
  XOR U36302 ( .A(n39110), .B(n39111), .Z(n36264) );
  NOR U36303 ( .A(n39112), .B(n39110), .Z(n39111) );
  XOR U36304 ( .A(n39113), .B(n39114), .Z(n36267) );
  NOR U36305 ( .A(n39115), .B(n39113), .Z(n39114) );
  XOR U36306 ( .A(n39116), .B(n39117), .Z(n36270) );
  NOR U36307 ( .A(n39118), .B(n39116), .Z(n39117) );
  XOR U36308 ( .A(n39119), .B(n39120), .Z(n36273) );
  NOR U36309 ( .A(n39121), .B(n39119), .Z(n39120) );
  XOR U36310 ( .A(n39122), .B(n39123), .Z(n36276) );
  NOR U36311 ( .A(n39124), .B(n39122), .Z(n39123) );
  XOR U36312 ( .A(n39125), .B(n39126), .Z(n36279) );
  NOR U36313 ( .A(n39127), .B(n39125), .Z(n39126) );
  XOR U36314 ( .A(n39128), .B(n39129), .Z(n36282) );
  NOR U36315 ( .A(n39130), .B(n39128), .Z(n39129) );
  XOR U36316 ( .A(n39131), .B(n39132), .Z(n36285) );
  NOR U36317 ( .A(n39133), .B(n39131), .Z(n39132) );
  XOR U36318 ( .A(n39134), .B(n39135), .Z(n36288) );
  NOR U36319 ( .A(n39136), .B(n39134), .Z(n39135) );
  XOR U36320 ( .A(n39137), .B(n39138), .Z(n36291) );
  NOR U36321 ( .A(n39139), .B(n39137), .Z(n39138) );
  XOR U36322 ( .A(n39140), .B(n39141), .Z(n36294) );
  NOR U36323 ( .A(n39142), .B(n39140), .Z(n39141) );
  XOR U36324 ( .A(n39143), .B(n39144), .Z(n36297) );
  NOR U36325 ( .A(n39145), .B(n39143), .Z(n39144) );
  XOR U36326 ( .A(n39146), .B(n39147), .Z(n36300) );
  NOR U36327 ( .A(n39148), .B(n39146), .Z(n39147) );
  XOR U36328 ( .A(n39149), .B(n39150), .Z(n36303) );
  NOR U36329 ( .A(n39151), .B(n39149), .Z(n39150) );
  XOR U36330 ( .A(n39152), .B(n39153), .Z(n36306) );
  NOR U36331 ( .A(n39154), .B(n39152), .Z(n39153) );
  XOR U36332 ( .A(n39155), .B(n39156), .Z(n36309) );
  NOR U36333 ( .A(n39157), .B(n39155), .Z(n39156) );
  XOR U36334 ( .A(n39158), .B(n39159), .Z(n36312) );
  NOR U36335 ( .A(n39160), .B(n39158), .Z(n39159) );
  XOR U36336 ( .A(n39161), .B(n39162), .Z(n36315) );
  NOR U36337 ( .A(n39163), .B(n39161), .Z(n39162) );
  XOR U36338 ( .A(n39164), .B(n39165), .Z(n36318) );
  NOR U36339 ( .A(n39166), .B(n39164), .Z(n39165) );
  XOR U36340 ( .A(n39167), .B(n39168), .Z(n36321) );
  NOR U36341 ( .A(n39169), .B(n39167), .Z(n39168) );
  XOR U36342 ( .A(n39170), .B(n39171), .Z(n36324) );
  NOR U36343 ( .A(n39172), .B(n39170), .Z(n39171) );
  XOR U36344 ( .A(n39173), .B(n39174), .Z(n36327) );
  NOR U36345 ( .A(n39175), .B(n39173), .Z(n39174) );
  XOR U36346 ( .A(n39176), .B(n39177), .Z(n36330) );
  NOR U36347 ( .A(n39178), .B(n39176), .Z(n39177) );
  XOR U36348 ( .A(n39179), .B(n39180), .Z(n36333) );
  NOR U36349 ( .A(n39181), .B(n39179), .Z(n39180) );
  XOR U36350 ( .A(n39182), .B(n39183), .Z(n36336) );
  NOR U36351 ( .A(n39184), .B(n39182), .Z(n39183) );
  XOR U36352 ( .A(n39185), .B(n39186), .Z(n36339) );
  NOR U36353 ( .A(n39187), .B(n39185), .Z(n39186) );
  XOR U36354 ( .A(n39188), .B(n39189), .Z(n36342) );
  NOR U36355 ( .A(n39190), .B(n39188), .Z(n39189) );
  XOR U36356 ( .A(n39191), .B(n39192), .Z(n36345) );
  NOR U36357 ( .A(n39193), .B(n39191), .Z(n39192) );
  XOR U36358 ( .A(n39194), .B(n39195), .Z(n36348) );
  NOR U36359 ( .A(n39196), .B(n39194), .Z(n39195) );
  XOR U36360 ( .A(n39197), .B(n39198), .Z(n36351) );
  NOR U36361 ( .A(n39199), .B(n39197), .Z(n39198) );
  XOR U36362 ( .A(n39200), .B(n39201), .Z(n36354) );
  NOR U36363 ( .A(n39202), .B(n39200), .Z(n39201) );
  XOR U36364 ( .A(n39203), .B(n39204), .Z(n36357) );
  NOR U36365 ( .A(n39205), .B(n39203), .Z(n39204) );
  XOR U36366 ( .A(n39206), .B(n39207), .Z(n36360) );
  NOR U36367 ( .A(n39208), .B(n39206), .Z(n39207) );
  XOR U36368 ( .A(n39209), .B(n39210), .Z(n36363) );
  NOR U36369 ( .A(n39211), .B(n39209), .Z(n39210) );
  XOR U36370 ( .A(n39212), .B(n39213), .Z(n36366) );
  NOR U36371 ( .A(n39214), .B(n39212), .Z(n39213) );
  XOR U36372 ( .A(n39215), .B(n39216), .Z(n36369) );
  NOR U36373 ( .A(n39217), .B(n39215), .Z(n39216) );
  XOR U36374 ( .A(n39218), .B(n39219), .Z(n36372) );
  NOR U36375 ( .A(n39220), .B(n39218), .Z(n39219) );
  XOR U36376 ( .A(n39221), .B(n39222), .Z(n36375) );
  NOR U36377 ( .A(n39223), .B(n39221), .Z(n39222) );
  XOR U36378 ( .A(n39224), .B(n39225), .Z(n36378) );
  NOR U36379 ( .A(n39226), .B(n39224), .Z(n39225) );
  XOR U36380 ( .A(n39227), .B(n39228), .Z(n36381) );
  NOR U36381 ( .A(n39229), .B(n39227), .Z(n39228) );
  XOR U36382 ( .A(n39230), .B(n39231), .Z(n36384) );
  NOR U36383 ( .A(n39232), .B(n39230), .Z(n39231) );
  XOR U36384 ( .A(n39233), .B(n39234), .Z(n36387) );
  NOR U36385 ( .A(n39235), .B(n39233), .Z(n39234) );
  XOR U36386 ( .A(n39236), .B(n39237), .Z(n36390) );
  NOR U36387 ( .A(n39238), .B(n39236), .Z(n39237) );
  XOR U36388 ( .A(n39239), .B(n39240), .Z(n36393) );
  NOR U36389 ( .A(n39241), .B(n39239), .Z(n39240) );
  XOR U36390 ( .A(n39242), .B(n39243), .Z(n36396) );
  NOR U36391 ( .A(n39244), .B(n39242), .Z(n39243) );
  XOR U36392 ( .A(n39245), .B(n39246), .Z(n36399) );
  NOR U36393 ( .A(n39247), .B(n39245), .Z(n39246) );
  XOR U36394 ( .A(n39248), .B(n39249), .Z(n36402) );
  NOR U36395 ( .A(n39250), .B(n39248), .Z(n39249) );
  XOR U36396 ( .A(n39251), .B(n39252), .Z(n36405) );
  NOR U36397 ( .A(n39253), .B(n39251), .Z(n39252) );
  XOR U36398 ( .A(n39254), .B(n39255), .Z(n36408) );
  NOR U36399 ( .A(n39256), .B(n39254), .Z(n39255) );
  XOR U36400 ( .A(n39257), .B(n39258), .Z(n36411) );
  NOR U36401 ( .A(n39259), .B(n39257), .Z(n39258) );
  XOR U36402 ( .A(n39260), .B(n39261), .Z(n36414) );
  NOR U36403 ( .A(n39262), .B(n39260), .Z(n39261) );
  XOR U36404 ( .A(n39263), .B(n39264), .Z(n36417) );
  NOR U36405 ( .A(n39265), .B(n39263), .Z(n39264) );
  XOR U36406 ( .A(n39266), .B(n39267), .Z(n36420) );
  NOR U36407 ( .A(n39268), .B(n39266), .Z(n39267) );
  XOR U36408 ( .A(n39269), .B(n39270), .Z(n36423) );
  NOR U36409 ( .A(n39271), .B(n39269), .Z(n39270) );
  XOR U36410 ( .A(n39272), .B(n39273), .Z(n36426) );
  NOR U36411 ( .A(n39274), .B(n39272), .Z(n39273) );
  XOR U36412 ( .A(n39275), .B(n39276), .Z(n36429) );
  NOR U36413 ( .A(n39277), .B(n39275), .Z(n39276) );
  XOR U36414 ( .A(n39278), .B(n39279), .Z(n36432) );
  NOR U36415 ( .A(n39280), .B(n39278), .Z(n39279) );
  XOR U36416 ( .A(n39281), .B(n39282), .Z(n36435) );
  NOR U36417 ( .A(n39283), .B(n39281), .Z(n39282) );
  XOR U36418 ( .A(n39284), .B(n39285), .Z(n36438) );
  NOR U36419 ( .A(n39286), .B(n39284), .Z(n39285) );
  XOR U36420 ( .A(n39287), .B(n39288), .Z(n36441) );
  NOR U36421 ( .A(n39289), .B(n39287), .Z(n39288) );
  XOR U36422 ( .A(n39290), .B(n39291), .Z(n36444) );
  NOR U36423 ( .A(n39292), .B(n39290), .Z(n39291) );
  XOR U36424 ( .A(n39293), .B(n39294), .Z(n36447) );
  NOR U36425 ( .A(n39295), .B(n39293), .Z(n39294) );
  XOR U36426 ( .A(n39296), .B(n39297), .Z(n36450) );
  NOR U36427 ( .A(n39298), .B(n39296), .Z(n39297) );
  XOR U36428 ( .A(n39299), .B(n39300), .Z(n36453) );
  NOR U36429 ( .A(n39301), .B(n39299), .Z(n39300) );
  XOR U36430 ( .A(n39302), .B(n39303), .Z(n36456) );
  NOR U36431 ( .A(n39304), .B(n39302), .Z(n39303) );
  XOR U36432 ( .A(n39305), .B(n39306), .Z(n36459) );
  NOR U36433 ( .A(n39307), .B(n39305), .Z(n39306) );
  XOR U36434 ( .A(n39308), .B(n39309), .Z(n36462) );
  NOR U36435 ( .A(n39310), .B(n39308), .Z(n39309) );
  XOR U36436 ( .A(n39311), .B(n39312), .Z(n36465) );
  NOR U36437 ( .A(n39313), .B(n39311), .Z(n39312) );
  XOR U36438 ( .A(n39314), .B(n39315), .Z(n36468) );
  NOR U36439 ( .A(n39316), .B(n39314), .Z(n39315) );
  XOR U36440 ( .A(n39317), .B(n39318), .Z(n36471) );
  NOR U36441 ( .A(n39319), .B(n39317), .Z(n39318) );
  XOR U36442 ( .A(n39320), .B(n39321), .Z(n36474) );
  NOR U36443 ( .A(n39322), .B(n39320), .Z(n39321) );
  XOR U36444 ( .A(n39323), .B(n39324), .Z(n36477) );
  NOR U36445 ( .A(n39325), .B(n39323), .Z(n39324) );
  XOR U36446 ( .A(n39326), .B(n39327), .Z(n36480) );
  NOR U36447 ( .A(n39328), .B(n39326), .Z(n39327) );
  XOR U36448 ( .A(n39329), .B(n39330), .Z(n36483) );
  NOR U36449 ( .A(n39331), .B(n39329), .Z(n39330) );
  XOR U36450 ( .A(n39332), .B(n39333), .Z(n36486) );
  NOR U36451 ( .A(n39334), .B(n39332), .Z(n39333) );
  XOR U36452 ( .A(n39335), .B(n39336), .Z(n36489) );
  NOR U36453 ( .A(n39337), .B(n39335), .Z(n39336) );
  XOR U36454 ( .A(n39338), .B(n39339), .Z(n36492) );
  NOR U36455 ( .A(n39340), .B(n39338), .Z(n39339) );
  XOR U36456 ( .A(n39341), .B(n39342), .Z(n36495) );
  NOR U36457 ( .A(n39343), .B(n39341), .Z(n39342) );
  XOR U36458 ( .A(n39344), .B(n39345), .Z(n36498) );
  NOR U36459 ( .A(n39346), .B(n39344), .Z(n39345) );
  XOR U36460 ( .A(n39347), .B(n39348), .Z(n36501) );
  NOR U36461 ( .A(n39349), .B(n39347), .Z(n39348) );
  XOR U36462 ( .A(n39350), .B(n39351), .Z(n36504) );
  NOR U36463 ( .A(n39352), .B(n39350), .Z(n39351) );
  XOR U36464 ( .A(n39353), .B(n39354), .Z(n36507) );
  NOR U36465 ( .A(n39355), .B(n39353), .Z(n39354) );
  XOR U36466 ( .A(n39356), .B(n39357), .Z(n36510) );
  NOR U36467 ( .A(n39358), .B(n39356), .Z(n39357) );
  XOR U36468 ( .A(n39359), .B(n39360), .Z(n36513) );
  NOR U36469 ( .A(n39361), .B(n39359), .Z(n39360) );
  XOR U36470 ( .A(n39362), .B(n39363), .Z(n36516) );
  NOR U36471 ( .A(n39364), .B(n39362), .Z(n39363) );
  XOR U36472 ( .A(n39365), .B(n39366), .Z(n36519) );
  NOR U36473 ( .A(n39367), .B(n39365), .Z(n39366) );
  XOR U36474 ( .A(n39368), .B(n39369), .Z(n36522) );
  NOR U36475 ( .A(n39370), .B(n39368), .Z(n39369) );
  XOR U36476 ( .A(n39371), .B(n39372), .Z(n36525) );
  NOR U36477 ( .A(n39373), .B(n39371), .Z(n39372) );
  XOR U36478 ( .A(n39374), .B(n39375), .Z(n36528) );
  NOR U36479 ( .A(n39376), .B(n39374), .Z(n39375) );
  XOR U36480 ( .A(n39377), .B(n39378), .Z(n36531) );
  NOR U36481 ( .A(n39379), .B(n39377), .Z(n39378) );
  XOR U36482 ( .A(n39380), .B(n39381), .Z(n36534) );
  NOR U36483 ( .A(n39382), .B(n39380), .Z(n39381) );
  XOR U36484 ( .A(n39383), .B(n39384), .Z(n36537) );
  NOR U36485 ( .A(n39385), .B(n39383), .Z(n39384) );
  XOR U36486 ( .A(n39386), .B(n39387), .Z(n36540) );
  NOR U36487 ( .A(n39388), .B(n39386), .Z(n39387) );
  XOR U36488 ( .A(n39389), .B(n39390), .Z(n36543) );
  NOR U36489 ( .A(n39391), .B(n39389), .Z(n39390) );
  XOR U36490 ( .A(n39392), .B(n39393), .Z(n36546) );
  NOR U36491 ( .A(n39394), .B(n39392), .Z(n39393) );
  XOR U36492 ( .A(n39395), .B(n39396), .Z(n36549) );
  NOR U36493 ( .A(n39397), .B(n39395), .Z(n39396) );
  XOR U36494 ( .A(n39398), .B(n39399), .Z(n36552) );
  NOR U36495 ( .A(n39400), .B(n39398), .Z(n39399) );
  XOR U36496 ( .A(n39401), .B(n39402), .Z(n36555) );
  NOR U36497 ( .A(n39403), .B(n39401), .Z(n39402) );
  XOR U36498 ( .A(n39404), .B(n39405), .Z(n36558) );
  NOR U36499 ( .A(n39406), .B(n39404), .Z(n39405) );
  XOR U36500 ( .A(n39407), .B(n39408), .Z(n36561) );
  NOR U36501 ( .A(n39409), .B(n39407), .Z(n39408) );
  XOR U36502 ( .A(n39410), .B(n39411), .Z(n36564) );
  NOR U36503 ( .A(n39412), .B(n39410), .Z(n39411) );
  XOR U36504 ( .A(n39413), .B(n39414), .Z(n36567) );
  NOR U36505 ( .A(n39415), .B(n39413), .Z(n39414) );
  XOR U36506 ( .A(n39416), .B(n39417), .Z(n36570) );
  NOR U36507 ( .A(n39418), .B(n39416), .Z(n39417) );
  XOR U36508 ( .A(n39419), .B(n39420), .Z(n36573) );
  NOR U36509 ( .A(n39421), .B(n39419), .Z(n39420) );
  XOR U36510 ( .A(n39422), .B(n39423), .Z(n36576) );
  NOR U36511 ( .A(n39424), .B(n39422), .Z(n39423) );
  XOR U36512 ( .A(n39425), .B(n39426), .Z(n36579) );
  NOR U36513 ( .A(n39427), .B(n39425), .Z(n39426) );
  XOR U36514 ( .A(n39428), .B(n39429), .Z(n36582) );
  NOR U36515 ( .A(n39430), .B(n39428), .Z(n39429) );
  XOR U36516 ( .A(n39431), .B(n39432), .Z(n36585) );
  NOR U36517 ( .A(n39433), .B(n39431), .Z(n39432) );
  XOR U36518 ( .A(n39434), .B(n39435), .Z(n36588) );
  NOR U36519 ( .A(n39436), .B(n39434), .Z(n39435) );
  XOR U36520 ( .A(n39437), .B(n39438), .Z(n36591) );
  NOR U36521 ( .A(n39439), .B(n39437), .Z(n39438) );
  XOR U36522 ( .A(n39440), .B(n39441), .Z(n36594) );
  NOR U36523 ( .A(n39442), .B(n39440), .Z(n39441) );
  XOR U36524 ( .A(n39443), .B(n39444), .Z(n36597) );
  NOR U36525 ( .A(n39445), .B(n39443), .Z(n39444) );
  XOR U36526 ( .A(n39446), .B(n39447), .Z(n36600) );
  NOR U36527 ( .A(n39448), .B(n39446), .Z(n39447) );
  XOR U36528 ( .A(n39449), .B(n39450), .Z(n36603) );
  NOR U36529 ( .A(n39451), .B(n39449), .Z(n39450) );
  XOR U36530 ( .A(n39452), .B(n39453), .Z(n36606) );
  NOR U36531 ( .A(n39454), .B(n39452), .Z(n39453) );
  XOR U36532 ( .A(n39455), .B(n39456), .Z(n36609) );
  NOR U36533 ( .A(n39457), .B(n39455), .Z(n39456) );
  XOR U36534 ( .A(n39458), .B(n39459), .Z(n36612) );
  NOR U36535 ( .A(n39460), .B(n39458), .Z(n39459) );
  XOR U36536 ( .A(n39461), .B(n39462), .Z(n36615) );
  NOR U36537 ( .A(n39463), .B(n39461), .Z(n39462) );
  XOR U36538 ( .A(n39464), .B(n39465), .Z(n36618) );
  NOR U36539 ( .A(n39466), .B(n39464), .Z(n39465) );
  XOR U36540 ( .A(n39467), .B(n39468), .Z(n36621) );
  NOR U36541 ( .A(n39469), .B(n39467), .Z(n39468) );
  XOR U36542 ( .A(n39470), .B(n39471), .Z(n36624) );
  NOR U36543 ( .A(n39472), .B(n39470), .Z(n39471) );
  XOR U36544 ( .A(n39473), .B(n39474), .Z(n36627) );
  NOR U36545 ( .A(n39475), .B(n39473), .Z(n39474) );
  XOR U36546 ( .A(n39476), .B(n39477), .Z(n36630) );
  NOR U36547 ( .A(n39478), .B(n39476), .Z(n39477) );
  XOR U36548 ( .A(n39479), .B(n39480), .Z(n36633) );
  NOR U36549 ( .A(n39481), .B(n39479), .Z(n39480) );
  XOR U36550 ( .A(n39482), .B(n39483), .Z(n36636) );
  NOR U36551 ( .A(n39484), .B(n39482), .Z(n39483) );
  XOR U36552 ( .A(n39485), .B(n39486), .Z(n36639) );
  NOR U36553 ( .A(n39487), .B(n39485), .Z(n39486) );
  XOR U36554 ( .A(n39488), .B(n39489), .Z(n36642) );
  NOR U36555 ( .A(n39490), .B(n39488), .Z(n39489) );
  XOR U36556 ( .A(n39491), .B(n39492), .Z(n36645) );
  NOR U36557 ( .A(n39493), .B(n39491), .Z(n39492) );
  XOR U36558 ( .A(n39494), .B(n39495), .Z(n36648) );
  NOR U36559 ( .A(n39496), .B(n39494), .Z(n39495) );
  XOR U36560 ( .A(n39497), .B(n39498), .Z(n36651) );
  NOR U36561 ( .A(n39499), .B(n39497), .Z(n39498) );
  XOR U36562 ( .A(n39500), .B(n39501), .Z(n36654) );
  NOR U36563 ( .A(n39502), .B(n39500), .Z(n39501) );
  XOR U36564 ( .A(n39503), .B(n39504), .Z(n36657) );
  NOR U36565 ( .A(n39505), .B(n39503), .Z(n39504) );
  XOR U36566 ( .A(n39506), .B(n39507), .Z(n36660) );
  NOR U36567 ( .A(n39508), .B(n39506), .Z(n39507) );
  XOR U36568 ( .A(n39509), .B(n39510), .Z(n36663) );
  NOR U36569 ( .A(n39511), .B(n39509), .Z(n39510) );
  XOR U36570 ( .A(n39512), .B(n39513), .Z(n36666) );
  NOR U36571 ( .A(n39514), .B(n39512), .Z(n39513) );
  XOR U36572 ( .A(n39515), .B(n39516), .Z(n36669) );
  NOR U36573 ( .A(n39517), .B(n39515), .Z(n39516) );
  XOR U36574 ( .A(n39518), .B(n39519), .Z(n36672) );
  NOR U36575 ( .A(n39520), .B(n39518), .Z(n39519) );
  XOR U36576 ( .A(n39521), .B(n39522), .Z(n36675) );
  NOR U36577 ( .A(n39523), .B(n39521), .Z(n39522) );
  XOR U36578 ( .A(n39524), .B(n39525), .Z(n36678) );
  NOR U36579 ( .A(n39526), .B(n39524), .Z(n39525) );
  XOR U36580 ( .A(n39527), .B(n39528), .Z(n36681) );
  NOR U36581 ( .A(n39529), .B(n39527), .Z(n39528) );
  XOR U36582 ( .A(n39530), .B(n39531), .Z(n36684) );
  NOR U36583 ( .A(n39532), .B(n39530), .Z(n39531) );
  XOR U36584 ( .A(n39533), .B(n39534), .Z(n36687) );
  NOR U36585 ( .A(n39535), .B(n39533), .Z(n39534) );
  XOR U36586 ( .A(n39536), .B(n39537), .Z(n36690) );
  NOR U36587 ( .A(n39538), .B(n39536), .Z(n39537) );
  XOR U36588 ( .A(n39539), .B(n39540), .Z(n36693) );
  NOR U36589 ( .A(n39541), .B(n39539), .Z(n39540) );
  XOR U36590 ( .A(n39542), .B(n39543), .Z(n36696) );
  NOR U36591 ( .A(n39544), .B(n39542), .Z(n39543) );
  XOR U36592 ( .A(n39545), .B(n39546), .Z(n36699) );
  NOR U36593 ( .A(n39547), .B(n39545), .Z(n39546) );
  XOR U36594 ( .A(n39548), .B(n39549), .Z(n36702) );
  NOR U36595 ( .A(n39550), .B(n39548), .Z(n39549) );
  XOR U36596 ( .A(n39551), .B(n39552), .Z(n36705) );
  NOR U36597 ( .A(n39553), .B(n39551), .Z(n39552) );
  XOR U36598 ( .A(n39554), .B(n39555), .Z(n36708) );
  NOR U36599 ( .A(n39556), .B(n39554), .Z(n39555) );
  XOR U36600 ( .A(n39557), .B(n39558), .Z(n36711) );
  NOR U36601 ( .A(n39559), .B(n39557), .Z(n39558) );
  XOR U36602 ( .A(n39560), .B(n39561), .Z(n36714) );
  NOR U36603 ( .A(n39562), .B(n39560), .Z(n39561) );
  XOR U36604 ( .A(n39563), .B(n39564), .Z(n36717) );
  NOR U36605 ( .A(n39565), .B(n39563), .Z(n39564) );
  XOR U36606 ( .A(n39566), .B(n39567), .Z(n36720) );
  NOR U36607 ( .A(n39568), .B(n39566), .Z(n39567) );
  XOR U36608 ( .A(n39569), .B(n39570), .Z(n36723) );
  NOR U36609 ( .A(n39571), .B(n39569), .Z(n39570) );
  XOR U36610 ( .A(n39572), .B(n39573), .Z(n36726) );
  NOR U36611 ( .A(n39574), .B(n39572), .Z(n39573) );
  XOR U36612 ( .A(n39575), .B(n39576), .Z(n36729) );
  NOR U36613 ( .A(n39577), .B(n39575), .Z(n39576) );
  XOR U36614 ( .A(n39578), .B(n39579), .Z(n36732) );
  NOR U36615 ( .A(n39580), .B(n39578), .Z(n39579) );
  XOR U36616 ( .A(n39581), .B(n39582), .Z(n36735) );
  NOR U36617 ( .A(n39583), .B(n39581), .Z(n39582) );
  XOR U36618 ( .A(n39584), .B(n39585), .Z(n36738) );
  NOR U36619 ( .A(n39586), .B(n39584), .Z(n39585) );
  XOR U36620 ( .A(n39587), .B(n39588), .Z(n36741) );
  NOR U36621 ( .A(n39589), .B(n39587), .Z(n39588) );
  XOR U36622 ( .A(n39590), .B(n39591), .Z(n36744) );
  NOR U36623 ( .A(n39592), .B(n39590), .Z(n39591) );
  XOR U36624 ( .A(n39593), .B(n39594), .Z(n36747) );
  NOR U36625 ( .A(n39595), .B(n39593), .Z(n39594) );
  XOR U36626 ( .A(n39596), .B(n39597), .Z(n36750) );
  NOR U36627 ( .A(n39598), .B(n39596), .Z(n39597) );
  XOR U36628 ( .A(n39599), .B(n39600), .Z(n36753) );
  NOR U36629 ( .A(n39601), .B(n39599), .Z(n39600) );
  XOR U36630 ( .A(n39602), .B(n39603), .Z(n36756) );
  NOR U36631 ( .A(n39604), .B(n39602), .Z(n39603) );
  XOR U36632 ( .A(n39605), .B(n39606), .Z(n36759) );
  NOR U36633 ( .A(n39607), .B(n39605), .Z(n39606) );
  XOR U36634 ( .A(n39608), .B(n39609), .Z(n36762) );
  NOR U36635 ( .A(n39610), .B(n39608), .Z(n39609) );
  XOR U36636 ( .A(n39611), .B(n39612), .Z(n36765) );
  NOR U36637 ( .A(n39613), .B(n39611), .Z(n39612) );
  XOR U36638 ( .A(n39614), .B(n39615), .Z(n36768) );
  NOR U36639 ( .A(n39616), .B(n39614), .Z(n39615) );
  XOR U36640 ( .A(n39617), .B(n39618), .Z(n36771) );
  NOR U36641 ( .A(n39619), .B(n39617), .Z(n39618) );
  XOR U36642 ( .A(n39620), .B(n39621), .Z(n36774) );
  NOR U36643 ( .A(n39622), .B(n39620), .Z(n39621) );
  XOR U36644 ( .A(n39623), .B(n39624), .Z(n36777) );
  NOR U36645 ( .A(n39625), .B(n39623), .Z(n39624) );
  XOR U36646 ( .A(n39626), .B(n39627), .Z(n36780) );
  NOR U36647 ( .A(n39628), .B(n39626), .Z(n39627) );
  XOR U36648 ( .A(n39629), .B(n39630), .Z(n36783) );
  NOR U36649 ( .A(n39631), .B(n39629), .Z(n39630) );
  XOR U36650 ( .A(n39632), .B(n39633), .Z(n36786) );
  NOR U36651 ( .A(n39634), .B(n39632), .Z(n39633) );
  XOR U36652 ( .A(n39635), .B(n39636), .Z(n36789) );
  NOR U36653 ( .A(n39637), .B(n39635), .Z(n39636) );
  XOR U36654 ( .A(n39638), .B(n39639), .Z(n36792) );
  NOR U36655 ( .A(n39640), .B(n39638), .Z(n39639) );
  XOR U36656 ( .A(n39641), .B(n39642), .Z(n36795) );
  NOR U36657 ( .A(n39643), .B(n39641), .Z(n39642) );
  XOR U36658 ( .A(n39644), .B(n39645), .Z(n36798) );
  NOR U36659 ( .A(n39646), .B(n39644), .Z(n39645) );
  XOR U36660 ( .A(n39647), .B(n39648), .Z(n36801) );
  NOR U36661 ( .A(n39649), .B(n39647), .Z(n39648) );
  XOR U36662 ( .A(n39650), .B(n39651), .Z(n36804) );
  NOR U36663 ( .A(n39652), .B(n39650), .Z(n39651) );
  XOR U36664 ( .A(n39653), .B(n39654), .Z(n36807) );
  NOR U36665 ( .A(n39655), .B(n39653), .Z(n39654) );
  XOR U36666 ( .A(n39656), .B(n39657), .Z(n36810) );
  NOR U36667 ( .A(n39658), .B(n39656), .Z(n39657) );
  XOR U36668 ( .A(n39659), .B(n39660), .Z(n36813) );
  NOR U36669 ( .A(n39661), .B(n39659), .Z(n39660) );
  XOR U36670 ( .A(n39662), .B(n39663), .Z(n36816) );
  NOR U36671 ( .A(n39664), .B(n39662), .Z(n39663) );
  XOR U36672 ( .A(n39665), .B(n39666), .Z(n36819) );
  NOR U36673 ( .A(n39667), .B(n39665), .Z(n39666) );
  XOR U36674 ( .A(n39668), .B(n39669), .Z(n36822) );
  NOR U36675 ( .A(n39670), .B(n39668), .Z(n39669) );
  XOR U36676 ( .A(n39671), .B(n39672), .Z(n36825) );
  NOR U36677 ( .A(n39673), .B(n39671), .Z(n39672) );
  XOR U36678 ( .A(n39674), .B(n39675), .Z(n36828) );
  NOR U36679 ( .A(n39676), .B(n39674), .Z(n39675) );
  XOR U36680 ( .A(n39677), .B(n39678), .Z(n36831) );
  NOR U36681 ( .A(n39679), .B(n39677), .Z(n39678) );
  XOR U36682 ( .A(n39680), .B(n39681), .Z(n36834) );
  NOR U36683 ( .A(n39682), .B(n39680), .Z(n39681) );
  XOR U36684 ( .A(n39683), .B(n39684), .Z(n36837) );
  NOR U36685 ( .A(n39685), .B(n39683), .Z(n39684) );
  XOR U36686 ( .A(n39686), .B(n39687), .Z(n36840) );
  NOR U36687 ( .A(n39688), .B(n39686), .Z(n39687) );
  XOR U36688 ( .A(n39689), .B(n39690), .Z(n36843) );
  NOR U36689 ( .A(n39691), .B(n39689), .Z(n39690) );
  XOR U36690 ( .A(n39692), .B(n39693), .Z(n36846) );
  NOR U36691 ( .A(n39694), .B(n39692), .Z(n39693) );
  XOR U36692 ( .A(n39695), .B(n39696), .Z(n36849) );
  NOR U36693 ( .A(n39697), .B(n39695), .Z(n39696) );
  XOR U36694 ( .A(n39698), .B(n39699), .Z(n36852) );
  NOR U36695 ( .A(n39700), .B(n39698), .Z(n39699) );
  XOR U36696 ( .A(n39701), .B(n39702), .Z(n36855) );
  NOR U36697 ( .A(n39703), .B(n39701), .Z(n39702) );
  XOR U36698 ( .A(n39704), .B(n39705), .Z(n36858) );
  NOR U36699 ( .A(n39706), .B(n39704), .Z(n39705) );
  XOR U36700 ( .A(n39707), .B(n39708), .Z(n36861) );
  NOR U36701 ( .A(n39709), .B(n39707), .Z(n39708) );
  XOR U36702 ( .A(n39710), .B(n39711), .Z(n36864) );
  NOR U36703 ( .A(n39712), .B(n39710), .Z(n39711) );
  XOR U36704 ( .A(n39713), .B(n39714), .Z(n36867) );
  NOR U36705 ( .A(n39715), .B(n39713), .Z(n39714) );
  XOR U36706 ( .A(n39716), .B(n39717), .Z(n36870) );
  NOR U36707 ( .A(n39718), .B(n39716), .Z(n39717) );
  XOR U36708 ( .A(n39719), .B(n39720), .Z(n36873) );
  NOR U36709 ( .A(n39721), .B(n39719), .Z(n39720) );
  XOR U36710 ( .A(n39722), .B(n39723), .Z(n36876) );
  NOR U36711 ( .A(n39724), .B(n39722), .Z(n39723) );
  XOR U36712 ( .A(n39725), .B(n39726), .Z(n36879) );
  NOR U36713 ( .A(n39727), .B(n39725), .Z(n39726) );
  XOR U36714 ( .A(n39728), .B(n39729), .Z(n36882) );
  NOR U36715 ( .A(n39730), .B(n39728), .Z(n39729) );
  XOR U36716 ( .A(n39731), .B(n39732), .Z(n36885) );
  NOR U36717 ( .A(n39733), .B(n39731), .Z(n39732) );
  XOR U36718 ( .A(n39734), .B(n39735), .Z(n36888) );
  NOR U36719 ( .A(n39736), .B(n39734), .Z(n39735) );
  XOR U36720 ( .A(n39737), .B(n39738), .Z(n36891) );
  NOR U36721 ( .A(n39739), .B(n39737), .Z(n39738) );
  XOR U36722 ( .A(n39740), .B(n39741), .Z(n36894) );
  NOR U36723 ( .A(n39742), .B(n39740), .Z(n39741) );
  XOR U36724 ( .A(n39743), .B(n39744), .Z(n36897) );
  NOR U36725 ( .A(n39745), .B(n39743), .Z(n39744) );
  XOR U36726 ( .A(n39746), .B(n39747), .Z(n36900) );
  NOR U36727 ( .A(n39748), .B(n39746), .Z(n39747) );
  XOR U36728 ( .A(n39749), .B(n39750), .Z(n36903) );
  NOR U36729 ( .A(n39751), .B(n39749), .Z(n39750) );
  XOR U36730 ( .A(n39752), .B(n39753), .Z(n36906) );
  NOR U36731 ( .A(n39754), .B(n39752), .Z(n39753) );
  XOR U36732 ( .A(n39755), .B(n39756), .Z(n36909) );
  NOR U36733 ( .A(n39757), .B(n39755), .Z(n39756) );
  XOR U36734 ( .A(n39758), .B(n39759), .Z(n36912) );
  NOR U36735 ( .A(n39760), .B(n39758), .Z(n39759) );
  XOR U36736 ( .A(n39761), .B(n39762), .Z(n36915) );
  NOR U36737 ( .A(n39763), .B(n39761), .Z(n39762) );
  XOR U36738 ( .A(n39764), .B(n39765), .Z(n36918) );
  NOR U36739 ( .A(n39766), .B(n39764), .Z(n39765) );
  XOR U36740 ( .A(n39767), .B(n39768), .Z(n36921) );
  NOR U36741 ( .A(n39769), .B(n39767), .Z(n39768) );
  XOR U36742 ( .A(n39770), .B(n39771), .Z(n36924) );
  NOR U36743 ( .A(n39772), .B(n39770), .Z(n39771) );
  XOR U36744 ( .A(n39773), .B(n39774), .Z(n36927) );
  NOR U36745 ( .A(n39775), .B(n39773), .Z(n39774) );
  XOR U36746 ( .A(n39776), .B(n39777), .Z(n36930) );
  NOR U36747 ( .A(n39778), .B(n39776), .Z(n39777) );
  XOR U36748 ( .A(n39779), .B(n39780), .Z(n36933) );
  NOR U36749 ( .A(n39781), .B(n39779), .Z(n39780) );
  XOR U36750 ( .A(n39782), .B(n39783), .Z(n36936) );
  NOR U36751 ( .A(n39784), .B(n39782), .Z(n39783) );
  XOR U36752 ( .A(n39785), .B(n39786), .Z(n36939) );
  NOR U36753 ( .A(n39787), .B(n39785), .Z(n39786) );
  XOR U36754 ( .A(n39788), .B(n39789), .Z(n36942) );
  NOR U36755 ( .A(n39790), .B(n39788), .Z(n39789) );
  XOR U36756 ( .A(n39791), .B(n39792), .Z(n36945) );
  NOR U36757 ( .A(n39793), .B(n39791), .Z(n39792) );
  XOR U36758 ( .A(n39794), .B(n39795), .Z(n36948) );
  NOR U36759 ( .A(n39796), .B(n39794), .Z(n39795) );
  XOR U36760 ( .A(n39797), .B(n39798), .Z(n36951) );
  NOR U36761 ( .A(n39799), .B(n39797), .Z(n39798) );
  XOR U36762 ( .A(n39800), .B(n39801), .Z(n36954) );
  NOR U36763 ( .A(n39802), .B(n39800), .Z(n39801) );
  XOR U36764 ( .A(n39803), .B(n39804), .Z(n36957) );
  NOR U36765 ( .A(n39805), .B(n39803), .Z(n39804) );
  XOR U36766 ( .A(n39806), .B(n39807), .Z(n36960) );
  NOR U36767 ( .A(n121), .B(n39808), .Z(n39807) );
  XOR U36768 ( .A(n39809), .B(n39810), .Z(n36963) );
  AND U36769 ( .A(n39811), .B(n39812), .Z(n39810) );
  XOR U36770 ( .A(n39809), .B(n124), .Z(n39812) );
  XNOR U36771 ( .A(n38386), .B(n38385), .Z(n124) );
  XNOR U36772 ( .A(n38383), .B(n38382), .Z(n38385) );
  XNOR U36773 ( .A(n38380), .B(n38379), .Z(n38382) );
  XNOR U36774 ( .A(n38377), .B(n38376), .Z(n38379) );
  XNOR U36775 ( .A(n38374), .B(n38373), .Z(n38376) );
  XNOR U36776 ( .A(n38371), .B(n38370), .Z(n38373) );
  XNOR U36777 ( .A(n38368), .B(n38367), .Z(n38370) );
  XNOR U36778 ( .A(n38365), .B(n38364), .Z(n38367) );
  XNOR U36779 ( .A(n38362), .B(n38361), .Z(n38364) );
  XNOR U36780 ( .A(n38359), .B(n38358), .Z(n38361) );
  XNOR U36781 ( .A(n38356), .B(n38355), .Z(n38358) );
  XNOR U36782 ( .A(n38353), .B(n38352), .Z(n38355) );
  XNOR U36783 ( .A(n38350), .B(n38349), .Z(n38352) );
  XNOR U36784 ( .A(n38347), .B(n38346), .Z(n38349) );
  XNOR U36785 ( .A(n38344), .B(n38343), .Z(n38346) );
  XNOR U36786 ( .A(n38341), .B(n38340), .Z(n38343) );
  XNOR U36787 ( .A(n38338), .B(n38337), .Z(n38340) );
  XNOR U36788 ( .A(n38335), .B(n38334), .Z(n38337) );
  XNOR U36789 ( .A(n38332), .B(n38331), .Z(n38334) );
  XNOR U36790 ( .A(n38329), .B(n38328), .Z(n38331) );
  XNOR U36791 ( .A(n38326), .B(n38325), .Z(n38328) );
  XNOR U36792 ( .A(n38323), .B(n38322), .Z(n38325) );
  XNOR U36793 ( .A(n38320), .B(n38319), .Z(n38322) );
  XNOR U36794 ( .A(n38317), .B(n38316), .Z(n38319) );
  XNOR U36795 ( .A(n38314), .B(n38313), .Z(n38316) );
  XNOR U36796 ( .A(n38311), .B(n38310), .Z(n38313) );
  XNOR U36797 ( .A(n38308), .B(n38307), .Z(n38310) );
  XNOR U36798 ( .A(n38305), .B(n38304), .Z(n38307) );
  XNOR U36799 ( .A(n38302), .B(n38301), .Z(n38304) );
  XNOR U36800 ( .A(n38299), .B(n38298), .Z(n38301) );
  XNOR U36801 ( .A(n38296), .B(n38295), .Z(n38298) );
  XNOR U36802 ( .A(n38293), .B(n38292), .Z(n38295) );
  XNOR U36803 ( .A(n38290), .B(n38289), .Z(n38292) );
  XNOR U36804 ( .A(n38287), .B(n38286), .Z(n38289) );
  XNOR U36805 ( .A(n38284), .B(n38283), .Z(n38286) );
  XNOR U36806 ( .A(n38281), .B(n38280), .Z(n38283) );
  XNOR U36807 ( .A(n38278), .B(n38277), .Z(n38280) );
  XNOR U36808 ( .A(n38275), .B(n38274), .Z(n38277) );
  XNOR U36809 ( .A(n38272), .B(n38271), .Z(n38274) );
  XNOR U36810 ( .A(n38269), .B(n38268), .Z(n38271) );
  XNOR U36811 ( .A(n38266), .B(n38265), .Z(n38268) );
  XNOR U36812 ( .A(n38263), .B(n38262), .Z(n38265) );
  XNOR U36813 ( .A(n38260), .B(n38259), .Z(n38262) );
  XNOR U36814 ( .A(n38257), .B(n38256), .Z(n38259) );
  XNOR U36815 ( .A(n38254), .B(n38253), .Z(n38256) );
  XNOR U36816 ( .A(n38251), .B(n38250), .Z(n38253) );
  XNOR U36817 ( .A(n38248), .B(n38247), .Z(n38250) );
  XNOR U36818 ( .A(n38245), .B(n38244), .Z(n38247) );
  XNOR U36819 ( .A(n38242), .B(n38241), .Z(n38244) );
  XNOR U36820 ( .A(n38239), .B(n38238), .Z(n38241) );
  XNOR U36821 ( .A(n38236), .B(n38235), .Z(n38238) );
  XNOR U36822 ( .A(n38233), .B(n38232), .Z(n38235) );
  XNOR U36823 ( .A(n38230), .B(n38229), .Z(n38232) );
  XNOR U36824 ( .A(n38227), .B(n38226), .Z(n38229) );
  XNOR U36825 ( .A(n38224), .B(n38223), .Z(n38226) );
  XNOR U36826 ( .A(n38221), .B(n38220), .Z(n38223) );
  XNOR U36827 ( .A(n38218), .B(n38217), .Z(n38220) );
  XNOR U36828 ( .A(n38215), .B(n38214), .Z(n38217) );
  XNOR U36829 ( .A(n38212), .B(n38211), .Z(n38214) );
  XNOR U36830 ( .A(n38209), .B(n38208), .Z(n38211) );
  XNOR U36831 ( .A(n38206), .B(n38205), .Z(n38208) );
  XNOR U36832 ( .A(n38203), .B(n38202), .Z(n38205) );
  XNOR U36833 ( .A(n38200), .B(n38199), .Z(n38202) );
  XNOR U36834 ( .A(n38197), .B(n38196), .Z(n38199) );
  XNOR U36835 ( .A(n38194), .B(n38193), .Z(n38196) );
  XNOR U36836 ( .A(n38191), .B(n38190), .Z(n38193) );
  XNOR U36837 ( .A(n38188), .B(n38187), .Z(n38190) );
  XNOR U36838 ( .A(n38185), .B(n38184), .Z(n38187) );
  XNOR U36839 ( .A(n38182), .B(n38181), .Z(n38184) );
  XNOR U36840 ( .A(n38179), .B(n38178), .Z(n38181) );
  XNOR U36841 ( .A(n38176), .B(n38175), .Z(n38178) );
  XNOR U36842 ( .A(n38173), .B(n38172), .Z(n38175) );
  XNOR U36843 ( .A(n38170), .B(n38169), .Z(n38172) );
  XNOR U36844 ( .A(n38167), .B(n38166), .Z(n38169) );
  XNOR U36845 ( .A(n38164), .B(n38163), .Z(n38166) );
  XNOR U36846 ( .A(n38161), .B(n38160), .Z(n38163) );
  XNOR U36847 ( .A(n38158), .B(n38157), .Z(n38160) );
  XNOR U36848 ( .A(n38155), .B(n38154), .Z(n38157) );
  XNOR U36849 ( .A(n38152), .B(n38151), .Z(n38154) );
  XNOR U36850 ( .A(n38149), .B(n38148), .Z(n38151) );
  XNOR U36851 ( .A(n38146), .B(n38145), .Z(n38148) );
  XNOR U36852 ( .A(n38143), .B(n38142), .Z(n38145) );
  XNOR U36853 ( .A(n38140), .B(n38139), .Z(n38142) );
  XNOR U36854 ( .A(n38137), .B(n38136), .Z(n38139) );
  XNOR U36855 ( .A(n38134), .B(n38133), .Z(n38136) );
  XNOR U36856 ( .A(n38131), .B(n38130), .Z(n38133) );
  XNOR U36857 ( .A(n38128), .B(n38127), .Z(n38130) );
  XNOR U36858 ( .A(n38125), .B(n38124), .Z(n38127) );
  XNOR U36859 ( .A(n38122), .B(n38121), .Z(n38124) );
  XNOR U36860 ( .A(n38119), .B(n38118), .Z(n38121) );
  XNOR U36861 ( .A(n38116), .B(n38115), .Z(n38118) );
  XNOR U36862 ( .A(n38113), .B(n38112), .Z(n38115) );
  XNOR U36863 ( .A(n38110), .B(n38109), .Z(n38112) );
  XNOR U36864 ( .A(n38107), .B(n38106), .Z(n38109) );
  XNOR U36865 ( .A(n38104), .B(n38103), .Z(n38106) );
  XNOR U36866 ( .A(n38101), .B(n38100), .Z(n38103) );
  XNOR U36867 ( .A(n38098), .B(n38097), .Z(n38100) );
  XNOR U36868 ( .A(n38095), .B(n38094), .Z(n38097) );
  XNOR U36869 ( .A(n38092), .B(n38091), .Z(n38094) );
  XNOR U36870 ( .A(n38089), .B(n38088), .Z(n38091) );
  XNOR U36871 ( .A(n38086), .B(n38085), .Z(n38088) );
  XNOR U36872 ( .A(n38083), .B(n38082), .Z(n38085) );
  XNOR U36873 ( .A(n38080), .B(n38079), .Z(n38082) );
  XNOR U36874 ( .A(n38077), .B(n38076), .Z(n38079) );
  XNOR U36875 ( .A(n38074), .B(n38073), .Z(n38076) );
  XNOR U36876 ( .A(n38071), .B(n38070), .Z(n38073) );
  XNOR U36877 ( .A(n38068), .B(n38067), .Z(n38070) );
  XNOR U36878 ( .A(n38065), .B(n38064), .Z(n38067) );
  XNOR U36879 ( .A(n38062), .B(n38061), .Z(n38064) );
  XNOR U36880 ( .A(n38059), .B(n38058), .Z(n38061) );
  XNOR U36881 ( .A(n38056), .B(n38055), .Z(n38058) );
  XNOR U36882 ( .A(n38053), .B(n38052), .Z(n38055) );
  XNOR U36883 ( .A(n38050), .B(n38049), .Z(n38052) );
  XNOR U36884 ( .A(n38047), .B(n38046), .Z(n38049) );
  XNOR U36885 ( .A(n38044), .B(n38043), .Z(n38046) );
  XNOR U36886 ( .A(n38041), .B(n38040), .Z(n38043) );
  XNOR U36887 ( .A(n38038), .B(n38037), .Z(n38040) );
  XNOR U36888 ( .A(n38035), .B(n38034), .Z(n38037) );
  XNOR U36889 ( .A(n38032), .B(n38031), .Z(n38034) );
  XNOR U36890 ( .A(n38029), .B(n38028), .Z(n38031) );
  XNOR U36891 ( .A(n38026), .B(n38025), .Z(n38028) );
  XNOR U36892 ( .A(n38023), .B(n38022), .Z(n38025) );
  XNOR U36893 ( .A(n38020), .B(n38019), .Z(n38022) );
  XNOR U36894 ( .A(n38017), .B(n38016), .Z(n38019) );
  XNOR U36895 ( .A(n38014), .B(n38013), .Z(n38016) );
  XNOR U36896 ( .A(n38011), .B(n38010), .Z(n38013) );
  XNOR U36897 ( .A(n38008), .B(n38007), .Z(n38010) );
  XNOR U36898 ( .A(n38005), .B(n38004), .Z(n38007) );
  XNOR U36899 ( .A(n38002), .B(n38001), .Z(n38004) );
  XNOR U36900 ( .A(n37999), .B(n37998), .Z(n38001) );
  XNOR U36901 ( .A(n37996), .B(n37995), .Z(n37998) );
  XNOR U36902 ( .A(n37993), .B(n37992), .Z(n37995) );
  XNOR U36903 ( .A(n37990), .B(n37989), .Z(n37992) );
  XNOR U36904 ( .A(n37987), .B(n37986), .Z(n37989) );
  XNOR U36905 ( .A(n37984), .B(n37983), .Z(n37986) );
  XNOR U36906 ( .A(n37981), .B(n37980), .Z(n37983) );
  XNOR U36907 ( .A(n37978), .B(n37977), .Z(n37980) );
  XNOR U36908 ( .A(n37975), .B(n37974), .Z(n37977) );
  XNOR U36909 ( .A(n37972), .B(n37971), .Z(n37974) );
  XNOR U36910 ( .A(n37969), .B(n37968), .Z(n37971) );
  XNOR U36911 ( .A(n37966), .B(n37965), .Z(n37968) );
  XNOR U36912 ( .A(n37963), .B(n37962), .Z(n37965) );
  XNOR U36913 ( .A(n37960), .B(n37959), .Z(n37962) );
  XNOR U36914 ( .A(n37957), .B(n37956), .Z(n37959) );
  XNOR U36915 ( .A(n37954), .B(n37953), .Z(n37956) );
  XNOR U36916 ( .A(n37951), .B(n37950), .Z(n37953) );
  XNOR U36917 ( .A(n37948), .B(n37947), .Z(n37950) );
  XNOR U36918 ( .A(n37945), .B(n37944), .Z(n37947) );
  XNOR U36919 ( .A(n37942), .B(n37941), .Z(n37944) );
  XNOR U36920 ( .A(n37939), .B(n37938), .Z(n37941) );
  XNOR U36921 ( .A(n37936), .B(n37935), .Z(n37938) );
  XNOR U36922 ( .A(n37933), .B(n37932), .Z(n37935) );
  XNOR U36923 ( .A(n37930), .B(n37929), .Z(n37932) );
  XNOR U36924 ( .A(n37927), .B(n37926), .Z(n37929) );
  XNOR U36925 ( .A(n37924), .B(n37923), .Z(n37926) );
  XNOR U36926 ( .A(n37921), .B(n37920), .Z(n37923) );
  XNOR U36927 ( .A(n37918), .B(n37917), .Z(n37920) );
  XNOR U36928 ( .A(n37915), .B(n37914), .Z(n37917) );
  XNOR U36929 ( .A(n37912), .B(n37911), .Z(n37914) );
  XNOR U36930 ( .A(n37909), .B(n37908), .Z(n37911) );
  XNOR U36931 ( .A(n37906), .B(n37905), .Z(n37908) );
  XNOR U36932 ( .A(n37903), .B(n37902), .Z(n37905) );
  XNOR U36933 ( .A(n37900), .B(n37899), .Z(n37902) );
  XNOR U36934 ( .A(n37897), .B(n37896), .Z(n37899) );
  XNOR U36935 ( .A(n37894), .B(n37893), .Z(n37896) );
  XNOR U36936 ( .A(n37891), .B(n37890), .Z(n37893) );
  XNOR U36937 ( .A(n37888), .B(n37887), .Z(n37890) );
  XNOR U36938 ( .A(n37885), .B(n37884), .Z(n37887) );
  XNOR U36939 ( .A(n37882), .B(n37881), .Z(n37884) );
  XNOR U36940 ( .A(n37879), .B(n37878), .Z(n37881) );
  XNOR U36941 ( .A(n37876), .B(n37875), .Z(n37878) );
  XNOR U36942 ( .A(n37873), .B(n37872), .Z(n37875) );
  XNOR U36943 ( .A(n37870), .B(n37869), .Z(n37872) );
  XNOR U36944 ( .A(n37867), .B(n37866), .Z(n37869) );
  XNOR U36945 ( .A(n37864), .B(n37863), .Z(n37866) );
  XNOR U36946 ( .A(n37861), .B(n37860), .Z(n37863) );
  XNOR U36947 ( .A(n37858), .B(n37857), .Z(n37860) );
  XNOR U36948 ( .A(n37855), .B(n37854), .Z(n37857) );
  XNOR U36949 ( .A(n37852), .B(n37851), .Z(n37854) );
  XNOR U36950 ( .A(n37849), .B(n37848), .Z(n37851) );
  XNOR U36951 ( .A(n37846), .B(n37845), .Z(n37848) );
  XNOR U36952 ( .A(n37843), .B(n37842), .Z(n37845) );
  XNOR U36953 ( .A(n37840), .B(n37839), .Z(n37842) );
  XNOR U36954 ( .A(n37837), .B(n37836), .Z(n37839) );
  XNOR U36955 ( .A(n37834), .B(n37833), .Z(n37836) );
  XNOR U36956 ( .A(n37831), .B(n37830), .Z(n37833) );
  XNOR U36957 ( .A(n37828), .B(n37827), .Z(n37830) );
  XNOR U36958 ( .A(n37825), .B(n37824), .Z(n37827) );
  XNOR U36959 ( .A(n37822), .B(n37821), .Z(n37824) );
  XNOR U36960 ( .A(n37819), .B(n37818), .Z(n37821) );
  XNOR U36961 ( .A(n37816), .B(n37815), .Z(n37818) );
  XNOR U36962 ( .A(n37813), .B(n37812), .Z(n37815) );
  XNOR U36963 ( .A(n37810), .B(n37809), .Z(n37812) );
  XNOR U36964 ( .A(n37807), .B(n37806), .Z(n37809) );
  XNOR U36965 ( .A(n37804), .B(n37803), .Z(n37806) );
  XNOR U36966 ( .A(n37801), .B(n37800), .Z(n37803) );
  XNOR U36967 ( .A(n37798), .B(n37797), .Z(n37800) );
  XNOR U36968 ( .A(n37795), .B(n37794), .Z(n37797) );
  XNOR U36969 ( .A(n37792), .B(n37791), .Z(n37794) );
  XNOR U36970 ( .A(n37789), .B(n37788), .Z(n37791) );
  XNOR U36971 ( .A(n37786), .B(n37785), .Z(n37788) );
  XNOR U36972 ( .A(n37783), .B(n37782), .Z(n37785) );
  XNOR U36973 ( .A(n37780), .B(n37779), .Z(n37782) );
  XNOR U36974 ( .A(n37777), .B(n37776), .Z(n37779) );
  XNOR U36975 ( .A(n37774), .B(n37773), .Z(n37776) );
  XNOR U36976 ( .A(n37771), .B(n37770), .Z(n37773) );
  XNOR U36977 ( .A(n37768), .B(n37767), .Z(n37770) );
  XNOR U36978 ( .A(n37765), .B(n37764), .Z(n37767) );
  XNOR U36979 ( .A(n37762), .B(n37761), .Z(n37764) );
  XNOR U36980 ( .A(n37759), .B(n37758), .Z(n37761) );
  XNOR U36981 ( .A(n37756), .B(n37755), .Z(n37758) );
  XNOR U36982 ( .A(n37753), .B(n37752), .Z(n37755) );
  XNOR U36983 ( .A(n37750), .B(n37749), .Z(n37752) );
  XNOR U36984 ( .A(n37747), .B(n37746), .Z(n37749) );
  XNOR U36985 ( .A(n37744), .B(n37743), .Z(n37746) );
  XNOR U36986 ( .A(n37741), .B(n37740), .Z(n37743) );
  XNOR U36987 ( .A(n37738), .B(n37737), .Z(n37740) );
  XNOR U36988 ( .A(n37735), .B(n37734), .Z(n37737) );
  XNOR U36989 ( .A(n37732), .B(n37731), .Z(n37734) );
  XNOR U36990 ( .A(n37729), .B(n37728), .Z(n37731) );
  XNOR U36991 ( .A(n37726), .B(n37725), .Z(n37728) );
  XNOR U36992 ( .A(n37723), .B(n37722), .Z(n37725) );
  XNOR U36993 ( .A(n37720), .B(n37719), .Z(n37722) );
  XNOR U36994 ( .A(n37717), .B(n37716), .Z(n37719) );
  XNOR U36995 ( .A(n37714), .B(n37713), .Z(n37716) );
  XNOR U36996 ( .A(n37711), .B(n37710), .Z(n37713) );
  XNOR U36997 ( .A(n37708), .B(n37707), .Z(n37710) );
  XNOR U36998 ( .A(n37705), .B(n37704), .Z(n37707) );
  XNOR U36999 ( .A(n37702), .B(n37701), .Z(n37704) );
  XNOR U37000 ( .A(n37699), .B(n37698), .Z(n37701) );
  XNOR U37001 ( .A(n37696), .B(n37695), .Z(n37698) );
  XNOR U37002 ( .A(n37693), .B(n37692), .Z(n37695) );
  XNOR U37003 ( .A(n37690), .B(n37689), .Z(n37692) );
  XNOR U37004 ( .A(n37687), .B(n37686), .Z(n37689) );
  XNOR U37005 ( .A(n37684), .B(n37683), .Z(n37686) );
  XNOR U37006 ( .A(n37681), .B(n37680), .Z(n37683) );
  XNOR U37007 ( .A(n37678), .B(n37677), .Z(n37680) );
  XNOR U37008 ( .A(n37675), .B(n37674), .Z(n37677) );
  XNOR U37009 ( .A(n37672), .B(n37671), .Z(n37674) );
  XNOR U37010 ( .A(n37669), .B(n37668), .Z(n37671) );
  XNOR U37011 ( .A(n37666), .B(n37665), .Z(n37668) );
  XNOR U37012 ( .A(n37663), .B(n37662), .Z(n37665) );
  XNOR U37013 ( .A(n37660), .B(n37659), .Z(n37662) );
  XNOR U37014 ( .A(n37657), .B(n37656), .Z(n37659) );
  XNOR U37015 ( .A(n37654), .B(n37653), .Z(n37656) );
  XNOR U37016 ( .A(n37651), .B(n37650), .Z(n37653) );
  XNOR U37017 ( .A(n37648), .B(n37647), .Z(n37650) );
  XNOR U37018 ( .A(n37645), .B(n37644), .Z(n37647) );
  XNOR U37019 ( .A(n37642), .B(n37641), .Z(n37644) );
  XNOR U37020 ( .A(n37639), .B(n37638), .Z(n37641) );
  XNOR U37021 ( .A(n37636), .B(n37635), .Z(n37638) );
  XNOR U37022 ( .A(n37633), .B(n37632), .Z(n37635) );
  XNOR U37023 ( .A(n37630), .B(n37629), .Z(n37632) );
  XNOR U37024 ( .A(n37627), .B(n37626), .Z(n37629) );
  XNOR U37025 ( .A(n37624), .B(n37623), .Z(n37626) );
  XNOR U37026 ( .A(n37621), .B(n37620), .Z(n37623) );
  XNOR U37027 ( .A(n37618), .B(n37617), .Z(n37620) );
  XNOR U37028 ( .A(n37615), .B(n37614), .Z(n37617) );
  XNOR U37029 ( .A(n37612), .B(n37611), .Z(n37614) );
  XNOR U37030 ( .A(n37609), .B(n37608), .Z(n37611) );
  XNOR U37031 ( .A(n37606), .B(n37605), .Z(n37608) );
  XNOR U37032 ( .A(n37603), .B(n37602), .Z(n37605) );
  XNOR U37033 ( .A(n37600), .B(n37599), .Z(n37602) );
  XNOR U37034 ( .A(n37597), .B(n37596), .Z(n37599) );
  XNOR U37035 ( .A(n37594), .B(n37593), .Z(n37596) );
  XNOR U37036 ( .A(n37591), .B(n37590), .Z(n37593) );
  XNOR U37037 ( .A(n37588), .B(n37587), .Z(n37590) );
  XNOR U37038 ( .A(n37585), .B(n37584), .Z(n37587) );
  XNOR U37039 ( .A(n37582), .B(n37581), .Z(n37584) );
  XNOR U37040 ( .A(n37579), .B(n37578), .Z(n37581) );
  XNOR U37041 ( .A(n37576), .B(n37575), .Z(n37578) );
  XNOR U37042 ( .A(n37573), .B(n37572), .Z(n37575) );
  XNOR U37043 ( .A(n37570), .B(n37569), .Z(n37572) );
  XNOR U37044 ( .A(n37567), .B(n37566), .Z(n37569) );
  XNOR U37045 ( .A(n37564), .B(n37563), .Z(n37566) );
  XNOR U37046 ( .A(n37561), .B(n37560), .Z(n37563) );
  XNOR U37047 ( .A(n37558), .B(n37557), .Z(n37560) );
  XNOR U37048 ( .A(n37555), .B(n37554), .Z(n37557) );
  XNOR U37049 ( .A(n37552), .B(n37551), .Z(n37554) );
  XNOR U37050 ( .A(n37549), .B(n37548), .Z(n37551) );
  XNOR U37051 ( .A(n37546), .B(n37545), .Z(n37548) );
  XNOR U37052 ( .A(n37543), .B(n37542), .Z(n37545) );
  XNOR U37053 ( .A(n37540), .B(n37539), .Z(n37542) );
  XNOR U37054 ( .A(n37537), .B(n37536), .Z(n37539) );
  XNOR U37055 ( .A(n37534), .B(n37533), .Z(n37536) );
  XNOR U37056 ( .A(n37531), .B(n37530), .Z(n37533) );
  XNOR U37057 ( .A(n37528), .B(n37527), .Z(n37530) );
  XNOR U37058 ( .A(n37525), .B(n37524), .Z(n37527) );
  XNOR U37059 ( .A(n37522), .B(n37521), .Z(n37524) );
  XNOR U37060 ( .A(n37519), .B(n37518), .Z(n37521) );
  XNOR U37061 ( .A(n37516), .B(n37515), .Z(n37518) );
  XNOR U37062 ( .A(n37513), .B(n37512), .Z(n37515) );
  XNOR U37063 ( .A(n37510), .B(n37509), .Z(n37512) );
  XNOR U37064 ( .A(n37507), .B(n37506), .Z(n37509) );
  XNOR U37065 ( .A(n37504), .B(n37503), .Z(n37506) );
  XNOR U37066 ( .A(n37501), .B(n37500), .Z(n37503) );
  XNOR U37067 ( .A(n37498), .B(n37497), .Z(n37500) );
  XNOR U37068 ( .A(n37495), .B(n37494), .Z(n37497) );
  XNOR U37069 ( .A(n37492), .B(n37491), .Z(n37494) );
  XNOR U37070 ( .A(n37489), .B(n37488), .Z(n37491) );
  XNOR U37071 ( .A(n37486), .B(n37485), .Z(n37488) );
  XNOR U37072 ( .A(n37483), .B(n37482), .Z(n37485) );
  XNOR U37073 ( .A(n37480), .B(n37479), .Z(n37482) );
  XNOR U37074 ( .A(n37477), .B(n37476), .Z(n37479) );
  XNOR U37075 ( .A(n37474), .B(n37473), .Z(n37476) );
  XNOR U37076 ( .A(n37471), .B(n37470), .Z(n37473) );
  XNOR U37077 ( .A(n37468), .B(n37467), .Z(n37470) );
  XNOR U37078 ( .A(n37465), .B(n37464), .Z(n37467) );
  XNOR U37079 ( .A(n37462), .B(n37461), .Z(n37464) );
  XNOR U37080 ( .A(n37459), .B(n37458), .Z(n37461) );
  XNOR U37081 ( .A(n37456), .B(n37455), .Z(n37458) );
  XNOR U37082 ( .A(n37453), .B(n37452), .Z(n37455) );
  XNOR U37083 ( .A(n37450), .B(n37449), .Z(n37452) );
  XNOR U37084 ( .A(n37447), .B(n37446), .Z(n37449) );
  XNOR U37085 ( .A(n37444), .B(n37443), .Z(n37446) );
  XNOR U37086 ( .A(n37441), .B(n37440), .Z(n37443) );
  XNOR U37087 ( .A(n37438), .B(n37437), .Z(n37440) );
  XNOR U37088 ( .A(n37435), .B(n37434), .Z(n37437) );
  XNOR U37089 ( .A(n37432), .B(n37431), .Z(n37434) );
  XNOR U37090 ( .A(n37429), .B(n37428), .Z(n37431) );
  XNOR U37091 ( .A(n37426), .B(n37425), .Z(n37428) );
  XNOR U37092 ( .A(n37423), .B(n37422), .Z(n37425) );
  XNOR U37093 ( .A(n37420), .B(n37419), .Z(n37422) );
  XNOR U37094 ( .A(n37417), .B(n37416), .Z(n37419) );
  XNOR U37095 ( .A(n37414), .B(n37413), .Z(n37416) );
  XNOR U37096 ( .A(n37411), .B(n37410), .Z(n37413) );
  XNOR U37097 ( .A(n37408), .B(n37407), .Z(n37410) );
  XNOR U37098 ( .A(n37405), .B(n37404), .Z(n37407) );
  XNOR U37099 ( .A(n37402), .B(n37401), .Z(n37404) );
  XNOR U37100 ( .A(n37399), .B(n37398), .Z(n37401) );
  XNOR U37101 ( .A(n37396), .B(n37395), .Z(n37398) );
  XNOR U37102 ( .A(n37393), .B(n37392), .Z(n37395) );
  XNOR U37103 ( .A(n37390), .B(n37389), .Z(n37392) );
  XNOR U37104 ( .A(n37387), .B(n37386), .Z(n37389) );
  XNOR U37105 ( .A(n37384), .B(n37383), .Z(n37386) );
  XNOR U37106 ( .A(n37381), .B(n37380), .Z(n37383) );
  XNOR U37107 ( .A(n37378), .B(n37377), .Z(n37380) );
  XNOR U37108 ( .A(n37375), .B(n37374), .Z(n37377) );
  XNOR U37109 ( .A(n37372), .B(n37371), .Z(n37374) );
  XNOR U37110 ( .A(n37369), .B(n37368), .Z(n37371) );
  XNOR U37111 ( .A(n37366), .B(n37365), .Z(n37368) );
  XNOR U37112 ( .A(n37363), .B(n37362), .Z(n37365) );
  XNOR U37113 ( .A(n37360), .B(n37359), .Z(n37362) );
  XNOR U37114 ( .A(n37357), .B(n37356), .Z(n37359) );
  XNOR U37115 ( .A(n37354), .B(n37353), .Z(n37356) );
  XNOR U37116 ( .A(n37351), .B(n37350), .Z(n37353) );
  XNOR U37117 ( .A(n37348), .B(n37347), .Z(n37350) );
  XNOR U37118 ( .A(n37345), .B(n37344), .Z(n37347) );
  XNOR U37119 ( .A(n37342), .B(n37341), .Z(n37344) );
  XNOR U37120 ( .A(n37339), .B(n37338), .Z(n37341) );
  XNOR U37121 ( .A(n37336), .B(n37335), .Z(n37338) );
  XNOR U37122 ( .A(n37333), .B(n37332), .Z(n37335) );
  XNOR U37123 ( .A(n37330), .B(n37329), .Z(n37332) );
  XNOR U37124 ( .A(n37327), .B(n37326), .Z(n37329) );
  XNOR U37125 ( .A(n37324), .B(n37323), .Z(n37326) );
  XNOR U37126 ( .A(n37321), .B(n37320), .Z(n37323) );
  XNOR U37127 ( .A(n37318), .B(n37317), .Z(n37320) );
  XNOR U37128 ( .A(n37315), .B(n37314), .Z(n37317) );
  XNOR U37129 ( .A(n37312), .B(n37311), .Z(n37314) );
  XNOR U37130 ( .A(n37309), .B(n37308), .Z(n37311) );
  XNOR U37131 ( .A(n37306), .B(n37305), .Z(n37308) );
  XNOR U37132 ( .A(n37303), .B(n37302), .Z(n37305) );
  XNOR U37133 ( .A(n37300), .B(n37299), .Z(n37302) );
  XNOR U37134 ( .A(n37297), .B(n37296), .Z(n37299) );
  XNOR U37135 ( .A(n37294), .B(n37293), .Z(n37296) );
  XNOR U37136 ( .A(n37291), .B(n37290), .Z(n37293) );
  XNOR U37137 ( .A(n37288), .B(n37287), .Z(n37290) );
  XNOR U37138 ( .A(n37285), .B(n37284), .Z(n37287) );
  XNOR U37139 ( .A(n37282), .B(n37281), .Z(n37284) );
  XNOR U37140 ( .A(n37279), .B(n37278), .Z(n37281) );
  XNOR U37141 ( .A(n37276), .B(n37275), .Z(n37278) );
  XNOR U37142 ( .A(n37273), .B(n37272), .Z(n37275) );
  XNOR U37143 ( .A(n37270), .B(n37269), .Z(n37272) );
  XNOR U37144 ( .A(n37267), .B(n37266), .Z(n37269) );
  XNOR U37145 ( .A(n37264), .B(n37263), .Z(n37266) );
  XNOR U37146 ( .A(n37261), .B(n37260), .Z(n37263) );
  XNOR U37147 ( .A(n37258), .B(n37257), .Z(n37260) );
  XNOR U37148 ( .A(n37255), .B(n37254), .Z(n37257) );
  XNOR U37149 ( .A(n37252), .B(n37251), .Z(n37254) );
  XNOR U37150 ( .A(n37249), .B(n37248), .Z(n37251) );
  XNOR U37151 ( .A(n37246), .B(n37245), .Z(n37248) );
  XNOR U37152 ( .A(n37243), .B(n37242), .Z(n37245) );
  XNOR U37153 ( .A(n37240), .B(n37239), .Z(n37242) );
  XNOR U37154 ( .A(n37237), .B(n37236), .Z(n37239) );
  XNOR U37155 ( .A(n37234), .B(n37233), .Z(n37236) );
  XOR U37156 ( .A(n37231), .B(n37230), .Z(n37233) );
  XOR U37157 ( .A(n37228), .B(n37227), .Z(n37230) );
  XOR U37158 ( .A(n37224), .B(n37225), .Z(n37227) );
  AND U37159 ( .A(n39813), .B(n39814), .Z(n37225) );
  XOR U37160 ( .A(n37221), .B(n37222), .Z(n37224) );
  AND U37161 ( .A(n39815), .B(n39816), .Z(n37222) );
  XOR U37162 ( .A(n37218), .B(n37219), .Z(n37221) );
  AND U37163 ( .A(n39817), .B(n39818), .Z(n37219) );
  XNOR U37164 ( .A(n36967), .B(n37216), .Z(n37218) );
  AND U37165 ( .A(n39819), .B(n39820), .Z(n37216) );
  XOR U37166 ( .A(n36969), .B(n36968), .Z(n36967) );
  AND U37167 ( .A(n39821), .B(n39822), .Z(n36968) );
  XOR U37168 ( .A(n36971), .B(n36970), .Z(n36969) );
  AND U37169 ( .A(n39823), .B(n39824), .Z(n36970) );
  XOR U37170 ( .A(n36973), .B(n36972), .Z(n36971) );
  AND U37171 ( .A(n39825), .B(n39826), .Z(n36972) );
  XOR U37172 ( .A(n36975), .B(n36974), .Z(n36973) );
  AND U37173 ( .A(n39827), .B(n39828), .Z(n36974) );
  XOR U37174 ( .A(n36977), .B(n36976), .Z(n36975) );
  AND U37175 ( .A(n39829), .B(n39830), .Z(n36976) );
  XOR U37176 ( .A(n36979), .B(n36978), .Z(n36977) );
  AND U37177 ( .A(n39831), .B(n39832), .Z(n36978) );
  XOR U37178 ( .A(n36981), .B(n36980), .Z(n36979) );
  AND U37179 ( .A(n39833), .B(n39834), .Z(n36980) );
  XOR U37180 ( .A(n36983), .B(n36982), .Z(n36981) );
  AND U37181 ( .A(n39835), .B(n39836), .Z(n36982) );
  XOR U37182 ( .A(n36985), .B(n36984), .Z(n36983) );
  AND U37183 ( .A(n39837), .B(n39838), .Z(n36984) );
  XOR U37184 ( .A(n36987), .B(n36986), .Z(n36985) );
  AND U37185 ( .A(n39839), .B(n39840), .Z(n36986) );
  XOR U37186 ( .A(n36989), .B(n36988), .Z(n36987) );
  AND U37187 ( .A(n39841), .B(n39842), .Z(n36988) );
  XOR U37188 ( .A(n36991), .B(n36990), .Z(n36989) );
  AND U37189 ( .A(n39843), .B(n39844), .Z(n36990) );
  XOR U37190 ( .A(n36993), .B(n36992), .Z(n36991) );
  AND U37191 ( .A(n39845), .B(n39846), .Z(n36992) );
  XOR U37192 ( .A(n36995), .B(n36994), .Z(n36993) );
  AND U37193 ( .A(n39847), .B(n39848), .Z(n36994) );
  XOR U37194 ( .A(n36997), .B(n36996), .Z(n36995) );
  AND U37195 ( .A(n39849), .B(n39850), .Z(n36996) );
  XOR U37196 ( .A(n36999), .B(n36998), .Z(n36997) );
  AND U37197 ( .A(n39851), .B(n39852), .Z(n36998) );
  XOR U37198 ( .A(n37001), .B(n37000), .Z(n36999) );
  AND U37199 ( .A(n39853), .B(n39854), .Z(n37000) );
  XOR U37200 ( .A(n37003), .B(n37002), .Z(n37001) );
  AND U37201 ( .A(n39855), .B(n39856), .Z(n37002) );
  XOR U37202 ( .A(n37005), .B(n37004), .Z(n37003) );
  AND U37203 ( .A(n39857), .B(n39858), .Z(n37004) );
  XOR U37204 ( .A(n37007), .B(n37006), .Z(n37005) );
  AND U37205 ( .A(n39859), .B(n39860), .Z(n37006) );
  XOR U37206 ( .A(n37009), .B(n37008), .Z(n37007) );
  AND U37207 ( .A(n39861), .B(n39862), .Z(n37008) );
  XOR U37208 ( .A(n37011), .B(n37010), .Z(n37009) );
  AND U37209 ( .A(n39863), .B(n39864), .Z(n37010) );
  XOR U37210 ( .A(n37013), .B(n37012), .Z(n37011) );
  AND U37211 ( .A(n39865), .B(n39866), .Z(n37012) );
  XOR U37212 ( .A(n37015), .B(n37014), .Z(n37013) );
  AND U37213 ( .A(n39867), .B(n39868), .Z(n37014) );
  XOR U37214 ( .A(n37017), .B(n37016), .Z(n37015) );
  AND U37215 ( .A(n39869), .B(n39870), .Z(n37016) );
  XOR U37216 ( .A(n37019), .B(n37018), .Z(n37017) );
  AND U37217 ( .A(n39871), .B(n39872), .Z(n37018) );
  XOR U37218 ( .A(n37021), .B(n37020), .Z(n37019) );
  AND U37219 ( .A(n39873), .B(n39874), .Z(n37020) );
  XOR U37220 ( .A(n37023), .B(n37022), .Z(n37021) );
  AND U37221 ( .A(n39875), .B(n39876), .Z(n37022) );
  XOR U37222 ( .A(n37025), .B(n37024), .Z(n37023) );
  AND U37223 ( .A(n39877), .B(n39878), .Z(n37024) );
  XOR U37224 ( .A(n37027), .B(n37026), .Z(n37025) );
  AND U37225 ( .A(n39879), .B(n39880), .Z(n37026) );
  XOR U37226 ( .A(n37029), .B(n37028), .Z(n37027) );
  AND U37227 ( .A(n39881), .B(n39882), .Z(n37028) );
  XOR U37228 ( .A(n37031), .B(n37030), .Z(n37029) );
  AND U37229 ( .A(n39883), .B(n39884), .Z(n37030) );
  XOR U37230 ( .A(n37033), .B(n37032), .Z(n37031) );
  AND U37231 ( .A(n39885), .B(n39886), .Z(n37032) );
  XOR U37232 ( .A(n37035), .B(n37034), .Z(n37033) );
  AND U37233 ( .A(n39887), .B(n39888), .Z(n37034) );
  XOR U37234 ( .A(n37037), .B(n37036), .Z(n37035) );
  AND U37235 ( .A(n39889), .B(n39890), .Z(n37036) );
  XOR U37236 ( .A(n37039), .B(n37038), .Z(n37037) );
  AND U37237 ( .A(n39891), .B(n39892), .Z(n37038) );
  XOR U37238 ( .A(n37041), .B(n37040), .Z(n37039) );
  AND U37239 ( .A(n39893), .B(n39894), .Z(n37040) );
  XOR U37240 ( .A(n37043), .B(n37042), .Z(n37041) );
  AND U37241 ( .A(n39895), .B(n39896), .Z(n37042) );
  XOR U37242 ( .A(n37045), .B(n37044), .Z(n37043) );
  AND U37243 ( .A(n39897), .B(n39898), .Z(n37044) );
  XOR U37244 ( .A(n37047), .B(n37046), .Z(n37045) );
  AND U37245 ( .A(n39899), .B(n39900), .Z(n37046) );
  XOR U37246 ( .A(n37049), .B(n37048), .Z(n37047) );
  AND U37247 ( .A(n39901), .B(n39902), .Z(n37048) );
  XOR U37248 ( .A(n37051), .B(n37050), .Z(n37049) );
  AND U37249 ( .A(n39903), .B(n39904), .Z(n37050) );
  XOR U37250 ( .A(n37053), .B(n37052), .Z(n37051) );
  AND U37251 ( .A(n39905), .B(n39906), .Z(n37052) );
  XOR U37252 ( .A(n37055), .B(n37054), .Z(n37053) );
  AND U37253 ( .A(n39907), .B(n39908), .Z(n37054) );
  XOR U37254 ( .A(n37057), .B(n37056), .Z(n37055) );
  AND U37255 ( .A(n39909), .B(n39910), .Z(n37056) );
  XOR U37256 ( .A(n37059), .B(n37058), .Z(n37057) );
  AND U37257 ( .A(n39911), .B(n39912), .Z(n37058) );
  XOR U37258 ( .A(n37061), .B(n37060), .Z(n37059) );
  AND U37259 ( .A(n39913), .B(n39914), .Z(n37060) );
  XOR U37260 ( .A(n37063), .B(n37062), .Z(n37061) );
  AND U37261 ( .A(n39915), .B(n39916), .Z(n37062) );
  XOR U37262 ( .A(n37065), .B(n37064), .Z(n37063) );
  AND U37263 ( .A(n39917), .B(n39918), .Z(n37064) );
  XOR U37264 ( .A(n37067), .B(n37066), .Z(n37065) );
  AND U37265 ( .A(n39919), .B(n39920), .Z(n37066) );
  XOR U37266 ( .A(n37069), .B(n37068), .Z(n37067) );
  AND U37267 ( .A(n39921), .B(n39922), .Z(n37068) );
  XOR U37268 ( .A(n37071), .B(n37070), .Z(n37069) );
  AND U37269 ( .A(n39923), .B(n39924), .Z(n37070) );
  XOR U37270 ( .A(n37073), .B(n37072), .Z(n37071) );
  AND U37271 ( .A(n39925), .B(n39926), .Z(n37072) );
  XOR U37272 ( .A(n37075), .B(n37074), .Z(n37073) );
  AND U37273 ( .A(n39927), .B(n39928), .Z(n37074) );
  XOR U37274 ( .A(n37077), .B(n37076), .Z(n37075) );
  AND U37275 ( .A(n39929), .B(n39930), .Z(n37076) );
  XOR U37276 ( .A(n37079), .B(n37078), .Z(n37077) );
  AND U37277 ( .A(n39931), .B(n39932), .Z(n37078) );
  XOR U37278 ( .A(n37081), .B(n37080), .Z(n37079) );
  AND U37279 ( .A(n39933), .B(n39934), .Z(n37080) );
  XOR U37280 ( .A(n37083), .B(n37082), .Z(n37081) );
  AND U37281 ( .A(n39935), .B(n39936), .Z(n37082) );
  XOR U37282 ( .A(n37085), .B(n37084), .Z(n37083) );
  AND U37283 ( .A(n39937), .B(n39938), .Z(n37084) );
  XOR U37284 ( .A(n37087), .B(n37086), .Z(n37085) );
  AND U37285 ( .A(n39939), .B(n39940), .Z(n37086) );
  XOR U37286 ( .A(n37089), .B(n37088), .Z(n37087) );
  AND U37287 ( .A(n39941), .B(n39942), .Z(n37088) );
  XOR U37288 ( .A(n37091), .B(n37090), .Z(n37089) );
  AND U37289 ( .A(n39943), .B(n39944), .Z(n37090) );
  XOR U37290 ( .A(n37093), .B(n37092), .Z(n37091) );
  AND U37291 ( .A(n39945), .B(n39946), .Z(n37092) );
  XOR U37292 ( .A(n37095), .B(n37094), .Z(n37093) );
  AND U37293 ( .A(n39947), .B(n39948), .Z(n37094) );
  XOR U37294 ( .A(n37097), .B(n37096), .Z(n37095) );
  AND U37295 ( .A(n39949), .B(n39950), .Z(n37096) );
  XOR U37296 ( .A(n37099), .B(n37098), .Z(n37097) );
  AND U37297 ( .A(n39951), .B(n39952), .Z(n37098) );
  XOR U37298 ( .A(n37101), .B(n37100), .Z(n37099) );
  AND U37299 ( .A(n39953), .B(n39954), .Z(n37100) );
  XOR U37300 ( .A(n37103), .B(n37102), .Z(n37101) );
  AND U37301 ( .A(n39955), .B(n39956), .Z(n37102) );
  XOR U37302 ( .A(n37105), .B(n37104), .Z(n37103) );
  AND U37303 ( .A(n39957), .B(n39958), .Z(n37104) );
  XOR U37304 ( .A(n37107), .B(n37106), .Z(n37105) );
  AND U37305 ( .A(n39959), .B(n39960), .Z(n37106) );
  XOR U37306 ( .A(n37109), .B(n37108), .Z(n37107) );
  AND U37307 ( .A(n39961), .B(n39962), .Z(n37108) );
  XOR U37308 ( .A(n37111), .B(n37110), .Z(n37109) );
  AND U37309 ( .A(n39963), .B(n39964), .Z(n37110) );
  XOR U37310 ( .A(n37113), .B(n37112), .Z(n37111) );
  AND U37311 ( .A(n39965), .B(n39966), .Z(n37112) );
  XOR U37312 ( .A(n37115), .B(n37114), .Z(n37113) );
  AND U37313 ( .A(n39967), .B(n39968), .Z(n37114) );
  XOR U37314 ( .A(n37117), .B(n37116), .Z(n37115) );
  AND U37315 ( .A(n39969), .B(n39970), .Z(n37116) );
  XOR U37316 ( .A(n37119), .B(n37118), .Z(n37117) );
  AND U37317 ( .A(n39971), .B(n39972), .Z(n37118) );
  XOR U37318 ( .A(n37121), .B(n37120), .Z(n37119) );
  AND U37319 ( .A(n39973), .B(n39974), .Z(n37120) );
  XOR U37320 ( .A(n37123), .B(n37122), .Z(n37121) );
  AND U37321 ( .A(n39975), .B(n39976), .Z(n37122) );
  XOR U37322 ( .A(n37125), .B(n37124), .Z(n37123) );
  AND U37323 ( .A(n39977), .B(n39978), .Z(n37124) );
  XOR U37324 ( .A(n37127), .B(n37126), .Z(n37125) );
  AND U37325 ( .A(n39979), .B(n39980), .Z(n37126) );
  XOR U37326 ( .A(n37129), .B(n37128), .Z(n37127) );
  AND U37327 ( .A(n39981), .B(n39982), .Z(n37128) );
  XOR U37328 ( .A(n37131), .B(n37130), .Z(n37129) );
  AND U37329 ( .A(n39983), .B(n39984), .Z(n37130) );
  XOR U37330 ( .A(n37133), .B(n37132), .Z(n37131) );
  AND U37331 ( .A(n39985), .B(n39986), .Z(n37132) );
  XOR U37332 ( .A(n37135), .B(n37134), .Z(n37133) );
  AND U37333 ( .A(n39987), .B(n39988), .Z(n37134) );
  XOR U37334 ( .A(n37137), .B(n37136), .Z(n37135) );
  AND U37335 ( .A(n39989), .B(n39990), .Z(n37136) );
  XOR U37336 ( .A(n37139), .B(n37138), .Z(n37137) );
  AND U37337 ( .A(n39991), .B(n39992), .Z(n37138) );
  XOR U37338 ( .A(n37141), .B(n37140), .Z(n37139) );
  AND U37339 ( .A(n39993), .B(n39994), .Z(n37140) );
  XOR U37340 ( .A(n37143), .B(n37142), .Z(n37141) );
  AND U37341 ( .A(n39995), .B(n39996), .Z(n37142) );
  XOR U37342 ( .A(n37145), .B(n37144), .Z(n37143) );
  AND U37343 ( .A(n39997), .B(n39998), .Z(n37144) );
  XOR U37344 ( .A(n37147), .B(n37146), .Z(n37145) );
  AND U37345 ( .A(n39999), .B(n40000), .Z(n37146) );
  XOR U37346 ( .A(n37149), .B(n37148), .Z(n37147) );
  AND U37347 ( .A(n40001), .B(n40002), .Z(n37148) );
  XOR U37348 ( .A(n37151), .B(n37150), .Z(n37149) );
  AND U37349 ( .A(n40003), .B(n40004), .Z(n37150) );
  XOR U37350 ( .A(n37153), .B(n37152), .Z(n37151) );
  AND U37351 ( .A(n40005), .B(n40006), .Z(n37152) );
  XOR U37352 ( .A(n37155), .B(n37154), .Z(n37153) );
  AND U37353 ( .A(n40007), .B(n40008), .Z(n37154) );
  XOR U37354 ( .A(n37157), .B(n37156), .Z(n37155) );
  AND U37355 ( .A(n40009), .B(n40010), .Z(n37156) );
  XOR U37356 ( .A(n37159), .B(n37158), .Z(n37157) );
  AND U37357 ( .A(n40011), .B(n40012), .Z(n37158) );
  XOR U37358 ( .A(n37212), .B(n37160), .Z(n37159) );
  AND U37359 ( .A(n40013), .B(n40014), .Z(n37160) );
  XOR U37360 ( .A(n37214), .B(n37213), .Z(n37212) );
  AND U37361 ( .A(n40015), .B(n40016), .Z(n37213) );
  XOR U37362 ( .A(n37195), .B(n37215), .Z(n37214) );
  AND U37363 ( .A(n40017), .B(n40018), .Z(n37215) );
  XOR U37364 ( .A(n37197), .B(n37196), .Z(n37195) );
  AND U37365 ( .A(n40019), .B(n40020), .Z(n37196) );
  XOR U37366 ( .A(n37199), .B(n37198), .Z(n37197) );
  AND U37367 ( .A(n40021), .B(n40022), .Z(n37198) );
  XOR U37368 ( .A(n37203), .B(n37200), .Z(n37199) );
  AND U37369 ( .A(n40023), .B(n40024), .Z(n37200) );
  XOR U37370 ( .A(n37205), .B(n37204), .Z(n37203) );
  AND U37371 ( .A(n40025), .B(n40026), .Z(n37204) );
  XOR U37372 ( .A(n37208), .B(n37206), .Z(n37205) );
  AND U37373 ( .A(n40027), .B(n40028), .Z(n37206) );
  XOR U37374 ( .A(n37210), .B(n37209), .Z(n37208) );
  AND U37375 ( .A(n40029), .B(n40030), .Z(n37209) );
  XOR U37376 ( .A(n37175), .B(n37211), .Z(n37210) );
  AND U37377 ( .A(n40031), .B(n40032), .Z(n37211) );
  XNOR U37378 ( .A(n37182), .B(n37176), .Z(n37175) );
  AND U37379 ( .A(n40033), .B(n40034), .Z(n37176) );
  XOR U37380 ( .A(n37181), .B(n37173), .Z(n37182) );
  AND U37381 ( .A(n40035), .B(n40036), .Z(n37173) );
  XOR U37382 ( .A(n37194), .B(n37172), .Z(n37181) );
  AND U37383 ( .A(n40037), .B(n40038), .Z(n37172) );
  XNOR U37384 ( .A(n40039), .B(n40040), .Z(n37194) );
  XOR U37385 ( .A(n37192), .B(n40041), .Z(n40040) );
  XOR U37386 ( .A(n37190), .B(n37188), .Z(n40041) );
  AND U37387 ( .A(n40042), .B(n40043), .Z(n37188) );
  AND U37388 ( .A(n40044), .B(n40045), .Z(n37190) );
  AND U37389 ( .A(n40046), .B(n40047), .Z(n37192) );
  XNOR U37390 ( .A(n40048), .B(n37191), .Z(n40039) );
  XOR U37391 ( .A(n40049), .B(n40050), .Z(n37191) );
  XOR U37392 ( .A(n40051), .B(n40052), .Z(n40050) );
  AND U37393 ( .A(n40053), .B(n40054), .Z(n40052) );
  XNOR U37394 ( .A(n40055), .B(n40056), .Z(n40049) );
  NOR U37395 ( .A(n40057), .B(n40058), .Z(n40056) );
  AND U37396 ( .A(n40059), .B(n40060), .Z(n40058) );
  IV U37397 ( .A(n40061), .Z(n40057) );
  NOR U37398 ( .A(n40051), .B(n40062), .Z(n40061) );
  AND U37399 ( .A(n40063), .B(n40064), .Z(n40062) );
  NOR U37400 ( .A(n40053), .B(n40063), .Z(n40055) );
  XNOR U37401 ( .A(n37193), .B(n37171), .Z(n40048) );
  AND U37402 ( .A(n40065), .B(n40066), .Z(n37171) );
  AND U37403 ( .A(n40067), .B(n40068), .Z(n37193) );
  XOR U37404 ( .A(n40069), .B(n40070), .Z(n37228) );
  NOR U37405 ( .A(n40071), .B(n40072), .Z(n40070) );
  IV U37406 ( .A(n40069), .Z(n40071) );
  XOR U37407 ( .A(n40073), .B(n40074), .Z(n37231) );
  NOR U37408 ( .A(n40073), .B(n40075), .Z(n40074) );
  XNOR U37409 ( .A(n40076), .B(n40077), .Z(n37234) );
  AND U37410 ( .A(n40076), .B(n40078), .Z(n40077) );
  XNOR U37411 ( .A(n40079), .B(n40080), .Z(n37237) );
  AND U37412 ( .A(n40079), .B(n40081), .Z(n40080) );
  XNOR U37413 ( .A(n40082), .B(n40083), .Z(n37240) );
  AND U37414 ( .A(n40082), .B(n40084), .Z(n40083) );
  XNOR U37415 ( .A(n40085), .B(n40086), .Z(n37243) );
  AND U37416 ( .A(n40085), .B(n40087), .Z(n40086) );
  XNOR U37417 ( .A(n40088), .B(n40089), .Z(n37246) );
  AND U37418 ( .A(n40088), .B(n40090), .Z(n40089) );
  XNOR U37419 ( .A(n40091), .B(n40092), .Z(n37249) );
  AND U37420 ( .A(n40091), .B(n40093), .Z(n40092) );
  XNOR U37421 ( .A(n40094), .B(n40095), .Z(n37252) );
  AND U37422 ( .A(n40094), .B(n40096), .Z(n40095) );
  XNOR U37423 ( .A(n40097), .B(n40098), .Z(n37255) );
  AND U37424 ( .A(n40097), .B(n40099), .Z(n40098) );
  XNOR U37425 ( .A(n40100), .B(n40101), .Z(n37258) );
  AND U37426 ( .A(n40100), .B(n40102), .Z(n40101) );
  XNOR U37427 ( .A(n40103), .B(n40104), .Z(n37261) );
  AND U37428 ( .A(n40103), .B(n40105), .Z(n40104) );
  XNOR U37429 ( .A(n40106), .B(n40107), .Z(n37264) );
  AND U37430 ( .A(n40106), .B(n40108), .Z(n40107) );
  XNOR U37431 ( .A(n40109), .B(n40110), .Z(n37267) );
  AND U37432 ( .A(n40109), .B(n40111), .Z(n40110) );
  XNOR U37433 ( .A(n40112), .B(n40113), .Z(n37270) );
  AND U37434 ( .A(n40112), .B(n40114), .Z(n40113) );
  XNOR U37435 ( .A(n40115), .B(n40116), .Z(n37273) );
  AND U37436 ( .A(n40115), .B(n40117), .Z(n40116) );
  XNOR U37437 ( .A(n40118), .B(n40119), .Z(n37276) );
  AND U37438 ( .A(n40118), .B(n40120), .Z(n40119) );
  XNOR U37439 ( .A(n40121), .B(n40122), .Z(n37279) );
  AND U37440 ( .A(n40121), .B(n40123), .Z(n40122) );
  XNOR U37441 ( .A(n40124), .B(n40125), .Z(n37282) );
  AND U37442 ( .A(n40124), .B(n40126), .Z(n40125) );
  XNOR U37443 ( .A(n40127), .B(n40128), .Z(n37285) );
  AND U37444 ( .A(n40127), .B(n40129), .Z(n40128) );
  XNOR U37445 ( .A(n40130), .B(n40131), .Z(n37288) );
  AND U37446 ( .A(n40130), .B(n40132), .Z(n40131) );
  XNOR U37447 ( .A(n40133), .B(n40134), .Z(n37291) );
  AND U37448 ( .A(n40133), .B(n40135), .Z(n40134) );
  XNOR U37449 ( .A(n40136), .B(n40137), .Z(n37294) );
  AND U37450 ( .A(n40136), .B(n40138), .Z(n40137) );
  XNOR U37451 ( .A(n40139), .B(n40140), .Z(n37297) );
  AND U37452 ( .A(n40139), .B(n40141), .Z(n40140) );
  XNOR U37453 ( .A(n40142), .B(n40143), .Z(n37300) );
  AND U37454 ( .A(n40142), .B(n40144), .Z(n40143) );
  XNOR U37455 ( .A(n40145), .B(n40146), .Z(n37303) );
  AND U37456 ( .A(n40145), .B(n40147), .Z(n40146) );
  XNOR U37457 ( .A(n40148), .B(n40149), .Z(n37306) );
  AND U37458 ( .A(n40148), .B(n40150), .Z(n40149) );
  XNOR U37459 ( .A(n40151), .B(n40152), .Z(n37309) );
  AND U37460 ( .A(n40151), .B(n40153), .Z(n40152) );
  XNOR U37461 ( .A(n40154), .B(n40155), .Z(n37312) );
  AND U37462 ( .A(n40154), .B(n40156), .Z(n40155) );
  XNOR U37463 ( .A(n40157), .B(n40158), .Z(n37315) );
  AND U37464 ( .A(n40157), .B(n40159), .Z(n40158) );
  XNOR U37465 ( .A(n40160), .B(n40161), .Z(n37318) );
  AND U37466 ( .A(n40160), .B(n40162), .Z(n40161) );
  XNOR U37467 ( .A(n40163), .B(n40164), .Z(n37321) );
  AND U37468 ( .A(n40163), .B(n40165), .Z(n40164) );
  XNOR U37469 ( .A(n40166), .B(n40167), .Z(n37324) );
  AND U37470 ( .A(n40166), .B(n40168), .Z(n40167) );
  XNOR U37471 ( .A(n40169), .B(n40170), .Z(n37327) );
  AND U37472 ( .A(n40169), .B(n40171), .Z(n40170) );
  XNOR U37473 ( .A(n40172), .B(n40173), .Z(n37330) );
  AND U37474 ( .A(n40172), .B(n40174), .Z(n40173) );
  XNOR U37475 ( .A(n40175), .B(n40176), .Z(n37333) );
  AND U37476 ( .A(n40175), .B(n40177), .Z(n40176) );
  XNOR U37477 ( .A(n40178), .B(n40179), .Z(n37336) );
  AND U37478 ( .A(n40178), .B(n40180), .Z(n40179) );
  XNOR U37479 ( .A(n40181), .B(n40182), .Z(n37339) );
  AND U37480 ( .A(n40181), .B(n40183), .Z(n40182) );
  XNOR U37481 ( .A(n40184), .B(n40185), .Z(n37342) );
  AND U37482 ( .A(n40184), .B(n40186), .Z(n40185) );
  XNOR U37483 ( .A(n40187), .B(n40188), .Z(n37345) );
  AND U37484 ( .A(n40187), .B(n40189), .Z(n40188) );
  XNOR U37485 ( .A(n40190), .B(n40191), .Z(n37348) );
  AND U37486 ( .A(n40190), .B(n40192), .Z(n40191) );
  XNOR U37487 ( .A(n40193), .B(n40194), .Z(n37351) );
  AND U37488 ( .A(n40193), .B(n40195), .Z(n40194) );
  XNOR U37489 ( .A(n40196), .B(n40197), .Z(n37354) );
  AND U37490 ( .A(n40196), .B(n40198), .Z(n40197) );
  XNOR U37491 ( .A(n40199), .B(n40200), .Z(n37357) );
  AND U37492 ( .A(n40199), .B(n40201), .Z(n40200) );
  XNOR U37493 ( .A(n40202), .B(n40203), .Z(n37360) );
  AND U37494 ( .A(n40202), .B(n40204), .Z(n40203) );
  XNOR U37495 ( .A(n40205), .B(n40206), .Z(n37363) );
  AND U37496 ( .A(n40205), .B(n40207), .Z(n40206) );
  XNOR U37497 ( .A(n40208), .B(n40209), .Z(n37366) );
  AND U37498 ( .A(n40208), .B(n40210), .Z(n40209) );
  XNOR U37499 ( .A(n40211), .B(n40212), .Z(n37369) );
  AND U37500 ( .A(n40211), .B(n40213), .Z(n40212) );
  XNOR U37501 ( .A(n40214), .B(n40215), .Z(n37372) );
  AND U37502 ( .A(n40214), .B(n40216), .Z(n40215) );
  XNOR U37503 ( .A(n40217), .B(n40218), .Z(n37375) );
  AND U37504 ( .A(n40217), .B(n40219), .Z(n40218) );
  XNOR U37505 ( .A(n40220), .B(n40221), .Z(n37378) );
  AND U37506 ( .A(n40220), .B(n40222), .Z(n40221) );
  XNOR U37507 ( .A(n40223), .B(n40224), .Z(n37381) );
  AND U37508 ( .A(n40223), .B(n40225), .Z(n40224) );
  XNOR U37509 ( .A(n40226), .B(n40227), .Z(n37384) );
  AND U37510 ( .A(n40226), .B(n40228), .Z(n40227) );
  XNOR U37511 ( .A(n40229), .B(n40230), .Z(n37387) );
  AND U37512 ( .A(n40229), .B(n40231), .Z(n40230) );
  XNOR U37513 ( .A(n40232), .B(n40233), .Z(n37390) );
  AND U37514 ( .A(n40232), .B(n40234), .Z(n40233) );
  XNOR U37515 ( .A(n40235), .B(n40236), .Z(n37393) );
  AND U37516 ( .A(n40235), .B(n40237), .Z(n40236) );
  XNOR U37517 ( .A(n40238), .B(n40239), .Z(n37396) );
  AND U37518 ( .A(n40238), .B(n40240), .Z(n40239) );
  XNOR U37519 ( .A(n40241), .B(n40242), .Z(n37399) );
  AND U37520 ( .A(n40241), .B(n40243), .Z(n40242) );
  XNOR U37521 ( .A(n40244), .B(n40245), .Z(n37402) );
  AND U37522 ( .A(n40244), .B(n40246), .Z(n40245) );
  XNOR U37523 ( .A(n40247), .B(n40248), .Z(n37405) );
  AND U37524 ( .A(n40247), .B(n40249), .Z(n40248) );
  XNOR U37525 ( .A(n40250), .B(n40251), .Z(n37408) );
  AND U37526 ( .A(n40250), .B(n40252), .Z(n40251) );
  XNOR U37527 ( .A(n40253), .B(n40254), .Z(n37411) );
  AND U37528 ( .A(n40253), .B(n40255), .Z(n40254) );
  XNOR U37529 ( .A(n40256), .B(n40257), .Z(n37414) );
  AND U37530 ( .A(n40256), .B(n40258), .Z(n40257) );
  XNOR U37531 ( .A(n40259), .B(n40260), .Z(n37417) );
  AND U37532 ( .A(n40259), .B(n40261), .Z(n40260) );
  XNOR U37533 ( .A(n40262), .B(n40263), .Z(n37420) );
  AND U37534 ( .A(n40262), .B(n40264), .Z(n40263) );
  XNOR U37535 ( .A(n40265), .B(n40266), .Z(n37423) );
  AND U37536 ( .A(n40265), .B(n40267), .Z(n40266) );
  XNOR U37537 ( .A(n40268), .B(n40269), .Z(n37426) );
  AND U37538 ( .A(n40268), .B(n40270), .Z(n40269) );
  XNOR U37539 ( .A(n40271), .B(n40272), .Z(n37429) );
  AND U37540 ( .A(n40271), .B(n40273), .Z(n40272) );
  XNOR U37541 ( .A(n40274), .B(n40275), .Z(n37432) );
  AND U37542 ( .A(n40274), .B(n40276), .Z(n40275) );
  XNOR U37543 ( .A(n40277), .B(n40278), .Z(n37435) );
  AND U37544 ( .A(n40277), .B(n40279), .Z(n40278) );
  XNOR U37545 ( .A(n40280), .B(n40281), .Z(n37438) );
  AND U37546 ( .A(n40280), .B(n40282), .Z(n40281) );
  XNOR U37547 ( .A(n40283), .B(n40284), .Z(n37441) );
  AND U37548 ( .A(n40283), .B(n40285), .Z(n40284) );
  XNOR U37549 ( .A(n40286), .B(n40287), .Z(n37444) );
  AND U37550 ( .A(n40286), .B(n40288), .Z(n40287) );
  XNOR U37551 ( .A(n40289), .B(n40290), .Z(n37447) );
  AND U37552 ( .A(n40289), .B(n40291), .Z(n40290) );
  XNOR U37553 ( .A(n40292), .B(n40293), .Z(n37450) );
  AND U37554 ( .A(n40292), .B(n40294), .Z(n40293) );
  XNOR U37555 ( .A(n40295), .B(n40296), .Z(n37453) );
  AND U37556 ( .A(n40295), .B(n40297), .Z(n40296) );
  XNOR U37557 ( .A(n40298), .B(n40299), .Z(n37456) );
  AND U37558 ( .A(n40298), .B(n40300), .Z(n40299) );
  XNOR U37559 ( .A(n40301), .B(n40302), .Z(n37459) );
  AND U37560 ( .A(n40301), .B(n40303), .Z(n40302) );
  XNOR U37561 ( .A(n40304), .B(n40305), .Z(n37462) );
  AND U37562 ( .A(n40304), .B(n40306), .Z(n40305) );
  XNOR U37563 ( .A(n40307), .B(n40308), .Z(n37465) );
  AND U37564 ( .A(n40307), .B(n40309), .Z(n40308) );
  XNOR U37565 ( .A(n40310), .B(n40311), .Z(n37468) );
  AND U37566 ( .A(n40310), .B(n40312), .Z(n40311) );
  XNOR U37567 ( .A(n40313), .B(n40314), .Z(n37471) );
  AND U37568 ( .A(n40313), .B(n40315), .Z(n40314) );
  XNOR U37569 ( .A(n40316), .B(n40317), .Z(n37474) );
  AND U37570 ( .A(n40316), .B(n40318), .Z(n40317) );
  XNOR U37571 ( .A(n40319), .B(n40320), .Z(n37477) );
  AND U37572 ( .A(n40319), .B(n40321), .Z(n40320) );
  XNOR U37573 ( .A(n40322), .B(n40323), .Z(n37480) );
  AND U37574 ( .A(n40322), .B(n40324), .Z(n40323) );
  XNOR U37575 ( .A(n40325), .B(n40326), .Z(n37483) );
  AND U37576 ( .A(n40325), .B(n40327), .Z(n40326) );
  XNOR U37577 ( .A(n40328), .B(n40329), .Z(n37486) );
  AND U37578 ( .A(n40328), .B(n40330), .Z(n40329) );
  XNOR U37579 ( .A(n40331), .B(n40332), .Z(n37489) );
  AND U37580 ( .A(n40331), .B(n40333), .Z(n40332) );
  XNOR U37581 ( .A(n40334), .B(n40335), .Z(n37492) );
  AND U37582 ( .A(n40334), .B(n40336), .Z(n40335) );
  XNOR U37583 ( .A(n40337), .B(n40338), .Z(n37495) );
  AND U37584 ( .A(n40337), .B(n40339), .Z(n40338) );
  XNOR U37585 ( .A(n40340), .B(n40341), .Z(n37498) );
  AND U37586 ( .A(n40340), .B(n40342), .Z(n40341) );
  XNOR U37587 ( .A(n40343), .B(n40344), .Z(n37501) );
  AND U37588 ( .A(n40343), .B(n40345), .Z(n40344) );
  XNOR U37589 ( .A(n40346), .B(n40347), .Z(n37504) );
  AND U37590 ( .A(n40346), .B(n40348), .Z(n40347) );
  XNOR U37591 ( .A(n40349), .B(n40350), .Z(n37507) );
  AND U37592 ( .A(n40349), .B(n40351), .Z(n40350) );
  XNOR U37593 ( .A(n40352), .B(n40353), .Z(n37510) );
  AND U37594 ( .A(n40352), .B(n40354), .Z(n40353) );
  XNOR U37595 ( .A(n40355), .B(n40356), .Z(n37513) );
  AND U37596 ( .A(n40355), .B(n40357), .Z(n40356) );
  XNOR U37597 ( .A(n40358), .B(n40359), .Z(n37516) );
  AND U37598 ( .A(n40358), .B(n40360), .Z(n40359) );
  XNOR U37599 ( .A(n40361), .B(n40362), .Z(n37519) );
  AND U37600 ( .A(n40361), .B(n40363), .Z(n40362) );
  XNOR U37601 ( .A(n40364), .B(n40365), .Z(n37522) );
  AND U37602 ( .A(n40364), .B(n40366), .Z(n40365) );
  XNOR U37603 ( .A(n40367), .B(n40368), .Z(n37525) );
  AND U37604 ( .A(n40367), .B(n40369), .Z(n40368) );
  XNOR U37605 ( .A(n40370), .B(n40371), .Z(n37528) );
  AND U37606 ( .A(n40370), .B(n40372), .Z(n40371) );
  XNOR U37607 ( .A(n40373), .B(n40374), .Z(n37531) );
  AND U37608 ( .A(n40373), .B(n40375), .Z(n40374) );
  XNOR U37609 ( .A(n40376), .B(n40377), .Z(n37534) );
  AND U37610 ( .A(n40376), .B(n40378), .Z(n40377) );
  XNOR U37611 ( .A(n40379), .B(n40380), .Z(n37537) );
  AND U37612 ( .A(n40379), .B(n40381), .Z(n40380) );
  XNOR U37613 ( .A(n40382), .B(n40383), .Z(n37540) );
  AND U37614 ( .A(n40382), .B(n40384), .Z(n40383) );
  XNOR U37615 ( .A(n40385), .B(n40386), .Z(n37543) );
  AND U37616 ( .A(n40385), .B(n40387), .Z(n40386) );
  XNOR U37617 ( .A(n40388), .B(n40389), .Z(n37546) );
  AND U37618 ( .A(n40388), .B(n40390), .Z(n40389) );
  XNOR U37619 ( .A(n40391), .B(n40392), .Z(n37549) );
  AND U37620 ( .A(n40391), .B(n40393), .Z(n40392) );
  XNOR U37621 ( .A(n40394), .B(n40395), .Z(n37552) );
  AND U37622 ( .A(n40394), .B(n40396), .Z(n40395) );
  XNOR U37623 ( .A(n40397), .B(n40398), .Z(n37555) );
  AND U37624 ( .A(n40397), .B(n40399), .Z(n40398) );
  XNOR U37625 ( .A(n40400), .B(n40401), .Z(n37558) );
  AND U37626 ( .A(n40400), .B(n40402), .Z(n40401) );
  XNOR U37627 ( .A(n40403), .B(n40404), .Z(n37561) );
  AND U37628 ( .A(n40403), .B(n40405), .Z(n40404) );
  XNOR U37629 ( .A(n40406), .B(n40407), .Z(n37564) );
  AND U37630 ( .A(n40406), .B(n40408), .Z(n40407) );
  XNOR U37631 ( .A(n40409), .B(n40410), .Z(n37567) );
  AND U37632 ( .A(n40409), .B(n40411), .Z(n40410) );
  XNOR U37633 ( .A(n40412), .B(n40413), .Z(n37570) );
  AND U37634 ( .A(n40412), .B(n40414), .Z(n40413) );
  XNOR U37635 ( .A(n40415), .B(n40416), .Z(n37573) );
  AND U37636 ( .A(n40415), .B(n40417), .Z(n40416) );
  XNOR U37637 ( .A(n40418), .B(n40419), .Z(n37576) );
  AND U37638 ( .A(n40418), .B(n40420), .Z(n40419) );
  XNOR U37639 ( .A(n40421), .B(n40422), .Z(n37579) );
  AND U37640 ( .A(n40421), .B(n40423), .Z(n40422) );
  XNOR U37641 ( .A(n40424), .B(n40425), .Z(n37582) );
  AND U37642 ( .A(n40424), .B(n40426), .Z(n40425) );
  XNOR U37643 ( .A(n40427), .B(n40428), .Z(n37585) );
  AND U37644 ( .A(n40427), .B(n40429), .Z(n40428) );
  XNOR U37645 ( .A(n40430), .B(n40431), .Z(n37588) );
  AND U37646 ( .A(n40430), .B(n40432), .Z(n40431) );
  XNOR U37647 ( .A(n40433), .B(n40434), .Z(n37591) );
  AND U37648 ( .A(n40433), .B(n40435), .Z(n40434) );
  XNOR U37649 ( .A(n40436), .B(n40437), .Z(n37594) );
  AND U37650 ( .A(n40436), .B(n40438), .Z(n40437) );
  XNOR U37651 ( .A(n40439), .B(n40440), .Z(n37597) );
  AND U37652 ( .A(n40439), .B(n40441), .Z(n40440) );
  XNOR U37653 ( .A(n40442), .B(n40443), .Z(n37600) );
  AND U37654 ( .A(n40442), .B(n40444), .Z(n40443) );
  XNOR U37655 ( .A(n40445), .B(n40446), .Z(n37603) );
  AND U37656 ( .A(n40445), .B(n40447), .Z(n40446) );
  XNOR U37657 ( .A(n40448), .B(n40449), .Z(n37606) );
  AND U37658 ( .A(n40448), .B(n40450), .Z(n40449) );
  XNOR U37659 ( .A(n40451), .B(n40452), .Z(n37609) );
  AND U37660 ( .A(n40451), .B(n40453), .Z(n40452) );
  XNOR U37661 ( .A(n40454), .B(n40455), .Z(n37612) );
  AND U37662 ( .A(n40454), .B(n40456), .Z(n40455) );
  XNOR U37663 ( .A(n40457), .B(n40458), .Z(n37615) );
  AND U37664 ( .A(n40457), .B(n40459), .Z(n40458) );
  XNOR U37665 ( .A(n40460), .B(n40461), .Z(n37618) );
  AND U37666 ( .A(n40460), .B(n40462), .Z(n40461) );
  XNOR U37667 ( .A(n40463), .B(n40464), .Z(n37621) );
  AND U37668 ( .A(n40463), .B(n40465), .Z(n40464) );
  XNOR U37669 ( .A(n40466), .B(n40467), .Z(n37624) );
  AND U37670 ( .A(n40466), .B(n40468), .Z(n40467) );
  XNOR U37671 ( .A(n40469), .B(n40470), .Z(n37627) );
  AND U37672 ( .A(n40469), .B(n40471), .Z(n40470) );
  XNOR U37673 ( .A(n40472), .B(n40473), .Z(n37630) );
  AND U37674 ( .A(n40472), .B(n40474), .Z(n40473) );
  XNOR U37675 ( .A(n40475), .B(n40476), .Z(n37633) );
  AND U37676 ( .A(n40475), .B(n40477), .Z(n40476) );
  XNOR U37677 ( .A(n40478), .B(n40479), .Z(n37636) );
  AND U37678 ( .A(n40478), .B(n40480), .Z(n40479) );
  XNOR U37679 ( .A(n40481), .B(n40482), .Z(n37639) );
  AND U37680 ( .A(n40481), .B(n40483), .Z(n40482) );
  XNOR U37681 ( .A(n40484), .B(n40485), .Z(n37642) );
  AND U37682 ( .A(n40484), .B(n40486), .Z(n40485) );
  XNOR U37683 ( .A(n40487), .B(n40488), .Z(n37645) );
  AND U37684 ( .A(n40487), .B(n40489), .Z(n40488) );
  XNOR U37685 ( .A(n40490), .B(n40491), .Z(n37648) );
  AND U37686 ( .A(n40490), .B(n40492), .Z(n40491) );
  XNOR U37687 ( .A(n40493), .B(n40494), .Z(n37651) );
  AND U37688 ( .A(n40493), .B(n40495), .Z(n40494) );
  XNOR U37689 ( .A(n40496), .B(n40497), .Z(n37654) );
  AND U37690 ( .A(n40496), .B(n40498), .Z(n40497) );
  XNOR U37691 ( .A(n40499), .B(n40500), .Z(n37657) );
  AND U37692 ( .A(n40499), .B(n40501), .Z(n40500) );
  XNOR U37693 ( .A(n40502), .B(n40503), .Z(n37660) );
  AND U37694 ( .A(n40502), .B(n40504), .Z(n40503) );
  XNOR U37695 ( .A(n40505), .B(n40506), .Z(n37663) );
  AND U37696 ( .A(n40505), .B(n40507), .Z(n40506) );
  XNOR U37697 ( .A(n40508), .B(n40509), .Z(n37666) );
  AND U37698 ( .A(n40508), .B(n40510), .Z(n40509) );
  XNOR U37699 ( .A(n40511), .B(n40512), .Z(n37669) );
  AND U37700 ( .A(n40511), .B(n40513), .Z(n40512) );
  XNOR U37701 ( .A(n40514), .B(n40515), .Z(n37672) );
  AND U37702 ( .A(n40514), .B(n40516), .Z(n40515) );
  XNOR U37703 ( .A(n40517), .B(n40518), .Z(n37675) );
  AND U37704 ( .A(n40517), .B(n40519), .Z(n40518) );
  XNOR U37705 ( .A(n40520), .B(n40521), .Z(n37678) );
  AND U37706 ( .A(n40520), .B(n40522), .Z(n40521) );
  XNOR U37707 ( .A(n40523), .B(n40524), .Z(n37681) );
  AND U37708 ( .A(n40523), .B(n40525), .Z(n40524) );
  XNOR U37709 ( .A(n40526), .B(n40527), .Z(n37684) );
  AND U37710 ( .A(n40526), .B(n40528), .Z(n40527) );
  XNOR U37711 ( .A(n40529), .B(n40530), .Z(n37687) );
  AND U37712 ( .A(n40529), .B(n40531), .Z(n40530) );
  XNOR U37713 ( .A(n40532), .B(n40533), .Z(n37690) );
  AND U37714 ( .A(n40532), .B(n40534), .Z(n40533) );
  XNOR U37715 ( .A(n40535), .B(n40536), .Z(n37693) );
  AND U37716 ( .A(n40535), .B(n40537), .Z(n40536) );
  XNOR U37717 ( .A(n40538), .B(n40539), .Z(n37696) );
  AND U37718 ( .A(n40538), .B(n40540), .Z(n40539) );
  XNOR U37719 ( .A(n40541), .B(n40542), .Z(n37699) );
  AND U37720 ( .A(n40541), .B(n40543), .Z(n40542) );
  XNOR U37721 ( .A(n40544), .B(n40545), .Z(n37702) );
  AND U37722 ( .A(n40544), .B(n40546), .Z(n40545) );
  XNOR U37723 ( .A(n40547), .B(n40548), .Z(n37705) );
  AND U37724 ( .A(n40547), .B(n40549), .Z(n40548) );
  XNOR U37725 ( .A(n40550), .B(n40551), .Z(n37708) );
  AND U37726 ( .A(n40550), .B(n40552), .Z(n40551) );
  XNOR U37727 ( .A(n40553), .B(n40554), .Z(n37711) );
  AND U37728 ( .A(n40553), .B(n40555), .Z(n40554) );
  XNOR U37729 ( .A(n40556), .B(n40557), .Z(n37714) );
  AND U37730 ( .A(n40556), .B(n40558), .Z(n40557) );
  XNOR U37731 ( .A(n40559), .B(n40560), .Z(n37717) );
  AND U37732 ( .A(n40559), .B(n40561), .Z(n40560) );
  XNOR U37733 ( .A(n40562), .B(n40563), .Z(n37720) );
  AND U37734 ( .A(n40562), .B(n40564), .Z(n40563) );
  XNOR U37735 ( .A(n40565), .B(n40566), .Z(n37723) );
  AND U37736 ( .A(n40565), .B(n40567), .Z(n40566) );
  XNOR U37737 ( .A(n40568), .B(n40569), .Z(n37726) );
  AND U37738 ( .A(n40568), .B(n40570), .Z(n40569) );
  XNOR U37739 ( .A(n40571), .B(n40572), .Z(n37729) );
  AND U37740 ( .A(n40571), .B(n40573), .Z(n40572) );
  XNOR U37741 ( .A(n40574), .B(n40575), .Z(n37732) );
  AND U37742 ( .A(n40574), .B(n40576), .Z(n40575) );
  XNOR U37743 ( .A(n40577), .B(n40578), .Z(n37735) );
  AND U37744 ( .A(n40577), .B(n40579), .Z(n40578) );
  XNOR U37745 ( .A(n40580), .B(n40581), .Z(n37738) );
  AND U37746 ( .A(n40580), .B(n40582), .Z(n40581) );
  XNOR U37747 ( .A(n40583), .B(n40584), .Z(n37741) );
  AND U37748 ( .A(n40583), .B(n40585), .Z(n40584) );
  XNOR U37749 ( .A(n40586), .B(n40587), .Z(n37744) );
  AND U37750 ( .A(n40586), .B(n40588), .Z(n40587) );
  XNOR U37751 ( .A(n40589), .B(n40590), .Z(n37747) );
  AND U37752 ( .A(n40589), .B(n40591), .Z(n40590) );
  XNOR U37753 ( .A(n40592), .B(n40593), .Z(n37750) );
  AND U37754 ( .A(n40592), .B(n40594), .Z(n40593) );
  XNOR U37755 ( .A(n40595), .B(n40596), .Z(n37753) );
  AND U37756 ( .A(n40595), .B(n40597), .Z(n40596) );
  XNOR U37757 ( .A(n40598), .B(n40599), .Z(n37756) );
  AND U37758 ( .A(n40598), .B(n40600), .Z(n40599) );
  XNOR U37759 ( .A(n40601), .B(n40602), .Z(n37759) );
  AND U37760 ( .A(n40601), .B(n40603), .Z(n40602) );
  XNOR U37761 ( .A(n40604), .B(n40605), .Z(n37762) );
  AND U37762 ( .A(n40604), .B(n40606), .Z(n40605) );
  XNOR U37763 ( .A(n40607), .B(n40608), .Z(n37765) );
  AND U37764 ( .A(n40607), .B(n40609), .Z(n40608) );
  XNOR U37765 ( .A(n40610), .B(n40611), .Z(n37768) );
  AND U37766 ( .A(n40610), .B(n40612), .Z(n40611) );
  XNOR U37767 ( .A(n40613), .B(n40614), .Z(n37771) );
  AND U37768 ( .A(n40613), .B(n40615), .Z(n40614) );
  XNOR U37769 ( .A(n40616), .B(n40617), .Z(n37774) );
  AND U37770 ( .A(n40616), .B(n40618), .Z(n40617) );
  XNOR U37771 ( .A(n40619), .B(n40620), .Z(n37777) );
  AND U37772 ( .A(n40619), .B(n40621), .Z(n40620) );
  XNOR U37773 ( .A(n40622), .B(n40623), .Z(n37780) );
  AND U37774 ( .A(n40622), .B(n40624), .Z(n40623) );
  XNOR U37775 ( .A(n40625), .B(n40626), .Z(n37783) );
  AND U37776 ( .A(n40625), .B(n40627), .Z(n40626) );
  XNOR U37777 ( .A(n40628), .B(n40629), .Z(n37786) );
  AND U37778 ( .A(n40628), .B(n40630), .Z(n40629) );
  XNOR U37779 ( .A(n40631), .B(n40632), .Z(n37789) );
  AND U37780 ( .A(n40631), .B(n40633), .Z(n40632) );
  XNOR U37781 ( .A(n40634), .B(n40635), .Z(n37792) );
  AND U37782 ( .A(n40634), .B(n40636), .Z(n40635) );
  XNOR U37783 ( .A(n40637), .B(n40638), .Z(n37795) );
  AND U37784 ( .A(n40637), .B(n40639), .Z(n40638) );
  XNOR U37785 ( .A(n40640), .B(n40641), .Z(n37798) );
  AND U37786 ( .A(n40640), .B(n40642), .Z(n40641) );
  XNOR U37787 ( .A(n40643), .B(n40644), .Z(n37801) );
  AND U37788 ( .A(n40643), .B(n40645), .Z(n40644) );
  XNOR U37789 ( .A(n40646), .B(n40647), .Z(n37804) );
  AND U37790 ( .A(n40646), .B(n40648), .Z(n40647) );
  XNOR U37791 ( .A(n40649), .B(n40650), .Z(n37807) );
  AND U37792 ( .A(n40649), .B(n40651), .Z(n40650) );
  XNOR U37793 ( .A(n40652), .B(n40653), .Z(n37810) );
  AND U37794 ( .A(n40652), .B(n40654), .Z(n40653) );
  XNOR U37795 ( .A(n40655), .B(n40656), .Z(n37813) );
  AND U37796 ( .A(n40655), .B(n40657), .Z(n40656) );
  XNOR U37797 ( .A(n40658), .B(n40659), .Z(n37816) );
  AND U37798 ( .A(n40658), .B(n40660), .Z(n40659) );
  XNOR U37799 ( .A(n40661), .B(n40662), .Z(n37819) );
  AND U37800 ( .A(n40661), .B(n40663), .Z(n40662) );
  XNOR U37801 ( .A(n40664), .B(n40665), .Z(n37822) );
  AND U37802 ( .A(n40664), .B(n40666), .Z(n40665) );
  XNOR U37803 ( .A(n40667), .B(n40668), .Z(n37825) );
  AND U37804 ( .A(n40667), .B(n40669), .Z(n40668) );
  XNOR U37805 ( .A(n40670), .B(n40671), .Z(n37828) );
  AND U37806 ( .A(n40670), .B(n40672), .Z(n40671) );
  XNOR U37807 ( .A(n40673), .B(n40674), .Z(n37831) );
  AND U37808 ( .A(n40673), .B(n40675), .Z(n40674) );
  XNOR U37809 ( .A(n40676), .B(n40677), .Z(n37834) );
  AND U37810 ( .A(n40676), .B(n40678), .Z(n40677) );
  XNOR U37811 ( .A(n40679), .B(n40680), .Z(n37837) );
  AND U37812 ( .A(n40679), .B(n40681), .Z(n40680) );
  XNOR U37813 ( .A(n40682), .B(n40683), .Z(n37840) );
  AND U37814 ( .A(n40682), .B(n40684), .Z(n40683) );
  XNOR U37815 ( .A(n40685), .B(n40686), .Z(n37843) );
  AND U37816 ( .A(n40685), .B(n40687), .Z(n40686) );
  XNOR U37817 ( .A(n40688), .B(n40689), .Z(n37846) );
  AND U37818 ( .A(n40688), .B(n40690), .Z(n40689) );
  XNOR U37819 ( .A(n40691), .B(n40692), .Z(n37849) );
  AND U37820 ( .A(n40691), .B(n40693), .Z(n40692) );
  XNOR U37821 ( .A(n40694), .B(n40695), .Z(n37852) );
  AND U37822 ( .A(n40694), .B(n40696), .Z(n40695) );
  XNOR U37823 ( .A(n40697), .B(n40698), .Z(n37855) );
  AND U37824 ( .A(n40697), .B(n40699), .Z(n40698) );
  XNOR U37825 ( .A(n40700), .B(n40701), .Z(n37858) );
  AND U37826 ( .A(n40700), .B(n40702), .Z(n40701) );
  XNOR U37827 ( .A(n40703), .B(n40704), .Z(n37861) );
  AND U37828 ( .A(n40703), .B(n40705), .Z(n40704) );
  XNOR U37829 ( .A(n40706), .B(n40707), .Z(n37864) );
  AND U37830 ( .A(n40706), .B(n40708), .Z(n40707) );
  XNOR U37831 ( .A(n40709), .B(n40710), .Z(n37867) );
  AND U37832 ( .A(n40709), .B(n40711), .Z(n40710) );
  XNOR U37833 ( .A(n40712), .B(n40713), .Z(n37870) );
  AND U37834 ( .A(n40712), .B(n40714), .Z(n40713) );
  XNOR U37835 ( .A(n40715), .B(n40716), .Z(n37873) );
  AND U37836 ( .A(n40715), .B(n40717), .Z(n40716) );
  XNOR U37837 ( .A(n40718), .B(n40719), .Z(n37876) );
  AND U37838 ( .A(n40718), .B(n40720), .Z(n40719) );
  XNOR U37839 ( .A(n40721), .B(n40722), .Z(n37879) );
  AND U37840 ( .A(n40721), .B(n40723), .Z(n40722) );
  XNOR U37841 ( .A(n40724), .B(n40725), .Z(n37882) );
  AND U37842 ( .A(n40724), .B(n40726), .Z(n40725) );
  XNOR U37843 ( .A(n40727), .B(n40728), .Z(n37885) );
  AND U37844 ( .A(n40727), .B(n40729), .Z(n40728) );
  XNOR U37845 ( .A(n40730), .B(n40731), .Z(n37888) );
  AND U37846 ( .A(n40730), .B(n40732), .Z(n40731) );
  XNOR U37847 ( .A(n40733), .B(n40734), .Z(n37891) );
  AND U37848 ( .A(n40733), .B(n40735), .Z(n40734) );
  XNOR U37849 ( .A(n40736), .B(n40737), .Z(n37894) );
  AND U37850 ( .A(n40736), .B(n40738), .Z(n40737) );
  XNOR U37851 ( .A(n40739), .B(n40740), .Z(n37897) );
  AND U37852 ( .A(n40739), .B(n40741), .Z(n40740) );
  XNOR U37853 ( .A(n40742), .B(n40743), .Z(n37900) );
  AND U37854 ( .A(n40742), .B(n40744), .Z(n40743) );
  XNOR U37855 ( .A(n40745), .B(n40746), .Z(n37903) );
  AND U37856 ( .A(n40745), .B(n40747), .Z(n40746) );
  XNOR U37857 ( .A(n40748), .B(n40749), .Z(n37906) );
  AND U37858 ( .A(n40748), .B(n40750), .Z(n40749) );
  XNOR U37859 ( .A(n40751), .B(n40752), .Z(n37909) );
  AND U37860 ( .A(n40751), .B(n40753), .Z(n40752) );
  XNOR U37861 ( .A(n40754), .B(n40755), .Z(n37912) );
  AND U37862 ( .A(n40754), .B(n40756), .Z(n40755) );
  XNOR U37863 ( .A(n40757), .B(n40758), .Z(n37915) );
  AND U37864 ( .A(n40757), .B(n40759), .Z(n40758) );
  XNOR U37865 ( .A(n40760), .B(n40761), .Z(n37918) );
  AND U37866 ( .A(n40760), .B(n40762), .Z(n40761) );
  XNOR U37867 ( .A(n40763), .B(n40764), .Z(n37921) );
  AND U37868 ( .A(n40763), .B(n40765), .Z(n40764) );
  XNOR U37869 ( .A(n40766), .B(n40767), .Z(n37924) );
  AND U37870 ( .A(n40766), .B(n40768), .Z(n40767) );
  XNOR U37871 ( .A(n40769), .B(n40770), .Z(n37927) );
  AND U37872 ( .A(n40769), .B(n40771), .Z(n40770) );
  XNOR U37873 ( .A(n40772), .B(n40773), .Z(n37930) );
  AND U37874 ( .A(n40772), .B(n40774), .Z(n40773) );
  XNOR U37875 ( .A(n40775), .B(n40776), .Z(n37933) );
  AND U37876 ( .A(n40775), .B(n40777), .Z(n40776) );
  XNOR U37877 ( .A(n40778), .B(n40779), .Z(n37936) );
  AND U37878 ( .A(n40778), .B(n40780), .Z(n40779) );
  XNOR U37879 ( .A(n40781), .B(n40782), .Z(n37939) );
  AND U37880 ( .A(n40781), .B(n40783), .Z(n40782) );
  XNOR U37881 ( .A(n40784), .B(n40785), .Z(n37942) );
  AND U37882 ( .A(n40784), .B(n40786), .Z(n40785) );
  XNOR U37883 ( .A(n40787), .B(n40788), .Z(n37945) );
  AND U37884 ( .A(n40787), .B(n40789), .Z(n40788) );
  XNOR U37885 ( .A(n40790), .B(n40791), .Z(n37948) );
  AND U37886 ( .A(n40790), .B(n40792), .Z(n40791) );
  XNOR U37887 ( .A(n40793), .B(n40794), .Z(n37951) );
  AND U37888 ( .A(n40793), .B(n40795), .Z(n40794) );
  XNOR U37889 ( .A(n40796), .B(n40797), .Z(n37954) );
  AND U37890 ( .A(n40796), .B(n40798), .Z(n40797) );
  XNOR U37891 ( .A(n40799), .B(n40800), .Z(n37957) );
  AND U37892 ( .A(n40799), .B(n40801), .Z(n40800) );
  XNOR U37893 ( .A(n40802), .B(n40803), .Z(n37960) );
  AND U37894 ( .A(n40802), .B(n40804), .Z(n40803) );
  XNOR U37895 ( .A(n40805), .B(n40806), .Z(n37963) );
  AND U37896 ( .A(n40805), .B(n40807), .Z(n40806) );
  XNOR U37897 ( .A(n40808), .B(n40809), .Z(n37966) );
  AND U37898 ( .A(n40808), .B(n40810), .Z(n40809) );
  XNOR U37899 ( .A(n40811), .B(n40812), .Z(n37969) );
  AND U37900 ( .A(n40811), .B(n40813), .Z(n40812) );
  XNOR U37901 ( .A(n40814), .B(n40815), .Z(n37972) );
  AND U37902 ( .A(n40814), .B(n40816), .Z(n40815) );
  XNOR U37903 ( .A(n40817), .B(n40818), .Z(n37975) );
  AND U37904 ( .A(n40817), .B(n40819), .Z(n40818) );
  XNOR U37905 ( .A(n40820), .B(n40821), .Z(n37978) );
  AND U37906 ( .A(n40820), .B(n40822), .Z(n40821) );
  XNOR U37907 ( .A(n40823), .B(n40824), .Z(n37981) );
  AND U37908 ( .A(n40823), .B(n40825), .Z(n40824) );
  XNOR U37909 ( .A(n40826), .B(n40827), .Z(n37984) );
  AND U37910 ( .A(n40826), .B(n40828), .Z(n40827) );
  XNOR U37911 ( .A(n40829), .B(n40830), .Z(n37987) );
  AND U37912 ( .A(n40829), .B(n40831), .Z(n40830) );
  XNOR U37913 ( .A(n40832), .B(n40833), .Z(n37990) );
  AND U37914 ( .A(n40832), .B(n40834), .Z(n40833) );
  XNOR U37915 ( .A(n40835), .B(n40836), .Z(n37993) );
  AND U37916 ( .A(n40835), .B(n40837), .Z(n40836) );
  XNOR U37917 ( .A(n40838), .B(n40839), .Z(n37996) );
  AND U37918 ( .A(n40838), .B(n40840), .Z(n40839) );
  XNOR U37919 ( .A(n40841), .B(n40842), .Z(n37999) );
  AND U37920 ( .A(n40841), .B(n40843), .Z(n40842) );
  XNOR U37921 ( .A(n40844), .B(n40845), .Z(n38002) );
  AND U37922 ( .A(n40844), .B(n40846), .Z(n40845) );
  XNOR U37923 ( .A(n40847), .B(n40848), .Z(n38005) );
  AND U37924 ( .A(n40847), .B(n40849), .Z(n40848) );
  XNOR U37925 ( .A(n40850), .B(n40851), .Z(n38008) );
  AND U37926 ( .A(n40850), .B(n40852), .Z(n40851) );
  XNOR U37927 ( .A(n40853), .B(n40854), .Z(n38011) );
  AND U37928 ( .A(n40853), .B(n40855), .Z(n40854) );
  XNOR U37929 ( .A(n40856), .B(n40857), .Z(n38014) );
  AND U37930 ( .A(n40856), .B(n40858), .Z(n40857) );
  XNOR U37931 ( .A(n40859), .B(n40860), .Z(n38017) );
  AND U37932 ( .A(n40859), .B(n40861), .Z(n40860) );
  XNOR U37933 ( .A(n40862), .B(n40863), .Z(n38020) );
  AND U37934 ( .A(n40862), .B(n40864), .Z(n40863) );
  XNOR U37935 ( .A(n40865), .B(n40866), .Z(n38023) );
  AND U37936 ( .A(n40865), .B(n40867), .Z(n40866) );
  XNOR U37937 ( .A(n40868), .B(n40869), .Z(n38026) );
  AND U37938 ( .A(n40868), .B(n40870), .Z(n40869) );
  XNOR U37939 ( .A(n40871), .B(n40872), .Z(n38029) );
  AND U37940 ( .A(n40871), .B(n40873), .Z(n40872) );
  XNOR U37941 ( .A(n40874), .B(n40875), .Z(n38032) );
  AND U37942 ( .A(n40874), .B(n40876), .Z(n40875) );
  XNOR U37943 ( .A(n40877), .B(n40878), .Z(n38035) );
  AND U37944 ( .A(n40877), .B(n40879), .Z(n40878) );
  XNOR U37945 ( .A(n40880), .B(n40881), .Z(n38038) );
  AND U37946 ( .A(n40880), .B(n40882), .Z(n40881) );
  XNOR U37947 ( .A(n40883), .B(n40884), .Z(n38041) );
  AND U37948 ( .A(n40883), .B(n40885), .Z(n40884) );
  XNOR U37949 ( .A(n40886), .B(n40887), .Z(n38044) );
  AND U37950 ( .A(n40886), .B(n40888), .Z(n40887) );
  XNOR U37951 ( .A(n40889), .B(n40890), .Z(n38047) );
  AND U37952 ( .A(n40889), .B(n40891), .Z(n40890) );
  XNOR U37953 ( .A(n40892), .B(n40893), .Z(n38050) );
  AND U37954 ( .A(n40892), .B(n40894), .Z(n40893) );
  XNOR U37955 ( .A(n40895), .B(n40896), .Z(n38053) );
  AND U37956 ( .A(n40895), .B(n40897), .Z(n40896) );
  XNOR U37957 ( .A(n40898), .B(n40899), .Z(n38056) );
  AND U37958 ( .A(n40898), .B(n40900), .Z(n40899) );
  XNOR U37959 ( .A(n40901), .B(n40902), .Z(n38059) );
  AND U37960 ( .A(n40901), .B(n40903), .Z(n40902) );
  XNOR U37961 ( .A(n40904), .B(n40905), .Z(n38062) );
  AND U37962 ( .A(n40904), .B(n40906), .Z(n40905) );
  XNOR U37963 ( .A(n40907), .B(n40908), .Z(n38065) );
  AND U37964 ( .A(n40907), .B(n40909), .Z(n40908) );
  XNOR U37965 ( .A(n40910), .B(n40911), .Z(n38068) );
  AND U37966 ( .A(n40910), .B(n40912), .Z(n40911) );
  XNOR U37967 ( .A(n40913), .B(n40914), .Z(n38071) );
  AND U37968 ( .A(n40913), .B(n40915), .Z(n40914) );
  XNOR U37969 ( .A(n40916), .B(n40917), .Z(n38074) );
  AND U37970 ( .A(n40916), .B(n40918), .Z(n40917) );
  XNOR U37971 ( .A(n40919), .B(n40920), .Z(n38077) );
  AND U37972 ( .A(n40919), .B(n40921), .Z(n40920) );
  XNOR U37973 ( .A(n40922), .B(n40923), .Z(n38080) );
  AND U37974 ( .A(n40922), .B(n40924), .Z(n40923) );
  XNOR U37975 ( .A(n40925), .B(n40926), .Z(n38083) );
  AND U37976 ( .A(n40925), .B(n40927), .Z(n40926) );
  XNOR U37977 ( .A(n40928), .B(n40929), .Z(n38086) );
  AND U37978 ( .A(n40928), .B(n40930), .Z(n40929) );
  XNOR U37979 ( .A(n40931), .B(n40932), .Z(n38089) );
  AND U37980 ( .A(n40931), .B(n40933), .Z(n40932) );
  XNOR U37981 ( .A(n40934), .B(n40935), .Z(n38092) );
  AND U37982 ( .A(n40934), .B(n40936), .Z(n40935) );
  XNOR U37983 ( .A(n40937), .B(n40938), .Z(n38095) );
  AND U37984 ( .A(n40937), .B(n40939), .Z(n40938) );
  XNOR U37985 ( .A(n40940), .B(n40941), .Z(n38098) );
  AND U37986 ( .A(n40940), .B(n40942), .Z(n40941) );
  XNOR U37987 ( .A(n40943), .B(n40944), .Z(n38101) );
  AND U37988 ( .A(n40943), .B(n40945), .Z(n40944) );
  XNOR U37989 ( .A(n40946), .B(n40947), .Z(n38104) );
  AND U37990 ( .A(n40946), .B(n40948), .Z(n40947) );
  XNOR U37991 ( .A(n40949), .B(n40950), .Z(n38107) );
  AND U37992 ( .A(n40949), .B(n40951), .Z(n40950) );
  XNOR U37993 ( .A(n40952), .B(n40953), .Z(n38110) );
  AND U37994 ( .A(n40952), .B(n40954), .Z(n40953) );
  XNOR U37995 ( .A(n40955), .B(n40956), .Z(n38113) );
  AND U37996 ( .A(n40955), .B(n40957), .Z(n40956) );
  XNOR U37997 ( .A(n40958), .B(n40959), .Z(n38116) );
  AND U37998 ( .A(n40958), .B(n40960), .Z(n40959) );
  XNOR U37999 ( .A(n40961), .B(n40962), .Z(n38119) );
  AND U38000 ( .A(n40961), .B(n40963), .Z(n40962) );
  XNOR U38001 ( .A(n40964), .B(n40965), .Z(n38122) );
  AND U38002 ( .A(n40964), .B(n40966), .Z(n40965) );
  XNOR U38003 ( .A(n40967), .B(n40968), .Z(n38125) );
  AND U38004 ( .A(n40967), .B(n40969), .Z(n40968) );
  XNOR U38005 ( .A(n40970), .B(n40971), .Z(n38128) );
  AND U38006 ( .A(n40970), .B(n40972), .Z(n40971) );
  XNOR U38007 ( .A(n40973), .B(n40974), .Z(n38131) );
  AND U38008 ( .A(n40973), .B(n40975), .Z(n40974) );
  XNOR U38009 ( .A(n40976), .B(n40977), .Z(n38134) );
  AND U38010 ( .A(n40976), .B(n40978), .Z(n40977) );
  XNOR U38011 ( .A(n40979), .B(n40980), .Z(n38137) );
  AND U38012 ( .A(n40979), .B(n40981), .Z(n40980) );
  XNOR U38013 ( .A(n40982), .B(n40983), .Z(n38140) );
  AND U38014 ( .A(n40982), .B(n40984), .Z(n40983) );
  XNOR U38015 ( .A(n40985), .B(n40986), .Z(n38143) );
  AND U38016 ( .A(n40985), .B(n40987), .Z(n40986) );
  XNOR U38017 ( .A(n40988), .B(n40989), .Z(n38146) );
  AND U38018 ( .A(n40988), .B(n40990), .Z(n40989) );
  XNOR U38019 ( .A(n40991), .B(n40992), .Z(n38149) );
  AND U38020 ( .A(n40991), .B(n40993), .Z(n40992) );
  XNOR U38021 ( .A(n40994), .B(n40995), .Z(n38152) );
  AND U38022 ( .A(n40994), .B(n40996), .Z(n40995) );
  XNOR U38023 ( .A(n40997), .B(n40998), .Z(n38155) );
  AND U38024 ( .A(n40997), .B(n40999), .Z(n40998) );
  XNOR U38025 ( .A(n41000), .B(n41001), .Z(n38158) );
  AND U38026 ( .A(n41000), .B(n41002), .Z(n41001) );
  XNOR U38027 ( .A(n41003), .B(n41004), .Z(n38161) );
  AND U38028 ( .A(n41003), .B(n41005), .Z(n41004) );
  XNOR U38029 ( .A(n41006), .B(n41007), .Z(n38164) );
  AND U38030 ( .A(n41006), .B(n41008), .Z(n41007) );
  XNOR U38031 ( .A(n41009), .B(n41010), .Z(n38167) );
  AND U38032 ( .A(n41009), .B(n41011), .Z(n41010) );
  XNOR U38033 ( .A(n41012), .B(n41013), .Z(n38170) );
  AND U38034 ( .A(n41012), .B(n41014), .Z(n41013) );
  XNOR U38035 ( .A(n41015), .B(n41016), .Z(n38173) );
  AND U38036 ( .A(n41015), .B(n41017), .Z(n41016) );
  XNOR U38037 ( .A(n41018), .B(n41019), .Z(n38176) );
  AND U38038 ( .A(n41018), .B(n41020), .Z(n41019) );
  XNOR U38039 ( .A(n41021), .B(n41022), .Z(n38179) );
  AND U38040 ( .A(n41021), .B(n41023), .Z(n41022) );
  XNOR U38041 ( .A(n41024), .B(n41025), .Z(n38182) );
  AND U38042 ( .A(n41024), .B(n41026), .Z(n41025) );
  XNOR U38043 ( .A(n41027), .B(n41028), .Z(n38185) );
  AND U38044 ( .A(n41027), .B(n41029), .Z(n41028) );
  XNOR U38045 ( .A(n41030), .B(n41031), .Z(n38188) );
  AND U38046 ( .A(n41030), .B(n41032), .Z(n41031) );
  XNOR U38047 ( .A(n41033), .B(n41034), .Z(n38191) );
  AND U38048 ( .A(n41033), .B(n41035), .Z(n41034) );
  XNOR U38049 ( .A(n41036), .B(n41037), .Z(n38194) );
  AND U38050 ( .A(n41036), .B(n41038), .Z(n41037) );
  XNOR U38051 ( .A(n41039), .B(n41040), .Z(n38197) );
  AND U38052 ( .A(n41039), .B(n41041), .Z(n41040) );
  XNOR U38053 ( .A(n41042), .B(n41043), .Z(n38200) );
  AND U38054 ( .A(n41042), .B(n41044), .Z(n41043) );
  XNOR U38055 ( .A(n41045), .B(n41046), .Z(n38203) );
  AND U38056 ( .A(n41045), .B(n41047), .Z(n41046) );
  XNOR U38057 ( .A(n41048), .B(n41049), .Z(n38206) );
  AND U38058 ( .A(n41048), .B(n41050), .Z(n41049) );
  XNOR U38059 ( .A(n41051), .B(n41052), .Z(n38209) );
  AND U38060 ( .A(n41051), .B(n41053), .Z(n41052) );
  XNOR U38061 ( .A(n41054), .B(n41055), .Z(n38212) );
  AND U38062 ( .A(n41054), .B(n41056), .Z(n41055) );
  XNOR U38063 ( .A(n41057), .B(n41058), .Z(n38215) );
  AND U38064 ( .A(n41057), .B(n41059), .Z(n41058) );
  XNOR U38065 ( .A(n41060), .B(n41061), .Z(n38218) );
  AND U38066 ( .A(n41060), .B(n41062), .Z(n41061) );
  XNOR U38067 ( .A(n41063), .B(n41064), .Z(n38221) );
  AND U38068 ( .A(n41063), .B(n41065), .Z(n41064) );
  XNOR U38069 ( .A(n41066), .B(n41067), .Z(n38224) );
  AND U38070 ( .A(n41066), .B(n41068), .Z(n41067) );
  XNOR U38071 ( .A(n41069), .B(n41070), .Z(n38227) );
  AND U38072 ( .A(n41069), .B(n41071), .Z(n41070) );
  XNOR U38073 ( .A(n41072), .B(n41073), .Z(n38230) );
  AND U38074 ( .A(n41072), .B(n41074), .Z(n41073) );
  XNOR U38075 ( .A(n41075), .B(n41076), .Z(n38233) );
  AND U38076 ( .A(n41075), .B(n41077), .Z(n41076) );
  XNOR U38077 ( .A(n41078), .B(n41079), .Z(n38236) );
  AND U38078 ( .A(n41078), .B(n41080), .Z(n41079) );
  XNOR U38079 ( .A(n41081), .B(n41082), .Z(n38239) );
  AND U38080 ( .A(n41081), .B(n41083), .Z(n41082) );
  XNOR U38081 ( .A(n41084), .B(n41085), .Z(n38242) );
  AND U38082 ( .A(n41084), .B(n41086), .Z(n41085) );
  XNOR U38083 ( .A(n41087), .B(n41088), .Z(n38245) );
  AND U38084 ( .A(n41087), .B(n41089), .Z(n41088) );
  XNOR U38085 ( .A(n41090), .B(n41091), .Z(n38248) );
  AND U38086 ( .A(n41090), .B(n41092), .Z(n41091) );
  XNOR U38087 ( .A(n41093), .B(n41094), .Z(n38251) );
  AND U38088 ( .A(n41093), .B(n41095), .Z(n41094) );
  XNOR U38089 ( .A(n41096), .B(n41097), .Z(n38254) );
  AND U38090 ( .A(n41096), .B(n41098), .Z(n41097) );
  XNOR U38091 ( .A(n41099), .B(n41100), .Z(n38257) );
  AND U38092 ( .A(n41099), .B(n41101), .Z(n41100) );
  XNOR U38093 ( .A(n41102), .B(n41103), .Z(n38260) );
  AND U38094 ( .A(n41102), .B(n41104), .Z(n41103) );
  XNOR U38095 ( .A(n41105), .B(n41106), .Z(n38263) );
  AND U38096 ( .A(n41105), .B(n41107), .Z(n41106) );
  XNOR U38097 ( .A(n41108), .B(n41109), .Z(n38266) );
  AND U38098 ( .A(n41108), .B(n41110), .Z(n41109) );
  XNOR U38099 ( .A(n41111), .B(n41112), .Z(n38269) );
  AND U38100 ( .A(n41111), .B(n41113), .Z(n41112) );
  XNOR U38101 ( .A(n41114), .B(n41115), .Z(n38272) );
  AND U38102 ( .A(n41114), .B(n41116), .Z(n41115) );
  XNOR U38103 ( .A(n41117), .B(n41118), .Z(n38275) );
  AND U38104 ( .A(n41117), .B(n41119), .Z(n41118) );
  XNOR U38105 ( .A(n41120), .B(n41121), .Z(n38278) );
  AND U38106 ( .A(n41120), .B(n41122), .Z(n41121) );
  XNOR U38107 ( .A(n41123), .B(n41124), .Z(n38281) );
  AND U38108 ( .A(n41123), .B(n41125), .Z(n41124) );
  XNOR U38109 ( .A(n41126), .B(n41127), .Z(n38284) );
  AND U38110 ( .A(n41126), .B(n41128), .Z(n41127) );
  XNOR U38111 ( .A(n41129), .B(n41130), .Z(n38287) );
  AND U38112 ( .A(n41129), .B(n41131), .Z(n41130) );
  XNOR U38113 ( .A(n41132), .B(n41133), .Z(n38290) );
  AND U38114 ( .A(n41132), .B(n41134), .Z(n41133) );
  XNOR U38115 ( .A(n41135), .B(n41136), .Z(n38293) );
  AND U38116 ( .A(n41135), .B(n41137), .Z(n41136) );
  XNOR U38117 ( .A(n41138), .B(n41139), .Z(n38296) );
  AND U38118 ( .A(n41138), .B(n41140), .Z(n41139) );
  XNOR U38119 ( .A(n41141), .B(n41142), .Z(n38299) );
  AND U38120 ( .A(n41141), .B(n41143), .Z(n41142) );
  XNOR U38121 ( .A(n41144), .B(n41145), .Z(n38302) );
  AND U38122 ( .A(n41144), .B(n41146), .Z(n41145) );
  XNOR U38123 ( .A(n41147), .B(n41148), .Z(n38305) );
  AND U38124 ( .A(n41147), .B(n41149), .Z(n41148) );
  XNOR U38125 ( .A(n41150), .B(n41151), .Z(n38308) );
  AND U38126 ( .A(n41150), .B(n41152), .Z(n41151) );
  XNOR U38127 ( .A(n41153), .B(n41154), .Z(n38311) );
  AND U38128 ( .A(n41153), .B(n41155), .Z(n41154) );
  XNOR U38129 ( .A(n41156), .B(n41157), .Z(n38314) );
  AND U38130 ( .A(n41156), .B(n41158), .Z(n41157) );
  XNOR U38131 ( .A(n41159), .B(n41160), .Z(n38317) );
  AND U38132 ( .A(n41159), .B(n41161), .Z(n41160) );
  XNOR U38133 ( .A(n41162), .B(n41163), .Z(n38320) );
  AND U38134 ( .A(n41162), .B(n41164), .Z(n41163) );
  XNOR U38135 ( .A(n41165), .B(n41166), .Z(n38323) );
  AND U38136 ( .A(n41165), .B(n41167), .Z(n41166) );
  XNOR U38137 ( .A(n41168), .B(n41169), .Z(n38326) );
  AND U38138 ( .A(n41168), .B(n41170), .Z(n41169) );
  XNOR U38139 ( .A(n41171), .B(n41172), .Z(n38329) );
  AND U38140 ( .A(n41171), .B(n41173), .Z(n41172) );
  XNOR U38141 ( .A(n41174), .B(n41175), .Z(n38332) );
  AND U38142 ( .A(n41174), .B(n41176), .Z(n41175) );
  XNOR U38143 ( .A(n41177), .B(n41178), .Z(n38335) );
  AND U38144 ( .A(n41177), .B(n41179), .Z(n41178) );
  XNOR U38145 ( .A(n41180), .B(n41181), .Z(n38338) );
  AND U38146 ( .A(n41180), .B(n41182), .Z(n41181) );
  XNOR U38147 ( .A(n41183), .B(n41184), .Z(n38341) );
  AND U38148 ( .A(n41183), .B(n41185), .Z(n41184) );
  XNOR U38149 ( .A(n41186), .B(n41187), .Z(n38344) );
  AND U38150 ( .A(n41186), .B(n41188), .Z(n41187) );
  XNOR U38151 ( .A(n41189), .B(n41190), .Z(n38347) );
  AND U38152 ( .A(n41189), .B(n41191), .Z(n41190) );
  XNOR U38153 ( .A(n41192), .B(n41193), .Z(n38350) );
  AND U38154 ( .A(n41192), .B(n41194), .Z(n41193) );
  XNOR U38155 ( .A(n41195), .B(n41196), .Z(n38353) );
  AND U38156 ( .A(n41195), .B(n41197), .Z(n41196) );
  XNOR U38157 ( .A(n41198), .B(n41199), .Z(n38356) );
  AND U38158 ( .A(n41198), .B(n41200), .Z(n41199) );
  XNOR U38159 ( .A(n41201), .B(n41202), .Z(n38359) );
  AND U38160 ( .A(n41201), .B(n41203), .Z(n41202) );
  XNOR U38161 ( .A(n41204), .B(n41205), .Z(n38362) );
  AND U38162 ( .A(n41204), .B(n41206), .Z(n41205) );
  XNOR U38163 ( .A(n41207), .B(n41208), .Z(n38365) );
  AND U38164 ( .A(n41207), .B(n41209), .Z(n41208) );
  XNOR U38165 ( .A(n41210), .B(n41211), .Z(n38368) );
  AND U38166 ( .A(n41210), .B(n41212), .Z(n41211) );
  XNOR U38167 ( .A(n41213), .B(n41214), .Z(n38371) );
  AND U38168 ( .A(n41213), .B(n41215), .Z(n41214) );
  XNOR U38169 ( .A(n41216), .B(n41217), .Z(n38374) );
  AND U38170 ( .A(n41216), .B(n41218), .Z(n41217) );
  XNOR U38171 ( .A(n41219), .B(n41220), .Z(n38377) );
  AND U38172 ( .A(n41219), .B(n41221), .Z(n41220) );
  XNOR U38173 ( .A(n41222), .B(n41223), .Z(n38380) );
  AND U38174 ( .A(n41222), .B(n41224), .Z(n41223) );
  XNOR U38175 ( .A(n41225), .B(n41226), .Z(n38383) );
  AND U38176 ( .A(n41225), .B(n41227), .Z(n41226) );
  XOR U38177 ( .A(n41228), .B(n41229), .Z(n38386) );
  AND U38178 ( .A(n41228), .B(n139), .Z(n41229) );
  XOR U38179 ( .A(n121), .B(n39809), .Z(n39811) );
  XOR U38180 ( .A(n39806), .B(n39805), .Z(n121) );
  XNOR U38181 ( .A(n39803), .B(n39802), .Z(n39805) );
  XNOR U38182 ( .A(n39800), .B(n39799), .Z(n39802) );
  XNOR U38183 ( .A(n39797), .B(n39796), .Z(n39799) );
  XNOR U38184 ( .A(n39794), .B(n39793), .Z(n39796) );
  XNOR U38185 ( .A(n39791), .B(n39790), .Z(n39793) );
  XNOR U38186 ( .A(n39788), .B(n39787), .Z(n39790) );
  XNOR U38187 ( .A(n39785), .B(n39784), .Z(n39787) );
  XNOR U38188 ( .A(n39782), .B(n39781), .Z(n39784) );
  XNOR U38189 ( .A(n39779), .B(n39778), .Z(n39781) );
  XNOR U38190 ( .A(n39776), .B(n39775), .Z(n39778) );
  XNOR U38191 ( .A(n39773), .B(n39772), .Z(n39775) );
  XNOR U38192 ( .A(n39770), .B(n39769), .Z(n39772) );
  XNOR U38193 ( .A(n39767), .B(n39766), .Z(n39769) );
  XNOR U38194 ( .A(n39764), .B(n39763), .Z(n39766) );
  XNOR U38195 ( .A(n39761), .B(n39760), .Z(n39763) );
  XNOR U38196 ( .A(n39758), .B(n39757), .Z(n39760) );
  XNOR U38197 ( .A(n39755), .B(n39754), .Z(n39757) );
  XNOR U38198 ( .A(n39752), .B(n39751), .Z(n39754) );
  XNOR U38199 ( .A(n39749), .B(n39748), .Z(n39751) );
  XNOR U38200 ( .A(n39746), .B(n39745), .Z(n39748) );
  XNOR U38201 ( .A(n39743), .B(n39742), .Z(n39745) );
  XNOR U38202 ( .A(n39740), .B(n39739), .Z(n39742) );
  XNOR U38203 ( .A(n39737), .B(n39736), .Z(n39739) );
  XNOR U38204 ( .A(n39734), .B(n39733), .Z(n39736) );
  XNOR U38205 ( .A(n39731), .B(n39730), .Z(n39733) );
  XNOR U38206 ( .A(n39728), .B(n39727), .Z(n39730) );
  XNOR U38207 ( .A(n39725), .B(n39724), .Z(n39727) );
  XNOR U38208 ( .A(n39722), .B(n39721), .Z(n39724) );
  XNOR U38209 ( .A(n39719), .B(n39718), .Z(n39721) );
  XNOR U38210 ( .A(n39716), .B(n39715), .Z(n39718) );
  XNOR U38211 ( .A(n39713), .B(n39712), .Z(n39715) );
  XNOR U38212 ( .A(n39710), .B(n39709), .Z(n39712) );
  XNOR U38213 ( .A(n39707), .B(n39706), .Z(n39709) );
  XNOR U38214 ( .A(n39704), .B(n39703), .Z(n39706) );
  XNOR U38215 ( .A(n39701), .B(n39700), .Z(n39703) );
  XNOR U38216 ( .A(n39698), .B(n39697), .Z(n39700) );
  XNOR U38217 ( .A(n39695), .B(n39694), .Z(n39697) );
  XNOR U38218 ( .A(n39692), .B(n39691), .Z(n39694) );
  XNOR U38219 ( .A(n39689), .B(n39688), .Z(n39691) );
  XNOR U38220 ( .A(n39686), .B(n39685), .Z(n39688) );
  XNOR U38221 ( .A(n39683), .B(n39682), .Z(n39685) );
  XNOR U38222 ( .A(n39680), .B(n39679), .Z(n39682) );
  XNOR U38223 ( .A(n39677), .B(n39676), .Z(n39679) );
  XNOR U38224 ( .A(n39674), .B(n39673), .Z(n39676) );
  XNOR U38225 ( .A(n39671), .B(n39670), .Z(n39673) );
  XNOR U38226 ( .A(n39668), .B(n39667), .Z(n39670) );
  XNOR U38227 ( .A(n39665), .B(n39664), .Z(n39667) );
  XNOR U38228 ( .A(n39662), .B(n39661), .Z(n39664) );
  XNOR U38229 ( .A(n39659), .B(n39658), .Z(n39661) );
  XNOR U38230 ( .A(n39656), .B(n39655), .Z(n39658) );
  XNOR U38231 ( .A(n39653), .B(n39652), .Z(n39655) );
  XNOR U38232 ( .A(n39650), .B(n39649), .Z(n39652) );
  XNOR U38233 ( .A(n39647), .B(n39646), .Z(n39649) );
  XNOR U38234 ( .A(n39644), .B(n39643), .Z(n39646) );
  XNOR U38235 ( .A(n39641), .B(n39640), .Z(n39643) );
  XNOR U38236 ( .A(n39638), .B(n39637), .Z(n39640) );
  XNOR U38237 ( .A(n39635), .B(n39634), .Z(n39637) );
  XNOR U38238 ( .A(n39632), .B(n39631), .Z(n39634) );
  XNOR U38239 ( .A(n39629), .B(n39628), .Z(n39631) );
  XNOR U38240 ( .A(n39626), .B(n39625), .Z(n39628) );
  XNOR U38241 ( .A(n39623), .B(n39622), .Z(n39625) );
  XNOR U38242 ( .A(n39620), .B(n39619), .Z(n39622) );
  XNOR U38243 ( .A(n39617), .B(n39616), .Z(n39619) );
  XNOR U38244 ( .A(n39614), .B(n39613), .Z(n39616) );
  XNOR U38245 ( .A(n39611), .B(n39610), .Z(n39613) );
  XNOR U38246 ( .A(n39608), .B(n39607), .Z(n39610) );
  XNOR U38247 ( .A(n39605), .B(n39604), .Z(n39607) );
  XNOR U38248 ( .A(n39602), .B(n39601), .Z(n39604) );
  XNOR U38249 ( .A(n39599), .B(n39598), .Z(n39601) );
  XNOR U38250 ( .A(n39596), .B(n39595), .Z(n39598) );
  XNOR U38251 ( .A(n39593), .B(n39592), .Z(n39595) );
  XNOR U38252 ( .A(n39590), .B(n39589), .Z(n39592) );
  XNOR U38253 ( .A(n39587), .B(n39586), .Z(n39589) );
  XNOR U38254 ( .A(n39584), .B(n39583), .Z(n39586) );
  XNOR U38255 ( .A(n39581), .B(n39580), .Z(n39583) );
  XNOR U38256 ( .A(n39578), .B(n39577), .Z(n39580) );
  XNOR U38257 ( .A(n39575), .B(n39574), .Z(n39577) );
  XNOR U38258 ( .A(n39572), .B(n39571), .Z(n39574) );
  XNOR U38259 ( .A(n39569), .B(n39568), .Z(n39571) );
  XNOR U38260 ( .A(n39566), .B(n39565), .Z(n39568) );
  XNOR U38261 ( .A(n39563), .B(n39562), .Z(n39565) );
  XNOR U38262 ( .A(n39560), .B(n39559), .Z(n39562) );
  XNOR U38263 ( .A(n39557), .B(n39556), .Z(n39559) );
  XNOR U38264 ( .A(n39554), .B(n39553), .Z(n39556) );
  XNOR U38265 ( .A(n39551), .B(n39550), .Z(n39553) );
  XNOR U38266 ( .A(n39548), .B(n39547), .Z(n39550) );
  XNOR U38267 ( .A(n39545), .B(n39544), .Z(n39547) );
  XNOR U38268 ( .A(n39542), .B(n39541), .Z(n39544) );
  XNOR U38269 ( .A(n39539), .B(n39538), .Z(n39541) );
  XNOR U38270 ( .A(n39536), .B(n39535), .Z(n39538) );
  XNOR U38271 ( .A(n39533), .B(n39532), .Z(n39535) );
  XNOR U38272 ( .A(n39530), .B(n39529), .Z(n39532) );
  XNOR U38273 ( .A(n39527), .B(n39526), .Z(n39529) );
  XNOR U38274 ( .A(n39524), .B(n39523), .Z(n39526) );
  XNOR U38275 ( .A(n39521), .B(n39520), .Z(n39523) );
  XNOR U38276 ( .A(n39518), .B(n39517), .Z(n39520) );
  XNOR U38277 ( .A(n39515), .B(n39514), .Z(n39517) );
  XNOR U38278 ( .A(n39512), .B(n39511), .Z(n39514) );
  XNOR U38279 ( .A(n39509), .B(n39508), .Z(n39511) );
  XNOR U38280 ( .A(n39506), .B(n39505), .Z(n39508) );
  XNOR U38281 ( .A(n39503), .B(n39502), .Z(n39505) );
  XNOR U38282 ( .A(n39500), .B(n39499), .Z(n39502) );
  XNOR U38283 ( .A(n39497), .B(n39496), .Z(n39499) );
  XNOR U38284 ( .A(n39494), .B(n39493), .Z(n39496) );
  XNOR U38285 ( .A(n39491), .B(n39490), .Z(n39493) );
  XNOR U38286 ( .A(n39488), .B(n39487), .Z(n39490) );
  XNOR U38287 ( .A(n39485), .B(n39484), .Z(n39487) );
  XNOR U38288 ( .A(n39482), .B(n39481), .Z(n39484) );
  XNOR U38289 ( .A(n39479), .B(n39478), .Z(n39481) );
  XNOR U38290 ( .A(n39476), .B(n39475), .Z(n39478) );
  XNOR U38291 ( .A(n39473), .B(n39472), .Z(n39475) );
  XNOR U38292 ( .A(n39470), .B(n39469), .Z(n39472) );
  XNOR U38293 ( .A(n39467), .B(n39466), .Z(n39469) );
  XNOR U38294 ( .A(n39464), .B(n39463), .Z(n39466) );
  XNOR U38295 ( .A(n39461), .B(n39460), .Z(n39463) );
  XNOR U38296 ( .A(n39458), .B(n39457), .Z(n39460) );
  XNOR U38297 ( .A(n39455), .B(n39454), .Z(n39457) );
  XNOR U38298 ( .A(n39452), .B(n39451), .Z(n39454) );
  XNOR U38299 ( .A(n39449), .B(n39448), .Z(n39451) );
  XNOR U38300 ( .A(n39446), .B(n39445), .Z(n39448) );
  XNOR U38301 ( .A(n39443), .B(n39442), .Z(n39445) );
  XNOR U38302 ( .A(n39440), .B(n39439), .Z(n39442) );
  XNOR U38303 ( .A(n39437), .B(n39436), .Z(n39439) );
  XNOR U38304 ( .A(n39434), .B(n39433), .Z(n39436) );
  XNOR U38305 ( .A(n39431), .B(n39430), .Z(n39433) );
  XNOR U38306 ( .A(n39428), .B(n39427), .Z(n39430) );
  XNOR U38307 ( .A(n39425), .B(n39424), .Z(n39427) );
  XNOR U38308 ( .A(n39422), .B(n39421), .Z(n39424) );
  XNOR U38309 ( .A(n39419), .B(n39418), .Z(n39421) );
  XNOR U38310 ( .A(n39416), .B(n39415), .Z(n39418) );
  XNOR U38311 ( .A(n39413), .B(n39412), .Z(n39415) );
  XNOR U38312 ( .A(n39410), .B(n39409), .Z(n39412) );
  XNOR U38313 ( .A(n39407), .B(n39406), .Z(n39409) );
  XNOR U38314 ( .A(n39404), .B(n39403), .Z(n39406) );
  XNOR U38315 ( .A(n39401), .B(n39400), .Z(n39403) );
  XNOR U38316 ( .A(n39398), .B(n39397), .Z(n39400) );
  XNOR U38317 ( .A(n39395), .B(n39394), .Z(n39397) );
  XNOR U38318 ( .A(n39392), .B(n39391), .Z(n39394) );
  XNOR U38319 ( .A(n39389), .B(n39388), .Z(n39391) );
  XNOR U38320 ( .A(n39386), .B(n39385), .Z(n39388) );
  XNOR U38321 ( .A(n39383), .B(n39382), .Z(n39385) );
  XNOR U38322 ( .A(n39380), .B(n39379), .Z(n39382) );
  XNOR U38323 ( .A(n39377), .B(n39376), .Z(n39379) );
  XNOR U38324 ( .A(n39374), .B(n39373), .Z(n39376) );
  XNOR U38325 ( .A(n39371), .B(n39370), .Z(n39373) );
  XNOR U38326 ( .A(n39368), .B(n39367), .Z(n39370) );
  XNOR U38327 ( .A(n39365), .B(n39364), .Z(n39367) );
  XNOR U38328 ( .A(n39362), .B(n39361), .Z(n39364) );
  XNOR U38329 ( .A(n39359), .B(n39358), .Z(n39361) );
  XNOR U38330 ( .A(n39356), .B(n39355), .Z(n39358) );
  XNOR U38331 ( .A(n39353), .B(n39352), .Z(n39355) );
  XNOR U38332 ( .A(n39350), .B(n39349), .Z(n39352) );
  XNOR U38333 ( .A(n39347), .B(n39346), .Z(n39349) );
  XNOR U38334 ( .A(n39344), .B(n39343), .Z(n39346) );
  XNOR U38335 ( .A(n39341), .B(n39340), .Z(n39343) );
  XNOR U38336 ( .A(n39338), .B(n39337), .Z(n39340) );
  XNOR U38337 ( .A(n39335), .B(n39334), .Z(n39337) );
  XNOR U38338 ( .A(n39332), .B(n39331), .Z(n39334) );
  XNOR U38339 ( .A(n39329), .B(n39328), .Z(n39331) );
  XNOR U38340 ( .A(n39326), .B(n39325), .Z(n39328) );
  XNOR U38341 ( .A(n39323), .B(n39322), .Z(n39325) );
  XNOR U38342 ( .A(n39320), .B(n39319), .Z(n39322) );
  XNOR U38343 ( .A(n39317), .B(n39316), .Z(n39319) );
  XNOR U38344 ( .A(n39314), .B(n39313), .Z(n39316) );
  XNOR U38345 ( .A(n39311), .B(n39310), .Z(n39313) );
  XNOR U38346 ( .A(n39308), .B(n39307), .Z(n39310) );
  XNOR U38347 ( .A(n39305), .B(n39304), .Z(n39307) );
  XNOR U38348 ( .A(n39302), .B(n39301), .Z(n39304) );
  XNOR U38349 ( .A(n39299), .B(n39298), .Z(n39301) );
  XNOR U38350 ( .A(n39296), .B(n39295), .Z(n39298) );
  XNOR U38351 ( .A(n39293), .B(n39292), .Z(n39295) );
  XNOR U38352 ( .A(n39290), .B(n39289), .Z(n39292) );
  XNOR U38353 ( .A(n39287), .B(n39286), .Z(n39289) );
  XNOR U38354 ( .A(n39284), .B(n39283), .Z(n39286) );
  XNOR U38355 ( .A(n39281), .B(n39280), .Z(n39283) );
  XNOR U38356 ( .A(n39278), .B(n39277), .Z(n39280) );
  XNOR U38357 ( .A(n39275), .B(n39274), .Z(n39277) );
  XNOR U38358 ( .A(n39272), .B(n39271), .Z(n39274) );
  XNOR U38359 ( .A(n39269), .B(n39268), .Z(n39271) );
  XNOR U38360 ( .A(n39266), .B(n39265), .Z(n39268) );
  XNOR U38361 ( .A(n39263), .B(n39262), .Z(n39265) );
  XNOR U38362 ( .A(n39260), .B(n39259), .Z(n39262) );
  XNOR U38363 ( .A(n39257), .B(n39256), .Z(n39259) );
  XNOR U38364 ( .A(n39254), .B(n39253), .Z(n39256) );
  XNOR U38365 ( .A(n39251), .B(n39250), .Z(n39253) );
  XNOR U38366 ( .A(n39248), .B(n39247), .Z(n39250) );
  XNOR U38367 ( .A(n39245), .B(n39244), .Z(n39247) );
  XNOR U38368 ( .A(n39242), .B(n39241), .Z(n39244) );
  XNOR U38369 ( .A(n39239), .B(n39238), .Z(n39241) );
  XNOR U38370 ( .A(n39236), .B(n39235), .Z(n39238) );
  XNOR U38371 ( .A(n39233), .B(n39232), .Z(n39235) );
  XNOR U38372 ( .A(n39230), .B(n39229), .Z(n39232) );
  XNOR U38373 ( .A(n39227), .B(n39226), .Z(n39229) );
  XNOR U38374 ( .A(n39224), .B(n39223), .Z(n39226) );
  XNOR U38375 ( .A(n39221), .B(n39220), .Z(n39223) );
  XNOR U38376 ( .A(n39218), .B(n39217), .Z(n39220) );
  XNOR U38377 ( .A(n39215), .B(n39214), .Z(n39217) );
  XNOR U38378 ( .A(n39212), .B(n39211), .Z(n39214) );
  XNOR U38379 ( .A(n39209), .B(n39208), .Z(n39211) );
  XNOR U38380 ( .A(n39206), .B(n39205), .Z(n39208) );
  XNOR U38381 ( .A(n39203), .B(n39202), .Z(n39205) );
  XNOR U38382 ( .A(n39200), .B(n39199), .Z(n39202) );
  XNOR U38383 ( .A(n39197), .B(n39196), .Z(n39199) );
  XNOR U38384 ( .A(n39194), .B(n39193), .Z(n39196) );
  XNOR U38385 ( .A(n39191), .B(n39190), .Z(n39193) );
  XNOR U38386 ( .A(n39188), .B(n39187), .Z(n39190) );
  XNOR U38387 ( .A(n39185), .B(n39184), .Z(n39187) );
  XNOR U38388 ( .A(n39182), .B(n39181), .Z(n39184) );
  XNOR U38389 ( .A(n39179), .B(n39178), .Z(n39181) );
  XNOR U38390 ( .A(n39176), .B(n39175), .Z(n39178) );
  XNOR U38391 ( .A(n39173), .B(n39172), .Z(n39175) );
  XNOR U38392 ( .A(n39170), .B(n39169), .Z(n39172) );
  XNOR U38393 ( .A(n39167), .B(n39166), .Z(n39169) );
  XNOR U38394 ( .A(n39164), .B(n39163), .Z(n39166) );
  XNOR U38395 ( .A(n39161), .B(n39160), .Z(n39163) );
  XNOR U38396 ( .A(n39158), .B(n39157), .Z(n39160) );
  XNOR U38397 ( .A(n39155), .B(n39154), .Z(n39157) );
  XNOR U38398 ( .A(n39152), .B(n39151), .Z(n39154) );
  XNOR U38399 ( .A(n39149), .B(n39148), .Z(n39151) );
  XNOR U38400 ( .A(n39146), .B(n39145), .Z(n39148) );
  XNOR U38401 ( .A(n39143), .B(n39142), .Z(n39145) );
  XNOR U38402 ( .A(n39140), .B(n39139), .Z(n39142) );
  XNOR U38403 ( .A(n39137), .B(n39136), .Z(n39139) );
  XNOR U38404 ( .A(n39134), .B(n39133), .Z(n39136) );
  XNOR U38405 ( .A(n39131), .B(n39130), .Z(n39133) );
  XNOR U38406 ( .A(n39128), .B(n39127), .Z(n39130) );
  XNOR U38407 ( .A(n39125), .B(n39124), .Z(n39127) );
  XNOR U38408 ( .A(n39122), .B(n39121), .Z(n39124) );
  XNOR U38409 ( .A(n39119), .B(n39118), .Z(n39121) );
  XNOR U38410 ( .A(n39116), .B(n39115), .Z(n39118) );
  XNOR U38411 ( .A(n39113), .B(n39112), .Z(n39115) );
  XNOR U38412 ( .A(n39110), .B(n39109), .Z(n39112) );
  XNOR U38413 ( .A(n39107), .B(n39106), .Z(n39109) );
  XNOR U38414 ( .A(n39104), .B(n39103), .Z(n39106) );
  XNOR U38415 ( .A(n39101), .B(n39100), .Z(n39103) );
  XNOR U38416 ( .A(n39098), .B(n39097), .Z(n39100) );
  XNOR U38417 ( .A(n39095), .B(n39094), .Z(n39097) );
  XNOR U38418 ( .A(n39092), .B(n39091), .Z(n39094) );
  XNOR U38419 ( .A(n39089), .B(n39088), .Z(n39091) );
  XNOR U38420 ( .A(n39086), .B(n39085), .Z(n39088) );
  XNOR U38421 ( .A(n39083), .B(n39082), .Z(n39085) );
  XNOR U38422 ( .A(n39080), .B(n39079), .Z(n39082) );
  XNOR U38423 ( .A(n39077), .B(n39076), .Z(n39079) );
  XNOR U38424 ( .A(n39074), .B(n39073), .Z(n39076) );
  XNOR U38425 ( .A(n39071), .B(n39070), .Z(n39073) );
  XNOR U38426 ( .A(n39068), .B(n39067), .Z(n39070) );
  XNOR U38427 ( .A(n39065), .B(n39064), .Z(n39067) );
  XNOR U38428 ( .A(n39062), .B(n39061), .Z(n39064) );
  XNOR U38429 ( .A(n39059), .B(n39058), .Z(n39061) );
  XNOR U38430 ( .A(n39056), .B(n39055), .Z(n39058) );
  XNOR U38431 ( .A(n39053), .B(n39052), .Z(n39055) );
  XNOR U38432 ( .A(n39050), .B(n39049), .Z(n39052) );
  XNOR U38433 ( .A(n39047), .B(n39046), .Z(n39049) );
  XNOR U38434 ( .A(n39044), .B(n39043), .Z(n39046) );
  XNOR U38435 ( .A(n39041), .B(n39040), .Z(n39043) );
  XNOR U38436 ( .A(n39038), .B(n39037), .Z(n39040) );
  XNOR U38437 ( .A(n39035), .B(n39034), .Z(n39037) );
  XNOR U38438 ( .A(n39032), .B(n39031), .Z(n39034) );
  XNOR U38439 ( .A(n39029), .B(n39028), .Z(n39031) );
  XNOR U38440 ( .A(n39026), .B(n39025), .Z(n39028) );
  XNOR U38441 ( .A(n39023), .B(n39022), .Z(n39025) );
  XNOR U38442 ( .A(n39020), .B(n39019), .Z(n39022) );
  XNOR U38443 ( .A(n39017), .B(n39016), .Z(n39019) );
  XNOR U38444 ( .A(n39014), .B(n39013), .Z(n39016) );
  XNOR U38445 ( .A(n39011), .B(n39010), .Z(n39013) );
  XNOR U38446 ( .A(n39008), .B(n39007), .Z(n39010) );
  XNOR U38447 ( .A(n39005), .B(n39004), .Z(n39007) );
  XNOR U38448 ( .A(n39002), .B(n39001), .Z(n39004) );
  XNOR U38449 ( .A(n38999), .B(n38998), .Z(n39001) );
  XNOR U38450 ( .A(n38996), .B(n38995), .Z(n38998) );
  XNOR U38451 ( .A(n38993), .B(n38992), .Z(n38995) );
  XNOR U38452 ( .A(n38990), .B(n38989), .Z(n38992) );
  XNOR U38453 ( .A(n38987), .B(n38986), .Z(n38989) );
  XNOR U38454 ( .A(n38984), .B(n38983), .Z(n38986) );
  XNOR U38455 ( .A(n38981), .B(n38980), .Z(n38983) );
  XNOR U38456 ( .A(n38978), .B(n38977), .Z(n38980) );
  XNOR U38457 ( .A(n38975), .B(n38974), .Z(n38977) );
  XNOR U38458 ( .A(n38972), .B(n38971), .Z(n38974) );
  XNOR U38459 ( .A(n38969), .B(n38968), .Z(n38971) );
  XNOR U38460 ( .A(n38966), .B(n38965), .Z(n38968) );
  XNOR U38461 ( .A(n38963), .B(n38962), .Z(n38965) );
  XNOR U38462 ( .A(n38960), .B(n38959), .Z(n38962) );
  XNOR U38463 ( .A(n38957), .B(n38956), .Z(n38959) );
  XNOR U38464 ( .A(n38954), .B(n38953), .Z(n38956) );
  XNOR U38465 ( .A(n38951), .B(n38950), .Z(n38953) );
  XNOR U38466 ( .A(n38948), .B(n38947), .Z(n38950) );
  XNOR U38467 ( .A(n38945), .B(n38944), .Z(n38947) );
  XNOR U38468 ( .A(n38942), .B(n38941), .Z(n38944) );
  XNOR U38469 ( .A(n38939), .B(n38938), .Z(n38941) );
  XNOR U38470 ( .A(n38936), .B(n38935), .Z(n38938) );
  XNOR U38471 ( .A(n38933), .B(n38932), .Z(n38935) );
  XNOR U38472 ( .A(n38930), .B(n38929), .Z(n38932) );
  XNOR U38473 ( .A(n38927), .B(n38926), .Z(n38929) );
  XNOR U38474 ( .A(n38924), .B(n38923), .Z(n38926) );
  XNOR U38475 ( .A(n38921), .B(n38920), .Z(n38923) );
  XNOR U38476 ( .A(n38918), .B(n38917), .Z(n38920) );
  XNOR U38477 ( .A(n38915), .B(n38914), .Z(n38917) );
  XNOR U38478 ( .A(n38912), .B(n38911), .Z(n38914) );
  XNOR U38479 ( .A(n38909), .B(n38908), .Z(n38911) );
  XNOR U38480 ( .A(n38906), .B(n38905), .Z(n38908) );
  XNOR U38481 ( .A(n38903), .B(n38902), .Z(n38905) );
  XNOR U38482 ( .A(n38900), .B(n38899), .Z(n38902) );
  XNOR U38483 ( .A(n38897), .B(n38896), .Z(n38899) );
  XNOR U38484 ( .A(n38894), .B(n38893), .Z(n38896) );
  XNOR U38485 ( .A(n38891), .B(n38890), .Z(n38893) );
  XNOR U38486 ( .A(n38888), .B(n38887), .Z(n38890) );
  XNOR U38487 ( .A(n38885), .B(n38884), .Z(n38887) );
  XNOR U38488 ( .A(n38882), .B(n38881), .Z(n38884) );
  XNOR U38489 ( .A(n38879), .B(n38878), .Z(n38881) );
  XNOR U38490 ( .A(n38876), .B(n38875), .Z(n38878) );
  XNOR U38491 ( .A(n38873), .B(n38872), .Z(n38875) );
  XNOR U38492 ( .A(n38870), .B(n38869), .Z(n38872) );
  XNOR U38493 ( .A(n38867), .B(n38866), .Z(n38869) );
  XNOR U38494 ( .A(n38864), .B(n38863), .Z(n38866) );
  XNOR U38495 ( .A(n38861), .B(n38860), .Z(n38863) );
  XNOR U38496 ( .A(n38858), .B(n38857), .Z(n38860) );
  XNOR U38497 ( .A(n38855), .B(n38854), .Z(n38857) );
  XNOR U38498 ( .A(n38852), .B(n38851), .Z(n38854) );
  XNOR U38499 ( .A(n38849), .B(n38848), .Z(n38851) );
  XNOR U38500 ( .A(n38846), .B(n38845), .Z(n38848) );
  XNOR U38501 ( .A(n38843), .B(n38842), .Z(n38845) );
  XNOR U38502 ( .A(n38840), .B(n38839), .Z(n38842) );
  XNOR U38503 ( .A(n38837), .B(n38836), .Z(n38839) );
  XNOR U38504 ( .A(n38834), .B(n38833), .Z(n38836) );
  XNOR U38505 ( .A(n38831), .B(n38830), .Z(n38833) );
  XNOR U38506 ( .A(n38828), .B(n38827), .Z(n38830) );
  XNOR U38507 ( .A(n38825), .B(n38824), .Z(n38827) );
  XNOR U38508 ( .A(n38822), .B(n38821), .Z(n38824) );
  XNOR U38509 ( .A(n38819), .B(n38818), .Z(n38821) );
  XNOR U38510 ( .A(n38816), .B(n38815), .Z(n38818) );
  XNOR U38511 ( .A(n38813), .B(n38812), .Z(n38815) );
  XNOR U38512 ( .A(n38810), .B(n38809), .Z(n38812) );
  XNOR U38513 ( .A(n38807), .B(n38806), .Z(n38809) );
  XNOR U38514 ( .A(n38804), .B(n38803), .Z(n38806) );
  XNOR U38515 ( .A(n38801), .B(n38800), .Z(n38803) );
  XNOR U38516 ( .A(n38798), .B(n38797), .Z(n38800) );
  XNOR U38517 ( .A(n38795), .B(n38794), .Z(n38797) );
  XNOR U38518 ( .A(n38792), .B(n38791), .Z(n38794) );
  XNOR U38519 ( .A(n38789), .B(n38788), .Z(n38791) );
  XNOR U38520 ( .A(n38786), .B(n38785), .Z(n38788) );
  XNOR U38521 ( .A(n38783), .B(n38782), .Z(n38785) );
  XNOR U38522 ( .A(n38780), .B(n38779), .Z(n38782) );
  XNOR U38523 ( .A(n38777), .B(n38776), .Z(n38779) );
  XNOR U38524 ( .A(n38774), .B(n38773), .Z(n38776) );
  XNOR U38525 ( .A(n38771), .B(n38770), .Z(n38773) );
  XNOR U38526 ( .A(n38768), .B(n38767), .Z(n38770) );
  XNOR U38527 ( .A(n38765), .B(n38764), .Z(n38767) );
  XNOR U38528 ( .A(n38762), .B(n38761), .Z(n38764) );
  XNOR U38529 ( .A(n38759), .B(n38758), .Z(n38761) );
  XNOR U38530 ( .A(n38756), .B(n38755), .Z(n38758) );
  XNOR U38531 ( .A(n38753), .B(n38752), .Z(n38755) );
  XNOR U38532 ( .A(n38750), .B(n38749), .Z(n38752) );
  XNOR U38533 ( .A(n38747), .B(n38746), .Z(n38749) );
  XNOR U38534 ( .A(n38744), .B(n38743), .Z(n38746) );
  XNOR U38535 ( .A(n38741), .B(n38740), .Z(n38743) );
  XNOR U38536 ( .A(n38738), .B(n38737), .Z(n38740) );
  XNOR U38537 ( .A(n38735), .B(n38734), .Z(n38737) );
  XNOR U38538 ( .A(n38732), .B(n38731), .Z(n38734) );
  XNOR U38539 ( .A(n38729), .B(n38728), .Z(n38731) );
  XNOR U38540 ( .A(n38726), .B(n38725), .Z(n38728) );
  XNOR U38541 ( .A(n38723), .B(n38722), .Z(n38725) );
  XNOR U38542 ( .A(n38720), .B(n38719), .Z(n38722) );
  XNOR U38543 ( .A(n38717), .B(n38716), .Z(n38719) );
  XNOR U38544 ( .A(n38714), .B(n38713), .Z(n38716) );
  XNOR U38545 ( .A(n38711), .B(n38710), .Z(n38713) );
  XNOR U38546 ( .A(n38708), .B(n38707), .Z(n38710) );
  XNOR U38547 ( .A(n38705), .B(n38704), .Z(n38707) );
  XNOR U38548 ( .A(n38702), .B(n38701), .Z(n38704) );
  XNOR U38549 ( .A(n38699), .B(n38698), .Z(n38701) );
  XNOR U38550 ( .A(n38696), .B(n38695), .Z(n38698) );
  XNOR U38551 ( .A(n38693), .B(n38692), .Z(n38695) );
  XNOR U38552 ( .A(n38690), .B(n38689), .Z(n38692) );
  XNOR U38553 ( .A(n38687), .B(n38686), .Z(n38689) );
  XNOR U38554 ( .A(n38684), .B(n38683), .Z(n38686) );
  XNOR U38555 ( .A(n38681), .B(n38680), .Z(n38683) );
  XNOR U38556 ( .A(n38678), .B(n38677), .Z(n38680) );
  XNOR U38557 ( .A(n38675), .B(n38674), .Z(n38677) );
  XNOR U38558 ( .A(n38672), .B(n38671), .Z(n38674) );
  XNOR U38559 ( .A(n38669), .B(n38668), .Z(n38671) );
  XNOR U38560 ( .A(n38666), .B(n38665), .Z(n38668) );
  XNOR U38561 ( .A(n38663), .B(n38662), .Z(n38665) );
  XNOR U38562 ( .A(n38660), .B(n38659), .Z(n38662) );
  XNOR U38563 ( .A(n38657), .B(n38656), .Z(n38659) );
  XNOR U38564 ( .A(n38654), .B(n38653), .Z(n38656) );
  XOR U38565 ( .A(n38651), .B(n38650), .Z(n38653) );
  XOR U38566 ( .A(n38648), .B(n38647), .Z(n38650) );
  XOR U38567 ( .A(n38644), .B(n38645), .Z(n38647) );
  AND U38568 ( .A(n41230), .B(n41231), .Z(n38645) );
  XOR U38569 ( .A(n38641), .B(n38642), .Z(n38644) );
  AND U38570 ( .A(n41232), .B(n41233), .Z(n38642) );
  XOR U38571 ( .A(n38638), .B(n38639), .Z(n38641) );
  AND U38572 ( .A(n41234), .B(n41235), .Z(n38639) );
  XNOR U38573 ( .A(n38388), .B(n38636), .Z(n38638) );
  AND U38574 ( .A(n41236), .B(n41237), .Z(n38636) );
  XOR U38575 ( .A(n38390), .B(n38389), .Z(n38388) );
  AND U38576 ( .A(n41238), .B(n41239), .Z(n38389) );
  XOR U38577 ( .A(n38392), .B(n38391), .Z(n38390) );
  AND U38578 ( .A(n41240), .B(n41241), .Z(n38391) );
  XOR U38579 ( .A(n38394), .B(n38393), .Z(n38392) );
  AND U38580 ( .A(n41242), .B(n41243), .Z(n38393) );
  XOR U38581 ( .A(n38396), .B(n38395), .Z(n38394) );
  AND U38582 ( .A(n41244), .B(n41245), .Z(n38395) );
  XOR U38583 ( .A(n38398), .B(n38397), .Z(n38396) );
  AND U38584 ( .A(n41246), .B(n41247), .Z(n38397) );
  XOR U38585 ( .A(n38400), .B(n38399), .Z(n38398) );
  AND U38586 ( .A(n41248), .B(n41249), .Z(n38399) );
  XOR U38587 ( .A(n38402), .B(n38401), .Z(n38400) );
  AND U38588 ( .A(n41250), .B(n41251), .Z(n38401) );
  XOR U38589 ( .A(n38404), .B(n38403), .Z(n38402) );
  AND U38590 ( .A(n41252), .B(n41253), .Z(n38403) );
  XOR U38591 ( .A(n38406), .B(n38405), .Z(n38404) );
  AND U38592 ( .A(n41254), .B(n41255), .Z(n38405) );
  XOR U38593 ( .A(n38408), .B(n38407), .Z(n38406) );
  AND U38594 ( .A(n41256), .B(n41257), .Z(n38407) );
  XOR U38595 ( .A(n38410), .B(n38409), .Z(n38408) );
  AND U38596 ( .A(n41258), .B(n41259), .Z(n38409) );
  XOR U38597 ( .A(n38412), .B(n38411), .Z(n38410) );
  AND U38598 ( .A(n41260), .B(n41261), .Z(n38411) );
  XOR U38599 ( .A(n38414), .B(n38413), .Z(n38412) );
  AND U38600 ( .A(n41262), .B(n41263), .Z(n38413) );
  XOR U38601 ( .A(n38416), .B(n38415), .Z(n38414) );
  AND U38602 ( .A(n41264), .B(n41265), .Z(n38415) );
  XOR U38603 ( .A(n38418), .B(n38417), .Z(n38416) );
  AND U38604 ( .A(n41266), .B(n41267), .Z(n38417) );
  XOR U38605 ( .A(n38420), .B(n38419), .Z(n38418) );
  AND U38606 ( .A(n41268), .B(n41269), .Z(n38419) );
  XOR U38607 ( .A(n38422), .B(n38421), .Z(n38420) );
  AND U38608 ( .A(n41270), .B(n41271), .Z(n38421) );
  XOR U38609 ( .A(n38424), .B(n38423), .Z(n38422) );
  AND U38610 ( .A(n41272), .B(n41273), .Z(n38423) );
  XOR U38611 ( .A(n38426), .B(n38425), .Z(n38424) );
  AND U38612 ( .A(n41274), .B(n41275), .Z(n38425) );
  XOR U38613 ( .A(n38428), .B(n38427), .Z(n38426) );
  AND U38614 ( .A(n41276), .B(n41277), .Z(n38427) );
  XOR U38615 ( .A(n38430), .B(n38429), .Z(n38428) );
  AND U38616 ( .A(n41278), .B(n41279), .Z(n38429) );
  XOR U38617 ( .A(n38432), .B(n38431), .Z(n38430) );
  AND U38618 ( .A(n41280), .B(n41281), .Z(n38431) );
  XOR U38619 ( .A(n38434), .B(n38433), .Z(n38432) );
  AND U38620 ( .A(n41282), .B(n41283), .Z(n38433) );
  XOR U38621 ( .A(n38436), .B(n38435), .Z(n38434) );
  AND U38622 ( .A(n41284), .B(n41285), .Z(n38435) );
  XOR U38623 ( .A(n38438), .B(n38437), .Z(n38436) );
  AND U38624 ( .A(n41286), .B(n41287), .Z(n38437) );
  XOR U38625 ( .A(n38440), .B(n38439), .Z(n38438) );
  AND U38626 ( .A(n41288), .B(n41289), .Z(n38439) );
  XOR U38627 ( .A(n38442), .B(n38441), .Z(n38440) );
  AND U38628 ( .A(n41290), .B(n41291), .Z(n38441) );
  XOR U38629 ( .A(n38444), .B(n38443), .Z(n38442) );
  AND U38630 ( .A(n41292), .B(n41293), .Z(n38443) );
  XOR U38631 ( .A(n38446), .B(n38445), .Z(n38444) );
  AND U38632 ( .A(n41294), .B(n41295), .Z(n38445) );
  XOR U38633 ( .A(n38448), .B(n38447), .Z(n38446) );
  AND U38634 ( .A(n41296), .B(n41297), .Z(n38447) );
  XOR U38635 ( .A(n38450), .B(n38449), .Z(n38448) );
  AND U38636 ( .A(n41298), .B(n41299), .Z(n38449) );
  XOR U38637 ( .A(n38452), .B(n38451), .Z(n38450) );
  AND U38638 ( .A(n41300), .B(n41301), .Z(n38451) );
  XOR U38639 ( .A(n38454), .B(n38453), .Z(n38452) );
  AND U38640 ( .A(n41302), .B(n41303), .Z(n38453) );
  XOR U38641 ( .A(n38456), .B(n38455), .Z(n38454) );
  AND U38642 ( .A(n41304), .B(n41305), .Z(n38455) );
  XOR U38643 ( .A(n38458), .B(n38457), .Z(n38456) );
  AND U38644 ( .A(n41306), .B(n41307), .Z(n38457) );
  XOR U38645 ( .A(n38460), .B(n38459), .Z(n38458) );
  AND U38646 ( .A(n41308), .B(n41309), .Z(n38459) );
  XOR U38647 ( .A(n38462), .B(n38461), .Z(n38460) );
  AND U38648 ( .A(n41310), .B(n41311), .Z(n38461) );
  XOR U38649 ( .A(n38464), .B(n38463), .Z(n38462) );
  AND U38650 ( .A(n41312), .B(n41313), .Z(n38463) );
  XOR U38651 ( .A(n38466), .B(n38465), .Z(n38464) );
  AND U38652 ( .A(n41314), .B(n41315), .Z(n38465) );
  XOR U38653 ( .A(n38468), .B(n38467), .Z(n38466) );
  AND U38654 ( .A(n41316), .B(n41317), .Z(n38467) );
  XOR U38655 ( .A(n38470), .B(n38469), .Z(n38468) );
  AND U38656 ( .A(n41318), .B(n41319), .Z(n38469) );
  XOR U38657 ( .A(n38472), .B(n38471), .Z(n38470) );
  AND U38658 ( .A(n41320), .B(n41321), .Z(n38471) );
  XOR U38659 ( .A(n38474), .B(n38473), .Z(n38472) );
  AND U38660 ( .A(n41322), .B(n41323), .Z(n38473) );
  XOR U38661 ( .A(n38476), .B(n38475), .Z(n38474) );
  AND U38662 ( .A(n41324), .B(n41325), .Z(n38475) );
  XOR U38663 ( .A(n38478), .B(n38477), .Z(n38476) );
  AND U38664 ( .A(n41326), .B(n41327), .Z(n38477) );
  XOR U38665 ( .A(n38480), .B(n38479), .Z(n38478) );
  AND U38666 ( .A(n41328), .B(n41329), .Z(n38479) );
  XOR U38667 ( .A(n38482), .B(n38481), .Z(n38480) );
  AND U38668 ( .A(n41330), .B(n41331), .Z(n38481) );
  XOR U38669 ( .A(n38484), .B(n38483), .Z(n38482) );
  AND U38670 ( .A(n41332), .B(n41333), .Z(n38483) );
  XOR U38671 ( .A(n38486), .B(n38485), .Z(n38484) );
  AND U38672 ( .A(n41334), .B(n41335), .Z(n38485) );
  XOR U38673 ( .A(n38488), .B(n38487), .Z(n38486) );
  AND U38674 ( .A(n41336), .B(n41337), .Z(n38487) );
  XOR U38675 ( .A(n38490), .B(n38489), .Z(n38488) );
  AND U38676 ( .A(n41338), .B(n41339), .Z(n38489) );
  XOR U38677 ( .A(n38492), .B(n38491), .Z(n38490) );
  AND U38678 ( .A(n41340), .B(n41341), .Z(n38491) );
  XOR U38679 ( .A(n38494), .B(n38493), .Z(n38492) );
  AND U38680 ( .A(n41342), .B(n41343), .Z(n38493) );
  XOR U38681 ( .A(n38496), .B(n38495), .Z(n38494) );
  AND U38682 ( .A(n41344), .B(n41345), .Z(n38495) );
  XOR U38683 ( .A(n38498), .B(n38497), .Z(n38496) );
  AND U38684 ( .A(n41346), .B(n41347), .Z(n38497) );
  XOR U38685 ( .A(n38500), .B(n38499), .Z(n38498) );
  AND U38686 ( .A(n41348), .B(n41349), .Z(n38499) );
  XOR U38687 ( .A(n38502), .B(n38501), .Z(n38500) );
  AND U38688 ( .A(n41350), .B(n41351), .Z(n38501) );
  XOR U38689 ( .A(n38504), .B(n38503), .Z(n38502) );
  AND U38690 ( .A(n41352), .B(n41353), .Z(n38503) );
  XOR U38691 ( .A(n38506), .B(n38505), .Z(n38504) );
  AND U38692 ( .A(n41354), .B(n41355), .Z(n38505) );
  XOR U38693 ( .A(n38508), .B(n38507), .Z(n38506) );
  AND U38694 ( .A(n41356), .B(n41357), .Z(n38507) );
  XOR U38695 ( .A(n38510), .B(n38509), .Z(n38508) );
  AND U38696 ( .A(n41358), .B(n41359), .Z(n38509) );
  XOR U38697 ( .A(n38512), .B(n38511), .Z(n38510) );
  AND U38698 ( .A(n41360), .B(n41361), .Z(n38511) );
  XOR U38699 ( .A(n38514), .B(n38513), .Z(n38512) );
  AND U38700 ( .A(n41362), .B(n41363), .Z(n38513) );
  XOR U38701 ( .A(n38516), .B(n38515), .Z(n38514) );
  AND U38702 ( .A(n41364), .B(n41365), .Z(n38515) );
  XOR U38703 ( .A(n38518), .B(n38517), .Z(n38516) );
  AND U38704 ( .A(n41366), .B(n41367), .Z(n38517) );
  XOR U38705 ( .A(n38520), .B(n38519), .Z(n38518) );
  AND U38706 ( .A(n41368), .B(n41369), .Z(n38519) );
  XOR U38707 ( .A(n38522), .B(n38521), .Z(n38520) );
  AND U38708 ( .A(n41370), .B(n41371), .Z(n38521) );
  XOR U38709 ( .A(n38524), .B(n38523), .Z(n38522) );
  AND U38710 ( .A(n41372), .B(n41373), .Z(n38523) );
  XOR U38711 ( .A(n38526), .B(n38525), .Z(n38524) );
  AND U38712 ( .A(n41374), .B(n41375), .Z(n38525) );
  XOR U38713 ( .A(n38528), .B(n38527), .Z(n38526) );
  AND U38714 ( .A(n41376), .B(n41377), .Z(n38527) );
  XOR U38715 ( .A(n38530), .B(n38529), .Z(n38528) );
  AND U38716 ( .A(n41378), .B(n41379), .Z(n38529) );
  XOR U38717 ( .A(n38532), .B(n38531), .Z(n38530) );
  AND U38718 ( .A(n41380), .B(n41381), .Z(n38531) );
  XOR U38719 ( .A(n38534), .B(n38533), .Z(n38532) );
  AND U38720 ( .A(n41382), .B(n41383), .Z(n38533) );
  XOR U38721 ( .A(n38536), .B(n38535), .Z(n38534) );
  AND U38722 ( .A(n41384), .B(n41385), .Z(n38535) );
  XOR U38723 ( .A(n38538), .B(n38537), .Z(n38536) );
  AND U38724 ( .A(n41386), .B(n41387), .Z(n38537) );
  XOR U38725 ( .A(n38540), .B(n38539), .Z(n38538) );
  AND U38726 ( .A(n41388), .B(n41389), .Z(n38539) );
  XOR U38727 ( .A(n38542), .B(n38541), .Z(n38540) );
  AND U38728 ( .A(n41390), .B(n41391), .Z(n38541) );
  XOR U38729 ( .A(n38544), .B(n38543), .Z(n38542) );
  AND U38730 ( .A(n41392), .B(n41393), .Z(n38543) );
  XOR U38731 ( .A(n38546), .B(n38545), .Z(n38544) );
  AND U38732 ( .A(n41394), .B(n41395), .Z(n38545) );
  XOR U38733 ( .A(n38548), .B(n38547), .Z(n38546) );
  AND U38734 ( .A(n41396), .B(n41397), .Z(n38547) );
  XOR U38735 ( .A(n38550), .B(n38549), .Z(n38548) );
  AND U38736 ( .A(n41398), .B(n41399), .Z(n38549) );
  XOR U38737 ( .A(n38552), .B(n38551), .Z(n38550) );
  AND U38738 ( .A(n41400), .B(n41401), .Z(n38551) );
  XOR U38739 ( .A(n38554), .B(n38553), .Z(n38552) );
  AND U38740 ( .A(n41402), .B(n41403), .Z(n38553) );
  XOR U38741 ( .A(n38556), .B(n38555), .Z(n38554) );
  AND U38742 ( .A(n41404), .B(n41405), .Z(n38555) );
  XOR U38743 ( .A(n38558), .B(n38557), .Z(n38556) );
  AND U38744 ( .A(n41406), .B(n41407), .Z(n38557) );
  XOR U38745 ( .A(n38560), .B(n38559), .Z(n38558) );
  AND U38746 ( .A(n41408), .B(n41409), .Z(n38559) );
  XOR U38747 ( .A(n38562), .B(n38561), .Z(n38560) );
  AND U38748 ( .A(n41410), .B(n41411), .Z(n38561) );
  XOR U38749 ( .A(n38564), .B(n38563), .Z(n38562) );
  AND U38750 ( .A(n41412), .B(n41413), .Z(n38563) );
  XOR U38751 ( .A(n38566), .B(n38565), .Z(n38564) );
  AND U38752 ( .A(n41414), .B(n41415), .Z(n38565) );
  XOR U38753 ( .A(n38568), .B(n38567), .Z(n38566) );
  AND U38754 ( .A(n41416), .B(n41417), .Z(n38567) );
  XOR U38755 ( .A(n38570), .B(n38569), .Z(n38568) );
  AND U38756 ( .A(n41418), .B(n41419), .Z(n38569) );
  XOR U38757 ( .A(n38572), .B(n38571), .Z(n38570) );
  AND U38758 ( .A(n41420), .B(n41421), .Z(n38571) );
  XOR U38759 ( .A(n38574), .B(n38573), .Z(n38572) );
  AND U38760 ( .A(n41422), .B(n41423), .Z(n38573) );
  XOR U38761 ( .A(n38576), .B(n38575), .Z(n38574) );
  AND U38762 ( .A(n41424), .B(n41425), .Z(n38575) );
  XOR U38763 ( .A(n38578), .B(n38577), .Z(n38576) );
  AND U38764 ( .A(n41426), .B(n41427), .Z(n38577) );
  XOR U38765 ( .A(n38580), .B(n38579), .Z(n38578) );
  AND U38766 ( .A(n41428), .B(n41429), .Z(n38579) );
  XOR U38767 ( .A(n38632), .B(n38581), .Z(n38580) );
  AND U38768 ( .A(n41430), .B(n41431), .Z(n38581) );
  XOR U38769 ( .A(n38634), .B(n38633), .Z(n38632) );
  AND U38770 ( .A(n41432), .B(n41433), .Z(n38633) );
  XOR U38771 ( .A(n38616), .B(n38635), .Z(n38634) );
  AND U38772 ( .A(n41434), .B(n41435), .Z(n38635) );
  XOR U38773 ( .A(n38618), .B(n38617), .Z(n38616) );
  AND U38774 ( .A(n41436), .B(n41437), .Z(n38617) );
  XOR U38775 ( .A(n38620), .B(n38619), .Z(n38618) );
  AND U38776 ( .A(n41438), .B(n41439), .Z(n38619) );
  XOR U38777 ( .A(n38624), .B(n38621), .Z(n38620) );
  AND U38778 ( .A(n41440), .B(n41441), .Z(n38621) );
  XOR U38779 ( .A(n38626), .B(n38625), .Z(n38624) );
  AND U38780 ( .A(n41442), .B(n41443), .Z(n38625) );
  XOR U38781 ( .A(n38628), .B(n38627), .Z(n38626) );
  AND U38782 ( .A(n41444), .B(n41445), .Z(n38627) );
  XOR U38783 ( .A(n38630), .B(n38629), .Z(n38628) );
  AND U38784 ( .A(n41446), .B(n41447), .Z(n38629) );
  XOR U38785 ( .A(n38605), .B(n38631), .Z(n38630) );
  AND U38786 ( .A(n41448), .B(n41449), .Z(n38631) );
  XNOR U38787 ( .A(n38602), .B(n38606), .Z(n38605) );
  AND U38788 ( .A(n41450), .B(n41451), .Z(n38606) );
  XOR U38789 ( .A(n38601), .B(n38593), .Z(n38602) );
  AND U38790 ( .A(n41452), .B(n41453), .Z(n38593) );
  XNOR U38791 ( .A(n38596), .B(n38592), .Z(n38601) );
  AND U38792 ( .A(n41454), .B(n41455), .Z(n38592) );
  XOR U38793 ( .A(n41456), .B(n41457), .Z(n38596) );
  XOR U38794 ( .A(n38614), .B(n41458), .Z(n41457) );
  XOR U38795 ( .A(n38612), .B(n38610), .Z(n41458) );
  AND U38796 ( .A(n41459), .B(n41460), .Z(n38610) );
  AND U38797 ( .A(n41461), .B(n41462), .Z(n38612) );
  AND U38798 ( .A(n41463), .B(n41464), .Z(n38614) );
  XNOR U38799 ( .A(n41465), .B(n38613), .Z(n41456) );
  XOR U38800 ( .A(n41466), .B(n41467), .Z(n38613) );
  XOR U38801 ( .A(n41468), .B(n41469), .Z(n41467) );
  AND U38802 ( .A(n41470), .B(n41471), .Z(n41469) );
  XNOR U38803 ( .A(n41472), .B(n41473), .Z(n41466) );
  NOR U38804 ( .A(n41474), .B(n41475), .Z(n41473) );
  AND U38805 ( .A(n41476), .B(n41477), .Z(n41475) );
  IV U38806 ( .A(n41478), .Z(n41474) );
  NOR U38807 ( .A(n41468), .B(n41479), .Z(n41478) );
  AND U38808 ( .A(n41480), .B(n41481), .Z(n41479) );
  NOR U38809 ( .A(n41470), .B(n41480), .Z(n41472) );
  XNOR U38810 ( .A(n38615), .B(n38597), .Z(n41465) );
  AND U38811 ( .A(n41482), .B(n41483), .Z(n38597) );
  AND U38812 ( .A(n41484), .B(n41485), .Z(n38615) );
  XOR U38813 ( .A(n41486), .B(n41487), .Z(n38648) );
  NOR U38814 ( .A(n41488), .B(n41489), .Z(n41487) );
  IV U38815 ( .A(n41486), .Z(n41488) );
  XOR U38816 ( .A(n41490), .B(n41491), .Z(n38651) );
  NOR U38817 ( .A(n41490), .B(n41492), .Z(n41491) );
  XNOR U38818 ( .A(n41493), .B(n41494), .Z(n38654) );
  AND U38819 ( .A(n41493), .B(n41495), .Z(n41494) );
  XNOR U38820 ( .A(n41496), .B(n41497), .Z(n38657) );
  AND U38821 ( .A(n41496), .B(n41498), .Z(n41497) );
  XNOR U38822 ( .A(n41499), .B(n41500), .Z(n38660) );
  AND U38823 ( .A(n41499), .B(n41501), .Z(n41500) );
  XNOR U38824 ( .A(n41502), .B(n41503), .Z(n38663) );
  AND U38825 ( .A(n41502), .B(n41504), .Z(n41503) );
  XNOR U38826 ( .A(n41505), .B(n41506), .Z(n38666) );
  AND U38827 ( .A(n41505), .B(n41507), .Z(n41506) );
  XNOR U38828 ( .A(n41508), .B(n41509), .Z(n38669) );
  AND U38829 ( .A(n41508), .B(n41510), .Z(n41509) );
  XNOR U38830 ( .A(n41511), .B(n41512), .Z(n38672) );
  AND U38831 ( .A(n41511), .B(n41513), .Z(n41512) );
  XNOR U38832 ( .A(n41514), .B(n41515), .Z(n38675) );
  AND U38833 ( .A(n41514), .B(n41516), .Z(n41515) );
  XNOR U38834 ( .A(n41517), .B(n41518), .Z(n38678) );
  AND U38835 ( .A(n41517), .B(n41519), .Z(n41518) );
  XNOR U38836 ( .A(n41520), .B(n41521), .Z(n38681) );
  AND U38837 ( .A(n41520), .B(n41522), .Z(n41521) );
  XNOR U38838 ( .A(n41523), .B(n41524), .Z(n38684) );
  AND U38839 ( .A(n41523), .B(n41525), .Z(n41524) );
  XNOR U38840 ( .A(n41526), .B(n41527), .Z(n38687) );
  AND U38841 ( .A(n41526), .B(n41528), .Z(n41527) );
  XNOR U38842 ( .A(n41529), .B(n41530), .Z(n38690) );
  AND U38843 ( .A(n41529), .B(n41531), .Z(n41530) );
  XNOR U38844 ( .A(n41532), .B(n41533), .Z(n38693) );
  AND U38845 ( .A(n41532), .B(n41534), .Z(n41533) );
  XNOR U38846 ( .A(n41535), .B(n41536), .Z(n38696) );
  AND U38847 ( .A(n41535), .B(n41537), .Z(n41536) );
  XNOR U38848 ( .A(n41538), .B(n41539), .Z(n38699) );
  AND U38849 ( .A(n41538), .B(n41540), .Z(n41539) );
  XNOR U38850 ( .A(n41541), .B(n41542), .Z(n38702) );
  AND U38851 ( .A(n41541), .B(n41543), .Z(n41542) );
  XNOR U38852 ( .A(n41544), .B(n41545), .Z(n38705) );
  AND U38853 ( .A(n41544), .B(n41546), .Z(n41545) );
  XNOR U38854 ( .A(n41547), .B(n41548), .Z(n38708) );
  AND U38855 ( .A(n41547), .B(n41549), .Z(n41548) );
  XNOR U38856 ( .A(n41550), .B(n41551), .Z(n38711) );
  AND U38857 ( .A(n41550), .B(n41552), .Z(n41551) );
  XNOR U38858 ( .A(n41553), .B(n41554), .Z(n38714) );
  AND U38859 ( .A(n41553), .B(n41555), .Z(n41554) );
  XNOR U38860 ( .A(n41556), .B(n41557), .Z(n38717) );
  AND U38861 ( .A(n41556), .B(n41558), .Z(n41557) );
  XNOR U38862 ( .A(n41559), .B(n41560), .Z(n38720) );
  AND U38863 ( .A(n41559), .B(n41561), .Z(n41560) );
  XNOR U38864 ( .A(n41562), .B(n41563), .Z(n38723) );
  AND U38865 ( .A(n41562), .B(n41564), .Z(n41563) );
  XNOR U38866 ( .A(n41565), .B(n41566), .Z(n38726) );
  AND U38867 ( .A(n41565), .B(n41567), .Z(n41566) );
  XNOR U38868 ( .A(n41568), .B(n41569), .Z(n38729) );
  AND U38869 ( .A(n41568), .B(n41570), .Z(n41569) );
  XNOR U38870 ( .A(n41571), .B(n41572), .Z(n38732) );
  AND U38871 ( .A(n41571), .B(n41573), .Z(n41572) );
  XNOR U38872 ( .A(n41574), .B(n41575), .Z(n38735) );
  AND U38873 ( .A(n41574), .B(n41576), .Z(n41575) );
  XNOR U38874 ( .A(n41577), .B(n41578), .Z(n38738) );
  AND U38875 ( .A(n41577), .B(n41579), .Z(n41578) );
  XNOR U38876 ( .A(n41580), .B(n41581), .Z(n38741) );
  AND U38877 ( .A(n41580), .B(n41582), .Z(n41581) );
  XNOR U38878 ( .A(n41583), .B(n41584), .Z(n38744) );
  AND U38879 ( .A(n41583), .B(n41585), .Z(n41584) );
  XNOR U38880 ( .A(n41586), .B(n41587), .Z(n38747) );
  AND U38881 ( .A(n41586), .B(n41588), .Z(n41587) );
  XNOR U38882 ( .A(n41589), .B(n41590), .Z(n38750) );
  AND U38883 ( .A(n41589), .B(n41591), .Z(n41590) );
  XNOR U38884 ( .A(n41592), .B(n41593), .Z(n38753) );
  AND U38885 ( .A(n41592), .B(n41594), .Z(n41593) );
  XNOR U38886 ( .A(n41595), .B(n41596), .Z(n38756) );
  AND U38887 ( .A(n41595), .B(n41597), .Z(n41596) );
  XNOR U38888 ( .A(n41598), .B(n41599), .Z(n38759) );
  AND U38889 ( .A(n41598), .B(n41600), .Z(n41599) );
  XNOR U38890 ( .A(n41601), .B(n41602), .Z(n38762) );
  AND U38891 ( .A(n41601), .B(n41603), .Z(n41602) );
  XNOR U38892 ( .A(n41604), .B(n41605), .Z(n38765) );
  AND U38893 ( .A(n41604), .B(n41606), .Z(n41605) );
  XNOR U38894 ( .A(n41607), .B(n41608), .Z(n38768) );
  AND U38895 ( .A(n41607), .B(n41609), .Z(n41608) );
  XNOR U38896 ( .A(n41610), .B(n41611), .Z(n38771) );
  AND U38897 ( .A(n41610), .B(n41612), .Z(n41611) );
  XNOR U38898 ( .A(n41613), .B(n41614), .Z(n38774) );
  AND U38899 ( .A(n41613), .B(n41615), .Z(n41614) );
  XNOR U38900 ( .A(n41616), .B(n41617), .Z(n38777) );
  AND U38901 ( .A(n41616), .B(n41618), .Z(n41617) );
  XNOR U38902 ( .A(n41619), .B(n41620), .Z(n38780) );
  AND U38903 ( .A(n41619), .B(n41621), .Z(n41620) );
  XNOR U38904 ( .A(n41622), .B(n41623), .Z(n38783) );
  AND U38905 ( .A(n41622), .B(n41624), .Z(n41623) );
  XNOR U38906 ( .A(n41625), .B(n41626), .Z(n38786) );
  AND U38907 ( .A(n41625), .B(n41627), .Z(n41626) );
  XNOR U38908 ( .A(n41628), .B(n41629), .Z(n38789) );
  AND U38909 ( .A(n41628), .B(n41630), .Z(n41629) );
  XNOR U38910 ( .A(n41631), .B(n41632), .Z(n38792) );
  AND U38911 ( .A(n41631), .B(n41633), .Z(n41632) );
  XNOR U38912 ( .A(n41634), .B(n41635), .Z(n38795) );
  AND U38913 ( .A(n41634), .B(n41636), .Z(n41635) );
  XNOR U38914 ( .A(n41637), .B(n41638), .Z(n38798) );
  AND U38915 ( .A(n41637), .B(n41639), .Z(n41638) );
  XNOR U38916 ( .A(n41640), .B(n41641), .Z(n38801) );
  AND U38917 ( .A(n41640), .B(n41642), .Z(n41641) );
  XNOR U38918 ( .A(n41643), .B(n41644), .Z(n38804) );
  AND U38919 ( .A(n41643), .B(n41645), .Z(n41644) );
  XNOR U38920 ( .A(n41646), .B(n41647), .Z(n38807) );
  AND U38921 ( .A(n41646), .B(n41648), .Z(n41647) );
  XNOR U38922 ( .A(n41649), .B(n41650), .Z(n38810) );
  AND U38923 ( .A(n41649), .B(n41651), .Z(n41650) );
  XNOR U38924 ( .A(n41652), .B(n41653), .Z(n38813) );
  AND U38925 ( .A(n41652), .B(n41654), .Z(n41653) );
  XNOR U38926 ( .A(n41655), .B(n41656), .Z(n38816) );
  AND U38927 ( .A(n41655), .B(n41657), .Z(n41656) );
  XNOR U38928 ( .A(n41658), .B(n41659), .Z(n38819) );
  AND U38929 ( .A(n41658), .B(n41660), .Z(n41659) );
  XNOR U38930 ( .A(n41661), .B(n41662), .Z(n38822) );
  AND U38931 ( .A(n41661), .B(n41663), .Z(n41662) );
  XNOR U38932 ( .A(n41664), .B(n41665), .Z(n38825) );
  AND U38933 ( .A(n41664), .B(n41666), .Z(n41665) );
  XNOR U38934 ( .A(n41667), .B(n41668), .Z(n38828) );
  AND U38935 ( .A(n41667), .B(n41669), .Z(n41668) );
  XNOR U38936 ( .A(n41670), .B(n41671), .Z(n38831) );
  AND U38937 ( .A(n41670), .B(n41672), .Z(n41671) );
  XNOR U38938 ( .A(n41673), .B(n41674), .Z(n38834) );
  AND U38939 ( .A(n41673), .B(n41675), .Z(n41674) );
  XNOR U38940 ( .A(n41676), .B(n41677), .Z(n38837) );
  AND U38941 ( .A(n41676), .B(n41678), .Z(n41677) );
  XNOR U38942 ( .A(n41679), .B(n41680), .Z(n38840) );
  AND U38943 ( .A(n41679), .B(n41681), .Z(n41680) );
  XNOR U38944 ( .A(n41682), .B(n41683), .Z(n38843) );
  AND U38945 ( .A(n41682), .B(n41684), .Z(n41683) );
  XNOR U38946 ( .A(n41685), .B(n41686), .Z(n38846) );
  AND U38947 ( .A(n41685), .B(n41687), .Z(n41686) );
  XNOR U38948 ( .A(n41688), .B(n41689), .Z(n38849) );
  AND U38949 ( .A(n41688), .B(n41690), .Z(n41689) );
  XNOR U38950 ( .A(n41691), .B(n41692), .Z(n38852) );
  AND U38951 ( .A(n41691), .B(n41693), .Z(n41692) );
  XNOR U38952 ( .A(n41694), .B(n41695), .Z(n38855) );
  AND U38953 ( .A(n41694), .B(n41696), .Z(n41695) );
  XNOR U38954 ( .A(n41697), .B(n41698), .Z(n38858) );
  AND U38955 ( .A(n41697), .B(n41699), .Z(n41698) );
  XNOR U38956 ( .A(n41700), .B(n41701), .Z(n38861) );
  AND U38957 ( .A(n41700), .B(n41702), .Z(n41701) );
  XNOR U38958 ( .A(n41703), .B(n41704), .Z(n38864) );
  AND U38959 ( .A(n41703), .B(n41705), .Z(n41704) );
  XNOR U38960 ( .A(n41706), .B(n41707), .Z(n38867) );
  AND U38961 ( .A(n41706), .B(n41708), .Z(n41707) );
  XNOR U38962 ( .A(n41709), .B(n41710), .Z(n38870) );
  AND U38963 ( .A(n41709), .B(n41711), .Z(n41710) );
  XNOR U38964 ( .A(n41712), .B(n41713), .Z(n38873) );
  AND U38965 ( .A(n41712), .B(n41714), .Z(n41713) );
  XNOR U38966 ( .A(n41715), .B(n41716), .Z(n38876) );
  AND U38967 ( .A(n41715), .B(n41717), .Z(n41716) );
  XNOR U38968 ( .A(n41718), .B(n41719), .Z(n38879) );
  AND U38969 ( .A(n41718), .B(n41720), .Z(n41719) );
  XNOR U38970 ( .A(n41721), .B(n41722), .Z(n38882) );
  AND U38971 ( .A(n41721), .B(n41723), .Z(n41722) );
  XNOR U38972 ( .A(n41724), .B(n41725), .Z(n38885) );
  AND U38973 ( .A(n41724), .B(n41726), .Z(n41725) );
  XNOR U38974 ( .A(n41727), .B(n41728), .Z(n38888) );
  AND U38975 ( .A(n41727), .B(n41729), .Z(n41728) );
  XNOR U38976 ( .A(n41730), .B(n41731), .Z(n38891) );
  AND U38977 ( .A(n41730), .B(n41732), .Z(n41731) );
  XNOR U38978 ( .A(n41733), .B(n41734), .Z(n38894) );
  AND U38979 ( .A(n41733), .B(n41735), .Z(n41734) );
  XNOR U38980 ( .A(n41736), .B(n41737), .Z(n38897) );
  AND U38981 ( .A(n41736), .B(n41738), .Z(n41737) );
  XNOR U38982 ( .A(n41739), .B(n41740), .Z(n38900) );
  AND U38983 ( .A(n41739), .B(n41741), .Z(n41740) );
  XNOR U38984 ( .A(n41742), .B(n41743), .Z(n38903) );
  AND U38985 ( .A(n41742), .B(n41744), .Z(n41743) );
  XNOR U38986 ( .A(n41745), .B(n41746), .Z(n38906) );
  AND U38987 ( .A(n41745), .B(n41747), .Z(n41746) );
  XNOR U38988 ( .A(n41748), .B(n41749), .Z(n38909) );
  AND U38989 ( .A(n41748), .B(n41750), .Z(n41749) );
  XNOR U38990 ( .A(n41751), .B(n41752), .Z(n38912) );
  AND U38991 ( .A(n41751), .B(n41753), .Z(n41752) );
  XNOR U38992 ( .A(n41754), .B(n41755), .Z(n38915) );
  AND U38993 ( .A(n41754), .B(n41756), .Z(n41755) );
  XNOR U38994 ( .A(n41757), .B(n41758), .Z(n38918) );
  AND U38995 ( .A(n41757), .B(n41759), .Z(n41758) );
  XNOR U38996 ( .A(n41760), .B(n41761), .Z(n38921) );
  AND U38997 ( .A(n41760), .B(n41762), .Z(n41761) );
  XNOR U38998 ( .A(n41763), .B(n41764), .Z(n38924) );
  AND U38999 ( .A(n41763), .B(n41765), .Z(n41764) );
  XNOR U39000 ( .A(n41766), .B(n41767), .Z(n38927) );
  AND U39001 ( .A(n41766), .B(n41768), .Z(n41767) );
  XNOR U39002 ( .A(n41769), .B(n41770), .Z(n38930) );
  AND U39003 ( .A(n41769), .B(n41771), .Z(n41770) );
  XNOR U39004 ( .A(n41772), .B(n41773), .Z(n38933) );
  AND U39005 ( .A(n41772), .B(n41774), .Z(n41773) );
  XNOR U39006 ( .A(n41775), .B(n41776), .Z(n38936) );
  AND U39007 ( .A(n41775), .B(n41777), .Z(n41776) );
  XNOR U39008 ( .A(n41778), .B(n41779), .Z(n38939) );
  AND U39009 ( .A(n41778), .B(n41780), .Z(n41779) );
  XNOR U39010 ( .A(n41781), .B(n41782), .Z(n38942) );
  AND U39011 ( .A(n41781), .B(n41783), .Z(n41782) );
  XNOR U39012 ( .A(n41784), .B(n41785), .Z(n38945) );
  AND U39013 ( .A(n41784), .B(n41786), .Z(n41785) );
  XNOR U39014 ( .A(n41787), .B(n41788), .Z(n38948) );
  AND U39015 ( .A(n41787), .B(n41789), .Z(n41788) );
  XNOR U39016 ( .A(n41790), .B(n41791), .Z(n38951) );
  AND U39017 ( .A(n41790), .B(n41792), .Z(n41791) );
  XNOR U39018 ( .A(n41793), .B(n41794), .Z(n38954) );
  AND U39019 ( .A(n41793), .B(n41795), .Z(n41794) );
  XNOR U39020 ( .A(n41796), .B(n41797), .Z(n38957) );
  AND U39021 ( .A(n41796), .B(n41798), .Z(n41797) );
  XNOR U39022 ( .A(n41799), .B(n41800), .Z(n38960) );
  AND U39023 ( .A(n41799), .B(n41801), .Z(n41800) );
  XNOR U39024 ( .A(n41802), .B(n41803), .Z(n38963) );
  AND U39025 ( .A(n41802), .B(n41804), .Z(n41803) );
  XNOR U39026 ( .A(n41805), .B(n41806), .Z(n38966) );
  AND U39027 ( .A(n41805), .B(n41807), .Z(n41806) );
  XNOR U39028 ( .A(n41808), .B(n41809), .Z(n38969) );
  AND U39029 ( .A(n41808), .B(n41810), .Z(n41809) );
  XNOR U39030 ( .A(n41811), .B(n41812), .Z(n38972) );
  AND U39031 ( .A(n41811), .B(n41813), .Z(n41812) );
  XNOR U39032 ( .A(n41814), .B(n41815), .Z(n38975) );
  AND U39033 ( .A(n41814), .B(n41816), .Z(n41815) );
  XNOR U39034 ( .A(n41817), .B(n41818), .Z(n38978) );
  AND U39035 ( .A(n41817), .B(n41819), .Z(n41818) );
  XNOR U39036 ( .A(n41820), .B(n41821), .Z(n38981) );
  AND U39037 ( .A(n41820), .B(n41822), .Z(n41821) );
  XNOR U39038 ( .A(n41823), .B(n41824), .Z(n38984) );
  AND U39039 ( .A(n41823), .B(n41825), .Z(n41824) );
  XNOR U39040 ( .A(n41826), .B(n41827), .Z(n38987) );
  AND U39041 ( .A(n41826), .B(n41828), .Z(n41827) );
  XNOR U39042 ( .A(n41829), .B(n41830), .Z(n38990) );
  AND U39043 ( .A(n41829), .B(n41831), .Z(n41830) );
  XNOR U39044 ( .A(n41832), .B(n41833), .Z(n38993) );
  AND U39045 ( .A(n41832), .B(n41834), .Z(n41833) );
  XNOR U39046 ( .A(n41835), .B(n41836), .Z(n38996) );
  AND U39047 ( .A(n41835), .B(n41837), .Z(n41836) );
  XNOR U39048 ( .A(n41838), .B(n41839), .Z(n38999) );
  AND U39049 ( .A(n41838), .B(n41840), .Z(n41839) );
  XNOR U39050 ( .A(n41841), .B(n41842), .Z(n39002) );
  AND U39051 ( .A(n41841), .B(n41843), .Z(n41842) );
  XNOR U39052 ( .A(n41844), .B(n41845), .Z(n39005) );
  AND U39053 ( .A(n41844), .B(n41846), .Z(n41845) );
  XNOR U39054 ( .A(n41847), .B(n41848), .Z(n39008) );
  AND U39055 ( .A(n41847), .B(n41849), .Z(n41848) );
  XNOR U39056 ( .A(n41850), .B(n41851), .Z(n39011) );
  AND U39057 ( .A(n41850), .B(n41852), .Z(n41851) );
  XNOR U39058 ( .A(n41853), .B(n41854), .Z(n39014) );
  AND U39059 ( .A(n41853), .B(n41855), .Z(n41854) );
  XNOR U39060 ( .A(n41856), .B(n41857), .Z(n39017) );
  AND U39061 ( .A(n41856), .B(n41858), .Z(n41857) );
  XNOR U39062 ( .A(n41859), .B(n41860), .Z(n39020) );
  AND U39063 ( .A(n41859), .B(n41861), .Z(n41860) );
  XNOR U39064 ( .A(n41862), .B(n41863), .Z(n39023) );
  AND U39065 ( .A(n41862), .B(n41864), .Z(n41863) );
  XNOR U39066 ( .A(n41865), .B(n41866), .Z(n39026) );
  AND U39067 ( .A(n41865), .B(n41867), .Z(n41866) );
  XNOR U39068 ( .A(n41868), .B(n41869), .Z(n39029) );
  AND U39069 ( .A(n41868), .B(n41870), .Z(n41869) );
  XNOR U39070 ( .A(n41871), .B(n41872), .Z(n39032) );
  AND U39071 ( .A(n41871), .B(n41873), .Z(n41872) );
  XNOR U39072 ( .A(n41874), .B(n41875), .Z(n39035) );
  AND U39073 ( .A(n41874), .B(n41876), .Z(n41875) );
  XNOR U39074 ( .A(n41877), .B(n41878), .Z(n39038) );
  AND U39075 ( .A(n41877), .B(n41879), .Z(n41878) );
  XNOR U39076 ( .A(n41880), .B(n41881), .Z(n39041) );
  AND U39077 ( .A(n41880), .B(n41882), .Z(n41881) );
  XNOR U39078 ( .A(n41883), .B(n41884), .Z(n39044) );
  AND U39079 ( .A(n41883), .B(n41885), .Z(n41884) );
  XNOR U39080 ( .A(n41886), .B(n41887), .Z(n39047) );
  AND U39081 ( .A(n41886), .B(n41888), .Z(n41887) );
  XNOR U39082 ( .A(n41889), .B(n41890), .Z(n39050) );
  AND U39083 ( .A(n41889), .B(n41891), .Z(n41890) );
  XNOR U39084 ( .A(n41892), .B(n41893), .Z(n39053) );
  AND U39085 ( .A(n41892), .B(n41894), .Z(n41893) );
  XNOR U39086 ( .A(n41895), .B(n41896), .Z(n39056) );
  AND U39087 ( .A(n41895), .B(n41897), .Z(n41896) );
  XNOR U39088 ( .A(n41898), .B(n41899), .Z(n39059) );
  AND U39089 ( .A(n41898), .B(n41900), .Z(n41899) );
  XNOR U39090 ( .A(n41901), .B(n41902), .Z(n39062) );
  AND U39091 ( .A(n41901), .B(n41903), .Z(n41902) );
  XNOR U39092 ( .A(n41904), .B(n41905), .Z(n39065) );
  AND U39093 ( .A(n41904), .B(n41906), .Z(n41905) );
  XNOR U39094 ( .A(n41907), .B(n41908), .Z(n39068) );
  AND U39095 ( .A(n41907), .B(n41909), .Z(n41908) );
  XNOR U39096 ( .A(n41910), .B(n41911), .Z(n39071) );
  AND U39097 ( .A(n41910), .B(n41912), .Z(n41911) );
  XNOR U39098 ( .A(n41913), .B(n41914), .Z(n39074) );
  AND U39099 ( .A(n41913), .B(n41915), .Z(n41914) );
  XNOR U39100 ( .A(n41916), .B(n41917), .Z(n39077) );
  AND U39101 ( .A(n41916), .B(n41918), .Z(n41917) );
  XNOR U39102 ( .A(n41919), .B(n41920), .Z(n39080) );
  AND U39103 ( .A(n41919), .B(n41921), .Z(n41920) );
  XNOR U39104 ( .A(n41922), .B(n41923), .Z(n39083) );
  AND U39105 ( .A(n41922), .B(n41924), .Z(n41923) );
  XNOR U39106 ( .A(n41925), .B(n41926), .Z(n39086) );
  AND U39107 ( .A(n41925), .B(n41927), .Z(n41926) );
  XNOR U39108 ( .A(n41928), .B(n41929), .Z(n39089) );
  AND U39109 ( .A(n41928), .B(n41930), .Z(n41929) );
  XNOR U39110 ( .A(n41931), .B(n41932), .Z(n39092) );
  AND U39111 ( .A(n41931), .B(n41933), .Z(n41932) );
  XNOR U39112 ( .A(n41934), .B(n41935), .Z(n39095) );
  AND U39113 ( .A(n41934), .B(n41936), .Z(n41935) );
  XNOR U39114 ( .A(n41937), .B(n41938), .Z(n39098) );
  AND U39115 ( .A(n41937), .B(n41939), .Z(n41938) );
  XNOR U39116 ( .A(n41940), .B(n41941), .Z(n39101) );
  AND U39117 ( .A(n41940), .B(n41942), .Z(n41941) );
  XNOR U39118 ( .A(n41943), .B(n41944), .Z(n39104) );
  AND U39119 ( .A(n41943), .B(n41945), .Z(n41944) );
  XNOR U39120 ( .A(n41946), .B(n41947), .Z(n39107) );
  AND U39121 ( .A(n41946), .B(n41948), .Z(n41947) );
  XNOR U39122 ( .A(n41949), .B(n41950), .Z(n39110) );
  AND U39123 ( .A(n41949), .B(n41951), .Z(n41950) );
  XNOR U39124 ( .A(n41952), .B(n41953), .Z(n39113) );
  AND U39125 ( .A(n41952), .B(n41954), .Z(n41953) );
  XNOR U39126 ( .A(n41955), .B(n41956), .Z(n39116) );
  AND U39127 ( .A(n41955), .B(n41957), .Z(n41956) );
  XNOR U39128 ( .A(n41958), .B(n41959), .Z(n39119) );
  AND U39129 ( .A(n41958), .B(n41960), .Z(n41959) );
  XNOR U39130 ( .A(n41961), .B(n41962), .Z(n39122) );
  AND U39131 ( .A(n41961), .B(n41963), .Z(n41962) );
  XNOR U39132 ( .A(n41964), .B(n41965), .Z(n39125) );
  AND U39133 ( .A(n41964), .B(n41966), .Z(n41965) );
  XNOR U39134 ( .A(n41967), .B(n41968), .Z(n39128) );
  AND U39135 ( .A(n41967), .B(n41969), .Z(n41968) );
  XNOR U39136 ( .A(n41970), .B(n41971), .Z(n39131) );
  AND U39137 ( .A(n41970), .B(n41972), .Z(n41971) );
  XNOR U39138 ( .A(n41973), .B(n41974), .Z(n39134) );
  AND U39139 ( .A(n41973), .B(n41975), .Z(n41974) );
  XNOR U39140 ( .A(n41976), .B(n41977), .Z(n39137) );
  AND U39141 ( .A(n41976), .B(n41978), .Z(n41977) );
  XNOR U39142 ( .A(n41979), .B(n41980), .Z(n39140) );
  AND U39143 ( .A(n41979), .B(n41981), .Z(n41980) );
  XNOR U39144 ( .A(n41982), .B(n41983), .Z(n39143) );
  AND U39145 ( .A(n41982), .B(n41984), .Z(n41983) );
  XNOR U39146 ( .A(n41985), .B(n41986), .Z(n39146) );
  AND U39147 ( .A(n41985), .B(n41987), .Z(n41986) );
  XNOR U39148 ( .A(n41988), .B(n41989), .Z(n39149) );
  AND U39149 ( .A(n41988), .B(n41990), .Z(n41989) );
  XNOR U39150 ( .A(n41991), .B(n41992), .Z(n39152) );
  AND U39151 ( .A(n41991), .B(n41993), .Z(n41992) );
  XNOR U39152 ( .A(n41994), .B(n41995), .Z(n39155) );
  AND U39153 ( .A(n41994), .B(n41996), .Z(n41995) );
  XNOR U39154 ( .A(n41997), .B(n41998), .Z(n39158) );
  AND U39155 ( .A(n41997), .B(n41999), .Z(n41998) );
  XNOR U39156 ( .A(n42000), .B(n42001), .Z(n39161) );
  AND U39157 ( .A(n42000), .B(n42002), .Z(n42001) );
  XNOR U39158 ( .A(n42003), .B(n42004), .Z(n39164) );
  AND U39159 ( .A(n42003), .B(n42005), .Z(n42004) );
  XNOR U39160 ( .A(n42006), .B(n42007), .Z(n39167) );
  AND U39161 ( .A(n42006), .B(n42008), .Z(n42007) );
  XNOR U39162 ( .A(n42009), .B(n42010), .Z(n39170) );
  AND U39163 ( .A(n42009), .B(n42011), .Z(n42010) );
  XNOR U39164 ( .A(n42012), .B(n42013), .Z(n39173) );
  AND U39165 ( .A(n42012), .B(n42014), .Z(n42013) );
  XNOR U39166 ( .A(n42015), .B(n42016), .Z(n39176) );
  AND U39167 ( .A(n42015), .B(n42017), .Z(n42016) );
  XNOR U39168 ( .A(n42018), .B(n42019), .Z(n39179) );
  AND U39169 ( .A(n42018), .B(n42020), .Z(n42019) );
  XNOR U39170 ( .A(n42021), .B(n42022), .Z(n39182) );
  AND U39171 ( .A(n42021), .B(n42023), .Z(n42022) );
  XNOR U39172 ( .A(n42024), .B(n42025), .Z(n39185) );
  AND U39173 ( .A(n42024), .B(n42026), .Z(n42025) );
  XNOR U39174 ( .A(n42027), .B(n42028), .Z(n39188) );
  AND U39175 ( .A(n42027), .B(n42029), .Z(n42028) );
  XNOR U39176 ( .A(n42030), .B(n42031), .Z(n39191) );
  AND U39177 ( .A(n42030), .B(n42032), .Z(n42031) );
  XNOR U39178 ( .A(n42033), .B(n42034), .Z(n39194) );
  AND U39179 ( .A(n42033), .B(n42035), .Z(n42034) );
  XNOR U39180 ( .A(n42036), .B(n42037), .Z(n39197) );
  AND U39181 ( .A(n42036), .B(n42038), .Z(n42037) );
  XNOR U39182 ( .A(n42039), .B(n42040), .Z(n39200) );
  AND U39183 ( .A(n42039), .B(n42041), .Z(n42040) );
  XNOR U39184 ( .A(n42042), .B(n42043), .Z(n39203) );
  AND U39185 ( .A(n42042), .B(n42044), .Z(n42043) );
  XNOR U39186 ( .A(n42045), .B(n42046), .Z(n39206) );
  AND U39187 ( .A(n42045), .B(n42047), .Z(n42046) );
  XNOR U39188 ( .A(n42048), .B(n42049), .Z(n39209) );
  AND U39189 ( .A(n42048), .B(n42050), .Z(n42049) );
  XNOR U39190 ( .A(n42051), .B(n42052), .Z(n39212) );
  AND U39191 ( .A(n42051), .B(n42053), .Z(n42052) );
  XNOR U39192 ( .A(n42054), .B(n42055), .Z(n39215) );
  AND U39193 ( .A(n42054), .B(n42056), .Z(n42055) );
  XNOR U39194 ( .A(n42057), .B(n42058), .Z(n39218) );
  AND U39195 ( .A(n42057), .B(n42059), .Z(n42058) );
  XNOR U39196 ( .A(n42060), .B(n42061), .Z(n39221) );
  AND U39197 ( .A(n42060), .B(n42062), .Z(n42061) );
  XNOR U39198 ( .A(n42063), .B(n42064), .Z(n39224) );
  AND U39199 ( .A(n42063), .B(n42065), .Z(n42064) );
  XNOR U39200 ( .A(n42066), .B(n42067), .Z(n39227) );
  AND U39201 ( .A(n42066), .B(n42068), .Z(n42067) );
  XNOR U39202 ( .A(n42069), .B(n42070), .Z(n39230) );
  AND U39203 ( .A(n42069), .B(n42071), .Z(n42070) );
  XNOR U39204 ( .A(n42072), .B(n42073), .Z(n39233) );
  AND U39205 ( .A(n42072), .B(n42074), .Z(n42073) );
  XNOR U39206 ( .A(n42075), .B(n42076), .Z(n39236) );
  AND U39207 ( .A(n42075), .B(n42077), .Z(n42076) );
  XNOR U39208 ( .A(n42078), .B(n42079), .Z(n39239) );
  AND U39209 ( .A(n42078), .B(n42080), .Z(n42079) );
  XNOR U39210 ( .A(n42081), .B(n42082), .Z(n39242) );
  AND U39211 ( .A(n42081), .B(n42083), .Z(n42082) );
  XNOR U39212 ( .A(n42084), .B(n42085), .Z(n39245) );
  AND U39213 ( .A(n42084), .B(n42086), .Z(n42085) );
  XNOR U39214 ( .A(n42087), .B(n42088), .Z(n39248) );
  AND U39215 ( .A(n42087), .B(n42089), .Z(n42088) );
  XNOR U39216 ( .A(n42090), .B(n42091), .Z(n39251) );
  AND U39217 ( .A(n42090), .B(n42092), .Z(n42091) );
  XNOR U39218 ( .A(n42093), .B(n42094), .Z(n39254) );
  AND U39219 ( .A(n42093), .B(n42095), .Z(n42094) );
  XNOR U39220 ( .A(n42096), .B(n42097), .Z(n39257) );
  AND U39221 ( .A(n42096), .B(n42098), .Z(n42097) );
  XNOR U39222 ( .A(n42099), .B(n42100), .Z(n39260) );
  AND U39223 ( .A(n42099), .B(n42101), .Z(n42100) );
  XNOR U39224 ( .A(n42102), .B(n42103), .Z(n39263) );
  AND U39225 ( .A(n42102), .B(n42104), .Z(n42103) );
  XNOR U39226 ( .A(n42105), .B(n42106), .Z(n39266) );
  AND U39227 ( .A(n42105), .B(n42107), .Z(n42106) );
  XNOR U39228 ( .A(n42108), .B(n42109), .Z(n39269) );
  AND U39229 ( .A(n42108), .B(n42110), .Z(n42109) );
  XNOR U39230 ( .A(n42111), .B(n42112), .Z(n39272) );
  AND U39231 ( .A(n42111), .B(n42113), .Z(n42112) );
  XNOR U39232 ( .A(n42114), .B(n42115), .Z(n39275) );
  AND U39233 ( .A(n42114), .B(n42116), .Z(n42115) );
  XNOR U39234 ( .A(n42117), .B(n42118), .Z(n39278) );
  AND U39235 ( .A(n42117), .B(n42119), .Z(n42118) );
  XNOR U39236 ( .A(n42120), .B(n42121), .Z(n39281) );
  AND U39237 ( .A(n42120), .B(n42122), .Z(n42121) );
  XNOR U39238 ( .A(n42123), .B(n42124), .Z(n39284) );
  AND U39239 ( .A(n42123), .B(n42125), .Z(n42124) );
  XNOR U39240 ( .A(n42126), .B(n42127), .Z(n39287) );
  AND U39241 ( .A(n42126), .B(n42128), .Z(n42127) );
  XNOR U39242 ( .A(n42129), .B(n42130), .Z(n39290) );
  AND U39243 ( .A(n42129), .B(n42131), .Z(n42130) );
  XNOR U39244 ( .A(n42132), .B(n42133), .Z(n39293) );
  AND U39245 ( .A(n42132), .B(n42134), .Z(n42133) );
  XNOR U39246 ( .A(n42135), .B(n42136), .Z(n39296) );
  AND U39247 ( .A(n42135), .B(n42137), .Z(n42136) );
  XNOR U39248 ( .A(n42138), .B(n42139), .Z(n39299) );
  AND U39249 ( .A(n42138), .B(n42140), .Z(n42139) );
  XNOR U39250 ( .A(n42141), .B(n42142), .Z(n39302) );
  AND U39251 ( .A(n42141), .B(n42143), .Z(n42142) );
  XNOR U39252 ( .A(n42144), .B(n42145), .Z(n39305) );
  AND U39253 ( .A(n42144), .B(n42146), .Z(n42145) );
  XNOR U39254 ( .A(n42147), .B(n42148), .Z(n39308) );
  AND U39255 ( .A(n42147), .B(n42149), .Z(n42148) );
  XNOR U39256 ( .A(n42150), .B(n42151), .Z(n39311) );
  AND U39257 ( .A(n42150), .B(n42152), .Z(n42151) );
  XNOR U39258 ( .A(n42153), .B(n42154), .Z(n39314) );
  AND U39259 ( .A(n42153), .B(n42155), .Z(n42154) );
  XNOR U39260 ( .A(n42156), .B(n42157), .Z(n39317) );
  AND U39261 ( .A(n42156), .B(n42158), .Z(n42157) );
  XNOR U39262 ( .A(n42159), .B(n42160), .Z(n39320) );
  AND U39263 ( .A(n42159), .B(n42161), .Z(n42160) );
  XNOR U39264 ( .A(n42162), .B(n42163), .Z(n39323) );
  AND U39265 ( .A(n42162), .B(n42164), .Z(n42163) );
  XNOR U39266 ( .A(n42165), .B(n42166), .Z(n39326) );
  AND U39267 ( .A(n42165), .B(n42167), .Z(n42166) );
  XNOR U39268 ( .A(n42168), .B(n42169), .Z(n39329) );
  AND U39269 ( .A(n42168), .B(n42170), .Z(n42169) );
  XNOR U39270 ( .A(n42171), .B(n42172), .Z(n39332) );
  AND U39271 ( .A(n42171), .B(n42173), .Z(n42172) );
  XNOR U39272 ( .A(n42174), .B(n42175), .Z(n39335) );
  AND U39273 ( .A(n42174), .B(n42176), .Z(n42175) );
  XNOR U39274 ( .A(n42177), .B(n42178), .Z(n39338) );
  AND U39275 ( .A(n42177), .B(n42179), .Z(n42178) );
  XNOR U39276 ( .A(n42180), .B(n42181), .Z(n39341) );
  AND U39277 ( .A(n42180), .B(n42182), .Z(n42181) );
  XNOR U39278 ( .A(n42183), .B(n42184), .Z(n39344) );
  AND U39279 ( .A(n42183), .B(n42185), .Z(n42184) );
  XNOR U39280 ( .A(n42186), .B(n42187), .Z(n39347) );
  AND U39281 ( .A(n42186), .B(n42188), .Z(n42187) );
  XNOR U39282 ( .A(n42189), .B(n42190), .Z(n39350) );
  AND U39283 ( .A(n42189), .B(n42191), .Z(n42190) );
  XNOR U39284 ( .A(n42192), .B(n42193), .Z(n39353) );
  AND U39285 ( .A(n42192), .B(n42194), .Z(n42193) );
  XNOR U39286 ( .A(n42195), .B(n42196), .Z(n39356) );
  AND U39287 ( .A(n42195), .B(n42197), .Z(n42196) );
  XNOR U39288 ( .A(n42198), .B(n42199), .Z(n39359) );
  AND U39289 ( .A(n42198), .B(n42200), .Z(n42199) );
  XNOR U39290 ( .A(n42201), .B(n42202), .Z(n39362) );
  AND U39291 ( .A(n42201), .B(n42203), .Z(n42202) );
  XNOR U39292 ( .A(n42204), .B(n42205), .Z(n39365) );
  AND U39293 ( .A(n42204), .B(n42206), .Z(n42205) );
  XNOR U39294 ( .A(n42207), .B(n42208), .Z(n39368) );
  AND U39295 ( .A(n42207), .B(n42209), .Z(n42208) );
  XNOR U39296 ( .A(n42210), .B(n42211), .Z(n39371) );
  AND U39297 ( .A(n42210), .B(n42212), .Z(n42211) );
  XNOR U39298 ( .A(n42213), .B(n42214), .Z(n39374) );
  AND U39299 ( .A(n42213), .B(n42215), .Z(n42214) );
  XNOR U39300 ( .A(n42216), .B(n42217), .Z(n39377) );
  AND U39301 ( .A(n42216), .B(n42218), .Z(n42217) );
  XNOR U39302 ( .A(n42219), .B(n42220), .Z(n39380) );
  AND U39303 ( .A(n42219), .B(n42221), .Z(n42220) );
  XNOR U39304 ( .A(n42222), .B(n42223), .Z(n39383) );
  AND U39305 ( .A(n42222), .B(n42224), .Z(n42223) );
  XNOR U39306 ( .A(n42225), .B(n42226), .Z(n39386) );
  AND U39307 ( .A(n42225), .B(n42227), .Z(n42226) );
  XNOR U39308 ( .A(n42228), .B(n42229), .Z(n39389) );
  AND U39309 ( .A(n42228), .B(n42230), .Z(n42229) );
  XNOR U39310 ( .A(n42231), .B(n42232), .Z(n39392) );
  AND U39311 ( .A(n42231), .B(n42233), .Z(n42232) );
  XNOR U39312 ( .A(n42234), .B(n42235), .Z(n39395) );
  AND U39313 ( .A(n42234), .B(n42236), .Z(n42235) );
  XNOR U39314 ( .A(n42237), .B(n42238), .Z(n39398) );
  AND U39315 ( .A(n42237), .B(n42239), .Z(n42238) );
  XNOR U39316 ( .A(n42240), .B(n42241), .Z(n39401) );
  AND U39317 ( .A(n42240), .B(n42242), .Z(n42241) );
  XNOR U39318 ( .A(n42243), .B(n42244), .Z(n39404) );
  AND U39319 ( .A(n42243), .B(n42245), .Z(n42244) );
  XNOR U39320 ( .A(n42246), .B(n42247), .Z(n39407) );
  AND U39321 ( .A(n42246), .B(n42248), .Z(n42247) );
  XNOR U39322 ( .A(n42249), .B(n42250), .Z(n39410) );
  AND U39323 ( .A(n42249), .B(n42251), .Z(n42250) );
  XNOR U39324 ( .A(n42252), .B(n42253), .Z(n39413) );
  AND U39325 ( .A(n42252), .B(n42254), .Z(n42253) );
  XNOR U39326 ( .A(n42255), .B(n42256), .Z(n39416) );
  AND U39327 ( .A(n42255), .B(n42257), .Z(n42256) );
  XNOR U39328 ( .A(n42258), .B(n42259), .Z(n39419) );
  AND U39329 ( .A(n42258), .B(n42260), .Z(n42259) );
  XNOR U39330 ( .A(n42261), .B(n42262), .Z(n39422) );
  AND U39331 ( .A(n42261), .B(n42263), .Z(n42262) );
  XNOR U39332 ( .A(n42264), .B(n42265), .Z(n39425) );
  AND U39333 ( .A(n42264), .B(n42266), .Z(n42265) );
  XNOR U39334 ( .A(n42267), .B(n42268), .Z(n39428) );
  AND U39335 ( .A(n42267), .B(n42269), .Z(n42268) );
  XNOR U39336 ( .A(n42270), .B(n42271), .Z(n39431) );
  AND U39337 ( .A(n42270), .B(n42272), .Z(n42271) );
  XNOR U39338 ( .A(n42273), .B(n42274), .Z(n39434) );
  AND U39339 ( .A(n42273), .B(n42275), .Z(n42274) );
  XNOR U39340 ( .A(n42276), .B(n42277), .Z(n39437) );
  AND U39341 ( .A(n42276), .B(n42278), .Z(n42277) );
  XNOR U39342 ( .A(n42279), .B(n42280), .Z(n39440) );
  AND U39343 ( .A(n42279), .B(n42281), .Z(n42280) );
  XNOR U39344 ( .A(n42282), .B(n42283), .Z(n39443) );
  AND U39345 ( .A(n42282), .B(n42284), .Z(n42283) );
  XNOR U39346 ( .A(n42285), .B(n42286), .Z(n39446) );
  AND U39347 ( .A(n42285), .B(n42287), .Z(n42286) );
  XNOR U39348 ( .A(n42288), .B(n42289), .Z(n39449) );
  AND U39349 ( .A(n42288), .B(n42290), .Z(n42289) );
  XNOR U39350 ( .A(n42291), .B(n42292), .Z(n39452) );
  AND U39351 ( .A(n42291), .B(n42293), .Z(n42292) );
  XNOR U39352 ( .A(n42294), .B(n42295), .Z(n39455) );
  AND U39353 ( .A(n42294), .B(n42296), .Z(n42295) );
  XNOR U39354 ( .A(n42297), .B(n42298), .Z(n39458) );
  AND U39355 ( .A(n42297), .B(n42299), .Z(n42298) );
  XNOR U39356 ( .A(n42300), .B(n42301), .Z(n39461) );
  AND U39357 ( .A(n42300), .B(n42302), .Z(n42301) );
  XNOR U39358 ( .A(n42303), .B(n42304), .Z(n39464) );
  AND U39359 ( .A(n42303), .B(n42305), .Z(n42304) );
  XNOR U39360 ( .A(n42306), .B(n42307), .Z(n39467) );
  AND U39361 ( .A(n42306), .B(n42308), .Z(n42307) );
  XNOR U39362 ( .A(n42309), .B(n42310), .Z(n39470) );
  AND U39363 ( .A(n42309), .B(n42311), .Z(n42310) );
  XNOR U39364 ( .A(n42312), .B(n42313), .Z(n39473) );
  AND U39365 ( .A(n42312), .B(n42314), .Z(n42313) );
  XNOR U39366 ( .A(n42315), .B(n42316), .Z(n39476) );
  AND U39367 ( .A(n42315), .B(n42317), .Z(n42316) );
  XNOR U39368 ( .A(n42318), .B(n42319), .Z(n39479) );
  AND U39369 ( .A(n42318), .B(n42320), .Z(n42319) );
  XNOR U39370 ( .A(n42321), .B(n42322), .Z(n39482) );
  AND U39371 ( .A(n42321), .B(n42323), .Z(n42322) );
  XNOR U39372 ( .A(n42324), .B(n42325), .Z(n39485) );
  AND U39373 ( .A(n42324), .B(n42326), .Z(n42325) );
  XNOR U39374 ( .A(n42327), .B(n42328), .Z(n39488) );
  AND U39375 ( .A(n42327), .B(n42329), .Z(n42328) );
  XNOR U39376 ( .A(n42330), .B(n42331), .Z(n39491) );
  AND U39377 ( .A(n42330), .B(n42332), .Z(n42331) );
  XNOR U39378 ( .A(n42333), .B(n42334), .Z(n39494) );
  AND U39379 ( .A(n42333), .B(n42335), .Z(n42334) );
  XNOR U39380 ( .A(n42336), .B(n42337), .Z(n39497) );
  AND U39381 ( .A(n42336), .B(n42338), .Z(n42337) );
  XNOR U39382 ( .A(n42339), .B(n42340), .Z(n39500) );
  AND U39383 ( .A(n42339), .B(n42341), .Z(n42340) );
  XNOR U39384 ( .A(n42342), .B(n42343), .Z(n39503) );
  AND U39385 ( .A(n42342), .B(n42344), .Z(n42343) );
  XNOR U39386 ( .A(n42345), .B(n42346), .Z(n39506) );
  AND U39387 ( .A(n42345), .B(n42347), .Z(n42346) );
  XNOR U39388 ( .A(n42348), .B(n42349), .Z(n39509) );
  AND U39389 ( .A(n42348), .B(n42350), .Z(n42349) );
  XNOR U39390 ( .A(n42351), .B(n42352), .Z(n39512) );
  AND U39391 ( .A(n42351), .B(n42353), .Z(n42352) );
  XNOR U39392 ( .A(n42354), .B(n42355), .Z(n39515) );
  AND U39393 ( .A(n42354), .B(n42356), .Z(n42355) );
  XNOR U39394 ( .A(n42357), .B(n42358), .Z(n39518) );
  AND U39395 ( .A(n42357), .B(n42359), .Z(n42358) );
  XNOR U39396 ( .A(n42360), .B(n42361), .Z(n39521) );
  AND U39397 ( .A(n42360), .B(n42362), .Z(n42361) );
  XNOR U39398 ( .A(n42363), .B(n42364), .Z(n39524) );
  AND U39399 ( .A(n42363), .B(n42365), .Z(n42364) );
  XNOR U39400 ( .A(n42366), .B(n42367), .Z(n39527) );
  AND U39401 ( .A(n42366), .B(n42368), .Z(n42367) );
  XNOR U39402 ( .A(n42369), .B(n42370), .Z(n39530) );
  AND U39403 ( .A(n42369), .B(n42371), .Z(n42370) );
  XNOR U39404 ( .A(n42372), .B(n42373), .Z(n39533) );
  AND U39405 ( .A(n42372), .B(n42374), .Z(n42373) );
  XNOR U39406 ( .A(n42375), .B(n42376), .Z(n39536) );
  AND U39407 ( .A(n42375), .B(n42377), .Z(n42376) );
  XNOR U39408 ( .A(n42378), .B(n42379), .Z(n39539) );
  AND U39409 ( .A(n42378), .B(n42380), .Z(n42379) );
  XNOR U39410 ( .A(n42381), .B(n42382), .Z(n39542) );
  AND U39411 ( .A(n42381), .B(n42383), .Z(n42382) );
  XNOR U39412 ( .A(n42384), .B(n42385), .Z(n39545) );
  AND U39413 ( .A(n42384), .B(n42386), .Z(n42385) );
  XNOR U39414 ( .A(n42387), .B(n42388), .Z(n39548) );
  AND U39415 ( .A(n42387), .B(n42389), .Z(n42388) );
  XNOR U39416 ( .A(n42390), .B(n42391), .Z(n39551) );
  AND U39417 ( .A(n42390), .B(n42392), .Z(n42391) );
  XNOR U39418 ( .A(n42393), .B(n42394), .Z(n39554) );
  AND U39419 ( .A(n42393), .B(n42395), .Z(n42394) );
  XNOR U39420 ( .A(n42396), .B(n42397), .Z(n39557) );
  AND U39421 ( .A(n42396), .B(n42398), .Z(n42397) );
  XNOR U39422 ( .A(n42399), .B(n42400), .Z(n39560) );
  AND U39423 ( .A(n42399), .B(n42401), .Z(n42400) );
  XNOR U39424 ( .A(n42402), .B(n42403), .Z(n39563) );
  AND U39425 ( .A(n42402), .B(n42404), .Z(n42403) );
  XNOR U39426 ( .A(n42405), .B(n42406), .Z(n39566) );
  AND U39427 ( .A(n42405), .B(n42407), .Z(n42406) );
  XNOR U39428 ( .A(n42408), .B(n42409), .Z(n39569) );
  AND U39429 ( .A(n42408), .B(n42410), .Z(n42409) );
  XNOR U39430 ( .A(n42411), .B(n42412), .Z(n39572) );
  AND U39431 ( .A(n42411), .B(n42413), .Z(n42412) );
  XNOR U39432 ( .A(n42414), .B(n42415), .Z(n39575) );
  AND U39433 ( .A(n42414), .B(n42416), .Z(n42415) );
  XNOR U39434 ( .A(n42417), .B(n42418), .Z(n39578) );
  AND U39435 ( .A(n42417), .B(n42419), .Z(n42418) );
  XNOR U39436 ( .A(n42420), .B(n42421), .Z(n39581) );
  AND U39437 ( .A(n42420), .B(n42422), .Z(n42421) );
  XNOR U39438 ( .A(n42423), .B(n42424), .Z(n39584) );
  AND U39439 ( .A(n42423), .B(n42425), .Z(n42424) );
  XNOR U39440 ( .A(n42426), .B(n42427), .Z(n39587) );
  AND U39441 ( .A(n42426), .B(n42428), .Z(n42427) );
  XNOR U39442 ( .A(n42429), .B(n42430), .Z(n39590) );
  AND U39443 ( .A(n42429), .B(n42431), .Z(n42430) );
  XNOR U39444 ( .A(n42432), .B(n42433), .Z(n39593) );
  AND U39445 ( .A(n42432), .B(n42434), .Z(n42433) );
  XNOR U39446 ( .A(n42435), .B(n42436), .Z(n39596) );
  AND U39447 ( .A(n42435), .B(n42437), .Z(n42436) );
  XNOR U39448 ( .A(n42438), .B(n42439), .Z(n39599) );
  AND U39449 ( .A(n42438), .B(n42440), .Z(n42439) );
  XNOR U39450 ( .A(n42441), .B(n42442), .Z(n39602) );
  AND U39451 ( .A(n42441), .B(n42443), .Z(n42442) );
  XNOR U39452 ( .A(n42444), .B(n42445), .Z(n39605) );
  AND U39453 ( .A(n42444), .B(n42446), .Z(n42445) );
  XNOR U39454 ( .A(n42447), .B(n42448), .Z(n39608) );
  AND U39455 ( .A(n42447), .B(n42449), .Z(n42448) );
  XNOR U39456 ( .A(n42450), .B(n42451), .Z(n39611) );
  AND U39457 ( .A(n42450), .B(n42452), .Z(n42451) );
  XNOR U39458 ( .A(n42453), .B(n42454), .Z(n39614) );
  AND U39459 ( .A(n42453), .B(n42455), .Z(n42454) );
  XNOR U39460 ( .A(n42456), .B(n42457), .Z(n39617) );
  AND U39461 ( .A(n42456), .B(n42458), .Z(n42457) );
  XNOR U39462 ( .A(n42459), .B(n42460), .Z(n39620) );
  AND U39463 ( .A(n42459), .B(n42461), .Z(n42460) );
  XNOR U39464 ( .A(n42462), .B(n42463), .Z(n39623) );
  AND U39465 ( .A(n42462), .B(n42464), .Z(n42463) );
  XNOR U39466 ( .A(n42465), .B(n42466), .Z(n39626) );
  AND U39467 ( .A(n42465), .B(n42467), .Z(n42466) );
  XNOR U39468 ( .A(n42468), .B(n42469), .Z(n39629) );
  AND U39469 ( .A(n42468), .B(n42470), .Z(n42469) );
  XNOR U39470 ( .A(n42471), .B(n42472), .Z(n39632) );
  AND U39471 ( .A(n42471), .B(n42473), .Z(n42472) );
  XNOR U39472 ( .A(n42474), .B(n42475), .Z(n39635) );
  AND U39473 ( .A(n42474), .B(n42476), .Z(n42475) );
  XNOR U39474 ( .A(n42477), .B(n42478), .Z(n39638) );
  AND U39475 ( .A(n42477), .B(n42479), .Z(n42478) );
  XNOR U39476 ( .A(n42480), .B(n42481), .Z(n39641) );
  AND U39477 ( .A(n42480), .B(n42482), .Z(n42481) );
  XNOR U39478 ( .A(n42483), .B(n42484), .Z(n39644) );
  AND U39479 ( .A(n42483), .B(n42485), .Z(n42484) );
  XNOR U39480 ( .A(n42486), .B(n42487), .Z(n39647) );
  AND U39481 ( .A(n42486), .B(n42488), .Z(n42487) );
  XNOR U39482 ( .A(n42489), .B(n42490), .Z(n39650) );
  AND U39483 ( .A(n42489), .B(n42491), .Z(n42490) );
  XNOR U39484 ( .A(n42492), .B(n42493), .Z(n39653) );
  AND U39485 ( .A(n42492), .B(n42494), .Z(n42493) );
  XNOR U39486 ( .A(n42495), .B(n42496), .Z(n39656) );
  AND U39487 ( .A(n42495), .B(n42497), .Z(n42496) );
  XNOR U39488 ( .A(n42498), .B(n42499), .Z(n39659) );
  AND U39489 ( .A(n42498), .B(n42500), .Z(n42499) );
  XNOR U39490 ( .A(n42501), .B(n42502), .Z(n39662) );
  AND U39491 ( .A(n42501), .B(n42503), .Z(n42502) );
  XNOR U39492 ( .A(n42504), .B(n42505), .Z(n39665) );
  AND U39493 ( .A(n42504), .B(n42506), .Z(n42505) );
  XNOR U39494 ( .A(n42507), .B(n42508), .Z(n39668) );
  AND U39495 ( .A(n42507), .B(n42509), .Z(n42508) );
  XNOR U39496 ( .A(n42510), .B(n42511), .Z(n39671) );
  AND U39497 ( .A(n42510), .B(n42512), .Z(n42511) );
  XNOR U39498 ( .A(n42513), .B(n42514), .Z(n39674) );
  AND U39499 ( .A(n42513), .B(n42515), .Z(n42514) );
  XNOR U39500 ( .A(n42516), .B(n42517), .Z(n39677) );
  AND U39501 ( .A(n42516), .B(n42518), .Z(n42517) );
  XNOR U39502 ( .A(n42519), .B(n42520), .Z(n39680) );
  AND U39503 ( .A(n42519), .B(n42521), .Z(n42520) );
  XNOR U39504 ( .A(n42522), .B(n42523), .Z(n39683) );
  AND U39505 ( .A(n42522), .B(n42524), .Z(n42523) );
  XNOR U39506 ( .A(n42525), .B(n42526), .Z(n39686) );
  AND U39507 ( .A(n42525), .B(n42527), .Z(n42526) );
  XNOR U39508 ( .A(n42528), .B(n42529), .Z(n39689) );
  AND U39509 ( .A(n42528), .B(n42530), .Z(n42529) );
  XNOR U39510 ( .A(n42531), .B(n42532), .Z(n39692) );
  AND U39511 ( .A(n42531), .B(n42533), .Z(n42532) );
  XNOR U39512 ( .A(n42534), .B(n42535), .Z(n39695) );
  AND U39513 ( .A(n42534), .B(n42536), .Z(n42535) );
  XNOR U39514 ( .A(n42537), .B(n42538), .Z(n39698) );
  AND U39515 ( .A(n42537), .B(n42539), .Z(n42538) );
  XNOR U39516 ( .A(n42540), .B(n42541), .Z(n39701) );
  AND U39517 ( .A(n42540), .B(n42542), .Z(n42541) );
  XNOR U39518 ( .A(n42543), .B(n42544), .Z(n39704) );
  AND U39519 ( .A(n42543), .B(n42545), .Z(n42544) );
  XNOR U39520 ( .A(n42546), .B(n42547), .Z(n39707) );
  AND U39521 ( .A(n42546), .B(n42548), .Z(n42547) );
  XNOR U39522 ( .A(n42549), .B(n42550), .Z(n39710) );
  AND U39523 ( .A(n42549), .B(n42551), .Z(n42550) );
  XNOR U39524 ( .A(n42552), .B(n42553), .Z(n39713) );
  AND U39525 ( .A(n42552), .B(n42554), .Z(n42553) );
  XNOR U39526 ( .A(n42555), .B(n42556), .Z(n39716) );
  AND U39527 ( .A(n42555), .B(n42557), .Z(n42556) );
  XNOR U39528 ( .A(n42558), .B(n42559), .Z(n39719) );
  AND U39529 ( .A(n42558), .B(n42560), .Z(n42559) );
  XNOR U39530 ( .A(n42561), .B(n42562), .Z(n39722) );
  AND U39531 ( .A(n42561), .B(n42563), .Z(n42562) );
  XNOR U39532 ( .A(n42564), .B(n42565), .Z(n39725) );
  AND U39533 ( .A(n42564), .B(n42566), .Z(n42565) );
  XNOR U39534 ( .A(n42567), .B(n42568), .Z(n39728) );
  AND U39535 ( .A(n42567), .B(n42569), .Z(n42568) );
  XNOR U39536 ( .A(n42570), .B(n42571), .Z(n39731) );
  AND U39537 ( .A(n42570), .B(n42572), .Z(n42571) );
  XNOR U39538 ( .A(n42573), .B(n42574), .Z(n39734) );
  AND U39539 ( .A(n42573), .B(n42575), .Z(n42574) );
  XNOR U39540 ( .A(n42576), .B(n42577), .Z(n39737) );
  AND U39541 ( .A(n42576), .B(n42578), .Z(n42577) );
  XNOR U39542 ( .A(n42579), .B(n42580), .Z(n39740) );
  AND U39543 ( .A(n42579), .B(n42581), .Z(n42580) );
  XNOR U39544 ( .A(n42582), .B(n42583), .Z(n39743) );
  AND U39545 ( .A(n42582), .B(n42584), .Z(n42583) );
  XNOR U39546 ( .A(n42585), .B(n42586), .Z(n39746) );
  AND U39547 ( .A(n42585), .B(n42587), .Z(n42586) );
  XNOR U39548 ( .A(n42588), .B(n42589), .Z(n39749) );
  AND U39549 ( .A(n42588), .B(n42590), .Z(n42589) );
  XNOR U39550 ( .A(n42591), .B(n42592), .Z(n39752) );
  AND U39551 ( .A(n42591), .B(n42593), .Z(n42592) );
  XNOR U39552 ( .A(n42594), .B(n42595), .Z(n39755) );
  AND U39553 ( .A(n42594), .B(n42596), .Z(n42595) );
  XNOR U39554 ( .A(n42597), .B(n42598), .Z(n39758) );
  AND U39555 ( .A(n42597), .B(n42599), .Z(n42598) );
  XNOR U39556 ( .A(n42600), .B(n42601), .Z(n39761) );
  AND U39557 ( .A(n42600), .B(n42602), .Z(n42601) );
  XNOR U39558 ( .A(n42603), .B(n42604), .Z(n39764) );
  AND U39559 ( .A(n42603), .B(n42605), .Z(n42604) );
  XNOR U39560 ( .A(n42606), .B(n42607), .Z(n39767) );
  AND U39561 ( .A(n42606), .B(n42608), .Z(n42607) );
  XNOR U39562 ( .A(n42609), .B(n42610), .Z(n39770) );
  AND U39563 ( .A(n42609), .B(n42611), .Z(n42610) );
  XNOR U39564 ( .A(n42612), .B(n42613), .Z(n39773) );
  AND U39565 ( .A(n42612), .B(n42614), .Z(n42613) );
  XNOR U39566 ( .A(n42615), .B(n42616), .Z(n39776) );
  AND U39567 ( .A(n42615), .B(n42617), .Z(n42616) );
  XNOR U39568 ( .A(n42618), .B(n42619), .Z(n39779) );
  AND U39569 ( .A(n42618), .B(n42620), .Z(n42619) );
  XNOR U39570 ( .A(n42621), .B(n42622), .Z(n39782) );
  AND U39571 ( .A(n42621), .B(n42623), .Z(n42622) );
  XNOR U39572 ( .A(n42624), .B(n42625), .Z(n39785) );
  AND U39573 ( .A(n42624), .B(n42626), .Z(n42625) );
  XNOR U39574 ( .A(n42627), .B(n42628), .Z(n39788) );
  AND U39575 ( .A(n42627), .B(n42629), .Z(n42628) );
  XNOR U39576 ( .A(n42630), .B(n42631), .Z(n39791) );
  AND U39577 ( .A(n42630), .B(n42632), .Z(n42631) );
  XNOR U39578 ( .A(n42633), .B(n42634), .Z(n39794) );
  AND U39579 ( .A(n42633), .B(n42635), .Z(n42634) );
  XNOR U39580 ( .A(n42636), .B(n42637), .Z(n39797) );
  AND U39581 ( .A(n42636), .B(n42638), .Z(n42637) );
  XNOR U39582 ( .A(n42639), .B(n42640), .Z(n39800) );
  AND U39583 ( .A(n42639), .B(n42641), .Z(n42640) );
  XNOR U39584 ( .A(n42642), .B(n42643), .Z(n39803) );
  AND U39585 ( .A(n42642), .B(n42644), .Z(n42643) );
  IV U39586 ( .A(n39808), .Z(n39806) );
  XNOR U39587 ( .A(n42645), .B(n42646), .Z(n39808) );
  AND U39588 ( .A(n42645), .B(n135), .Z(n42646) );
  XOR U39589 ( .A(n42647), .B(n42648), .Z(n39809) );
  AND U39590 ( .A(n42649), .B(n42650), .Z(n42648) );
  XOR U39591 ( .A(n139), .B(n42647), .Z(n42650) );
  XOR U39592 ( .A(n41227), .B(n41228), .Z(n139) );
  AND U39593 ( .A(n42651), .B(n42652), .Z(n41228) );
  XOR U39594 ( .A(n41224), .B(n41225), .Z(n41227) );
  AND U39595 ( .A(n42653), .B(n42654), .Z(n41225) );
  XOR U39596 ( .A(n41221), .B(n41222), .Z(n41224) );
  AND U39597 ( .A(n42655), .B(n42656), .Z(n41222) );
  XOR U39598 ( .A(n41218), .B(n41219), .Z(n41221) );
  AND U39599 ( .A(n42657), .B(n42658), .Z(n41219) );
  XOR U39600 ( .A(n41215), .B(n41216), .Z(n41218) );
  AND U39601 ( .A(n42659), .B(n42660), .Z(n41216) );
  XOR U39602 ( .A(n41212), .B(n41213), .Z(n41215) );
  AND U39603 ( .A(n42661), .B(n42662), .Z(n41213) );
  XOR U39604 ( .A(n41209), .B(n41210), .Z(n41212) );
  AND U39605 ( .A(n42663), .B(n42664), .Z(n41210) );
  XOR U39606 ( .A(n41206), .B(n41207), .Z(n41209) );
  AND U39607 ( .A(n42665), .B(n42666), .Z(n41207) );
  XOR U39608 ( .A(n41203), .B(n41204), .Z(n41206) );
  AND U39609 ( .A(n42667), .B(n42668), .Z(n41204) );
  XOR U39610 ( .A(n41200), .B(n41201), .Z(n41203) );
  AND U39611 ( .A(n42669), .B(n42670), .Z(n41201) );
  XOR U39612 ( .A(n41197), .B(n41198), .Z(n41200) );
  AND U39613 ( .A(n42671), .B(n42672), .Z(n41198) );
  XOR U39614 ( .A(n41194), .B(n41195), .Z(n41197) );
  AND U39615 ( .A(n42673), .B(n42674), .Z(n41195) );
  XOR U39616 ( .A(n41191), .B(n41192), .Z(n41194) );
  AND U39617 ( .A(n42675), .B(n42676), .Z(n41192) );
  XOR U39618 ( .A(n41188), .B(n41189), .Z(n41191) );
  AND U39619 ( .A(n42677), .B(n42678), .Z(n41189) );
  XOR U39620 ( .A(n41185), .B(n41186), .Z(n41188) );
  AND U39621 ( .A(n42679), .B(n42680), .Z(n41186) );
  XOR U39622 ( .A(n41182), .B(n41183), .Z(n41185) );
  AND U39623 ( .A(n42681), .B(n42682), .Z(n41183) );
  XOR U39624 ( .A(n41179), .B(n41180), .Z(n41182) );
  AND U39625 ( .A(n42683), .B(n42684), .Z(n41180) );
  XOR U39626 ( .A(n41176), .B(n41177), .Z(n41179) );
  AND U39627 ( .A(n42685), .B(n42686), .Z(n41177) );
  XOR U39628 ( .A(n41173), .B(n41174), .Z(n41176) );
  AND U39629 ( .A(n42687), .B(n42688), .Z(n41174) );
  XOR U39630 ( .A(n41170), .B(n41171), .Z(n41173) );
  AND U39631 ( .A(n42689), .B(n42690), .Z(n41171) );
  XOR U39632 ( .A(n41167), .B(n41168), .Z(n41170) );
  AND U39633 ( .A(n42691), .B(n42692), .Z(n41168) );
  XOR U39634 ( .A(n41164), .B(n41165), .Z(n41167) );
  AND U39635 ( .A(n42693), .B(n42694), .Z(n41165) );
  XOR U39636 ( .A(n41161), .B(n41162), .Z(n41164) );
  AND U39637 ( .A(n42695), .B(n42696), .Z(n41162) );
  XOR U39638 ( .A(n41158), .B(n41159), .Z(n41161) );
  AND U39639 ( .A(n42697), .B(n42698), .Z(n41159) );
  XOR U39640 ( .A(n41155), .B(n41156), .Z(n41158) );
  AND U39641 ( .A(n42699), .B(n42700), .Z(n41156) );
  XOR U39642 ( .A(n41152), .B(n41153), .Z(n41155) );
  AND U39643 ( .A(n42701), .B(n42702), .Z(n41153) );
  XOR U39644 ( .A(n41149), .B(n41150), .Z(n41152) );
  AND U39645 ( .A(n42703), .B(n42704), .Z(n41150) );
  XOR U39646 ( .A(n41146), .B(n41147), .Z(n41149) );
  AND U39647 ( .A(n42705), .B(n42706), .Z(n41147) );
  XOR U39648 ( .A(n41143), .B(n41144), .Z(n41146) );
  AND U39649 ( .A(n42707), .B(n42708), .Z(n41144) );
  XOR U39650 ( .A(n41140), .B(n41141), .Z(n41143) );
  AND U39651 ( .A(n42709), .B(n42710), .Z(n41141) );
  XOR U39652 ( .A(n41137), .B(n41138), .Z(n41140) );
  AND U39653 ( .A(n42711), .B(n42712), .Z(n41138) );
  XOR U39654 ( .A(n41134), .B(n41135), .Z(n41137) );
  AND U39655 ( .A(n42713), .B(n42714), .Z(n41135) );
  XOR U39656 ( .A(n41131), .B(n41132), .Z(n41134) );
  AND U39657 ( .A(n42715), .B(n42716), .Z(n41132) );
  XOR U39658 ( .A(n41128), .B(n41129), .Z(n41131) );
  AND U39659 ( .A(n42717), .B(n42718), .Z(n41129) );
  XOR U39660 ( .A(n41125), .B(n41126), .Z(n41128) );
  AND U39661 ( .A(n42719), .B(n42720), .Z(n41126) );
  XOR U39662 ( .A(n41122), .B(n41123), .Z(n41125) );
  AND U39663 ( .A(n42721), .B(n42722), .Z(n41123) );
  XOR U39664 ( .A(n41119), .B(n41120), .Z(n41122) );
  AND U39665 ( .A(n42723), .B(n42724), .Z(n41120) );
  XOR U39666 ( .A(n41116), .B(n41117), .Z(n41119) );
  AND U39667 ( .A(n42725), .B(n42726), .Z(n41117) );
  XOR U39668 ( .A(n41113), .B(n41114), .Z(n41116) );
  AND U39669 ( .A(n42727), .B(n42728), .Z(n41114) );
  XOR U39670 ( .A(n41110), .B(n41111), .Z(n41113) );
  AND U39671 ( .A(n42729), .B(n42730), .Z(n41111) );
  XOR U39672 ( .A(n41107), .B(n41108), .Z(n41110) );
  AND U39673 ( .A(n42731), .B(n42732), .Z(n41108) );
  XOR U39674 ( .A(n41104), .B(n41105), .Z(n41107) );
  AND U39675 ( .A(n42733), .B(n42734), .Z(n41105) );
  XOR U39676 ( .A(n41101), .B(n41102), .Z(n41104) );
  AND U39677 ( .A(n42735), .B(n42736), .Z(n41102) );
  XOR U39678 ( .A(n41098), .B(n41099), .Z(n41101) );
  AND U39679 ( .A(n42737), .B(n42738), .Z(n41099) );
  XOR U39680 ( .A(n41095), .B(n41096), .Z(n41098) );
  AND U39681 ( .A(n42739), .B(n42740), .Z(n41096) );
  XOR U39682 ( .A(n41092), .B(n41093), .Z(n41095) );
  AND U39683 ( .A(n42741), .B(n42742), .Z(n41093) );
  XOR U39684 ( .A(n41089), .B(n41090), .Z(n41092) );
  AND U39685 ( .A(n42743), .B(n42744), .Z(n41090) );
  XOR U39686 ( .A(n41086), .B(n41087), .Z(n41089) );
  AND U39687 ( .A(n42745), .B(n42746), .Z(n41087) );
  XOR U39688 ( .A(n41083), .B(n41084), .Z(n41086) );
  AND U39689 ( .A(n42747), .B(n42748), .Z(n41084) );
  XOR U39690 ( .A(n41080), .B(n41081), .Z(n41083) );
  AND U39691 ( .A(n42749), .B(n42750), .Z(n41081) );
  XOR U39692 ( .A(n41077), .B(n41078), .Z(n41080) );
  AND U39693 ( .A(n42751), .B(n42752), .Z(n41078) );
  XOR U39694 ( .A(n41074), .B(n41075), .Z(n41077) );
  AND U39695 ( .A(n42753), .B(n42754), .Z(n41075) );
  XOR U39696 ( .A(n41071), .B(n41072), .Z(n41074) );
  AND U39697 ( .A(n42755), .B(n42756), .Z(n41072) );
  XOR U39698 ( .A(n41068), .B(n41069), .Z(n41071) );
  AND U39699 ( .A(n42757), .B(n42758), .Z(n41069) );
  XOR U39700 ( .A(n41065), .B(n41066), .Z(n41068) );
  AND U39701 ( .A(n42759), .B(n42760), .Z(n41066) );
  XOR U39702 ( .A(n41062), .B(n41063), .Z(n41065) );
  AND U39703 ( .A(n42761), .B(n42762), .Z(n41063) );
  XOR U39704 ( .A(n41059), .B(n41060), .Z(n41062) );
  AND U39705 ( .A(n42763), .B(n42764), .Z(n41060) );
  XOR U39706 ( .A(n41056), .B(n41057), .Z(n41059) );
  AND U39707 ( .A(n42765), .B(n42766), .Z(n41057) );
  XOR U39708 ( .A(n41053), .B(n41054), .Z(n41056) );
  AND U39709 ( .A(n42767), .B(n42768), .Z(n41054) );
  XOR U39710 ( .A(n41050), .B(n41051), .Z(n41053) );
  AND U39711 ( .A(n42769), .B(n42770), .Z(n41051) );
  XOR U39712 ( .A(n41047), .B(n41048), .Z(n41050) );
  AND U39713 ( .A(n42771), .B(n42772), .Z(n41048) );
  XOR U39714 ( .A(n41044), .B(n41045), .Z(n41047) );
  AND U39715 ( .A(n42773), .B(n42774), .Z(n41045) );
  XOR U39716 ( .A(n41041), .B(n41042), .Z(n41044) );
  AND U39717 ( .A(n42775), .B(n42776), .Z(n41042) );
  XOR U39718 ( .A(n41038), .B(n41039), .Z(n41041) );
  AND U39719 ( .A(n42777), .B(n42778), .Z(n41039) );
  XOR U39720 ( .A(n41035), .B(n41036), .Z(n41038) );
  AND U39721 ( .A(n42779), .B(n42780), .Z(n41036) );
  XOR U39722 ( .A(n41032), .B(n41033), .Z(n41035) );
  AND U39723 ( .A(n42781), .B(n42782), .Z(n41033) );
  XOR U39724 ( .A(n41029), .B(n41030), .Z(n41032) );
  AND U39725 ( .A(n42783), .B(n42784), .Z(n41030) );
  XOR U39726 ( .A(n41026), .B(n41027), .Z(n41029) );
  AND U39727 ( .A(n42785), .B(n42786), .Z(n41027) );
  XOR U39728 ( .A(n41023), .B(n41024), .Z(n41026) );
  AND U39729 ( .A(n42787), .B(n42788), .Z(n41024) );
  XOR U39730 ( .A(n41020), .B(n41021), .Z(n41023) );
  AND U39731 ( .A(n42789), .B(n42790), .Z(n41021) );
  XOR U39732 ( .A(n41017), .B(n41018), .Z(n41020) );
  AND U39733 ( .A(n42791), .B(n42792), .Z(n41018) );
  XOR U39734 ( .A(n41014), .B(n41015), .Z(n41017) );
  AND U39735 ( .A(n42793), .B(n42794), .Z(n41015) );
  XOR U39736 ( .A(n41011), .B(n41012), .Z(n41014) );
  AND U39737 ( .A(n42795), .B(n42796), .Z(n41012) );
  XOR U39738 ( .A(n41008), .B(n41009), .Z(n41011) );
  AND U39739 ( .A(n42797), .B(n42798), .Z(n41009) );
  XOR U39740 ( .A(n41005), .B(n41006), .Z(n41008) );
  AND U39741 ( .A(n42799), .B(n42800), .Z(n41006) );
  XOR U39742 ( .A(n41002), .B(n41003), .Z(n41005) );
  AND U39743 ( .A(n42801), .B(n42802), .Z(n41003) );
  XOR U39744 ( .A(n40999), .B(n41000), .Z(n41002) );
  AND U39745 ( .A(n42803), .B(n42804), .Z(n41000) );
  XOR U39746 ( .A(n40996), .B(n40997), .Z(n40999) );
  AND U39747 ( .A(n42805), .B(n42806), .Z(n40997) );
  XOR U39748 ( .A(n40993), .B(n40994), .Z(n40996) );
  AND U39749 ( .A(n42807), .B(n42808), .Z(n40994) );
  XOR U39750 ( .A(n40990), .B(n40991), .Z(n40993) );
  AND U39751 ( .A(n42809), .B(n42810), .Z(n40991) );
  XOR U39752 ( .A(n40987), .B(n40988), .Z(n40990) );
  AND U39753 ( .A(n42811), .B(n42812), .Z(n40988) );
  XOR U39754 ( .A(n40984), .B(n40985), .Z(n40987) );
  AND U39755 ( .A(n42813), .B(n42814), .Z(n40985) );
  XOR U39756 ( .A(n40981), .B(n40982), .Z(n40984) );
  AND U39757 ( .A(n42815), .B(n42816), .Z(n40982) );
  XOR U39758 ( .A(n40978), .B(n40979), .Z(n40981) );
  AND U39759 ( .A(n42817), .B(n42818), .Z(n40979) );
  XOR U39760 ( .A(n40975), .B(n40976), .Z(n40978) );
  AND U39761 ( .A(n42819), .B(n42820), .Z(n40976) );
  XOR U39762 ( .A(n40972), .B(n40973), .Z(n40975) );
  AND U39763 ( .A(n42821), .B(n42822), .Z(n40973) );
  XOR U39764 ( .A(n40969), .B(n40970), .Z(n40972) );
  AND U39765 ( .A(n42823), .B(n42824), .Z(n40970) );
  XOR U39766 ( .A(n40966), .B(n40967), .Z(n40969) );
  AND U39767 ( .A(n42825), .B(n42826), .Z(n40967) );
  XOR U39768 ( .A(n40963), .B(n40964), .Z(n40966) );
  AND U39769 ( .A(n42827), .B(n42828), .Z(n40964) );
  XOR U39770 ( .A(n40960), .B(n40961), .Z(n40963) );
  AND U39771 ( .A(n42829), .B(n42830), .Z(n40961) );
  XOR U39772 ( .A(n40957), .B(n40958), .Z(n40960) );
  AND U39773 ( .A(n42831), .B(n42832), .Z(n40958) );
  XOR U39774 ( .A(n40954), .B(n40955), .Z(n40957) );
  AND U39775 ( .A(n42833), .B(n42834), .Z(n40955) );
  XOR U39776 ( .A(n40951), .B(n40952), .Z(n40954) );
  AND U39777 ( .A(n42835), .B(n42836), .Z(n40952) );
  XOR U39778 ( .A(n40948), .B(n40949), .Z(n40951) );
  AND U39779 ( .A(n42837), .B(n42838), .Z(n40949) );
  XOR U39780 ( .A(n40945), .B(n40946), .Z(n40948) );
  AND U39781 ( .A(n42839), .B(n42840), .Z(n40946) );
  XOR U39782 ( .A(n40942), .B(n40943), .Z(n40945) );
  AND U39783 ( .A(n42841), .B(n42842), .Z(n40943) );
  XOR U39784 ( .A(n40939), .B(n40940), .Z(n40942) );
  AND U39785 ( .A(n42843), .B(n42844), .Z(n40940) );
  XOR U39786 ( .A(n40936), .B(n40937), .Z(n40939) );
  AND U39787 ( .A(n42845), .B(n42846), .Z(n40937) );
  XOR U39788 ( .A(n40933), .B(n40934), .Z(n40936) );
  AND U39789 ( .A(n42847), .B(n42848), .Z(n40934) );
  XOR U39790 ( .A(n40930), .B(n40931), .Z(n40933) );
  AND U39791 ( .A(n42849), .B(n42850), .Z(n40931) );
  XOR U39792 ( .A(n40927), .B(n40928), .Z(n40930) );
  AND U39793 ( .A(n42851), .B(n42852), .Z(n40928) );
  XOR U39794 ( .A(n40924), .B(n40925), .Z(n40927) );
  AND U39795 ( .A(n42853), .B(n42854), .Z(n40925) );
  XOR U39796 ( .A(n40921), .B(n40922), .Z(n40924) );
  AND U39797 ( .A(n42855), .B(n42856), .Z(n40922) );
  XOR U39798 ( .A(n40918), .B(n40919), .Z(n40921) );
  AND U39799 ( .A(n42857), .B(n42858), .Z(n40919) );
  XOR U39800 ( .A(n40915), .B(n40916), .Z(n40918) );
  AND U39801 ( .A(n42859), .B(n42860), .Z(n40916) );
  XOR U39802 ( .A(n40912), .B(n40913), .Z(n40915) );
  AND U39803 ( .A(n42861), .B(n42862), .Z(n40913) );
  XOR U39804 ( .A(n40909), .B(n40910), .Z(n40912) );
  AND U39805 ( .A(n42863), .B(n42864), .Z(n40910) );
  XOR U39806 ( .A(n40906), .B(n40907), .Z(n40909) );
  AND U39807 ( .A(n42865), .B(n42866), .Z(n40907) );
  XOR U39808 ( .A(n40903), .B(n40904), .Z(n40906) );
  AND U39809 ( .A(n42867), .B(n42868), .Z(n40904) );
  XOR U39810 ( .A(n40900), .B(n40901), .Z(n40903) );
  AND U39811 ( .A(n42869), .B(n42870), .Z(n40901) );
  XOR U39812 ( .A(n40897), .B(n40898), .Z(n40900) );
  AND U39813 ( .A(n42871), .B(n42872), .Z(n40898) );
  XOR U39814 ( .A(n40894), .B(n40895), .Z(n40897) );
  AND U39815 ( .A(n42873), .B(n42874), .Z(n40895) );
  XOR U39816 ( .A(n40891), .B(n40892), .Z(n40894) );
  AND U39817 ( .A(n42875), .B(n42876), .Z(n40892) );
  XOR U39818 ( .A(n40888), .B(n40889), .Z(n40891) );
  AND U39819 ( .A(n42877), .B(n42878), .Z(n40889) );
  XOR U39820 ( .A(n40885), .B(n40886), .Z(n40888) );
  AND U39821 ( .A(n42879), .B(n42880), .Z(n40886) );
  XOR U39822 ( .A(n40882), .B(n40883), .Z(n40885) );
  AND U39823 ( .A(n42881), .B(n42882), .Z(n40883) );
  XOR U39824 ( .A(n40879), .B(n40880), .Z(n40882) );
  AND U39825 ( .A(n42883), .B(n42884), .Z(n40880) );
  XOR U39826 ( .A(n40876), .B(n40877), .Z(n40879) );
  AND U39827 ( .A(n42885), .B(n42886), .Z(n40877) );
  XOR U39828 ( .A(n40873), .B(n40874), .Z(n40876) );
  AND U39829 ( .A(n42887), .B(n42888), .Z(n40874) );
  XOR U39830 ( .A(n40870), .B(n40871), .Z(n40873) );
  AND U39831 ( .A(n42889), .B(n42890), .Z(n40871) );
  XOR U39832 ( .A(n40867), .B(n40868), .Z(n40870) );
  AND U39833 ( .A(n42891), .B(n42892), .Z(n40868) );
  XOR U39834 ( .A(n40864), .B(n40865), .Z(n40867) );
  AND U39835 ( .A(n42893), .B(n42894), .Z(n40865) );
  XOR U39836 ( .A(n40861), .B(n40862), .Z(n40864) );
  AND U39837 ( .A(n42895), .B(n42896), .Z(n40862) );
  XOR U39838 ( .A(n40858), .B(n40859), .Z(n40861) );
  AND U39839 ( .A(n42897), .B(n42898), .Z(n40859) );
  XOR U39840 ( .A(n40855), .B(n40856), .Z(n40858) );
  AND U39841 ( .A(n42899), .B(n42900), .Z(n40856) );
  XOR U39842 ( .A(n40852), .B(n40853), .Z(n40855) );
  AND U39843 ( .A(n42901), .B(n42902), .Z(n40853) );
  XOR U39844 ( .A(n40849), .B(n40850), .Z(n40852) );
  AND U39845 ( .A(n42903), .B(n42904), .Z(n40850) );
  XOR U39846 ( .A(n40846), .B(n40847), .Z(n40849) );
  AND U39847 ( .A(n42905), .B(n42906), .Z(n40847) );
  XOR U39848 ( .A(n40843), .B(n40844), .Z(n40846) );
  AND U39849 ( .A(n42907), .B(n42908), .Z(n40844) );
  XOR U39850 ( .A(n40840), .B(n40841), .Z(n40843) );
  AND U39851 ( .A(n42909), .B(n42910), .Z(n40841) );
  XOR U39852 ( .A(n40837), .B(n40838), .Z(n40840) );
  AND U39853 ( .A(n42911), .B(n42912), .Z(n40838) );
  XOR U39854 ( .A(n40834), .B(n40835), .Z(n40837) );
  AND U39855 ( .A(n42913), .B(n42914), .Z(n40835) );
  XOR U39856 ( .A(n40831), .B(n40832), .Z(n40834) );
  AND U39857 ( .A(n42915), .B(n42916), .Z(n40832) );
  XOR U39858 ( .A(n40828), .B(n40829), .Z(n40831) );
  AND U39859 ( .A(n42917), .B(n42918), .Z(n40829) );
  XOR U39860 ( .A(n40825), .B(n40826), .Z(n40828) );
  AND U39861 ( .A(n42919), .B(n42920), .Z(n40826) );
  XOR U39862 ( .A(n40822), .B(n40823), .Z(n40825) );
  AND U39863 ( .A(n42921), .B(n42922), .Z(n40823) );
  XOR U39864 ( .A(n40819), .B(n40820), .Z(n40822) );
  AND U39865 ( .A(n42923), .B(n42924), .Z(n40820) );
  XOR U39866 ( .A(n40816), .B(n40817), .Z(n40819) );
  AND U39867 ( .A(n42925), .B(n42926), .Z(n40817) );
  XOR U39868 ( .A(n40813), .B(n40814), .Z(n40816) );
  AND U39869 ( .A(n42927), .B(n42928), .Z(n40814) );
  XOR U39870 ( .A(n40810), .B(n40811), .Z(n40813) );
  AND U39871 ( .A(n42929), .B(n42930), .Z(n40811) );
  XOR U39872 ( .A(n40807), .B(n40808), .Z(n40810) );
  AND U39873 ( .A(n42931), .B(n42932), .Z(n40808) );
  XOR U39874 ( .A(n40804), .B(n40805), .Z(n40807) );
  AND U39875 ( .A(n42933), .B(n42934), .Z(n40805) );
  XOR U39876 ( .A(n40801), .B(n40802), .Z(n40804) );
  AND U39877 ( .A(n42935), .B(n42936), .Z(n40802) );
  XOR U39878 ( .A(n40798), .B(n40799), .Z(n40801) );
  AND U39879 ( .A(n42937), .B(n42938), .Z(n40799) );
  XOR U39880 ( .A(n40795), .B(n40796), .Z(n40798) );
  AND U39881 ( .A(n42939), .B(n42940), .Z(n40796) );
  XOR U39882 ( .A(n40792), .B(n40793), .Z(n40795) );
  AND U39883 ( .A(n42941), .B(n42942), .Z(n40793) );
  XOR U39884 ( .A(n40789), .B(n40790), .Z(n40792) );
  AND U39885 ( .A(n42943), .B(n42944), .Z(n40790) );
  XOR U39886 ( .A(n40786), .B(n40787), .Z(n40789) );
  AND U39887 ( .A(n42945), .B(n42946), .Z(n40787) );
  XOR U39888 ( .A(n40783), .B(n40784), .Z(n40786) );
  AND U39889 ( .A(n42947), .B(n42948), .Z(n40784) );
  XOR U39890 ( .A(n40780), .B(n40781), .Z(n40783) );
  AND U39891 ( .A(n42949), .B(n42950), .Z(n40781) );
  XOR U39892 ( .A(n40777), .B(n40778), .Z(n40780) );
  AND U39893 ( .A(n42951), .B(n42952), .Z(n40778) );
  XOR U39894 ( .A(n40774), .B(n40775), .Z(n40777) );
  AND U39895 ( .A(n42953), .B(n42954), .Z(n40775) );
  XOR U39896 ( .A(n40771), .B(n40772), .Z(n40774) );
  AND U39897 ( .A(n42955), .B(n42956), .Z(n40772) );
  XOR U39898 ( .A(n40768), .B(n40769), .Z(n40771) );
  AND U39899 ( .A(n42957), .B(n42958), .Z(n40769) );
  XOR U39900 ( .A(n40765), .B(n40766), .Z(n40768) );
  AND U39901 ( .A(n42959), .B(n42960), .Z(n40766) );
  XOR U39902 ( .A(n40762), .B(n40763), .Z(n40765) );
  AND U39903 ( .A(n42961), .B(n42962), .Z(n40763) );
  XOR U39904 ( .A(n40759), .B(n40760), .Z(n40762) );
  AND U39905 ( .A(n42963), .B(n42964), .Z(n40760) );
  XOR U39906 ( .A(n40756), .B(n40757), .Z(n40759) );
  AND U39907 ( .A(n42965), .B(n42966), .Z(n40757) );
  XOR U39908 ( .A(n40753), .B(n40754), .Z(n40756) );
  AND U39909 ( .A(n42967), .B(n42968), .Z(n40754) );
  XOR U39910 ( .A(n40750), .B(n40751), .Z(n40753) );
  AND U39911 ( .A(n42969), .B(n42970), .Z(n40751) );
  XOR U39912 ( .A(n40747), .B(n40748), .Z(n40750) );
  AND U39913 ( .A(n42971), .B(n42972), .Z(n40748) );
  XOR U39914 ( .A(n40744), .B(n40745), .Z(n40747) );
  AND U39915 ( .A(n42973), .B(n42974), .Z(n40745) );
  XOR U39916 ( .A(n40741), .B(n40742), .Z(n40744) );
  AND U39917 ( .A(n42975), .B(n42976), .Z(n40742) );
  XOR U39918 ( .A(n40738), .B(n40739), .Z(n40741) );
  AND U39919 ( .A(n42977), .B(n42978), .Z(n40739) );
  XOR U39920 ( .A(n40735), .B(n40736), .Z(n40738) );
  AND U39921 ( .A(n42979), .B(n42980), .Z(n40736) );
  XOR U39922 ( .A(n40732), .B(n40733), .Z(n40735) );
  AND U39923 ( .A(n42981), .B(n42982), .Z(n40733) );
  XOR U39924 ( .A(n40729), .B(n40730), .Z(n40732) );
  AND U39925 ( .A(n42983), .B(n42984), .Z(n40730) );
  XOR U39926 ( .A(n40726), .B(n40727), .Z(n40729) );
  AND U39927 ( .A(n42985), .B(n42986), .Z(n40727) );
  XOR U39928 ( .A(n40723), .B(n40724), .Z(n40726) );
  AND U39929 ( .A(n42987), .B(n42988), .Z(n40724) );
  XOR U39930 ( .A(n40720), .B(n40721), .Z(n40723) );
  AND U39931 ( .A(n42989), .B(n42990), .Z(n40721) );
  XOR U39932 ( .A(n40717), .B(n40718), .Z(n40720) );
  AND U39933 ( .A(n42991), .B(n42992), .Z(n40718) );
  XOR U39934 ( .A(n40714), .B(n40715), .Z(n40717) );
  AND U39935 ( .A(n42993), .B(n42994), .Z(n40715) );
  XOR U39936 ( .A(n40711), .B(n40712), .Z(n40714) );
  AND U39937 ( .A(n42995), .B(n42996), .Z(n40712) );
  XOR U39938 ( .A(n40708), .B(n40709), .Z(n40711) );
  AND U39939 ( .A(n42997), .B(n42998), .Z(n40709) );
  XOR U39940 ( .A(n40705), .B(n40706), .Z(n40708) );
  AND U39941 ( .A(n42999), .B(n43000), .Z(n40706) );
  XOR U39942 ( .A(n40702), .B(n40703), .Z(n40705) );
  AND U39943 ( .A(n43001), .B(n43002), .Z(n40703) );
  XOR U39944 ( .A(n40699), .B(n40700), .Z(n40702) );
  AND U39945 ( .A(n43003), .B(n43004), .Z(n40700) );
  XOR U39946 ( .A(n40696), .B(n40697), .Z(n40699) );
  AND U39947 ( .A(n43005), .B(n43006), .Z(n40697) );
  XOR U39948 ( .A(n40693), .B(n40694), .Z(n40696) );
  AND U39949 ( .A(n43007), .B(n43008), .Z(n40694) );
  XOR U39950 ( .A(n40690), .B(n40691), .Z(n40693) );
  AND U39951 ( .A(n43009), .B(n43010), .Z(n40691) );
  XOR U39952 ( .A(n40687), .B(n40688), .Z(n40690) );
  AND U39953 ( .A(n43011), .B(n43012), .Z(n40688) );
  XOR U39954 ( .A(n40684), .B(n40685), .Z(n40687) );
  AND U39955 ( .A(n43013), .B(n43014), .Z(n40685) );
  XOR U39956 ( .A(n40681), .B(n40682), .Z(n40684) );
  AND U39957 ( .A(n43015), .B(n43016), .Z(n40682) );
  XOR U39958 ( .A(n40678), .B(n40679), .Z(n40681) );
  AND U39959 ( .A(n43017), .B(n43018), .Z(n40679) );
  XOR U39960 ( .A(n40675), .B(n40676), .Z(n40678) );
  AND U39961 ( .A(n43019), .B(n43020), .Z(n40676) );
  XOR U39962 ( .A(n40672), .B(n40673), .Z(n40675) );
  AND U39963 ( .A(n43021), .B(n43022), .Z(n40673) );
  XOR U39964 ( .A(n40669), .B(n40670), .Z(n40672) );
  AND U39965 ( .A(n43023), .B(n43024), .Z(n40670) );
  XOR U39966 ( .A(n40666), .B(n40667), .Z(n40669) );
  AND U39967 ( .A(n43025), .B(n43026), .Z(n40667) );
  XOR U39968 ( .A(n40663), .B(n40664), .Z(n40666) );
  AND U39969 ( .A(n43027), .B(n43028), .Z(n40664) );
  XOR U39970 ( .A(n40660), .B(n40661), .Z(n40663) );
  AND U39971 ( .A(n43029), .B(n43030), .Z(n40661) );
  XOR U39972 ( .A(n40657), .B(n40658), .Z(n40660) );
  AND U39973 ( .A(n43031), .B(n43032), .Z(n40658) );
  XOR U39974 ( .A(n40654), .B(n40655), .Z(n40657) );
  AND U39975 ( .A(n43033), .B(n43034), .Z(n40655) );
  XOR U39976 ( .A(n40651), .B(n40652), .Z(n40654) );
  AND U39977 ( .A(n43035), .B(n43036), .Z(n40652) );
  XOR U39978 ( .A(n40648), .B(n40649), .Z(n40651) );
  AND U39979 ( .A(n43037), .B(n43038), .Z(n40649) );
  XOR U39980 ( .A(n40645), .B(n40646), .Z(n40648) );
  AND U39981 ( .A(n43039), .B(n43040), .Z(n40646) );
  XOR U39982 ( .A(n40642), .B(n40643), .Z(n40645) );
  AND U39983 ( .A(n43041), .B(n43042), .Z(n40643) );
  XOR U39984 ( .A(n40639), .B(n40640), .Z(n40642) );
  AND U39985 ( .A(n43043), .B(n43044), .Z(n40640) );
  XOR U39986 ( .A(n40636), .B(n40637), .Z(n40639) );
  AND U39987 ( .A(n43045), .B(n43046), .Z(n40637) );
  XOR U39988 ( .A(n40633), .B(n40634), .Z(n40636) );
  AND U39989 ( .A(n43047), .B(n43048), .Z(n40634) );
  XOR U39990 ( .A(n40630), .B(n40631), .Z(n40633) );
  AND U39991 ( .A(n43049), .B(n43050), .Z(n40631) );
  XOR U39992 ( .A(n40627), .B(n40628), .Z(n40630) );
  AND U39993 ( .A(n43051), .B(n43052), .Z(n40628) );
  XOR U39994 ( .A(n40624), .B(n40625), .Z(n40627) );
  AND U39995 ( .A(n43053), .B(n43054), .Z(n40625) );
  XOR U39996 ( .A(n40621), .B(n40622), .Z(n40624) );
  AND U39997 ( .A(n43055), .B(n43056), .Z(n40622) );
  XOR U39998 ( .A(n40618), .B(n40619), .Z(n40621) );
  AND U39999 ( .A(n43057), .B(n43058), .Z(n40619) );
  XOR U40000 ( .A(n40615), .B(n40616), .Z(n40618) );
  AND U40001 ( .A(n43059), .B(n43060), .Z(n40616) );
  XOR U40002 ( .A(n40612), .B(n40613), .Z(n40615) );
  AND U40003 ( .A(n43061), .B(n43062), .Z(n40613) );
  XOR U40004 ( .A(n40609), .B(n40610), .Z(n40612) );
  AND U40005 ( .A(n43063), .B(n43064), .Z(n40610) );
  XOR U40006 ( .A(n40606), .B(n40607), .Z(n40609) );
  AND U40007 ( .A(n43065), .B(n43066), .Z(n40607) );
  XOR U40008 ( .A(n40603), .B(n40604), .Z(n40606) );
  AND U40009 ( .A(n43067), .B(n43068), .Z(n40604) );
  XOR U40010 ( .A(n40600), .B(n40601), .Z(n40603) );
  AND U40011 ( .A(n43069), .B(n43070), .Z(n40601) );
  XOR U40012 ( .A(n40597), .B(n40598), .Z(n40600) );
  AND U40013 ( .A(n43071), .B(n43072), .Z(n40598) );
  XOR U40014 ( .A(n40594), .B(n40595), .Z(n40597) );
  AND U40015 ( .A(n43073), .B(n43074), .Z(n40595) );
  XOR U40016 ( .A(n40591), .B(n40592), .Z(n40594) );
  AND U40017 ( .A(n43075), .B(n43076), .Z(n40592) );
  XOR U40018 ( .A(n40588), .B(n40589), .Z(n40591) );
  AND U40019 ( .A(n43077), .B(n43078), .Z(n40589) );
  XOR U40020 ( .A(n40585), .B(n40586), .Z(n40588) );
  AND U40021 ( .A(n43079), .B(n43080), .Z(n40586) );
  XOR U40022 ( .A(n40582), .B(n40583), .Z(n40585) );
  AND U40023 ( .A(n43081), .B(n43082), .Z(n40583) );
  XOR U40024 ( .A(n40579), .B(n40580), .Z(n40582) );
  AND U40025 ( .A(n43083), .B(n43084), .Z(n40580) );
  XOR U40026 ( .A(n40576), .B(n40577), .Z(n40579) );
  AND U40027 ( .A(n43085), .B(n43086), .Z(n40577) );
  XOR U40028 ( .A(n40573), .B(n40574), .Z(n40576) );
  AND U40029 ( .A(n43087), .B(n43088), .Z(n40574) );
  XOR U40030 ( .A(n40570), .B(n40571), .Z(n40573) );
  AND U40031 ( .A(n43089), .B(n43090), .Z(n40571) );
  XOR U40032 ( .A(n40567), .B(n40568), .Z(n40570) );
  AND U40033 ( .A(n43091), .B(n43092), .Z(n40568) );
  XOR U40034 ( .A(n40564), .B(n40565), .Z(n40567) );
  AND U40035 ( .A(n43093), .B(n43094), .Z(n40565) );
  XOR U40036 ( .A(n40561), .B(n40562), .Z(n40564) );
  AND U40037 ( .A(n43095), .B(n43096), .Z(n40562) );
  XOR U40038 ( .A(n40558), .B(n40559), .Z(n40561) );
  AND U40039 ( .A(n43097), .B(n43098), .Z(n40559) );
  XOR U40040 ( .A(n40555), .B(n40556), .Z(n40558) );
  AND U40041 ( .A(n43099), .B(n43100), .Z(n40556) );
  XOR U40042 ( .A(n40552), .B(n40553), .Z(n40555) );
  AND U40043 ( .A(n43101), .B(n43102), .Z(n40553) );
  XOR U40044 ( .A(n40549), .B(n40550), .Z(n40552) );
  AND U40045 ( .A(n43103), .B(n43104), .Z(n40550) );
  XOR U40046 ( .A(n40546), .B(n40547), .Z(n40549) );
  AND U40047 ( .A(n43105), .B(n43106), .Z(n40547) );
  XOR U40048 ( .A(n40543), .B(n40544), .Z(n40546) );
  AND U40049 ( .A(n43107), .B(n43108), .Z(n40544) );
  XOR U40050 ( .A(n40540), .B(n40541), .Z(n40543) );
  AND U40051 ( .A(n43109), .B(n43110), .Z(n40541) );
  XOR U40052 ( .A(n40537), .B(n40538), .Z(n40540) );
  AND U40053 ( .A(n43111), .B(n43112), .Z(n40538) );
  XOR U40054 ( .A(n40534), .B(n40535), .Z(n40537) );
  AND U40055 ( .A(n43113), .B(n43114), .Z(n40535) );
  XOR U40056 ( .A(n40531), .B(n40532), .Z(n40534) );
  AND U40057 ( .A(n43115), .B(n43116), .Z(n40532) );
  XOR U40058 ( .A(n40528), .B(n40529), .Z(n40531) );
  AND U40059 ( .A(n43117), .B(n43118), .Z(n40529) );
  XOR U40060 ( .A(n40525), .B(n40526), .Z(n40528) );
  AND U40061 ( .A(n43119), .B(n43120), .Z(n40526) );
  XOR U40062 ( .A(n40522), .B(n40523), .Z(n40525) );
  AND U40063 ( .A(n43121), .B(n43122), .Z(n40523) );
  XOR U40064 ( .A(n40519), .B(n40520), .Z(n40522) );
  AND U40065 ( .A(n43123), .B(n43124), .Z(n40520) );
  XOR U40066 ( .A(n40516), .B(n40517), .Z(n40519) );
  AND U40067 ( .A(n43125), .B(n43126), .Z(n40517) );
  XOR U40068 ( .A(n40513), .B(n40514), .Z(n40516) );
  AND U40069 ( .A(n43127), .B(n43128), .Z(n40514) );
  XOR U40070 ( .A(n40510), .B(n40511), .Z(n40513) );
  AND U40071 ( .A(n43129), .B(n43130), .Z(n40511) );
  XOR U40072 ( .A(n40507), .B(n40508), .Z(n40510) );
  AND U40073 ( .A(n43131), .B(n43132), .Z(n40508) );
  XOR U40074 ( .A(n40504), .B(n40505), .Z(n40507) );
  AND U40075 ( .A(n43133), .B(n43134), .Z(n40505) );
  XOR U40076 ( .A(n40501), .B(n40502), .Z(n40504) );
  AND U40077 ( .A(n43135), .B(n43136), .Z(n40502) );
  XOR U40078 ( .A(n40498), .B(n40499), .Z(n40501) );
  AND U40079 ( .A(n43137), .B(n43138), .Z(n40499) );
  XOR U40080 ( .A(n40495), .B(n40496), .Z(n40498) );
  AND U40081 ( .A(n43139), .B(n43140), .Z(n40496) );
  XOR U40082 ( .A(n40492), .B(n40493), .Z(n40495) );
  AND U40083 ( .A(n43141), .B(n43142), .Z(n40493) );
  XOR U40084 ( .A(n40489), .B(n40490), .Z(n40492) );
  AND U40085 ( .A(n43143), .B(n43144), .Z(n40490) );
  XOR U40086 ( .A(n40486), .B(n40487), .Z(n40489) );
  AND U40087 ( .A(n43145), .B(n43146), .Z(n40487) );
  XOR U40088 ( .A(n40483), .B(n40484), .Z(n40486) );
  AND U40089 ( .A(n43147), .B(n43148), .Z(n40484) );
  XOR U40090 ( .A(n40480), .B(n40481), .Z(n40483) );
  AND U40091 ( .A(n43149), .B(n43150), .Z(n40481) );
  XOR U40092 ( .A(n40477), .B(n40478), .Z(n40480) );
  AND U40093 ( .A(n43151), .B(n43152), .Z(n40478) );
  XOR U40094 ( .A(n40474), .B(n40475), .Z(n40477) );
  AND U40095 ( .A(n43153), .B(n43154), .Z(n40475) );
  XOR U40096 ( .A(n40471), .B(n40472), .Z(n40474) );
  AND U40097 ( .A(n43155), .B(n43156), .Z(n40472) );
  XOR U40098 ( .A(n40468), .B(n40469), .Z(n40471) );
  AND U40099 ( .A(n43157), .B(n43158), .Z(n40469) );
  XOR U40100 ( .A(n40465), .B(n40466), .Z(n40468) );
  AND U40101 ( .A(n43159), .B(n43160), .Z(n40466) );
  XOR U40102 ( .A(n40462), .B(n40463), .Z(n40465) );
  AND U40103 ( .A(n43161), .B(n43162), .Z(n40463) );
  XOR U40104 ( .A(n40459), .B(n40460), .Z(n40462) );
  AND U40105 ( .A(n43163), .B(n43164), .Z(n40460) );
  XOR U40106 ( .A(n40456), .B(n40457), .Z(n40459) );
  AND U40107 ( .A(n43165), .B(n43166), .Z(n40457) );
  XOR U40108 ( .A(n40453), .B(n40454), .Z(n40456) );
  AND U40109 ( .A(n43167), .B(n43168), .Z(n40454) );
  XOR U40110 ( .A(n40450), .B(n40451), .Z(n40453) );
  AND U40111 ( .A(n43169), .B(n43170), .Z(n40451) );
  XOR U40112 ( .A(n40447), .B(n40448), .Z(n40450) );
  AND U40113 ( .A(n43171), .B(n43172), .Z(n40448) );
  XOR U40114 ( .A(n40444), .B(n40445), .Z(n40447) );
  AND U40115 ( .A(n43173), .B(n43174), .Z(n40445) );
  XOR U40116 ( .A(n40441), .B(n40442), .Z(n40444) );
  AND U40117 ( .A(n43175), .B(n43176), .Z(n40442) );
  XOR U40118 ( .A(n40438), .B(n40439), .Z(n40441) );
  AND U40119 ( .A(n43177), .B(n43178), .Z(n40439) );
  XOR U40120 ( .A(n40435), .B(n40436), .Z(n40438) );
  AND U40121 ( .A(n43179), .B(n43180), .Z(n40436) );
  XOR U40122 ( .A(n40432), .B(n40433), .Z(n40435) );
  AND U40123 ( .A(n43181), .B(n43182), .Z(n40433) );
  XOR U40124 ( .A(n40429), .B(n40430), .Z(n40432) );
  AND U40125 ( .A(n43183), .B(n43184), .Z(n40430) );
  XOR U40126 ( .A(n40426), .B(n40427), .Z(n40429) );
  AND U40127 ( .A(n43185), .B(n43186), .Z(n40427) );
  XOR U40128 ( .A(n40423), .B(n40424), .Z(n40426) );
  AND U40129 ( .A(n43187), .B(n43188), .Z(n40424) );
  XOR U40130 ( .A(n40420), .B(n40421), .Z(n40423) );
  AND U40131 ( .A(n43189), .B(n43190), .Z(n40421) );
  XOR U40132 ( .A(n40417), .B(n40418), .Z(n40420) );
  AND U40133 ( .A(n43191), .B(n43192), .Z(n40418) );
  XOR U40134 ( .A(n40414), .B(n40415), .Z(n40417) );
  AND U40135 ( .A(n43193), .B(n43194), .Z(n40415) );
  XOR U40136 ( .A(n40411), .B(n40412), .Z(n40414) );
  AND U40137 ( .A(n43195), .B(n43196), .Z(n40412) );
  XOR U40138 ( .A(n40408), .B(n40409), .Z(n40411) );
  AND U40139 ( .A(n43197), .B(n43198), .Z(n40409) );
  XOR U40140 ( .A(n40405), .B(n40406), .Z(n40408) );
  AND U40141 ( .A(n43199), .B(n43200), .Z(n40406) );
  XOR U40142 ( .A(n40402), .B(n40403), .Z(n40405) );
  AND U40143 ( .A(n43201), .B(n43202), .Z(n40403) );
  XOR U40144 ( .A(n40399), .B(n40400), .Z(n40402) );
  AND U40145 ( .A(n43203), .B(n43204), .Z(n40400) );
  XOR U40146 ( .A(n40396), .B(n40397), .Z(n40399) );
  AND U40147 ( .A(n43205), .B(n43206), .Z(n40397) );
  XOR U40148 ( .A(n40393), .B(n40394), .Z(n40396) );
  AND U40149 ( .A(n43207), .B(n43208), .Z(n40394) );
  XOR U40150 ( .A(n40390), .B(n40391), .Z(n40393) );
  AND U40151 ( .A(n43209), .B(n43210), .Z(n40391) );
  XOR U40152 ( .A(n40387), .B(n40388), .Z(n40390) );
  AND U40153 ( .A(n43211), .B(n43212), .Z(n40388) );
  XOR U40154 ( .A(n40384), .B(n40385), .Z(n40387) );
  AND U40155 ( .A(n43213), .B(n43214), .Z(n40385) );
  XOR U40156 ( .A(n40381), .B(n40382), .Z(n40384) );
  AND U40157 ( .A(n43215), .B(n43216), .Z(n40382) );
  XOR U40158 ( .A(n40378), .B(n40379), .Z(n40381) );
  AND U40159 ( .A(n43217), .B(n43218), .Z(n40379) );
  XOR U40160 ( .A(n40375), .B(n40376), .Z(n40378) );
  AND U40161 ( .A(n43219), .B(n43220), .Z(n40376) );
  XOR U40162 ( .A(n40372), .B(n40373), .Z(n40375) );
  AND U40163 ( .A(n43221), .B(n43222), .Z(n40373) );
  XOR U40164 ( .A(n40369), .B(n40370), .Z(n40372) );
  AND U40165 ( .A(n43223), .B(n43224), .Z(n40370) );
  XOR U40166 ( .A(n40366), .B(n40367), .Z(n40369) );
  AND U40167 ( .A(n43225), .B(n43226), .Z(n40367) );
  XOR U40168 ( .A(n40363), .B(n40364), .Z(n40366) );
  AND U40169 ( .A(n43227), .B(n43228), .Z(n40364) );
  XOR U40170 ( .A(n40360), .B(n40361), .Z(n40363) );
  AND U40171 ( .A(n43229), .B(n43230), .Z(n40361) );
  XOR U40172 ( .A(n40357), .B(n40358), .Z(n40360) );
  AND U40173 ( .A(n43231), .B(n43232), .Z(n40358) );
  XOR U40174 ( .A(n40354), .B(n40355), .Z(n40357) );
  AND U40175 ( .A(n43233), .B(n43234), .Z(n40355) );
  XOR U40176 ( .A(n40351), .B(n40352), .Z(n40354) );
  AND U40177 ( .A(n43235), .B(n43236), .Z(n40352) );
  XOR U40178 ( .A(n40348), .B(n40349), .Z(n40351) );
  AND U40179 ( .A(n43237), .B(n43238), .Z(n40349) );
  XOR U40180 ( .A(n40345), .B(n40346), .Z(n40348) );
  AND U40181 ( .A(n43239), .B(n43240), .Z(n40346) );
  XOR U40182 ( .A(n40342), .B(n40343), .Z(n40345) );
  AND U40183 ( .A(n43241), .B(n43242), .Z(n40343) );
  XOR U40184 ( .A(n40339), .B(n40340), .Z(n40342) );
  AND U40185 ( .A(n43243), .B(n43244), .Z(n40340) );
  XOR U40186 ( .A(n40336), .B(n40337), .Z(n40339) );
  AND U40187 ( .A(n43245), .B(n43246), .Z(n40337) );
  XOR U40188 ( .A(n40333), .B(n40334), .Z(n40336) );
  AND U40189 ( .A(n43247), .B(n43248), .Z(n40334) );
  XOR U40190 ( .A(n40330), .B(n40331), .Z(n40333) );
  AND U40191 ( .A(n43249), .B(n43250), .Z(n40331) );
  XOR U40192 ( .A(n40327), .B(n40328), .Z(n40330) );
  AND U40193 ( .A(n43251), .B(n43252), .Z(n40328) );
  XOR U40194 ( .A(n40324), .B(n40325), .Z(n40327) );
  AND U40195 ( .A(n43253), .B(n43254), .Z(n40325) );
  XOR U40196 ( .A(n40321), .B(n40322), .Z(n40324) );
  AND U40197 ( .A(n43255), .B(n43256), .Z(n40322) );
  XOR U40198 ( .A(n40318), .B(n40319), .Z(n40321) );
  AND U40199 ( .A(n43257), .B(n43258), .Z(n40319) );
  XOR U40200 ( .A(n40315), .B(n40316), .Z(n40318) );
  AND U40201 ( .A(n43259), .B(n43260), .Z(n40316) );
  XOR U40202 ( .A(n40312), .B(n40313), .Z(n40315) );
  AND U40203 ( .A(n43261), .B(n43262), .Z(n40313) );
  XOR U40204 ( .A(n40309), .B(n40310), .Z(n40312) );
  AND U40205 ( .A(n43263), .B(n43264), .Z(n40310) );
  XOR U40206 ( .A(n40306), .B(n40307), .Z(n40309) );
  AND U40207 ( .A(n43265), .B(n43266), .Z(n40307) );
  XOR U40208 ( .A(n40303), .B(n40304), .Z(n40306) );
  AND U40209 ( .A(n43267), .B(n43268), .Z(n40304) );
  XOR U40210 ( .A(n40300), .B(n40301), .Z(n40303) );
  AND U40211 ( .A(n43269), .B(n43270), .Z(n40301) );
  XOR U40212 ( .A(n40297), .B(n40298), .Z(n40300) );
  AND U40213 ( .A(n43271), .B(n43272), .Z(n40298) );
  XOR U40214 ( .A(n40294), .B(n40295), .Z(n40297) );
  AND U40215 ( .A(n43273), .B(n43274), .Z(n40295) );
  XOR U40216 ( .A(n40291), .B(n40292), .Z(n40294) );
  AND U40217 ( .A(n43275), .B(n43276), .Z(n40292) );
  XOR U40218 ( .A(n40288), .B(n40289), .Z(n40291) );
  AND U40219 ( .A(n43277), .B(n43278), .Z(n40289) );
  XOR U40220 ( .A(n40285), .B(n40286), .Z(n40288) );
  AND U40221 ( .A(n43279), .B(n43280), .Z(n40286) );
  XOR U40222 ( .A(n40282), .B(n40283), .Z(n40285) );
  AND U40223 ( .A(n43281), .B(n43282), .Z(n40283) );
  XOR U40224 ( .A(n40279), .B(n40280), .Z(n40282) );
  AND U40225 ( .A(n43283), .B(n43284), .Z(n40280) );
  XOR U40226 ( .A(n40276), .B(n40277), .Z(n40279) );
  AND U40227 ( .A(n43285), .B(n43286), .Z(n40277) );
  XOR U40228 ( .A(n40273), .B(n40274), .Z(n40276) );
  AND U40229 ( .A(n43287), .B(n43288), .Z(n40274) );
  XOR U40230 ( .A(n40270), .B(n40271), .Z(n40273) );
  AND U40231 ( .A(n43289), .B(n43290), .Z(n40271) );
  XOR U40232 ( .A(n40267), .B(n40268), .Z(n40270) );
  AND U40233 ( .A(n43291), .B(n43292), .Z(n40268) );
  XOR U40234 ( .A(n40264), .B(n40265), .Z(n40267) );
  AND U40235 ( .A(n43293), .B(n43294), .Z(n40265) );
  XOR U40236 ( .A(n40261), .B(n40262), .Z(n40264) );
  AND U40237 ( .A(n43295), .B(n43296), .Z(n40262) );
  XOR U40238 ( .A(n40258), .B(n40259), .Z(n40261) );
  AND U40239 ( .A(n43297), .B(n43298), .Z(n40259) );
  XOR U40240 ( .A(n40255), .B(n40256), .Z(n40258) );
  AND U40241 ( .A(n43299), .B(n43300), .Z(n40256) );
  XOR U40242 ( .A(n40252), .B(n40253), .Z(n40255) );
  AND U40243 ( .A(n43301), .B(n43302), .Z(n40253) );
  XOR U40244 ( .A(n40249), .B(n40250), .Z(n40252) );
  AND U40245 ( .A(n43303), .B(n43304), .Z(n40250) );
  XOR U40246 ( .A(n40246), .B(n40247), .Z(n40249) );
  AND U40247 ( .A(n43305), .B(n43306), .Z(n40247) );
  XOR U40248 ( .A(n40243), .B(n40244), .Z(n40246) );
  AND U40249 ( .A(n43307), .B(n43308), .Z(n40244) );
  XOR U40250 ( .A(n40240), .B(n40241), .Z(n40243) );
  AND U40251 ( .A(n43309), .B(n43310), .Z(n40241) );
  XOR U40252 ( .A(n40237), .B(n40238), .Z(n40240) );
  AND U40253 ( .A(n43311), .B(n43312), .Z(n40238) );
  XOR U40254 ( .A(n40234), .B(n40235), .Z(n40237) );
  AND U40255 ( .A(n43313), .B(n43314), .Z(n40235) );
  XOR U40256 ( .A(n40231), .B(n40232), .Z(n40234) );
  AND U40257 ( .A(n43315), .B(n43316), .Z(n40232) );
  XOR U40258 ( .A(n40228), .B(n40229), .Z(n40231) );
  AND U40259 ( .A(n43317), .B(n43318), .Z(n40229) );
  XOR U40260 ( .A(n40225), .B(n40226), .Z(n40228) );
  AND U40261 ( .A(n43319), .B(n43320), .Z(n40226) );
  XOR U40262 ( .A(n40222), .B(n40223), .Z(n40225) );
  AND U40263 ( .A(n43321), .B(n43322), .Z(n40223) );
  XOR U40264 ( .A(n40219), .B(n40220), .Z(n40222) );
  AND U40265 ( .A(n43323), .B(n43324), .Z(n40220) );
  XOR U40266 ( .A(n40216), .B(n40217), .Z(n40219) );
  AND U40267 ( .A(n43325), .B(n43326), .Z(n40217) );
  XOR U40268 ( .A(n40213), .B(n40214), .Z(n40216) );
  AND U40269 ( .A(n43327), .B(n43328), .Z(n40214) );
  XOR U40270 ( .A(n40210), .B(n40211), .Z(n40213) );
  AND U40271 ( .A(n43329), .B(n43330), .Z(n40211) );
  XOR U40272 ( .A(n40207), .B(n40208), .Z(n40210) );
  AND U40273 ( .A(n43331), .B(n43332), .Z(n40208) );
  XOR U40274 ( .A(n40204), .B(n40205), .Z(n40207) );
  AND U40275 ( .A(n43333), .B(n43334), .Z(n40205) );
  XOR U40276 ( .A(n40201), .B(n40202), .Z(n40204) );
  AND U40277 ( .A(n43335), .B(n43336), .Z(n40202) );
  XOR U40278 ( .A(n40198), .B(n40199), .Z(n40201) );
  AND U40279 ( .A(n43337), .B(n43338), .Z(n40199) );
  XOR U40280 ( .A(n40195), .B(n40196), .Z(n40198) );
  AND U40281 ( .A(n43339), .B(n43340), .Z(n40196) );
  XOR U40282 ( .A(n40192), .B(n40193), .Z(n40195) );
  AND U40283 ( .A(n43341), .B(n43342), .Z(n40193) );
  XOR U40284 ( .A(n40189), .B(n40190), .Z(n40192) );
  AND U40285 ( .A(n43343), .B(n43344), .Z(n40190) );
  XOR U40286 ( .A(n40186), .B(n40187), .Z(n40189) );
  AND U40287 ( .A(n43345), .B(n43346), .Z(n40187) );
  XOR U40288 ( .A(n40183), .B(n40184), .Z(n40186) );
  AND U40289 ( .A(n43347), .B(n43348), .Z(n40184) );
  XOR U40290 ( .A(n40180), .B(n40181), .Z(n40183) );
  AND U40291 ( .A(n43349), .B(n43350), .Z(n40181) );
  XOR U40292 ( .A(n40177), .B(n40178), .Z(n40180) );
  AND U40293 ( .A(n43351), .B(n43352), .Z(n40178) );
  XOR U40294 ( .A(n40174), .B(n40175), .Z(n40177) );
  AND U40295 ( .A(n43353), .B(n43354), .Z(n40175) );
  XOR U40296 ( .A(n40171), .B(n40172), .Z(n40174) );
  AND U40297 ( .A(n43355), .B(n43356), .Z(n40172) );
  XOR U40298 ( .A(n40168), .B(n40169), .Z(n40171) );
  AND U40299 ( .A(n43357), .B(n43358), .Z(n40169) );
  XOR U40300 ( .A(n40165), .B(n40166), .Z(n40168) );
  AND U40301 ( .A(n43359), .B(n43360), .Z(n40166) );
  XOR U40302 ( .A(n40162), .B(n40163), .Z(n40165) );
  AND U40303 ( .A(n43361), .B(n43362), .Z(n40163) );
  XOR U40304 ( .A(n40159), .B(n40160), .Z(n40162) );
  AND U40305 ( .A(n43363), .B(n43364), .Z(n40160) );
  XOR U40306 ( .A(n40156), .B(n40157), .Z(n40159) );
  AND U40307 ( .A(n43365), .B(n43366), .Z(n40157) );
  XOR U40308 ( .A(n40153), .B(n40154), .Z(n40156) );
  AND U40309 ( .A(n43367), .B(n43368), .Z(n40154) );
  XOR U40310 ( .A(n40150), .B(n40151), .Z(n40153) );
  AND U40311 ( .A(n43369), .B(n43370), .Z(n40151) );
  XOR U40312 ( .A(n40147), .B(n40148), .Z(n40150) );
  AND U40313 ( .A(n43371), .B(n43372), .Z(n40148) );
  XOR U40314 ( .A(n40144), .B(n40145), .Z(n40147) );
  AND U40315 ( .A(n43373), .B(n43374), .Z(n40145) );
  XOR U40316 ( .A(n40141), .B(n40142), .Z(n40144) );
  AND U40317 ( .A(n43375), .B(n43376), .Z(n40142) );
  XOR U40318 ( .A(n40138), .B(n40139), .Z(n40141) );
  AND U40319 ( .A(n43377), .B(n43378), .Z(n40139) );
  XOR U40320 ( .A(n40135), .B(n40136), .Z(n40138) );
  AND U40321 ( .A(n43379), .B(n43380), .Z(n40136) );
  XOR U40322 ( .A(n40132), .B(n40133), .Z(n40135) );
  AND U40323 ( .A(n43381), .B(n43382), .Z(n40133) );
  XOR U40324 ( .A(n40129), .B(n40130), .Z(n40132) );
  AND U40325 ( .A(n43383), .B(n43384), .Z(n40130) );
  XOR U40326 ( .A(n40126), .B(n40127), .Z(n40129) );
  AND U40327 ( .A(n43385), .B(n43386), .Z(n40127) );
  XOR U40328 ( .A(n40123), .B(n40124), .Z(n40126) );
  AND U40329 ( .A(n43387), .B(n43388), .Z(n40124) );
  XOR U40330 ( .A(n40120), .B(n40121), .Z(n40123) );
  AND U40331 ( .A(n43389), .B(n43390), .Z(n40121) );
  XOR U40332 ( .A(n40117), .B(n40118), .Z(n40120) );
  AND U40333 ( .A(n43391), .B(n43392), .Z(n40118) );
  XOR U40334 ( .A(n40114), .B(n40115), .Z(n40117) );
  AND U40335 ( .A(n43393), .B(n43394), .Z(n40115) );
  XOR U40336 ( .A(n40111), .B(n40112), .Z(n40114) );
  AND U40337 ( .A(n43395), .B(n43396), .Z(n40112) );
  XOR U40338 ( .A(n40108), .B(n40109), .Z(n40111) );
  AND U40339 ( .A(n43397), .B(n43398), .Z(n40109) );
  XOR U40340 ( .A(n40105), .B(n40106), .Z(n40108) );
  AND U40341 ( .A(n43399), .B(n43400), .Z(n40106) );
  XOR U40342 ( .A(n40102), .B(n40103), .Z(n40105) );
  AND U40343 ( .A(n43401), .B(n43402), .Z(n40103) );
  XOR U40344 ( .A(n40099), .B(n40100), .Z(n40102) );
  AND U40345 ( .A(n43403), .B(n43404), .Z(n40100) );
  XOR U40346 ( .A(n40096), .B(n40097), .Z(n40099) );
  AND U40347 ( .A(n43405), .B(n43406), .Z(n40097) );
  XOR U40348 ( .A(n40093), .B(n40094), .Z(n40096) );
  AND U40349 ( .A(n43407), .B(n43408), .Z(n40094) );
  XOR U40350 ( .A(n40090), .B(n40091), .Z(n40093) );
  AND U40351 ( .A(n43409), .B(n43410), .Z(n40091) );
  XOR U40352 ( .A(n40087), .B(n40088), .Z(n40090) );
  AND U40353 ( .A(n43411), .B(n43412), .Z(n40088) );
  XOR U40354 ( .A(n40084), .B(n40085), .Z(n40087) );
  AND U40355 ( .A(n43413), .B(n43414), .Z(n40085) );
  XOR U40356 ( .A(n40081), .B(n40082), .Z(n40084) );
  AND U40357 ( .A(n43415), .B(n43416), .Z(n40082) );
  XOR U40358 ( .A(n40078), .B(n40079), .Z(n40081) );
  AND U40359 ( .A(n43417), .B(n43418), .Z(n40079) );
  XNOR U40360 ( .A(n40075), .B(n40076), .Z(n40078) );
  AND U40361 ( .A(n43419), .B(n43420), .Z(n40076) );
  XOR U40362 ( .A(n43421), .B(n40073), .Z(n40075) );
  IV U40363 ( .A(n43422), .Z(n40073) );
  AND U40364 ( .A(n43423), .B(n43424), .Z(n43422) );
  IV U40365 ( .A(n40072), .Z(n43421) );
  XOR U40366 ( .A(n39813), .B(n40069), .Z(n40072) );
  AND U40367 ( .A(n43425), .B(n43426), .Z(n40069) );
  XOR U40368 ( .A(n39815), .B(n39814), .Z(n39813) );
  AND U40369 ( .A(n43427), .B(n43428), .Z(n39814) );
  XOR U40370 ( .A(n39817), .B(n39816), .Z(n39815) );
  AND U40371 ( .A(n43429), .B(n43430), .Z(n39816) );
  XOR U40372 ( .A(n39819), .B(n39818), .Z(n39817) );
  AND U40373 ( .A(n43431), .B(n43432), .Z(n39818) );
  XOR U40374 ( .A(n39821), .B(n39820), .Z(n39819) );
  AND U40375 ( .A(n43433), .B(n43434), .Z(n39820) );
  XOR U40376 ( .A(n39823), .B(n39822), .Z(n39821) );
  AND U40377 ( .A(n43435), .B(n43436), .Z(n39822) );
  XOR U40378 ( .A(n39825), .B(n39824), .Z(n39823) );
  AND U40379 ( .A(n43437), .B(n43438), .Z(n39824) );
  XOR U40380 ( .A(n39827), .B(n39826), .Z(n39825) );
  AND U40381 ( .A(n43439), .B(n43440), .Z(n39826) );
  XOR U40382 ( .A(n39829), .B(n39828), .Z(n39827) );
  AND U40383 ( .A(n43441), .B(n43442), .Z(n39828) );
  XOR U40384 ( .A(n39831), .B(n39830), .Z(n39829) );
  AND U40385 ( .A(n43443), .B(n43444), .Z(n39830) );
  XOR U40386 ( .A(n39833), .B(n39832), .Z(n39831) );
  AND U40387 ( .A(n43445), .B(n43446), .Z(n39832) );
  XOR U40388 ( .A(n39835), .B(n39834), .Z(n39833) );
  AND U40389 ( .A(n43447), .B(n43448), .Z(n39834) );
  XOR U40390 ( .A(n39837), .B(n39836), .Z(n39835) );
  AND U40391 ( .A(n43449), .B(n43450), .Z(n39836) );
  XOR U40392 ( .A(n39839), .B(n39838), .Z(n39837) );
  AND U40393 ( .A(n43451), .B(n43452), .Z(n39838) );
  XOR U40394 ( .A(n39841), .B(n39840), .Z(n39839) );
  AND U40395 ( .A(n43453), .B(n43454), .Z(n39840) );
  XOR U40396 ( .A(n39843), .B(n39842), .Z(n39841) );
  AND U40397 ( .A(n43455), .B(n43456), .Z(n39842) );
  XOR U40398 ( .A(n39845), .B(n39844), .Z(n39843) );
  AND U40399 ( .A(n43457), .B(n43458), .Z(n39844) );
  XOR U40400 ( .A(n39847), .B(n39846), .Z(n39845) );
  AND U40401 ( .A(n43459), .B(n43460), .Z(n39846) );
  XOR U40402 ( .A(n39849), .B(n39848), .Z(n39847) );
  AND U40403 ( .A(n43461), .B(n43462), .Z(n39848) );
  XOR U40404 ( .A(n39851), .B(n39850), .Z(n39849) );
  AND U40405 ( .A(n43463), .B(n43464), .Z(n39850) );
  XOR U40406 ( .A(n39853), .B(n39852), .Z(n39851) );
  AND U40407 ( .A(n43465), .B(n43466), .Z(n39852) );
  XOR U40408 ( .A(n39855), .B(n39854), .Z(n39853) );
  AND U40409 ( .A(n43467), .B(n43468), .Z(n39854) );
  XOR U40410 ( .A(n39857), .B(n39856), .Z(n39855) );
  AND U40411 ( .A(n43469), .B(n43470), .Z(n39856) );
  XOR U40412 ( .A(n39859), .B(n39858), .Z(n39857) );
  AND U40413 ( .A(n43471), .B(n43472), .Z(n39858) );
  XOR U40414 ( .A(n39861), .B(n39860), .Z(n39859) );
  AND U40415 ( .A(n43473), .B(n43474), .Z(n39860) );
  XOR U40416 ( .A(n39863), .B(n39862), .Z(n39861) );
  AND U40417 ( .A(n43475), .B(n43476), .Z(n39862) );
  XOR U40418 ( .A(n39865), .B(n39864), .Z(n39863) );
  AND U40419 ( .A(n43477), .B(n43478), .Z(n39864) );
  XOR U40420 ( .A(n39867), .B(n39866), .Z(n39865) );
  AND U40421 ( .A(n43479), .B(n43480), .Z(n39866) );
  XOR U40422 ( .A(n39869), .B(n39868), .Z(n39867) );
  AND U40423 ( .A(n43481), .B(n43482), .Z(n39868) );
  XOR U40424 ( .A(n39871), .B(n39870), .Z(n39869) );
  AND U40425 ( .A(n43483), .B(n43484), .Z(n39870) );
  XOR U40426 ( .A(n39873), .B(n39872), .Z(n39871) );
  AND U40427 ( .A(n43485), .B(n43486), .Z(n39872) );
  XOR U40428 ( .A(n39875), .B(n39874), .Z(n39873) );
  AND U40429 ( .A(n43487), .B(n43488), .Z(n39874) );
  XOR U40430 ( .A(n39877), .B(n39876), .Z(n39875) );
  AND U40431 ( .A(n43489), .B(n43490), .Z(n39876) );
  XOR U40432 ( .A(n39879), .B(n39878), .Z(n39877) );
  AND U40433 ( .A(n43491), .B(n43492), .Z(n39878) );
  XOR U40434 ( .A(n39881), .B(n39880), .Z(n39879) );
  AND U40435 ( .A(n43493), .B(n43494), .Z(n39880) );
  XOR U40436 ( .A(n39883), .B(n39882), .Z(n39881) );
  AND U40437 ( .A(n43495), .B(n43496), .Z(n39882) );
  XOR U40438 ( .A(n39885), .B(n39884), .Z(n39883) );
  AND U40439 ( .A(n43497), .B(n43498), .Z(n39884) );
  XOR U40440 ( .A(n39887), .B(n39886), .Z(n39885) );
  AND U40441 ( .A(n43499), .B(n43500), .Z(n39886) );
  XOR U40442 ( .A(n39889), .B(n39888), .Z(n39887) );
  AND U40443 ( .A(n43501), .B(n43502), .Z(n39888) );
  XOR U40444 ( .A(n39891), .B(n39890), .Z(n39889) );
  AND U40445 ( .A(n43503), .B(n43504), .Z(n39890) );
  XOR U40446 ( .A(n39893), .B(n39892), .Z(n39891) );
  AND U40447 ( .A(n43505), .B(n43506), .Z(n39892) );
  XOR U40448 ( .A(n39895), .B(n39894), .Z(n39893) );
  AND U40449 ( .A(n43507), .B(n43508), .Z(n39894) );
  XOR U40450 ( .A(n39897), .B(n39896), .Z(n39895) );
  AND U40451 ( .A(n43509), .B(n43510), .Z(n39896) );
  XOR U40452 ( .A(n39899), .B(n39898), .Z(n39897) );
  AND U40453 ( .A(n43511), .B(n43512), .Z(n39898) );
  XOR U40454 ( .A(n39901), .B(n39900), .Z(n39899) );
  AND U40455 ( .A(n43513), .B(n43514), .Z(n39900) );
  XOR U40456 ( .A(n39903), .B(n39902), .Z(n39901) );
  AND U40457 ( .A(n43515), .B(n43516), .Z(n39902) );
  XOR U40458 ( .A(n39905), .B(n39904), .Z(n39903) );
  AND U40459 ( .A(n43517), .B(n43518), .Z(n39904) );
  XOR U40460 ( .A(n39907), .B(n39906), .Z(n39905) );
  AND U40461 ( .A(n43519), .B(n43520), .Z(n39906) );
  XOR U40462 ( .A(n39909), .B(n39908), .Z(n39907) );
  AND U40463 ( .A(n43521), .B(n43522), .Z(n39908) );
  XOR U40464 ( .A(n39911), .B(n39910), .Z(n39909) );
  AND U40465 ( .A(n43523), .B(n43524), .Z(n39910) );
  XOR U40466 ( .A(n39913), .B(n39912), .Z(n39911) );
  AND U40467 ( .A(n43525), .B(n43526), .Z(n39912) );
  XOR U40468 ( .A(n39915), .B(n39914), .Z(n39913) );
  AND U40469 ( .A(n43527), .B(n43528), .Z(n39914) );
  XOR U40470 ( .A(n39917), .B(n39916), .Z(n39915) );
  AND U40471 ( .A(n43529), .B(n43530), .Z(n39916) );
  XOR U40472 ( .A(n39919), .B(n39918), .Z(n39917) );
  AND U40473 ( .A(n43531), .B(n43532), .Z(n39918) );
  XOR U40474 ( .A(n39921), .B(n39920), .Z(n39919) );
  AND U40475 ( .A(n43533), .B(n43534), .Z(n39920) );
  XOR U40476 ( .A(n39923), .B(n39922), .Z(n39921) );
  AND U40477 ( .A(n43535), .B(n43536), .Z(n39922) );
  XOR U40478 ( .A(n39925), .B(n39924), .Z(n39923) );
  AND U40479 ( .A(n43537), .B(n43538), .Z(n39924) );
  XOR U40480 ( .A(n39927), .B(n39926), .Z(n39925) );
  AND U40481 ( .A(n43539), .B(n43540), .Z(n39926) );
  XOR U40482 ( .A(n39929), .B(n39928), .Z(n39927) );
  AND U40483 ( .A(n43541), .B(n43542), .Z(n39928) );
  XOR U40484 ( .A(n39931), .B(n39930), .Z(n39929) );
  AND U40485 ( .A(n43543), .B(n43544), .Z(n39930) );
  XOR U40486 ( .A(n39933), .B(n39932), .Z(n39931) );
  AND U40487 ( .A(n43545), .B(n43546), .Z(n39932) );
  XOR U40488 ( .A(n39935), .B(n39934), .Z(n39933) );
  AND U40489 ( .A(n43547), .B(n43548), .Z(n39934) );
  XOR U40490 ( .A(n39937), .B(n39936), .Z(n39935) );
  AND U40491 ( .A(n43549), .B(n43550), .Z(n39936) );
  XOR U40492 ( .A(n39939), .B(n39938), .Z(n39937) );
  AND U40493 ( .A(n43551), .B(n43552), .Z(n39938) );
  XOR U40494 ( .A(n39941), .B(n39940), .Z(n39939) );
  AND U40495 ( .A(n43553), .B(n43554), .Z(n39940) );
  XOR U40496 ( .A(n39943), .B(n39942), .Z(n39941) );
  AND U40497 ( .A(n43555), .B(n43556), .Z(n39942) );
  XOR U40498 ( .A(n39945), .B(n39944), .Z(n39943) );
  AND U40499 ( .A(n43557), .B(n43558), .Z(n39944) );
  XOR U40500 ( .A(n39947), .B(n39946), .Z(n39945) );
  AND U40501 ( .A(n43559), .B(n43560), .Z(n39946) );
  XOR U40502 ( .A(n39949), .B(n39948), .Z(n39947) );
  AND U40503 ( .A(n43561), .B(n43562), .Z(n39948) );
  XOR U40504 ( .A(n39951), .B(n39950), .Z(n39949) );
  AND U40505 ( .A(n43563), .B(n43564), .Z(n39950) );
  XOR U40506 ( .A(n39953), .B(n39952), .Z(n39951) );
  AND U40507 ( .A(n43565), .B(n43566), .Z(n39952) );
  XOR U40508 ( .A(n39955), .B(n39954), .Z(n39953) );
  AND U40509 ( .A(n43567), .B(n43568), .Z(n39954) );
  XOR U40510 ( .A(n39957), .B(n39956), .Z(n39955) );
  AND U40511 ( .A(n43569), .B(n43570), .Z(n39956) );
  XOR U40512 ( .A(n39959), .B(n39958), .Z(n39957) );
  AND U40513 ( .A(n43571), .B(n43572), .Z(n39958) );
  XOR U40514 ( .A(n39961), .B(n39960), .Z(n39959) );
  AND U40515 ( .A(n43573), .B(n43574), .Z(n39960) );
  XOR U40516 ( .A(n39963), .B(n39962), .Z(n39961) );
  AND U40517 ( .A(n43575), .B(n43576), .Z(n39962) );
  XOR U40518 ( .A(n39965), .B(n39964), .Z(n39963) );
  AND U40519 ( .A(n43577), .B(n43578), .Z(n39964) );
  XOR U40520 ( .A(n39967), .B(n39966), .Z(n39965) );
  AND U40521 ( .A(n43579), .B(n43580), .Z(n39966) );
  XOR U40522 ( .A(n39969), .B(n39968), .Z(n39967) );
  AND U40523 ( .A(n43581), .B(n43582), .Z(n39968) );
  XOR U40524 ( .A(n39971), .B(n39970), .Z(n39969) );
  AND U40525 ( .A(n43583), .B(n43584), .Z(n39970) );
  XOR U40526 ( .A(n39973), .B(n39972), .Z(n39971) );
  AND U40527 ( .A(n43585), .B(n43586), .Z(n39972) );
  XOR U40528 ( .A(n39975), .B(n39974), .Z(n39973) );
  AND U40529 ( .A(n43587), .B(n43588), .Z(n39974) );
  XOR U40530 ( .A(n39977), .B(n39976), .Z(n39975) );
  AND U40531 ( .A(n43589), .B(n43590), .Z(n39976) );
  XOR U40532 ( .A(n39979), .B(n39978), .Z(n39977) );
  AND U40533 ( .A(n43591), .B(n43592), .Z(n39978) );
  XOR U40534 ( .A(n39981), .B(n39980), .Z(n39979) );
  AND U40535 ( .A(n43593), .B(n43594), .Z(n39980) );
  XOR U40536 ( .A(n39983), .B(n39982), .Z(n39981) );
  AND U40537 ( .A(n43595), .B(n43596), .Z(n39982) );
  XOR U40538 ( .A(n39985), .B(n39984), .Z(n39983) );
  AND U40539 ( .A(n43597), .B(n43598), .Z(n39984) );
  XOR U40540 ( .A(n39987), .B(n39986), .Z(n39985) );
  AND U40541 ( .A(n43599), .B(n43600), .Z(n39986) );
  XOR U40542 ( .A(n39989), .B(n39988), .Z(n39987) );
  AND U40543 ( .A(n43601), .B(n43602), .Z(n39988) );
  XOR U40544 ( .A(n39991), .B(n39990), .Z(n39989) );
  AND U40545 ( .A(n43603), .B(n43604), .Z(n39990) );
  XOR U40546 ( .A(n39993), .B(n39992), .Z(n39991) );
  AND U40547 ( .A(n43605), .B(n43606), .Z(n39992) );
  XOR U40548 ( .A(n39995), .B(n39994), .Z(n39993) );
  AND U40549 ( .A(n43607), .B(n43608), .Z(n39994) );
  XOR U40550 ( .A(n39997), .B(n39996), .Z(n39995) );
  AND U40551 ( .A(n43609), .B(n43610), .Z(n39996) );
  XOR U40552 ( .A(n39999), .B(n39998), .Z(n39997) );
  AND U40553 ( .A(n43611), .B(n43612), .Z(n39998) );
  XOR U40554 ( .A(n40001), .B(n40000), .Z(n39999) );
  AND U40555 ( .A(n43613), .B(n43614), .Z(n40000) );
  XOR U40556 ( .A(n40003), .B(n40002), .Z(n40001) );
  AND U40557 ( .A(n43615), .B(n43616), .Z(n40002) );
  XOR U40558 ( .A(n40005), .B(n40004), .Z(n40003) );
  AND U40559 ( .A(n43617), .B(n43618), .Z(n40004) );
  XOR U40560 ( .A(n40007), .B(n40006), .Z(n40005) );
  AND U40561 ( .A(n43619), .B(n43620), .Z(n40006) );
  XOR U40562 ( .A(n40009), .B(n40008), .Z(n40007) );
  AND U40563 ( .A(n43621), .B(n43622), .Z(n40008) );
  XOR U40564 ( .A(n40011), .B(n40010), .Z(n40009) );
  AND U40565 ( .A(n43623), .B(n43624), .Z(n40010) );
  XOR U40566 ( .A(n40013), .B(n40012), .Z(n40011) );
  AND U40567 ( .A(n43625), .B(n43626), .Z(n40012) );
  XOR U40568 ( .A(n40015), .B(n40014), .Z(n40013) );
  AND U40569 ( .A(n43627), .B(n43628), .Z(n40014) );
  XOR U40570 ( .A(n40017), .B(n40016), .Z(n40015) );
  AND U40571 ( .A(n43629), .B(n43630), .Z(n40016) );
  XOR U40572 ( .A(n40019), .B(n40018), .Z(n40017) );
  AND U40573 ( .A(n43631), .B(n43632), .Z(n40018) );
  XOR U40574 ( .A(n40021), .B(n40020), .Z(n40019) );
  AND U40575 ( .A(n43633), .B(n43634), .Z(n40020) );
  XOR U40576 ( .A(n40023), .B(n40022), .Z(n40021) );
  AND U40577 ( .A(n43635), .B(n43636), .Z(n40022) );
  XOR U40578 ( .A(n40025), .B(n40024), .Z(n40023) );
  AND U40579 ( .A(n43637), .B(n43638), .Z(n40024) );
  XOR U40580 ( .A(n40027), .B(n40026), .Z(n40025) );
  AND U40581 ( .A(n43639), .B(n43640), .Z(n40026) );
  XOR U40582 ( .A(n40029), .B(n40028), .Z(n40027) );
  AND U40583 ( .A(n43641), .B(n43642), .Z(n40028) );
  XOR U40584 ( .A(n40031), .B(n40030), .Z(n40029) );
  AND U40585 ( .A(n43643), .B(n43644), .Z(n40030) );
  XOR U40586 ( .A(n40033), .B(n40032), .Z(n40031) );
  AND U40587 ( .A(n43645), .B(n43646), .Z(n40032) );
  XOR U40588 ( .A(n40035), .B(n40034), .Z(n40033) );
  AND U40589 ( .A(n43647), .B(n43648), .Z(n40034) );
  XOR U40590 ( .A(n40037), .B(n40036), .Z(n40035) );
  AND U40591 ( .A(n43649), .B(n43650), .Z(n40036) );
  XOR U40592 ( .A(n40065), .B(n40038), .Z(n40037) );
  AND U40593 ( .A(n43651), .B(n43652), .Z(n40038) );
  XOR U40594 ( .A(n40067), .B(n40066), .Z(n40065) );
  AND U40595 ( .A(n43653), .B(n43654), .Z(n40066) );
  XOR U40596 ( .A(n40046), .B(n40068), .Z(n40067) );
  AND U40597 ( .A(n43655), .B(n43656), .Z(n40068) );
  XOR U40598 ( .A(n40042), .B(n40047), .Z(n40046) );
  AND U40599 ( .A(n43657), .B(n43658), .Z(n40047) );
  XOR U40600 ( .A(n40044), .B(n40043), .Z(n40042) );
  AND U40601 ( .A(n43659), .B(n43660), .Z(n40043) );
  XNOR U40602 ( .A(n40054), .B(n40045), .Z(n40044) );
  AND U40603 ( .A(n43661), .B(n43662), .Z(n40045) );
  XOR U40604 ( .A(n40064), .B(n40053), .Z(n40054) );
  AND U40605 ( .A(n43663), .B(n43664), .Z(n40053) );
  XNOR U40606 ( .A(n43665), .B(n40059), .Z(n40064) );
  XOR U40607 ( .A(n40060), .B(n43666), .Z(n40059) );
  AND U40608 ( .A(n43667), .B(n43668), .Z(n43666) );
  XOR U40609 ( .A(n43669), .B(n43670), .Z(n40060) );
  NOR U40610 ( .A(n43671), .B(n43672), .Z(n43670) );
  AND U40611 ( .A(n43673), .B(n43674), .Z(n43672) );
  AND U40612 ( .A(n43675), .B(n43676), .Z(n43671) );
  XNOR U40613 ( .A(n43673), .B(n43674), .Z(n43669) );
  XNOR U40614 ( .A(n40051), .B(n40063), .Z(n43665) );
  AND U40615 ( .A(n43677), .B(n43678), .Z(n40063) );
  AND U40616 ( .A(n43679), .B(n43680), .Z(n40051) );
  XNOR U40617 ( .A(n42647), .B(n135), .Z(n42649) );
  XOR U40618 ( .A(n42644), .B(n42645), .Z(n135) );
  AND U40619 ( .A(n43681), .B(n43682), .Z(n42645) );
  XOR U40620 ( .A(n42641), .B(n42642), .Z(n42644) );
  AND U40621 ( .A(n43683), .B(n43684), .Z(n42642) );
  XOR U40622 ( .A(n42638), .B(n42639), .Z(n42641) );
  AND U40623 ( .A(n43685), .B(n43686), .Z(n42639) );
  XOR U40624 ( .A(n42635), .B(n42636), .Z(n42638) );
  AND U40625 ( .A(n43687), .B(n43688), .Z(n42636) );
  XOR U40626 ( .A(n42632), .B(n42633), .Z(n42635) );
  AND U40627 ( .A(n43689), .B(n43690), .Z(n42633) );
  XOR U40628 ( .A(n42629), .B(n42630), .Z(n42632) );
  AND U40629 ( .A(n43691), .B(n43692), .Z(n42630) );
  XOR U40630 ( .A(n42626), .B(n42627), .Z(n42629) );
  AND U40631 ( .A(n43693), .B(n43694), .Z(n42627) );
  XOR U40632 ( .A(n42623), .B(n42624), .Z(n42626) );
  AND U40633 ( .A(n43695), .B(n43696), .Z(n42624) );
  XOR U40634 ( .A(n42620), .B(n42621), .Z(n42623) );
  AND U40635 ( .A(n43697), .B(n43698), .Z(n42621) );
  XOR U40636 ( .A(n42617), .B(n42618), .Z(n42620) );
  AND U40637 ( .A(n43699), .B(n43700), .Z(n42618) );
  XOR U40638 ( .A(n42614), .B(n42615), .Z(n42617) );
  AND U40639 ( .A(n43701), .B(n43702), .Z(n42615) );
  XOR U40640 ( .A(n42611), .B(n42612), .Z(n42614) );
  AND U40641 ( .A(n43703), .B(n43704), .Z(n42612) );
  XOR U40642 ( .A(n42608), .B(n42609), .Z(n42611) );
  AND U40643 ( .A(n43705), .B(n43706), .Z(n42609) );
  XOR U40644 ( .A(n42605), .B(n42606), .Z(n42608) );
  AND U40645 ( .A(n43707), .B(n43708), .Z(n42606) );
  XOR U40646 ( .A(n42602), .B(n42603), .Z(n42605) );
  AND U40647 ( .A(n43709), .B(n43710), .Z(n42603) );
  XOR U40648 ( .A(n42599), .B(n42600), .Z(n42602) );
  AND U40649 ( .A(n43711), .B(n43712), .Z(n42600) );
  XOR U40650 ( .A(n42596), .B(n42597), .Z(n42599) );
  AND U40651 ( .A(n43713), .B(n43714), .Z(n42597) );
  XOR U40652 ( .A(n42593), .B(n42594), .Z(n42596) );
  AND U40653 ( .A(n43715), .B(n43716), .Z(n42594) );
  XOR U40654 ( .A(n42590), .B(n42591), .Z(n42593) );
  AND U40655 ( .A(n43717), .B(n43718), .Z(n42591) );
  XOR U40656 ( .A(n42587), .B(n42588), .Z(n42590) );
  AND U40657 ( .A(n43719), .B(n43720), .Z(n42588) );
  XOR U40658 ( .A(n42584), .B(n42585), .Z(n42587) );
  AND U40659 ( .A(n43721), .B(n43722), .Z(n42585) );
  XOR U40660 ( .A(n42581), .B(n42582), .Z(n42584) );
  AND U40661 ( .A(n43723), .B(n43724), .Z(n42582) );
  XOR U40662 ( .A(n42578), .B(n42579), .Z(n42581) );
  AND U40663 ( .A(n43725), .B(n43726), .Z(n42579) );
  XOR U40664 ( .A(n42575), .B(n42576), .Z(n42578) );
  AND U40665 ( .A(n43727), .B(n43728), .Z(n42576) );
  XOR U40666 ( .A(n42572), .B(n42573), .Z(n42575) );
  AND U40667 ( .A(n43729), .B(n43730), .Z(n42573) );
  XOR U40668 ( .A(n42569), .B(n42570), .Z(n42572) );
  AND U40669 ( .A(n43731), .B(n43732), .Z(n42570) );
  XOR U40670 ( .A(n42566), .B(n42567), .Z(n42569) );
  AND U40671 ( .A(n43733), .B(n43734), .Z(n42567) );
  XOR U40672 ( .A(n42563), .B(n42564), .Z(n42566) );
  AND U40673 ( .A(n43735), .B(n43736), .Z(n42564) );
  XOR U40674 ( .A(n42560), .B(n42561), .Z(n42563) );
  AND U40675 ( .A(n43737), .B(n43738), .Z(n42561) );
  XOR U40676 ( .A(n42557), .B(n42558), .Z(n42560) );
  AND U40677 ( .A(n43739), .B(n43740), .Z(n42558) );
  XOR U40678 ( .A(n42554), .B(n42555), .Z(n42557) );
  AND U40679 ( .A(n43741), .B(n43742), .Z(n42555) );
  XOR U40680 ( .A(n42551), .B(n42552), .Z(n42554) );
  AND U40681 ( .A(n43743), .B(n43744), .Z(n42552) );
  XOR U40682 ( .A(n42548), .B(n42549), .Z(n42551) );
  AND U40683 ( .A(n43745), .B(n43746), .Z(n42549) );
  XOR U40684 ( .A(n42545), .B(n42546), .Z(n42548) );
  AND U40685 ( .A(n43747), .B(n43748), .Z(n42546) );
  XOR U40686 ( .A(n42542), .B(n42543), .Z(n42545) );
  AND U40687 ( .A(n43749), .B(n43750), .Z(n42543) );
  XOR U40688 ( .A(n42539), .B(n42540), .Z(n42542) );
  AND U40689 ( .A(n43751), .B(n43752), .Z(n42540) );
  XOR U40690 ( .A(n42536), .B(n42537), .Z(n42539) );
  AND U40691 ( .A(n43753), .B(n43754), .Z(n42537) );
  XOR U40692 ( .A(n42533), .B(n42534), .Z(n42536) );
  AND U40693 ( .A(n43755), .B(n43756), .Z(n42534) );
  XOR U40694 ( .A(n42530), .B(n42531), .Z(n42533) );
  AND U40695 ( .A(n43757), .B(n43758), .Z(n42531) );
  XOR U40696 ( .A(n42527), .B(n42528), .Z(n42530) );
  AND U40697 ( .A(n43759), .B(n43760), .Z(n42528) );
  XOR U40698 ( .A(n42524), .B(n42525), .Z(n42527) );
  AND U40699 ( .A(n43761), .B(n43762), .Z(n42525) );
  XOR U40700 ( .A(n42521), .B(n42522), .Z(n42524) );
  AND U40701 ( .A(n43763), .B(n43764), .Z(n42522) );
  XOR U40702 ( .A(n42518), .B(n42519), .Z(n42521) );
  AND U40703 ( .A(n43765), .B(n43766), .Z(n42519) );
  XOR U40704 ( .A(n42515), .B(n42516), .Z(n42518) );
  AND U40705 ( .A(n43767), .B(n43768), .Z(n42516) );
  XOR U40706 ( .A(n42512), .B(n42513), .Z(n42515) );
  AND U40707 ( .A(n43769), .B(n43770), .Z(n42513) );
  XOR U40708 ( .A(n42509), .B(n42510), .Z(n42512) );
  AND U40709 ( .A(n43771), .B(n43772), .Z(n42510) );
  XOR U40710 ( .A(n42506), .B(n42507), .Z(n42509) );
  AND U40711 ( .A(n43773), .B(n43774), .Z(n42507) );
  XOR U40712 ( .A(n42503), .B(n42504), .Z(n42506) );
  AND U40713 ( .A(n43775), .B(n43776), .Z(n42504) );
  XOR U40714 ( .A(n42500), .B(n42501), .Z(n42503) );
  AND U40715 ( .A(n43777), .B(n43778), .Z(n42501) );
  XOR U40716 ( .A(n42497), .B(n42498), .Z(n42500) );
  AND U40717 ( .A(n43779), .B(n43780), .Z(n42498) );
  XOR U40718 ( .A(n42494), .B(n42495), .Z(n42497) );
  AND U40719 ( .A(n43781), .B(n43782), .Z(n42495) );
  XOR U40720 ( .A(n42491), .B(n42492), .Z(n42494) );
  AND U40721 ( .A(n43783), .B(n43784), .Z(n42492) );
  XOR U40722 ( .A(n42488), .B(n42489), .Z(n42491) );
  AND U40723 ( .A(n43785), .B(n43786), .Z(n42489) );
  XOR U40724 ( .A(n42485), .B(n42486), .Z(n42488) );
  AND U40725 ( .A(n43787), .B(n43788), .Z(n42486) );
  XOR U40726 ( .A(n42482), .B(n42483), .Z(n42485) );
  AND U40727 ( .A(n43789), .B(n43790), .Z(n42483) );
  XOR U40728 ( .A(n42479), .B(n42480), .Z(n42482) );
  AND U40729 ( .A(n43791), .B(n43792), .Z(n42480) );
  XOR U40730 ( .A(n42476), .B(n42477), .Z(n42479) );
  AND U40731 ( .A(n43793), .B(n43794), .Z(n42477) );
  XOR U40732 ( .A(n42473), .B(n42474), .Z(n42476) );
  AND U40733 ( .A(n43795), .B(n43796), .Z(n42474) );
  XOR U40734 ( .A(n42470), .B(n42471), .Z(n42473) );
  AND U40735 ( .A(n43797), .B(n43798), .Z(n42471) );
  XOR U40736 ( .A(n42467), .B(n42468), .Z(n42470) );
  AND U40737 ( .A(n43799), .B(n43800), .Z(n42468) );
  XOR U40738 ( .A(n42464), .B(n42465), .Z(n42467) );
  AND U40739 ( .A(n43801), .B(n43802), .Z(n42465) );
  XOR U40740 ( .A(n42461), .B(n42462), .Z(n42464) );
  AND U40741 ( .A(n43803), .B(n43804), .Z(n42462) );
  XOR U40742 ( .A(n42458), .B(n42459), .Z(n42461) );
  AND U40743 ( .A(n43805), .B(n43806), .Z(n42459) );
  XOR U40744 ( .A(n42455), .B(n42456), .Z(n42458) );
  AND U40745 ( .A(n43807), .B(n43808), .Z(n42456) );
  XOR U40746 ( .A(n42452), .B(n42453), .Z(n42455) );
  AND U40747 ( .A(n43809), .B(n43810), .Z(n42453) );
  XOR U40748 ( .A(n42449), .B(n42450), .Z(n42452) );
  AND U40749 ( .A(n43811), .B(n43812), .Z(n42450) );
  XOR U40750 ( .A(n42446), .B(n42447), .Z(n42449) );
  AND U40751 ( .A(n43813), .B(n43814), .Z(n42447) );
  XOR U40752 ( .A(n42443), .B(n42444), .Z(n42446) );
  AND U40753 ( .A(n43815), .B(n43816), .Z(n42444) );
  XOR U40754 ( .A(n42440), .B(n42441), .Z(n42443) );
  AND U40755 ( .A(n43817), .B(n43818), .Z(n42441) );
  XOR U40756 ( .A(n42437), .B(n42438), .Z(n42440) );
  AND U40757 ( .A(n43819), .B(n43820), .Z(n42438) );
  XOR U40758 ( .A(n42434), .B(n42435), .Z(n42437) );
  AND U40759 ( .A(n43821), .B(n43822), .Z(n42435) );
  XOR U40760 ( .A(n42431), .B(n42432), .Z(n42434) );
  AND U40761 ( .A(n43823), .B(n43824), .Z(n42432) );
  XOR U40762 ( .A(n42428), .B(n42429), .Z(n42431) );
  AND U40763 ( .A(n43825), .B(n43826), .Z(n42429) );
  XOR U40764 ( .A(n42425), .B(n42426), .Z(n42428) );
  AND U40765 ( .A(n43827), .B(n43828), .Z(n42426) );
  XOR U40766 ( .A(n42422), .B(n42423), .Z(n42425) );
  AND U40767 ( .A(n43829), .B(n43830), .Z(n42423) );
  XOR U40768 ( .A(n42419), .B(n42420), .Z(n42422) );
  AND U40769 ( .A(n43831), .B(n43832), .Z(n42420) );
  XOR U40770 ( .A(n42416), .B(n42417), .Z(n42419) );
  AND U40771 ( .A(n43833), .B(n43834), .Z(n42417) );
  XOR U40772 ( .A(n42413), .B(n42414), .Z(n42416) );
  AND U40773 ( .A(n43835), .B(n43836), .Z(n42414) );
  XOR U40774 ( .A(n42410), .B(n42411), .Z(n42413) );
  AND U40775 ( .A(n43837), .B(n43838), .Z(n42411) );
  XOR U40776 ( .A(n42407), .B(n42408), .Z(n42410) );
  AND U40777 ( .A(n43839), .B(n43840), .Z(n42408) );
  XOR U40778 ( .A(n42404), .B(n42405), .Z(n42407) );
  AND U40779 ( .A(n43841), .B(n43842), .Z(n42405) );
  XOR U40780 ( .A(n42401), .B(n42402), .Z(n42404) );
  AND U40781 ( .A(n43843), .B(n43844), .Z(n42402) );
  XOR U40782 ( .A(n42398), .B(n42399), .Z(n42401) );
  AND U40783 ( .A(n43845), .B(n43846), .Z(n42399) );
  XOR U40784 ( .A(n42395), .B(n42396), .Z(n42398) );
  AND U40785 ( .A(n43847), .B(n43848), .Z(n42396) );
  XOR U40786 ( .A(n42392), .B(n42393), .Z(n42395) );
  AND U40787 ( .A(n43849), .B(n43850), .Z(n42393) );
  XOR U40788 ( .A(n42389), .B(n42390), .Z(n42392) );
  AND U40789 ( .A(n43851), .B(n43852), .Z(n42390) );
  XOR U40790 ( .A(n42386), .B(n42387), .Z(n42389) );
  AND U40791 ( .A(n43853), .B(n43854), .Z(n42387) );
  XOR U40792 ( .A(n42383), .B(n42384), .Z(n42386) );
  AND U40793 ( .A(n43855), .B(n43856), .Z(n42384) );
  XOR U40794 ( .A(n42380), .B(n42381), .Z(n42383) );
  AND U40795 ( .A(n43857), .B(n43858), .Z(n42381) );
  XOR U40796 ( .A(n42377), .B(n42378), .Z(n42380) );
  AND U40797 ( .A(n43859), .B(n43860), .Z(n42378) );
  XOR U40798 ( .A(n42374), .B(n42375), .Z(n42377) );
  AND U40799 ( .A(n43861), .B(n43862), .Z(n42375) );
  XOR U40800 ( .A(n42371), .B(n42372), .Z(n42374) );
  AND U40801 ( .A(n43863), .B(n43864), .Z(n42372) );
  XOR U40802 ( .A(n42368), .B(n42369), .Z(n42371) );
  AND U40803 ( .A(n43865), .B(n43866), .Z(n42369) );
  XOR U40804 ( .A(n42365), .B(n42366), .Z(n42368) );
  AND U40805 ( .A(n43867), .B(n43868), .Z(n42366) );
  XOR U40806 ( .A(n42362), .B(n42363), .Z(n42365) );
  AND U40807 ( .A(n43869), .B(n43870), .Z(n42363) );
  XOR U40808 ( .A(n42359), .B(n42360), .Z(n42362) );
  AND U40809 ( .A(n43871), .B(n43872), .Z(n42360) );
  XOR U40810 ( .A(n42356), .B(n42357), .Z(n42359) );
  AND U40811 ( .A(n43873), .B(n43874), .Z(n42357) );
  XOR U40812 ( .A(n42353), .B(n42354), .Z(n42356) );
  AND U40813 ( .A(n43875), .B(n43876), .Z(n42354) );
  XOR U40814 ( .A(n42350), .B(n42351), .Z(n42353) );
  AND U40815 ( .A(n43877), .B(n43878), .Z(n42351) );
  XOR U40816 ( .A(n42347), .B(n42348), .Z(n42350) );
  AND U40817 ( .A(n43879), .B(n43880), .Z(n42348) );
  XOR U40818 ( .A(n42344), .B(n42345), .Z(n42347) );
  AND U40819 ( .A(n43881), .B(n43882), .Z(n42345) );
  XOR U40820 ( .A(n42341), .B(n42342), .Z(n42344) );
  AND U40821 ( .A(n43883), .B(n43884), .Z(n42342) );
  XOR U40822 ( .A(n42338), .B(n42339), .Z(n42341) );
  AND U40823 ( .A(n43885), .B(n43886), .Z(n42339) );
  XOR U40824 ( .A(n42335), .B(n42336), .Z(n42338) );
  AND U40825 ( .A(n43887), .B(n43888), .Z(n42336) );
  XOR U40826 ( .A(n42332), .B(n42333), .Z(n42335) );
  AND U40827 ( .A(n43889), .B(n43890), .Z(n42333) );
  XOR U40828 ( .A(n42329), .B(n42330), .Z(n42332) );
  AND U40829 ( .A(n43891), .B(n43892), .Z(n42330) );
  XOR U40830 ( .A(n42326), .B(n42327), .Z(n42329) );
  AND U40831 ( .A(n43893), .B(n43894), .Z(n42327) );
  XOR U40832 ( .A(n42323), .B(n42324), .Z(n42326) );
  AND U40833 ( .A(n43895), .B(n43896), .Z(n42324) );
  XOR U40834 ( .A(n42320), .B(n42321), .Z(n42323) );
  AND U40835 ( .A(n43897), .B(n43898), .Z(n42321) );
  XOR U40836 ( .A(n42317), .B(n42318), .Z(n42320) );
  AND U40837 ( .A(n43899), .B(n43900), .Z(n42318) );
  XOR U40838 ( .A(n42314), .B(n42315), .Z(n42317) );
  AND U40839 ( .A(n43901), .B(n43902), .Z(n42315) );
  XOR U40840 ( .A(n42311), .B(n42312), .Z(n42314) );
  AND U40841 ( .A(n43903), .B(n43904), .Z(n42312) );
  XOR U40842 ( .A(n42308), .B(n42309), .Z(n42311) );
  AND U40843 ( .A(n43905), .B(n43906), .Z(n42309) );
  XOR U40844 ( .A(n42305), .B(n42306), .Z(n42308) );
  AND U40845 ( .A(n43907), .B(n43908), .Z(n42306) );
  XOR U40846 ( .A(n42302), .B(n42303), .Z(n42305) );
  AND U40847 ( .A(n43909), .B(n43910), .Z(n42303) );
  XOR U40848 ( .A(n42299), .B(n42300), .Z(n42302) );
  AND U40849 ( .A(n43911), .B(n43912), .Z(n42300) );
  XOR U40850 ( .A(n42296), .B(n42297), .Z(n42299) );
  AND U40851 ( .A(n43913), .B(n43914), .Z(n42297) );
  XOR U40852 ( .A(n42293), .B(n42294), .Z(n42296) );
  AND U40853 ( .A(n43915), .B(n43916), .Z(n42294) );
  XOR U40854 ( .A(n42290), .B(n42291), .Z(n42293) );
  AND U40855 ( .A(n43917), .B(n43918), .Z(n42291) );
  XOR U40856 ( .A(n42287), .B(n42288), .Z(n42290) );
  AND U40857 ( .A(n43919), .B(n43920), .Z(n42288) );
  XOR U40858 ( .A(n42284), .B(n42285), .Z(n42287) );
  AND U40859 ( .A(n43921), .B(n43922), .Z(n42285) );
  XOR U40860 ( .A(n42281), .B(n42282), .Z(n42284) );
  AND U40861 ( .A(n43923), .B(n43924), .Z(n42282) );
  XOR U40862 ( .A(n42278), .B(n42279), .Z(n42281) );
  AND U40863 ( .A(n43925), .B(n43926), .Z(n42279) );
  XOR U40864 ( .A(n42275), .B(n42276), .Z(n42278) );
  AND U40865 ( .A(n43927), .B(n43928), .Z(n42276) );
  XOR U40866 ( .A(n42272), .B(n42273), .Z(n42275) );
  AND U40867 ( .A(n43929), .B(n43930), .Z(n42273) );
  XOR U40868 ( .A(n42269), .B(n42270), .Z(n42272) );
  AND U40869 ( .A(n43931), .B(n43932), .Z(n42270) );
  XOR U40870 ( .A(n42266), .B(n42267), .Z(n42269) );
  AND U40871 ( .A(n43933), .B(n43934), .Z(n42267) );
  XOR U40872 ( .A(n42263), .B(n42264), .Z(n42266) );
  AND U40873 ( .A(n43935), .B(n43936), .Z(n42264) );
  XOR U40874 ( .A(n42260), .B(n42261), .Z(n42263) );
  AND U40875 ( .A(n43937), .B(n43938), .Z(n42261) );
  XOR U40876 ( .A(n42257), .B(n42258), .Z(n42260) );
  AND U40877 ( .A(n43939), .B(n43940), .Z(n42258) );
  XOR U40878 ( .A(n42254), .B(n42255), .Z(n42257) );
  AND U40879 ( .A(n43941), .B(n43942), .Z(n42255) );
  XOR U40880 ( .A(n42251), .B(n42252), .Z(n42254) );
  AND U40881 ( .A(n43943), .B(n43944), .Z(n42252) );
  XOR U40882 ( .A(n42248), .B(n42249), .Z(n42251) );
  AND U40883 ( .A(n43945), .B(n43946), .Z(n42249) );
  XOR U40884 ( .A(n42245), .B(n42246), .Z(n42248) );
  AND U40885 ( .A(n43947), .B(n43948), .Z(n42246) );
  XOR U40886 ( .A(n42242), .B(n42243), .Z(n42245) );
  AND U40887 ( .A(n43949), .B(n43950), .Z(n42243) );
  XOR U40888 ( .A(n42239), .B(n42240), .Z(n42242) );
  AND U40889 ( .A(n43951), .B(n43952), .Z(n42240) );
  XOR U40890 ( .A(n42236), .B(n42237), .Z(n42239) );
  AND U40891 ( .A(n43953), .B(n43954), .Z(n42237) );
  XOR U40892 ( .A(n42233), .B(n42234), .Z(n42236) );
  AND U40893 ( .A(n43955), .B(n43956), .Z(n42234) );
  XOR U40894 ( .A(n42230), .B(n42231), .Z(n42233) );
  AND U40895 ( .A(n43957), .B(n43958), .Z(n42231) );
  XOR U40896 ( .A(n42227), .B(n42228), .Z(n42230) );
  AND U40897 ( .A(n43959), .B(n43960), .Z(n42228) );
  XOR U40898 ( .A(n42224), .B(n42225), .Z(n42227) );
  AND U40899 ( .A(n43961), .B(n43962), .Z(n42225) );
  XOR U40900 ( .A(n42221), .B(n42222), .Z(n42224) );
  AND U40901 ( .A(n43963), .B(n43964), .Z(n42222) );
  XOR U40902 ( .A(n42218), .B(n42219), .Z(n42221) );
  AND U40903 ( .A(n43965), .B(n43966), .Z(n42219) );
  XOR U40904 ( .A(n42215), .B(n42216), .Z(n42218) );
  AND U40905 ( .A(n43967), .B(n43968), .Z(n42216) );
  XOR U40906 ( .A(n42212), .B(n42213), .Z(n42215) );
  AND U40907 ( .A(n43969), .B(n43970), .Z(n42213) );
  XOR U40908 ( .A(n42209), .B(n42210), .Z(n42212) );
  AND U40909 ( .A(n43971), .B(n43972), .Z(n42210) );
  XOR U40910 ( .A(n42206), .B(n42207), .Z(n42209) );
  AND U40911 ( .A(n43973), .B(n43974), .Z(n42207) );
  XOR U40912 ( .A(n42203), .B(n42204), .Z(n42206) );
  AND U40913 ( .A(n43975), .B(n43976), .Z(n42204) );
  XOR U40914 ( .A(n42200), .B(n42201), .Z(n42203) );
  AND U40915 ( .A(n43977), .B(n43978), .Z(n42201) );
  XOR U40916 ( .A(n42197), .B(n42198), .Z(n42200) );
  AND U40917 ( .A(n43979), .B(n43980), .Z(n42198) );
  XOR U40918 ( .A(n42194), .B(n42195), .Z(n42197) );
  AND U40919 ( .A(n43981), .B(n43982), .Z(n42195) );
  XOR U40920 ( .A(n42191), .B(n42192), .Z(n42194) );
  AND U40921 ( .A(n43983), .B(n43984), .Z(n42192) );
  XOR U40922 ( .A(n42188), .B(n42189), .Z(n42191) );
  AND U40923 ( .A(n43985), .B(n43986), .Z(n42189) );
  XOR U40924 ( .A(n42185), .B(n42186), .Z(n42188) );
  AND U40925 ( .A(n43987), .B(n43988), .Z(n42186) );
  XOR U40926 ( .A(n42182), .B(n42183), .Z(n42185) );
  AND U40927 ( .A(n43989), .B(n43990), .Z(n42183) );
  XOR U40928 ( .A(n42179), .B(n42180), .Z(n42182) );
  AND U40929 ( .A(n43991), .B(n43992), .Z(n42180) );
  XOR U40930 ( .A(n42176), .B(n42177), .Z(n42179) );
  AND U40931 ( .A(n43993), .B(n43994), .Z(n42177) );
  XOR U40932 ( .A(n42173), .B(n42174), .Z(n42176) );
  AND U40933 ( .A(n43995), .B(n43996), .Z(n42174) );
  XOR U40934 ( .A(n42170), .B(n42171), .Z(n42173) );
  AND U40935 ( .A(n43997), .B(n43998), .Z(n42171) );
  XOR U40936 ( .A(n42167), .B(n42168), .Z(n42170) );
  AND U40937 ( .A(n43999), .B(n44000), .Z(n42168) );
  XOR U40938 ( .A(n42164), .B(n42165), .Z(n42167) );
  AND U40939 ( .A(n44001), .B(n44002), .Z(n42165) );
  XOR U40940 ( .A(n42161), .B(n42162), .Z(n42164) );
  AND U40941 ( .A(n44003), .B(n44004), .Z(n42162) );
  XOR U40942 ( .A(n42158), .B(n42159), .Z(n42161) );
  AND U40943 ( .A(n44005), .B(n44006), .Z(n42159) );
  XOR U40944 ( .A(n42155), .B(n42156), .Z(n42158) );
  AND U40945 ( .A(n44007), .B(n44008), .Z(n42156) );
  XOR U40946 ( .A(n42152), .B(n42153), .Z(n42155) );
  AND U40947 ( .A(n44009), .B(n44010), .Z(n42153) );
  XOR U40948 ( .A(n42149), .B(n42150), .Z(n42152) );
  AND U40949 ( .A(n44011), .B(n44012), .Z(n42150) );
  XOR U40950 ( .A(n42146), .B(n42147), .Z(n42149) );
  AND U40951 ( .A(n44013), .B(n44014), .Z(n42147) );
  XOR U40952 ( .A(n42143), .B(n42144), .Z(n42146) );
  AND U40953 ( .A(n44015), .B(n44016), .Z(n42144) );
  XOR U40954 ( .A(n42140), .B(n42141), .Z(n42143) );
  AND U40955 ( .A(n44017), .B(n44018), .Z(n42141) );
  XOR U40956 ( .A(n42137), .B(n42138), .Z(n42140) );
  AND U40957 ( .A(n44019), .B(n44020), .Z(n42138) );
  XOR U40958 ( .A(n42134), .B(n42135), .Z(n42137) );
  AND U40959 ( .A(n44021), .B(n44022), .Z(n42135) );
  XOR U40960 ( .A(n42131), .B(n42132), .Z(n42134) );
  AND U40961 ( .A(n44023), .B(n44024), .Z(n42132) );
  XOR U40962 ( .A(n42128), .B(n42129), .Z(n42131) );
  AND U40963 ( .A(n44025), .B(n44026), .Z(n42129) );
  XOR U40964 ( .A(n42125), .B(n42126), .Z(n42128) );
  AND U40965 ( .A(n44027), .B(n44028), .Z(n42126) );
  XOR U40966 ( .A(n42122), .B(n42123), .Z(n42125) );
  AND U40967 ( .A(n44029), .B(n44030), .Z(n42123) );
  XOR U40968 ( .A(n42119), .B(n42120), .Z(n42122) );
  AND U40969 ( .A(n44031), .B(n44032), .Z(n42120) );
  XOR U40970 ( .A(n42116), .B(n42117), .Z(n42119) );
  AND U40971 ( .A(n44033), .B(n44034), .Z(n42117) );
  XOR U40972 ( .A(n42113), .B(n42114), .Z(n42116) );
  AND U40973 ( .A(n44035), .B(n44036), .Z(n42114) );
  XOR U40974 ( .A(n42110), .B(n42111), .Z(n42113) );
  AND U40975 ( .A(n44037), .B(n44038), .Z(n42111) );
  XOR U40976 ( .A(n42107), .B(n42108), .Z(n42110) );
  AND U40977 ( .A(n44039), .B(n44040), .Z(n42108) );
  XOR U40978 ( .A(n42104), .B(n42105), .Z(n42107) );
  AND U40979 ( .A(n44041), .B(n44042), .Z(n42105) );
  XOR U40980 ( .A(n42101), .B(n42102), .Z(n42104) );
  AND U40981 ( .A(n44043), .B(n44044), .Z(n42102) );
  XOR U40982 ( .A(n42098), .B(n42099), .Z(n42101) );
  AND U40983 ( .A(n44045), .B(n44046), .Z(n42099) );
  XOR U40984 ( .A(n42095), .B(n42096), .Z(n42098) );
  AND U40985 ( .A(n44047), .B(n44048), .Z(n42096) );
  XOR U40986 ( .A(n42092), .B(n42093), .Z(n42095) );
  AND U40987 ( .A(n44049), .B(n44050), .Z(n42093) );
  XOR U40988 ( .A(n42089), .B(n42090), .Z(n42092) );
  AND U40989 ( .A(n44051), .B(n44052), .Z(n42090) );
  XOR U40990 ( .A(n42086), .B(n42087), .Z(n42089) );
  AND U40991 ( .A(n44053), .B(n44054), .Z(n42087) );
  XOR U40992 ( .A(n42083), .B(n42084), .Z(n42086) );
  AND U40993 ( .A(n44055), .B(n44056), .Z(n42084) );
  XOR U40994 ( .A(n42080), .B(n42081), .Z(n42083) );
  AND U40995 ( .A(n44057), .B(n44058), .Z(n42081) );
  XOR U40996 ( .A(n42077), .B(n42078), .Z(n42080) );
  AND U40997 ( .A(n44059), .B(n44060), .Z(n42078) );
  XOR U40998 ( .A(n42074), .B(n42075), .Z(n42077) );
  AND U40999 ( .A(n44061), .B(n44062), .Z(n42075) );
  XOR U41000 ( .A(n42071), .B(n42072), .Z(n42074) );
  AND U41001 ( .A(n44063), .B(n44064), .Z(n42072) );
  XOR U41002 ( .A(n42068), .B(n42069), .Z(n42071) );
  AND U41003 ( .A(n44065), .B(n44066), .Z(n42069) );
  XOR U41004 ( .A(n42065), .B(n42066), .Z(n42068) );
  AND U41005 ( .A(n44067), .B(n44068), .Z(n42066) );
  XOR U41006 ( .A(n42062), .B(n42063), .Z(n42065) );
  AND U41007 ( .A(n44069), .B(n44070), .Z(n42063) );
  XOR U41008 ( .A(n42059), .B(n42060), .Z(n42062) );
  AND U41009 ( .A(n44071), .B(n44072), .Z(n42060) );
  XOR U41010 ( .A(n42056), .B(n42057), .Z(n42059) );
  AND U41011 ( .A(n44073), .B(n44074), .Z(n42057) );
  XOR U41012 ( .A(n42053), .B(n42054), .Z(n42056) );
  AND U41013 ( .A(n44075), .B(n44076), .Z(n42054) );
  XOR U41014 ( .A(n42050), .B(n42051), .Z(n42053) );
  AND U41015 ( .A(n44077), .B(n44078), .Z(n42051) );
  XOR U41016 ( .A(n42047), .B(n42048), .Z(n42050) );
  AND U41017 ( .A(n44079), .B(n44080), .Z(n42048) );
  XOR U41018 ( .A(n42044), .B(n42045), .Z(n42047) );
  AND U41019 ( .A(n44081), .B(n44082), .Z(n42045) );
  XOR U41020 ( .A(n42041), .B(n42042), .Z(n42044) );
  AND U41021 ( .A(n44083), .B(n44084), .Z(n42042) );
  XOR U41022 ( .A(n42038), .B(n42039), .Z(n42041) );
  AND U41023 ( .A(n44085), .B(n44086), .Z(n42039) );
  XOR U41024 ( .A(n42035), .B(n42036), .Z(n42038) );
  AND U41025 ( .A(n44087), .B(n44088), .Z(n42036) );
  XOR U41026 ( .A(n42032), .B(n42033), .Z(n42035) );
  AND U41027 ( .A(n44089), .B(n44090), .Z(n42033) );
  XOR U41028 ( .A(n42029), .B(n42030), .Z(n42032) );
  AND U41029 ( .A(n44091), .B(n44092), .Z(n42030) );
  XOR U41030 ( .A(n42026), .B(n42027), .Z(n42029) );
  AND U41031 ( .A(n44093), .B(n44094), .Z(n42027) );
  XOR U41032 ( .A(n42023), .B(n42024), .Z(n42026) );
  AND U41033 ( .A(n44095), .B(n44096), .Z(n42024) );
  XOR U41034 ( .A(n42020), .B(n42021), .Z(n42023) );
  AND U41035 ( .A(n44097), .B(n44098), .Z(n42021) );
  XOR U41036 ( .A(n42017), .B(n42018), .Z(n42020) );
  AND U41037 ( .A(n44099), .B(n44100), .Z(n42018) );
  XOR U41038 ( .A(n42014), .B(n42015), .Z(n42017) );
  AND U41039 ( .A(n44101), .B(n44102), .Z(n42015) );
  XOR U41040 ( .A(n42011), .B(n42012), .Z(n42014) );
  AND U41041 ( .A(n44103), .B(n44104), .Z(n42012) );
  XOR U41042 ( .A(n42008), .B(n42009), .Z(n42011) );
  AND U41043 ( .A(n44105), .B(n44106), .Z(n42009) );
  XOR U41044 ( .A(n42005), .B(n42006), .Z(n42008) );
  AND U41045 ( .A(n44107), .B(n44108), .Z(n42006) );
  XOR U41046 ( .A(n42002), .B(n42003), .Z(n42005) );
  AND U41047 ( .A(n44109), .B(n44110), .Z(n42003) );
  XOR U41048 ( .A(n41999), .B(n42000), .Z(n42002) );
  AND U41049 ( .A(n44111), .B(n44112), .Z(n42000) );
  XOR U41050 ( .A(n41996), .B(n41997), .Z(n41999) );
  AND U41051 ( .A(n44113), .B(n44114), .Z(n41997) );
  XOR U41052 ( .A(n41993), .B(n41994), .Z(n41996) );
  AND U41053 ( .A(n44115), .B(n44116), .Z(n41994) );
  XOR U41054 ( .A(n41990), .B(n41991), .Z(n41993) );
  AND U41055 ( .A(n44117), .B(n44118), .Z(n41991) );
  XOR U41056 ( .A(n41987), .B(n41988), .Z(n41990) );
  AND U41057 ( .A(n44119), .B(n44120), .Z(n41988) );
  XOR U41058 ( .A(n41984), .B(n41985), .Z(n41987) );
  AND U41059 ( .A(n44121), .B(n44122), .Z(n41985) );
  XOR U41060 ( .A(n41981), .B(n41982), .Z(n41984) );
  AND U41061 ( .A(n44123), .B(n44124), .Z(n41982) );
  XOR U41062 ( .A(n41978), .B(n41979), .Z(n41981) );
  AND U41063 ( .A(n44125), .B(n44126), .Z(n41979) );
  XOR U41064 ( .A(n41975), .B(n41976), .Z(n41978) );
  AND U41065 ( .A(n44127), .B(n44128), .Z(n41976) );
  XOR U41066 ( .A(n41972), .B(n41973), .Z(n41975) );
  AND U41067 ( .A(n44129), .B(n44130), .Z(n41973) );
  XOR U41068 ( .A(n41969), .B(n41970), .Z(n41972) );
  AND U41069 ( .A(n44131), .B(n44132), .Z(n41970) );
  XOR U41070 ( .A(n41966), .B(n41967), .Z(n41969) );
  AND U41071 ( .A(n44133), .B(n44134), .Z(n41967) );
  XOR U41072 ( .A(n41963), .B(n41964), .Z(n41966) );
  AND U41073 ( .A(n44135), .B(n44136), .Z(n41964) );
  XOR U41074 ( .A(n41960), .B(n41961), .Z(n41963) );
  AND U41075 ( .A(n44137), .B(n44138), .Z(n41961) );
  XOR U41076 ( .A(n41957), .B(n41958), .Z(n41960) );
  AND U41077 ( .A(n44139), .B(n44140), .Z(n41958) );
  XOR U41078 ( .A(n41954), .B(n41955), .Z(n41957) );
  AND U41079 ( .A(n44141), .B(n44142), .Z(n41955) );
  XOR U41080 ( .A(n41951), .B(n41952), .Z(n41954) );
  AND U41081 ( .A(n44143), .B(n44144), .Z(n41952) );
  XOR U41082 ( .A(n41948), .B(n41949), .Z(n41951) );
  AND U41083 ( .A(n44145), .B(n44146), .Z(n41949) );
  XOR U41084 ( .A(n41945), .B(n41946), .Z(n41948) );
  AND U41085 ( .A(n44147), .B(n44148), .Z(n41946) );
  XOR U41086 ( .A(n41942), .B(n41943), .Z(n41945) );
  AND U41087 ( .A(n44149), .B(n44150), .Z(n41943) );
  XOR U41088 ( .A(n41939), .B(n41940), .Z(n41942) );
  AND U41089 ( .A(n44151), .B(n44152), .Z(n41940) );
  XOR U41090 ( .A(n41936), .B(n41937), .Z(n41939) );
  AND U41091 ( .A(n44153), .B(n44154), .Z(n41937) );
  XOR U41092 ( .A(n41933), .B(n41934), .Z(n41936) );
  AND U41093 ( .A(n44155), .B(n44156), .Z(n41934) );
  XOR U41094 ( .A(n41930), .B(n41931), .Z(n41933) );
  AND U41095 ( .A(n44157), .B(n44158), .Z(n41931) );
  XOR U41096 ( .A(n41927), .B(n41928), .Z(n41930) );
  AND U41097 ( .A(n44159), .B(n44160), .Z(n41928) );
  XOR U41098 ( .A(n41924), .B(n41925), .Z(n41927) );
  AND U41099 ( .A(n44161), .B(n44162), .Z(n41925) );
  XOR U41100 ( .A(n41921), .B(n41922), .Z(n41924) );
  AND U41101 ( .A(n44163), .B(n44164), .Z(n41922) );
  XOR U41102 ( .A(n41918), .B(n41919), .Z(n41921) );
  AND U41103 ( .A(n44165), .B(n44166), .Z(n41919) );
  XOR U41104 ( .A(n41915), .B(n41916), .Z(n41918) );
  AND U41105 ( .A(n44167), .B(n44168), .Z(n41916) );
  XOR U41106 ( .A(n41912), .B(n41913), .Z(n41915) );
  AND U41107 ( .A(n44169), .B(n44170), .Z(n41913) );
  XOR U41108 ( .A(n41909), .B(n41910), .Z(n41912) );
  AND U41109 ( .A(n44171), .B(n44172), .Z(n41910) );
  XOR U41110 ( .A(n41906), .B(n41907), .Z(n41909) );
  AND U41111 ( .A(n44173), .B(n44174), .Z(n41907) );
  XOR U41112 ( .A(n41903), .B(n41904), .Z(n41906) );
  AND U41113 ( .A(n44175), .B(n44176), .Z(n41904) );
  XOR U41114 ( .A(n41900), .B(n41901), .Z(n41903) );
  AND U41115 ( .A(n44177), .B(n44178), .Z(n41901) );
  XOR U41116 ( .A(n41897), .B(n41898), .Z(n41900) );
  AND U41117 ( .A(n44179), .B(n44180), .Z(n41898) );
  XOR U41118 ( .A(n41894), .B(n41895), .Z(n41897) );
  AND U41119 ( .A(n44181), .B(n44182), .Z(n41895) );
  XOR U41120 ( .A(n41891), .B(n41892), .Z(n41894) );
  AND U41121 ( .A(n44183), .B(n44184), .Z(n41892) );
  XOR U41122 ( .A(n41888), .B(n41889), .Z(n41891) );
  AND U41123 ( .A(n44185), .B(n44186), .Z(n41889) );
  XOR U41124 ( .A(n41885), .B(n41886), .Z(n41888) );
  AND U41125 ( .A(n44187), .B(n44188), .Z(n41886) );
  XOR U41126 ( .A(n41882), .B(n41883), .Z(n41885) );
  AND U41127 ( .A(n44189), .B(n44190), .Z(n41883) );
  XOR U41128 ( .A(n41879), .B(n41880), .Z(n41882) );
  AND U41129 ( .A(n44191), .B(n44192), .Z(n41880) );
  XOR U41130 ( .A(n41876), .B(n41877), .Z(n41879) );
  AND U41131 ( .A(n44193), .B(n44194), .Z(n41877) );
  XOR U41132 ( .A(n41873), .B(n41874), .Z(n41876) );
  AND U41133 ( .A(n44195), .B(n44196), .Z(n41874) );
  XOR U41134 ( .A(n41870), .B(n41871), .Z(n41873) );
  AND U41135 ( .A(n44197), .B(n44198), .Z(n41871) );
  XOR U41136 ( .A(n41867), .B(n41868), .Z(n41870) );
  AND U41137 ( .A(n44199), .B(n44200), .Z(n41868) );
  XOR U41138 ( .A(n41864), .B(n41865), .Z(n41867) );
  AND U41139 ( .A(n44201), .B(n44202), .Z(n41865) );
  XOR U41140 ( .A(n41861), .B(n41862), .Z(n41864) );
  AND U41141 ( .A(n44203), .B(n44204), .Z(n41862) );
  XOR U41142 ( .A(n41858), .B(n41859), .Z(n41861) );
  AND U41143 ( .A(n44205), .B(n44206), .Z(n41859) );
  XOR U41144 ( .A(n41855), .B(n41856), .Z(n41858) );
  AND U41145 ( .A(n44207), .B(n44208), .Z(n41856) );
  XOR U41146 ( .A(n41852), .B(n41853), .Z(n41855) );
  AND U41147 ( .A(n44209), .B(n44210), .Z(n41853) );
  XOR U41148 ( .A(n41849), .B(n41850), .Z(n41852) );
  AND U41149 ( .A(n44211), .B(n44212), .Z(n41850) );
  XOR U41150 ( .A(n41846), .B(n41847), .Z(n41849) );
  AND U41151 ( .A(n44213), .B(n44214), .Z(n41847) );
  XOR U41152 ( .A(n41843), .B(n41844), .Z(n41846) );
  AND U41153 ( .A(n44215), .B(n44216), .Z(n41844) );
  XOR U41154 ( .A(n41840), .B(n41841), .Z(n41843) );
  AND U41155 ( .A(n44217), .B(n44218), .Z(n41841) );
  XOR U41156 ( .A(n41837), .B(n41838), .Z(n41840) );
  AND U41157 ( .A(n44219), .B(n44220), .Z(n41838) );
  XOR U41158 ( .A(n41834), .B(n41835), .Z(n41837) );
  AND U41159 ( .A(n44221), .B(n44222), .Z(n41835) );
  XOR U41160 ( .A(n41831), .B(n41832), .Z(n41834) );
  AND U41161 ( .A(n44223), .B(n44224), .Z(n41832) );
  XOR U41162 ( .A(n41828), .B(n41829), .Z(n41831) );
  AND U41163 ( .A(n44225), .B(n44226), .Z(n41829) );
  XOR U41164 ( .A(n41825), .B(n41826), .Z(n41828) );
  AND U41165 ( .A(n44227), .B(n44228), .Z(n41826) );
  XOR U41166 ( .A(n41822), .B(n41823), .Z(n41825) );
  AND U41167 ( .A(n44229), .B(n44230), .Z(n41823) );
  XOR U41168 ( .A(n41819), .B(n41820), .Z(n41822) );
  AND U41169 ( .A(n44231), .B(n44232), .Z(n41820) );
  XOR U41170 ( .A(n41816), .B(n41817), .Z(n41819) );
  AND U41171 ( .A(n44233), .B(n44234), .Z(n41817) );
  XOR U41172 ( .A(n41813), .B(n41814), .Z(n41816) );
  AND U41173 ( .A(n44235), .B(n44236), .Z(n41814) );
  XOR U41174 ( .A(n41810), .B(n41811), .Z(n41813) );
  AND U41175 ( .A(n44237), .B(n44238), .Z(n41811) );
  XOR U41176 ( .A(n41807), .B(n41808), .Z(n41810) );
  AND U41177 ( .A(n44239), .B(n44240), .Z(n41808) );
  XOR U41178 ( .A(n41804), .B(n41805), .Z(n41807) );
  AND U41179 ( .A(n44241), .B(n44242), .Z(n41805) );
  XOR U41180 ( .A(n41801), .B(n41802), .Z(n41804) );
  AND U41181 ( .A(n44243), .B(n44244), .Z(n41802) );
  XOR U41182 ( .A(n41798), .B(n41799), .Z(n41801) );
  AND U41183 ( .A(n44245), .B(n44246), .Z(n41799) );
  XOR U41184 ( .A(n41795), .B(n41796), .Z(n41798) );
  AND U41185 ( .A(n44247), .B(n44248), .Z(n41796) );
  XOR U41186 ( .A(n41792), .B(n41793), .Z(n41795) );
  AND U41187 ( .A(n44249), .B(n44250), .Z(n41793) );
  XOR U41188 ( .A(n41789), .B(n41790), .Z(n41792) );
  AND U41189 ( .A(n44251), .B(n44252), .Z(n41790) );
  XOR U41190 ( .A(n41786), .B(n41787), .Z(n41789) );
  AND U41191 ( .A(n44253), .B(n44254), .Z(n41787) );
  XOR U41192 ( .A(n41783), .B(n41784), .Z(n41786) );
  AND U41193 ( .A(n44255), .B(n44256), .Z(n41784) );
  XOR U41194 ( .A(n41780), .B(n41781), .Z(n41783) );
  AND U41195 ( .A(n44257), .B(n44258), .Z(n41781) );
  XOR U41196 ( .A(n41777), .B(n41778), .Z(n41780) );
  AND U41197 ( .A(n44259), .B(n44260), .Z(n41778) );
  XOR U41198 ( .A(n41774), .B(n41775), .Z(n41777) );
  AND U41199 ( .A(n44261), .B(n44262), .Z(n41775) );
  XOR U41200 ( .A(n41771), .B(n41772), .Z(n41774) );
  AND U41201 ( .A(n44263), .B(n44264), .Z(n41772) );
  XOR U41202 ( .A(n41768), .B(n41769), .Z(n41771) );
  AND U41203 ( .A(n44265), .B(n44266), .Z(n41769) );
  XOR U41204 ( .A(n41765), .B(n41766), .Z(n41768) );
  AND U41205 ( .A(n44267), .B(n44268), .Z(n41766) );
  XOR U41206 ( .A(n41762), .B(n41763), .Z(n41765) );
  AND U41207 ( .A(n44269), .B(n44270), .Z(n41763) );
  XOR U41208 ( .A(n41759), .B(n41760), .Z(n41762) );
  AND U41209 ( .A(n44271), .B(n44272), .Z(n41760) );
  XOR U41210 ( .A(n41756), .B(n41757), .Z(n41759) );
  AND U41211 ( .A(n44273), .B(n44274), .Z(n41757) );
  XOR U41212 ( .A(n41753), .B(n41754), .Z(n41756) );
  AND U41213 ( .A(n44275), .B(n44276), .Z(n41754) );
  XOR U41214 ( .A(n41750), .B(n41751), .Z(n41753) );
  AND U41215 ( .A(n44277), .B(n44278), .Z(n41751) );
  XOR U41216 ( .A(n41747), .B(n41748), .Z(n41750) );
  AND U41217 ( .A(n44279), .B(n44280), .Z(n41748) );
  XOR U41218 ( .A(n41744), .B(n41745), .Z(n41747) );
  AND U41219 ( .A(n44281), .B(n44282), .Z(n41745) );
  XOR U41220 ( .A(n41741), .B(n41742), .Z(n41744) );
  AND U41221 ( .A(n44283), .B(n44284), .Z(n41742) );
  XOR U41222 ( .A(n41738), .B(n41739), .Z(n41741) );
  AND U41223 ( .A(n44285), .B(n44286), .Z(n41739) );
  XOR U41224 ( .A(n41735), .B(n41736), .Z(n41738) );
  AND U41225 ( .A(n44287), .B(n44288), .Z(n41736) );
  XOR U41226 ( .A(n41732), .B(n41733), .Z(n41735) );
  AND U41227 ( .A(n44289), .B(n44290), .Z(n41733) );
  XOR U41228 ( .A(n41729), .B(n41730), .Z(n41732) );
  AND U41229 ( .A(n44291), .B(n44292), .Z(n41730) );
  XOR U41230 ( .A(n41726), .B(n41727), .Z(n41729) );
  AND U41231 ( .A(n44293), .B(n44294), .Z(n41727) );
  XOR U41232 ( .A(n41723), .B(n41724), .Z(n41726) );
  AND U41233 ( .A(n44295), .B(n44296), .Z(n41724) );
  XOR U41234 ( .A(n41720), .B(n41721), .Z(n41723) );
  AND U41235 ( .A(n44297), .B(n44298), .Z(n41721) );
  XOR U41236 ( .A(n41717), .B(n41718), .Z(n41720) );
  AND U41237 ( .A(n44299), .B(n44300), .Z(n41718) );
  XOR U41238 ( .A(n41714), .B(n41715), .Z(n41717) );
  AND U41239 ( .A(n44301), .B(n44302), .Z(n41715) );
  XOR U41240 ( .A(n41711), .B(n41712), .Z(n41714) );
  AND U41241 ( .A(n44303), .B(n44304), .Z(n41712) );
  XOR U41242 ( .A(n41708), .B(n41709), .Z(n41711) );
  AND U41243 ( .A(n44305), .B(n44306), .Z(n41709) );
  XOR U41244 ( .A(n41705), .B(n41706), .Z(n41708) );
  AND U41245 ( .A(n44307), .B(n44308), .Z(n41706) );
  XOR U41246 ( .A(n41702), .B(n41703), .Z(n41705) );
  AND U41247 ( .A(n44309), .B(n44310), .Z(n41703) );
  XOR U41248 ( .A(n41699), .B(n41700), .Z(n41702) );
  AND U41249 ( .A(n44311), .B(n44312), .Z(n41700) );
  XOR U41250 ( .A(n41696), .B(n41697), .Z(n41699) );
  AND U41251 ( .A(n44313), .B(n44314), .Z(n41697) );
  XOR U41252 ( .A(n41693), .B(n41694), .Z(n41696) );
  AND U41253 ( .A(n44315), .B(n44316), .Z(n41694) );
  XOR U41254 ( .A(n41690), .B(n41691), .Z(n41693) );
  AND U41255 ( .A(n44317), .B(n44318), .Z(n41691) );
  XOR U41256 ( .A(n41687), .B(n41688), .Z(n41690) );
  AND U41257 ( .A(n44319), .B(n44320), .Z(n41688) );
  XOR U41258 ( .A(n41684), .B(n41685), .Z(n41687) );
  AND U41259 ( .A(n44321), .B(n44322), .Z(n41685) );
  XOR U41260 ( .A(n41681), .B(n41682), .Z(n41684) );
  AND U41261 ( .A(n44323), .B(n44324), .Z(n41682) );
  XOR U41262 ( .A(n41678), .B(n41679), .Z(n41681) );
  AND U41263 ( .A(n44325), .B(n44326), .Z(n41679) );
  XOR U41264 ( .A(n41675), .B(n41676), .Z(n41678) );
  AND U41265 ( .A(n44327), .B(n44328), .Z(n41676) );
  XOR U41266 ( .A(n41672), .B(n41673), .Z(n41675) );
  AND U41267 ( .A(n44329), .B(n44330), .Z(n41673) );
  XOR U41268 ( .A(n41669), .B(n41670), .Z(n41672) );
  AND U41269 ( .A(n44331), .B(n44332), .Z(n41670) );
  XOR U41270 ( .A(n41666), .B(n41667), .Z(n41669) );
  AND U41271 ( .A(n44333), .B(n44334), .Z(n41667) );
  XOR U41272 ( .A(n41663), .B(n41664), .Z(n41666) );
  AND U41273 ( .A(n44335), .B(n44336), .Z(n41664) );
  XOR U41274 ( .A(n41660), .B(n41661), .Z(n41663) );
  AND U41275 ( .A(n44337), .B(n44338), .Z(n41661) );
  XOR U41276 ( .A(n41657), .B(n41658), .Z(n41660) );
  AND U41277 ( .A(n44339), .B(n44340), .Z(n41658) );
  XOR U41278 ( .A(n41654), .B(n41655), .Z(n41657) );
  AND U41279 ( .A(n44341), .B(n44342), .Z(n41655) );
  XOR U41280 ( .A(n41651), .B(n41652), .Z(n41654) );
  AND U41281 ( .A(n44343), .B(n44344), .Z(n41652) );
  XOR U41282 ( .A(n41648), .B(n41649), .Z(n41651) );
  AND U41283 ( .A(n44345), .B(n44346), .Z(n41649) );
  XOR U41284 ( .A(n41645), .B(n41646), .Z(n41648) );
  AND U41285 ( .A(n44347), .B(n44348), .Z(n41646) );
  XOR U41286 ( .A(n41642), .B(n41643), .Z(n41645) );
  AND U41287 ( .A(n44349), .B(n44350), .Z(n41643) );
  XOR U41288 ( .A(n41639), .B(n41640), .Z(n41642) );
  AND U41289 ( .A(n44351), .B(n44352), .Z(n41640) );
  XOR U41290 ( .A(n41636), .B(n41637), .Z(n41639) );
  AND U41291 ( .A(n44353), .B(n44354), .Z(n41637) );
  XOR U41292 ( .A(n41633), .B(n41634), .Z(n41636) );
  AND U41293 ( .A(n44355), .B(n44356), .Z(n41634) );
  XOR U41294 ( .A(n41630), .B(n41631), .Z(n41633) );
  AND U41295 ( .A(n44357), .B(n44358), .Z(n41631) );
  XOR U41296 ( .A(n41627), .B(n41628), .Z(n41630) );
  AND U41297 ( .A(n44359), .B(n44360), .Z(n41628) );
  XOR U41298 ( .A(n41624), .B(n41625), .Z(n41627) );
  AND U41299 ( .A(n44361), .B(n44362), .Z(n41625) );
  XOR U41300 ( .A(n41621), .B(n41622), .Z(n41624) );
  AND U41301 ( .A(n44363), .B(n44364), .Z(n41622) );
  XOR U41302 ( .A(n41618), .B(n41619), .Z(n41621) );
  AND U41303 ( .A(n44365), .B(n44366), .Z(n41619) );
  XOR U41304 ( .A(n41615), .B(n41616), .Z(n41618) );
  AND U41305 ( .A(n44367), .B(n44368), .Z(n41616) );
  XOR U41306 ( .A(n41612), .B(n41613), .Z(n41615) );
  AND U41307 ( .A(n44369), .B(n44370), .Z(n41613) );
  XOR U41308 ( .A(n41609), .B(n41610), .Z(n41612) );
  AND U41309 ( .A(n44371), .B(n44372), .Z(n41610) );
  XOR U41310 ( .A(n41606), .B(n41607), .Z(n41609) );
  AND U41311 ( .A(n44373), .B(n44374), .Z(n41607) );
  XOR U41312 ( .A(n41603), .B(n41604), .Z(n41606) );
  AND U41313 ( .A(n44375), .B(n44376), .Z(n41604) );
  XOR U41314 ( .A(n41600), .B(n41601), .Z(n41603) );
  AND U41315 ( .A(n44377), .B(n44378), .Z(n41601) );
  XOR U41316 ( .A(n41597), .B(n41598), .Z(n41600) );
  AND U41317 ( .A(n44379), .B(n44380), .Z(n41598) );
  XOR U41318 ( .A(n41594), .B(n41595), .Z(n41597) );
  AND U41319 ( .A(n44381), .B(n44382), .Z(n41595) );
  XOR U41320 ( .A(n41591), .B(n41592), .Z(n41594) );
  AND U41321 ( .A(n44383), .B(n44384), .Z(n41592) );
  XOR U41322 ( .A(n41588), .B(n41589), .Z(n41591) );
  AND U41323 ( .A(n44385), .B(n44386), .Z(n41589) );
  XOR U41324 ( .A(n41585), .B(n41586), .Z(n41588) );
  AND U41325 ( .A(n44387), .B(n44388), .Z(n41586) );
  XOR U41326 ( .A(n41582), .B(n41583), .Z(n41585) );
  AND U41327 ( .A(n44389), .B(n44390), .Z(n41583) );
  XOR U41328 ( .A(n41579), .B(n41580), .Z(n41582) );
  AND U41329 ( .A(n44391), .B(n44392), .Z(n41580) );
  XOR U41330 ( .A(n41576), .B(n41577), .Z(n41579) );
  AND U41331 ( .A(n44393), .B(n44394), .Z(n41577) );
  XOR U41332 ( .A(n41573), .B(n41574), .Z(n41576) );
  AND U41333 ( .A(n44395), .B(n44396), .Z(n41574) );
  XOR U41334 ( .A(n41570), .B(n41571), .Z(n41573) );
  AND U41335 ( .A(n44397), .B(n44398), .Z(n41571) );
  XOR U41336 ( .A(n41567), .B(n41568), .Z(n41570) );
  AND U41337 ( .A(n44399), .B(n44400), .Z(n41568) );
  XOR U41338 ( .A(n41564), .B(n41565), .Z(n41567) );
  AND U41339 ( .A(n44401), .B(n44402), .Z(n41565) );
  XOR U41340 ( .A(n41561), .B(n41562), .Z(n41564) );
  AND U41341 ( .A(n44403), .B(n44404), .Z(n41562) );
  XOR U41342 ( .A(n41558), .B(n41559), .Z(n41561) );
  AND U41343 ( .A(n44405), .B(n44406), .Z(n41559) );
  XOR U41344 ( .A(n41555), .B(n41556), .Z(n41558) );
  AND U41345 ( .A(n44407), .B(n44408), .Z(n41556) );
  XOR U41346 ( .A(n41552), .B(n41553), .Z(n41555) );
  AND U41347 ( .A(n44409), .B(n44410), .Z(n41553) );
  XOR U41348 ( .A(n41549), .B(n41550), .Z(n41552) );
  AND U41349 ( .A(n44411), .B(n44412), .Z(n41550) );
  XOR U41350 ( .A(n41546), .B(n41547), .Z(n41549) );
  AND U41351 ( .A(n44413), .B(n44414), .Z(n41547) );
  XOR U41352 ( .A(n41543), .B(n41544), .Z(n41546) );
  AND U41353 ( .A(n44415), .B(n44416), .Z(n41544) );
  XOR U41354 ( .A(n41540), .B(n41541), .Z(n41543) );
  AND U41355 ( .A(n44417), .B(n44418), .Z(n41541) );
  XOR U41356 ( .A(n41537), .B(n41538), .Z(n41540) );
  AND U41357 ( .A(n44419), .B(n44420), .Z(n41538) );
  XOR U41358 ( .A(n41534), .B(n41535), .Z(n41537) );
  AND U41359 ( .A(n44421), .B(n44422), .Z(n41535) );
  XOR U41360 ( .A(n41531), .B(n41532), .Z(n41534) );
  AND U41361 ( .A(n44423), .B(n44424), .Z(n41532) );
  XOR U41362 ( .A(n41528), .B(n41529), .Z(n41531) );
  AND U41363 ( .A(n44425), .B(n44426), .Z(n41529) );
  XOR U41364 ( .A(n41525), .B(n41526), .Z(n41528) );
  AND U41365 ( .A(n44427), .B(n44428), .Z(n41526) );
  XOR U41366 ( .A(n41522), .B(n41523), .Z(n41525) );
  AND U41367 ( .A(n44429), .B(n44430), .Z(n41523) );
  XOR U41368 ( .A(n41519), .B(n41520), .Z(n41522) );
  AND U41369 ( .A(n44431), .B(n44432), .Z(n41520) );
  XOR U41370 ( .A(n41516), .B(n41517), .Z(n41519) );
  AND U41371 ( .A(n44433), .B(n44434), .Z(n41517) );
  XOR U41372 ( .A(n41513), .B(n41514), .Z(n41516) );
  AND U41373 ( .A(n44435), .B(n44436), .Z(n41514) );
  XOR U41374 ( .A(n41510), .B(n41511), .Z(n41513) );
  AND U41375 ( .A(n44437), .B(n44438), .Z(n41511) );
  XOR U41376 ( .A(n41507), .B(n41508), .Z(n41510) );
  AND U41377 ( .A(n44439), .B(n44440), .Z(n41508) );
  XOR U41378 ( .A(n41504), .B(n41505), .Z(n41507) );
  AND U41379 ( .A(n44441), .B(n44442), .Z(n41505) );
  XOR U41380 ( .A(n41501), .B(n41502), .Z(n41504) );
  AND U41381 ( .A(n44443), .B(n44444), .Z(n41502) );
  XOR U41382 ( .A(n41498), .B(n41499), .Z(n41501) );
  AND U41383 ( .A(n44445), .B(n44446), .Z(n41499) );
  XOR U41384 ( .A(n41495), .B(n41496), .Z(n41498) );
  AND U41385 ( .A(n44447), .B(n44448), .Z(n41496) );
  XNOR U41386 ( .A(n41492), .B(n41493), .Z(n41495) );
  AND U41387 ( .A(n44449), .B(n44450), .Z(n41493) );
  XOR U41388 ( .A(n44451), .B(n41490), .Z(n41492) );
  IV U41389 ( .A(n44452), .Z(n41490) );
  AND U41390 ( .A(n44453), .B(n44454), .Z(n44452) );
  IV U41391 ( .A(n41489), .Z(n44451) );
  XOR U41392 ( .A(n41230), .B(n41486), .Z(n41489) );
  AND U41393 ( .A(n44455), .B(n44456), .Z(n41486) );
  XOR U41394 ( .A(n41232), .B(n41231), .Z(n41230) );
  AND U41395 ( .A(n44457), .B(n44458), .Z(n41231) );
  XOR U41396 ( .A(n41234), .B(n41233), .Z(n41232) );
  AND U41397 ( .A(n44459), .B(n44460), .Z(n41233) );
  XOR U41398 ( .A(n41236), .B(n41235), .Z(n41234) );
  AND U41399 ( .A(n44461), .B(n44462), .Z(n41235) );
  XOR U41400 ( .A(n41238), .B(n41237), .Z(n41236) );
  AND U41401 ( .A(n44463), .B(n44464), .Z(n41237) );
  XOR U41402 ( .A(n41240), .B(n41239), .Z(n41238) );
  AND U41403 ( .A(n44465), .B(n44466), .Z(n41239) );
  XOR U41404 ( .A(n41242), .B(n41241), .Z(n41240) );
  AND U41405 ( .A(n44467), .B(n44468), .Z(n41241) );
  XOR U41406 ( .A(n41244), .B(n41243), .Z(n41242) );
  AND U41407 ( .A(n44469), .B(n44470), .Z(n41243) );
  XOR U41408 ( .A(n41246), .B(n41245), .Z(n41244) );
  AND U41409 ( .A(n44471), .B(n44472), .Z(n41245) );
  XOR U41410 ( .A(n41248), .B(n41247), .Z(n41246) );
  AND U41411 ( .A(n44473), .B(n44474), .Z(n41247) );
  XOR U41412 ( .A(n41250), .B(n41249), .Z(n41248) );
  AND U41413 ( .A(n44475), .B(n44476), .Z(n41249) );
  XOR U41414 ( .A(n41252), .B(n41251), .Z(n41250) );
  AND U41415 ( .A(n44477), .B(n44478), .Z(n41251) );
  XOR U41416 ( .A(n41254), .B(n41253), .Z(n41252) );
  AND U41417 ( .A(n44479), .B(n44480), .Z(n41253) );
  XOR U41418 ( .A(n41256), .B(n41255), .Z(n41254) );
  AND U41419 ( .A(n44481), .B(n44482), .Z(n41255) );
  XOR U41420 ( .A(n41258), .B(n41257), .Z(n41256) );
  AND U41421 ( .A(n44483), .B(n44484), .Z(n41257) );
  XOR U41422 ( .A(n41260), .B(n41259), .Z(n41258) );
  AND U41423 ( .A(n44485), .B(n44486), .Z(n41259) );
  XOR U41424 ( .A(n41262), .B(n41261), .Z(n41260) );
  AND U41425 ( .A(n44487), .B(n44488), .Z(n41261) );
  XOR U41426 ( .A(n41264), .B(n41263), .Z(n41262) );
  AND U41427 ( .A(n44489), .B(n44490), .Z(n41263) );
  XOR U41428 ( .A(n41266), .B(n41265), .Z(n41264) );
  AND U41429 ( .A(n44491), .B(n44492), .Z(n41265) );
  XOR U41430 ( .A(n41268), .B(n41267), .Z(n41266) );
  AND U41431 ( .A(n44493), .B(n44494), .Z(n41267) );
  XOR U41432 ( .A(n41270), .B(n41269), .Z(n41268) );
  AND U41433 ( .A(n44495), .B(n44496), .Z(n41269) );
  XOR U41434 ( .A(n41272), .B(n41271), .Z(n41270) );
  AND U41435 ( .A(n44497), .B(n44498), .Z(n41271) );
  XOR U41436 ( .A(n41274), .B(n41273), .Z(n41272) );
  AND U41437 ( .A(n44499), .B(n44500), .Z(n41273) );
  XOR U41438 ( .A(n41276), .B(n41275), .Z(n41274) );
  AND U41439 ( .A(n44501), .B(n44502), .Z(n41275) );
  XOR U41440 ( .A(n41278), .B(n41277), .Z(n41276) );
  AND U41441 ( .A(n44503), .B(n44504), .Z(n41277) );
  XOR U41442 ( .A(n41280), .B(n41279), .Z(n41278) );
  AND U41443 ( .A(n44505), .B(n44506), .Z(n41279) );
  XOR U41444 ( .A(n41282), .B(n41281), .Z(n41280) );
  AND U41445 ( .A(n44507), .B(n44508), .Z(n41281) );
  XOR U41446 ( .A(n41284), .B(n41283), .Z(n41282) );
  AND U41447 ( .A(n44509), .B(n44510), .Z(n41283) );
  XOR U41448 ( .A(n41286), .B(n41285), .Z(n41284) );
  AND U41449 ( .A(n44511), .B(n44512), .Z(n41285) );
  XOR U41450 ( .A(n41288), .B(n41287), .Z(n41286) );
  AND U41451 ( .A(n44513), .B(n44514), .Z(n41287) );
  XOR U41452 ( .A(n41290), .B(n41289), .Z(n41288) );
  AND U41453 ( .A(n44515), .B(n44516), .Z(n41289) );
  XOR U41454 ( .A(n41292), .B(n41291), .Z(n41290) );
  AND U41455 ( .A(n44517), .B(n44518), .Z(n41291) );
  XOR U41456 ( .A(n41294), .B(n41293), .Z(n41292) );
  AND U41457 ( .A(n44519), .B(n44520), .Z(n41293) );
  XOR U41458 ( .A(n41296), .B(n41295), .Z(n41294) );
  AND U41459 ( .A(n44521), .B(n44522), .Z(n41295) );
  XOR U41460 ( .A(n41298), .B(n41297), .Z(n41296) );
  AND U41461 ( .A(n44523), .B(n44524), .Z(n41297) );
  XOR U41462 ( .A(n41300), .B(n41299), .Z(n41298) );
  AND U41463 ( .A(n44525), .B(n44526), .Z(n41299) );
  XOR U41464 ( .A(n41302), .B(n41301), .Z(n41300) );
  AND U41465 ( .A(n44527), .B(n44528), .Z(n41301) );
  XOR U41466 ( .A(n41304), .B(n41303), .Z(n41302) );
  AND U41467 ( .A(n44529), .B(n44530), .Z(n41303) );
  XOR U41468 ( .A(n41306), .B(n41305), .Z(n41304) );
  AND U41469 ( .A(n44531), .B(n44532), .Z(n41305) );
  XOR U41470 ( .A(n41308), .B(n41307), .Z(n41306) );
  AND U41471 ( .A(n44533), .B(n44534), .Z(n41307) );
  XOR U41472 ( .A(n41310), .B(n41309), .Z(n41308) );
  AND U41473 ( .A(n44535), .B(n44536), .Z(n41309) );
  XOR U41474 ( .A(n41312), .B(n41311), .Z(n41310) );
  AND U41475 ( .A(n44537), .B(n44538), .Z(n41311) );
  XOR U41476 ( .A(n41314), .B(n41313), .Z(n41312) );
  AND U41477 ( .A(n44539), .B(n44540), .Z(n41313) );
  XOR U41478 ( .A(n41316), .B(n41315), .Z(n41314) );
  AND U41479 ( .A(n44541), .B(n44542), .Z(n41315) );
  XOR U41480 ( .A(n41318), .B(n41317), .Z(n41316) );
  AND U41481 ( .A(n44543), .B(n44544), .Z(n41317) );
  XOR U41482 ( .A(n41320), .B(n41319), .Z(n41318) );
  AND U41483 ( .A(n44545), .B(n44546), .Z(n41319) );
  XOR U41484 ( .A(n41322), .B(n41321), .Z(n41320) );
  AND U41485 ( .A(n44547), .B(n44548), .Z(n41321) );
  XOR U41486 ( .A(n41324), .B(n41323), .Z(n41322) );
  AND U41487 ( .A(n44549), .B(n44550), .Z(n41323) );
  XOR U41488 ( .A(n41326), .B(n41325), .Z(n41324) );
  AND U41489 ( .A(n44551), .B(n44552), .Z(n41325) );
  XOR U41490 ( .A(n41328), .B(n41327), .Z(n41326) );
  AND U41491 ( .A(n44553), .B(n44554), .Z(n41327) );
  XOR U41492 ( .A(n41330), .B(n41329), .Z(n41328) );
  AND U41493 ( .A(n44555), .B(n44556), .Z(n41329) );
  XOR U41494 ( .A(n41332), .B(n41331), .Z(n41330) );
  AND U41495 ( .A(n44557), .B(n44558), .Z(n41331) );
  XOR U41496 ( .A(n41334), .B(n41333), .Z(n41332) );
  AND U41497 ( .A(n44559), .B(n44560), .Z(n41333) );
  XOR U41498 ( .A(n41336), .B(n41335), .Z(n41334) );
  AND U41499 ( .A(n44561), .B(n44562), .Z(n41335) );
  XOR U41500 ( .A(n41338), .B(n41337), .Z(n41336) );
  AND U41501 ( .A(n44563), .B(n44564), .Z(n41337) );
  XOR U41502 ( .A(n41340), .B(n41339), .Z(n41338) );
  AND U41503 ( .A(n44565), .B(n44566), .Z(n41339) );
  XOR U41504 ( .A(n41342), .B(n41341), .Z(n41340) );
  AND U41505 ( .A(n44567), .B(n44568), .Z(n41341) );
  XOR U41506 ( .A(n41344), .B(n41343), .Z(n41342) );
  AND U41507 ( .A(n44569), .B(n44570), .Z(n41343) );
  XOR U41508 ( .A(n41346), .B(n41345), .Z(n41344) );
  AND U41509 ( .A(n44571), .B(n44572), .Z(n41345) );
  XOR U41510 ( .A(n41348), .B(n41347), .Z(n41346) );
  AND U41511 ( .A(n44573), .B(n44574), .Z(n41347) );
  XOR U41512 ( .A(n41350), .B(n41349), .Z(n41348) );
  AND U41513 ( .A(n44575), .B(n44576), .Z(n41349) );
  XOR U41514 ( .A(n41352), .B(n41351), .Z(n41350) );
  AND U41515 ( .A(n44577), .B(n44578), .Z(n41351) );
  XOR U41516 ( .A(n41354), .B(n41353), .Z(n41352) );
  AND U41517 ( .A(n44579), .B(n44580), .Z(n41353) );
  XOR U41518 ( .A(n41356), .B(n41355), .Z(n41354) );
  AND U41519 ( .A(n44581), .B(n44582), .Z(n41355) );
  XOR U41520 ( .A(n41358), .B(n41357), .Z(n41356) );
  AND U41521 ( .A(n44583), .B(n44584), .Z(n41357) );
  XOR U41522 ( .A(n41360), .B(n41359), .Z(n41358) );
  AND U41523 ( .A(n44585), .B(n44586), .Z(n41359) );
  XOR U41524 ( .A(n41362), .B(n41361), .Z(n41360) );
  AND U41525 ( .A(n44587), .B(n44588), .Z(n41361) );
  XOR U41526 ( .A(n41364), .B(n41363), .Z(n41362) );
  AND U41527 ( .A(n44589), .B(n44590), .Z(n41363) );
  XOR U41528 ( .A(n41366), .B(n41365), .Z(n41364) );
  AND U41529 ( .A(n44591), .B(n44592), .Z(n41365) );
  XOR U41530 ( .A(n41368), .B(n41367), .Z(n41366) );
  AND U41531 ( .A(n44593), .B(n44594), .Z(n41367) );
  XOR U41532 ( .A(n41370), .B(n41369), .Z(n41368) );
  AND U41533 ( .A(n44595), .B(n44596), .Z(n41369) );
  XOR U41534 ( .A(n41372), .B(n41371), .Z(n41370) );
  AND U41535 ( .A(n44597), .B(n44598), .Z(n41371) );
  XOR U41536 ( .A(n41374), .B(n41373), .Z(n41372) );
  AND U41537 ( .A(n44599), .B(n44600), .Z(n41373) );
  XOR U41538 ( .A(n41376), .B(n41375), .Z(n41374) );
  AND U41539 ( .A(n44601), .B(n44602), .Z(n41375) );
  XOR U41540 ( .A(n41378), .B(n41377), .Z(n41376) );
  AND U41541 ( .A(n44603), .B(n44604), .Z(n41377) );
  XOR U41542 ( .A(n41380), .B(n41379), .Z(n41378) );
  AND U41543 ( .A(n44605), .B(n44606), .Z(n41379) );
  XOR U41544 ( .A(n41382), .B(n41381), .Z(n41380) );
  AND U41545 ( .A(n44607), .B(n44608), .Z(n41381) );
  XOR U41546 ( .A(n41384), .B(n41383), .Z(n41382) );
  AND U41547 ( .A(n44609), .B(n44610), .Z(n41383) );
  XOR U41548 ( .A(n41386), .B(n41385), .Z(n41384) );
  AND U41549 ( .A(n44611), .B(n44612), .Z(n41385) );
  XOR U41550 ( .A(n41388), .B(n41387), .Z(n41386) );
  AND U41551 ( .A(n44613), .B(n44614), .Z(n41387) );
  XOR U41552 ( .A(n41390), .B(n41389), .Z(n41388) );
  AND U41553 ( .A(n44615), .B(n44616), .Z(n41389) );
  XOR U41554 ( .A(n41392), .B(n41391), .Z(n41390) );
  AND U41555 ( .A(n44617), .B(n44618), .Z(n41391) );
  XOR U41556 ( .A(n41394), .B(n41393), .Z(n41392) );
  AND U41557 ( .A(n44619), .B(n44620), .Z(n41393) );
  XOR U41558 ( .A(n41396), .B(n41395), .Z(n41394) );
  AND U41559 ( .A(n44621), .B(n44622), .Z(n41395) );
  XOR U41560 ( .A(n41398), .B(n41397), .Z(n41396) );
  AND U41561 ( .A(n44623), .B(n44624), .Z(n41397) );
  XOR U41562 ( .A(n41400), .B(n41399), .Z(n41398) );
  AND U41563 ( .A(n44625), .B(n44626), .Z(n41399) );
  XOR U41564 ( .A(n41402), .B(n41401), .Z(n41400) );
  AND U41565 ( .A(n44627), .B(n44628), .Z(n41401) );
  XOR U41566 ( .A(n41404), .B(n41403), .Z(n41402) );
  AND U41567 ( .A(n44629), .B(n44630), .Z(n41403) );
  XOR U41568 ( .A(n41406), .B(n41405), .Z(n41404) );
  AND U41569 ( .A(n44631), .B(n44632), .Z(n41405) );
  XOR U41570 ( .A(n41408), .B(n41407), .Z(n41406) );
  AND U41571 ( .A(n44633), .B(n44634), .Z(n41407) );
  XOR U41572 ( .A(n41410), .B(n41409), .Z(n41408) );
  AND U41573 ( .A(n44635), .B(n44636), .Z(n41409) );
  XOR U41574 ( .A(n41412), .B(n41411), .Z(n41410) );
  AND U41575 ( .A(n44637), .B(n44638), .Z(n41411) );
  XOR U41576 ( .A(n41414), .B(n41413), .Z(n41412) );
  AND U41577 ( .A(n44639), .B(n44640), .Z(n41413) );
  XOR U41578 ( .A(n41416), .B(n41415), .Z(n41414) );
  AND U41579 ( .A(n44641), .B(n44642), .Z(n41415) );
  XOR U41580 ( .A(n41418), .B(n41417), .Z(n41416) );
  AND U41581 ( .A(n44643), .B(n44644), .Z(n41417) );
  XOR U41582 ( .A(n41420), .B(n41419), .Z(n41418) );
  AND U41583 ( .A(n44645), .B(n44646), .Z(n41419) );
  XOR U41584 ( .A(n41422), .B(n41421), .Z(n41420) );
  AND U41585 ( .A(n44647), .B(n44648), .Z(n41421) );
  XOR U41586 ( .A(n41424), .B(n41423), .Z(n41422) );
  AND U41587 ( .A(n44649), .B(n44650), .Z(n41423) );
  XOR U41588 ( .A(n41426), .B(n41425), .Z(n41424) );
  AND U41589 ( .A(n44651), .B(n44652), .Z(n41425) );
  XOR U41590 ( .A(n41428), .B(n41427), .Z(n41426) );
  AND U41591 ( .A(n44653), .B(n44654), .Z(n41427) );
  XOR U41592 ( .A(n41430), .B(n41429), .Z(n41428) );
  AND U41593 ( .A(n44655), .B(n44656), .Z(n41429) );
  XOR U41594 ( .A(n41432), .B(n41431), .Z(n41430) );
  AND U41595 ( .A(n44657), .B(n44658), .Z(n41431) );
  XOR U41596 ( .A(n41434), .B(n41433), .Z(n41432) );
  AND U41597 ( .A(n44659), .B(n44660), .Z(n41433) );
  XOR U41598 ( .A(n41436), .B(n41435), .Z(n41434) );
  AND U41599 ( .A(n44661), .B(n44662), .Z(n41435) );
  XOR U41600 ( .A(n41438), .B(n41437), .Z(n41436) );
  AND U41601 ( .A(n44663), .B(n44664), .Z(n41437) );
  XOR U41602 ( .A(n41440), .B(n41439), .Z(n41438) );
  AND U41603 ( .A(n44665), .B(n44666), .Z(n41439) );
  XOR U41604 ( .A(n41442), .B(n41441), .Z(n41440) );
  AND U41605 ( .A(n44667), .B(n44668), .Z(n41441) );
  XOR U41606 ( .A(n41444), .B(n41443), .Z(n41442) );
  AND U41607 ( .A(n44669), .B(n44670), .Z(n41443) );
  XOR U41608 ( .A(n41446), .B(n41445), .Z(n41444) );
  AND U41609 ( .A(n44671), .B(n44672), .Z(n41445) );
  XOR U41610 ( .A(n41448), .B(n41447), .Z(n41446) );
  AND U41611 ( .A(n44673), .B(n44674), .Z(n41447) );
  XOR U41612 ( .A(n41450), .B(n41449), .Z(n41448) );
  AND U41613 ( .A(n44675), .B(n44676), .Z(n41449) );
  XOR U41614 ( .A(n41452), .B(n41451), .Z(n41450) );
  AND U41615 ( .A(n44677), .B(n44678), .Z(n41451) );
  XOR U41616 ( .A(n41454), .B(n41453), .Z(n41452) );
  AND U41617 ( .A(n44679), .B(n44680), .Z(n41453) );
  XOR U41618 ( .A(n41482), .B(n41455), .Z(n41454) );
  AND U41619 ( .A(n44681), .B(n44682), .Z(n41455) );
  XOR U41620 ( .A(n41484), .B(n41483), .Z(n41482) );
  AND U41621 ( .A(n44683), .B(n44684), .Z(n41483) );
  XOR U41622 ( .A(n41463), .B(n41485), .Z(n41484) );
  AND U41623 ( .A(n44685), .B(n44686), .Z(n41485) );
  XOR U41624 ( .A(n41459), .B(n41464), .Z(n41463) );
  AND U41625 ( .A(n44687), .B(n44688), .Z(n41464) );
  XOR U41626 ( .A(n41461), .B(n41460), .Z(n41459) );
  AND U41627 ( .A(n44689), .B(n44690), .Z(n41460) );
  XNOR U41628 ( .A(n41471), .B(n41462), .Z(n41461) );
  AND U41629 ( .A(n44691), .B(n44692), .Z(n41462) );
  XOR U41630 ( .A(n41481), .B(n41470), .Z(n41471) );
  AND U41631 ( .A(n44693), .B(n44694), .Z(n41470) );
  XNOR U41632 ( .A(n44695), .B(n41476), .Z(n41481) );
  XOR U41633 ( .A(n41477), .B(n44696), .Z(n41476) );
  AND U41634 ( .A(n44697), .B(n44698), .Z(n44696) );
  XOR U41635 ( .A(n44699), .B(n44700), .Z(n41477) );
  NOR U41636 ( .A(n44701), .B(n44702), .Z(n44700) );
  AND U41637 ( .A(n44703), .B(n44704), .Z(n44702) );
  AND U41638 ( .A(n44705), .B(n44706), .Z(n44701) );
  XNOR U41639 ( .A(n44703), .B(n44704), .Z(n44699) );
  XNOR U41640 ( .A(n41468), .B(n41480), .Z(n44695) );
  AND U41641 ( .A(n44707), .B(n44708), .Z(n41480) );
  AND U41642 ( .A(n44709), .B(n44710), .Z(n41468) );
  NOR U41643 ( .A(n22942), .B(n22945), .Z(n42647) );
  XNOR U41644 ( .A(n42652), .B(n42651), .Z(n22945) );
  NOR U41645 ( .A(n21919), .B(p_input[1023]), .Z(n42651) );
  XOR U41646 ( .A(n42654), .B(n42653), .Z(n42652) );
  NOR U41647 ( .A(n21921), .B(p_input[1021]), .Z(n42653) );
  XOR U41648 ( .A(n42656), .B(n42655), .Z(n42654) );
  NOR U41649 ( .A(n21923), .B(p_input[1019]), .Z(n42655) );
  XOR U41650 ( .A(n42658), .B(n42657), .Z(n42656) );
  NOR U41651 ( .A(n21925), .B(p_input[1017]), .Z(n42657) );
  XOR U41652 ( .A(n42660), .B(n42659), .Z(n42658) );
  NOR U41653 ( .A(n21927), .B(p_input[1015]), .Z(n42659) );
  XOR U41654 ( .A(n42662), .B(n42661), .Z(n42660) );
  NOR U41655 ( .A(n21929), .B(p_input[1013]), .Z(n42661) );
  XOR U41656 ( .A(n42664), .B(n42663), .Z(n42662) );
  NOR U41657 ( .A(n21931), .B(p_input[1011]), .Z(n42663) );
  XOR U41658 ( .A(n42666), .B(n42665), .Z(n42664) );
  NOR U41659 ( .A(n21933), .B(p_input[1009]), .Z(n42665) );
  XOR U41660 ( .A(n42668), .B(n42667), .Z(n42666) );
  NOR U41661 ( .A(n21935), .B(p_input[1007]), .Z(n42667) );
  XOR U41662 ( .A(n42670), .B(n42669), .Z(n42668) );
  NOR U41663 ( .A(n21937), .B(p_input[1005]), .Z(n42669) );
  XOR U41664 ( .A(n42672), .B(n42671), .Z(n42670) );
  NOR U41665 ( .A(n21939), .B(p_input[1003]), .Z(n42671) );
  XOR U41666 ( .A(n42674), .B(n42673), .Z(n42672) );
  NOR U41667 ( .A(n21941), .B(p_input[1001]), .Z(n42673) );
  XOR U41668 ( .A(n42676), .B(n42675), .Z(n42674) );
  NOR U41669 ( .A(n21943), .B(p_input[999]), .Z(n42675) );
  XOR U41670 ( .A(n42678), .B(n42677), .Z(n42676) );
  NOR U41671 ( .A(n21945), .B(p_input[997]), .Z(n42677) );
  XOR U41672 ( .A(n42680), .B(n42679), .Z(n42678) );
  NOR U41673 ( .A(n21947), .B(p_input[995]), .Z(n42679) );
  XOR U41674 ( .A(n42682), .B(n42681), .Z(n42680) );
  NOR U41675 ( .A(n21949), .B(p_input[993]), .Z(n42681) );
  XOR U41676 ( .A(n42684), .B(n42683), .Z(n42682) );
  NOR U41677 ( .A(n21951), .B(p_input[991]), .Z(n42683) );
  XOR U41678 ( .A(n42686), .B(n42685), .Z(n42684) );
  NOR U41679 ( .A(n21953), .B(p_input[989]), .Z(n42685) );
  XOR U41680 ( .A(n42688), .B(n42687), .Z(n42686) );
  NOR U41681 ( .A(n21955), .B(p_input[987]), .Z(n42687) );
  XOR U41682 ( .A(n42690), .B(n42689), .Z(n42688) );
  NOR U41683 ( .A(n21957), .B(p_input[985]), .Z(n42689) );
  XOR U41684 ( .A(n42692), .B(n42691), .Z(n42690) );
  NOR U41685 ( .A(n21959), .B(p_input[983]), .Z(n42691) );
  XOR U41686 ( .A(n42694), .B(n42693), .Z(n42692) );
  NOR U41687 ( .A(n21961), .B(p_input[981]), .Z(n42693) );
  XOR U41688 ( .A(n42696), .B(n42695), .Z(n42694) );
  NOR U41689 ( .A(n21963), .B(p_input[979]), .Z(n42695) );
  XOR U41690 ( .A(n42698), .B(n42697), .Z(n42696) );
  NOR U41691 ( .A(n21965), .B(p_input[977]), .Z(n42697) );
  XOR U41692 ( .A(n42700), .B(n42699), .Z(n42698) );
  NOR U41693 ( .A(n21967), .B(p_input[975]), .Z(n42699) );
  XOR U41694 ( .A(n42702), .B(n42701), .Z(n42700) );
  NOR U41695 ( .A(n21969), .B(p_input[973]), .Z(n42701) );
  XOR U41696 ( .A(n42704), .B(n42703), .Z(n42702) );
  NOR U41697 ( .A(n21971), .B(p_input[971]), .Z(n42703) );
  XOR U41698 ( .A(n42706), .B(n42705), .Z(n42704) );
  NOR U41699 ( .A(n21973), .B(p_input[969]), .Z(n42705) );
  XOR U41700 ( .A(n42708), .B(n42707), .Z(n42706) );
  NOR U41701 ( .A(n21975), .B(p_input[967]), .Z(n42707) );
  XOR U41702 ( .A(n42710), .B(n42709), .Z(n42708) );
  NOR U41703 ( .A(n21977), .B(p_input[965]), .Z(n42709) );
  XOR U41704 ( .A(n42712), .B(n42711), .Z(n42710) );
  NOR U41705 ( .A(n21979), .B(p_input[963]), .Z(n42711) );
  XOR U41706 ( .A(n42714), .B(n42713), .Z(n42712) );
  NOR U41707 ( .A(n21981), .B(p_input[961]), .Z(n42713) );
  XOR U41708 ( .A(n42716), .B(n42715), .Z(n42714) );
  NOR U41709 ( .A(n21983), .B(p_input[959]), .Z(n42715) );
  XOR U41710 ( .A(n42718), .B(n42717), .Z(n42716) );
  NOR U41711 ( .A(n21985), .B(p_input[957]), .Z(n42717) );
  XOR U41712 ( .A(n42720), .B(n42719), .Z(n42718) );
  NOR U41713 ( .A(n21987), .B(p_input[955]), .Z(n42719) );
  XOR U41714 ( .A(n42722), .B(n42721), .Z(n42720) );
  NOR U41715 ( .A(n21989), .B(p_input[953]), .Z(n42721) );
  XOR U41716 ( .A(n42724), .B(n42723), .Z(n42722) );
  NOR U41717 ( .A(n21991), .B(p_input[951]), .Z(n42723) );
  XOR U41718 ( .A(n42726), .B(n42725), .Z(n42724) );
  NOR U41719 ( .A(n21993), .B(p_input[949]), .Z(n42725) );
  XOR U41720 ( .A(n42728), .B(n42727), .Z(n42726) );
  NOR U41721 ( .A(n21995), .B(p_input[947]), .Z(n42727) );
  XOR U41722 ( .A(n42730), .B(n42729), .Z(n42728) );
  NOR U41723 ( .A(n21997), .B(p_input[945]), .Z(n42729) );
  XOR U41724 ( .A(n42732), .B(n42731), .Z(n42730) );
  NOR U41725 ( .A(n21999), .B(p_input[943]), .Z(n42731) );
  XOR U41726 ( .A(n42734), .B(n42733), .Z(n42732) );
  NOR U41727 ( .A(n22001), .B(p_input[941]), .Z(n42733) );
  XOR U41728 ( .A(n42736), .B(n42735), .Z(n42734) );
  NOR U41729 ( .A(n22003), .B(p_input[939]), .Z(n42735) );
  XOR U41730 ( .A(n42738), .B(n42737), .Z(n42736) );
  NOR U41731 ( .A(n22005), .B(p_input[937]), .Z(n42737) );
  XOR U41732 ( .A(n42740), .B(n42739), .Z(n42738) );
  NOR U41733 ( .A(n22007), .B(p_input[935]), .Z(n42739) );
  XOR U41734 ( .A(n42742), .B(n42741), .Z(n42740) );
  NOR U41735 ( .A(n22009), .B(p_input[933]), .Z(n42741) );
  XOR U41736 ( .A(n42744), .B(n42743), .Z(n42742) );
  NOR U41737 ( .A(n22011), .B(p_input[931]), .Z(n42743) );
  XOR U41738 ( .A(n42746), .B(n42745), .Z(n42744) );
  NOR U41739 ( .A(n22013), .B(p_input[929]), .Z(n42745) );
  XOR U41740 ( .A(n42748), .B(n42747), .Z(n42746) );
  NOR U41741 ( .A(n22015), .B(p_input[927]), .Z(n42747) );
  XOR U41742 ( .A(n42750), .B(n42749), .Z(n42748) );
  NOR U41743 ( .A(n22017), .B(p_input[925]), .Z(n42749) );
  XOR U41744 ( .A(n42752), .B(n42751), .Z(n42750) );
  NOR U41745 ( .A(n22019), .B(p_input[923]), .Z(n42751) );
  XOR U41746 ( .A(n42754), .B(n42753), .Z(n42752) );
  NOR U41747 ( .A(n22021), .B(p_input[921]), .Z(n42753) );
  XOR U41748 ( .A(n42756), .B(n42755), .Z(n42754) );
  NOR U41749 ( .A(n22023), .B(p_input[919]), .Z(n42755) );
  XOR U41750 ( .A(n42758), .B(n42757), .Z(n42756) );
  NOR U41751 ( .A(n22025), .B(p_input[917]), .Z(n42757) );
  XOR U41752 ( .A(n42760), .B(n42759), .Z(n42758) );
  NOR U41753 ( .A(n22027), .B(p_input[915]), .Z(n42759) );
  XOR U41754 ( .A(n42762), .B(n42761), .Z(n42760) );
  NOR U41755 ( .A(n22029), .B(p_input[913]), .Z(n42761) );
  XOR U41756 ( .A(n42764), .B(n42763), .Z(n42762) );
  NOR U41757 ( .A(n22031), .B(p_input[911]), .Z(n42763) );
  XOR U41758 ( .A(n42766), .B(n42765), .Z(n42764) );
  NOR U41759 ( .A(n22033), .B(p_input[909]), .Z(n42765) );
  XOR U41760 ( .A(n42768), .B(n42767), .Z(n42766) );
  NOR U41761 ( .A(n22035), .B(p_input[907]), .Z(n42767) );
  XOR U41762 ( .A(n42770), .B(n42769), .Z(n42768) );
  NOR U41763 ( .A(n22037), .B(p_input[905]), .Z(n42769) );
  XOR U41764 ( .A(n42772), .B(n42771), .Z(n42770) );
  NOR U41765 ( .A(n22039), .B(p_input[903]), .Z(n42771) );
  XOR U41766 ( .A(n42774), .B(n42773), .Z(n42772) );
  NOR U41767 ( .A(n22041), .B(p_input[901]), .Z(n42773) );
  XOR U41768 ( .A(n42776), .B(n42775), .Z(n42774) );
  NOR U41769 ( .A(n22043), .B(p_input[899]), .Z(n42775) );
  XOR U41770 ( .A(n42778), .B(n42777), .Z(n42776) );
  NOR U41771 ( .A(n22045), .B(p_input[897]), .Z(n42777) );
  XOR U41772 ( .A(n42780), .B(n42779), .Z(n42778) );
  NOR U41773 ( .A(n22047), .B(p_input[895]), .Z(n42779) );
  XOR U41774 ( .A(n42782), .B(n42781), .Z(n42780) );
  NOR U41775 ( .A(n22049), .B(p_input[893]), .Z(n42781) );
  XOR U41776 ( .A(n42784), .B(n42783), .Z(n42782) );
  NOR U41777 ( .A(n22051), .B(p_input[891]), .Z(n42783) );
  XOR U41778 ( .A(n42786), .B(n42785), .Z(n42784) );
  NOR U41779 ( .A(n22053), .B(p_input[889]), .Z(n42785) );
  XOR U41780 ( .A(n42788), .B(n42787), .Z(n42786) );
  NOR U41781 ( .A(n22055), .B(p_input[887]), .Z(n42787) );
  XOR U41782 ( .A(n42790), .B(n42789), .Z(n42788) );
  NOR U41783 ( .A(n22057), .B(p_input[885]), .Z(n42789) );
  XOR U41784 ( .A(n42792), .B(n42791), .Z(n42790) );
  NOR U41785 ( .A(n22059), .B(p_input[883]), .Z(n42791) );
  XOR U41786 ( .A(n42794), .B(n42793), .Z(n42792) );
  NOR U41787 ( .A(n22061), .B(p_input[881]), .Z(n42793) );
  XOR U41788 ( .A(n42796), .B(n42795), .Z(n42794) );
  NOR U41789 ( .A(n22063), .B(p_input[879]), .Z(n42795) );
  XOR U41790 ( .A(n42798), .B(n42797), .Z(n42796) );
  NOR U41791 ( .A(n22065), .B(p_input[877]), .Z(n42797) );
  XOR U41792 ( .A(n42800), .B(n42799), .Z(n42798) );
  NOR U41793 ( .A(n22067), .B(p_input[875]), .Z(n42799) );
  XOR U41794 ( .A(n42802), .B(n42801), .Z(n42800) );
  NOR U41795 ( .A(n22069), .B(p_input[873]), .Z(n42801) );
  XOR U41796 ( .A(n42804), .B(n42803), .Z(n42802) );
  NOR U41797 ( .A(n22071), .B(p_input[871]), .Z(n42803) );
  XOR U41798 ( .A(n42806), .B(n42805), .Z(n42804) );
  NOR U41799 ( .A(n22073), .B(p_input[869]), .Z(n42805) );
  XOR U41800 ( .A(n42808), .B(n42807), .Z(n42806) );
  NOR U41801 ( .A(n22075), .B(p_input[867]), .Z(n42807) );
  XOR U41802 ( .A(n42810), .B(n42809), .Z(n42808) );
  NOR U41803 ( .A(n22077), .B(p_input[865]), .Z(n42809) );
  XOR U41804 ( .A(n42812), .B(n42811), .Z(n42810) );
  NOR U41805 ( .A(n22079), .B(p_input[863]), .Z(n42811) );
  XOR U41806 ( .A(n42814), .B(n42813), .Z(n42812) );
  NOR U41807 ( .A(n22081), .B(p_input[861]), .Z(n42813) );
  XOR U41808 ( .A(n42816), .B(n42815), .Z(n42814) );
  NOR U41809 ( .A(n22083), .B(p_input[859]), .Z(n42815) );
  XOR U41810 ( .A(n42818), .B(n42817), .Z(n42816) );
  NOR U41811 ( .A(n22085), .B(p_input[857]), .Z(n42817) );
  XOR U41812 ( .A(n42820), .B(n42819), .Z(n42818) );
  NOR U41813 ( .A(n22087), .B(p_input[855]), .Z(n42819) );
  XOR U41814 ( .A(n42822), .B(n42821), .Z(n42820) );
  NOR U41815 ( .A(n22089), .B(p_input[853]), .Z(n42821) );
  XOR U41816 ( .A(n42824), .B(n42823), .Z(n42822) );
  NOR U41817 ( .A(n22091), .B(p_input[851]), .Z(n42823) );
  XOR U41818 ( .A(n42826), .B(n42825), .Z(n42824) );
  NOR U41819 ( .A(n22093), .B(p_input[849]), .Z(n42825) );
  XOR U41820 ( .A(n42828), .B(n42827), .Z(n42826) );
  NOR U41821 ( .A(n22095), .B(p_input[847]), .Z(n42827) );
  XOR U41822 ( .A(n42830), .B(n42829), .Z(n42828) );
  NOR U41823 ( .A(n22097), .B(p_input[845]), .Z(n42829) );
  XOR U41824 ( .A(n42832), .B(n42831), .Z(n42830) );
  NOR U41825 ( .A(n22099), .B(p_input[843]), .Z(n42831) );
  XOR U41826 ( .A(n42834), .B(n42833), .Z(n42832) );
  NOR U41827 ( .A(n22101), .B(p_input[841]), .Z(n42833) );
  XOR U41828 ( .A(n42836), .B(n42835), .Z(n42834) );
  NOR U41829 ( .A(n22103), .B(p_input[839]), .Z(n42835) );
  XOR U41830 ( .A(n42838), .B(n42837), .Z(n42836) );
  NOR U41831 ( .A(n22105), .B(p_input[837]), .Z(n42837) );
  XOR U41832 ( .A(n42840), .B(n42839), .Z(n42838) );
  NOR U41833 ( .A(n22107), .B(p_input[835]), .Z(n42839) );
  XOR U41834 ( .A(n42842), .B(n42841), .Z(n42840) );
  NOR U41835 ( .A(n22109), .B(p_input[833]), .Z(n42841) );
  XOR U41836 ( .A(n42844), .B(n42843), .Z(n42842) );
  NOR U41837 ( .A(n22111), .B(p_input[831]), .Z(n42843) );
  XOR U41838 ( .A(n42846), .B(n42845), .Z(n42844) );
  NOR U41839 ( .A(n22113), .B(p_input[829]), .Z(n42845) );
  XOR U41840 ( .A(n42848), .B(n42847), .Z(n42846) );
  NOR U41841 ( .A(n22115), .B(p_input[827]), .Z(n42847) );
  XOR U41842 ( .A(n42850), .B(n42849), .Z(n42848) );
  NOR U41843 ( .A(n22117), .B(p_input[825]), .Z(n42849) );
  XOR U41844 ( .A(n42852), .B(n42851), .Z(n42850) );
  NOR U41845 ( .A(n22119), .B(p_input[823]), .Z(n42851) );
  XOR U41846 ( .A(n42854), .B(n42853), .Z(n42852) );
  NOR U41847 ( .A(n22121), .B(p_input[821]), .Z(n42853) );
  XOR U41848 ( .A(n42856), .B(n42855), .Z(n42854) );
  NOR U41849 ( .A(n22123), .B(p_input[819]), .Z(n42855) );
  XOR U41850 ( .A(n42858), .B(n42857), .Z(n42856) );
  NOR U41851 ( .A(n22125), .B(p_input[817]), .Z(n42857) );
  XOR U41852 ( .A(n42860), .B(n42859), .Z(n42858) );
  NOR U41853 ( .A(n22127), .B(p_input[815]), .Z(n42859) );
  XOR U41854 ( .A(n42862), .B(n42861), .Z(n42860) );
  NOR U41855 ( .A(n22129), .B(p_input[813]), .Z(n42861) );
  XOR U41856 ( .A(n42864), .B(n42863), .Z(n42862) );
  NOR U41857 ( .A(n22131), .B(p_input[811]), .Z(n42863) );
  XOR U41858 ( .A(n42866), .B(n42865), .Z(n42864) );
  NOR U41859 ( .A(n22133), .B(p_input[809]), .Z(n42865) );
  XOR U41860 ( .A(n42868), .B(n42867), .Z(n42866) );
  NOR U41861 ( .A(n22135), .B(p_input[807]), .Z(n42867) );
  XOR U41862 ( .A(n42870), .B(n42869), .Z(n42868) );
  NOR U41863 ( .A(n22137), .B(p_input[805]), .Z(n42869) );
  XOR U41864 ( .A(n42872), .B(n42871), .Z(n42870) );
  NOR U41865 ( .A(n22139), .B(p_input[803]), .Z(n42871) );
  XOR U41866 ( .A(n42874), .B(n42873), .Z(n42872) );
  NOR U41867 ( .A(n22141), .B(p_input[801]), .Z(n42873) );
  XOR U41868 ( .A(n42876), .B(n42875), .Z(n42874) );
  NOR U41869 ( .A(n22143), .B(p_input[799]), .Z(n42875) );
  XOR U41870 ( .A(n42878), .B(n42877), .Z(n42876) );
  NOR U41871 ( .A(n22145), .B(p_input[797]), .Z(n42877) );
  XOR U41872 ( .A(n42880), .B(n42879), .Z(n42878) );
  NOR U41873 ( .A(n22147), .B(p_input[795]), .Z(n42879) );
  XOR U41874 ( .A(n42882), .B(n42881), .Z(n42880) );
  NOR U41875 ( .A(n22149), .B(p_input[793]), .Z(n42881) );
  XOR U41876 ( .A(n42884), .B(n42883), .Z(n42882) );
  NOR U41877 ( .A(n22151), .B(p_input[791]), .Z(n42883) );
  XOR U41878 ( .A(n42886), .B(n42885), .Z(n42884) );
  NOR U41879 ( .A(n22153), .B(p_input[789]), .Z(n42885) );
  XOR U41880 ( .A(n42888), .B(n42887), .Z(n42886) );
  NOR U41881 ( .A(n22155), .B(p_input[787]), .Z(n42887) );
  XOR U41882 ( .A(n42890), .B(n42889), .Z(n42888) );
  NOR U41883 ( .A(n22157), .B(p_input[785]), .Z(n42889) );
  XOR U41884 ( .A(n42892), .B(n42891), .Z(n42890) );
  NOR U41885 ( .A(n22159), .B(p_input[783]), .Z(n42891) );
  XOR U41886 ( .A(n42894), .B(n42893), .Z(n42892) );
  NOR U41887 ( .A(n22161), .B(p_input[781]), .Z(n42893) );
  XOR U41888 ( .A(n42896), .B(n42895), .Z(n42894) );
  NOR U41889 ( .A(n22163), .B(p_input[779]), .Z(n42895) );
  XOR U41890 ( .A(n42898), .B(n42897), .Z(n42896) );
  NOR U41891 ( .A(n22165), .B(p_input[777]), .Z(n42897) );
  XOR U41892 ( .A(n42900), .B(n42899), .Z(n42898) );
  NOR U41893 ( .A(n22167), .B(p_input[775]), .Z(n42899) );
  XOR U41894 ( .A(n42902), .B(n42901), .Z(n42900) );
  NOR U41895 ( .A(n22169), .B(p_input[773]), .Z(n42901) );
  XOR U41896 ( .A(n42904), .B(n42903), .Z(n42902) );
  NOR U41897 ( .A(n22171), .B(p_input[771]), .Z(n42903) );
  XOR U41898 ( .A(n42906), .B(n42905), .Z(n42904) );
  NOR U41899 ( .A(n22173), .B(p_input[769]), .Z(n42905) );
  XOR U41900 ( .A(n42908), .B(n42907), .Z(n42906) );
  NOR U41901 ( .A(n22175), .B(p_input[767]), .Z(n42907) );
  XOR U41902 ( .A(n42910), .B(n42909), .Z(n42908) );
  NOR U41903 ( .A(n22177), .B(p_input[765]), .Z(n42909) );
  XOR U41904 ( .A(n42912), .B(n42911), .Z(n42910) );
  NOR U41905 ( .A(n22179), .B(p_input[763]), .Z(n42911) );
  XOR U41906 ( .A(n42914), .B(n42913), .Z(n42912) );
  NOR U41907 ( .A(n22181), .B(p_input[761]), .Z(n42913) );
  XOR U41908 ( .A(n42916), .B(n42915), .Z(n42914) );
  NOR U41909 ( .A(n22183), .B(p_input[759]), .Z(n42915) );
  XOR U41910 ( .A(n42918), .B(n42917), .Z(n42916) );
  NOR U41911 ( .A(n22185), .B(p_input[757]), .Z(n42917) );
  XOR U41912 ( .A(n42920), .B(n42919), .Z(n42918) );
  NOR U41913 ( .A(n22187), .B(p_input[755]), .Z(n42919) );
  XOR U41914 ( .A(n42922), .B(n42921), .Z(n42920) );
  NOR U41915 ( .A(n22189), .B(p_input[753]), .Z(n42921) );
  XOR U41916 ( .A(n42924), .B(n42923), .Z(n42922) );
  NOR U41917 ( .A(n22191), .B(p_input[751]), .Z(n42923) );
  XOR U41918 ( .A(n42926), .B(n42925), .Z(n42924) );
  NOR U41919 ( .A(n22193), .B(p_input[749]), .Z(n42925) );
  XOR U41920 ( .A(n42928), .B(n42927), .Z(n42926) );
  NOR U41921 ( .A(n22195), .B(p_input[747]), .Z(n42927) );
  XOR U41922 ( .A(n42930), .B(n42929), .Z(n42928) );
  NOR U41923 ( .A(n22197), .B(p_input[745]), .Z(n42929) );
  XOR U41924 ( .A(n42932), .B(n42931), .Z(n42930) );
  NOR U41925 ( .A(n22199), .B(p_input[743]), .Z(n42931) );
  XOR U41926 ( .A(n42934), .B(n42933), .Z(n42932) );
  NOR U41927 ( .A(n22201), .B(p_input[741]), .Z(n42933) );
  XOR U41928 ( .A(n42936), .B(n42935), .Z(n42934) );
  NOR U41929 ( .A(n22203), .B(p_input[739]), .Z(n42935) );
  XOR U41930 ( .A(n42938), .B(n42937), .Z(n42936) );
  NOR U41931 ( .A(n22205), .B(p_input[737]), .Z(n42937) );
  XOR U41932 ( .A(n42940), .B(n42939), .Z(n42938) );
  NOR U41933 ( .A(n22207), .B(p_input[735]), .Z(n42939) );
  XOR U41934 ( .A(n42942), .B(n42941), .Z(n42940) );
  NOR U41935 ( .A(n22209), .B(p_input[733]), .Z(n42941) );
  XOR U41936 ( .A(n42944), .B(n42943), .Z(n42942) );
  NOR U41937 ( .A(n22211), .B(p_input[731]), .Z(n42943) );
  XOR U41938 ( .A(n42946), .B(n42945), .Z(n42944) );
  NOR U41939 ( .A(n22213), .B(p_input[729]), .Z(n42945) );
  XOR U41940 ( .A(n42948), .B(n42947), .Z(n42946) );
  NOR U41941 ( .A(n22215), .B(p_input[727]), .Z(n42947) );
  XOR U41942 ( .A(n42950), .B(n42949), .Z(n42948) );
  NOR U41943 ( .A(n22217), .B(p_input[725]), .Z(n42949) );
  XOR U41944 ( .A(n42952), .B(n42951), .Z(n42950) );
  NOR U41945 ( .A(n22219), .B(p_input[723]), .Z(n42951) );
  XOR U41946 ( .A(n42954), .B(n42953), .Z(n42952) );
  NOR U41947 ( .A(n22221), .B(p_input[721]), .Z(n42953) );
  XOR U41948 ( .A(n42956), .B(n42955), .Z(n42954) );
  NOR U41949 ( .A(n22223), .B(p_input[719]), .Z(n42955) );
  XOR U41950 ( .A(n42958), .B(n42957), .Z(n42956) );
  NOR U41951 ( .A(n22225), .B(p_input[717]), .Z(n42957) );
  XOR U41952 ( .A(n42960), .B(n42959), .Z(n42958) );
  NOR U41953 ( .A(n22227), .B(p_input[715]), .Z(n42959) );
  XOR U41954 ( .A(n42962), .B(n42961), .Z(n42960) );
  NOR U41955 ( .A(n22229), .B(p_input[713]), .Z(n42961) );
  XOR U41956 ( .A(n42964), .B(n42963), .Z(n42962) );
  NOR U41957 ( .A(n22231), .B(p_input[711]), .Z(n42963) );
  XOR U41958 ( .A(n42966), .B(n42965), .Z(n42964) );
  NOR U41959 ( .A(n22233), .B(p_input[709]), .Z(n42965) );
  XOR U41960 ( .A(n42968), .B(n42967), .Z(n42966) );
  NOR U41961 ( .A(n22235), .B(p_input[707]), .Z(n42967) );
  XOR U41962 ( .A(n42970), .B(n42969), .Z(n42968) );
  NOR U41963 ( .A(n22237), .B(p_input[705]), .Z(n42969) );
  XOR U41964 ( .A(n42972), .B(n42971), .Z(n42970) );
  NOR U41965 ( .A(n22239), .B(p_input[703]), .Z(n42971) );
  XOR U41966 ( .A(n42974), .B(n42973), .Z(n42972) );
  NOR U41967 ( .A(n22241), .B(p_input[701]), .Z(n42973) );
  XOR U41968 ( .A(n42976), .B(n42975), .Z(n42974) );
  NOR U41969 ( .A(n22243), .B(p_input[699]), .Z(n42975) );
  XOR U41970 ( .A(n42978), .B(n42977), .Z(n42976) );
  NOR U41971 ( .A(n22245), .B(p_input[697]), .Z(n42977) );
  XOR U41972 ( .A(n42980), .B(n42979), .Z(n42978) );
  NOR U41973 ( .A(n22247), .B(p_input[695]), .Z(n42979) );
  XOR U41974 ( .A(n42982), .B(n42981), .Z(n42980) );
  NOR U41975 ( .A(n22249), .B(p_input[693]), .Z(n42981) );
  XOR U41976 ( .A(n42984), .B(n42983), .Z(n42982) );
  NOR U41977 ( .A(n22251), .B(p_input[691]), .Z(n42983) );
  XOR U41978 ( .A(n42986), .B(n42985), .Z(n42984) );
  NOR U41979 ( .A(n22253), .B(p_input[689]), .Z(n42985) );
  XOR U41980 ( .A(n42988), .B(n42987), .Z(n42986) );
  NOR U41981 ( .A(n22255), .B(p_input[687]), .Z(n42987) );
  XOR U41982 ( .A(n42990), .B(n42989), .Z(n42988) );
  NOR U41983 ( .A(n22257), .B(p_input[685]), .Z(n42989) );
  XOR U41984 ( .A(n42992), .B(n42991), .Z(n42990) );
  NOR U41985 ( .A(n22259), .B(p_input[683]), .Z(n42991) );
  XOR U41986 ( .A(n42994), .B(n42993), .Z(n42992) );
  NOR U41987 ( .A(n22261), .B(p_input[681]), .Z(n42993) );
  XOR U41988 ( .A(n42996), .B(n42995), .Z(n42994) );
  NOR U41989 ( .A(n22263), .B(p_input[679]), .Z(n42995) );
  XOR U41990 ( .A(n42998), .B(n42997), .Z(n42996) );
  NOR U41991 ( .A(n22265), .B(p_input[677]), .Z(n42997) );
  XOR U41992 ( .A(n43000), .B(n42999), .Z(n42998) );
  NOR U41993 ( .A(n22267), .B(p_input[675]), .Z(n42999) );
  XOR U41994 ( .A(n43002), .B(n43001), .Z(n43000) );
  NOR U41995 ( .A(n22269), .B(p_input[673]), .Z(n43001) );
  XOR U41996 ( .A(n43004), .B(n43003), .Z(n43002) );
  NOR U41997 ( .A(n22271), .B(p_input[671]), .Z(n43003) );
  XOR U41998 ( .A(n43006), .B(n43005), .Z(n43004) );
  NOR U41999 ( .A(n22273), .B(p_input[669]), .Z(n43005) );
  XOR U42000 ( .A(n43008), .B(n43007), .Z(n43006) );
  NOR U42001 ( .A(n22275), .B(p_input[667]), .Z(n43007) );
  XOR U42002 ( .A(n43010), .B(n43009), .Z(n43008) );
  NOR U42003 ( .A(n22277), .B(p_input[665]), .Z(n43009) );
  XOR U42004 ( .A(n43012), .B(n43011), .Z(n43010) );
  NOR U42005 ( .A(n22279), .B(p_input[663]), .Z(n43011) );
  XOR U42006 ( .A(n43014), .B(n43013), .Z(n43012) );
  NOR U42007 ( .A(n22281), .B(p_input[661]), .Z(n43013) );
  XOR U42008 ( .A(n43016), .B(n43015), .Z(n43014) );
  NOR U42009 ( .A(n22283), .B(p_input[659]), .Z(n43015) );
  XOR U42010 ( .A(n43018), .B(n43017), .Z(n43016) );
  NOR U42011 ( .A(n22285), .B(p_input[657]), .Z(n43017) );
  XOR U42012 ( .A(n43020), .B(n43019), .Z(n43018) );
  NOR U42013 ( .A(n22287), .B(p_input[655]), .Z(n43019) );
  XOR U42014 ( .A(n43022), .B(n43021), .Z(n43020) );
  NOR U42015 ( .A(n22289), .B(p_input[653]), .Z(n43021) );
  XOR U42016 ( .A(n43024), .B(n43023), .Z(n43022) );
  NOR U42017 ( .A(n22291), .B(p_input[651]), .Z(n43023) );
  XOR U42018 ( .A(n43026), .B(n43025), .Z(n43024) );
  NOR U42019 ( .A(n22293), .B(p_input[649]), .Z(n43025) );
  XOR U42020 ( .A(n43028), .B(n43027), .Z(n43026) );
  NOR U42021 ( .A(n22295), .B(p_input[647]), .Z(n43027) );
  XOR U42022 ( .A(n43030), .B(n43029), .Z(n43028) );
  NOR U42023 ( .A(n22297), .B(p_input[645]), .Z(n43029) );
  XOR U42024 ( .A(n43032), .B(n43031), .Z(n43030) );
  NOR U42025 ( .A(n22299), .B(p_input[643]), .Z(n43031) );
  XOR U42026 ( .A(n43034), .B(n43033), .Z(n43032) );
  NOR U42027 ( .A(n22301), .B(p_input[641]), .Z(n43033) );
  XOR U42028 ( .A(n43036), .B(n43035), .Z(n43034) );
  NOR U42029 ( .A(n22303), .B(p_input[639]), .Z(n43035) );
  XOR U42030 ( .A(n43038), .B(n43037), .Z(n43036) );
  NOR U42031 ( .A(n22305), .B(p_input[637]), .Z(n43037) );
  XOR U42032 ( .A(n43040), .B(n43039), .Z(n43038) );
  NOR U42033 ( .A(n22307), .B(p_input[635]), .Z(n43039) );
  XOR U42034 ( .A(n43042), .B(n43041), .Z(n43040) );
  NOR U42035 ( .A(n22309), .B(p_input[633]), .Z(n43041) );
  XOR U42036 ( .A(n43044), .B(n43043), .Z(n43042) );
  NOR U42037 ( .A(n22311), .B(p_input[631]), .Z(n43043) );
  XOR U42038 ( .A(n43046), .B(n43045), .Z(n43044) );
  NOR U42039 ( .A(n22313), .B(p_input[629]), .Z(n43045) );
  XOR U42040 ( .A(n43048), .B(n43047), .Z(n43046) );
  NOR U42041 ( .A(n22315), .B(p_input[627]), .Z(n43047) );
  XOR U42042 ( .A(n43050), .B(n43049), .Z(n43048) );
  NOR U42043 ( .A(n22317), .B(p_input[625]), .Z(n43049) );
  XOR U42044 ( .A(n43052), .B(n43051), .Z(n43050) );
  NOR U42045 ( .A(n22319), .B(p_input[623]), .Z(n43051) );
  XOR U42046 ( .A(n43054), .B(n43053), .Z(n43052) );
  NOR U42047 ( .A(n22321), .B(p_input[621]), .Z(n43053) );
  XOR U42048 ( .A(n43056), .B(n43055), .Z(n43054) );
  NOR U42049 ( .A(n22323), .B(p_input[619]), .Z(n43055) );
  XOR U42050 ( .A(n43058), .B(n43057), .Z(n43056) );
  NOR U42051 ( .A(n22325), .B(p_input[617]), .Z(n43057) );
  XOR U42052 ( .A(n43060), .B(n43059), .Z(n43058) );
  NOR U42053 ( .A(n22327), .B(p_input[615]), .Z(n43059) );
  XOR U42054 ( .A(n43062), .B(n43061), .Z(n43060) );
  NOR U42055 ( .A(n22329), .B(p_input[613]), .Z(n43061) );
  XOR U42056 ( .A(n43064), .B(n43063), .Z(n43062) );
  NOR U42057 ( .A(n22331), .B(p_input[611]), .Z(n43063) );
  XOR U42058 ( .A(n43066), .B(n43065), .Z(n43064) );
  NOR U42059 ( .A(n22333), .B(p_input[609]), .Z(n43065) );
  XOR U42060 ( .A(n43068), .B(n43067), .Z(n43066) );
  NOR U42061 ( .A(n22335), .B(p_input[607]), .Z(n43067) );
  XOR U42062 ( .A(n43070), .B(n43069), .Z(n43068) );
  NOR U42063 ( .A(n22337), .B(p_input[605]), .Z(n43069) );
  XOR U42064 ( .A(n43072), .B(n43071), .Z(n43070) );
  NOR U42065 ( .A(n22339), .B(p_input[603]), .Z(n43071) );
  XOR U42066 ( .A(n43074), .B(n43073), .Z(n43072) );
  NOR U42067 ( .A(n22341), .B(p_input[601]), .Z(n43073) );
  XOR U42068 ( .A(n43076), .B(n43075), .Z(n43074) );
  NOR U42069 ( .A(n22343), .B(p_input[599]), .Z(n43075) );
  XOR U42070 ( .A(n43078), .B(n43077), .Z(n43076) );
  NOR U42071 ( .A(n22345), .B(p_input[597]), .Z(n43077) );
  XOR U42072 ( .A(n43080), .B(n43079), .Z(n43078) );
  NOR U42073 ( .A(n22347), .B(p_input[595]), .Z(n43079) );
  XOR U42074 ( .A(n43082), .B(n43081), .Z(n43080) );
  NOR U42075 ( .A(n22349), .B(p_input[593]), .Z(n43081) );
  XOR U42076 ( .A(n43084), .B(n43083), .Z(n43082) );
  NOR U42077 ( .A(n22351), .B(p_input[591]), .Z(n43083) );
  XOR U42078 ( .A(n43086), .B(n43085), .Z(n43084) );
  NOR U42079 ( .A(n22353), .B(p_input[589]), .Z(n43085) );
  XOR U42080 ( .A(n43088), .B(n43087), .Z(n43086) );
  NOR U42081 ( .A(n22355), .B(p_input[587]), .Z(n43087) );
  XOR U42082 ( .A(n43090), .B(n43089), .Z(n43088) );
  NOR U42083 ( .A(n22357), .B(p_input[585]), .Z(n43089) );
  XOR U42084 ( .A(n43092), .B(n43091), .Z(n43090) );
  NOR U42085 ( .A(n22359), .B(p_input[583]), .Z(n43091) );
  XOR U42086 ( .A(n43094), .B(n43093), .Z(n43092) );
  NOR U42087 ( .A(n22361), .B(p_input[581]), .Z(n43093) );
  XOR U42088 ( .A(n43096), .B(n43095), .Z(n43094) );
  NOR U42089 ( .A(n22363), .B(p_input[579]), .Z(n43095) );
  XOR U42090 ( .A(n43098), .B(n43097), .Z(n43096) );
  NOR U42091 ( .A(n22365), .B(p_input[577]), .Z(n43097) );
  XOR U42092 ( .A(n43100), .B(n43099), .Z(n43098) );
  NOR U42093 ( .A(n22367), .B(p_input[575]), .Z(n43099) );
  XOR U42094 ( .A(n43102), .B(n43101), .Z(n43100) );
  NOR U42095 ( .A(n22369), .B(p_input[573]), .Z(n43101) );
  XOR U42096 ( .A(n43104), .B(n43103), .Z(n43102) );
  NOR U42097 ( .A(n22371), .B(p_input[571]), .Z(n43103) );
  XOR U42098 ( .A(n43106), .B(n43105), .Z(n43104) );
  NOR U42099 ( .A(n22373), .B(p_input[569]), .Z(n43105) );
  XOR U42100 ( .A(n43108), .B(n43107), .Z(n43106) );
  NOR U42101 ( .A(n22375), .B(p_input[567]), .Z(n43107) );
  XOR U42102 ( .A(n43110), .B(n43109), .Z(n43108) );
  NOR U42103 ( .A(n22377), .B(p_input[565]), .Z(n43109) );
  XOR U42104 ( .A(n43112), .B(n43111), .Z(n43110) );
  NOR U42105 ( .A(n22379), .B(p_input[563]), .Z(n43111) );
  XOR U42106 ( .A(n43114), .B(n43113), .Z(n43112) );
  NOR U42107 ( .A(n22381), .B(p_input[561]), .Z(n43113) );
  XOR U42108 ( .A(n43116), .B(n43115), .Z(n43114) );
  NOR U42109 ( .A(n22383), .B(p_input[559]), .Z(n43115) );
  XOR U42110 ( .A(n43118), .B(n43117), .Z(n43116) );
  NOR U42111 ( .A(n22385), .B(p_input[557]), .Z(n43117) );
  XOR U42112 ( .A(n43120), .B(n43119), .Z(n43118) );
  NOR U42113 ( .A(n22387), .B(p_input[555]), .Z(n43119) );
  XOR U42114 ( .A(n43122), .B(n43121), .Z(n43120) );
  NOR U42115 ( .A(n22389), .B(p_input[553]), .Z(n43121) );
  XOR U42116 ( .A(n43124), .B(n43123), .Z(n43122) );
  NOR U42117 ( .A(n22391), .B(p_input[551]), .Z(n43123) );
  XOR U42118 ( .A(n43126), .B(n43125), .Z(n43124) );
  NOR U42119 ( .A(n22393), .B(p_input[549]), .Z(n43125) );
  XOR U42120 ( .A(n43128), .B(n43127), .Z(n43126) );
  NOR U42121 ( .A(n22395), .B(p_input[547]), .Z(n43127) );
  XOR U42122 ( .A(n43130), .B(n43129), .Z(n43128) );
  NOR U42123 ( .A(n22397), .B(p_input[545]), .Z(n43129) );
  XOR U42124 ( .A(n43132), .B(n43131), .Z(n43130) );
  NOR U42125 ( .A(n22399), .B(p_input[543]), .Z(n43131) );
  XOR U42126 ( .A(n43134), .B(n43133), .Z(n43132) );
  NOR U42127 ( .A(n22401), .B(p_input[541]), .Z(n43133) );
  XOR U42128 ( .A(n43136), .B(n43135), .Z(n43134) );
  NOR U42129 ( .A(n22403), .B(p_input[539]), .Z(n43135) );
  XOR U42130 ( .A(n43138), .B(n43137), .Z(n43136) );
  NOR U42131 ( .A(n22405), .B(p_input[537]), .Z(n43137) );
  XOR U42132 ( .A(n43140), .B(n43139), .Z(n43138) );
  NOR U42133 ( .A(n22407), .B(p_input[535]), .Z(n43139) );
  XOR U42134 ( .A(n43142), .B(n43141), .Z(n43140) );
  NOR U42135 ( .A(n22409), .B(p_input[533]), .Z(n43141) );
  XOR U42136 ( .A(n43144), .B(n43143), .Z(n43142) );
  NOR U42137 ( .A(n22411), .B(p_input[531]), .Z(n43143) );
  XOR U42138 ( .A(n43146), .B(n43145), .Z(n43144) );
  NOR U42139 ( .A(n22413), .B(p_input[529]), .Z(n43145) );
  XOR U42140 ( .A(n43148), .B(n43147), .Z(n43146) );
  NOR U42141 ( .A(n22415), .B(p_input[527]), .Z(n43147) );
  XOR U42142 ( .A(n43150), .B(n43149), .Z(n43148) );
  NOR U42143 ( .A(n22417), .B(p_input[525]), .Z(n43149) );
  XOR U42144 ( .A(n43152), .B(n43151), .Z(n43150) );
  NOR U42145 ( .A(n22419), .B(p_input[523]), .Z(n43151) );
  XOR U42146 ( .A(n43154), .B(n43153), .Z(n43152) );
  NOR U42147 ( .A(n22421), .B(p_input[521]), .Z(n43153) );
  XOR U42148 ( .A(n43156), .B(n43155), .Z(n43154) );
  NOR U42149 ( .A(n22423), .B(p_input[519]), .Z(n43155) );
  XOR U42150 ( .A(n43158), .B(n43157), .Z(n43156) );
  NOR U42151 ( .A(n22425), .B(p_input[517]), .Z(n43157) );
  XOR U42152 ( .A(n43160), .B(n43159), .Z(n43158) );
  NOR U42153 ( .A(n22427), .B(p_input[515]), .Z(n43159) );
  XOR U42154 ( .A(n43162), .B(n43161), .Z(n43160) );
  NOR U42155 ( .A(n22429), .B(p_input[513]), .Z(n43161) );
  XOR U42156 ( .A(n43164), .B(n43163), .Z(n43162) );
  NOR U42157 ( .A(n22431), .B(p_input[511]), .Z(n43163) );
  XOR U42158 ( .A(n43166), .B(n43165), .Z(n43164) );
  NOR U42159 ( .A(n22433), .B(p_input[509]), .Z(n43165) );
  XOR U42160 ( .A(n43168), .B(n43167), .Z(n43166) );
  NOR U42161 ( .A(n22435), .B(p_input[507]), .Z(n43167) );
  XOR U42162 ( .A(n43170), .B(n43169), .Z(n43168) );
  NOR U42163 ( .A(n22437), .B(p_input[505]), .Z(n43169) );
  XOR U42164 ( .A(n43172), .B(n43171), .Z(n43170) );
  NOR U42165 ( .A(n22439), .B(p_input[503]), .Z(n43171) );
  XOR U42166 ( .A(n43174), .B(n43173), .Z(n43172) );
  NOR U42167 ( .A(n22441), .B(p_input[501]), .Z(n43173) );
  XOR U42168 ( .A(n43176), .B(n43175), .Z(n43174) );
  NOR U42169 ( .A(n22443), .B(p_input[499]), .Z(n43175) );
  XOR U42170 ( .A(n43178), .B(n43177), .Z(n43176) );
  NOR U42171 ( .A(n22445), .B(p_input[497]), .Z(n43177) );
  XOR U42172 ( .A(n43180), .B(n43179), .Z(n43178) );
  NOR U42173 ( .A(n22447), .B(p_input[495]), .Z(n43179) );
  XOR U42174 ( .A(n43182), .B(n43181), .Z(n43180) );
  NOR U42175 ( .A(n22449), .B(p_input[493]), .Z(n43181) );
  XOR U42176 ( .A(n43184), .B(n43183), .Z(n43182) );
  NOR U42177 ( .A(n22451), .B(p_input[491]), .Z(n43183) );
  XOR U42178 ( .A(n43186), .B(n43185), .Z(n43184) );
  NOR U42179 ( .A(n22453), .B(p_input[489]), .Z(n43185) );
  XOR U42180 ( .A(n43188), .B(n43187), .Z(n43186) );
  NOR U42181 ( .A(n22455), .B(p_input[487]), .Z(n43187) );
  XOR U42182 ( .A(n43190), .B(n43189), .Z(n43188) );
  NOR U42183 ( .A(n22457), .B(p_input[485]), .Z(n43189) );
  XOR U42184 ( .A(n43192), .B(n43191), .Z(n43190) );
  NOR U42185 ( .A(n22459), .B(p_input[483]), .Z(n43191) );
  XOR U42186 ( .A(n43194), .B(n43193), .Z(n43192) );
  NOR U42187 ( .A(n22461), .B(p_input[481]), .Z(n43193) );
  XOR U42188 ( .A(n43196), .B(n43195), .Z(n43194) );
  NOR U42189 ( .A(n22463), .B(p_input[479]), .Z(n43195) );
  XOR U42190 ( .A(n43198), .B(n43197), .Z(n43196) );
  NOR U42191 ( .A(n22465), .B(p_input[477]), .Z(n43197) );
  XOR U42192 ( .A(n43200), .B(n43199), .Z(n43198) );
  NOR U42193 ( .A(n22467), .B(p_input[475]), .Z(n43199) );
  XOR U42194 ( .A(n43202), .B(n43201), .Z(n43200) );
  NOR U42195 ( .A(n22469), .B(p_input[473]), .Z(n43201) );
  XOR U42196 ( .A(n43204), .B(n43203), .Z(n43202) );
  NOR U42197 ( .A(n22471), .B(p_input[471]), .Z(n43203) );
  XOR U42198 ( .A(n43206), .B(n43205), .Z(n43204) );
  NOR U42199 ( .A(n22473), .B(p_input[469]), .Z(n43205) );
  XOR U42200 ( .A(n43208), .B(n43207), .Z(n43206) );
  NOR U42201 ( .A(n22475), .B(p_input[467]), .Z(n43207) );
  XOR U42202 ( .A(n43210), .B(n43209), .Z(n43208) );
  NOR U42203 ( .A(n22477), .B(p_input[465]), .Z(n43209) );
  XOR U42204 ( .A(n43212), .B(n43211), .Z(n43210) );
  NOR U42205 ( .A(n22479), .B(p_input[463]), .Z(n43211) );
  XOR U42206 ( .A(n43214), .B(n43213), .Z(n43212) );
  NOR U42207 ( .A(n22481), .B(p_input[461]), .Z(n43213) );
  XOR U42208 ( .A(n43216), .B(n43215), .Z(n43214) );
  NOR U42209 ( .A(n22483), .B(p_input[459]), .Z(n43215) );
  XOR U42210 ( .A(n43218), .B(n43217), .Z(n43216) );
  NOR U42211 ( .A(n22485), .B(p_input[457]), .Z(n43217) );
  XOR U42212 ( .A(n43220), .B(n43219), .Z(n43218) );
  NOR U42213 ( .A(n22487), .B(p_input[455]), .Z(n43219) );
  XOR U42214 ( .A(n43222), .B(n43221), .Z(n43220) );
  NOR U42215 ( .A(n22489), .B(p_input[453]), .Z(n43221) );
  XOR U42216 ( .A(n43224), .B(n43223), .Z(n43222) );
  NOR U42217 ( .A(n22491), .B(p_input[451]), .Z(n43223) );
  XOR U42218 ( .A(n43226), .B(n43225), .Z(n43224) );
  NOR U42219 ( .A(n22493), .B(p_input[449]), .Z(n43225) );
  XOR U42220 ( .A(n43228), .B(n43227), .Z(n43226) );
  NOR U42221 ( .A(n22495), .B(p_input[447]), .Z(n43227) );
  XOR U42222 ( .A(n43230), .B(n43229), .Z(n43228) );
  NOR U42223 ( .A(n22497), .B(p_input[445]), .Z(n43229) );
  XOR U42224 ( .A(n43232), .B(n43231), .Z(n43230) );
  NOR U42225 ( .A(n22499), .B(p_input[443]), .Z(n43231) );
  XOR U42226 ( .A(n43234), .B(n43233), .Z(n43232) );
  NOR U42227 ( .A(n22501), .B(p_input[441]), .Z(n43233) );
  XOR U42228 ( .A(n43236), .B(n43235), .Z(n43234) );
  NOR U42229 ( .A(n22503), .B(p_input[439]), .Z(n43235) );
  XOR U42230 ( .A(n43238), .B(n43237), .Z(n43236) );
  NOR U42231 ( .A(n22505), .B(p_input[437]), .Z(n43237) );
  XOR U42232 ( .A(n43240), .B(n43239), .Z(n43238) );
  NOR U42233 ( .A(n22507), .B(p_input[435]), .Z(n43239) );
  XOR U42234 ( .A(n43242), .B(n43241), .Z(n43240) );
  NOR U42235 ( .A(n22509), .B(p_input[433]), .Z(n43241) );
  XOR U42236 ( .A(n43244), .B(n43243), .Z(n43242) );
  NOR U42237 ( .A(n22511), .B(p_input[431]), .Z(n43243) );
  XOR U42238 ( .A(n43246), .B(n43245), .Z(n43244) );
  NOR U42239 ( .A(n22513), .B(p_input[429]), .Z(n43245) );
  XOR U42240 ( .A(n43248), .B(n43247), .Z(n43246) );
  NOR U42241 ( .A(n22515), .B(p_input[427]), .Z(n43247) );
  XOR U42242 ( .A(n43250), .B(n43249), .Z(n43248) );
  NOR U42243 ( .A(n22517), .B(p_input[425]), .Z(n43249) );
  XOR U42244 ( .A(n43252), .B(n43251), .Z(n43250) );
  NOR U42245 ( .A(n22519), .B(p_input[423]), .Z(n43251) );
  XOR U42246 ( .A(n43254), .B(n43253), .Z(n43252) );
  NOR U42247 ( .A(n22521), .B(p_input[421]), .Z(n43253) );
  XOR U42248 ( .A(n43256), .B(n43255), .Z(n43254) );
  NOR U42249 ( .A(n22523), .B(p_input[419]), .Z(n43255) );
  XOR U42250 ( .A(n43258), .B(n43257), .Z(n43256) );
  NOR U42251 ( .A(n22525), .B(p_input[417]), .Z(n43257) );
  XOR U42252 ( .A(n43260), .B(n43259), .Z(n43258) );
  NOR U42253 ( .A(n22527), .B(p_input[415]), .Z(n43259) );
  XOR U42254 ( .A(n43262), .B(n43261), .Z(n43260) );
  NOR U42255 ( .A(n22529), .B(p_input[413]), .Z(n43261) );
  XOR U42256 ( .A(n43264), .B(n43263), .Z(n43262) );
  NOR U42257 ( .A(n22531), .B(p_input[411]), .Z(n43263) );
  XOR U42258 ( .A(n43266), .B(n43265), .Z(n43264) );
  NOR U42259 ( .A(n22533), .B(p_input[409]), .Z(n43265) );
  XOR U42260 ( .A(n43268), .B(n43267), .Z(n43266) );
  NOR U42261 ( .A(n22535), .B(p_input[407]), .Z(n43267) );
  XOR U42262 ( .A(n43270), .B(n43269), .Z(n43268) );
  NOR U42263 ( .A(n22537), .B(p_input[405]), .Z(n43269) );
  XOR U42264 ( .A(n43272), .B(n43271), .Z(n43270) );
  NOR U42265 ( .A(n22539), .B(p_input[403]), .Z(n43271) );
  XOR U42266 ( .A(n43274), .B(n43273), .Z(n43272) );
  NOR U42267 ( .A(n22541), .B(p_input[401]), .Z(n43273) );
  XOR U42268 ( .A(n43276), .B(n43275), .Z(n43274) );
  NOR U42269 ( .A(n22543), .B(p_input[399]), .Z(n43275) );
  XOR U42270 ( .A(n43278), .B(n43277), .Z(n43276) );
  NOR U42271 ( .A(n22545), .B(p_input[397]), .Z(n43277) );
  XOR U42272 ( .A(n43280), .B(n43279), .Z(n43278) );
  NOR U42273 ( .A(n22547), .B(p_input[395]), .Z(n43279) );
  XOR U42274 ( .A(n43282), .B(n43281), .Z(n43280) );
  NOR U42275 ( .A(n22549), .B(p_input[393]), .Z(n43281) );
  XOR U42276 ( .A(n43284), .B(n43283), .Z(n43282) );
  NOR U42277 ( .A(n22551), .B(p_input[391]), .Z(n43283) );
  XOR U42278 ( .A(n43286), .B(n43285), .Z(n43284) );
  NOR U42279 ( .A(n22553), .B(p_input[389]), .Z(n43285) );
  XOR U42280 ( .A(n43288), .B(n43287), .Z(n43286) );
  NOR U42281 ( .A(n22555), .B(p_input[387]), .Z(n43287) );
  XOR U42282 ( .A(n43290), .B(n43289), .Z(n43288) );
  NOR U42283 ( .A(n22557), .B(p_input[385]), .Z(n43289) );
  XOR U42284 ( .A(n43292), .B(n43291), .Z(n43290) );
  NOR U42285 ( .A(n22559), .B(p_input[383]), .Z(n43291) );
  XOR U42286 ( .A(n43294), .B(n43293), .Z(n43292) );
  NOR U42287 ( .A(n22561), .B(p_input[381]), .Z(n43293) );
  XOR U42288 ( .A(n43296), .B(n43295), .Z(n43294) );
  NOR U42289 ( .A(n22563), .B(p_input[379]), .Z(n43295) );
  XOR U42290 ( .A(n43298), .B(n43297), .Z(n43296) );
  NOR U42291 ( .A(n22565), .B(p_input[377]), .Z(n43297) );
  XOR U42292 ( .A(n43300), .B(n43299), .Z(n43298) );
  NOR U42293 ( .A(n22567), .B(p_input[375]), .Z(n43299) );
  XOR U42294 ( .A(n43302), .B(n43301), .Z(n43300) );
  NOR U42295 ( .A(n22569), .B(p_input[373]), .Z(n43301) );
  XOR U42296 ( .A(n43304), .B(n43303), .Z(n43302) );
  NOR U42297 ( .A(n22571), .B(p_input[371]), .Z(n43303) );
  XOR U42298 ( .A(n43306), .B(n43305), .Z(n43304) );
  NOR U42299 ( .A(n22573), .B(p_input[369]), .Z(n43305) );
  XOR U42300 ( .A(n43308), .B(n43307), .Z(n43306) );
  NOR U42301 ( .A(n22575), .B(p_input[367]), .Z(n43307) );
  XOR U42302 ( .A(n43310), .B(n43309), .Z(n43308) );
  NOR U42303 ( .A(n22577), .B(p_input[365]), .Z(n43309) );
  XOR U42304 ( .A(n43312), .B(n43311), .Z(n43310) );
  NOR U42305 ( .A(n22579), .B(p_input[363]), .Z(n43311) );
  XOR U42306 ( .A(n43314), .B(n43313), .Z(n43312) );
  NOR U42307 ( .A(n22581), .B(p_input[361]), .Z(n43313) );
  XOR U42308 ( .A(n43316), .B(n43315), .Z(n43314) );
  NOR U42309 ( .A(n22583), .B(p_input[359]), .Z(n43315) );
  XOR U42310 ( .A(n43318), .B(n43317), .Z(n43316) );
  NOR U42311 ( .A(n22585), .B(p_input[357]), .Z(n43317) );
  XOR U42312 ( .A(n43320), .B(n43319), .Z(n43318) );
  NOR U42313 ( .A(n22587), .B(p_input[355]), .Z(n43319) );
  XOR U42314 ( .A(n43322), .B(n43321), .Z(n43320) );
  NOR U42315 ( .A(n22589), .B(p_input[353]), .Z(n43321) );
  XOR U42316 ( .A(n43324), .B(n43323), .Z(n43322) );
  NOR U42317 ( .A(n22591), .B(p_input[351]), .Z(n43323) );
  XOR U42318 ( .A(n43326), .B(n43325), .Z(n43324) );
  NOR U42319 ( .A(n22593), .B(p_input[349]), .Z(n43325) );
  XOR U42320 ( .A(n43328), .B(n43327), .Z(n43326) );
  NOR U42321 ( .A(n22595), .B(p_input[347]), .Z(n43327) );
  XOR U42322 ( .A(n43330), .B(n43329), .Z(n43328) );
  NOR U42323 ( .A(n22597), .B(p_input[345]), .Z(n43329) );
  XOR U42324 ( .A(n43332), .B(n43331), .Z(n43330) );
  NOR U42325 ( .A(n22599), .B(p_input[343]), .Z(n43331) );
  XOR U42326 ( .A(n43334), .B(n43333), .Z(n43332) );
  NOR U42327 ( .A(n22601), .B(p_input[341]), .Z(n43333) );
  XOR U42328 ( .A(n43336), .B(n43335), .Z(n43334) );
  NOR U42329 ( .A(n22603), .B(p_input[339]), .Z(n43335) );
  XOR U42330 ( .A(n43338), .B(n43337), .Z(n43336) );
  NOR U42331 ( .A(n22605), .B(p_input[337]), .Z(n43337) );
  XOR U42332 ( .A(n43340), .B(n43339), .Z(n43338) );
  NOR U42333 ( .A(n22607), .B(p_input[335]), .Z(n43339) );
  XOR U42334 ( .A(n43342), .B(n43341), .Z(n43340) );
  NOR U42335 ( .A(n22609), .B(p_input[333]), .Z(n43341) );
  XOR U42336 ( .A(n43344), .B(n43343), .Z(n43342) );
  NOR U42337 ( .A(n22611), .B(p_input[331]), .Z(n43343) );
  XOR U42338 ( .A(n43346), .B(n43345), .Z(n43344) );
  NOR U42339 ( .A(n22613), .B(p_input[329]), .Z(n43345) );
  XOR U42340 ( .A(n43348), .B(n43347), .Z(n43346) );
  NOR U42341 ( .A(n22615), .B(p_input[327]), .Z(n43347) );
  XOR U42342 ( .A(n43350), .B(n43349), .Z(n43348) );
  NOR U42343 ( .A(n22617), .B(p_input[325]), .Z(n43349) );
  XOR U42344 ( .A(n43352), .B(n43351), .Z(n43350) );
  NOR U42345 ( .A(n22619), .B(p_input[323]), .Z(n43351) );
  XOR U42346 ( .A(n43354), .B(n43353), .Z(n43352) );
  NOR U42347 ( .A(n22621), .B(p_input[321]), .Z(n43353) );
  XOR U42348 ( .A(n43356), .B(n43355), .Z(n43354) );
  NOR U42349 ( .A(n22623), .B(p_input[319]), .Z(n43355) );
  XOR U42350 ( .A(n43358), .B(n43357), .Z(n43356) );
  NOR U42351 ( .A(n22625), .B(p_input[317]), .Z(n43357) );
  XOR U42352 ( .A(n43360), .B(n43359), .Z(n43358) );
  NOR U42353 ( .A(n22627), .B(p_input[315]), .Z(n43359) );
  XOR U42354 ( .A(n43362), .B(n43361), .Z(n43360) );
  NOR U42355 ( .A(n22629), .B(p_input[313]), .Z(n43361) );
  XOR U42356 ( .A(n43364), .B(n43363), .Z(n43362) );
  NOR U42357 ( .A(n22631), .B(p_input[311]), .Z(n43363) );
  XOR U42358 ( .A(n43366), .B(n43365), .Z(n43364) );
  NOR U42359 ( .A(n22633), .B(p_input[309]), .Z(n43365) );
  XOR U42360 ( .A(n43368), .B(n43367), .Z(n43366) );
  NOR U42361 ( .A(n22635), .B(p_input[307]), .Z(n43367) );
  XOR U42362 ( .A(n43370), .B(n43369), .Z(n43368) );
  NOR U42363 ( .A(n22637), .B(p_input[305]), .Z(n43369) );
  XOR U42364 ( .A(n43372), .B(n43371), .Z(n43370) );
  NOR U42365 ( .A(n22639), .B(p_input[303]), .Z(n43371) );
  XOR U42366 ( .A(n43374), .B(n43373), .Z(n43372) );
  NOR U42367 ( .A(n22641), .B(p_input[301]), .Z(n43373) );
  XOR U42368 ( .A(n43376), .B(n43375), .Z(n43374) );
  NOR U42369 ( .A(n22643), .B(p_input[299]), .Z(n43375) );
  XOR U42370 ( .A(n43378), .B(n43377), .Z(n43376) );
  NOR U42371 ( .A(n22645), .B(p_input[297]), .Z(n43377) );
  XOR U42372 ( .A(n43380), .B(n43379), .Z(n43378) );
  NOR U42373 ( .A(n22647), .B(p_input[295]), .Z(n43379) );
  XOR U42374 ( .A(n43382), .B(n43381), .Z(n43380) );
  NOR U42375 ( .A(n22649), .B(p_input[293]), .Z(n43381) );
  XOR U42376 ( .A(n43384), .B(n43383), .Z(n43382) );
  NOR U42377 ( .A(n22651), .B(p_input[291]), .Z(n43383) );
  XOR U42378 ( .A(n43386), .B(n43385), .Z(n43384) );
  NOR U42379 ( .A(n22653), .B(p_input[289]), .Z(n43385) );
  XOR U42380 ( .A(n43388), .B(n43387), .Z(n43386) );
  NOR U42381 ( .A(n22655), .B(p_input[287]), .Z(n43387) );
  XOR U42382 ( .A(n43390), .B(n43389), .Z(n43388) );
  NOR U42383 ( .A(n22657), .B(p_input[285]), .Z(n43389) );
  XOR U42384 ( .A(n43392), .B(n43391), .Z(n43390) );
  NOR U42385 ( .A(n22659), .B(p_input[283]), .Z(n43391) );
  XOR U42386 ( .A(n43394), .B(n43393), .Z(n43392) );
  NOR U42387 ( .A(n22661), .B(p_input[281]), .Z(n43393) );
  XOR U42388 ( .A(n43396), .B(n43395), .Z(n43394) );
  NOR U42389 ( .A(n22663), .B(p_input[279]), .Z(n43395) );
  XOR U42390 ( .A(n43398), .B(n43397), .Z(n43396) );
  NOR U42391 ( .A(n22665), .B(p_input[277]), .Z(n43397) );
  XOR U42392 ( .A(n43400), .B(n43399), .Z(n43398) );
  NOR U42393 ( .A(n22667), .B(p_input[275]), .Z(n43399) );
  XOR U42394 ( .A(n43402), .B(n43401), .Z(n43400) );
  NOR U42395 ( .A(n22669), .B(p_input[273]), .Z(n43401) );
  XOR U42396 ( .A(n43404), .B(n43403), .Z(n43402) );
  NOR U42397 ( .A(n22671), .B(p_input[271]), .Z(n43403) );
  XOR U42398 ( .A(n43406), .B(n43405), .Z(n43404) );
  NOR U42399 ( .A(n22673), .B(p_input[269]), .Z(n43405) );
  XOR U42400 ( .A(n43408), .B(n43407), .Z(n43406) );
  NOR U42401 ( .A(n22675), .B(p_input[267]), .Z(n43407) );
  XOR U42402 ( .A(n43410), .B(n43409), .Z(n43408) );
  NOR U42403 ( .A(n22677), .B(p_input[265]), .Z(n43409) );
  XOR U42404 ( .A(n43412), .B(n43411), .Z(n43410) );
  NOR U42405 ( .A(n22679), .B(p_input[263]), .Z(n43411) );
  XOR U42406 ( .A(n43414), .B(n43413), .Z(n43412) );
  NOR U42407 ( .A(n22681), .B(p_input[261]), .Z(n43413) );
  XOR U42408 ( .A(n43416), .B(n43415), .Z(n43414) );
  NOR U42409 ( .A(n22683), .B(p_input[259]), .Z(n43415) );
  XOR U42410 ( .A(n43418), .B(n43417), .Z(n43416) );
  NOR U42411 ( .A(n22685), .B(p_input[257]), .Z(n43417) );
  XOR U42412 ( .A(n43420), .B(n43419), .Z(n43418) );
  NOR U42413 ( .A(n22687), .B(p_input[255]), .Z(n43419) );
  XOR U42414 ( .A(n43424), .B(n43423), .Z(n43420) );
  NOR U42415 ( .A(n22689), .B(p_input[253]), .Z(n43423) );
  XOR U42416 ( .A(n43426), .B(n43425), .Z(n43424) );
  NOR U42417 ( .A(n22691), .B(p_input[251]), .Z(n43425) );
  XOR U42418 ( .A(n43428), .B(n43427), .Z(n43426) );
  NOR U42419 ( .A(n22693), .B(p_input[249]), .Z(n43427) );
  XOR U42420 ( .A(n43430), .B(n43429), .Z(n43428) );
  NOR U42421 ( .A(n22695), .B(p_input[247]), .Z(n43429) );
  XOR U42422 ( .A(n43432), .B(n43431), .Z(n43430) );
  NOR U42423 ( .A(n22697), .B(p_input[245]), .Z(n43431) );
  XOR U42424 ( .A(n43434), .B(n43433), .Z(n43432) );
  NOR U42425 ( .A(n22699), .B(p_input[243]), .Z(n43433) );
  XOR U42426 ( .A(n43436), .B(n43435), .Z(n43434) );
  NOR U42427 ( .A(n22701), .B(p_input[241]), .Z(n43435) );
  XOR U42428 ( .A(n43438), .B(n43437), .Z(n43436) );
  NOR U42429 ( .A(n22703), .B(p_input[239]), .Z(n43437) );
  XOR U42430 ( .A(n43440), .B(n43439), .Z(n43438) );
  NOR U42431 ( .A(n22705), .B(p_input[237]), .Z(n43439) );
  XOR U42432 ( .A(n43442), .B(n43441), .Z(n43440) );
  NOR U42433 ( .A(n22707), .B(p_input[235]), .Z(n43441) );
  XOR U42434 ( .A(n43444), .B(n43443), .Z(n43442) );
  NOR U42435 ( .A(n22709), .B(p_input[233]), .Z(n43443) );
  XOR U42436 ( .A(n43446), .B(n43445), .Z(n43444) );
  NOR U42437 ( .A(n22711), .B(p_input[231]), .Z(n43445) );
  XOR U42438 ( .A(n43448), .B(n43447), .Z(n43446) );
  NOR U42439 ( .A(n22713), .B(p_input[229]), .Z(n43447) );
  XOR U42440 ( .A(n43450), .B(n43449), .Z(n43448) );
  NOR U42441 ( .A(n22715), .B(p_input[227]), .Z(n43449) );
  XOR U42442 ( .A(n43452), .B(n43451), .Z(n43450) );
  NOR U42443 ( .A(n22717), .B(p_input[225]), .Z(n43451) );
  XOR U42444 ( .A(n43454), .B(n43453), .Z(n43452) );
  NOR U42445 ( .A(n22719), .B(p_input[223]), .Z(n43453) );
  XOR U42446 ( .A(n43456), .B(n43455), .Z(n43454) );
  NOR U42447 ( .A(n22721), .B(p_input[221]), .Z(n43455) );
  XOR U42448 ( .A(n43458), .B(n43457), .Z(n43456) );
  NOR U42449 ( .A(n22723), .B(p_input[219]), .Z(n43457) );
  XOR U42450 ( .A(n43460), .B(n43459), .Z(n43458) );
  NOR U42451 ( .A(n22725), .B(p_input[217]), .Z(n43459) );
  XOR U42452 ( .A(n43462), .B(n43461), .Z(n43460) );
  NOR U42453 ( .A(n22727), .B(p_input[215]), .Z(n43461) );
  XOR U42454 ( .A(n43464), .B(n43463), .Z(n43462) );
  NOR U42455 ( .A(n22729), .B(p_input[213]), .Z(n43463) );
  XOR U42456 ( .A(n43466), .B(n43465), .Z(n43464) );
  NOR U42457 ( .A(n22731), .B(p_input[211]), .Z(n43465) );
  XOR U42458 ( .A(n43468), .B(n43467), .Z(n43466) );
  NOR U42459 ( .A(n22733), .B(p_input[209]), .Z(n43467) );
  XOR U42460 ( .A(n43470), .B(n43469), .Z(n43468) );
  NOR U42461 ( .A(n22735), .B(p_input[207]), .Z(n43469) );
  XOR U42462 ( .A(n43472), .B(n43471), .Z(n43470) );
  NOR U42463 ( .A(n22737), .B(p_input[205]), .Z(n43471) );
  XOR U42464 ( .A(n43474), .B(n43473), .Z(n43472) );
  NOR U42465 ( .A(n22739), .B(p_input[203]), .Z(n43473) );
  XOR U42466 ( .A(n43476), .B(n43475), .Z(n43474) );
  NOR U42467 ( .A(n22741), .B(p_input[201]), .Z(n43475) );
  XOR U42468 ( .A(n43478), .B(n43477), .Z(n43476) );
  NOR U42469 ( .A(n22743), .B(p_input[199]), .Z(n43477) );
  XOR U42470 ( .A(n43480), .B(n43479), .Z(n43478) );
  NOR U42471 ( .A(n22745), .B(p_input[197]), .Z(n43479) );
  XOR U42472 ( .A(n43482), .B(n43481), .Z(n43480) );
  NOR U42473 ( .A(n22747), .B(p_input[195]), .Z(n43481) );
  XOR U42474 ( .A(n43484), .B(n43483), .Z(n43482) );
  NOR U42475 ( .A(n22749), .B(p_input[193]), .Z(n43483) );
  XOR U42476 ( .A(n43486), .B(n43485), .Z(n43484) );
  NOR U42477 ( .A(n22751), .B(p_input[191]), .Z(n43485) );
  XOR U42478 ( .A(n43488), .B(n43487), .Z(n43486) );
  NOR U42479 ( .A(n22753), .B(p_input[189]), .Z(n43487) );
  XOR U42480 ( .A(n43490), .B(n43489), .Z(n43488) );
  NOR U42481 ( .A(n22755), .B(p_input[187]), .Z(n43489) );
  XOR U42482 ( .A(n43492), .B(n43491), .Z(n43490) );
  NOR U42483 ( .A(n22757), .B(p_input[185]), .Z(n43491) );
  XOR U42484 ( .A(n43494), .B(n43493), .Z(n43492) );
  NOR U42485 ( .A(n22759), .B(p_input[183]), .Z(n43493) );
  XOR U42486 ( .A(n43496), .B(n43495), .Z(n43494) );
  NOR U42487 ( .A(n22761), .B(p_input[181]), .Z(n43495) );
  XOR U42488 ( .A(n43498), .B(n43497), .Z(n43496) );
  NOR U42489 ( .A(n22763), .B(p_input[179]), .Z(n43497) );
  XOR U42490 ( .A(n43500), .B(n43499), .Z(n43498) );
  NOR U42491 ( .A(n22765), .B(p_input[177]), .Z(n43499) );
  XOR U42492 ( .A(n43502), .B(n43501), .Z(n43500) );
  NOR U42493 ( .A(n22767), .B(p_input[175]), .Z(n43501) );
  XOR U42494 ( .A(n43504), .B(n43503), .Z(n43502) );
  NOR U42495 ( .A(n22769), .B(p_input[173]), .Z(n43503) );
  XOR U42496 ( .A(n43506), .B(n43505), .Z(n43504) );
  NOR U42497 ( .A(n22771), .B(p_input[171]), .Z(n43505) );
  XOR U42498 ( .A(n43508), .B(n43507), .Z(n43506) );
  NOR U42499 ( .A(n22773), .B(p_input[169]), .Z(n43507) );
  XOR U42500 ( .A(n43510), .B(n43509), .Z(n43508) );
  NOR U42501 ( .A(n22775), .B(p_input[167]), .Z(n43509) );
  XOR U42502 ( .A(n43512), .B(n43511), .Z(n43510) );
  NOR U42503 ( .A(n22777), .B(p_input[165]), .Z(n43511) );
  XOR U42504 ( .A(n43514), .B(n43513), .Z(n43512) );
  NOR U42505 ( .A(n22779), .B(p_input[163]), .Z(n43513) );
  XOR U42506 ( .A(n43516), .B(n43515), .Z(n43514) );
  NOR U42507 ( .A(n22781), .B(p_input[161]), .Z(n43515) );
  XOR U42508 ( .A(n43518), .B(n43517), .Z(n43516) );
  NOR U42509 ( .A(n22783), .B(p_input[159]), .Z(n43517) );
  XOR U42510 ( .A(n43520), .B(n43519), .Z(n43518) );
  NOR U42511 ( .A(n22785), .B(p_input[157]), .Z(n43519) );
  XOR U42512 ( .A(n43522), .B(n43521), .Z(n43520) );
  NOR U42513 ( .A(n22787), .B(p_input[155]), .Z(n43521) );
  XOR U42514 ( .A(n43524), .B(n43523), .Z(n43522) );
  NOR U42515 ( .A(n22789), .B(p_input[153]), .Z(n43523) );
  XOR U42516 ( .A(n43526), .B(n43525), .Z(n43524) );
  NOR U42517 ( .A(n22791), .B(p_input[151]), .Z(n43525) );
  XOR U42518 ( .A(n43528), .B(n43527), .Z(n43526) );
  NOR U42519 ( .A(n22793), .B(p_input[149]), .Z(n43527) );
  XOR U42520 ( .A(n43530), .B(n43529), .Z(n43528) );
  NOR U42521 ( .A(n22795), .B(p_input[147]), .Z(n43529) );
  XOR U42522 ( .A(n43532), .B(n43531), .Z(n43530) );
  NOR U42523 ( .A(n22797), .B(p_input[145]), .Z(n43531) );
  XOR U42524 ( .A(n43534), .B(n43533), .Z(n43532) );
  NOR U42525 ( .A(n22799), .B(p_input[143]), .Z(n43533) );
  XOR U42526 ( .A(n43536), .B(n43535), .Z(n43534) );
  NOR U42527 ( .A(n22801), .B(p_input[141]), .Z(n43535) );
  XOR U42528 ( .A(n43538), .B(n43537), .Z(n43536) );
  NOR U42529 ( .A(n22803), .B(p_input[139]), .Z(n43537) );
  XOR U42530 ( .A(n43540), .B(n43539), .Z(n43538) );
  NOR U42531 ( .A(n22805), .B(p_input[137]), .Z(n43539) );
  XOR U42532 ( .A(n43542), .B(n43541), .Z(n43540) );
  NOR U42533 ( .A(n22807), .B(p_input[135]), .Z(n43541) );
  XOR U42534 ( .A(n43544), .B(n43543), .Z(n43542) );
  NOR U42535 ( .A(n22809), .B(p_input[133]), .Z(n43543) );
  XOR U42536 ( .A(n43546), .B(n43545), .Z(n43544) );
  NOR U42537 ( .A(n22811), .B(p_input[131]), .Z(n43545) );
  XOR U42538 ( .A(n43548), .B(n43547), .Z(n43546) );
  NOR U42539 ( .A(n22813), .B(p_input[129]), .Z(n43547) );
  XOR U42540 ( .A(n43550), .B(n43549), .Z(n43548) );
  NOR U42541 ( .A(n22815), .B(p_input[127]), .Z(n43549) );
  XOR U42542 ( .A(n43552), .B(n43551), .Z(n43550) );
  NOR U42543 ( .A(n22817), .B(p_input[125]), .Z(n43551) );
  XOR U42544 ( .A(n43554), .B(n43553), .Z(n43552) );
  NOR U42545 ( .A(n22819), .B(p_input[123]), .Z(n43553) );
  XOR U42546 ( .A(n43556), .B(n43555), .Z(n43554) );
  NOR U42547 ( .A(n22821), .B(p_input[121]), .Z(n43555) );
  XOR U42548 ( .A(n43558), .B(n43557), .Z(n43556) );
  NOR U42549 ( .A(n22823), .B(p_input[119]), .Z(n43557) );
  XOR U42550 ( .A(n43560), .B(n43559), .Z(n43558) );
  NOR U42551 ( .A(n22825), .B(p_input[117]), .Z(n43559) );
  XOR U42552 ( .A(n43562), .B(n43561), .Z(n43560) );
  NOR U42553 ( .A(n22827), .B(p_input[115]), .Z(n43561) );
  XOR U42554 ( .A(n43564), .B(n43563), .Z(n43562) );
  NOR U42555 ( .A(n22829), .B(p_input[113]), .Z(n43563) );
  XOR U42556 ( .A(n43566), .B(n43565), .Z(n43564) );
  NOR U42557 ( .A(n22831), .B(p_input[111]), .Z(n43565) );
  XOR U42558 ( .A(n43568), .B(n43567), .Z(n43566) );
  NOR U42559 ( .A(n22833), .B(p_input[109]), .Z(n43567) );
  XOR U42560 ( .A(n43570), .B(n43569), .Z(n43568) );
  NOR U42561 ( .A(n22835), .B(p_input[107]), .Z(n43569) );
  XOR U42562 ( .A(n43572), .B(n43571), .Z(n43570) );
  NOR U42563 ( .A(n22837), .B(p_input[105]), .Z(n43571) );
  XOR U42564 ( .A(n43574), .B(n43573), .Z(n43572) );
  NOR U42565 ( .A(n22839), .B(p_input[103]), .Z(n43573) );
  XOR U42566 ( .A(n43576), .B(n43575), .Z(n43574) );
  NOR U42567 ( .A(n22841), .B(p_input[101]), .Z(n43575) );
  XOR U42568 ( .A(n43578), .B(n43577), .Z(n43576) );
  NOR U42569 ( .A(n22843), .B(p_input[99]), .Z(n43577) );
  XOR U42570 ( .A(n43580), .B(n43579), .Z(n43578) );
  NOR U42571 ( .A(n22845), .B(p_input[97]), .Z(n43579) );
  XOR U42572 ( .A(n43582), .B(n43581), .Z(n43580) );
  NOR U42573 ( .A(n22847), .B(p_input[95]), .Z(n43581) );
  XOR U42574 ( .A(n43584), .B(n43583), .Z(n43582) );
  NOR U42575 ( .A(n22849), .B(p_input[93]), .Z(n43583) );
  XOR U42576 ( .A(n43586), .B(n43585), .Z(n43584) );
  NOR U42577 ( .A(n22851), .B(p_input[91]), .Z(n43585) );
  XOR U42578 ( .A(n43588), .B(n43587), .Z(n43586) );
  NOR U42579 ( .A(n22853), .B(p_input[89]), .Z(n43587) );
  XOR U42580 ( .A(n43590), .B(n43589), .Z(n43588) );
  NOR U42581 ( .A(n22855), .B(p_input[87]), .Z(n43589) );
  XOR U42582 ( .A(n43592), .B(n43591), .Z(n43590) );
  NOR U42583 ( .A(n22857), .B(p_input[85]), .Z(n43591) );
  XOR U42584 ( .A(n43594), .B(n43593), .Z(n43592) );
  NOR U42585 ( .A(n22859), .B(p_input[83]), .Z(n43593) );
  XOR U42586 ( .A(n43596), .B(n43595), .Z(n43594) );
  NOR U42587 ( .A(n22861), .B(p_input[81]), .Z(n43595) );
  XOR U42588 ( .A(n43598), .B(n43597), .Z(n43596) );
  NOR U42589 ( .A(n22863), .B(p_input[79]), .Z(n43597) );
  XOR U42590 ( .A(n43600), .B(n43599), .Z(n43598) );
  NOR U42591 ( .A(n22865), .B(p_input[77]), .Z(n43599) );
  XOR U42592 ( .A(n43602), .B(n43601), .Z(n43600) );
  NOR U42593 ( .A(n22867), .B(p_input[75]), .Z(n43601) );
  XOR U42594 ( .A(n43604), .B(n43603), .Z(n43602) );
  NOR U42595 ( .A(n22869), .B(p_input[73]), .Z(n43603) );
  XOR U42596 ( .A(n43606), .B(n43605), .Z(n43604) );
  NOR U42597 ( .A(n22871), .B(p_input[71]), .Z(n43605) );
  XOR U42598 ( .A(n43608), .B(n43607), .Z(n43606) );
  NOR U42599 ( .A(n22873), .B(p_input[69]), .Z(n43607) );
  XOR U42600 ( .A(n43610), .B(n43609), .Z(n43608) );
  NOR U42601 ( .A(n22875), .B(p_input[67]), .Z(n43609) );
  XOR U42602 ( .A(n43612), .B(n43611), .Z(n43610) );
  NOR U42603 ( .A(n22877), .B(p_input[65]), .Z(n43611) );
  XOR U42604 ( .A(n43614), .B(n43613), .Z(n43612) );
  NOR U42605 ( .A(n22879), .B(p_input[63]), .Z(n43613) );
  XOR U42606 ( .A(n43616), .B(n43615), .Z(n43614) );
  NOR U42607 ( .A(n22881), .B(p_input[61]), .Z(n43615) );
  XOR U42608 ( .A(n43618), .B(n43617), .Z(n43616) );
  NOR U42609 ( .A(n22883), .B(p_input[59]), .Z(n43617) );
  XOR U42610 ( .A(n43620), .B(n43619), .Z(n43618) );
  NOR U42611 ( .A(n22885), .B(p_input[57]), .Z(n43619) );
  XOR U42612 ( .A(n43622), .B(n43621), .Z(n43620) );
  NOR U42613 ( .A(n22887), .B(p_input[55]), .Z(n43621) );
  XOR U42614 ( .A(n43624), .B(n43623), .Z(n43622) );
  NOR U42615 ( .A(n22889), .B(p_input[53]), .Z(n43623) );
  XOR U42616 ( .A(n43626), .B(n43625), .Z(n43624) );
  NOR U42617 ( .A(n22891), .B(p_input[51]), .Z(n43625) );
  XOR U42618 ( .A(n43628), .B(n43627), .Z(n43626) );
  NOR U42619 ( .A(n22893), .B(p_input[49]), .Z(n43627) );
  XOR U42620 ( .A(n43630), .B(n43629), .Z(n43628) );
  NOR U42621 ( .A(n22895), .B(p_input[47]), .Z(n43629) );
  XOR U42622 ( .A(n43632), .B(n43631), .Z(n43630) );
  NOR U42623 ( .A(n22897), .B(p_input[45]), .Z(n43631) );
  XOR U42624 ( .A(n43634), .B(n43633), .Z(n43632) );
  NOR U42625 ( .A(n22899), .B(p_input[43]), .Z(n43633) );
  XOR U42626 ( .A(n43636), .B(n43635), .Z(n43634) );
  NOR U42627 ( .A(n22901), .B(p_input[41]), .Z(n43635) );
  XOR U42628 ( .A(n43638), .B(n43637), .Z(n43636) );
  NOR U42629 ( .A(n22903), .B(p_input[39]), .Z(n43637) );
  XOR U42630 ( .A(n43640), .B(n43639), .Z(n43638) );
  NOR U42631 ( .A(n22905), .B(p_input[37]), .Z(n43639) );
  XOR U42632 ( .A(n43642), .B(n43641), .Z(n43640) );
  NOR U42633 ( .A(n22907), .B(p_input[35]), .Z(n43641) );
  XOR U42634 ( .A(n43644), .B(n43643), .Z(n43642) );
  NOR U42635 ( .A(n22909), .B(p_input[33]), .Z(n43643) );
  XOR U42636 ( .A(n43646), .B(n43645), .Z(n43644) );
  NOR U42637 ( .A(n22911), .B(p_input[31]), .Z(n43645) );
  XOR U42638 ( .A(n43648), .B(n43647), .Z(n43646) );
  NOR U42639 ( .A(n22913), .B(p_input[29]), .Z(n43647) );
  XOR U42640 ( .A(n43650), .B(n43649), .Z(n43648) );
  NOR U42641 ( .A(n22915), .B(p_input[27]), .Z(n43649) );
  XOR U42642 ( .A(n43652), .B(n43651), .Z(n43650) );
  NOR U42643 ( .A(n22917), .B(p_input[25]), .Z(n43651) );
  XOR U42644 ( .A(n43654), .B(n43653), .Z(n43652) );
  NOR U42645 ( .A(n22919), .B(p_input[23]), .Z(n43653) );
  XOR U42646 ( .A(n43656), .B(n43655), .Z(n43654) );
  NOR U42647 ( .A(n22921), .B(p_input[21]), .Z(n43655) );
  XOR U42648 ( .A(n43658), .B(n43657), .Z(n43656) );
  NOR U42649 ( .A(n22923), .B(p_input[19]), .Z(n43657) );
  XOR U42650 ( .A(n43660), .B(n43659), .Z(n43658) );
  NOR U42651 ( .A(n22925), .B(p_input[17]), .Z(n43659) );
  XOR U42652 ( .A(n43662), .B(n43661), .Z(n43660) );
  NOR U42653 ( .A(n22927), .B(p_input[15]), .Z(n43661) );
  XOR U42654 ( .A(n43664), .B(n43663), .Z(n43662) );
  NOR U42655 ( .A(n22929), .B(p_input[13]), .Z(n43663) );
  XOR U42656 ( .A(n43678), .B(n43677), .Z(n43664) );
  NOR U42657 ( .A(n22931), .B(p_input[11]), .Z(n43677) );
  XOR U42658 ( .A(n43680), .B(n43679), .Z(n43678) );
  NOR U42659 ( .A(n22933), .B(p_input[9]), .Z(n43679) );
  XOR U42660 ( .A(n43668), .B(n43667), .Z(n43680) );
  NOR U42661 ( .A(n22935), .B(p_input[7]), .Z(n43667) );
  XOR U42662 ( .A(n43675), .B(n43676), .Z(n43668) );
  XOR U42663 ( .A(n43673), .B(n43674), .Z(n43676) );
  NOR U42664 ( .A(n22937), .B(p_input[3]), .Z(n43674) );
  NOR U42665 ( .A(n22939), .B(p_input[1]), .Z(n43673) );
  NOR U42666 ( .A(n22941), .B(p_input[5]), .Z(n43675) );
  XOR U42667 ( .A(n43682), .B(n43681), .Z(n22942) );
  AND U42668 ( .A(n21918), .B(n21919), .Z(n43681) );
  IV U42669 ( .A(p_input[1022]), .Z(n21919) );
  IV U42670 ( .A(p_input[1023]), .Z(n21918) );
  XOR U42671 ( .A(n43684), .B(n43683), .Z(n43682) );
  AND U42672 ( .A(n21920), .B(n21921), .Z(n43683) );
  IV U42673 ( .A(p_input[1020]), .Z(n21921) );
  IV U42674 ( .A(p_input[1021]), .Z(n21920) );
  XOR U42675 ( .A(n43686), .B(n43685), .Z(n43684) );
  AND U42676 ( .A(n21922), .B(n21923), .Z(n43685) );
  IV U42677 ( .A(p_input[1018]), .Z(n21923) );
  IV U42678 ( .A(p_input[1019]), .Z(n21922) );
  XOR U42679 ( .A(n43688), .B(n43687), .Z(n43686) );
  AND U42680 ( .A(n21924), .B(n21925), .Z(n43687) );
  IV U42681 ( .A(p_input[1016]), .Z(n21925) );
  IV U42682 ( .A(p_input[1017]), .Z(n21924) );
  XOR U42683 ( .A(n43690), .B(n43689), .Z(n43688) );
  AND U42684 ( .A(n21926), .B(n21927), .Z(n43689) );
  IV U42685 ( .A(p_input[1014]), .Z(n21927) );
  IV U42686 ( .A(p_input[1015]), .Z(n21926) );
  XOR U42687 ( .A(n43692), .B(n43691), .Z(n43690) );
  AND U42688 ( .A(n21928), .B(n21929), .Z(n43691) );
  IV U42689 ( .A(p_input[1012]), .Z(n21929) );
  IV U42690 ( .A(p_input[1013]), .Z(n21928) );
  XOR U42691 ( .A(n43694), .B(n43693), .Z(n43692) );
  AND U42692 ( .A(n21930), .B(n21931), .Z(n43693) );
  IV U42693 ( .A(p_input[1010]), .Z(n21931) );
  IV U42694 ( .A(p_input[1011]), .Z(n21930) );
  XOR U42695 ( .A(n43696), .B(n43695), .Z(n43694) );
  AND U42696 ( .A(n21932), .B(n21933), .Z(n43695) );
  IV U42697 ( .A(p_input[1008]), .Z(n21933) );
  IV U42698 ( .A(p_input[1009]), .Z(n21932) );
  XOR U42699 ( .A(n43698), .B(n43697), .Z(n43696) );
  AND U42700 ( .A(n21934), .B(n21935), .Z(n43697) );
  IV U42701 ( .A(p_input[1006]), .Z(n21935) );
  IV U42702 ( .A(p_input[1007]), .Z(n21934) );
  XOR U42703 ( .A(n43700), .B(n43699), .Z(n43698) );
  AND U42704 ( .A(n21936), .B(n21937), .Z(n43699) );
  IV U42705 ( .A(p_input[1004]), .Z(n21937) );
  IV U42706 ( .A(p_input[1005]), .Z(n21936) );
  XOR U42707 ( .A(n43702), .B(n43701), .Z(n43700) );
  AND U42708 ( .A(n21938), .B(n21939), .Z(n43701) );
  IV U42709 ( .A(p_input[1002]), .Z(n21939) );
  IV U42710 ( .A(p_input[1003]), .Z(n21938) );
  XOR U42711 ( .A(n43704), .B(n43703), .Z(n43702) );
  AND U42712 ( .A(n21940), .B(n21941), .Z(n43703) );
  IV U42713 ( .A(p_input[1000]), .Z(n21941) );
  IV U42714 ( .A(p_input[1001]), .Z(n21940) );
  XOR U42715 ( .A(n43706), .B(n43705), .Z(n43704) );
  AND U42716 ( .A(n21942), .B(n21943), .Z(n43705) );
  IV U42717 ( .A(p_input[998]), .Z(n21943) );
  IV U42718 ( .A(p_input[999]), .Z(n21942) );
  XOR U42719 ( .A(n43708), .B(n43707), .Z(n43706) );
  AND U42720 ( .A(n21944), .B(n21945), .Z(n43707) );
  IV U42721 ( .A(p_input[996]), .Z(n21945) );
  IV U42722 ( .A(p_input[997]), .Z(n21944) );
  XOR U42723 ( .A(n43710), .B(n43709), .Z(n43708) );
  AND U42724 ( .A(n21946), .B(n21947), .Z(n43709) );
  IV U42725 ( .A(p_input[994]), .Z(n21947) );
  IV U42726 ( .A(p_input[995]), .Z(n21946) );
  XOR U42727 ( .A(n43712), .B(n43711), .Z(n43710) );
  AND U42728 ( .A(n21948), .B(n21949), .Z(n43711) );
  IV U42729 ( .A(p_input[992]), .Z(n21949) );
  IV U42730 ( .A(p_input[993]), .Z(n21948) );
  XOR U42731 ( .A(n43714), .B(n43713), .Z(n43712) );
  AND U42732 ( .A(n21950), .B(n21951), .Z(n43713) );
  IV U42733 ( .A(p_input[990]), .Z(n21951) );
  IV U42734 ( .A(p_input[991]), .Z(n21950) );
  XOR U42735 ( .A(n43716), .B(n43715), .Z(n43714) );
  AND U42736 ( .A(n21952), .B(n21953), .Z(n43715) );
  IV U42737 ( .A(p_input[988]), .Z(n21953) );
  IV U42738 ( .A(p_input[989]), .Z(n21952) );
  XOR U42739 ( .A(n43718), .B(n43717), .Z(n43716) );
  AND U42740 ( .A(n21954), .B(n21955), .Z(n43717) );
  IV U42741 ( .A(p_input[986]), .Z(n21955) );
  IV U42742 ( .A(p_input[987]), .Z(n21954) );
  XOR U42743 ( .A(n43720), .B(n43719), .Z(n43718) );
  AND U42744 ( .A(n21956), .B(n21957), .Z(n43719) );
  IV U42745 ( .A(p_input[984]), .Z(n21957) );
  IV U42746 ( .A(p_input[985]), .Z(n21956) );
  XOR U42747 ( .A(n43722), .B(n43721), .Z(n43720) );
  AND U42748 ( .A(n21958), .B(n21959), .Z(n43721) );
  IV U42749 ( .A(p_input[982]), .Z(n21959) );
  IV U42750 ( .A(p_input[983]), .Z(n21958) );
  XOR U42751 ( .A(n43724), .B(n43723), .Z(n43722) );
  AND U42752 ( .A(n21960), .B(n21961), .Z(n43723) );
  IV U42753 ( .A(p_input[980]), .Z(n21961) );
  IV U42754 ( .A(p_input[981]), .Z(n21960) );
  XOR U42755 ( .A(n43726), .B(n43725), .Z(n43724) );
  AND U42756 ( .A(n21962), .B(n21963), .Z(n43725) );
  IV U42757 ( .A(p_input[978]), .Z(n21963) );
  IV U42758 ( .A(p_input[979]), .Z(n21962) );
  XOR U42759 ( .A(n43728), .B(n43727), .Z(n43726) );
  AND U42760 ( .A(n21964), .B(n21965), .Z(n43727) );
  IV U42761 ( .A(p_input[976]), .Z(n21965) );
  IV U42762 ( .A(p_input[977]), .Z(n21964) );
  XOR U42763 ( .A(n43730), .B(n43729), .Z(n43728) );
  AND U42764 ( .A(n21966), .B(n21967), .Z(n43729) );
  IV U42765 ( .A(p_input[974]), .Z(n21967) );
  IV U42766 ( .A(p_input[975]), .Z(n21966) );
  XOR U42767 ( .A(n43732), .B(n43731), .Z(n43730) );
  AND U42768 ( .A(n21968), .B(n21969), .Z(n43731) );
  IV U42769 ( .A(p_input[972]), .Z(n21969) );
  IV U42770 ( .A(p_input[973]), .Z(n21968) );
  XOR U42771 ( .A(n43734), .B(n43733), .Z(n43732) );
  AND U42772 ( .A(n21970), .B(n21971), .Z(n43733) );
  IV U42773 ( .A(p_input[970]), .Z(n21971) );
  IV U42774 ( .A(p_input[971]), .Z(n21970) );
  XOR U42775 ( .A(n43736), .B(n43735), .Z(n43734) );
  AND U42776 ( .A(n21972), .B(n21973), .Z(n43735) );
  IV U42777 ( .A(p_input[968]), .Z(n21973) );
  IV U42778 ( .A(p_input[969]), .Z(n21972) );
  XOR U42779 ( .A(n43738), .B(n43737), .Z(n43736) );
  AND U42780 ( .A(n21974), .B(n21975), .Z(n43737) );
  IV U42781 ( .A(p_input[966]), .Z(n21975) );
  IV U42782 ( .A(p_input[967]), .Z(n21974) );
  XOR U42783 ( .A(n43740), .B(n43739), .Z(n43738) );
  AND U42784 ( .A(n21976), .B(n21977), .Z(n43739) );
  IV U42785 ( .A(p_input[964]), .Z(n21977) );
  IV U42786 ( .A(p_input[965]), .Z(n21976) );
  XOR U42787 ( .A(n43742), .B(n43741), .Z(n43740) );
  AND U42788 ( .A(n21978), .B(n21979), .Z(n43741) );
  IV U42789 ( .A(p_input[962]), .Z(n21979) );
  IV U42790 ( .A(p_input[963]), .Z(n21978) );
  XOR U42791 ( .A(n43744), .B(n43743), .Z(n43742) );
  AND U42792 ( .A(n21980), .B(n21981), .Z(n43743) );
  IV U42793 ( .A(p_input[960]), .Z(n21981) );
  IV U42794 ( .A(p_input[961]), .Z(n21980) );
  XOR U42795 ( .A(n43746), .B(n43745), .Z(n43744) );
  AND U42796 ( .A(n21982), .B(n21983), .Z(n43745) );
  IV U42797 ( .A(p_input[958]), .Z(n21983) );
  IV U42798 ( .A(p_input[959]), .Z(n21982) );
  XOR U42799 ( .A(n43748), .B(n43747), .Z(n43746) );
  AND U42800 ( .A(n21984), .B(n21985), .Z(n43747) );
  IV U42801 ( .A(p_input[956]), .Z(n21985) );
  IV U42802 ( .A(p_input[957]), .Z(n21984) );
  XOR U42803 ( .A(n43750), .B(n43749), .Z(n43748) );
  AND U42804 ( .A(n21986), .B(n21987), .Z(n43749) );
  IV U42805 ( .A(p_input[954]), .Z(n21987) );
  IV U42806 ( .A(p_input[955]), .Z(n21986) );
  XOR U42807 ( .A(n43752), .B(n43751), .Z(n43750) );
  AND U42808 ( .A(n21988), .B(n21989), .Z(n43751) );
  IV U42809 ( .A(p_input[952]), .Z(n21989) );
  IV U42810 ( .A(p_input[953]), .Z(n21988) );
  XOR U42811 ( .A(n43754), .B(n43753), .Z(n43752) );
  AND U42812 ( .A(n21990), .B(n21991), .Z(n43753) );
  IV U42813 ( .A(p_input[950]), .Z(n21991) );
  IV U42814 ( .A(p_input[951]), .Z(n21990) );
  XOR U42815 ( .A(n43756), .B(n43755), .Z(n43754) );
  AND U42816 ( .A(n21992), .B(n21993), .Z(n43755) );
  IV U42817 ( .A(p_input[948]), .Z(n21993) );
  IV U42818 ( .A(p_input[949]), .Z(n21992) );
  XOR U42819 ( .A(n43758), .B(n43757), .Z(n43756) );
  AND U42820 ( .A(n21994), .B(n21995), .Z(n43757) );
  IV U42821 ( .A(p_input[946]), .Z(n21995) );
  IV U42822 ( .A(p_input[947]), .Z(n21994) );
  XOR U42823 ( .A(n43760), .B(n43759), .Z(n43758) );
  AND U42824 ( .A(n21996), .B(n21997), .Z(n43759) );
  IV U42825 ( .A(p_input[944]), .Z(n21997) );
  IV U42826 ( .A(p_input[945]), .Z(n21996) );
  XOR U42827 ( .A(n43762), .B(n43761), .Z(n43760) );
  AND U42828 ( .A(n21998), .B(n21999), .Z(n43761) );
  IV U42829 ( .A(p_input[942]), .Z(n21999) );
  IV U42830 ( .A(p_input[943]), .Z(n21998) );
  XOR U42831 ( .A(n43764), .B(n43763), .Z(n43762) );
  AND U42832 ( .A(n22000), .B(n22001), .Z(n43763) );
  IV U42833 ( .A(p_input[940]), .Z(n22001) );
  IV U42834 ( .A(p_input[941]), .Z(n22000) );
  XOR U42835 ( .A(n43766), .B(n43765), .Z(n43764) );
  AND U42836 ( .A(n22002), .B(n22003), .Z(n43765) );
  IV U42837 ( .A(p_input[938]), .Z(n22003) );
  IV U42838 ( .A(p_input[939]), .Z(n22002) );
  XOR U42839 ( .A(n43768), .B(n43767), .Z(n43766) );
  AND U42840 ( .A(n22004), .B(n22005), .Z(n43767) );
  IV U42841 ( .A(p_input[936]), .Z(n22005) );
  IV U42842 ( .A(p_input[937]), .Z(n22004) );
  XOR U42843 ( .A(n43770), .B(n43769), .Z(n43768) );
  AND U42844 ( .A(n22006), .B(n22007), .Z(n43769) );
  IV U42845 ( .A(p_input[934]), .Z(n22007) );
  IV U42846 ( .A(p_input[935]), .Z(n22006) );
  XOR U42847 ( .A(n43772), .B(n43771), .Z(n43770) );
  AND U42848 ( .A(n22008), .B(n22009), .Z(n43771) );
  IV U42849 ( .A(p_input[932]), .Z(n22009) );
  IV U42850 ( .A(p_input[933]), .Z(n22008) );
  XOR U42851 ( .A(n43774), .B(n43773), .Z(n43772) );
  AND U42852 ( .A(n22010), .B(n22011), .Z(n43773) );
  IV U42853 ( .A(p_input[930]), .Z(n22011) );
  IV U42854 ( .A(p_input[931]), .Z(n22010) );
  XOR U42855 ( .A(n43776), .B(n43775), .Z(n43774) );
  AND U42856 ( .A(n22012), .B(n22013), .Z(n43775) );
  IV U42857 ( .A(p_input[928]), .Z(n22013) );
  IV U42858 ( .A(p_input[929]), .Z(n22012) );
  XOR U42859 ( .A(n43778), .B(n43777), .Z(n43776) );
  AND U42860 ( .A(n22014), .B(n22015), .Z(n43777) );
  IV U42861 ( .A(p_input[926]), .Z(n22015) );
  IV U42862 ( .A(p_input[927]), .Z(n22014) );
  XOR U42863 ( .A(n43780), .B(n43779), .Z(n43778) );
  AND U42864 ( .A(n22016), .B(n22017), .Z(n43779) );
  IV U42865 ( .A(p_input[924]), .Z(n22017) );
  IV U42866 ( .A(p_input[925]), .Z(n22016) );
  XOR U42867 ( .A(n43782), .B(n43781), .Z(n43780) );
  AND U42868 ( .A(n22018), .B(n22019), .Z(n43781) );
  IV U42869 ( .A(p_input[922]), .Z(n22019) );
  IV U42870 ( .A(p_input[923]), .Z(n22018) );
  XOR U42871 ( .A(n43784), .B(n43783), .Z(n43782) );
  AND U42872 ( .A(n22020), .B(n22021), .Z(n43783) );
  IV U42873 ( .A(p_input[920]), .Z(n22021) );
  IV U42874 ( .A(p_input[921]), .Z(n22020) );
  XOR U42875 ( .A(n43786), .B(n43785), .Z(n43784) );
  AND U42876 ( .A(n22022), .B(n22023), .Z(n43785) );
  IV U42877 ( .A(p_input[918]), .Z(n22023) );
  IV U42878 ( .A(p_input[919]), .Z(n22022) );
  XOR U42879 ( .A(n43788), .B(n43787), .Z(n43786) );
  AND U42880 ( .A(n22024), .B(n22025), .Z(n43787) );
  IV U42881 ( .A(p_input[916]), .Z(n22025) );
  IV U42882 ( .A(p_input[917]), .Z(n22024) );
  XOR U42883 ( .A(n43790), .B(n43789), .Z(n43788) );
  AND U42884 ( .A(n22026), .B(n22027), .Z(n43789) );
  IV U42885 ( .A(p_input[914]), .Z(n22027) );
  IV U42886 ( .A(p_input[915]), .Z(n22026) );
  XOR U42887 ( .A(n43792), .B(n43791), .Z(n43790) );
  AND U42888 ( .A(n22028), .B(n22029), .Z(n43791) );
  IV U42889 ( .A(p_input[912]), .Z(n22029) );
  IV U42890 ( .A(p_input[913]), .Z(n22028) );
  XOR U42891 ( .A(n43794), .B(n43793), .Z(n43792) );
  AND U42892 ( .A(n22030), .B(n22031), .Z(n43793) );
  IV U42893 ( .A(p_input[910]), .Z(n22031) );
  IV U42894 ( .A(p_input[911]), .Z(n22030) );
  XOR U42895 ( .A(n43796), .B(n43795), .Z(n43794) );
  AND U42896 ( .A(n22032), .B(n22033), .Z(n43795) );
  IV U42897 ( .A(p_input[908]), .Z(n22033) );
  IV U42898 ( .A(p_input[909]), .Z(n22032) );
  XOR U42899 ( .A(n43798), .B(n43797), .Z(n43796) );
  AND U42900 ( .A(n22034), .B(n22035), .Z(n43797) );
  IV U42901 ( .A(p_input[906]), .Z(n22035) );
  IV U42902 ( .A(p_input[907]), .Z(n22034) );
  XOR U42903 ( .A(n43800), .B(n43799), .Z(n43798) );
  AND U42904 ( .A(n22036), .B(n22037), .Z(n43799) );
  IV U42905 ( .A(p_input[904]), .Z(n22037) );
  IV U42906 ( .A(p_input[905]), .Z(n22036) );
  XOR U42907 ( .A(n43802), .B(n43801), .Z(n43800) );
  AND U42908 ( .A(n22038), .B(n22039), .Z(n43801) );
  IV U42909 ( .A(p_input[902]), .Z(n22039) );
  IV U42910 ( .A(p_input[903]), .Z(n22038) );
  XOR U42911 ( .A(n43804), .B(n43803), .Z(n43802) );
  AND U42912 ( .A(n22040), .B(n22041), .Z(n43803) );
  IV U42913 ( .A(p_input[900]), .Z(n22041) );
  IV U42914 ( .A(p_input[901]), .Z(n22040) );
  XOR U42915 ( .A(n43806), .B(n43805), .Z(n43804) );
  AND U42916 ( .A(n22042), .B(n22043), .Z(n43805) );
  IV U42917 ( .A(p_input[898]), .Z(n22043) );
  IV U42918 ( .A(p_input[899]), .Z(n22042) );
  XOR U42919 ( .A(n43808), .B(n43807), .Z(n43806) );
  AND U42920 ( .A(n22044), .B(n22045), .Z(n43807) );
  IV U42921 ( .A(p_input[896]), .Z(n22045) );
  IV U42922 ( .A(p_input[897]), .Z(n22044) );
  XOR U42923 ( .A(n43810), .B(n43809), .Z(n43808) );
  AND U42924 ( .A(n22046), .B(n22047), .Z(n43809) );
  IV U42925 ( .A(p_input[894]), .Z(n22047) );
  IV U42926 ( .A(p_input[895]), .Z(n22046) );
  XOR U42927 ( .A(n43812), .B(n43811), .Z(n43810) );
  AND U42928 ( .A(n22048), .B(n22049), .Z(n43811) );
  IV U42929 ( .A(p_input[892]), .Z(n22049) );
  IV U42930 ( .A(p_input[893]), .Z(n22048) );
  XOR U42931 ( .A(n43814), .B(n43813), .Z(n43812) );
  AND U42932 ( .A(n22050), .B(n22051), .Z(n43813) );
  IV U42933 ( .A(p_input[890]), .Z(n22051) );
  IV U42934 ( .A(p_input[891]), .Z(n22050) );
  XOR U42935 ( .A(n43816), .B(n43815), .Z(n43814) );
  AND U42936 ( .A(n22052), .B(n22053), .Z(n43815) );
  IV U42937 ( .A(p_input[888]), .Z(n22053) );
  IV U42938 ( .A(p_input[889]), .Z(n22052) );
  XOR U42939 ( .A(n43818), .B(n43817), .Z(n43816) );
  AND U42940 ( .A(n22054), .B(n22055), .Z(n43817) );
  IV U42941 ( .A(p_input[886]), .Z(n22055) );
  IV U42942 ( .A(p_input[887]), .Z(n22054) );
  XOR U42943 ( .A(n43820), .B(n43819), .Z(n43818) );
  AND U42944 ( .A(n22056), .B(n22057), .Z(n43819) );
  IV U42945 ( .A(p_input[884]), .Z(n22057) );
  IV U42946 ( .A(p_input[885]), .Z(n22056) );
  XOR U42947 ( .A(n43822), .B(n43821), .Z(n43820) );
  AND U42948 ( .A(n22058), .B(n22059), .Z(n43821) );
  IV U42949 ( .A(p_input[882]), .Z(n22059) );
  IV U42950 ( .A(p_input[883]), .Z(n22058) );
  XOR U42951 ( .A(n43824), .B(n43823), .Z(n43822) );
  AND U42952 ( .A(n22060), .B(n22061), .Z(n43823) );
  IV U42953 ( .A(p_input[880]), .Z(n22061) );
  IV U42954 ( .A(p_input[881]), .Z(n22060) );
  XOR U42955 ( .A(n43826), .B(n43825), .Z(n43824) );
  AND U42956 ( .A(n22062), .B(n22063), .Z(n43825) );
  IV U42957 ( .A(p_input[878]), .Z(n22063) );
  IV U42958 ( .A(p_input[879]), .Z(n22062) );
  XOR U42959 ( .A(n43828), .B(n43827), .Z(n43826) );
  AND U42960 ( .A(n22064), .B(n22065), .Z(n43827) );
  IV U42961 ( .A(p_input[876]), .Z(n22065) );
  IV U42962 ( .A(p_input[877]), .Z(n22064) );
  XOR U42963 ( .A(n43830), .B(n43829), .Z(n43828) );
  AND U42964 ( .A(n22066), .B(n22067), .Z(n43829) );
  IV U42965 ( .A(p_input[874]), .Z(n22067) );
  IV U42966 ( .A(p_input[875]), .Z(n22066) );
  XOR U42967 ( .A(n43832), .B(n43831), .Z(n43830) );
  AND U42968 ( .A(n22068), .B(n22069), .Z(n43831) );
  IV U42969 ( .A(p_input[872]), .Z(n22069) );
  IV U42970 ( .A(p_input[873]), .Z(n22068) );
  XOR U42971 ( .A(n43834), .B(n43833), .Z(n43832) );
  AND U42972 ( .A(n22070), .B(n22071), .Z(n43833) );
  IV U42973 ( .A(p_input[870]), .Z(n22071) );
  IV U42974 ( .A(p_input[871]), .Z(n22070) );
  XOR U42975 ( .A(n43836), .B(n43835), .Z(n43834) );
  AND U42976 ( .A(n22072), .B(n22073), .Z(n43835) );
  IV U42977 ( .A(p_input[868]), .Z(n22073) );
  IV U42978 ( .A(p_input[869]), .Z(n22072) );
  XOR U42979 ( .A(n43838), .B(n43837), .Z(n43836) );
  AND U42980 ( .A(n22074), .B(n22075), .Z(n43837) );
  IV U42981 ( .A(p_input[866]), .Z(n22075) );
  IV U42982 ( .A(p_input[867]), .Z(n22074) );
  XOR U42983 ( .A(n43840), .B(n43839), .Z(n43838) );
  AND U42984 ( .A(n22076), .B(n22077), .Z(n43839) );
  IV U42985 ( .A(p_input[864]), .Z(n22077) );
  IV U42986 ( .A(p_input[865]), .Z(n22076) );
  XOR U42987 ( .A(n43842), .B(n43841), .Z(n43840) );
  AND U42988 ( .A(n22078), .B(n22079), .Z(n43841) );
  IV U42989 ( .A(p_input[862]), .Z(n22079) );
  IV U42990 ( .A(p_input[863]), .Z(n22078) );
  XOR U42991 ( .A(n43844), .B(n43843), .Z(n43842) );
  AND U42992 ( .A(n22080), .B(n22081), .Z(n43843) );
  IV U42993 ( .A(p_input[860]), .Z(n22081) );
  IV U42994 ( .A(p_input[861]), .Z(n22080) );
  XOR U42995 ( .A(n43846), .B(n43845), .Z(n43844) );
  AND U42996 ( .A(n22082), .B(n22083), .Z(n43845) );
  IV U42997 ( .A(p_input[858]), .Z(n22083) );
  IV U42998 ( .A(p_input[859]), .Z(n22082) );
  XOR U42999 ( .A(n43848), .B(n43847), .Z(n43846) );
  AND U43000 ( .A(n22084), .B(n22085), .Z(n43847) );
  IV U43001 ( .A(p_input[856]), .Z(n22085) );
  IV U43002 ( .A(p_input[857]), .Z(n22084) );
  XOR U43003 ( .A(n43850), .B(n43849), .Z(n43848) );
  AND U43004 ( .A(n22086), .B(n22087), .Z(n43849) );
  IV U43005 ( .A(p_input[854]), .Z(n22087) );
  IV U43006 ( .A(p_input[855]), .Z(n22086) );
  XOR U43007 ( .A(n43852), .B(n43851), .Z(n43850) );
  AND U43008 ( .A(n22088), .B(n22089), .Z(n43851) );
  IV U43009 ( .A(p_input[852]), .Z(n22089) );
  IV U43010 ( .A(p_input[853]), .Z(n22088) );
  XOR U43011 ( .A(n43854), .B(n43853), .Z(n43852) );
  AND U43012 ( .A(n22090), .B(n22091), .Z(n43853) );
  IV U43013 ( .A(p_input[850]), .Z(n22091) );
  IV U43014 ( .A(p_input[851]), .Z(n22090) );
  XOR U43015 ( .A(n43856), .B(n43855), .Z(n43854) );
  AND U43016 ( .A(n22092), .B(n22093), .Z(n43855) );
  IV U43017 ( .A(p_input[848]), .Z(n22093) );
  IV U43018 ( .A(p_input[849]), .Z(n22092) );
  XOR U43019 ( .A(n43858), .B(n43857), .Z(n43856) );
  AND U43020 ( .A(n22094), .B(n22095), .Z(n43857) );
  IV U43021 ( .A(p_input[846]), .Z(n22095) );
  IV U43022 ( .A(p_input[847]), .Z(n22094) );
  XOR U43023 ( .A(n43860), .B(n43859), .Z(n43858) );
  AND U43024 ( .A(n22096), .B(n22097), .Z(n43859) );
  IV U43025 ( .A(p_input[844]), .Z(n22097) );
  IV U43026 ( .A(p_input[845]), .Z(n22096) );
  XOR U43027 ( .A(n43862), .B(n43861), .Z(n43860) );
  AND U43028 ( .A(n22098), .B(n22099), .Z(n43861) );
  IV U43029 ( .A(p_input[842]), .Z(n22099) );
  IV U43030 ( .A(p_input[843]), .Z(n22098) );
  XOR U43031 ( .A(n43864), .B(n43863), .Z(n43862) );
  AND U43032 ( .A(n22100), .B(n22101), .Z(n43863) );
  IV U43033 ( .A(p_input[840]), .Z(n22101) );
  IV U43034 ( .A(p_input[841]), .Z(n22100) );
  XOR U43035 ( .A(n43866), .B(n43865), .Z(n43864) );
  AND U43036 ( .A(n22102), .B(n22103), .Z(n43865) );
  IV U43037 ( .A(p_input[838]), .Z(n22103) );
  IV U43038 ( .A(p_input[839]), .Z(n22102) );
  XOR U43039 ( .A(n43868), .B(n43867), .Z(n43866) );
  AND U43040 ( .A(n22104), .B(n22105), .Z(n43867) );
  IV U43041 ( .A(p_input[836]), .Z(n22105) );
  IV U43042 ( .A(p_input[837]), .Z(n22104) );
  XOR U43043 ( .A(n43870), .B(n43869), .Z(n43868) );
  AND U43044 ( .A(n22106), .B(n22107), .Z(n43869) );
  IV U43045 ( .A(p_input[834]), .Z(n22107) );
  IV U43046 ( .A(p_input[835]), .Z(n22106) );
  XOR U43047 ( .A(n43872), .B(n43871), .Z(n43870) );
  AND U43048 ( .A(n22108), .B(n22109), .Z(n43871) );
  IV U43049 ( .A(p_input[832]), .Z(n22109) );
  IV U43050 ( .A(p_input[833]), .Z(n22108) );
  XOR U43051 ( .A(n43874), .B(n43873), .Z(n43872) );
  AND U43052 ( .A(n22110), .B(n22111), .Z(n43873) );
  IV U43053 ( .A(p_input[830]), .Z(n22111) );
  IV U43054 ( .A(p_input[831]), .Z(n22110) );
  XOR U43055 ( .A(n43876), .B(n43875), .Z(n43874) );
  AND U43056 ( .A(n22112), .B(n22113), .Z(n43875) );
  IV U43057 ( .A(p_input[828]), .Z(n22113) );
  IV U43058 ( .A(p_input[829]), .Z(n22112) );
  XOR U43059 ( .A(n43878), .B(n43877), .Z(n43876) );
  AND U43060 ( .A(n22114), .B(n22115), .Z(n43877) );
  IV U43061 ( .A(p_input[826]), .Z(n22115) );
  IV U43062 ( .A(p_input[827]), .Z(n22114) );
  XOR U43063 ( .A(n43880), .B(n43879), .Z(n43878) );
  AND U43064 ( .A(n22116), .B(n22117), .Z(n43879) );
  IV U43065 ( .A(p_input[824]), .Z(n22117) );
  IV U43066 ( .A(p_input[825]), .Z(n22116) );
  XOR U43067 ( .A(n43882), .B(n43881), .Z(n43880) );
  AND U43068 ( .A(n22118), .B(n22119), .Z(n43881) );
  IV U43069 ( .A(p_input[822]), .Z(n22119) );
  IV U43070 ( .A(p_input[823]), .Z(n22118) );
  XOR U43071 ( .A(n43884), .B(n43883), .Z(n43882) );
  AND U43072 ( .A(n22120), .B(n22121), .Z(n43883) );
  IV U43073 ( .A(p_input[820]), .Z(n22121) );
  IV U43074 ( .A(p_input[821]), .Z(n22120) );
  XOR U43075 ( .A(n43886), .B(n43885), .Z(n43884) );
  AND U43076 ( .A(n22122), .B(n22123), .Z(n43885) );
  IV U43077 ( .A(p_input[818]), .Z(n22123) );
  IV U43078 ( .A(p_input[819]), .Z(n22122) );
  XOR U43079 ( .A(n43888), .B(n43887), .Z(n43886) );
  AND U43080 ( .A(n22124), .B(n22125), .Z(n43887) );
  IV U43081 ( .A(p_input[816]), .Z(n22125) );
  IV U43082 ( .A(p_input[817]), .Z(n22124) );
  XOR U43083 ( .A(n43890), .B(n43889), .Z(n43888) );
  AND U43084 ( .A(n22126), .B(n22127), .Z(n43889) );
  IV U43085 ( .A(p_input[814]), .Z(n22127) );
  IV U43086 ( .A(p_input[815]), .Z(n22126) );
  XOR U43087 ( .A(n43892), .B(n43891), .Z(n43890) );
  AND U43088 ( .A(n22128), .B(n22129), .Z(n43891) );
  IV U43089 ( .A(p_input[812]), .Z(n22129) );
  IV U43090 ( .A(p_input[813]), .Z(n22128) );
  XOR U43091 ( .A(n43894), .B(n43893), .Z(n43892) );
  AND U43092 ( .A(n22130), .B(n22131), .Z(n43893) );
  IV U43093 ( .A(p_input[810]), .Z(n22131) );
  IV U43094 ( .A(p_input[811]), .Z(n22130) );
  XOR U43095 ( .A(n43896), .B(n43895), .Z(n43894) );
  AND U43096 ( .A(n22132), .B(n22133), .Z(n43895) );
  IV U43097 ( .A(p_input[808]), .Z(n22133) );
  IV U43098 ( .A(p_input[809]), .Z(n22132) );
  XOR U43099 ( .A(n43898), .B(n43897), .Z(n43896) );
  AND U43100 ( .A(n22134), .B(n22135), .Z(n43897) );
  IV U43101 ( .A(p_input[806]), .Z(n22135) );
  IV U43102 ( .A(p_input[807]), .Z(n22134) );
  XOR U43103 ( .A(n43900), .B(n43899), .Z(n43898) );
  AND U43104 ( .A(n22136), .B(n22137), .Z(n43899) );
  IV U43105 ( .A(p_input[804]), .Z(n22137) );
  IV U43106 ( .A(p_input[805]), .Z(n22136) );
  XOR U43107 ( .A(n43902), .B(n43901), .Z(n43900) );
  AND U43108 ( .A(n22138), .B(n22139), .Z(n43901) );
  IV U43109 ( .A(p_input[802]), .Z(n22139) );
  IV U43110 ( .A(p_input[803]), .Z(n22138) );
  XOR U43111 ( .A(n43904), .B(n43903), .Z(n43902) );
  AND U43112 ( .A(n22140), .B(n22141), .Z(n43903) );
  IV U43113 ( .A(p_input[800]), .Z(n22141) );
  IV U43114 ( .A(p_input[801]), .Z(n22140) );
  XOR U43115 ( .A(n43906), .B(n43905), .Z(n43904) );
  AND U43116 ( .A(n22142), .B(n22143), .Z(n43905) );
  IV U43117 ( .A(p_input[798]), .Z(n22143) );
  IV U43118 ( .A(p_input[799]), .Z(n22142) );
  XOR U43119 ( .A(n43908), .B(n43907), .Z(n43906) );
  AND U43120 ( .A(n22144), .B(n22145), .Z(n43907) );
  IV U43121 ( .A(p_input[796]), .Z(n22145) );
  IV U43122 ( .A(p_input[797]), .Z(n22144) );
  XOR U43123 ( .A(n43910), .B(n43909), .Z(n43908) );
  AND U43124 ( .A(n22146), .B(n22147), .Z(n43909) );
  IV U43125 ( .A(p_input[794]), .Z(n22147) );
  IV U43126 ( .A(p_input[795]), .Z(n22146) );
  XOR U43127 ( .A(n43912), .B(n43911), .Z(n43910) );
  AND U43128 ( .A(n22148), .B(n22149), .Z(n43911) );
  IV U43129 ( .A(p_input[792]), .Z(n22149) );
  IV U43130 ( .A(p_input[793]), .Z(n22148) );
  XOR U43131 ( .A(n43914), .B(n43913), .Z(n43912) );
  AND U43132 ( .A(n22150), .B(n22151), .Z(n43913) );
  IV U43133 ( .A(p_input[790]), .Z(n22151) );
  IV U43134 ( .A(p_input[791]), .Z(n22150) );
  XOR U43135 ( .A(n43916), .B(n43915), .Z(n43914) );
  AND U43136 ( .A(n22152), .B(n22153), .Z(n43915) );
  IV U43137 ( .A(p_input[788]), .Z(n22153) );
  IV U43138 ( .A(p_input[789]), .Z(n22152) );
  XOR U43139 ( .A(n43918), .B(n43917), .Z(n43916) );
  AND U43140 ( .A(n22154), .B(n22155), .Z(n43917) );
  IV U43141 ( .A(p_input[786]), .Z(n22155) );
  IV U43142 ( .A(p_input[787]), .Z(n22154) );
  XOR U43143 ( .A(n43920), .B(n43919), .Z(n43918) );
  AND U43144 ( .A(n22156), .B(n22157), .Z(n43919) );
  IV U43145 ( .A(p_input[784]), .Z(n22157) );
  IV U43146 ( .A(p_input[785]), .Z(n22156) );
  XOR U43147 ( .A(n43922), .B(n43921), .Z(n43920) );
  AND U43148 ( .A(n22158), .B(n22159), .Z(n43921) );
  IV U43149 ( .A(p_input[782]), .Z(n22159) );
  IV U43150 ( .A(p_input[783]), .Z(n22158) );
  XOR U43151 ( .A(n43924), .B(n43923), .Z(n43922) );
  AND U43152 ( .A(n22160), .B(n22161), .Z(n43923) );
  IV U43153 ( .A(p_input[780]), .Z(n22161) );
  IV U43154 ( .A(p_input[781]), .Z(n22160) );
  XOR U43155 ( .A(n43926), .B(n43925), .Z(n43924) );
  AND U43156 ( .A(n22162), .B(n22163), .Z(n43925) );
  IV U43157 ( .A(p_input[778]), .Z(n22163) );
  IV U43158 ( .A(p_input[779]), .Z(n22162) );
  XOR U43159 ( .A(n43928), .B(n43927), .Z(n43926) );
  AND U43160 ( .A(n22164), .B(n22165), .Z(n43927) );
  IV U43161 ( .A(p_input[776]), .Z(n22165) );
  IV U43162 ( .A(p_input[777]), .Z(n22164) );
  XOR U43163 ( .A(n43930), .B(n43929), .Z(n43928) );
  AND U43164 ( .A(n22166), .B(n22167), .Z(n43929) );
  IV U43165 ( .A(p_input[774]), .Z(n22167) );
  IV U43166 ( .A(p_input[775]), .Z(n22166) );
  XOR U43167 ( .A(n43932), .B(n43931), .Z(n43930) );
  AND U43168 ( .A(n22168), .B(n22169), .Z(n43931) );
  IV U43169 ( .A(p_input[772]), .Z(n22169) );
  IV U43170 ( .A(p_input[773]), .Z(n22168) );
  XOR U43171 ( .A(n43934), .B(n43933), .Z(n43932) );
  AND U43172 ( .A(n22170), .B(n22171), .Z(n43933) );
  IV U43173 ( .A(p_input[770]), .Z(n22171) );
  IV U43174 ( .A(p_input[771]), .Z(n22170) );
  XOR U43175 ( .A(n43936), .B(n43935), .Z(n43934) );
  AND U43176 ( .A(n22172), .B(n22173), .Z(n43935) );
  IV U43177 ( .A(p_input[768]), .Z(n22173) );
  IV U43178 ( .A(p_input[769]), .Z(n22172) );
  XOR U43179 ( .A(n43938), .B(n43937), .Z(n43936) );
  AND U43180 ( .A(n22174), .B(n22175), .Z(n43937) );
  IV U43181 ( .A(p_input[766]), .Z(n22175) );
  IV U43182 ( .A(p_input[767]), .Z(n22174) );
  XOR U43183 ( .A(n43940), .B(n43939), .Z(n43938) );
  AND U43184 ( .A(n22176), .B(n22177), .Z(n43939) );
  IV U43185 ( .A(p_input[764]), .Z(n22177) );
  IV U43186 ( .A(p_input[765]), .Z(n22176) );
  XOR U43187 ( .A(n43942), .B(n43941), .Z(n43940) );
  AND U43188 ( .A(n22178), .B(n22179), .Z(n43941) );
  IV U43189 ( .A(p_input[762]), .Z(n22179) );
  IV U43190 ( .A(p_input[763]), .Z(n22178) );
  XOR U43191 ( .A(n43944), .B(n43943), .Z(n43942) );
  AND U43192 ( .A(n22180), .B(n22181), .Z(n43943) );
  IV U43193 ( .A(p_input[760]), .Z(n22181) );
  IV U43194 ( .A(p_input[761]), .Z(n22180) );
  XOR U43195 ( .A(n43946), .B(n43945), .Z(n43944) );
  AND U43196 ( .A(n22182), .B(n22183), .Z(n43945) );
  IV U43197 ( .A(p_input[758]), .Z(n22183) );
  IV U43198 ( .A(p_input[759]), .Z(n22182) );
  XOR U43199 ( .A(n43948), .B(n43947), .Z(n43946) );
  AND U43200 ( .A(n22184), .B(n22185), .Z(n43947) );
  IV U43201 ( .A(p_input[756]), .Z(n22185) );
  IV U43202 ( .A(p_input[757]), .Z(n22184) );
  XOR U43203 ( .A(n43950), .B(n43949), .Z(n43948) );
  AND U43204 ( .A(n22186), .B(n22187), .Z(n43949) );
  IV U43205 ( .A(p_input[754]), .Z(n22187) );
  IV U43206 ( .A(p_input[755]), .Z(n22186) );
  XOR U43207 ( .A(n43952), .B(n43951), .Z(n43950) );
  AND U43208 ( .A(n22188), .B(n22189), .Z(n43951) );
  IV U43209 ( .A(p_input[752]), .Z(n22189) );
  IV U43210 ( .A(p_input[753]), .Z(n22188) );
  XOR U43211 ( .A(n43954), .B(n43953), .Z(n43952) );
  AND U43212 ( .A(n22190), .B(n22191), .Z(n43953) );
  IV U43213 ( .A(p_input[750]), .Z(n22191) );
  IV U43214 ( .A(p_input[751]), .Z(n22190) );
  XOR U43215 ( .A(n43956), .B(n43955), .Z(n43954) );
  AND U43216 ( .A(n22192), .B(n22193), .Z(n43955) );
  IV U43217 ( .A(p_input[748]), .Z(n22193) );
  IV U43218 ( .A(p_input[749]), .Z(n22192) );
  XOR U43219 ( .A(n43958), .B(n43957), .Z(n43956) );
  AND U43220 ( .A(n22194), .B(n22195), .Z(n43957) );
  IV U43221 ( .A(p_input[746]), .Z(n22195) );
  IV U43222 ( .A(p_input[747]), .Z(n22194) );
  XOR U43223 ( .A(n43960), .B(n43959), .Z(n43958) );
  AND U43224 ( .A(n22196), .B(n22197), .Z(n43959) );
  IV U43225 ( .A(p_input[744]), .Z(n22197) );
  IV U43226 ( .A(p_input[745]), .Z(n22196) );
  XOR U43227 ( .A(n43962), .B(n43961), .Z(n43960) );
  AND U43228 ( .A(n22198), .B(n22199), .Z(n43961) );
  IV U43229 ( .A(p_input[742]), .Z(n22199) );
  IV U43230 ( .A(p_input[743]), .Z(n22198) );
  XOR U43231 ( .A(n43964), .B(n43963), .Z(n43962) );
  AND U43232 ( .A(n22200), .B(n22201), .Z(n43963) );
  IV U43233 ( .A(p_input[740]), .Z(n22201) );
  IV U43234 ( .A(p_input[741]), .Z(n22200) );
  XOR U43235 ( .A(n43966), .B(n43965), .Z(n43964) );
  AND U43236 ( .A(n22202), .B(n22203), .Z(n43965) );
  IV U43237 ( .A(p_input[738]), .Z(n22203) );
  IV U43238 ( .A(p_input[739]), .Z(n22202) );
  XOR U43239 ( .A(n43968), .B(n43967), .Z(n43966) );
  AND U43240 ( .A(n22204), .B(n22205), .Z(n43967) );
  IV U43241 ( .A(p_input[736]), .Z(n22205) );
  IV U43242 ( .A(p_input[737]), .Z(n22204) );
  XOR U43243 ( .A(n43970), .B(n43969), .Z(n43968) );
  AND U43244 ( .A(n22206), .B(n22207), .Z(n43969) );
  IV U43245 ( .A(p_input[734]), .Z(n22207) );
  IV U43246 ( .A(p_input[735]), .Z(n22206) );
  XOR U43247 ( .A(n43972), .B(n43971), .Z(n43970) );
  AND U43248 ( .A(n22208), .B(n22209), .Z(n43971) );
  IV U43249 ( .A(p_input[732]), .Z(n22209) );
  IV U43250 ( .A(p_input[733]), .Z(n22208) );
  XOR U43251 ( .A(n43974), .B(n43973), .Z(n43972) );
  AND U43252 ( .A(n22210), .B(n22211), .Z(n43973) );
  IV U43253 ( .A(p_input[730]), .Z(n22211) );
  IV U43254 ( .A(p_input[731]), .Z(n22210) );
  XOR U43255 ( .A(n43976), .B(n43975), .Z(n43974) );
  AND U43256 ( .A(n22212), .B(n22213), .Z(n43975) );
  IV U43257 ( .A(p_input[728]), .Z(n22213) );
  IV U43258 ( .A(p_input[729]), .Z(n22212) );
  XOR U43259 ( .A(n43978), .B(n43977), .Z(n43976) );
  AND U43260 ( .A(n22214), .B(n22215), .Z(n43977) );
  IV U43261 ( .A(p_input[726]), .Z(n22215) );
  IV U43262 ( .A(p_input[727]), .Z(n22214) );
  XOR U43263 ( .A(n43980), .B(n43979), .Z(n43978) );
  AND U43264 ( .A(n22216), .B(n22217), .Z(n43979) );
  IV U43265 ( .A(p_input[724]), .Z(n22217) );
  IV U43266 ( .A(p_input[725]), .Z(n22216) );
  XOR U43267 ( .A(n43982), .B(n43981), .Z(n43980) );
  AND U43268 ( .A(n22218), .B(n22219), .Z(n43981) );
  IV U43269 ( .A(p_input[722]), .Z(n22219) );
  IV U43270 ( .A(p_input[723]), .Z(n22218) );
  XOR U43271 ( .A(n43984), .B(n43983), .Z(n43982) );
  AND U43272 ( .A(n22220), .B(n22221), .Z(n43983) );
  IV U43273 ( .A(p_input[720]), .Z(n22221) );
  IV U43274 ( .A(p_input[721]), .Z(n22220) );
  XOR U43275 ( .A(n43986), .B(n43985), .Z(n43984) );
  AND U43276 ( .A(n22222), .B(n22223), .Z(n43985) );
  IV U43277 ( .A(p_input[718]), .Z(n22223) );
  IV U43278 ( .A(p_input[719]), .Z(n22222) );
  XOR U43279 ( .A(n43988), .B(n43987), .Z(n43986) );
  AND U43280 ( .A(n22224), .B(n22225), .Z(n43987) );
  IV U43281 ( .A(p_input[716]), .Z(n22225) );
  IV U43282 ( .A(p_input[717]), .Z(n22224) );
  XOR U43283 ( .A(n43990), .B(n43989), .Z(n43988) );
  AND U43284 ( .A(n22226), .B(n22227), .Z(n43989) );
  IV U43285 ( .A(p_input[714]), .Z(n22227) );
  IV U43286 ( .A(p_input[715]), .Z(n22226) );
  XOR U43287 ( .A(n43992), .B(n43991), .Z(n43990) );
  AND U43288 ( .A(n22228), .B(n22229), .Z(n43991) );
  IV U43289 ( .A(p_input[712]), .Z(n22229) );
  IV U43290 ( .A(p_input[713]), .Z(n22228) );
  XOR U43291 ( .A(n43994), .B(n43993), .Z(n43992) );
  AND U43292 ( .A(n22230), .B(n22231), .Z(n43993) );
  IV U43293 ( .A(p_input[710]), .Z(n22231) );
  IV U43294 ( .A(p_input[711]), .Z(n22230) );
  XOR U43295 ( .A(n43996), .B(n43995), .Z(n43994) );
  AND U43296 ( .A(n22232), .B(n22233), .Z(n43995) );
  IV U43297 ( .A(p_input[708]), .Z(n22233) );
  IV U43298 ( .A(p_input[709]), .Z(n22232) );
  XOR U43299 ( .A(n43998), .B(n43997), .Z(n43996) );
  AND U43300 ( .A(n22234), .B(n22235), .Z(n43997) );
  IV U43301 ( .A(p_input[706]), .Z(n22235) );
  IV U43302 ( .A(p_input[707]), .Z(n22234) );
  XOR U43303 ( .A(n44000), .B(n43999), .Z(n43998) );
  AND U43304 ( .A(n22236), .B(n22237), .Z(n43999) );
  IV U43305 ( .A(p_input[704]), .Z(n22237) );
  IV U43306 ( .A(p_input[705]), .Z(n22236) );
  XOR U43307 ( .A(n44002), .B(n44001), .Z(n44000) );
  AND U43308 ( .A(n22238), .B(n22239), .Z(n44001) );
  IV U43309 ( .A(p_input[702]), .Z(n22239) );
  IV U43310 ( .A(p_input[703]), .Z(n22238) );
  XOR U43311 ( .A(n44004), .B(n44003), .Z(n44002) );
  AND U43312 ( .A(n22240), .B(n22241), .Z(n44003) );
  IV U43313 ( .A(p_input[700]), .Z(n22241) );
  IV U43314 ( .A(p_input[701]), .Z(n22240) );
  XOR U43315 ( .A(n44006), .B(n44005), .Z(n44004) );
  AND U43316 ( .A(n22242), .B(n22243), .Z(n44005) );
  IV U43317 ( .A(p_input[698]), .Z(n22243) );
  IV U43318 ( .A(p_input[699]), .Z(n22242) );
  XOR U43319 ( .A(n44008), .B(n44007), .Z(n44006) );
  AND U43320 ( .A(n22244), .B(n22245), .Z(n44007) );
  IV U43321 ( .A(p_input[696]), .Z(n22245) );
  IV U43322 ( .A(p_input[697]), .Z(n22244) );
  XOR U43323 ( .A(n44010), .B(n44009), .Z(n44008) );
  AND U43324 ( .A(n22246), .B(n22247), .Z(n44009) );
  IV U43325 ( .A(p_input[694]), .Z(n22247) );
  IV U43326 ( .A(p_input[695]), .Z(n22246) );
  XOR U43327 ( .A(n44012), .B(n44011), .Z(n44010) );
  AND U43328 ( .A(n22248), .B(n22249), .Z(n44011) );
  IV U43329 ( .A(p_input[692]), .Z(n22249) );
  IV U43330 ( .A(p_input[693]), .Z(n22248) );
  XOR U43331 ( .A(n44014), .B(n44013), .Z(n44012) );
  AND U43332 ( .A(n22250), .B(n22251), .Z(n44013) );
  IV U43333 ( .A(p_input[690]), .Z(n22251) );
  IV U43334 ( .A(p_input[691]), .Z(n22250) );
  XOR U43335 ( .A(n44016), .B(n44015), .Z(n44014) );
  AND U43336 ( .A(n22252), .B(n22253), .Z(n44015) );
  IV U43337 ( .A(p_input[688]), .Z(n22253) );
  IV U43338 ( .A(p_input[689]), .Z(n22252) );
  XOR U43339 ( .A(n44018), .B(n44017), .Z(n44016) );
  AND U43340 ( .A(n22254), .B(n22255), .Z(n44017) );
  IV U43341 ( .A(p_input[686]), .Z(n22255) );
  IV U43342 ( .A(p_input[687]), .Z(n22254) );
  XOR U43343 ( .A(n44020), .B(n44019), .Z(n44018) );
  AND U43344 ( .A(n22256), .B(n22257), .Z(n44019) );
  IV U43345 ( .A(p_input[684]), .Z(n22257) );
  IV U43346 ( .A(p_input[685]), .Z(n22256) );
  XOR U43347 ( .A(n44022), .B(n44021), .Z(n44020) );
  AND U43348 ( .A(n22258), .B(n22259), .Z(n44021) );
  IV U43349 ( .A(p_input[682]), .Z(n22259) );
  IV U43350 ( .A(p_input[683]), .Z(n22258) );
  XOR U43351 ( .A(n44024), .B(n44023), .Z(n44022) );
  AND U43352 ( .A(n22260), .B(n22261), .Z(n44023) );
  IV U43353 ( .A(p_input[680]), .Z(n22261) );
  IV U43354 ( .A(p_input[681]), .Z(n22260) );
  XOR U43355 ( .A(n44026), .B(n44025), .Z(n44024) );
  AND U43356 ( .A(n22262), .B(n22263), .Z(n44025) );
  IV U43357 ( .A(p_input[678]), .Z(n22263) );
  IV U43358 ( .A(p_input[679]), .Z(n22262) );
  XOR U43359 ( .A(n44028), .B(n44027), .Z(n44026) );
  AND U43360 ( .A(n22264), .B(n22265), .Z(n44027) );
  IV U43361 ( .A(p_input[676]), .Z(n22265) );
  IV U43362 ( .A(p_input[677]), .Z(n22264) );
  XOR U43363 ( .A(n44030), .B(n44029), .Z(n44028) );
  AND U43364 ( .A(n22266), .B(n22267), .Z(n44029) );
  IV U43365 ( .A(p_input[674]), .Z(n22267) );
  IV U43366 ( .A(p_input[675]), .Z(n22266) );
  XOR U43367 ( .A(n44032), .B(n44031), .Z(n44030) );
  AND U43368 ( .A(n22268), .B(n22269), .Z(n44031) );
  IV U43369 ( .A(p_input[672]), .Z(n22269) );
  IV U43370 ( .A(p_input[673]), .Z(n22268) );
  XOR U43371 ( .A(n44034), .B(n44033), .Z(n44032) );
  AND U43372 ( .A(n22270), .B(n22271), .Z(n44033) );
  IV U43373 ( .A(p_input[670]), .Z(n22271) );
  IV U43374 ( .A(p_input[671]), .Z(n22270) );
  XOR U43375 ( .A(n44036), .B(n44035), .Z(n44034) );
  AND U43376 ( .A(n22272), .B(n22273), .Z(n44035) );
  IV U43377 ( .A(p_input[668]), .Z(n22273) );
  IV U43378 ( .A(p_input[669]), .Z(n22272) );
  XOR U43379 ( .A(n44038), .B(n44037), .Z(n44036) );
  AND U43380 ( .A(n22274), .B(n22275), .Z(n44037) );
  IV U43381 ( .A(p_input[666]), .Z(n22275) );
  IV U43382 ( .A(p_input[667]), .Z(n22274) );
  XOR U43383 ( .A(n44040), .B(n44039), .Z(n44038) );
  AND U43384 ( .A(n22276), .B(n22277), .Z(n44039) );
  IV U43385 ( .A(p_input[664]), .Z(n22277) );
  IV U43386 ( .A(p_input[665]), .Z(n22276) );
  XOR U43387 ( .A(n44042), .B(n44041), .Z(n44040) );
  AND U43388 ( .A(n22278), .B(n22279), .Z(n44041) );
  IV U43389 ( .A(p_input[662]), .Z(n22279) );
  IV U43390 ( .A(p_input[663]), .Z(n22278) );
  XOR U43391 ( .A(n44044), .B(n44043), .Z(n44042) );
  AND U43392 ( .A(n22280), .B(n22281), .Z(n44043) );
  IV U43393 ( .A(p_input[660]), .Z(n22281) );
  IV U43394 ( .A(p_input[661]), .Z(n22280) );
  XOR U43395 ( .A(n44046), .B(n44045), .Z(n44044) );
  AND U43396 ( .A(n22282), .B(n22283), .Z(n44045) );
  IV U43397 ( .A(p_input[658]), .Z(n22283) );
  IV U43398 ( .A(p_input[659]), .Z(n22282) );
  XOR U43399 ( .A(n44048), .B(n44047), .Z(n44046) );
  AND U43400 ( .A(n22284), .B(n22285), .Z(n44047) );
  IV U43401 ( .A(p_input[656]), .Z(n22285) );
  IV U43402 ( .A(p_input[657]), .Z(n22284) );
  XOR U43403 ( .A(n44050), .B(n44049), .Z(n44048) );
  AND U43404 ( .A(n22286), .B(n22287), .Z(n44049) );
  IV U43405 ( .A(p_input[654]), .Z(n22287) );
  IV U43406 ( .A(p_input[655]), .Z(n22286) );
  XOR U43407 ( .A(n44052), .B(n44051), .Z(n44050) );
  AND U43408 ( .A(n22288), .B(n22289), .Z(n44051) );
  IV U43409 ( .A(p_input[652]), .Z(n22289) );
  IV U43410 ( .A(p_input[653]), .Z(n22288) );
  XOR U43411 ( .A(n44054), .B(n44053), .Z(n44052) );
  AND U43412 ( .A(n22290), .B(n22291), .Z(n44053) );
  IV U43413 ( .A(p_input[650]), .Z(n22291) );
  IV U43414 ( .A(p_input[651]), .Z(n22290) );
  XOR U43415 ( .A(n44056), .B(n44055), .Z(n44054) );
  AND U43416 ( .A(n22292), .B(n22293), .Z(n44055) );
  IV U43417 ( .A(p_input[648]), .Z(n22293) );
  IV U43418 ( .A(p_input[649]), .Z(n22292) );
  XOR U43419 ( .A(n44058), .B(n44057), .Z(n44056) );
  AND U43420 ( .A(n22294), .B(n22295), .Z(n44057) );
  IV U43421 ( .A(p_input[646]), .Z(n22295) );
  IV U43422 ( .A(p_input[647]), .Z(n22294) );
  XOR U43423 ( .A(n44060), .B(n44059), .Z(n44058) );
  AND U43424 ( .A(n22296), .B(n22297), .Z(n44059) );
  IV U43425 ( .A(p_input[644]), .Z(n22297) );
  IV U43426 ( .A(p_input[645]), .Z(n22296) );
  XOR U43427 ( .A(n44062), .B(n44061), .Z(n44060) );
  AND U43428 ( .A(n22298), .B(n22299), .Z(n44061) );
  IV U43429 ( .A(p_input[642]), .Z(n22299) );
  IV U43430 ( .A(p_input[643]), .Z(n22298) );
  XOR U43431 ( .A(n44064), .B(n44063), .Z(n44062) );
  AND U43432 ( .A(n22300), .B(n22301), .Z(n44063) );
  IV U43433 ( .A(p_input[640]), .Z(n22301) );
  IV U43434 ( .A(p_input[641]), .Z(n22300) );
  XOR U43435 ( .A(n44066), .B(n44065), .Z(n44064) );
  AND U43436 ( .A(n22302), .B(n22303), .Z(n44065) );
  IV U43437 ( .A(p_input[638]), .Z(n22303) );
  IV U43438 ( .A(p_input[639]), .Z(n22302) );
  XOR U43439 ( .A(n44068), .B(n44067), .Z(n44066) );
  AND U43440 ( .A(n22304), .B(n22305), .Z(n44067) );
  IV U43441 ( .A(p_input[636]), .Z(n22305) );
  IV U43442 ( .A(p_input[637]), .Z(n22304) );
  XOR U43443 ( .A(n44070), .B(n44069), .Z(n44068) );
  AND U43444 ( .A(n22306), .B(n22307), .Z(n44069) );
  IV U43445 ( .A(p_input[634]), .Z(n22307) );
  IV U43446 ( .A(p_input[635]), .Z(n22306) );
  XOR U43447 ( .A(n44072), .B(n44071), .Z(n44070) );
  AND U43448 ( .A(n22308), .B(n22309), .Z(n44071) );
  IV U43449 ( .A(p_input[632]), .Z(n22309) );
  IV U43450 ( .A(p_input[633]), .Z(n22308) );
  XOR U43451 ( .A(n44074), .B(n44073), .Z(n44072) );
  AND U43452 ( .A(n22310), .B(n22311), .Z(n44073) );
  IV U43453 ( .A(p_input[630]), .Z(n22311) );
  IV U43454 ( .A(p_input[631]), .Z(n22310) );
  XOR U43455 ( .A(n44076), .B(n44075), .Z(n44074) );
  AND U43456 ( .A(n22312), .B(n22313), .Z(n44075) );
  IV U43457 ( .A(p_input[628]), .Z(n22313) );
  IV U43458 ( .A(p_input[629]), .Z(n22312) );
  XOR U43459 ( .A(n44078), .B(n44077), .Z(n44076) );
  AND U43460 ( .A(n22314), .B(n22315), .Z(n44077) );
  IV U43461 ( .A(p_input[626]), .Z(n22315) );
  IV U43462 ( .A(p_input[627]), .Z(n22314) );
  XOR U43463 ( .A(n44080), .B(n44079), .Z(n44078) );
  AND U43464 ( .A(n22316), .B(n22317), .Z(n44079) );
  IV U43465 ( .A(p_input[624]), .Z(n22317) );
  IV U43466 ( .A(p_input[625]), .Z(n22316) );
  XOR U43467 ( .A(n44082), .B(n44081), .Z(n44080) );
  AND U43468 ( .A(n22318), .B(n22319), .Z(n44081) );
  IV U43469 ( .A(p_input[622]), .Z(n22319) );
  IV U43470 ( .A(p_input[623]), .Z(n22318) );
  XOR U43471 ( .A(n44084), .B(n44083), .Z(n44082) );
  AND U43472 ( .A(n22320), .B(n22321), .Z(n44083) );
  IV U43473 ( .A(p_input[620]), .Z(n22321) );
  IV U43474 ( .A(p_input[621]), .Z(n22320) );
  XOR U43475 ( .A(n44086), .B(n44085), .Z(n44084) );
  AND U43476 ( .A(n22322), .B(n22323), .Z(n44085) );
  IV U43477 ( .A(p_input[618]), .Z(n22323) );
  IV U43478 ( .A(p_input[619]), .Z(n22322) );
  XOR U43479 ( .A(n44088), .B(n44087), .Z(n44086) );
  AND U43480 ( .A(n22324), .B(n22325), .Z(n44087) );
  IV U43481 ( .A(p_input[616]), .Z(n22325) );
  IV U43482 ( .A(p_input[617]), .Z(n22324) );
  XOR U43483 ( .A(n44090), .B(n44089), .Z(n44088) );
  AND U43484 ( .A(n22326), .B(n22327), .Z(n44089) );
  IV U43485 ( .A(p_input[614]), .Z(n22327) );
  IV U43486 ( .A(p_input[615]), .Z(n22326) );
  XOR U43487 ( .A(n44092), .B(n44091), .Z(n44090) );
  AND U43488 ( .A(n22328), .B(n22329), .Z(n44091) );
  IV U43489 ( .A(p_input[612]), .Z(n22329) );
  IV U43490 ( .A(p_input[613]), .Z(n22328) );
  XOR U43491 ( .A(n44094), .B(n44093), .Z(n44092) );
  AND U43492 ( .A(n22330), .B(n22331), .Z(n44093) );
  IV U43493 ( .A(p_input[610]), .Z(n22331) );
  IV U43494 ( .A(p_input[611]), .Z(n22330) );
  XOR U43495 ( .A(n44096), .B(n44095), .Z(n44094) );
  AND U43496 ( .A(n22332), .B(n22333), .Z(n44095) );
  IV U43497 ( .A(p_input[608]), .Z(n22333) );
  IV U43498 ( .A(p_input[609]), .Z(n22332) );
  XOR U43499 ( .A(n44098), .B(n44097), .Z(n44096) );
  AND U43500 ( .A(n22334), .B(n22335), .Z(n44097) );
  IV U43501 ( .A(p_input[606]), .Z(n22335) );
  IV U43502 ( .A(p_input[607]), .Z(n22334) );
  XOR U43503 ( .A(n44100), .B(n44099), .Z(n44098) );
  AND U43504 ( .A(n22336), .B(n22337), .Z(n44099) );
  IV U43505 ( .A(p_input[604]), .Z(n22337) );
  IV U43506 ( .A(p_input[605]), .Z(n22336) );
  XOR U43507 ( .A(n44102), .B(n44101), .Z(n44100) );
  AND U43508 ( .A(n22338), .B(n22339), .Z(n44101) );
  IV U43509 ( .A(p_input[602]), .Z(n22339) );
  IV U43510 ( .A(p_input[603]), .Z(n22338) );
  XOR U43511 ( .A(n44104), .B(n44103), .Z(n44102) );
  AND U43512 ( .A(n22340), .B(n22341), .Z(n44103) );
  IV U43513 ( .A(p_input[600]), .Z(n22341) );
  IV U43514 ( .A(p_input[601]), .Z(n22340) );
  XOR U43515 ( .A(n44106), .B(n44105), .Z(n44104) );
  AND U43516 ( .A(n22342), .B(n22343), .Z(n44105) );
  IV U43517 ( .A(p_input[598]), .Z(n22343) );
  IV U43518 ( .A(p_input[599]), .Z(n22342) );
  XOR U43519 ( .A(n44108), .B(n44107), .Z(n44106) );
  AND U43520 ( .A(n22344), .B(n22345), .Z(n44107) );
  IV U43521 ( .A(p_input[596]), .Z(n22345) );
  IV U43522 ( .A(p_input[597]), .Z(n22344) );
  XOR U43523 ( .A(n44110), .B(n44109), .Z(n44108) );
  AND U43524 ( .A(n22346), .B(n22347), .Z(n44109) );
  IV U43525 ( .A(p_input[594]), .Z(n22347) );
  IV U43526 ( .A(p_input[595]), .Z(n22346) );
  XOR U43527 ( .A(n44112), .B(n44111), .Z(n44110) );
  AND U43528 ( .A(n22348), .B(n22349), .Z(n44111) );
  IV U43529 ( .A(p_input[592]), .Z(n22349) );
  IV U43530 ( .A(p_input[593]), .Z(n22348) );
  XOR U43531 ( .A(n44114), .B(n44113), .Z(n44112) );
  AND U43532 ( .A(n22350), .B(n22351), .Z(n44113) );
  IV U43533 ( .A(p_input[590]), .Z(n22351) );
  IV U43534 ( .A(p_input[591]), .Z(n22350) );
  XOR U43535 ( .A(n44116), .B(n44115), .Z(n44114) );
  AND U43536 ( .A(n22352), .B(n22353), .Z(n44115) );
  IV U43537 ( .A(p_input[588]), .Z(n22353) );
  IV U43538 ( .A(p_input[589]), .Z(n22352) );
  XOR U43539 ( .A(n44118), .B(n44117), .Z(n44116) );
  AND U43540 ( .A(n22354), .B(n22355), .Z(n44117) );
  IV U43541 ( .A(p_input[586]), .Z(n22355) );
  IV U43542 ( .A(p_input[587]), .Z(n22354) );
  XOR U43543 ( .A(n44120), .B(n44119), .Z(n44118) );
  AND U43544 ( .A(n22356), .B(n22357), .Z(n44119) );
  IV U43545 ( .A(p_input[584]), .Z(n22357) );
  IV U43546 ( .A(p_input[585]), .Z(n22356) );
  XOR U43547 ( .A(n44122), .B(n44121), .Z(n44120) );
  AND U43548 ( .A(n22358), .B(n22359), .Z(n44121) );
  IV U43549 ( .A(p_input[582]), .Z(n22359) );
  IV U43550 ( .A(p_input[583]), .Z(n22358) );
  XOR U43551 ( .A(n44124), .B(n44123), .Z(n44122) );
  AND U43552 ( .A(n22360), .B(n22361), .Z(n44123) );
  IV U43553 ( .A(p_input[580]), .Z(n22361) );
  IV U43554 ( .A(p_input[581]), .Z(n22360) );
  XOR U43555 ( .A(n44126), .B(n44125), .Z(n44124) );
  AND U43556 ( .A(n22362), .B(n22363), .Z(n44125) );
  IV U43557 ( .A(p_input[578]), .Z(n22363) );
  IV U43558 ( .A(p_input[579]), .Z(n22362) );
  XOR U43559 ( .A(n44128), .B(n44127), .Z(n44126) );
  AND U43560 ( .A(n22364), .B(n22365), .Z(n44127) );
  IV U43561 ( .A(p_input[576]), .Z(n22365) );
  IV U43562 ( .A(p_input[577]), .Z(n22364) );
  XOR U43563 ( .A(n44130), .B(n44129), .Z(n44128) );
  AND U43564 ( .A(n22366), .B(n22367), .Z(n44129) );
  IV U43565 ( .A(p_input[574]), .Z(n22367) );
  IV U43566 ( .A(p_input[575]), .Z(n22366) );
  XOR U43567 ( .A(n44132), .B(n44131), .Z(n44130) );
  AND U43568 ( .A(n22368), .B(n22369), .Z(n44131) );
  IV U43569 ( .A(p_input[572]), .Z(n22369) );
  IV U43570 ( .A(p_input[573]), .Z(n22368) );
  XOR U43571 ( .A(n44134), .B(n44133), .Z(n44132) );
  AND U43572 ( .A(n22370), .B(n22371), .Z(n44133) );
  IV U43573 ( .A(p_input[570]), .Z(n22371) );
  IV U43574 ( .A(p_input[571]), .Z(n22370) );
  XOR U43575 ( .A(n44136), .B(n44135), .Z(n44134) );
  AND U43576 ( .A(n22372), .B(n22373), .Z(n44135) );
  IV U43577 ( .A(p_input[568]), .Z(n22373) );
  IV U43578 ( .A(p_input[569]), .Z(n22372) );
  XOR U43579 ( .A(n44138), .B(n44137), .Z(n44136) );
  AND U43580 ( .A(n22374), .B(n22375), .Z(n44137) );
  IV U43581 ( .A(p_input[566]), .Z(n22375) );
  IV U43582 ( .A(p_input[567]), .Z(n22374) );
  XOR U43583 ( .A(n44140), .B(n44139), .Z(n44138) );
  AND U43584 ( .A(n22376), .B(n22377), .Z(n44139) );
  IV U43585 ( .A(p_input[564]), .Z(n22377) );
  IV U43586 ( .A(p_input[565]), .Z(n22376) );
  XOR U43587 ( .A(n44142), .B(n44141), .Z(n44140) );
  AND U43588 ( .A(n22378), .B(n22379), .Z(n44141) );
  IV U43589 ( .A(p_input[562]), .Z(n22379) );
  IV U43590 ( .A(p_input[563]), .Z(n22378) );
  XOR U43591 ( .A(n44144), .B(n44143), .Z(n44142) );
  AND U43592 ( .A(n22380), .B(n22381), .Z(n44143) );
  IV U43593 ( .A(p_input[560]), .Z(n22381) );
  IV U43594 ( .A(p_input[561]), .Z(n22380) );
  XOR U43595 ( .A(n44146), .B(n44145), .Z(n44144) );
  AND U43596 ( .A(n22382), .B(n22383), .Z(n44145) );
  IV U43597 ( .A(p_input[558]), .Z(n22383) );
  IV U43598 ( .A(p_input[559]), .Z(n22382) );
  XOR U43599 ( .A(n44148), .B(n44147), .Z(n44146) );
  AND U43600 ( .A(n22384), .B(n22385), .Z(n44147) );
  IV U43601 ( .A(p_input[556]), .Z(n22385) );
  IV U43602 ( .A(p_input[557]), .Z(n22384) );
  XOR U43603 ( .A(n44150), .B(n44149), .Z(n44148) );
  AND U43604 ( .A(n22386), .B(n22387), .Z(n44149) );
  IV U43605 ( .A(p_input[554]), .Z(n22387) );
  IV U43606 ( .A(p_input[555]), .Z(n22386) );
  XOR U43607 ( .A(n44152), .B(n44151), .Z(n44150) );
  AND U43608 ( .A(n22388), .B(n22389), .Z(n44151) );
  IV U43609 ( .A(p_input[552]), .Z(n22389) );
  IV U43610 ( .A(p_input[553]), .Z(n22388) );
  XOR U43611 ( .A(n44154), .B(n44153), .Z(n44152) );
  AND U43612 ( .A(n22390), .B(n22391), .Z(n44153) );
  IV U43613 ( .A(p_input[550]), .Z(n22391) );
  IV U43614 ( .A(p_input[551]), .Z(n22390) );
  XOR U43615 ( .A(n44156), .B(n44155), .Z(n44154) );
  AND U43616 ( .A(n22392), .B(n22393), .Z(n44155) );
  IV U43617 ( .A(p_input[548]), .Z(n22393) );
  IV U43618 ( .A(p_input[549]), .Z(n22392) );
  XOR U43619 ( .A(n44158), .B(n44157), .Z(n44156) );
  AND U43620 ( .A(n22394), .B(n22395), .Z(n44157) );
  IV U43621 ( .A(p_input[546]), .Z(n22395) );
  IV U43622 ( .A(p_input[547]), .Z(n22394) );
  XOR U43623 ( .A(n44160), .B(n44159), .Z(n44158) );
  AND U43624 ( .A(n22396), .B(n22397), .Z(n44159) );
  IV U43625 ( .A(p_input[544]), .Z(n22397) );
  IV U43626 ( .A(p_input[545]), .Z(n22396) );
  XOR U43627 ( .A(n44162), .B(n44161), .Z(n44160) );
  AND U43628 ( .A(n22398), .B(n22399), .Z(n44161) );
  IV U43629 ( .A(p_input[542]), .Z(n22399) );
  IV U43630 ( .A(p_input[543]), .Z(n22398) );
  XOR U43631 ( .A(n44164), .B(n44163), .Z(n44162) );
  AND U43632 ( .A(n22400), .B(n22401), .Z(n44163) );
  IV U43633 ( .A(p_input[540]), .Z(n22401) );
  IV U43634 ( .A(p_input[541]), .Z(n22400) );
  XOR U43635 ( .A(n44166), .B(n44165), .Z(n44164) );
  AND U43636 ( .A(n22402), .B(n22403), .Z(n44165) );
  IV U43637 ( .A(p_input[538]), .Z(n22403) );
  IV U43638 ( .A(p_input[539]), .Z(n22402) );
  XOR U43639 ( .A(n44168), .B(n44167), .Z(n44166) );
  AND U43640 ( .A(n22404), .B(n22405), .Z(n44167) );
  IV U43641 ( .A(p_input[536]), .Z(n22405) );
  IV U43642 ( .A(p_input[537]), .Z(n22404) );
  XOR U43643 ( .A(n44170), .B(n44169), .Z(n44168) );
  AND U43644 ( .A(n22406), .B(n22407), .Z(n44169) );
  IV U43645 ( .A(p_input[534]), .Z(n22407) );
  IV U43646 ( .A(p_input[535]), .Z(n22406) );
  XOR U43647 ( .A(n44172), .B(n44171), .Z(n44170) );
  AND U43648 ( .A(n22408), .B(n22409), .Z(n44171) );
  IV U43649 ( .A(p_input[532]), .Z(n22409) );
  IV U43650 ( .A(p_input[533]), .Z(n22408) );
  XOR U43651 ( .A(n44174), .B(n44173), .Z(n44172) );
  AND U43652 ( .A(n22410), .B(n22411), .Z(n44173) );
  IV U43653 ( .A(p_input[530]), .Z(n22411) );
  IV U43654 ( .A(p_input[531]), .Z(n22410) );
  XOR U43655 ( .A(n44176), .B(n44175), .Z(n44174) );
  AND U43656 ( .A(n22412), .B(n22413), .Z(n44175) );
  IV U43657 ( .A(p_input[528]), .Z(n22413) );
  IV U43658 ( .A(p_input[529]), .Z(n22412) );
  XOR U43659 ( .A(n44178), .B(n44177), .Z(n44176) );
  AND U43660 ( .A(n22414), .B(n22415), .Z(n44177) );
  IV U43661 ( .A(p_input[526]), .Z(n22415) );
  IV U43662 ( .A(p_input[527]), .Z(n22414) );
  XOR U43663 ( .A(n44180), .B(n44179), .Z(n44178) );
  AND U43664 ( .A(n22416), .B(n22417), .Z(n44179) );
  IV U43665 ( .A(p_input[524]), .Z(n22417) );
  IV U43666 ( .A(p_input[525]), .Z(n22416) );
  XOR U43667 ( .A(n44182), .B(n44181), .Z(n44180) );
  AND U43668 ( .A(n22418), .B(n22419), .Z(n44181) );
  IV U43669 ( .A(p_input[522]), .Z(n22419) );
  IV U43670 ( .A(p_input[523]), .Z(n22418) );
  XOR U43671 ( .A(n44184), .B(n44183), .Z(n44182) );
  AND U43672 ( .A(n22420), .B(n22421), .Z(n44183) );
  IV U43673 ( .A(p_input[520]), .Z(n22421) );
  IV U43674 ( .A(p_input[521]), .Z(n22420) );
  XOR U43675 ( .A(n44186), .B(n44185), .Z(n44184) );
  AND U43676 ( .A(n22422), .B(n22423), .Z(n44185) );
  IV U43677 ( .A(p_input[518]), .Z(n22423) );
  IV U43678 ( .A(p_input[519]), .Z(n22422) );
  XOR U43679 ( .A(n44188), .B(n44187), .Z(n44186) );
  AND U43680 ( .A(n22424), .B(n22425), .Z(n44187) );
  IV U43681 ( .A(p_input[516]), .Z(n22425) );
  IV U43682 ( .A(p_input[517]), .Z(n22424) );
  XOR U43683 ( .A(n44190), .B(n44189), .Z(n44188) );
  AND U43684 ( .A(n22426), .B(n22427), .Z(n44189) );
  IV U43685 ( .A(p_input[514]), .Z(n22427) );
  IV U43686 ( .A(p_input[515]), .Z(n22426) );
  XOR U43687 ( .A(n44192), .B(n44191), .Z(n44190) );
  AND U43688 ( .A(n22428), .B(n22429), .Z(n44191) );
  IV U43689 ( .A(p_input[512]), .Z(n22429) );
  IV U43690 ( .A(p_input[513]), .Z(n22428) );
  XOR U43691 ( .A(n44194), .B(n44193), .Z(n44192) );
  AND U43692 ( .A(n22430), .B(n22431), .Z(n44193) );
  IV U43693 ( .A(p_input[510]), .Z(n22431) );
  IV U43694 ( .A(p_input[511]), .Z(n22430) );
  XOR U43695 ( .A(n44196), .B(n44195), .Z(n44194) );
  AND U43696 ( .A(n22432), .B(n22433), .Z(n44195) );
  IV U43697 ( .A(p_input[508]), .Z(n22433) );
  IV U43698 ( .A(p_input[509]), .Z(n22432) );
  XOR U43699 ( .A(n44198), .B(n44197), .Z(n44196) );
  AND U43700 ( .A(n22434), .B(n22435), .Z(n44197) );
  IV U43701 ( .A(p_input[506]), .Z(n22435) );
  IV U43702 ( .A(p_input[507]), .Z(n22434) );
  XOR U43703 ( .A(n44200), .B(n44199), .Z(n44198) );
  AND U43704 ( .A(n22436), .B(n22437), .Z(n44199) );
  IV U43705 ( .A(p_input[504]), .Z(n22437) );
  IV U43706 ( .A(p_input[505]), .Z(n22436) );
  XOR U43707 ( .A(n44202), .B(n44201), .Z(n44200) );
  AND U43708 ( .A(n22438), .B(n22439), .Z(n44201) );
  IV U43709 ( .A(p_input[502]), .Z(n22439) );
  IV U43710 ( .A(p_input[503]), .Z(n22438) );
  XOR U43711 ( .A(n44204), .B(n44203), .Z(n44202) );
  AND U43712 ( .A(n22440), .B(n22441), .Z(n44203) );
  IV U43713 ( .A(p_input[500]), .Z(n22441) );
  IV U43714 ( .A(p_input[501]), .Z(n22440) );
  XOR U43715 ( .A(n44206), .B(n44205), .Z(n44204) );
  AND U43716 ( .A(n22442), .B(n22443), .Z(n44205) );
  IV U43717 ( .A(p_input[498]), .Z(n22443) );
  IV U43718 ( .A(p_input[499]), .Z(n22442) );
  XOR U43719 ( .A(n44208), .B(n44207), .Z(n44206) );
  AND U43720 ( .A(n22444), .B(n22445), .Z(n44207) );
  IV U43721 ( .A(p_input[496]), .Z(n22445) );
  IV U43722 ( .A(p_input[497]), .Z(n22444) );
  XOR U43723 ( .A(n44210), .B(n44209), .Z(n44208) );
  AND U43724 ( .A(n22446), .B(n22447), .Z(n44209) );
  IV U43725 ( .A(p_input[494]), .Z(n22447) );
  IV U43726 ( .A(p_input[495]), .Z(n22446) );
  XOR U43727 ( .A(n44212), .B(n44211), .Z(n44210) );
  AND U43728 ( .A(n22448), .B(n22449), .Z(n44211) );
  IV U43729 ( .A(p_input[492]), .Z(n22449) );
  IV U43730 ( .A(p_input[493]), .Z(n22448) );
  XOR U43731 ( .A(n44214), .B(n44213), .Z(n44212) );
  AND U43732 ( .A(n22450), .B(n22451), .Z(n44213) );
  IV U43733 ( .A(p_input[490]), .Z(n22451) );
  IV U43734 ( .A(p_input[491]), .Z(n22450) );
  XOR U43735 ( .A(n44216), .B(n44215), .Z(n44214) );
  AND U43736 ( .A(n22452), .B(n22453), .Z(n44215) );
  IV U43737 ( .A(p_input[488]), .Z(n22453) );
  IV U43738 ( .A(p_input[489]), .Z(n22452) );
  XOR U43739 ( .A(n44218), .B(n44217), .Z(n44216) );
  AND U43740 ( .A(n22454), .B(n22455), .Z(n44217) );
  IV U43741 ( .A(p_input[486]), .Z(n22455) );
  IV U43742 ( .A(p_input[487]), .Z(n22454) );
  XOR U43743 ( .A(n44220), .B(n44219), .Z(n44218) );
  AND U43744 ( .A(n22456), .B(n22457), .Z(n44219) );
  IV U43745 ( .A(p_input[484]), .Z(n22457) );
  IV U43746 ( .A(p_input[485]), .Z(n22456) );
  XOR U43747 ( .A(n44222), .B(n44221), .Z(n44220) );
  AND U43748 ( .A(n22458), .B(n22459), .Z(n44221) );
  IV U43749 ( .A(p_input[482]), .Z(n22459) );
  IV U43750 ( .A(p_input[483]), .Z(n22458) );
  XOR U43751 ( .A(n44224), .B(n44223), .Z(n44222) );
  AND U43752 ( .A(n22460), .B(n22461), .Z(n44223) );
  IV U43753 ( .A(p_input[480]), .Z(n22461) );
  IV U43754 ( .A(p_input[481]), .Z(n22460) );
  XOR U43755 ( .A(n44226), .B(n44225), .Z(n44224) );
  AND U43756 ( .A(n22462), .B(n22463), .Z(n44225) );
  IV U43757 ( .A(p_input[478]), .Z(n22463) );
  IV U43758 ( .A(p_input[479]), .Z(n22462) );
  XOR U43759 ( .A(n44228), .B(n44227), .Z(n44226) );
  AND U43760 ( .A(n22464), .B(n22465), .Z(n44227) );
  IV U43761 ( .A(p_input[476]), .Z(n22465) );
  IV U43762 ( .A(p_input[477]), .Z(n22464) );
  XOR U43763 ( .A(n44230), .B(n44229), .Z(n44228) );
  AND U43764 ( .A(n22466), .B(n22467), .Z(n44229) );
  IV U43765 ( .A(p_input[474]), .Z(n22467) );
  IV U43766 ( .A(p_input[475]), .Z(n22466) );
  XOR U43767 ( .A(n44232), .B(n44231), .Z(n44230) );
  AND U43768 ( .A(n22468), .B(n22469), .Z(n44231) );
  IV U43769 ( .A(p_input[472]), .Z(n22469) );
  IV U43770 ( .A(p_input[473]), .Z(n22468) );
  XOR U43771 ( .A(n44234), .B(n44233), .Z(n44232) );
  AND U43772 ( .A(n22470), .B(n22471), .Z(n44233) );
  IV U43773 ( .A(p_input[470]), .Z(n22471) );
  IV U43774 ( .A(p_input[471]), .Z(n22470) );
  XOR U43775 ( .A(n44236), .B(n44235), .Z(n44234) );
  AND U43776 ( .A(n22472), .B(n22473), .Z(n44235) );
  IV U43777 ( .A(p_input[468]), .Z(n22473) );
  IV U43778 ( .A(p_input[469]), .Z(n22472) );
  XOR U43779 ( .A(n44238), .B(n44237), .Z(n44236) );
  AND U43780 ( .A(n22474), .B(n22475), .Z(n44237) );
  IV U43781 ( .A(p_input[466]), .Z(n22475) );
  IV U43782 ( .A(p_input[467]), .Z(n22474) );
  XOR U43783 ( .A(n44240), .B(n44239), .Z(n44238) );
  AND U43784 ( .A(n22476), .B(n22477), .Z(n44239) );
  IV U43785 ( .A(p_input[464]), .Z(n22477) );
  IV U43786 ( .A(p_input[465]), .Z(n22476) );
  XOR U43787 ( .A(n44242), .B(n44241), .Z(n44240) );
  AND U43788 ( .A(n22478), .B(n22479), .Z(n44241) );
  IV U43789 ( .A(p_input[462]), .Z(n22479) );
  IV U43790 ( .A(p_input[463]), .Z(n22478) );
  XOR U43791 ( .A(n44244), .B(n44243), .Z(n44242) );
  AND U43792 ( .A(n22480), .B(n22481), .Z(n44243) );
  IV U43793 ( .A(p_input[460]), .Z(n22481) );
  IV U43794 ( .A(p_input[461]), .Z(n22480) );
  XOR U43795 ( .A(n44246), .B(n44245), .Z(n44244) );
  AND U43796 ( .A(n22482), .B(n22483), .Z(n44245) );
  IV U43797 ( .A(p_input[458]), .Z(n22483) );
  IV U43798 ( .A(p_input[459]), .Z(n22482) );
  XOR U43799 ( .A(n44248), .B(n44247), .Z(n44246) );
  AND U43800 ( .A(n22484), .B(n22485), .Z(n44247) );
  IV U43801 ( .A(p_input[456]), .Z(n22485) );
  IV U43802 ( .A(p_input[457]), .Z(n22484) );
  XOR U43803 ( .A(n44250), .B(n44249), .Z(n44248) );
  AND U43804 ( .A(n22486), .B(n22487), .Z(n44249) );
  IV U43805 ( .A(p_input[454]), .Z(n22487) );
  IV U43806 ( .A(p_input[455]), .Z(n22486) );
  XOR U43807 ( .A(n44252), .B(n44251), .Z(n44250) );
  AND U43808 ( .A(n22488), .B(n22489), .Z(n44251) );
  IV U43809 ( .A(p_input[452]), .Z(n22489) );
  IV U43810 ( .A(p_input[453]), .Z(n22488) );
  XOR U43811 ( .A(n44254), .B(n44253), .Z(n44252) );
  AND U43812 ( .A(n22490), .B(n22491), .Z(n44253) );
  IV U43813 ( .A(p_input[450]), .Z(n22491) );
  IV U43814 ( .A(p_input[451]), .Z(n22490) );
  XOR U43815 ( .A(n44256), .B(n44255), .Z(n44254) );
  AND U43816 ( .A(n22492), .B(n22493), .Z(n44255) );
  IV U43817 ( .A(p_input[448]), .Z(n22493) );
  IV U43818 ( .A(p_input[449]), .Z(n22492) );
  XOR U43819 ( .A(n44258), .B(n44257), .Z(n44256) );
  AND U43820 ( .A(n22494), .B(n22495), .Z(n44257) );
  IV U43821 ( .A(p_input[446]), .Z(n22495) );
  IV U43822 ( .A(p_input[447]), .Z(n22494) );
  XOR U43823 ( .A(n44260), .B(n44259), .Z(n44258) );
  AND U43824 ( .A(n22496), .B(n22497), .Z(n44259) );
  IV U43825 ( .A(p_input[444]), .Z(n22497) );
  IV U43826 ( .A(p_input[445]), .Z(n22496) );
  XOR U43827 ( .A(n44262), .B(n44261), .Z(n44260) );
  AND U43828 ( .A(n22498), .B(n22499), .Z(n44261) );
  IV U43829 ( .A(p_input[442]), .Z(n22499) );
  IV U43830 ( .A(p_input[443]), .Z(n22498) );
  XOR U43831 ( .A(n44264), .B(n44263), .Z(n44262) );
  AND U43832 ( .A(n22500), .B(n22501), .Z(n44263) );
  IV U43833 ( .A(p_input[440]), .Z(n22501) );
  IV U43834 ( .A(p_input[441]), .Z(n22500) );
  XOR U43835 ( .A(n44266), .B(n44265), .Z(n44264) );
  AND U43836 ( .A(n22502), .B(n22503), .Z(n44265) );
  IV U43837 ( .A(p_input[438]), .Z(n22503) );
  IV U43838 ( .A(p_input[439]), .Z(n22502) );
  XOR U43839 ( .A(n44268), .B(n44267), .Z(n44266) );
  AND U43840 ( .A(n22504), .B(n22505), .Z(n44267) );
  IV U43841 ( .A(p_input[436]), .Z(n22505) );
  IV U43842 ( .A(p_input[437]), .Z(n22504) );
  XOR U43843 ( .A(n44270), .B(n44269), .Z(n44268) );
  AND U43844 ( .A(n22506), .B(n22507), .Z(n44269) );
  IV U43845 ( .A(p_input[434]), .Z(n22507) );
  IV U43846 ( .A(p_input[435]), .Z(n22506) );
  XOR U43847 ( .A(n44272), .B(n44271), .Z(n44270) );
  AND U43848 ( .A(n22508), .B(n22509), .Z(n44271) );
  IV U43849 ( .A(p_input[432]), .Z(n22509) );
  IV U43850 ( .A(p_input[433]), .Z(n22508) );
  XOR U43851 ( .A(n44274), .B(n44273), .Z(n44272) );
  AND U43852 ( .A(n22510), .B(n22511), .Z(n44273) );
  IV U43853 ( .A(p_input[430]), .Z(n22511) );
  IV U43854 ( .A(p_input[431]), .Z(n22510) );
  XOR U43855 ( .A(n44276), .B(n44275), .Z(n44274) );
  AND U43856 ( .A(n22512), .B(n22513), .Z(n44275) );
  IV U43857 ( .A(p_input[428]), .Z(n22513) );
  IV U43858 ( .A(p_input[429]), .Z(n22512) );
  XOR U43859 ( .A(n44278), .B(n44277), .Z(n44276) );
  AND U43860 ( .A(n22514), .B(n22515), .Z(n44277) );
  IV U43861 ( .A(p_input[426]), .Z(n22515) );
  IV U43862 ( .A(p_input[427]), .Z(n22514) );
  XOR U43863 ( .A(n44280), .B(n44279), .Z(n44278) );
  AND U43864 ( .A(n22516), .B(n22517), .Z(n44279) );
  IV U43865 ( .A(p_input[424]), .Z(n22517) );
  IV U43866 ( .A(p_input[425]), .Z(n22516) );
  XOR U43867 ( .A(n44282), .B(n44281), .Z(n44280) );
  AND U43868 ( .A(n22518), .B(n22519), .Z(n44281) );
  IV U43869 ( .A(p_input[422]), .Z(n22519) );
  IV U43870 ( .A(p_input[423]), .Z(n22518) );
  XOR U43871 ( .A(n44284), .B(n44283), .Z(n44282) );
  AND U43872 ( .A(n22520), .B(n22521), .Z(n44283) );
  IV U43873 ( .A(p_input[420]), .Z(n22521) );
  IV U43874 ( .A(p_input[421]), .Z(n22520) );
  XOR U43875 ( .A(n44286), .B(n44285), .Z(n44284) );
  AND U43876 ( .A(n22522), .B(n22523), .Z(n44285) );
  IV U43877 ( .A(p_input[418]), .Z(n22523) );
  IV U43878 ( .A(p_input[419]), .Z(n22522) );
  XOR U43879 ( .A(n44288), .B(n44287), .Z(n44286) );
  AND U43880 ( .A(n22524), .B(n22525), .Z(n44287) );
  IV U43881 ( .A(p_input[416]), .Z(n22525) );
  IV U43882 ( .A(p_input[417]), .Z(n22524) );
  XOR U43883 ( .A(n44290), .B(n44289), .Z(n44288) );
  AND U43884 ( .A(n22526), .B(n22527), .Z(n44289) );
  IV U43885 ( .A(p_input[414]), .Z(n22527) );
  IV U43886 ( .A(p_input[415]), .Z(n22526) );
  XOR U43887 ( .A(n44292), .B(n44291), .Z(n44290) );
  AND U43888 ( .A(n22528), .B(n22529), .Z(n44291) );
  IV U43889 ( .A(p_input[412]), .Z(n22529) );
  IV U43890 ( .A(p_input[413]), .Z(n22528) );
  XOR U43891 ( .A(n44294), .B(n44293), .Z(n44292) );
  AND U43892 ( .A(n22530), .B(n22531), .Z(n44293) );
  IV U43893 ( .A(p_input[410]), .Z(n22531) );
  IV U43894 ( .A(p_input[411]), .Z(n22530) );
  XOR U43895 ( .A(n44296), .B(n44295), .Z(n44294) );
  AND U43896 ( .A(n22532), .B(n22533), .Z(n44295) );
  IV U43897 ( .A(p_input[408]), .Z(n22533) );
  IV U43898 ( .A(p_input[409]), .Z(n22532) );
  XOR U43899 ( .A(n44298), .B(n44297), .Z(n44296) );
  AND U43900 ( .A(n22534), .B(n22535), .Z(n44297) );
  IV U43901 ( .A(p_input[406]), .Z(n22535) );
  IV U43902 ( .A(p_input[407]), .Z(n22534) );
  XOR U43903 ( .A(n44300), .B(n44299), .Z(n44298) );
  AND U43904 ( .A(n22536), .B(n22537), .Z(n44299) );
  IV U43905 ( .A(p_input[404]), .Z(n22537) );
  IV U43906 ( .A(p_input[405]), .Z(n22536) );
  XOR U43907 ( .A(n44302), .B(n44301), .Z(n44300) );
  AND U43908 ( .A(n22538), .B(n22539), .Z(n44301) );
  IV U43909 ( .A(p_input[402]), .Z(n22539) );
  IV U43910 ( .A(p_input[403]), .Z(n22538) );
  XOR U43911 ( .A(n44304), .B(n44303), .Z(n44302) );
  AND U43912 ( .A(n22540), .B(n22541), .Z(n44303) );
  IV U43913 ( .A(p_input[400]), .Z(n22541) );
  IV U43914 ( .A(p_input[401]), .Z(n22540) );
  XOR U43915 ( .A(n44306), .B(n44305), .Z(n44304) );
  AND U43916 ( .A(n22542), .B(n22543), .Z(n44305) );
  IV U43917 ( .A(p_input[398]), .Z(n22543) );
  IV U43918 ( .A(p_input[399]), .Z(n22542) );
  XOR U43919 ( .A(n44308), .B(n44307), .Z(n44306) );
  AND U43920 ( .A(n22544), .B(n22545), .Z(n44307) );
  IV U43921 ( .A(p_input[396]), .Z(n22545) );
  IV U43922 ( .A(p_input[397]), .Z(n22544) );
  XOR U43923 ( .A(n44310), .B(n44309), .Z(n44308) );
  AND U43924 ( .A(n22546), .B(n22547), .Z(n44309) );
  IV U43925 ( .A(p_input[394]), .Z(n22547) );
  IV U43926 ( .A(p_input[395]), .Z(n22546) );
  XOR U43927 ( .A(n44312), .B(n44311), .Z(n44310) );
  AND U43928 ( .A(n22548), .B(n22549), .Z(n44311) );
  IV U43929 ( .A(p_input[392]), .Z(n22549) );
  IV U43930 ( .A(p_input[393]), .Z(n22548) );
  XOR U43931 ( .A(n44314), .B(n44313), .Z(n44312) );
  AND U43932 ( .A(n22550), .B(n22551), .Z(n44313) );
  IV U43933 ( .A(p_input[390]), .Z(n22551) );
  IV U43934 ( .A(p_input[391]), .Z(n22550) );
  XOR U43935 ( .A(n44316), .B(n44315), .Z(n44314) );
  AND U43936 ( .A(n22552), .B(n22553), .Z(n44315) );
  IV U43937 ( .A(p_input[388]), .Z(n22553) );
  IV U43938 ( .A(p_input[389]), .Z(n22552) );
  XOR U43939 ( .A(n44318), .B(n44317), .Z(n44316) );
  AND U43940 ( .A(n22554), .B(n22555), .Z(n44317) );
  IV U43941 ( .A(p_input[386]), .Z(n22555) );
  IV U43942 ( .A(p_input[387]), .Z(n22554) );
  XOR U43943 ( .A(n44320), .B(n44319), .Z(n44318) );
  AND U43944 ( .A(n22556), .B(n22557), .Z(n44319) );
  IV U43945 ( .A(p_input[384]), .Z(n22557) );
  IV U43946 ( .A(p_input[385]), .Z(n22556) );
  XOR U43947 ( .A(n44322), .B(n44321), .Z(n44320) );
  AND U43948 ( .A(n22558), .B(n22559), .Z(n44321) );
  IV U43949 ( .A(p_input[382]), .Z(n22559) );
  IV U43950 ( .A(p_input[383]), .Z(n22558) );
  XOR U43951 ( .A(n44324), .B(n44323), .Z(n44322) );
  AND U43952 ( .A(n22560), .B(n22561), .Z(n44323) );
  IV U43953 ( .A(p_input[380]), .Z(n22561) );
  IV U43954 ( .A(p_input[381]), .Z(n22560) );
  XOR U43955 ( .A(n44326), .B(n44325), .Z(n44324) );
  AND U43956 ( .A(n22562), .B(n22563), .Z(n44325) );
  IV U43957 ( .A(p_input[378]), .Z(n22563) );
  IV U43958 ( .A(p_input[379]), .Z(n22562) );
  XOR U43959 ( .A(n44328), .B(n44327), .Z(n44326) );
  AND U43960 ( .A(n22564), .B(n22565), .Z(n44327) );
  IV U43961 ( .A(p_input[376]), .Z(n22565) );
  IV U43962 ( .A(p_input[377]), .Z(n22564) );
  XOR U43963 ( .A(n44330), .B(n44329), .Z(n44328) );
  AND U43964 ( .A(n22566), .B(n22567), .Z(n44329) );
  IV U43965 ( .A(p_input[374]), .Z(n22567) );
  IV U43966 ( .A(p_input[375]), .Z(n22566) );
  XOR U43967 ( .A(n44332), .B(n44331), .Z(n44330) );
  AND U43968 ( .A(n22568), .B(n22569), .Z(n44331) );
  IV U43969 ( .A(p_input[372]), .Z(n22569) );
  IV U43970 ( .A(p_input[373]), .Z(n22568) );
  XOR U43971 ( .A(n44334), .B(n44333), .Z(n44332) );
  AND U43972 ( .A(n22570), .B(n22571), .Z(n44333) );
  IV U43973 ( .A(p_input[370]), .Z(n22571) );
  IV U43974 ( .A(p_input[371]), .Z(n22570) );
  XOR U43975 ( .A(n44336), .B(n44335), .Z(n44334) );
  AND U43976 ( .A(n22572), .B(n22573), .Z(n44335) );
  IV U43977 ( .A(p_input[368]), .Z(n22573) );
  IV U43978 ( .A(p_input[369]), .Z(n22572) );
  XOR U43979 ( .A(n44338), .B(n44337), .Z(n44336) );
  AND U43980 ( .A(n22574), .B(n22575), .Z(n44337) );
  IV U43981 ( .A(p_input[366]), .Z(n22575) );
  IV U43982 ( .A(p_input[367]), .Z(n22574) );
  XOR U43983 ( .A(n44340), .B(n44339), .Z(n44338) );
  AND U43984 ( .A(n22576), .B(n22577), .Z(n44339) );
  IV U43985 ( .A(p_input[364]), .Z(n22577) );
  IV U43986 ( .A(p_input[365]), .Z(n22576) );
  XOR U43987 ( .A(n44342), .B(n44341), .Z(n44340) );
  AND U43988 ( .A(n22578), .B(n22579), .Z(n44341) );
  IV U43989 ( .A(p_input[362]), .Z(n22579) );
  IV U43990 ( .A(p_input[363]), .Z(n22578) );
  XOR U43991 ( .A(n44344), .B(n44343), .Z(n44342) );
  AND U43992 ( .A(n22580), .B(n22581), .Z(n44343) );
  IV U43993 ( .A(p_input[360]), .Z(n22581) );
  IV U43994 ( .A(p_input[361]), .Z(n22580) );
  XOR U43995 ( .A(n44346), .B(n44345), .Z(n44344) );
  AND U43996 ( .A(n22582), .B(n22583), .Z(n44345) );
  IV U43997 ( .A(p_input[358]), .Z(n22583) );
  IV U43998 ( .A(p_input[359]), .Z(n22582) );
  XOR U43999 ( .A(n44348), .B(n44347), .Z(n44346) );
  AND U44000 ( .A(n22584), .B(n22585), .Z(n44347) );
  IV U44001 ( .A(p_input[356]), .Z(n22585) );
  IV U44002 ( .A(p_input[357]), .Z(n22584) );
  XOR U44003 ( .A(n44350), .B(n44349), .Z(n44348) );
  AND U44004 ( .A(n22586), .B(n22587), .Z(n44349) );
  IV U44005 ( .A(p_input[354]), .Z(n22587) );
  IV U44006 ( .A(p_input[355]), .Z(n22586) );
  XOR U44007 ( .A(n44352), .B(n44351), .Z(n44350) );
  AND U44008 ( .A(n22588), .B(n22589), .Z(n44351) );
  IV U44009 ( .A(p_input[352]), .Z(n22589) );
  IV U44010 ( .A(p_input[353]), .Z(n22588) );
  XOR U44011 ( .A(n44354), .B(n44353), .Z(n44352) );
  AND U44012 ( .A(n22590), .B(n22591), .Z(n44353) );
  IV U44013 ( .A(p_input[350]), .Z(n22591) );
  IV U44014 ( .A(p_input[351]), .Z(n22590) );
  XOR U44015 ( .A(n44356), .B(n44355), .Z(n44354) );
  AND U44016 ( .A(n22592), .B(n22593), .Z(n44355) );
  IV U44017 ( .A(p_input[348]), .Z(n22593) );
  IV U44018 ( .A(p_input[349]), .Z(n22592) );
  XOR U44019 ( .A(n44358), .B(n44357), .Z(n44356) );
  AND U44020 ( .A(n22594), .B(n22595), .Z(n44357) );
  IV U44021 ( .A(p_input[346]), .Z(n22595) );
  IV U44022 ( .A(p_input[347]), .Z(n22594) );
  XOR U44023 ( .A(n44360), .B(n44359), .Z(n44358) );
  AND U44024 ( .A(n22596), .B(n22597), .Z(n44359) );
  IV U44025 ( .A(p_input[344]), .Z(n22597) );
  IV U44026 ( .A(p_input[345]), .Z(n22596) );
  XOR U44027 ( .A(n44362), .B(n44361), .Z(n44360) );
  AND U44028 ( .A(n22598), .B(n22599), .Z(n44361) );
  IV U44029 ( .A(p_input[342]), .Z(n22599) );
  IV U44030 ( .A(p_input[343]), .Z(n22598) );
  XOR U44031 ( .A(n44364), .B(n44363), .Z(n44362) );
  AND U44032 ( .A(n22600), .B(n22601), .Z(n44363) );
  IV U44033 ( .A(p_input[340]), .Z(n22601) );
  IV U44034 ( .A(p_input[341]), .Z(n22600) );
  XOR U44035 ( .A(n44366), .B(n44365), .Z(n44364) );
  AND U44036 ( .A(n22602), .B(n22603), .Z(n44365) );
  IV U44037 ( .A(p_input[338]), .Z(n22603) );
  IV U44038 ( .A(p_input[339]), .Z(n22602) );
  XOR U44039 ( .A(n44368), .B(n44367), .Z(n44366) );
  AND U44040 ( .A(n22604), .B(n22605), .Z(n44367) );
  IV U44041 ( .A(p_input[336]), .Z(n22605) );
  IV U44042 ( .A(p_input[337]), .Z(n22604) );
  XOR U44043 ( .A(n44370), .B(n44369), .Z(n44368) );
  AND U44044 ( .A(n22606), .B(n22607), .Z(n44369) );
  IV U44045 ( .A(p_input[334]), .Z(n22607) );
  IV U44046 ( .A(p_input[335]), .Z(n22606) );
  XOR U44047 ( .A(n44372), .B(n44371), .Z(n44370) );
  AND U44048 ( .A(n22608), .B(n22609), .Z(n44371) );
  IV U44049 ( .A(p_input[332]), .Z(n22609) );
  IV U44050 ( .A(p_input[333]), .Z(n22608) );
  XOR U44051 ( .A(n44374), .B(n44373), .Z(n44372) );
  AND U44052 ( .A(n22610), .B(n22611), .Z(n44373) );
  IV U44053 ( .A(p_input[330]), .Z(n22611) );
  IV U44054 ( .A(p_input[331]), .Z(n22610) );
  XOR U44055 ( .A(n44376), .B(n44375), .Z(n44374) );
  AND U44056 ( .A(n22612), .B(n22613), .Z(n44375) );
  IV U44057 ( .A(p_input[328]), .Z(n22613) );
  IV U44058 ( .A(p_input[329]), .Z(n22612) );
  XOR U44059 ( .A(n44378), .B(n44377), .Z(n44376) );
  AND U44060 ( .A(n22614), .B(n22615), .Z(n44377) );
  IV U44061 ( .A(p_input[326]), .Z(n22615) );
  IV U44062 ( .A(p_input[327]), .Z(n22614) );
  XOR U44063 ( .A(n44380), .B(n44379), .Z(n44378) );
  AND U44064 ( .A(n22616), .B(n22617), .Z(n44379) );
  IV U44065 ( .A(p_input[324]), .Z(n22617) );
  IV U44066 ( .A(p_input[325]), .Z(n22616) );
  XOR U44067 ( .A(n44382), .B(n44381), .Z(n44380) );
  AND U44068 ( .A(n22618), .B(n22619), .Z(n44381) );
  IV U44069 ( .A(p_input[322]), .Z(n22619) );
  IV U44070 ( .A(p_input[323]), .Z(n22618) );
  XOR U44071 ( .A(n44384), .B(n44383), .Z(n44382) );
  AND U44072 ( .A(n22620), .B(n22621), .Z(n44383) );
  IV U44073 ( .A(p_input[320]), .Z(n22621) );
  IV U44074 ( .A(p_input[321]), .Z(n22620) );
  XOR U44075 ( .A(n44386), .B(n44385), .Z(n44384) );
  AND U44076 ( .A(n22622), .B(n22623), .Z(n44385) );
  IV U44077 ( .A(p_input[318]), .Z(n22623) );
  IV U44078 ( .A(p_input[319]), .Z(n22622) );
  XOR U44079 ( .A(n44388), .B(n44387), .Z(n44386) );
  AND U44080 ( .A(n22624), .B(n22625), .Z(n44387) );
  IV U44081 ( .A(p_input[316]), .Z(n22625) );
  IV U44082 ( .A(p_input[317]), .Z(n22624) );
  XOR U44083 ( .A(n44390), .B(n44389), .Z(n44388) );
  AND U44084 ( .A(n22626), .B(n22627), .Z(n44389) );
  IV U44085 ( .A(p_input[314]), .Z(n22627) );
  IV U44086 ( .A(p_input[315]), .Z(n22626) );
  XOR U44087 ( .A(n44392), .B(n44391), .Z(n44390) );
  AND U44088 ( .A(n22628), .B(n22629), .Z(n44391) );
  IV U44089 ( .A(p_input[312]), .Z(n22629) );
  IV U44090 ( .A(p_input[313]), .Z(n22628) );
  XOR U44091 ( .A(n44394), .B(n44393), .Z(n44392) );
  AND U44092 ( .A(n22630), .B(n22631), .Z(n44393) );
  IV U44093 ( .A(p_input[310]), .Z(n22631) );
  IV U44094 ( .A(p_input[311]), .Z(n22630) );
  XOR U44095 ( .A(n44396), .B(n44395), .Z(n44394) );
  AND U44096 ( .A(n22632), .B(n22633), .Z(n44395) );
  IV U44097 ( .A(p_input[308]), .Z(n22633) );
  IV U44098 ( .A(p_input[309]), .Z(n22632) );
  XOR U44099 ( .A(n44398), .B(n44397), .Z(n44396) );
  AND U44100 ( .A(n22634), .B(n22635), .Z(n44397) );
  IV U44101 ( .A(p_input[306]), .Z(n22635) );
  IV U44102 ( .A(p_input[307]), .Z(n22634) );
  XOR U44103 ( .A(n44400), .B(n44399), .Z(n44398) );
  AND U44104 ( .A(n22636), .B(n22637), .Z(n44399) );
  IV U44105 ( .A(p_input[304]), .Z(n22637) );
  IV U44106 ( .A(p_input[305]), .Z(n22636) );
  XOR U44107 ( .A(n44402), .B(n44401), .Z(n44400) );
  AND U44108 ( .A(n22638), .B(n22639), .Z(n44401) );
  IV U44109 ( .A(p_input[302]), .Z(n22639) );
  IV U44110 ( .A(p_input[303]), .Z(n22638) );
  XOR U44111 ( .A(n44404), .B(n44403), .Z(n44402) );
  AND U44112 ( .A(n22640), .B(n22641), .Z(n44403) );
  IV U44113 ( .A(p_input[300]), .Z(n22641) );
  IV U44114 ( .A(p_input[301]), .Z(n22640) );
  XOR U44115 ( .A(n44406), .B(n44405), .Z(n44404) );
  AND U44116 ( .A(n22642), .B(n22643), .Z(n44405) );
  IV U44117 ( .A(p_input[298]), .Z(n22643) );
  IV U44118 ( .A(p_input[299]), .Z(n22642) );
  XOR U44119 ( .A(n44408), .B(n44407), .Z(n44406) );
  AND U44120 ( .A(n22644), .B(n22645), .Z(n44407) );
  IV U44121 ( .A(p_input[296]), .Z(n22645) );
  IV U44122 ( .A(p_input[297]), .Z(n22644) );
  XOR U44123 ( .A(n44410), .B(n44409), .Z(n44408) );
  AND U44124 ( .A(n22646), .B(n22647), .Z(n44409) );
  IV U44125 ( .A(p_input[294]), .Z(n22647) );
  IV U44126 ( .A(p_input[295]), .Z(n22646) );
  XOR U44127 ( .A(n44412), .B(n44411), .Z(n44410) );
  AND U44128 ( .A(n22648), .B(n22649), .Z(n44411) );
  IV U44129 ( .A(p_input[292]), .Z(n22649) );
  IV U44130 ( .A(p_input[293]), .Z(n22648) );
  XOR U44131 ( .A(n44414), .B(n44413), .Z(n44412) );
  AND U44132 ( .A(n22650), .B(n22651), .Z(n44413) );
  IV U44133 ( .A(p_input[290]), .Z(n22651) );
  IV U44134 ( .A(p_input[291]), .Z(n22650) );
  XOR U44135 ( .A(n44416), .B(n44415), .Z(n44414) );
  AND U44136 ( .A(n22652), .B(n22653), .Z(n44415) );
  IV U44137 ( .A(p_input[288]), .Z(n22653) );
  IV U44138 ( .A(p_input[289]), .Z(n22652) );
  XOR U44139 ( .A(n44418), .B(n44417), .Z(n44416) );
  AND U44140 ( .A(n22654), .B(n22655), .Z(n44417) );
  IV U44141 ( .A(p_input[286]), .Z(n22655) );
  IV U44142 ( .A(p_input[287]), .Z(n22654) );
  XOR U44143 ( .A(n44420), .B(n44419), .Z(n44418) );
  AND U44144 ( .A(n22656), .B(n22657), .Z(n44419) );
  IV U44145 ( .A(p_input[284]), .Z(n22657) );
  IV U44146 ( .A(p_input[285]), .Z(n22656) );
  XOR U44147 ( .A(n44422), .B(n44421), .Z(n44420) );
  AND U44148 ( .A(n22658), .B(n22659), .Z(n44421) );
  IV U44149 ( .A(p_input[282]), .Z(n22659) );
  IV U44150 ( .A(p_input[283]), .Z(n22658) );
  XOR U44151 ( .A(n44424), .B(n44423), .Z(n44422) );
  AND U44152 ( .A(n22660), .B(n22661), .Z(n44423) );
  IV U44153 ( .A(p_input[280]), .Z(n22661) );
  IV U44154 ( .A(p_input[281]), .Z(n22660) );
  XOR U44155 ( .A(n44426), .B(n44425), .Z(n44424) );
  AND U44156 ( .A(n22662), .B(n22663), .Z(n44425) );
  IV U44157 ( .A(p_input[278]), .Z(n22663) );
  IV U44158 ( .A(p_input[279]), .Z(n22662) );
  XOR U44159 ( .A(n44428), .B(n44427), .Z(n44426) );
  AND U44160 ( .A(n22664), .B(n22665), .Z(n44427) );
  IV U44161 ( .A(p_input[276]), .Z(n22665) );
  IV U44162 ( .A(p_input[277]), .Z(n22664) );
  XOR U44163 ( .A(n44430), .B(n44429), .Z(n44428) );
  AND U44164 ( .A(n22666), .B(n22667), .Z(n44429) );
  IV U44165 ( .A(p_input[274]), .Z(n22667) );
  IV U44166 ( .A(p_input[275]), .Z(n22666) );
  XOR U44167 ( .A(n44432), .B(n44431), .Z(n44430) );
  AND U44168 ( .A(n22668), .B(n22669), .Z(n44431) );
  IV U44169 ( .A(p_input[272]), .Z(n22669) );
  IV U44170 ( .A(p_input[273]), .Z(n22668) );
  XOR U44171 ( .A(n44434), .B(n44433), .Z(n44432) );
  AND U44172 ( .A(n22670), .B(n22671), .Z(n44433) );
  IV U44173 ( .A(p_input[270]), .Z(n22671) );
  IV U44174 ( .A(p_input[271]), .Z(n22670) );
  XOR U44175 ( .A(n44436), .B(n44435), .Z(n44434) );
  AND U44176 ( .A(n22672), .B(n22673), .Z(n44435) );
  IV U44177 ( .A(p_input[268]), .Z(n22673) );
  IV U44178 ( .A(p_input[269]), .Z(n22672) );
  XOR U44179 ( .A(n44438), .B(n44437), .Z(n44436) );
  AND U44180 ( .A(n22674), .B(n22675), .Z(n44437) );
  IV U44181 ( .A(p_input[266]), .Z(n22675) );
  IV U44182 ( .A(p_input[267]), .Z(n22674) );
  XOR U44183 ( .A(n44440), .B(n44439), .Z(n44438) );
  AND U44184 ( .A(n22676), .B(n22677), .Z(n44439) );
  IV U44185 ( .A(p_input[264]), .Z(n22677) );
  IV U44186 ( .A(p_input[265]), .Z(n22676) );
  XOR U44187 ( .A(n44442), .B(n44441), .Z(n44440) );
  AND U44188 ( .A(n22678), .B(n22679), .Z(n44441) );
  IV U44189 ( .A(p_input[262]), .Z(n22679) );
  IV U44190 ( .A(p_input[263]), .Z(n22678) );
  XOR U44191 ( .A(n44444), .B(n44443), .Z(n44442) );
  AND U44192 ( .A(n22680), .B(n22681), .Z(n44443) );
  IV U44193 ( .A(p_input[260]), .Z(n22681) );
  IV U44194 ( .A(p_input[261]), .Z(n22680) );
  XOR U44195 ( .A(n44446), .B(n44445), .Z(n44444) );
  AND U44196 ( .A(n22682), .B(n22683), .Z(n44445) );
  IV U44197 ( .A(p_input[258]), .Z(n22683) );
  IV U44198 ( .A(p_input[259]), .Z(n22682) );
  XOR U44199 ( .A(n44448), .B(n44447), .Z(n44446) );
  AND U44200 ( .A(n22684), .B(n22685), .Z(n44447) );
  IV U44201 ( .A(p_input[256]), .Z(n22685) );
  IV U44202 ( .A(p_input[257]), .Z(n22684) );
  XOR U44203 ( .A(n44450), .B(n44449), .Z(n44448) );
  AND U44204 ( .A(n22686), .B(n22687), .Z(n44449) );
  IV U44205 ( .A(p_input[254]), .Z(n22687) );
  IV U44206 ( .A(p_input[255]), .Z(n22686) );
  XOR U44207 ( .A(n44454), .B(n44453), .Z(n44450) );
  AND U44208 ( .A(n22688), .B(n22689), .Z(n44453) );
  IV U44209 ( .A(p_input[252]), .Z(n22689) );
  IV U44210 ( .A(p_input[253]), .Z(n22688) );
  XOR U44211 ( .A(n44456), .B(n44455), .Z(n44454) );
  AND U44212 ( .A(n22690), .B(n22691), .Z(n44455) );
  IV U44213 ( .A(p_input[250]), .Z(n22691) );
  IV U44214 ( .A(p_input[251]), .Z(n22690) );
  XOR U44215 ( .A(n44458), .B(n44457), .Z(n44456) );
  AND U44216 ( .A(n22692), .B(n22693), .Z(n44457) );
  IV U44217 ( .A(p_input[248]), .Z(n22693) );
  IV U44218 ( .A(p_input[249]), .Z(n22692) );
  XOR U44219 ( .A(n44460), .B(n44459), .Z(n44458) );
  AND U44220 ( .A(n22694), .B(n22695), .Z(n44459) );
  IV U44221 ( .A(p_input[246]), .Z(n22695) );
  IV U44222 ( .A(p_input[247]), .Z(n22694) );
  XOR U44223 ( .A(n44462), .B(n44461), .Z(n44460) );
  AND U44224 ( .A(n22696), .B(n22697), .Z(n44461) );
  IV U44225 ( .A(p_input[244]), .Z(n22697) );
  IV U44226 ( .A(p_input[245]), .Z(n22696) );
  XOR U44227 ( .A(n44464), .B(n44463), .Z(n44462) );
  AND U44228 ( .A(n22698), .B(n22699), .Z(n44463) );
  IV U44229 ( .A(p_input[242]), .Z(n22699) );
  IV U44230 ( .A(p_input[243]), .Z(n22698) );
  XOR U44231 ( .A(n44466), .B(n44465), .Z(n44464) );
  AND U44232 ( .A(n22700), .B(n22701), .Z(n44465) );
  IV U44233 ( .A(p_input[240]), .Z(n22701) );
  IV U44234 ( .A(p_input[241]), .Z(n22700) );
  XOR U44235 ( .A(n44468), .B(n44467), .Z(n44466) );
  AND U44236 ( .A(n22702), .B(n22703), .Z(n44467) );
  IV U44237 ( .A(p_input[238]), .Z(n22703) );
  IV U44238 ( .A(p_input[239]), .Z(n22702) );
  XOR U44239 ( .A(n44470), .B(n44469), .Z(n44468) );
  AND U44240 ( .A(n22704), .B(n22705), .Z(n44469) );
  IV U44241 ( .A(p_input[236]), .Z(n22705) );
  IV U44242 ( .A(p_input[237]), .Z(n22704) );
  XOR U44243 ( .A(n44472), .B(n44471), .Z(n44470) );
  AND U44244 ( .A(n22706), .B(n22707), .Z(n44471) );
  IV U44245 ( .A(p_input[234]), .Z(n22707) );
  IV U44246 ( .A(p_input[235]), .Z(n22706) );
  XOR U44247 ( .A(n44474), .B(n44473), .Z(n44472) );
  AND U44248 ( .A(n22708), .B(n22709), .Z(n44473) );
  IV U44249 ( .A(p_input[232]), .Z(n22709) );
  IV U44250 ( .A(p_input[233]), .Z(n22708) );
  XOR U44251 ( .A(n44476), .B(n44475), .Z(n44474) );
  AND U44252 ( .A(n22710), .B(n22711), .Z(n44475) );
  IV U44253 ( .A(p_input[230]), .Z(n22711) );
  IV U44254 ( .A(p_input[231]), .Z(n22710) );
  XOR U44255 ( .A(n44478), .B(n44477), .Z(n44476) );
  AND U44256 ( .A(n22712), .B(n22713), .Z(n44477) );
  IV U44257 ( .A(p_input[228]), .Z(n22713) );
  IV U44258 ( .A(p_input[229]), .Z(n22712) );
  XOR U44259 ( .A(n44480), .B(n44479), .Z(n44478) );
  AND U44260 ( .A(n22714), .B(n22715), .Z(n44479) );
  IV U44261 ( .A(p_input[226]), .Z(n22715) );
  IV U44262 ( .A(p_input[227]), .Z(n22714) );
  XOR U44263 ( .A(n44482), .B(n44481), .Z(n44480) );
  AND U44264 ( .A(n22716), .B(n22717), .Z(n44481) );
  IV U44265 ( .A(p_input[224]), .Z(n22717) );
  IV U44266 ( .A(p_input[225]), .Z(n22716) );
  XOR U44267 ( .A(n44484), .B(n44483), .Z(n44482) );
  AND U44268 ( .A(n22718), .B(n22719), .Z(n44483) );
  IV U44269 ( .A(p_input[222]), .Z(n22719) );
  IV U44270 ( .A(p_input[223]), .Z(n22718) );
  XOR U44271 ( .A(n44486), .B(n44485), .Z(n44484) );
  AND U44272 ( .A(n22720), .B(n22721), .Z(n44485) );
  IV U44273 ( .A(p_input[220]), .Z(n22721) );
  IV U44274 ( .A(p_input[221]), .Z(n22720) );
  XOR U44275 ( .A(n44488), .B(n44487), .Z(n44486) );
  AND U44276 ( .A(n22722), .B(n22723), .Z(n44487) );
  IV U44277 ( .A(p_input[218]), .Z(n22723) );
  IV U44278 ( .A(p_input[219]), .Z(n22722) );
  XOR U44279 ( .A(n44490), .B(n44489), .Z(n44488) );
  AND U44280 ( .A(n22724), .B(n22725), .Z(n44489) );
  IV U44281 ( .A(p_input[216]), .Z(n22725) );
  IV U44282 ( .A(p_input[217]), .Z(n22724) );
  XOR U44283 ( .A(n44492), .B(n44491), .Z(n44490) );
  AND U44284 ( .A(n22726), .B(n22727), .Z(n44491) );
  IV U44285 ( .A(p_input[214]), .Z(n22727) );
  IV U44286 ( .A(p_input[215]), .Z(n22726) );
  XOR U44287 ( .A(n44494), .B(n44493), .Z(n44492) );
  AND U44288 ( .A(n22728), .B(n22729), .Z(n44493) );
  IV U44289 ( .A(p_input[212]), .Z(n22729) );
  IV U44290 ( .A(p_input[213]), .Z(n22728) );
  XOR U44291 ( .A(n44496), .B(n44495), .Z(n44494) );
  AND U44292 ( .A(n22730), .B(n22731), .Z(n44495) );
  IV U44293 ( .A(p_input[210]), .Z(n22731) );
  IV U44294 ( .A(p_input[211]), .Z(n22730) );
  XOR U44295 ( .A(n44498), .B(n44497), .Z(n44496) );
  AND U44296 ( .A(n22732), .B(n22733), .Z(n44497) );
  IV U44297 ( .A(p_input[208]), .Z(n22733) );
  IV U44298 ( .A(p_input[209]), .Z(n22732) );
  XOR U44299 ( .A(n44500), .B(n44499), .Z(n44498) );
  AND U44300 ( .A(n22734), .B(n22735), .Z(n44499) );
  IV U44301 ( .A(p_input[206]), .Z(n22735) );
  IV U44302 ( .A(p_input[207]), .Z(n22734) );
  XOR U44303 ( .A(n44502), .B(n44501), .Z(n44500) );
  AND U44304 ( .A(n22736), .B(n22737), .Z(n44501) );
  IV U44305 ( .A(p_input[204]), .Z(n22737) );
  IV U44306 ( .A(p_input[205]), .Z(n22736) );
  XOR U44307 ( .A(n44504), .B(n44503), .Z(n44502) );
  AND U44308 ( .A(n22738), .B(n22739), .Z(n44503) );
  IV U44309 ( .A(p_input[202]), .Z(n22739) );
  IV U44310 ( .A(p_input[203]), .Z(n22738) );
  XOR U44311 ( .A(n44506), .B(n44505), .Z(n44504) );
  AND U44312 ( .A(n22740), .B(n22741), .Z(n44505) );
  IV U44313 ( .A(p_input[200]), .Z(n22741) );
  IV U44314 ( .A(p_input[201]), .Z(n22740) );
  XOR U44315 ( .A(n44508), .B(n44507), .Z(n44506) );
  AND U44316 ( .A(n22742), .B(n22743), .Z(n44507) );
  IV U44317 ( .A(p_input[198]), .Z(n22743) );
  IV U44318 ( .A(p_input[199]), .Z(n22742) );
  XOR U44319 ( .A(n44510), .B(n44509), .Z(n44508) );
  AND U44320 ( .A(n22744), .B(n22745), .Z(n44509) );
  IV U44321 ( .A(p_input[196]), .Z(n22745) );
  IV U44322 ( .A(p_input[197]), .Z(n22744) );
  XOR U44323 ( .A(n44512), .B(n44511), .Z(n44510) );
  AND U44324 ( .A(n22746), .B(n22747), .Z(n44511) );
  IV U44325 ( .A(p_input[194]), .Z(n22747) );
  IV U44326 ( .A(p_input[195]), .Z(n22746) );
  XOR U44327 ( .A(n44514), .B(n44513), .Z(n44512) );
  AND U44328 ( .A(n22748), .B(n22749), .Z(n44513) );
  IV U44329 ( .A(p_input[192]), .Z(n22749) );
  IV U44330 ( .A(p_input[193]), .Z(n22748) );
  XOR U44331 ( .A(n44516), .B(n44515), .Z(n44514) );
  AND U44332 ( .A(n22750), .B(n22751), .Z(n44515) );
  IV U44333 ( .A(p_input[190]), .Z(n22751) );
  IV U44334 ( .A(p_input[191]), .Z(n22750) );
  XOR U44335 ( .A(n44518), .B(n44517), .Z(n44516) );
  AND U44336 ( .A(n22752), .B(n22753), .Z(n44517) );
  IV U44337 ( .A(p_input[188]), .Z(n22753) );
  IV U44338 ( .A(p_input[189]), .Z(n22752) );
  XOR U44339 ( .A(n44520), .B(n44519), .Z(n44518) );
  AND U44340 ( .A(n22754), .B(n22755), .Z(n44519) );
  IV U44341 ( .A(p_input[186]), .Z(n22755) );
  IV U44342 ( .A(p_input[187]), .Z(n22754) );
  XOR U44343 ( .A(n44522), .B(n44521), .Z(n44520) );
  AND U44344 ( .A(n22756), .B(n22757), .Z(n44521) );
  IV U44345 ( .A(p_input[184]), .Z(n22757) );
  IV U44346 ( .A(p_input[185]), .Z(n22756) );
  XOR U44347 ( .A(n44524), .B(n44523), .Z(n44522) );
  AND U44348 ( .A(n22758), .B(n22759), .Z(n44523) );
  IV U44349 ( .A(p_input[182]), .Z(n22759) );
  IV U44350 ( .A(p_input[183]), .Z(n22758) );
  XOR U44351 ( .A(n44526), .B(n44525), .Z(n44524) );
  AND U44352 ( .A(n22760), .B(n22761), .Z(n44525) );
  IV U44353 ( .A(p_input[180]), .Z(n22761) );
  IV U44354 ( .A(p_input[181]), .Z(n22760) );
  XOR U44355 ( .A(n44528), .B(n44527), .Z(n44526) );
  AND U44356 ( .A(n22762), .B(n22763), .Z(n44527) );
  IV U44357 ( .A(p_input[178]), .Z(n22763) );
  IV U44358 ( .A(p_input[179]), .Z(n22762) );
  XOR U44359 ( .A(n44530), .B(n44529), .Z(n44528) );
  AND U44360 ( .A(n22764), .B(n22765), .Z(n44529) );
  IV U44361 ( .A(p_input[176]), .Z(n22765) );
  IV U44362 ( .A(p_input[177]), .Z(n22764) );
  XOR U44363 ( .A(n44532), .B(n44531), .Z(n44530) );
  AND U44364 ( .A(n22766), .B(n22767), .Z(n44531) );
  IV U44365 ( .A(p_input[174]), .Z(n22767) );
  IV U44366 ( .A(p_input[175]), .Z(n22766) );
  XOR U44367 ( .A(n44534), .B(n44533), .Z(n44532) );
  AND U44368 ( .A(n22768), .B(n22769), .Z(n44533) );
  IV U44369 ( .A(p_input[172]), .Z(n22769) );
  IV U44370 ( .A(p_input[173]), .Z(n22768) );
  XOR U44371 ( .A(n44536), .B(n44535), .Z(n44534) );
  AND U44372 ( .A(n22770), .B(n22771), .Z(n44535) );
  IV U44373 ( .A(p_input[170]), .Z(n22771) );
  IV U44374 ( .A(p_input[171]), .Z(n22770) );
  XOR U44375 ( .A(n44538), .B(n44537), .Z(n44536) );
  AND U44376 ( .A(n22772), .B(n22773), .Z(n44537) );
  IV U44377 ( .A(p_input[168]), .Z(n22773) );
  IV U44378 ( .A(p_input[169]), .Z(n22772) );
  XOR U44379 ( .A(n44540), .B(n44539), .Z(n44538) );
  AND U44380 ( .A(n22774), .B(n22775), .Z(n44539) );
  IV U44381 ( .A(p_input[166]), .Z(n22775) );
  IV U44382 ( .A(p_input[167]), .Z(n22774) );
  XOR U44383 ( .A(n44542), .B(n44541), .Z(n44540) );
  AND U44384 ( .A(n22776), .B(n22777), .Z(n44541) );
  IV U44385 ( .A(p_input[164]), .Z(n22777) );
  IV U44386 ( .A(p_input[165]), .Z(n22776) );
  XOR U44387 ( .A(n44544), .B(n44543), .Z(n44542) );
  AND U44388 ( .A(n22778), .B(n22779), .Z(n44543) );
  IV U44389 ( .A(p_input[162]), .Z(n22779) );
  IV U44390 ( .A(p_input[163]), .Z(n22778) );
  XOR U44391 ( .A(n44546), .B(n44545), .Z(n44544) );
  AND U44392 ( .A(n22780), .B(n22781), .Z(n44545) );
  IV U44393 ( .A(p_input[160]), .Z(n22781) );
  IV U44394 ( .A(p_input[161]), .Z(n22780) );
  XOR U44395 ( .A(n44548), .B(n44547), .Z(n44546) );
  AND U44396 ( .A(n22782), .B(n22783), .Z(n44547) );
  IV U44397 ( .A(p_input[158]), .Z(n22783) );
  IV U44398 ( .A(p_input[159]), .Z(n22782) );
  XOR U44399 ( .A(n44550), .B(n44549), .Z(n44548) );
  AND U44400 ( .A(n22784), .B(n22785), .Z(n44549) );
  IV U44401 ( .A(p_input[156]), .Z(n22785) );
  IV U44402 ( .A(p_input[157]), .Z(n22784) );
  XOR U44403 ( .A(n44552), .B(n44551), .Z(n44550) );
  AND U44404 ( .A(n22786), .B(n22787), .Z(n44551) );
  IV U44405 ( .A(p_input[154]), .Z(n22787) );
  IV U44406 ( .A(p_input[155]), .Z(n22786) );
  XOR U44407 ( .A(n44554), .B(n44553), .Z(n44552) );
  AND U44408 ( .A(n22788), .B(n22789), .Z(n44553) );
  IV U44409 ( .A(p_input[152]), .Z(n22789) );
  IV U44410 ( .A(p_input[153]), .Z(n22788) );
  XOR U44411 ( .A(n44556), .B(n44555), .Z(n44554) );
  AND U44412 ( .A(n22790), .B(n22791), .Z(n44555) );
  IV U44413 ( .A(p_input[150]), .Z(n22791) );
  IV U44414 ( .A(p_input[151]), .Z(n22790) );
  XOR U44415 ( .A(n44558), .B(n44557), .Z(n44556) );
  AND U44416 ( .A(n22792), .B(n22793), .Z(n44557) );
  IV U44417 ( .A(p_input[148]), .Z(n22793) );
  IV U44418 ( .A(p_input[149]), .Z(n22792) );
  XOR U44419 ( .A(n44560), .B(n44559), .Z(n44558) );
  AND U44420 ( .A(n22794), .B(n22795), .Z(n44559) );
  IV U44421 ( .A(p_input[146]), .Z(n22795) );
  IV U44422 ( .A(p_input[147]), .Z(n22794) );
  XOR U44423 ( .A(n44562), .B(n44561), .Z(n44560) );
  AND U44424 ( .A(n22796), .B(n22797), .Z(n44561) );
  IV U44425 ( .A(p_input[144]), .Z(n22797) );
  IV U44426 ( .A(p_input[145]), .Z(n22796) );
  XOR U44427 ( .A(n44564), .B(n44563), .Z(n44562) );
  AND U44428 ( .A(n22798), .B(n22799), .Z(n44563) );
  IV U44429 ( .A(p_input[142]), .Z(n22799) );
  IV U44430 ( .A(p_input[143]), .Z(n22798) );
  XOR U44431 ( .A(n44566), .B(n44565), .Z(n44564) );
  AND U44432 ( .A(n22800), .B(n22801), .Z(n44565) );
  IV U44433 ( .A(p_input[140]), .Z(n22801) );
  IV U44434 ( .A(p_input[141]), .Z(n22800) );
  XOR U44435 ( .A(n44568), .B(n44567), .Z(n44566) );
  AND U44436 ( .A(n22802), .B(n22803), .Z(n44567) );
  IV U44437 ( .A(p_input[138]), .Z(n22803) );
  IV U44438 ( .A(p_input[139]), .Z(n22802) );
  XOR U44439 ( .A(n44570), .B(n44569), .Z(n44568) );
  AND U44440 ( .A(n22804), .B(n22805), .Z(n44569) );
  IV U44441 ( .A(p_input[136]), .Z(n22805) );
  IV U44442 ( .A(p_input[137]), .Z(n22804) );
  XOR U44443 ( .A(n44572), .B(n44571), .Z(n44570) );
  AND U44444 ( .A(n22806), .B(n22807), .Z(n44571) );
  IV U44445 ( .A(p_input[134]), .Z(n22807) );
  IV U44446 ( .A(p_input[135]), .Z(n22806) );
  XOR U44447 ( .A(n44574), .B(n44573), .Z(n44572) );
  AND U44448 ( .A(n22808), .B(n22809), .Z(n44573) );
  IV U44449 ( .A(p_input[132]), .Z(n22809) );
  IV U44450 ( .A(p_input[133]), .Z(n22808) );
  XOR U44451 ( .A(n44576), .B(n44575), .Z(n44574) );
  AND U44452 ( .A(n22810), .B(n22811), .Z(n44575) );
  IV U44453 ( .A(p_input[130]), .Z(n22811) );
  IV U44454 ( .A(p_input[131]), .Z(n22810) );
  XOR U44455 ( .A(n44578), .B(n44577), .Z(n44576) );
  AND U44456 ( .A(n22812), .B(n22813), .Z(n44577) );
  IV U44457 ( .A(p_input[128]), .Z(n22813) );
  IV U44458 ( .A(p_input[129]), .Z(n22812) );
  XOR U44459 ( .A(n44580), .B(n44579), .Z(n44578) );
  AND U44460 ( .A(n22814), .B(n22815), .Z(n44579) );
  IV U44461 ( .A(p_input[126]), .Z(n22815) );
  IV U44462 ( .A(p_input[127]), .Z(n22814) );
  XOR U44463 ( .A(n44582), .B(n44581), .Z(n44580) );
  AND U44464 ( .A(n22816), .B(n22817), .Z(n44581) );
  IV U44465 ( .A(p_input[124]), .Z(n22817) );
  IV U44466 ( .A(p_input[125]), .Z(n22816) );
  XOR U44467 ( .A(n44584), .B(n44583), .Z(n44582) );
  AND U44468 ( .A(n22818), .B(n22819), .Z(n44583) );
  IV U44469 ( .A(p_input[122]), .Z(n22819) );
  IV U44470 ( .A(p_input[123]), .Z(n22818) );
  XOR U44471 ( .A(n44586), .B(n44585), .Z(n44584) );
  AND U44472 ( .A(n22820), .B(n22821), .Z(n44585) );
  IV U44473 ( .A(p_input[120]), .Z(n22821) );
  IV U44474 ( .A(p_input[121]), .Z(n22820) );
  XOR U44475 ( .A(n44588), .B(n44587), .Z(n44586) );
  AND U44476 ( .A(n22822), .B(n22823), .Z(n44587) );
  IV U44477 ( .A(p_input[118]), .Z(n22823) );
  IV U44478 ( .A(p_input[119]), .Z(n22822) );
  XOR U44479 ( .A(n44590), .B(n44589), .Z(n44588) );
  AND U44480 ( .A(n22824), .B(n22825), .Z(n44589) );
  IV U44481 ( .A(p_input[116]), .Z(n22825) );
  IV U44482 ( .A(p_input[117]), .Z(n22824) );
  XOR U44483 ( .A(n44592), .B(n44591), .Z(n44590) );
  AND U44484 ( .A(n22826), .B(n22827), .Z(n44591) );
  IV U44485 ( .A(p_input[114]), .Z(n22827) );
  IV U44486 ( .A(p_input[115]), .Z(n22826) );
  XOR U44487 ( .A(n44594), .B(n44593), .Z(n44592) );
  AND U44488 ( .A(n22828), .B(n22829), .Z(n44593) );
  IV U44489 ( .A(p_input[112]), .Z(n22829) );
  IV U44490 ( .A(p_input[113]), .Z(n22828) );
  XOR U44491 ( .A(n44596), .B(n44595), .Z(n44594) );
  AND U44492 ( .A(n22830), .B(n22831), .Z(n44595) );
  IV U44493 ( .A(p_input[110]), .Z(n22831) );
  IV U44494 ( .A(p_input[111]), .Z(n22830) );
  XOR U44495 ( .A(n44598), .B(n44597), .Z(n44596) );
  AND U44496 ( .A(n22832), .B(n22833), .Z(n44597) );
  IV U44497 ( .A(p_input[108]), .Z(n22833) );
  IV U44498 ( .A(p_input[109]), .Z(n22832) );
  XOR U44499 ( .A(n44600), .B(n44599), .Z(n44598) );
  AND U44500 ( .A(n22834), .B(n22835), .Z(n44599) );
  IV U44501 ( .A(p_input[106]), .Z(n22835) );
  IV U44502 ( .A(p_input[107]), .Z(n22834) );
  XOR U44503 ( .A(n44602), .B(n44601), .Z(n44600) );
  AND U44504 ( .A(n22836), .B(n22837), .Z(n44601) );
  IV U44505 ( .A(p_input[104]), .Z(n22837) );
  IV U44506 ( .A(p_input[105]), .Z(n22836) );
  XOR U44507 ( .A(n44604), .B(n44603), .Z(n44602) );
  AND U44508 ( .A(n22838), .B(n22839), .Z(n44603) );
  IV U44509 ( .A(p_input[102]), .Z(n22839) );
  IV U44510 ( .A(p_input[103]), .Z(n22838) );
  XOR U44511 ( .A(n44606), .B(n44605), .Z(n44604) );
  AND U44512 ( .A(n22840), .B(n22841), .Z(n44605) );
  IV U44513 ( .A(p_input[100]), .Z(n22841) );
  IV U44514 ( .A(p_input[101]), .Z(n22840) );
  XOR U44515 ( .A(n44608), .B(n44607), .Z(n44606) );
  AND U44516 ( .A(n22842), .B(n22843), .Z(n44607) );
  IV U44517 ( .A(p_input[98]), .Z(n22843) );
  IV U44518 ( .A(p_input[99]), .Z(n22842) );
  XOR U44519 ( .A(n44610), .B(n44609), .Z(n44608) );
  AND U44520 ( .A(n22844), .B(n22845), .Z(n44609) );
  IV U44521 ( .A(p_input[96]), .Z(n22845) );
  IV U44522 ( .A(p_input[97]), .Z(n22844) );
  XOR U44523 ( .A(n44612), .B(n44611), .Z(n44610) );
  AND U44524 ( .A(n22846), .B(n22847), .Z(n44611) );
  IV U44525 ( .A(p_input[94]), .Z(n22847) );
  IV U44526 ( .A(p_input[95]), .Z(n22846) );
  XOR U44527 ( .A(n44614), .B(n44613), .Z(n44612) );
  AND U44528 ( .A(n22848), .B(n22849), .Z(n44613) );
  IV U44529 ( .A(p_input[92]), .Z(n22849) );
  IV U44530 ( .A(p_input[93]), .Z(n22848) );
  XOR U44531 ( .A(n44616), .B(n44615), .Z(n44614) );
  AND U44532 ( .A(n22850), .B(n22851), .Z(n44615) );
  IV U44533 ( .A(p_input[90]), .Z(n22851) );
  IV U44534 ( .A(p_input[91]), .Z(n22850) );
  XOR U44535 ( .A(n44618), .B(n44617), .Z(n44616) );
  AND U44536 ( .A(n22852), .B(n22853), .Z(n44617) );
  IV U44537 ( .A(p_input[88]), .Z(n22853) );
  IV U44538 ( .A(p_input[89]), .Z(n22852) );
  XOR U44539 ( .A(n44620), .B(n44619), .Z(n44618) );
  AND U44540 ( .A(n22854), .B(n22855), .Z(n44619) );
  IV U44541 ( .A(p_input[86]), .Z(n22855) );
  IV U44542 ( .A(p_input[87]), .Z(n22854) );
  XOR U44543 ( .A(n44622), .B(n44621), .Z(n44620) );
  AND U44544 ( .A(n22856), .B(n22857), .Z(n44621) );
  IV U44545 ( .A(p_input[84]), .Z(n22857) );
  IV U44546 ( .A(p_input[85]), .Z(n22856) );
  XOR U44547 ( .A(n44624), .B(n44623), .Z(n44622) );
  AND U44548 ( .A(n22858), .B(n22859), .Z(n44623) );
  IV U44549 ( .A(p_input[82]), .Z(n22859) );
  IV U44550 ( .A(p_input[83]), .Z(n22858) );
  XOR U44551 ( .A(n44626), .B(n44625), .Z(n44624) );
  AND U44552 ( .A(n22860), .B(n22861), .Z(n44625) );
  IV U44553 ( .A(p_input[80]), .Z(n22861) );
  IV U44554 ( .A(p_input[81]), .Z(n22860) );
  XOR U44555 ( .A(n44628), .B(n44627), .Z(n44626) );
  AND U44556 ( .A(n22862), .B(n22863), .Z(n44627) );
  IV U44557 ( .A(p_input[78]), .Z(n22863) );
  IV U44558 ( .A(p_input[79]), .Z(n22862) );
  XOR U44559 ( .A(n44630), .B(n44629), .Z(n44628) );
  AND U44560 ( .A(n22864), .B(n22865), .Z(n44629) );
  IV U44561 ( .A(p_input[76]), .Z(n22865) );
  IV U44562 ( .A(p_input[77]), .Z(n22864) );
  XOR U44563 ( .A(n44632), .B(n44631), .Z(n44630) );
  AND U44564 ( .A(n22866), .B(n22867), .Z(n44631) );
  IV U44565 ( .A(p_input[74]), .Z(n22867) );
  IV U44566 ( .A(p_input[75]), .Z(n22866) );
  XOR U44567 ( .A(n44634), .B(n44633), .Z(n44632) );
  AND U44568 ( .A(n22868), .B(n22869), .Z(n44633) );
  IV U44569 ( .A(p_input[72]), .Z(n22869) );
  IV U44570 ( .A(p_input[73]), .Z(n22868) );
  XOR U44571 ( .A(n44636), .B(n44635), .Z(n44634) );
  AND U44572 ( .A(n22870), .B(n22871), .Z(n44635) );
  IV U44573 ( .A(p_input[70]), .Z(n22871) );
  IV U44574 ( .A(p_input[71]), .Z(n22870) );
  XOR U44575 ( .A(n44638), .B(n44637), .Z(n44636) );
  AND U44576 ( .A(n22872), .B(n22873), .Z(n44637) );
  IV U44577 ( .A(p_input[68]), .Z(n22873) );
  IV U44578 ( .A(p_input[69]), .Z(n22872) );
  XOR U44579 ( .A(n44640), .B(n44639), .Z(n44638) );
  AND U44580 ( .A(n22874), .B(n22875), .Z(n44639) );
  IV U44581 ( .A(p_input[66]), .Z(n22875) );
  IV U44582 ( .A(p_input[67]), .Z(n22874) );
  XOR U44583 ( .A(n44642), .B(n44641), .Z(n44640) );
  AND U44584 ( .A(n22876), .B(n22877), .Z(n44641) );
  IV U44585 ( .A(p_input[64]), .Z(n22877) );
  IV U44586 ( .A(p_input[65]), .Z(n22876) );
  XOR U44587 ( .A(n44644), .B(n44643), .Z(n44642) );
  AND U44588 ( .A(n22878), .B(n22879), .Z(n44643) );
  IV U44589 ( .A(p_input[62]), .Z(n22879) );
  IV U44590 ( .A(p_input[63]), .Z(n22878) );
  XOR U44591 ( .A(n44646), .B(n44645), .Z(n44644) );
  AND U44592 ( .A(n22880), .B(n22881), .Z(n44645) );
  IV U44593 ( .A(p_input[60]), .Z(n22881) );
  IV U44594 ( .A(p_input[61]), .Z(n22880) );
  XOR U44595 ( .A(n44648), .B(n44647), .Z(n44646) );
  AND U44596 ( .A(n22882), .B(n22883), .Z(n44647) );
  IV U44597 ( .A(p_input[58]), .Z(n22883) );
  IV U44598 ( .A(p_input[59]), .Z(n22882) );
  XOR U44599 ( .A(n44650), .B(n44649), .Z(n44648) );
  AND U44600 ( .A(n22884), .B(n22885), .Z(n44649) );
  IV U44601 ( .A(p_input[56]), .Z(n22885) );
  IV U44602 ( .A(p_input[57]), .Z(n22884) );
  XOR U44603 ( .A(n44652), .B(n44651), .Z(n44650) );
  AND U44604 ( .A(n22886), .B(n22887), .Z(n44651) );
  IV U44605 ( .A(p_input[54]), .Z(n22887) );
  IV U44606 ( .A(p_input[55]), .Z(n22886) );
  XOR U44607 ( .A(n44654), .B(n44653), .Z(n44652) );
  AND U44608 ( .A(n22888), .B(n22889), .Z(n44653) );
  IV U44609 ( .A(p_input[52]), .Z(n22889) );
  IV U44610 ( .A(p_input[53]), .Z(n22888) );
  XOR U44611 ( .A(n44656), .B(n44655), .Z(n44654) );
  AND U44612 ( .A(n22890), .B(n22891), .Z(n44655) );
  IV U44613 ( .A(p_input[50]), .Z(n22891) );
  IV U44614 ( .A(p_input[51]), .Z(n22890) );
  XOR U44615 ( .A(n44658), .B(n44657), .Z(n44656) );
  AND U44616 ( .A(n22892), .B(n22893), .Z(n44657) );
  IV U44617 ( .A(p_input[48]), .Z(n22893) );
  IV U44618 ( .A(p_input[49]), .Z(n22892) );
  XOR U44619 ( .A(n44660), .B(n44659), .Z(n44658) );
  AND U44620 ( .A(n22894), .B(n22895), .Z(n44659) );
  IV U44621 ( .A(p_input[46]), .Z(n22895) );
  IV U44622 ( .A(p_input[47]), .Z(n22894) );
  XOR U44623 ( .A(n44662), .B(n44661), .Z(n44660) );
  AND U44624 ( .A(n22896), .B(n22897), .Z(n44661) );
  IV U44625 ( .A(p_input[44]), .Z(n22897) );
  IV U44626 ( .A(p_input[45]), .Z(n22896) );
  XOR U44627 ( .A(n44664), .B(n44663), .Z(n44662) );
  AND U44628 ( .A(n22898), .B(n22899), .Z(n44663) );
  IV U44629 ( .A(p_input[42]), .Z(n22899) );
  IV U44630 ( .A(p_input[43]), .Z(n22898) );
  XOR U44631 ( .A(n44666), .B(n44665), .Z(n44664) );
  AND U44632 ( .A(n22900), .B(n22901), .Z(n44665) );
  IV U44633 ( .A(p_input[40]), .Z(n22901) );
  IV U44634 ( .A(p_input[41]), .Z(n22900) );
  XOR U44635 ( .A(n44668), .B(n44667), .Z(n44666) );
  AND U44636 ( .A(n22902), .B(n22903), .Z(n44667) );
  IV U44637 ( .A(p_input[38]), .Z(n22903) );
  IV U44638 ( .A(p_input[39]), .Z(n22902) );
  XOR U44639 ( .A(n44670), .B(n44669), .Z(n44668) );
  AND U44640 ( .A(n22904), .B(n22905), .Z(n44669) );
  IV U44641 ( .A(p_input[36]), .Z(n22905) );
  IV U44642 ( .A(p_input[37]), .Z(n22904) );
  XOR U44643 ( .A(n44672), .B(n44671), .Z(n44670) );
  AND U44644 ( .A(n22906), .B(n22907), .Z(n44671) );
  IV U44645 ( .A(p_input[34]), .Z(n22907) );
  IV U44646 ( .A(p_input[35]), .Z(n22906) );
  XOR U44647 ( .A(n44674), .B(n44673), .Z(n44672) );
  AND U44648 ( .A(n22908), .B(n22909), .Z(n44673) );
  IV U44649 ( .A(p_input[32]), .Z(n22909) );
  IV U44650 ( .A(p_input[33]), .Z(n22908) );
  XOR U44651 ( .A(n44676), .B(n44675), .Z(n44674) );
  AND U44652 ( .A(n22910), .B(n22911), .Z(n44675) );
  IV U44653 ( .A(p_input[30]), .Z(n22911) );
  IV U44654 ( .A(p_input[31]), .Z(n22910) );
  XOR U44655 ( .A(n44678), .B(n44677), .Z(n44676) );
  AND U44656 ( .A(n22912), .B(n22913), .Z(n44677) );
  IV U44657 ( .A(p_input[28]), .Z(n22913) );
  IV U44658 ( .A(p_input[29]), .Z(n22912) );
  XOR U44659 ( .A(n44680), .B(n44679), .Z(n44678) );
  AND U44660 ( .A(n22914), .B(n22915), .Z(n44679) );
  IV U44661 ( .A(p_input[26]), .Z(n22915) );
  IV U44662 ( .A(p_input[27]), .Z(n22914) );
  XOR U44663 ( .A(n44682), .B(n44681), .Z(n44680) );
  AND U44664 ( .A(n22916), .B(n22917), .Z(n44681) );
  IV U44665 ( .A(p_input[24]), .Z(n22917) );
  IV U44666 ( .A(p_input[25]), .Z(n22916) );
  XOR U44667 ( .A(n44684), .B(n44683), .Z(n44682) );
  AND U44668 ( .A(n22918), .B(n22919), .Z(n44683) );
  IV U44669 ( .A(p_input[22]), .Z(n22919) );
  IV U44670 ( .A(p_input[23]), .Z(n22918) );
  XOR U44671 ( .A(n44686), .B(n44685), .Z(n44684) );
  AND U44672 ( .A(n22920), .B(n22921), .Z(n44685) );
  IV U44673 ( .A(p_input[20]), .Z(n22921) );
  IV U44674 ( .A(p_input[21]), .Z(n22920) );
  XOR U44675 ( .A(n44688), .B(n44687), .Z(n44686) );
  AND U44676 ( .A(n22922), .B(n22923), .Z(n44687) );
  IV U44677 ( .A(p_input[18]), .Z(n22923) );
  IV U44678 ( .A(p_input[19]), .Z(n22922) );
  XOR U44679 ( .A(n44690), .B(n44689), .Z(n44688) );
  AND U44680 ( .A(n22924), .B(n22925), .Z(n44689) );
  IV U44681 ( .A(p_input[16]), .Z(n22925) );
  IV U44682 ( .A(p_input[17]), .Z(n22924) );
  XOR U44683 ( .A(n44692), .B(n44691), .Z(n44690) );
  AND U44684 ( .A(n22926), .B(n22927), .Z(n44691) );
  IV U44685 ( .A(p_input[14]), .Z(n22927) );
  IV U44686 ( .A(p_input[15]), .Z(n22926) );
  XOR U44687 ( .A(n44694), .B(n44693), .Z(n44692) );
  AND U44688 ( .A(n22928), .B(n22929), .Z(n44693) );
  IV U44689 ( .A(p_input[12]), .Z(n22929) );
  IV U44690 ( .A(p_input[13]), .Z(n22928) );
  XOR U44691 ( .A(n44708), .B(n44707), .Z(n44694) );
  AND U44692 ( .A(n22930), .B(n22931), .Z(n44707) );
  IV U44693 ( .A(p_input[10]), .Z(n22931) );
  IV U44694 ( .A(p_input[11]), .Z(n22930) );
  XOR U44695 ( .A(n44710), .B(n44709), .Z(n44708) );
  AND U44696 ( .A(n22932), .B(n22933), .Z(n44709) );
  IV U44697 ( .A(p_input[8]), .Z(n22933) );
  IV U44698 ( .A(p_input[9]), .Z(n22932) );
  XOR U44699 ( .A(n44698), .B(n44697), .Z(n44710) );
  AND U44700 ( .A(n22934), .B(n22935), .Z(n44697) );
  IV U44701 ( .A(p_input[6]), .Z(n22935) );
  IV U44702 ( .A(p_input[7]), .Z(n22934) );
  XOR U44703 ( .A(n44705), .B(n44706), .Z(n44698) );
  XOR U44704 ( .A(n44703), .B(n44704), .Z(n44706) );
  AND U44705 ( .A(n22936), .B(n22937), .Z(n44704) );
  IV U44706 ( .A(p_input[2]), .Z(n22937) );
  IV U44707 ( .A(p_input[3]), .Z(n22936) );
  AND U44708 ( .A(n22938), .B(n22939), .Z(n44703) );
  IV U44709 ( .A(p_input[0]), .Z(n22939) );
  IV U44710 ( .A(p_input[1]), .Z(n22938) );
  AND U44711 ( .A(n22940), .B(n22941), .Z(n44705) );
  IV U44712 ( .A(p_input[4]), .Z(n22941) );
  IV U44713 ( .A(p_input[5]), .Z(n22940) );
endmodule

