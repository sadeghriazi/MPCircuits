
module voting_N2_M8 ( p_input, o );
  input [511:0] p_input;
  output [1:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529;

  XOR U2 ( .A(n1), .B(n2), .Z(o[0]) );
  AND U3 ( .A(o[1]), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(n5), .Z(n3) );
  IV U5 ( .A(n1), .Z(n5) );
  XNOR U6 ( .A(n6), .B(n7), .Z(o[1]) );
  AND U7 ( .A(n8), .B(n9), .Z(n7) );
  XOR U8 ( .A(n6), .B(n10), .Z(n9) );
  XOR U9 ( .A(n11), .B(n12), .Z(n10) );
  AND U10 ( .A(n4), .B(n13), .Z(n11) );
  XNOR U11 ( .A(n14), .B(n12), .Z(n13) );
  XOR U12 ( .A(n15), .B(n6), .Z(n8) );
  XOR U13 ( .A(n16), .B(n17), .Z(n15) );
  AND U14 ( .A(n1), .B(n18), .Z(n17) );
  XNOR U15 ( .A(n19), .B(n20), .Z(n18) );
  XOR U16 ( .A(n21), .B(n22), .Z(n6) );
  AND U17 ( .A(n23), .B(n24), .Z(n22) );
  XOR U18 ( .A(n21), .B(n25), .Z(n24) );
  XNOR U19 ( .A(n26), .B(n27), .Z(n25) );
  AND U20 ( .A(n4), .B(n28), .Z(n26) );
  XNOR U21 ( .A(n29), .B(n27), .Z(n28) );
  XOR U22 ( .A(n30), .B(n21), .Z(n23) );
  XOR U23 ( .A(n31), .B(n32), .Z(n30) );
  AND U24 ( .A(n1), .B(n33), .Z(n32) );
  XOR U25 ( .A(n34), .B(n35), .Z(n33) );
  XOR U26 ( .A(n36), .B(n37), .Z(n21) );
  AND U27 ( .A(n38), .B(n39), .Z(n37) );
  XOR U28 ( .A(n40), .B(n36), .Z(n39) );
  XNOR U29 ( .A(n41), .B(n42), .Z(n40) );
  AND U30 ( .A(n4), .B(n43), .Z(n42) );
  XOR U31 ( .A(n44), .B(n41), .Z(n43) );
  XOR U32 ( .A(n36), .B(n45), .Z(n38) );
  XNOR U33 ( .A(n46), .B(n47), .Z(n45) );
  AND U34 ( .A(n1), .B(n48), .Z(n46) );
  XNOR U35 ( .A(n49), .B(n47), .Z(n48) );
  XOR U36 ( .A(n50), .B(n51), .Z(n36) );
  AND U37 ( .A(n52), .B(n53), .Z(n51) );
  XOR U38 ( .A(n50), .B(n54), .Z(n53) );
  XNOR U39 ( .A(n55), .B(n56), .Z(n54) );
  AND U40 ( .A(n4), .B(n57), .Z(n55) );
  XNOR U41 ( .A(n58), .B(n56), .Z(n57) );
  XOR U42 ( .A(n59), .B(n50), .Z(n52) );
  XOR U43 ( .A(n60), .B(n61), .Z(n59) );
  AND U44 ( .A(n1), .B(n62), .Z(n61) );
  XOR U45 ( .A(n63), .B(n64), .Z(n62) );
  IV U46 ( .A(n60), .Z(n64) );
  XOR U47 ( .A(n65), .B(n66), .Z(n50) );
  AND U48 ( .A(n67), .B(n68), .Z(n66) );
  XOR U49 ( .A(n65), .B(n69), .Z(n68) );
  XNOR U50 ( .A(n70), .B(n71), .Z(n69) );
  AND U51 ( .A(n4), .B(n72), .Z(n70) );
  XNOR U52 ( .A(n73), .B(n71), .Z(n72) );
  XOR U53 ( .A(n74), .B(n65), .Z(n67) );
  XOR U54 ( .A(n75), .B(n76), .Z(n74) );
  AND U55 ( .A(n1), .B(n77), .Z(n76) );
  XOR U56 ( .A(n78), .B(n79), .Z(n77) );
  IV U57 ( .A(n75), .Z(n79) );
  XOR U58 ( .A(n80), .B(n81), .Z(n65) );
  AND U59 ( .A(n82), .B(n83), .Z(n81) );
  XOR U60 ( .A(n80), .B(n84), .Z(n83) );
  XNOR U61 ( .A(n85), .B(n86), .Z(n84) );
  AND U62 ( .A(n4), .B(n87), .Z(n85) );
  XNOR U63 ( .A(n88), .B(n86), .Z(n87) );
  XOR U64 ( .A(n89), .B(n80), .Z(n82) );
  XOR U65 ( .A(n90), .B(n91), .Z(n89) );
  AND U66 ( .A(n1), .B(n92), .Z(n91) );
  XOR U67 ( .A(n93), .B(n94), .Z(n92) );
  IV U68 ( .A(n90), .Z(n94) );
  XOR U69 ( .A(n95), .B(n96), .Z(n80) );
  AND U70 ( .A(n97), .B(n98), .Z(n96) );
  XOR U71 ( .A(n95), .B(n99), .Z(n98) );
  XNOR U72 ( .A(n100), .B(n101), .Z(n99) );
  AND U73 ( .A(n4), .B(n102), .Z(n100) );
  XNOR U74 ( .A(n103), .B(n101), .Z(n102) );
  XOR U75 ( .A(n104), .B(n95), .Z(n97) );
  XOR U76 ( .A(n105), .B(n106), .Z(n104) );
  AND U77 ( .A(n1), .B(n107), .Z(n106) );
  XOR U78 ( .A(n108), .B(n109), .Z(n107) );
  IV U79 ( .A(n105), .Z(n109) );
  XOR U80 ( .A(n110), .B(n111), .Z(n95) );
  AND U81 ( .A(n112), .B(n113), .Z(n111) );
  XOR U82 ( .A(n114), .B(n115), .Z(n113) );
  XOR U83 ( .A(n110), .B(n116), .Z(n115) );
  AND U84 ( .A(n4), .B(n117), .Z(n116) );
  XOR U85 ( .A(n114), .B(n118), .Z(n117) );
  XNOR U86 ( .A(n119), .B(n120), .Z(n112) );
  XOR U87 ( .A(n110), .B(n121), .Z(n120) );
  AND U88 ( .A(n1), .B(n122), .Z(n121) );
  XOR U89 ( .A(n123), .B(n119), .Z(n122) );
  AND U90 ( .A(n124), .B(n125), .Z(n110) );
  XNOR U91 ( .A(n126), .B(n127), .Z(n125) );
  AND U92 ( .A(n4), .B(n128), .Z(n126) );
  XNOR U93 ( .A(n129), .B(n127), .Z(n128) );
  XNOR U94 ( .A(n130), .B(n131), .Z(n4) );
  AND U95 ( .A(n132), .B(n133), .Z(n131) );
  XNOR U96 ( .A(n130), .B(n14), .Z(n133) );
  XOR U97 ( .A(n134), .B(n135), .Z(n14) );
  AND U98 ( .A(n136), .B(n137), .Z(n135) );
  XNOR U99 ( .A(n29), .B(n134), .Z(n136) );
  XNOR U100 ( .A(n138), .B(n139), .Z(n134) );
  AND U101 ( .A(n29), .B(n138), .Z(n139) );
  XNOR U102 ( .A(n12), .B(n130), .Z(n132) );
  XOR U103 ( .A(n140), .B(n141), .Z(n12) );
  AND U104 ( .A(n142), .B(n143), .Z(n141) );
  XOR U105 ( .A(n144), .B(n140), .Z(n142) );
  XOR U106 ( .A(n145), .B(n146), .Z(n140) );
  NOR U107 ( .A(n27), .B(n147), .Z(n146) );
  IV U108 ( .A(n145), .Z(n147) );
  IV U109 ( .A(n144), .Z(n27) );
  XOR U110 ( .A(n148), .B(n149), .Z(n130) );
  AND U111 ( .A(n150), .B(n151), .Z(n149) );
  XOR U112 ( .A(n148), .B(n29), .Z(n151) );
  XOR U113 ( .A(n138), .B(n137), .Z(n29) );
  XNOR U114 ( .A(n152), .B(n153), .Z(n137) );
  XOR U115 ( .A(n154), .B(n155), .Z(n153) );
  XOR U116 ( .A(n156), .B(n157), .Z(n155) );
  NOR U117 ( .A(n158), .B(n159), .Z(n157) );
  NOR U118 ( .A(n160), .B(n161), .Z(n156) );
  NOR U119 ( .A(n162), .B(n163), .Z(n154) );
  XOR U120 ( .A(n164), .B(n165), .Z(n152) );
  XOR U121 ( .A(n166), .B(n167), .Z(n165) );
  XOR U122 ( .A(n168), .B(n169), .Z(n167) );
  XNOR U123 ( .A(n170), .B(n171), .Z(n169) );
  XOR U124 ( .A(n172), .B(n173), .Z(n171) );
  XOR U125 ( .A(n174), .B(n175), .Z(n173) );
  XOR U126 ( .A(n176), .B(n177), .Z(n175) );
  XOR U127 ( .A(n178), .B(n179), .Z(n174) );
  XOR U128 ( .A(n180), .B(n181), .Z(n179) );
  XOR U129 ( .A(n182), .B(n183), .Z(n181) );
  XOR U130 ( .A(n184), .B(n185), .Z(n183) );
  XOR U131 ( .A(n186), .B(n187), .Z(n185) );
  XNOR U132 ( .A(n188), .B(n189), .Z(n184) );
  XNOR U133 ( .A(n190), .B(n191), .Z(n189) );
  NOR U134 ( .A(n192), .B(n187), .Z(n190) );
  XOR U135 ( .A(n193), .B(n194), .Z(n182) );
  XOR U136 ( .A(n195), .B(n196), .Z(n194) );
  XNOR U137 ( .A(n197), .B(n198), .Z(n196) );
  XOR U138 ( .A(n199), .B(n200), .Z(n198) );
  XOR U139 ( .A(n201), .B(n202), .Z(n200) );
  XOR U140 ( .A(n203), .B(n204), .Z(n202) );
  XOR U141 ( .A(n205), .B(n206), .Z(n201) );
  XOR U142 ( .A(n207), .B(n208), .Z(n206) );
  XOR U143 ( .A(n209), .B(n210), .Z(n208) );
  XOR U144 ( .A(n211), .B(n212), .Z(n210) );
  XOR U145 ( .A(n213), .B(n214), .Z(n212) );
  XNOR U146 ( .A(n215), .B(n216), .Z(n211) );
  XNOR U147 ( .A(n217), .B(n218), .Z(n216) );
  NOR U148 ( .A(n219), .B(n214), .Z(n217) );
  XOR U149 ( .A(n220), .B(n221), .Z(n209) );
  XOR U150 ( .A(n222), .B(n223), .Z(n221) );
  XNOR U151 ( .A(n224), .B(n225), .Z(n223) );
  XOR U152 ( .A(n226), .B(n227), .Z(n225) );
  XOR U153 ( .A(n228), .B(n229), .Z(n227) );
  XOR U154 ( .A(n230), .B(n231), .Z(n229) );
  XOR U155 ( .A(n232), .B(n233), .Z(n228) );
  XOR U156 ( .A(n234), .B(n235), .Z(n233) );
  XOR U157 ( .A(n236), .B(n237), .Z(n235) );
  XOR U158 ( .A(n238), .B(n239), .Z(n237) );
  XOR U159 ( .A(n240), .B(n241), .Z(n239) );
  XNOR U160 ( .A(n242), .B(n243), .Z(n238) );
  XNOR U161 ( .A(n244), .B(n245), .Z(n243) );
  NOR U162 ( .A(n246), .B(n241), .Z(n244) );
  XOR U163 ( .A(n247), .B(n248), .Z(n236) );
  XOR U164 ( .A(n249), .B(n250), .Z(n248) );
  XNOR U165 ( .A(n251), .B(n252), .Z(n250) );
  XOR U166 ( .A(n253), .B(n254), .Z(n252) );
  XOR U167 ( .A(n255), .B(n256), .Z(n254) );
  XOR U168 ( .A(n257), .B(n258), .Z(n256) );
  XOR U169 ( .A(n259), .B(n260), .Z(n255) );
  XOR U170 ( .A(n261), .B(n262), .Z(n260) );
  XOR U171 ( .A(n263), .B(n264), .Z(n262) );
  XOR U172 ( .A(n265), .B(n266), .Z(n264) );
  XOR U173 ( .A(n267), .B(n268), .Z(n266) );
  XNOR U174 ( .A(n269), .B(n270), .Z(n265) );
  XNOR U175 ( .A(n271), .B(n272), .Z(n270) );
  NOR U176 ( .A(n273), .B(n268), .Z(n271) );
  XOR U177 ( .A(n274), .B(n275), .Z(n263) );
  XOR U178 ( .A(n276), .B(n277), .Z(n275) );
  XNOR U179 ( .A(n278), .B(n279), .Z(n277) );
  XOR U180 ( .A(n280), .B(n281), .Z(n279) );
  XOR U181 ( .A(n282), .B(n283), .Z(n281) );
  XOR U182 ( .A(n284), .B(n285), .Z(n283) );
  XOR U183 ( .A(n286), .B(n287), .Z(n282) );
  XOR U184 ( .A(n288), .B(n289), .Z(n287) );
  XOR U185 ( .A(n290), .B(n291), .Z(n289) );
  XOR U186 ( .A(n292), .B(n293), .Z(n291) );
  XOR U187 ( .A(n294), .B(n295), .Z(n293) );
  XNOR U188 ( .A(n296), .B(n297), .Z(n292) );
  XNOR U189 ( .A(n298), .B(n299), .Z(n297) );
  NOR U190 ( .A(n300), .B(n295), .Z(n298) );
  XOR U191 ( .A(n301), .B(n302), .Z(n290) );
  XOR U192 ( .A(n303), .B(n304), .Z(n302) );
  XNOR U193 ( .A(n305), .B(n306), .Z(n304) );
  XOR U194 ( .A(n307), .B(n308), .Z(n306) );
  XOR U195 ( .A(n309), .B(n310), .Z(n308) );
  XOR U196 ( .A(n311), .B(n312), .Z(n310) );
  XOR U197 ( .A(n313), .B(n314), .Z(n309) );
  XOR U198 ( .A(n315), .B(n316), .Z(n314) );
  XOR U199 ( .A(n317), .B(n318), .Z(n316) );
  XOR U200 ( .A(n319), .B(n320), .Z(n318) );
  XOR U201 ( .A(n321), .B(n322), .Z(n320) );
  XNOR U202 ( .A(n323), .B(n324), .Z(n319) );
  XNOR U203 ( .A(n325), .B(n326), .Z(n324) );
  NOR U204 ( .A(n327), .B(n322), .Z(n325) );
  XOR U205 ( .A(n328), .B(n329), .Z(n317) );
  XOR U206 ( .A(n330), .B(n331), .Z(n329) );
  XNOR U207 ( .A(n332), .B(n333), .Z(n331) );
  XOR U208 ( .A(n334), .B(n335), .Z(n333) );
  XOR U209 ( .A(n336), .B(n337), .Z(n335) );
  XOR U210 ( .A(n338), .B(n339), .Z(n337) );
  XOR U211 ( .A(n340), .B(n341), .Z(n336) );
  XOR U212 ( .A(n342), .B(n343), .Z(n341) );
  XOR U213 ( .A(n344), .B(n345), .Z(n343) );
  XOR U214 ( .A(n346), .B(n347), .Z(n345) );
  XOR U215 ( .A(n348), .B(n349), .Z(n347) );
  XNOR U216 ( .A(n350), .B(n351), .Z(n346) );
  XNOR U217 ( .A(n352), .B(n353), .Z(n351) );
  NOR U218 ( .A(n354), .B(n349), .Z(n352) );
  XOR U219 ( .A(n355), .B(n356), .Z(n344) );
  XOR U220 ( .A(n357), .B(n358), .Z(n356) );
  XNOR U221 ( .A(n359), .B(n360), .Z(n358) );
  XOR U222 ( .A(n361), .B(n362), .Z(n360) );
  XOR U223 ( .A(n363), .B(n364), .Z(n362) );
  XOR U224 ( .A(n365), .B(n366), .Z(n364) );
  XOR U225 ( .A(n367), .B(n368), .Z(n363) );
  XOR U226 ( .A(n369), .B(n370), .Z(n368) );
  XOR U227 ( .A(n371), .B(n372), .Z(n370) );
  XOR U228 ( .A(n373), .B(n374), .Z(n372) );
  XOR U229 ( .A(n375), .B(n376), .Z(n374) );
  XNOR U230 ( .A(n377), .B(n378), .Z(n373) );
  XNOR U231 ( .A(n379), .B(n380), .Z(n378) );
  NOR U232 ( .A(n381), .B(n376), .Z(n379) );
  XOR U233 ( .A(n382), .B(n383), .Z(n371) );
  XOR U234 ( .A(n384), .B(n385), .Z(n383) );
  XNOR U235 ( .A(n386), .B(n387), .Z(n385) );
  XOR U236 ( .A(n388), .B(n389), .Z(n387) );
  XOR U237 ( .A(n390), .B(n391), .Z(n389) );
  XOR U238 ( .A(n392), .B(n393), .Z(n391) );
  XOR U239 ( .A(n394), .B(n395), .Z(n390) );
  XOR U240 ( .A(n396), .B(n397), .Z(n395) );
  XOR U241 ( .A(n398), .B(n399), .Z(n397) );
  XOR U242 ( .A(n400), .B(n401), .Z(n399) );
  XOR U243 ( .A(n402), .B(n403), .Z(n401) );
  XNOR U244 ( .A(n404), .B(n405), .Z(n400) );
  XNOR U245 ( .A(n406), .B(n407), .Z(n405) );
  NOR U246 ( .A(n408), .B(n403), .Z(n406) );
  XOR U247 ( .A(n409), .B(n410), .Z(n398) );
  XOR U248 ( .A(n411), .B(n412), .Z(n410) );
  XNOR U249 ( .A(n413), .B(n414), .Z(n412) );
  XOR U250 ( .A(n415), .B(n416), .Z(n414) );
  XOR U251 ( .A(n417), .B(n418), .Z(n416) );
  XOR U252 ( .A(n419), .B(n420), .Z(n418) );
  XOR U253 ( .A(n421), .B(n422), .Z(n417) );
  XOR U254 ( .A(n423), .B(n424), .Z(n422) );
  XOR U255 ( .A(n425), .B(n426), .Z(n424) );
  XOR U256 ( .A(n427), .B(n428), .Z(n426) );
  XOR U257 ( .A(n429), .B(n430), .Z(n428) );
  XNOR U258 ( .A(n431), .B(n432), .Z(n427) );
  XNOR U259 ( .A(n433), .B(n434), .Z(n432) );
  NOR U260 ( .A(n435), .B(n430), .Z(n433) );
  XOR U261 ( .A(n436), .B(n437), .Z(n425) );
  XOR U262 ( .A(n438), .B(n439), .Z(n437) );
  XNOR U263 ( .A(n440), .B(n441), .Z(n439) );
  XOR U264 ( .A(n442), .B(n443), .Z(n438) );
  XOR U265 ( .A(n444), .B(n445), .Z(n436) );
  XOR U266 ( .A(n446), .B(n447), .Z(n445) );
  AND U267 ( .A(n448), .B(n449), .Z(n447) );
  XOR U268 ( .A(n441), .B(n450), .Z(n448) );
  XOR U269 ( .A(n451), .B(n452), .Z(n441) );
  AND U270 ( .A(n450), .B(n451), .Z(n452) );
  NOR U271 ( .A(n453), .B(n442), .Z(n446) );
  XOR U272 ( .A(n454), .B(n455), .Z(n444) );
  NOR U273 ( .A(n456), .B(n443), .Z(n455) );
  NOR U274 ( .A(n457), .B(n440), .Z(n454) );
  XOR U275 ( .A(n458), .B(n459), .Z(n423) );
  NOR U276 ( .A(n460), .B(n434), .Z(n459) );
  NOR U277 ( .A(n461), .B(n431), .Z(n458) );
  XOR U278 ( .A(n462), .B(n463), .Z(n421) );
  XOR U279 ( .A(n464), .B(n465), .Z(n463) );
  NOR U280 ( .A(n466), .B(n429), .Z(n465) );
  NOR U281 ( .A(n467), .B(n468), .Z(n464) );
  XOR U282 ( .A(n469), .B(n470), .Z(n462) );
  AND U283 ( .A(n471), .B(n472), .Z(n470) );
  NOR U284 ( .A(n473), .B(n419), .Z(n469) );
  XOR U285 ( .A(n474), .B(n475), .Z(n415) );
  XNOR U286 ( .A(n468), .B(n472), .Z(n475) );
  XOR U287 ( .A(n476), .B(n477), .Z(n474) );
  NOR U288 ( .A(n478), .B(n420), .Z(n477) );
  NOR U289 ( .A(n479), .B(n480), .Z(n476) );
  XOR U290 ( .A(n481), .B(n482), .Z(n411) );
  XOR U291 ( .A(n483), .B(n484), .Z(n409) );
  XNOR U292 ( .A(n485), .B(n480), .Z(n484) );
  NOR U293 ( .A(n486), .B(n481), .Z(n485) );
  XOR U294 ( .A(n487), .B(n488), .Z(n483) );
  NOR U295 ( .A(n489), .B(n482), .Z(n488) );
  NOR U296 ( .A(n490), .B(n413), .Z(n487) );
  XOR U297 ( .A(n491), .B(n492), .Z(n396) );
  NOR U298 ( .A(n493), .B(n407), .Z(n492) );
  NOR U299 ( .A(n494), .B(n404), .Z(n491) );
  XOR U300 ( .A(n495), .B(n496), .Z(n394) );
  XOR U301 ( .A(n497), .B(n498), .Z(n496) );
  NOR U302 ( .A(n499), .B(n402), .Z(n498) );
  NOR U303 ( .A(n500), .B(n501), .Z(n497) );
  XOR U304 ( .A(n502), .B(n503), .Z(n495) );
  AND U305 ( .A(n504), .B(n505), .Z(n503) );
  NOR U306 ( .A(n506), .B(n392), .Z(n502) );
  XOR U307 ( .A(n507), .B(n508), .Z(n388) );
  XNOR U308 ( .A(n501), .B(n505), .Z(n508) );
  XOR U309 ( .A(n509), .B(n510), .Z(n507) );
  NOR U310 ( .A(n511), .B(n393), .Z(n510) );
  NOR U311 ( .A(n512), .B(n513), .Z(n509) );
  XOR U312 ( .A(n514), .B(n515), .Z(n384) );
  XOR U313 ( .A(n516), .B(n517), .Z(n382) );
  XNOR U314 ( .A(n518), .B(n513), .Z(n517) );
  NOR U315 ( .A(n519), .B(n514), .Z(n518) );
  XOR U316 ( .A(n520), .B(n521), .Z(n516) );
  NOR U317 ( .A(n522), .B(n515), .Z(n521) );
  NOR U318 ( .A(n523), .B(n386), .Z(n520) );
  XOR U319 ( .A(n524), .B(n525), .Z(n369) );
  NOR U320 ( .A(n526), .B(n380), .Z(n525) );
  NOR U321 ( .A(n527), .B(n377), .Z(n524) );
  XOR U322 ( .A(n528), .B(n529), .Z(n367) );
  XOR U323 ( .A(n530), .B(n531), .Z(n529) );
  NOR U324 ( .A(n532), .B(n375), .Z(n531) );
  NOR U325 ( .A(n533), .B(n534), .Z(n530) );
  XOR U326 ( .A(n535), .B(n536), .Z(n528) );
  AND U327 ( .A(n537), .B(n538), .Z(n536) );
  NOR U328 ( .A(n539), .B(n365), .Z(n535) );
  XOR U329 ( .A(n540), .B(n541), .Z(n361) );
  XNOR U330 ( .A(n534), .B(n538), .Z(n541) );
  XOR U331 ( .A(n542), .B(n543), .Z(n540) );
  NOR U332 ( .A(n544), .B(n366), .Z(n543) );
  NOR U333 ( .A(n545), .B(n546), .Z(n542) );
  XOR U334 ( .A(n547), .B(n548), .Z(n357) );
  XOR U335 ( .A(n549), .B(n550), .Z(n355) );
  XNOR U336 ( .A(n551), .B(n546), .Z(n550) );
  NOR U337 ( .A(n552), .B(n547), .Z(n551) );
  XOR U338 ( .A(n553), .B(n554), .Z(n549) );
  NOR U339 ( .A(n555), .B(n548), .Z(n554) );
  NOR U340 ( .A(n556), .B(n359), .Z(n553) );
  XOR U341 ( .A(n557), .B(n558), .Z(n342) );
  NOR U342 ( .A(n559), .B(n353), .Z(n558) );
  NOR U343 ( .A(n560), .B(n350), .Z(n557) );
  XOR U344 ( .A(n561), .B(n562), .Z(n340) );
  XOR U345 ( .A(n563), .B(n564), .Z(n562) );
  NOR U346 ( .A(n565), .B(n348), .Z(n564) );
  NOR U347 ( .A(n566), .B(n567), .Z(n563) );
  XOR U348 ( .A(n568), .B(n569), .Z(n561) );
  AND U349 ( .A(n570), .B(n571), .Z(n569) );
  NOR U350 ( .A(n572), .B(n338), .Z(n568) );
  XOR U351 ( .A(n573), .B(n574), .Z(n334) );
  XNOR U352 ( .A(n567), .B(n571), .Z(n574) );
  XOR U353 ( .A(n575), .B(n576), .Z(n573) );
  NOR U354 ( .A(n577), .B(n339), .Z(n576) );
  NOR U355 ( .A(n578), .B(n579), .Z(n575) );
  XOR U356 ( .A(n580), .B(n581), .Z(n330) );
  XOR U357 ( .A(n582), .B(n583), .Z(n328) );
  XNOR U358 ( .A(n584), .B(n579), .Z(n583) );
  NOR U359 ( .A(n585), .B(n580), .Z(n584) );
  XOR U360 ( .A(n586), .B(n587), .Z(n582) );
  NOR U361 ( .A(n588), .B(n581), .Z(n587) );
  NOR U362 ( .A(n589), .B(n332), .Z(n586) );
  XOR U363 ( .A(n590), .B(n591), .Z(n315) );
  NOR U364 ( .A(n592), .B(n326), .Z(n591) );
  NOR U365 ( .A(n593), .B(n323), .Z(n590) );
  XOR U366 ( .A(n594), .B(n595), .Z(n313) );
  XOR U367 ( .A(n596), .B(n597), .Z(n595) );
  NOR U368 ( .A(n598), .B(n321), .Z(n597) );
  NOR U369 ( .A(n599), .B(n600), .Z(n596) );
  XOR U370 ( .A(n601), .B(n602), .Z(n594) );
  AND U371 ( .A(n603), .B(n604), .Z(n602) );
  NOR U372 ( .A(n605), .B(n311), .Z(n601) );
  XOR U373 ( .A(n606), .B(n607), .Z(n307) );
  XNOR U374 ( .A(n600), .B(n604), .Z(n607) );
  XOR U375 ( .A(n608), .B(n609), .Z(n606) );
  NOR U376 ( .A(n610), .B(n312), .Z(n609) );
  NOR U377 ( .A(n611), .B(n612), .Z(n608) );
  XOR U378 ( .A(n613), .B(n614), .Z(n303) );
  XOR U379 ( .A(n615), .B(n616), .Z(n301) );
  XNOR U380 ( .A(n617), .B(n612), .Z(n616) );
  NOR U381 ( .A(n618), .B(n613), .Z(n617) );
  XOR U382 ( .A(n619), .B(n620), .Z(n615) );
  NOR U383 ( .A(n621), .B(n614), .Z(n620) );
  NOR U384 ( .A(n622), .B(n305), .Z(n619) );
  XOR U385 ( .A(n623), .B(n624), .Z(n288) );
  NOR U386 ( .A(n625), .B(n299), .Z(n624) );
  NOR U387 ( .A(n626), .B(n296), .Z(n623) );
  XOR U388 ( .A(n627), .B(n628), .Z(n286) );
  XOR U389 ( .A(n629), .B(n630), .Z(n628) );
  NOR U390 ( .A(n631), .B(n294), .Z(n630) );
  NOR U391 ( .A(n632), .B(n633), .Z(n629) );
  XOR U392 ( .A(n634), .B(n635), .Z(n627) );
  AND U393 ( .A(n636), .B(n637), .Z(n635) );
  NOR U394 ( .A(n638), .B(n284), .Z(n634) );
  XOR U395 ( .A(n639), .B(n640), .Z(n280) );
  XNOR U396 ( .A(n633), .B(n637), .Z(n640) );
  XOR U397 ( .A(n641), .B(n642), .Z(n639) );
  NOR U398 ( .A(n643), .B(n285), .Z(n642) );
  NOR U399 ( .A(n644), .B(n645), .Z(n641) );
  XOR U400 ( .A(n646), .B(n647), .Z(n276) );
  XOR U401 ( .A(n648), .B(n649), .Z(n274) );
  XNOR U402 ( .A(n650), .B(n645), .Z(n649) );
  NOR U403 ( .A(n651), .B(n646), .Z(n650) );
  XOR U404 ( .A(n652), .B(n653), .Z(n648) );
  NOR U405 ( .A(n654), .B(n647), .Z(n653) );
  NOR U406 ( .A(n655), .B(n278), .Z(n652) );
  XOR U407 ( .A(n656), .B(n657), .Z(n261) );
  NOR U408 ( .A(n658), .B(n272), .Z(n657) );
  NOR U409 ( .A(n659), .B(n269), .Z(n656) );
  XOR U410 ( .A(n660), .B(n661), .Z(n259) );
  XOR U411 ( .A(n662), .B(n663), .Z(n661) );
  NOR U412 ( .A(n664), .B(n267), .Z(n663) );
  NOR U413 ( .A(n665), .B(n666), .Z(n662) );
  XOR U414 ( .A(n667), .B(n668), .Z(n660) );
  AND U415 ( .A(n669), .B(n670), .Z(n668) );
  NOR U416 ( .A(n671), .B(n257), .Z(n667) );
  XOR U417 ( .A(n672), .B(n673), .Z(n253) );
  XNOR U418 ( .A(n666), .B(n670), .Z(n673) );
  XOR U419 ( .A(n674), .B(n675), .Z(n672) );
  NOR U420 ( .A(n676), .B(n258), .Z(n675) );
  NOR U421 ( .A(n677), .B(n678), .Z(n674) );
  XOR U422 ( .A(n679), .B(n680), .Z(n249) );
  XOR U423 ( .A(n681), .B(n682), .Z(n247) );
  XNOR U424 ( .A(n683), .B(n678), .Z(n682) );
  NOR U425 ( .A(n684), .B(n679), .Z(n683) );
  XOR U426 ( .A(n685), .B(n686), .Z(n681) );
  NOR U427 ( .A(n687), .B(n680), .Z(n686) );
  NOR U428 ( .A(n688), .B(n251), .Z(n685) );
  XOR U429 ( .A(n689), .B(n690), .Z(n234) );
  NOR U430 ( .A(n691), .B(n245), .Z(n690) );
  NOR U431 ( .A(n692), .B(n242), .Z(n689) );
  XOR U432 ( .A(n693), .B(n694), .Z(n232) );
  XOR U433 ( .A(n695), .B(n696), .Z(n694) );
  NOR U434 ( .A(n697), .B(n240), .Z(n696) );
  NOR U435 ( .A(n698), .B(n699), .Z(n695) );
  XOR U436 ( .A(n700), .B(n701), .Z(n693) );
  AND U437 ( .A(n702), .B(n703), .Z(n701) );
  NOR U438 ( .A(n704), .B(n230), .Z(n700) );
  XOR U439 ( .A(n705), .B(n706), .Z(n226) );
  XNOR U440 ( .A(n699), .B(n703), .Z(n706) );
  XOR U441 ( .A(n707), .B(n708), .Z(n705) );
  NOR U442 ( .A(n709), .B(n231), .Z(n708) );
  NOR U443 ( .A(n710), .B(n711), .Z(n707) );
  XOR U444 ( .A(n712), .B(n713), .Z(n222) );
  XOR U445 ( .A(n714), .B(n715), .Z(n220) );
  XNOR U446 ( .A(n716), .B(n711), .Z(n715) );
  NOR U447 ( .A(n717), .B(n712), .Z(n716) );
  XOR U448 ( .A(n718), .B(n719), .Z(n714) );
  NOR U449 ( .A(n720), .B(n713), .Z(n719) );
  NOR U450 ( .A(n721), .B(n224), .Z(n718) );
  XOR U451 ( .A(n722), .B(n723), .Z(n207) );
  NOR U452 ( .A(n724), .B(n218), .Z(n723) );
  NOR U453 ( .A(n725), .B(n215), .Z(n722) );
  XOR U454 ( .A(n726), .B(n727), .Z(n205) );
  XOR U455 ( .A(n728), .B(n729), .Z(n727) );
  NOR U456 ( .A(n730), .B(n213), .Z(n729) );
  NOR U457 ( .A(n731), .B(n732), .Z(n728) );
  XOR U458 ( .A(n733), .B(n734), .Z(n726) );
  AND U459 ( .A(n735), .B(n736), .Z(n734) );
  NOR U460 ( .A(n737), .B(n203), .Z(n733) );
  XOR U461 ( .A(n738), .B(n739), .Z(n199) );
  XNOR U462 ( .A(n732), .B(n736), .Z(n739) );
  XOR U463 ( .A(n740), .B(n741), .Z(n738) );
  NOR U464 ( .A(n742), .B(n204), .Z(n741) );
  NOR U465 ( .A(n743), .B(n744), .Z(n740) );
  XOR U466 ( .A(n745), .B(n746), .Z(n195) );
  XOR U467 ( .A(n747), .B(n748), .Z(n193) );
  XNOR U468 ( .A(n749), .B(n744), .Z(n748) );
  NOR U469 ( .A(n750), .B(n745), .Z(n749) );
  XOR U470 ( .A(n751), .B(n752), .Z(n747) );
  NOR U471 ( .A(n753), .B(n746), .Z(n752) );
  NOR U472 ( .A(n754), .B(n197), .Z(n751) );
  XOR U473 ( .A(n755), .B(n756), .Z(n180) );
  NOR U474 ( .A(n757), .B(n191), .Z(n756) );
  NOR U475 ( .A(n758), .B(n188), .Z(n755) );
  XOR U476 ( .A(n759), .B(n760), .Z(n178) );
  XOR U477 ( .A(n761), .B(n762), .Z(n760) );
  NOR U478 ( .A(n763), .B(n186), .Z(n762) );
  NOR U479 ( .A(n764), .B(n765), .Z(n761) );
  XOR U480 ( .A(n766), .B(n767), .Z(n759) );
  AND U481 ( .A(n768), .B(n769), .Z(n767) );
  NOR U482 ( .A(n770), .B(n176), .Z(n766) );
  XOR U483 ( .A(n771), .B(n772), .Z(n172) );
  XNOR U484 ( .A(n765), .B(n769), .Z(n772) );
  XOR U485 ( .A(n773), .B(n774), .Z(n771) );
  NOR U486 ( .A(n775), .B(n177), .Z(n774) );
  NOR U487 ( .A(n776), .B(n777), .Z(n773) );
  XOR U488 ( .A(n778), .B(n779), .Z(n168) );
  XOR U489 ( .A(n780), .B(n781), .Z(n166) );
  XNOR U490 ( .A(n782), .B(n777), .Z(n781) );
  NOR U491 ( .A(n783), .B(n778), .Z(n782) );
  XOR U492 ( .A(n784), .B(n785), .Z(n780) );
  NOR U493 ( .A(n786), .B(n779), .Z(n785) );
  NOR U494 ( .A(n787), .B(n170), .Z(n784) );
  XOR U495 ( .A(n788), .B(n789), .Z(n164) );
  XNOR U496 ( .A(n159), .B(n790), .Z(n789) );
  XNOR U497 ( .A(n791), .B(n163), .Z(n790) );
  AND U498 ( .A(n792), .B(n793), .Z(n791) );
  XOR U499 ( .A(n793), .B(n161), .Z(n788) );
  XNOR U500 ( .A(n794), .B(n795), .Z(n138) );
  NOR U501 ( .A(n44), .B(n794), .Z(n795) );
  XNOR U502 ( .A(n144), .B(n148), .Z(n150) );
  XOR U503 ( .A(n145), .B(n143), .Z(n144) );
  XNOR U504 ( .A(n796), .B(n797), .Z(n143) );
  XOR U505 ( .A(n798), .B(n799), .Z(n797) );
  XNOR U506 ( .A(n800), .B(n801), .Z(n799) );
  NOR U507 ( .A(n802), .B(n801), .Z(n800) );
  XOR U508 ( .A(n803), .B(n804), .Z(n798) );
  NOR U509 ( .A(n805), .B(n806), .Z(n804) );
  AND U510 ( .A(n807), .B(n808), .Z(n803) );
  XOR U511 ( .A(n809), .B(n810), .Z(n796) );
  XOR U512 ( .A(n811), .B(n812), .Z(n810) );
  XOR U513 ( .A(n813), .B(n814), .Z(n812) );
  XOR U514 ( .A(n815), .B(n816), .Z(n814) );
  XNOR U515 ( .A(n817), .B(n818), .Z(n816) );
  NOR U516 ( .A(n819), .B(n818), .Z(n817) );
  XOR U517 ( .A(n820), .B(n821), .Z(n815) );
  XOR U518 ( .A(n822), .B(n823), .Z(n821) );
  XOR U519 ( .A(n824), .B(n825), .Z(n823) );
  XNOR U520 ( .A(n826), .B(n827), .Z(n825) );
  NOR U521 ( .A(n828), .B(n827), .Z(n826) );
  XOR U522 ( .A(n829), .B(n830), .Z(n824) );
  XOR U523 ( .A(n831), .B(n832), .Z(n830) );
  XOR U524 ( .A(n833), .B(n834), .Z(n832) );
  XNOR U525 ( .A(n835), .B(n836), .Z(n834) );
  NOR U526 ( .A(n837), .B(n836), .Z(n835) );
  XOR U527 ( .A(n838), .B(n839), .Z(n833) );
  XOR U528 ( .A(n840), .B(n841), .Z(n839) );
  XOR U529 ( .A(n842), .B(n843), .Z(n841) );
  XNOR U530 ( .A(n844), .B(n845), .Z(n843) );
  NOR U531 ( .A(n846), .B(n845), .Z(n844) );
  XOR U532 ( .A(n847), .B(n848), .Z(n842) );
  XOR U533 ( .A(n849), .B(n850), .Z(n848) );
  XOR U534 ( .A(n851), .B(n852), .Z(n850) );
  XNOR U535 ( .A(n853), .B(n854), .Z(n852) );
  NOR U536 ( .A(n855), .B(n854), .Z(n853) );
  XOR U537 ( .A(n856), .B(n857), .Z(n851) );
  XOR U538 ( .A(n858), .B(n859), .Z(n857) );
  XOR U539 ( .A(n860), .B(n861), .Z(n859) );
  XNOR U540 ( .A(n862), .B(n863), .Z(n861) );
  NOR U541 ( .A(n864), .B(n863), .Z(n862) );
  XOR U542 ( .A(n865), .B(n866), .Z(n860) );
  XOR U543 ( .A(n867), .B(n868), .Z(n866) );
  XOR U544 ( .A(n869), .B(n870), .Z(n868) );
  XNOR U545 ( .A(n871), .B(n872), .Z(n870) );
  NOR U546 ( .A(n873), .B(n872), .Z(n871) );
  XOR U547 ( .A(n874), .B(n875), .Z(n869) );
  XOR U548 ( .A(n876), .B(n877), .Z(n875) );
  XOR U549 ( .A(n878), .B(n879), .Z(n877) );
  XNOR U550 ( .A(n880), .B(n881), .Z(n879) );
  NOR U551 ( .A(n882), .B(n881), .Z(n880) );
  XOR U552 ( .A(n883), .B(n884), .Z(n878) );
  XOR U553 ( .A(n885), .B(n886), .Z(n884) );
  XOR U554 ( .A(n887), .B(n888), .Z(n886) );
  XNOR U555 ( .A(n889), .B(n890), .Z(n888) );
  NOR U556 ( .A(n891), .B(n890), .Z(n889) );
  XOR U557 ( .A(n892), .B(n893), .Z(n887) );
  XOR U558 ( .A(n894), .B(n895), .Z(n893) );
  XOR U559 ( .A(n896), .B(n897), .Z(n895) );
  XNOR U560 ( .A(n898), .B(n899), .Z(n897) );
  NOR U561 ( .A(n900), .B(n899), .Z(n898) );
  XOR U562 ( .A(n901), .B(n902), .Z(n896) );
  XOR U563 ( .A(n903), .B(n904), .Z(n902) );
  XOR U564 ( .A(n905), .B(n906), .Z(n904) );
  XNOR U565 ( .A(n907), .B(n908), .Z(n906) );
  NOR U566 ( .A(n909), .B(n908), .Z(n907) );
  XOR U567 ( .A(n910), .B(n911), .Z(n905) );
  XOR U568 ( .A(n912), .B(n913), .Z(n911) );
  XOR U569 ( .A(n914), .B(n915), .Z(n913) );
  XNOR U570 ( .A(n916), .B(n917), .Z(n915) );
  NOR U571 ( .A(n918), .B(n917), .Z(n916) );
  XOR U572 ( .A(n919), .B(n920), .Z(n914) );
  XOR U573 ( .A(n921), .B(n922), .Z(n920) );
  XOR U574 ( .A(n923), .B(n924), .Z(n922) );
  XNOR U575 ( .A(n925), .B(n926), .Z(n924) );
  NOR U576 ( .A(n927), .B(n926), .Z(n925) );
  XOR U577 ( .A(n928), .B(n929), .Z(n923) );
  XOR U578 ( .A(n930), .B(n931), .Z(n929) );
  XOR U579 ( .A(n932), .B(n933), .Z(n931) );
  XNOR U580 ( .A(n934), .B(n935), .Z(n933) );
  NOR U581 ( .A(n936), .B(n935), .Z(n934) );
  XOR U582 ( .A(n937), .B(n938), .Z(n932) );
  XOR U583 ( .A(n939), .B(n940), .Z(n938) );
  XOR U584 ( .A(n941), .B(n942), .Z(n940) );
  XNOR U585 ( .A(n943), .B(n944), .Z(n942) );
  NOR U586 ( .A(n945), .B(n944), .Z(n943) );
  XOR U587 ( .A(n946), .B(n947), .Z(n941) );
  XOR U588 ( .A(n948), .B(n949), .Z(n947) );
  XOR U589 ( .A(n950), .B(n951), .Z(n949) );
  XNOR U590 ( .A(n952), .B(n953), .Z(n951) );
  NOR U591 ( .A(n954), .B(n953), .Z(n952) );
  XOR U592 ( .A(n955), .B(n956), .Z(n950) );
  XOR U593 ( .A(n957), .B(n958), .Z(n956) );
  XOR U594 ( .A(n959), .B(n960), .Z(n958) );
  XNOR U595 ( .A(n961), .B(n962), .Z(n960) );
  NOR U596 ( .A(n963), .B(n962), .Z(n961) );
  XOR U597 ( .A(n964), .B(n965), .Z(n959) );
  XOR U598 ( .A(n966), .B(n967), .Z(n965) );
  XOR U599 ( .A(n968), .B(n969), .Z(n967) );
  XNOR U600 ( .A(n970), .B(n971), .Z(n969) );
  NOR U601 ( .A(n972), .B(n971), .Z(n970) );
  XOR U602 ( .A(n973), .B(n974), .Z(n968) );
  XOR U603 ( .A(n975), .B(n976), .Z(n974) );
  XOR U604 ( .A(n977), .B(n978), .Z(n976) );
  XNOR U605 ( .A(n979), .B(n980), .Z(n978) );
  NOR U606 ( .A(n981), .B(n980), .Z(n979) );
  XOR U607 ( .A(n982), .B(n983), .Z(n977) );
  XOR U608 ( .A(n984), .B(n985), .Z(n983) );
  XOR U609 ( .A(n986), .B(n987), .Z(n985) );
  XNOR U610 ( .A(n988), .B(n989), .Z(n987) );
  NOR U611 ( .A(n990), .B(n989), .Z(n988) );
  XOR U612 ( .A(n991), .B(n992), .Z(n986) );
  XOR U613 ( .A(n993), .B(n994), .Z(n992) );
  XOR U614 ( .A(n995), .B(n996), .Z(n994) );
  XNOR U615 ( .A(n997), .B(n998), .Z(n996) );
  NOR U616 ( .A(n999), .B(n998), .Z(n997) );
  XOR U617 ( .A(n1000), .B(n1001), .Z(n995) );
  XOR U618 ( .A(n1002), .B(n1003), .Z(n1001) );
  XOR U619 ( .A(n1004), .B(n1005), .Z(n1003) );
  XNOR U620 ( .A(n1006), .B(n1007), .Z(n1005) );
  NOR U621 ( .A(n1008), .B(n1007), .Z(n1006) );
  XOR U622 ( .A(n1009), .B(n1010), .Z(n1004) );
  XOR U623 ( .A(n1011), .B(n1012), .Z(n1010) );
  XOR U624 ( .A(n1013), .B(n1014), .Z(n1012) );
  XNOR U625 ( .A(n1015), .B(n1016), .Z(n1014) );
  NOR U626 ( .A(n1017), .B(n1016), .Z(n1015) );
  XOR U627 ( .A(n1018), .B(n1019), .Z(n1013) );
  XOR U628 ( .A(n1020), .B(n1021), .Z(n1019) );
  XOR U629 ( .A(n1022), .B(n1023), .Z(n1021) );
  XNOR U630 ( .A(n1024), .B(n1025), .Z(n1023) );
  NOR U631 ( .A(n1026), .B(n1025), .Z(n1024) );
  XOR U632 ( .A(n1027), .B(n1028), .Z(n1022) );
  XOR U633 ( .A(n1029), .B(n1030), .Z(n1028) );
  XOR U634 ( .A(n1031), .B(n1032), .Z(n1030) );
  XNOR U635 ( .A(n1033), .B(n1034), .Z(n1032) );
  NOR U636 ( .A(n1035), .B(n1034), .Z(n1033) );
  XOR U637 ( .A(n1036), .B(n1037), .Z(n1031) );
  XOR U638 ( .A(n1038), .B(n1039), .Z(n1037) );
  XOR U639 ( .A(n1040), .B(n1041), .Z(n1039) );
  XNOR U640 ( .A(n1042), .B(n1043), .Z(n1041) );
  NOR U641 ( .A(n1044), .B(n1043), .Z(n1042) );
  XOR U642 ( .A(n1045), .B(n1046), .Z(n1040) );
  XOR U643 ( .A(n1047), .B(n1048), .Z(n1046) );
  XOR U644 ( .A(n1049), .B(n1050), .Z(n1048) );
  XNOR U645 ( .A(n1051), .B(n1052), .Z(n1050) );
  NOR U646 ( .A(n1053), .B(n1052), .Z(n1051) );
  XOR U647 ( .A(n1054), .B(n1055), .Z(n1049) );
  XOR U648 ( .A(n1056), .B(n1057), .Z(n1055) );
  XOR U649 ( .A(n1058), .B(n1059), .Z(n1057) );
  XNOR U650 ( .A(n1060), .B(n1061), .Z(n1059) );
  NOR U651 ( .A(n1062), .B(n1061), .Z(n1060) );
  XOR U652 ( .A(n1063), .B(n1064), .Z(n1058) );
  XOR U653 ( .A(n1065), .B(n1066), .Z(n1064) );
  XOR U654 ( .A(n1067), .B(n1068), .Z(n1066) );
  XNOR U655 ( .A(n1069), .B(n1070), .Z(n1068) );
  NOR U656 ( .A(n1071), .B(n1070), .Z(n1069) );
  XOR U657 ( .A(n1072), .B(n1073), .Z(n1067) );
  XOR U658 ( .A(n1074), .B(n1075), .Z(n1073) );
  XOR U659 ( .A(n1076), .B(n1077), .Z(n1075) );
  XOR U660 ( .A(n1078), .B(n1079), .Z(n1074) );
  XNOR U661 ( .A(n1080), .B(n1081), .Z(n1079) );
  XOR U662 ( .A(n1082), .B(n1083), .Z(n1081) );
  XOR U663 ( .A(n1084), .B(n1085), .Z(n1083) );
  XNOR U664 ( .A(n1086), .B(n1087), .Z(n1085) );
  XOR U665 ( .A(n1088), .B(n1089), .Z(n1084) );
  XOR U666 ( .A(n1090), .B(n1091), .Z(n1082) );
  XOR U667 ( .A(n1092), .B(n1093), .Z(n1091) );
  AND U668 ( .A(n1094), .B(n1095), .Z(n1093) );
  XOR U669 ( .A(n1087), .B(n1096), .Z(n1094) );
  XOR U670 ( .A(n1097), .B(n1098), .Z(n1087) );
  AND U671 ( .A(n1096), .B(n1097), .Z(n1098) );
  NOR U672 ( .A(n1099), .B(n1088), .Z(n1092) );
  XOR U673 ( .A(n1100), .B(n1101), .Z(n1090) );
  NOR U674 ( .A(n1102), .B(n1089), .Z(n1101) );
  NOR U675 ( .A(n1103), .B(n1086), .Z(n1100) );
  XNOR U676 ( .A(n1104), .B(n1105), .Z(n1078) );
  XNOR U677 ( .A(n1106), .B(n1107), .Z(n1105) );
  NOR U678 ( .A(n1108), .B(n1080), .Z(n1106) );
  XOR U679 ( .A(n1109), .B(n1110), .Z(n1072) );
  XOR U680 ( .A(n1111), .B(n1112), .Z(n1110) );
  NOR U681 ( .A(n1113), .B(n1076), .Z(n1112) );
  NOR U682 ( .A(n1114), .B(n1107), .Z(n1111) );
  XOR U683 ( .A(n1115), .B(n1116), .Z(n1109) );
  NOR U684 ( .A(n1117), .B(n1104), .Z(n1116) );
  NOR U685 ( .A(n1118), .B(n1077), .Z(n1115) );
  XOR U686 ( .A(n1119), .B(n1120), .Z(n1065) );
  XOR U687 ( .A(n1121), .B(n1122), .Z(n1063) );
  XNOR U688 ( .A(n1123), .B(n1124), .Z(n1122) );
  NOR U689 ( .A(n1125), .B(n1124), .Z(n1123) );
  XOR U690 ( .A(n1126), .B(n1127), .Z(n1121) );
  NOR U691 ( .A(n1128), .B(n1119), .Z(n1127) );
  NOR U692 ( .A(n1129), .B(n1120), .Z(n1126) );
  XOR U693 ( .A(n1130), .B(n1131), .Z(n1056) );
  XOR U694 ( .A(n1132), .B(n1133), .Z(n1054) );
  XNOR U695 ( .A(n1134), .B(n1135), .Z(n1133) );
  NOR U696 ( .A(n1136), .B(n1135), .Z(n1134) );
  XOR U697 ( .A(n1137), .B(n1138), .Z(n1132) );
  NOR U698 ( .A(n1139), .B(n1130), .Z(n1138) );
  NOR U699 ( .A(n1140), .B(n1131), .Z(n1137) );
  XOR U700 ( .A(n1141), .B(n1142), .Z(n1047) );
  XOR U701 ( .A(n1143), .B(n1144), .Z(n1045) );
  XNOR U702 ( .A(n1145), .B(n1146), .Z(n1144) );
  NOR U703 ( .A(n1147), .B(n1146), .Z(n1145) );
  XOR U704 ( .A(n1148), .B(n1149), .Z(n1143) );
  NOR U705 ( .A(n1150), .B(n1141), .Z(n1149) );
  NOR U706 ( .A(n1151), .B(n1142), .Z(n1148) );
  XOR U707 ( .A(n1152), .B(n1153), .Z(n1038) );
  XOR U708 ( .A(n1154), .B(n1155), .Z(n1036) );
  XNOR U709 ( .A(n1156), .B(n1157), .Z(n1155) );
  NOR U710 ( .A(n1158), .B(n1157), .Z(n1156) );
  XOR U711 ( .A(n1159), .B(n1160), .Z(n1154) );
  NOR U712 ( .A(n1161), .B(n1152), .Z(n1160) );
  NOR U713 ( .A(n1162), .B(n1153), .Z(n1159) );
  XOR U714 ( .A(n1163), .B(n1164), .Z(n1029) );
  XOR U715 ( .A(n1165), .B(n1166), .Z(n1027) );
  XNOR U716 ( .A(n1167), .B(n1168), .Z(n1166) );
  NOR U717 ( .A(n1169), .B(n1168), .Z(n1167) );
  XOR U718 ( .A(n1170), .B(n1171), .Z(n1165) );
  NOR U719 ( .A(n1172), .B(n1163), .Z(n1171) );
  NOR U720 ( .A(n1173), .B(n1164), .Z(n1170) );
  XOR U721 ( .A(n1174), .B(n1175), .Z(n1020) );
  XOR U722 ( .A(n1176), .B(n1177), .Z(n1018) );
  XNOR U723 ( .A(n1178), .B(n1179), .Z(n1177) );
  NOR U724 ( .A(n1180), .B(n1179), .Z(n1178) );
  XOR U725 ( .A(n1181), .B(n1182), .Z(n1176) );
  NOR U726 ( .A(n1183), .B(n1174), .Z(n1182) );
  NOR U727 ( .A(n1184), .B(n1175), .Z(n1181) );
  XOR U728 ( .A(n1185), .B(n1186), .Z(n1011) );
  XOR U729 ( .A(n1187), .B(n1188), .Z(n1009) );
  XNOR U730 ( .A(n1189), .B(n1190), .Z(n1188) );
  NOR U731 ( .A(n1191), .B(n1190), .Z(n1189) );
  XOR U732 ( .A(n1192), .B(n1193), .Z(n1187) );
  NOR U733 ( .A(n1194), .B(n1185), .Z(n1193) );
  NOR U734 ( .A(n1195), .B(n1186), .Z(n1192) );
  XOR U735 ( .A(n1196), .B(n1197), .Z(n1002) );
  XOR U736 ( .A(n1198), .B(n1199), .Z(n1000) );
  XNOR U737 ( .A(n1200), .B(n1201), .Z(n1199) );
  NOR U738 ( .A(n1202), .B(n1201), .Z(n1200) );
  XOR U739 ( .A(n1203), .B(n1204), .Z(n1198) );
  NOR U740 ( .A(n1205), .B(n1196), .Z(n1204) );
  NOR U741 ( .A(n1206), .B(n1197), .Z(n1203) );
  XOR U742 ( .A(n1207), .B(n1208), .Z(n993) );
  XOR U743 ( .A(n1209), .B(n1210), .Z(n991) );
  XNOR U744 ( .A(n1211), .B(n1212), .Z(n1210) );
  NOR U745 ( .A(n1213), .B(n1212), .Z(n1211) );
  XOR U746 ( .A(n1214), .B(n1215), .Z(n1209) );
  NOR U747 ( .A(n1216), .B(n1207), .Z(n1215) );
  NOR U748 ( .A(n1217), .B(n1208), .Z(n1214) );
  XOR U749 ( .A(n1218), .B(n1219), .Z(n984) );
  XOR U750 ( .A(n1220), .B(n1221), .Z(n982) );
  XNOR U751 ( .A(n1222), .B(n1223), .Z(n1221) );
  NOR U752 ( .A(n1224), .B(n1223), .Z(n1222) );
  XOR U753 ( .A(n1225), .B(n1226), .Z(n1220) );
  NOR U754 ( .A(n1227), .B(n1218), .Z(n1226) );
  NOR U755 ( .A(n1228), .B(n1219), .Z(n1225) );
  XOR U756 ( .A(n1229), .B(n1230), .Z(n975) );
  XOR U757 ( .A(n1231), .B(n1232), .Z(n973) );
  XNOR U758 ( .A(n1233), .B(n1234), .Z(n1232) );
  NOR U759 ( .A(n1235), .B(n1234), .Z(n1233) );
  XOR U760 ( .A(n1236), .B(n1237), .Z(n1231) );
  NOR U761 ( .A(n1238), .B(n1229), .Z(n1237) );
  NOR U762 ( .A(n1239), .B(n1230), .Z(n1236) );
  XOR U763 ( .A(n1240), .B(n1241), .Z(n966) );
  XOR U764 ( .A(n1242), .B(n1243), .Z(n964) );
  XNOR U765 ( .A(n1244), .B(n1245), .Z(n1243) );
  NOR U766 ( .A(n1246), .B(n1245), .Z(n1244) );
  XOR U767 ( .A(n1247), .B(n1248), .Z(n1242) );
  NOR U768 ( .A(n1249), .B(n1240), .Z(n1248) );
  NOR U769 ( .A(n1250), .B(n1241), .Z(n1247) );
  XOR U770 ( .A(n1251), .B(n1252), .Z(n957) );
  XOR U771 ( .A(n1253), .B(n1254), .Z(n955) );
  XNOR U772 ( .A(n1255), .B(n1256), .Z(n1254) );
  NOR U773 ( .A(n1257), .B(n1256), .Z(n1255) );
  XOR U774 ( .A(n1258), .B(n1259), .Z(n1253) );
  NOR U775 ( .A(n1260), .B(n1251), .Z(n1259) );
  NOR U776 ( .A(n1261), .B(n1252), .Z(n1258) );
  XOR U777 ( .A(n1262), .B(n1263), .Z(n948) );
  XOR U778 ( .A(n1264), .B(n1265), .Z(n946) );
  XNOR U779 ( .A(n1266), .B(n1267), .Z(n1265) );
  NOR U780 ( .A(n1268), .B(n1267), .Z(n1266) );
  XOR U781 ( .A(n1269), .B(n1270), .Z(n1264) );
  NOR U782 ( .A(n1271), .B(n1262), .Z(n1270) );
  NOR U783 ( .A(n1272), .B(n1263), .Z(n1269) );
  XOR U784 ( .A(n1273), .B(n1274), .Z(n939) );
  XOR U785 ( .A(n1275), .B(n1276), .Z(n937) );
  XNOR U786 ( .A(n1277), .B(n1278), .Z(n1276) );
  NOR U787 ( .A(n1279), .B(n1278), .Z(n1277) );
  XOR U788 ( .A(n1280), .B(n1281), .Z(n1275) );
  NOR U789 ( .A(n1282), .B(n1273), .Z(n1281) );
  NOR U790 ( .A(n1283), .B(n1274), .Z(n1280) );
  XOR U791 ( .A(n1284), .B(n1285), .Z(n930) );
  XOR U792 ( .A(n1286), .B(n1287), .Z(n928) );
  XNOR U793 ( .A(n1288), .B(n1289), .Z(n1287) );
  NOR U794 ( .A(n1290), .B(n1289), .Z(n1288) );
  XOR U795 ( .A(n1291), .B(n1292), .Z(n1286) );
  NOR U796 ( .A(n1293), .B(n1284), .Z(n1292) );
  NOR U797 ( .A(n1294), .B(n1285), .Z(n1291) );
  XOR U798 ( .A(n1295), .B(n1296), .Z(n921) );
  XOR U799 ( .A(n1297), .B(n1298), .Z(n919) );
  XNOR U800 ( .A(n1299), .B(n1300), .Z(n1298) );
  NOR U801 ( .A(n1301), .B(n1300), .Z(n1299) );
  XOR U802 ( .A(n1302), .B(n1303), .Z(n1297) );
  NOR U803 ( .A(n1304), .B(n1295), .Z(n1303) );
  NOR U804 ( .A(n1305), .B(n1296), .Z(n1302) );
  XOR U805 ( .A(n1306), .B(n1307), .Z(n912) );
  XOR U806 ( .A(n1308), .B(n1309), .Z(n910) );
  XNOR U807 ( .A(n1310), .B(n1311), .Z(n1309) );
  NOR U808 ( .A(n1312), .B(n1311), .Z(n1310) );
  XOR U809 ( .A(n1313), .B(n1314), .Z(n1308) );
  NOR U810 ( .A(n1315), .B(n1306), .Z(n1314) );
  NOR U811 ( .A(n1316), .B(n1307), .Z(n1313) );
  XOR U812 ( .A(n1317), .B(n1318), .Z(n903) );
  XOR U813 ( .A(n1319), .B(n1320), .Z(n901) );
  XNOR U814 ( .A(n1321), .B(n1322), .Z(n1320) );
  NOR U815 ( .A(n1323), .B(n1322), .Z(n1321) );
  XOR U816 ( .A(n1324), .B(n1325), .Z(n1319) );
  NOR U817 ( .A(n1326), .B(n1317), .Z(n1325) );
  NOR U818 ( .A(n1327), .B(n1318), .Z(n1324) );
  XOR U819 ( .A(n1328), .B(n1329), .Z(n894) );
  XOR U820 ( .A(n1330), .B(n1331), .Z(n892) );
  XNOR U821 ( .A(n1332), .B(n1333), .Z(n1331) );
  NOR U822 ( .A(n1334), .B(n1333), .Z(n1332) );
  XOR U823 ( .A(n1335), .B(n1336), .Z(n1330) );
  NOR U824 ( .A(n1337), .B(n1328), .Z(n1336) );
  NOR U825 ( .A(n1338), .B(n1329), .Z(n1335) );
  XOR U826 ( .A(n1339), .B(n1340), .Z(n885) );
  XOR U827 ( .A(n1341), .B(n1342), .Z(n883) );
  XNOR U828 ( .A(n1343), .B(n1344), .Z(n1342) );
  NOR U829 ( .A(n1345), .B(n1344), .Z(n1343) );
  XOR U830 ( .A(n1346), .B(n1347), .Z(n1341) );
  NOR U831 ( .A(n1348), .B(n1339), .Z(n1347) );
  NOR U832 ( .A(n1349), .B(n1340), .Z(n1346) );
  XOR U833 ( .A(n1350), .B(n1351), .Z(n876) );
  XOR U834 ( .A(n1352), .B(n1353), .Z(n874) );
  XNOR U835 ( .A(n1354), .B(n1355), .Z(n1353) );
  NOR U836 ( .A(n1356), .B(n1355), .Z(n1354) );
  XOR U837 ( .A(n1357), .B(n1358), .Z(n1352) );
  NOR U838 ( .A(n1359), .B(n1350), .Z(n1358) );
  NOR U839 ( .A(n1360), .B(n1351), .Z(n1357) );
  XOR U840 ( .A(n1361), .B(n1362), .Z(n867) );
  XOR U841 ( .A(n1363), .B(n1364), .Z(n865) );
  XNOR U842 ( .A(n1365), .B(n1366), .Z(n1364) );
  NOR U843 ( .A(n1367), .B(n1366), .Z(n1365) );
  XOR U844 ( .A(n1368), .B(n1369), .Z(n1363) );
  NOR U845 ( .A(n1370), .B(n1361), .Z(n1369) );
  NOR U846 ( .A(n1371), .B(n1362), .Z(n1368) );
  XOR U847 ( .A(n1372), .B(n1373), .Z(n858) );
  XOR U848 ( .A(n1374), .B(n1375), .Z(n856) );
  XNOR U849 ( .A(n1376), .B(n1377), .Z(n1375) );
  NOR U850 ( .A(n1378), .B(n1377), .Z(n1376) );
  XOR U851 ( .A(n1379), .B(n1380), .Z(n1374) );
  NOR U852 ( .A(n1381), .B(n1372), .Z(n1380) );
  NOR U853 ( .A(n1382), .B(n1373), .Z(n1379) );
  XOR U854 ( .A(n1383), .B(n1384), .Z(n849) );
  XOR U855 ( .A(n1385), .B(n1386), .Z(n847) );
  XNOR U856 ( .A(n1387), .B(n1388), .Z(n1386) );
  NOR U857 ( .A(n1389), .B(n1388), .Z(n1387) );
  XOR U858 ( .A(n1390), .B(n1391), .Z(n1385) );
  NOR U859 ( .A(n1392), .B(n1383), .Z(n1391) );
  NOR U860 ( .A(n1393), .B(n1384), .Z(n1390) );
  XOR U861 ( .A(n1394), .B(n1395), .Z(n840) );
  XOR U862 ( .A(n1396), .B(n1397), .Z(n838) );
  XNOR U863 ( .A(n1398), .B(n1399), .Z(n1397) );
  NOR U864 ( .A(n1400), .B(n1399), .Z(n1398) );
  XOR U865 ( .A(n1401), .B(n1402), .Z(n1396) );
  NOR U866 ( .A(n1403), .B(n1394), .Z(n1402) );
  NOR U867 ( .A(n1404), .B(n1395), .Z(n1401) );
  XOR U868 ( .A(n1405), .B(n1406), .Z(n831) );
  XOR U869 ( .A(n1407), .B(n1408), .Z(n829) );
  XNOR U870 ( .A(n1409), .B(n1410), .Z(n1408) );
  NOR U871 ( .A(n1411), .B(n1410), .Z(n1409) );
  XOR U872 ( .A(n1412), .B(n1413), .Z(n1407) );
  NOR U873 ( .A(n1414), .B(n1405), .Z(n1413) );
  NOR U874 ( .A(n1415), .B(n1406), .Z(n1412) );
  XOR U875 ( .A(n1416), .B(n1417), .Z(n822) );
  XOR U876 ( .A(n1418), .B(n1419), .Z(n820) );
  XNOR U877 ( .A(n1420), .B(n1421), .Z(n1419) );
  NOR U878 ( .A(n1422), .B(n1421), .Z(n1420) );
  XOR U879 ( .A(n1423), .B(n1424), .Z(n1418) );
  NOR U880 ( .A(n1425), .B(n1416), .Z(n1424) );
  NOR U881 ( .A(n1426), .B(n1417), .Z(n1423) );
  XOR U882 ( .A(n1427), .B(n1428), .Z(n813) );
  XOR U883 ( .A(n1429), .B(n1430), .Z(n811) );
  XNOR U884 ( .A(n1431), .B(n1432), .Z(n1430) );
  NOR U885 ( .A(n1433), .B(n1432), .Z(n1431) );
  XOR U886 ( .A(n1434), .B(n1435), .Z(n1429) );
  NOR U887 ( .A(n1436), .B(n1427), .Z(n1435) );
  NOR U888 ( .A(n1437), .B(n1428), .Z(n1434) );
  XOR U889 ( .A(n808), .B(n806), .Z(n809) );
  XNOR U890 ( .A(n1438), .B(n1439), .Z(n145) );
  NOR U891 ( .A(n41), .B(n1438), .Z(n1439) );
  XOR U892 ( .A(n1440), .B(n1441), .Z(n148) );
  AND U893 ( .A(n1442), .B(n1443), .Z(n1441) );
  XNOR U894 ( .A(n44), .B(n1440), .Z(n1443) );
  XOR U895 ( .A(n794), .B(n792), .Z(n44) );
  XOR U896 ( .A(n1444), .B(n160), .Z(n792) );
  XNOR U897 ( .A(n161), .B(n158), .Z(n160) );
  XNOR U898 ( .A(n159), .B(n162), .Z(n158) );
  XNOR U899 ( .A(n163), .B(n787), .Z(n162) );
  XNOR U900 ( .A(n170), .B(n786), .Z(n787) );
  XNOR U901 ( .A(n779), .B(n783), .Z(n786) );
  XNOR U902 ( .A(n778), .B(n776), .Z(n783) );
  XNOR U903 ( .A(n777), .B(n775), .Z(n776) );
  XNOR U904 ( .A(n177), .B(n770), .Z(n775) );
  XOR U905 ( .A(n176), .B(n768), .Z(n770) );
  XNOR U906 ( .A(n769), .B(n764), .Z(n768) );
  XNOR U907 ( .A(n765), .B(n192), .Z(n764) );
  XNOR U908 ( .A(n187), .B(n763), .Z(n192) );
  XNOR U909 ( .A(n186), .B(n758), .Z(n763) );
  XNOR U910 ( .A(n188), .B(n757), .Z(n758) );
  XNOR U911 ( .A(n191), .B(n754), .Z(n757) );
  XNOR U912 ( .A(n197), .B(n753), .Z(n754) );
  XNOR U913 ( .A(n746), .B(n750), .Z(n753) );
  XNOR U914 ( .A(n745), .B(n743), .Z(n750) );
  XNOR U915 ( .A(n744), .B(n742), .Z(n743) );
  XNOR U916 ( .A(n204), .B(n737), .Z(n742) );
  XOR U917 ( .A(n203), .B(n735), .Z(n737) );
  XNOR U918 ( .A(n736), .B(n731), .Z(n735) );
  XNOR U919 ( .A(n732), .B(n219), .Z(n731) );
  XNOR U920 ( .A(n214), .B(n730), .Z(n219) );
  XNOR U921 ( .A(n213), .B(n725), .Z(n730) );
  XNOR U922 ( .A(n215), .B(n724), .Z(n725) );
  XNOR U923 ( .A(n218), .B(n721), .Z(n724) );
  XNOR U924 ( .A(n224), .B(n720), .Z(n721) );
  XNOR U925 ( .A(n713), .B(n717), .Z(n720) );
  XNOR U926 ( .A(n712), .B(n710), .Z(n717) );
  XNOR U927 ( .A(n711), .B(n709), .Z(n710) );
  XNOR U928 ( .A(n231), .B(n704), .Z(n709) );
  XOR U929 ( .A(n230), .B(n702), .Z(n704) );
  XNOR U930 ( .A(n703), .B(n698), .Z(n702) );
  XNOR U931 ( .A(n699), .B(n246), .Z(n698) );
  XNOR U932 ( .A(n241), .B(n697), .Z(n246) );
  XNOR U933 ( .A(n240), .B(n692), .Z(n697) );
  XNOR U934 ( .A(n242), .B(n691), .Z(n692) );
  XNOR U935 ( .A(n245), .B(n688), .Z(n691) );
  XNOR U936 ( .A(n251), .B(n687), .Z(n688) );
  XNOR U937 ( .A(n680), .B(n684), .Z(n687) );
  XNOR U938 ( .A(n679), .B(n677), .Z(n684) );
  XNOR U939 ( .A(n678), .B(n676), .Z(n677) );
  XNOR U940 ( .A(n258), .B(n671), .Z(n676) );
  XOR U941 ( .A(n257), .B(n669), .Z(n671) );
  XNOR U942 ( .A(n670), .B(n665), .Z(n669) );
  XNOR U943 ( .A(n666), .B(n273), .Z(n665) );
  XNOR U944 ( .A(n268), .B(n664), .Z(n273) );
  XNOR U945 ( .A(n267), .B(n659), .Z(n664) );
  XNOR U946 ( .A(n269), .B(n658), .Z(n659) );
  XNOR U947 ( .A(n272), .B(n655), .Z(n658) );
  XNOR U948 ( .A(n278), .B(n654), .Z(n655) );
  XNOR U949 ( .A(n647), .B(n651), .Z(n654) );
  XNOR U950 ( .A(n646), .B(n644), .Z(n651) );
  XNOR U951 ( .A(n645), .B(n643), .Z(n644) );
  XNOR U952 ( .A(n285), .B(n638), .Z(n643) );
  XOR U953 ( .A(n284), .B(n636), .Z(n638) );
  XNOR U954 ( .A(n637), .B(n632), .Z(n636) );
  XNOR U955 ( .A(n633), .B(n300), .Z(n632) );
  XNOR U956 ( .A(n295), .B(n631), .Z(n300) );
  XNOR U957 ( .A(n294), .B(n626), .Z(n631) );
  XNOR U958 ( .A(n296), .B(n625), .Z(n626) );
  XNOR U959 ( .A(n299), .B(n622), .Z(n625) );
  XNOR U960 ( .A(n305), .B(n621), .Z(n622) );
  XNOR U961 ( .A(n614), .B(n618), .Z(n621) );
  XNOR U962 ( .A(n613), .B(n611), .Z(n618) );
  XNOR U963 ( .A(n612), .B(n610), .Z(n611) );
  XNOR U964 ( .A(n312), .B(n605), .Z(n610) );
  XOR U965 ( .A(n311), .B(n603), .Z(n605) );
  XNOR U966 ( .A(n604), .B(n599), .Z(n603) );
  XNOR U967 ( .A(n600), .B(n327), .Z(n599) );
  XNOR U968 ( .A(n322), .B(n598), .Z(n327) );
  XNOR U969 ( .A(n321), .B(n593), .Z(n598) );
  XNOR U970 ( .A(n323), .B(n592), .Z(n593) );
  XNOR U971 ( .A(n326), .B(n589), .Z(n592) );
  XNOR U972 ( .A(n332), .B(n588), .Z(n589) );
  XNOR U973 ( .A(n581), .B(n585), .Z(n588) );
  XNOR U974 ( .A(n580), .B(n578), .Z(n585) );
  XNOR U975 ( .A(n579), .B(n577), .Z(n578) );
  XNOR U976 ( .A(n339), .B(n572), .Z(n577) );
  XOR U977 ( .A(n338), .B(n570), .Z(n572) );
  XNOR U978 ( .A(n571), .B(n566), .Z(n570) );
  XNOR U979 ( .A(n567), .B(n354), .Z(n566) );
  XNOR U980 ( .A(n349), .B(n565), .Z(n354) );
  XNOR U981 ( .A(n348), .B(n560), .Z(n565) );
  XNOR U982 ( .A(n350), .B(n559), .Z(n560) );
  XNOR U983 ( .A(n353), .B(n556), .Z(n559) );
  XNOR U984 ( .A(n359), .B(n555), .Z(n556) );
  XNOR U985 ( .A(n548), .B(n552), .Z(n555) );
  XNOR U986 ( .A(n547), .B(n545), .Z(n552) );
  XNOR U987 ( .A(n546), .B(n544), .Z(n545) );
  XNOR U988 ( .A(n366), .B(n539), .Z(n544) );
  XOR U989 ( .A(n365), .B(n537), .Z(n539) );
  XNOR U990 ( .A(n538), .B(n533), .Z(n537) );
  XNOR U991 ( .A(n534), .B(n381), .Z(n533) );
  XNOR U992 ( .A(n376), .B(n532), .Z(n381) );
  XNOR U993 ( .A(n375), .B(n527), .Z(n532) );
  XNOR U994 ( .A(n377), .B(n526), .Z(n527) );
  XNOR U995 ( .A(n380), .B(n523), .Z(n526) );
  XNOR U996 ( .A(n386), .B(n522), .Z(n523) );
  XNOR U997 ( .A(n515), .B(n519), .Z(n522) );
  XNOR U998 ( .A(n514), .B(n512), .Z(n519) );
  XNOR U999 ( .A(n513), .B(n511), .Z(n512) );
  XNOR U1000 ( .A(n393), .B(n506), .Z(n511) );
  XOR U1001 ( .A(n392), .B(n504), .Z(n506) );
  XNOR U1002 ( .A(n505), .B(n500), .Z(n504) );
  XNOR U1003 ( .A(n501), .B(n408), .Z(n500) );
  XNOR U1004 ( .A(n403), .B(n499), .Z(n408) );
  XNOR U1005 ( .A(n402), .B(n494), .Z(n499) );
  XNOR U1006 ( .A(n404), .B(n493), .Z(n494) );
  XNOR U1007 ( .A(n407), .B(n490), .Z(n493) );
  XNOR U1008 ( .A(n413), .B(n489), .Z(n490) );
  XNOR U1009 ( .A(n482), .B(n486), .Z(n489) );
  XNOR U1010 ( .A(n481), .B(n479), .Z(n486) );
  XNOR U1011 ( .A(n480), .B(n478), .Z(n479) );
  XNOR U1012 ( .A(n420), .B(n473), .Z(n478) );
  XOR U1013 ( .A(n419), .B(n471), .Z(n473) );
  XNOR U1014 ( .A(n472), .B(n467), .Z(n471) );
  XNOR U1015 ( .A(n468), .B(n435), .Z(n467) );
  XNOR U1016 ( .A(n430), .B(n466), .Z(n435) );
  XNOR U1017 ( .A(n429), .B(n461), .Z(n466) );
  XNOR U1018 ( .A(n431), .B(n460), .Z(n461) );
  XNOR U1019 ( .A(n434), .B(n457), .Z(n460) );
  XNOR U1020 ( .A(n440), .B(n456), .Z(n457) );
  XNOR U1021 ( .A(n443), .B(n453), .Z(n456) );
  XOR U1022 ( .A(n442), .B(n450), .Z(n453) );
  XOR U1023 ( .A(n451), .B(n449), .Z(n450) );
  XOR U1024 ( .A(n1445), .B(n1446), .Z(n449) );
  XOR U1025 ( .A(n1447), .B(n1448), .Z(n1446) );
  XOR U1026 ( .A(n1449), .B(n1450), .Z(n1448) );
  NOR U1027 ( .A(n1451), .B(n1452), .Z(n1450) );
  NOR U1028 ( .A(n1453), .B(n1454), .Z(n1449) );
  NOR U1029 ( .A(n1455), .B(n1456), .Z(n1447) );
  XOR U1030 ( .A(n1457), .B(n1458), .Z(n1445) );
  XOR U1031 ( .A(n1459), .B(n1460), .Z(n1458) );
  XOR U1032 ( .A(n1461), .B(n1462), .Z(n1460) );
  XNOR U1033 ( .A(n1463), .B(n1464), .Z(n1462) );
  XOR U1034 ( .A(n1465), .B(n1466), .Z(n1464) );
  XOR U1035 ( .A(n1467), .B(n1468), .Z(n1466) );
  XOR U1036 ( .A(n1469), .B(n1470), .Z(n1468) );
  XOR U1037 ( .A(n1471), .B(n1472), .Z(n1467) );
  XOR U1038 ( .A(n1473), .B(n1474), .Z(n1472) );
  XOR U1039 ( .A(n1475), .B(n1476), .Z(n1474) );
  XOR U1040 ( .A(n1477), .B(n1478), .Z(n1476) );
  XNOR U1041 ( .A(n1479), .B(n1480), .Z(n1478) );
  XOR U1042 ( .A(n1481), .B(n1482), .Z(n1477) );
  XOR U1043 ( .A(n1483), .B(n1484), .Z(n1482) );
  AND U1044 ( .A(n1485), .B(n1486), .Z(n1483) );
  XOR U1045 ( .A(n1487), .B(n1488), .Z(n1475) );
  XOR U1046 ( .A(n1489), .B(n1490), .Z(n1488) );
  XOR U1047 ( .A(n1491), .B(n1492), .Z(n1490) );
  XOR U1048 ( .A(n1493), .B(n1494), .Z(n1492) );
  XOR U1049 ( .A(n1495), .B(n1496), .Z(n1494) );
  XOR U1050 ( .A(n1497), .B(n1498), .Z(n1496) );
  XOR U1051 ( .A(n1499), .B(n1500), .Z(n1498) );
  XOR U1052 ( .A(n1501), .B(n1502), .Z(n1500) );
  XOR U1053 ( .A(n1503), .B(n1504), .Z(n1502) );
  XOR U1054 ( .A(n1505), .B(n1506), .Z(n1504) );
  XOR U1055 ( .A(n1507), .B(n1508), .Z(n1506) );
  XOR U1056 ( .A(n1509), .B(n1510), .Z(n1508) );
  AND U1057 ( .A(n1511), .B(n1512), .Z(n1510) );
  NOR U1058 ( .A(n1513), .B(n1514), .Z(n1512) );
  NOR U1059 ( .A(n1515), .B(n1516), .Z(n1511) );
  AND U1060 ( .A(n1517), .B(n1518), .Z(n1516) );
  AND U1061 ( .A(n1519), .B(n1520), .Z(n1509) );
  NOR U1062 ( .A(n1521), .B(n1522), .Z(n1520) );
  NOR U1063 ( .A(n1523), .B(n1524), .Z(n1519) );
  AND U1064 ( .A(n1525), .B(n1526), .Z(n1524) );
  XOR U1065 ( .A(n1527), .B(n1528), .Z(n1507) );
  NOR U1066 ( .A(n1529), .B(n1530), .Z(n1528) );
  XOR U1067 ( .A(n1531), .B(n1532), .Z(n1530) );
  AND U1068 ( .A(n1533), .B(n1534), .Z(n1532) );
  NOR U1069 ( .A(n1535), .B(n1536), .Z(n1534) );
  NOR U1070 ( .A(n1537), .B(n1538), .Z(n1533) );
  AND U1071 ( .A(n1539), .B(n1540), .Z(n1538) );
  AND U1072 ( .A(n1541), .B(n1542), .Z(n1531) );
  NOR U1073 ( .A(n1543), .B(n1544), .Z(n1542) );
  AND U1074 ( .A(n1536), .B(n1545), .Z(n1544) );
  AND U1075 ( .A(n1537), .B(n1546), .Z(n1543) );
  NOR U1076 ( .A(n1547), .B(n1548), .Z(n1541) );
  XOR U1077 ( .A(n1549), .B(n1550), .Z(n1548) );
  AND U1078 ( .A(n1551), .B(n1552), .Z(n1550) );
  NOR U1079 ( .A(n1553), .B(n1554), .Z(n1552) );
  NOR U1080 ( .A(n1555), .B(n1556), .Z(n1551) );
  AND U1081 ( .A(n1557), .B(n1558), .Z(n1556) );
  AND U1082 ( .A(n1559), .B(n1560), .Z(n1549) );
  NOR U1083 ( .A(n1561), .B(n1562), .Z(n1560) );
  AND U1084 ( .A(n1554), .B(n1563), .Z(n1562) );
  AND U1085 ( .A(n1555), .B(n1564), .Z(n1561) );
  NOR U1086 ( .A(n1565), .B(n1566), .Z(n1559) );
  AND U1087 ( .A(n1567), .B(n1568), .Z(n1566) );
  AND U1088 ( .A(n1569), .B(n1570), .Z(n1568) );
  AND U1089 ( .A(n1571), .B(n1572), .Z(n1570) );
  NOR U1090 ( .A(n1573), .B(n1574), .Z(n1571) );
  NOR U1091 ( .A(n1575), .B(n1576), .Z(n1569) );
  AND U1092 ( .A(n1577), .B(n1578), .Z(n1567) );
  NOR U1093 ( .A(n1579), .B(n1580), .Z(n1578) );
  NOR U1094 ( .A(n1581), .B(n1582), .Z(n1577) );
  AND U1095 ( .A(n1553), .B(n1583), .Z(n1565) );
  AND U1096 ( .A(n1535), .B(n1584), .Z(n1547) );
  AND U1097 ( .A(n1521), .B(n1585), .Z(n1529) );
  NOR U1098 ( .A(n1586), .B(n1587), .Z(n1527) );
  AND U1099 ( .A(n1522), .B(n1588), .Z(n1587) );
  AND U1100 ( .A(n1523), .B(n1589), .Z(n1586) );
  XOR U1101 ( .A(n1590), .B(n1591), .Z(n1505) );
  XOR U1102 ( .A(n1592), .B(n1593), .Z(n1591) );
  NOR U1103 ( .A(n1594), .B(n1595), .Z(n1593) );
  AND U1104 ( .A(n1514), .B(n1596), .Z(n1595) );
  AND U1105 ( .A(n1515), .B(n1597), .Z(n1594) );
  NOR U1106 ( .A(n1598), .B(n1599), .Z(n1592) );
  AND U1107 ( .A(n1600), .B(n1601), .Z(n1599) );
  AND U1108 ( .A(n1602), .B(n1603), .Z(n1598) );
  XOR U1109 ( .A(n1604), .B(n1605), .Z(n1590) );
  AND U1110 ( .A(n1513), .B(n1606), .Z(n1605) );
  AND U1111 ( .A(n1607), .B(n1608), .Z(n1604) );
  AND U1112 ( .A(n1609), .B(n1610), .Z(n1503) );
  NOR U1113 ( .A(n1611), .B(n1612), .Z(n1610) );
  NOR U1114 ( .A(n1613), .B(n1614), .Z(n1609) );
  AND U1115 ( .A(n1615), .B(n1616), .Z(n1614) );
  XOR U1116 ( .A(n1617), .B(n1618), .Z(n1501) );
  AND U1117 ( .A(n1619), .B(n1620), .Z(n1618) );
  NOR U1118 ( .A(n1621), .B(n1622), .Z(n1620) );
  NOR U1119 ( .A(n1623), .B(n1624), .Z(n1619) );
  AND U1120 ( .A(n1625), .B(n1626), .Z(n1624) );
  AND U1121 ( .A(n1627), .B(n1628), .Z(n1617) );
  NOR U1122 ( .A(n1607), .B(n1600), .Z(n1628) );
  NOR U1123 ( .A(n1602), .B(n1629), .Z(n1627) );
  AND U1124 ( .A(n1630), .B(n1631), .Z(n1629) );
  XOR U1125 ( .A(n1632), .B(n1633), .Z(n1499) );
  XOR U1126 ( .A(n1634), .B(n1635), .Z(n1633) );
  NOR U1127 ( .A(n1636), .B(n1637), .Z(n1635) );
  AND U1128 ( .A(n1622), .B(n1638), .Z(n1637) );
  AND U1129 ( .A(n1623), .B(n1639), .Z(n1636) );
  NOR U1130 ( .A(n1640), .B(n1641), .Z(n1634) );
  AND U1131 ( .A(n1612), .B(n1642), .Z(n1641) );
  AND U1132 ( .A(n1613), .B(n1643), .Z(n1640) );
  XOR U1133 ( .A(n1644), .B(n1645), .Z(n1632) );
  AND U1134 ( .A(n1621), .B(n1646), .Z(n1645) );
  AND U1135 ( .A(n1611), .B(n1647), .Z(n1644) );
  NOR U1136 ( .A(n1648), .B(n1649), .Z(n1497) );
  AND U1137 ( .A(n1650), .B(n1651), .Z(n1649) );
  XOR U1138 ( .A(n1652), .B(n1653), .Z(n1495) );
  NOR U1139 ( .A(n1654), .B(n1655), .Z(n1653) );
  AND U1140 ( .A(n1656), .B(n1657), .Z(n1652) );
  NOR U1141 ( .A(n1658), .B(n1659), .Z(n1657) );
  NOR U1142 ( .A(n1660), .B(n1661), .Z(n1656) );
  AND U1143 ( .A(n1662), .B(n1663), .Z(n1661) );
  XOR U1144 ( .A(n1664), .B(n1665), .Z(n1493) );
  XOR U1145 ( .A(n1666), .B(n1667), .Z(n1665) );
  NOR U1146 ( .A(n1668), .B(n1669), .Z(n1667) );
  AND U1147 ( .A(n1659), .B(n1670), .Z(n1669) );
  AND U1148 ( .A(n1660), .B(n1671), .Z(n1668) );
  NOR U1149 ( .A(n1672), .B(n1673), .Z(n1666) );
  AND U1150 ( .A(n1655), .B(n1674), .Z(n1673) );
  AND U1151 ( .A(n1648), .B(n1675), .Z(n1672) );
  XOR U1152 ( .A(n1676), .B(n1677), .Z(n1664) );
  AND U1153 ( .A(n1658), .B(n1678), .Z(n1677) );
  AND U1154 ( .A(n1654), .B(n1679), .Z(n1676) );
  NOR U1155 ( .A(n1680), .B(n1681), .Z(n1491) );
  XOR U1156 ( .A(n1682), .B(n1683), .Z(n1489) );
  XOR U1157 ( .A(n1684), .B(n1685), .Z(n1487) );
  XOR U1158 ( .A(n1686), .B(n1687), .Z(n1685) );
  AND U1159 ( .A(n1680), .B(n1688), .Z(n1687) );
  AND U1160 ( .A(n1681), .B(n1689), .Z(n1686) );
  XOR U1161 ( .A(n1690), .B(n1691), .Z(n1684) );
  AND U1162 ( .A(n1682), .B(n1692), .Z(n1691) );
  AND U1163 ( .A(n1683), .B(n1693), .Z(n1690) );
  XOR U1164 ( .A(n1694), .B(n1695), .Z(n1473) );
  AND U1165 ( .A(n1484), .B(n1696), .Z(n1695) );
  AND U1166 ( .A(n1697), .B(n1481), .Z(n1694) );
  XOR U1167 ( .A(n1698), .B(n1699), .Z(n1471) );
  XOR U1168 ( .A(n1700), .B(n1701), .Z(n1699) );
  AND U1169 ( .A(n1702), .B(n1479), .Z(n1701) );
  NOR U1170 ( .A(n1703), .B(n1704), .Z(n1700) );
  XOR U1171 ( .A(n1705), .B(n1706), .Z(n1698) );
  AND U1172 ( .A(n1707), .B(n1708), .Z(n1706) );
  NOR U1173 ( .A(n1709), .B(n1469), .Z(n1705) );
  XOR U1174 ( .A(n1710), .B(n1711), .Z(n1465) );
  XNOR U1175 ( .A(n1704), .B(n1708), .Z(n1711) );
  XOR U1176 ( .A(n1712), .B(n1713), .Z(n1710) );
  NOR U1177 ( .A(n1714), .B(n1470), .Z(n1713) );
  NOR U1178 ( .A(n1715), .B(n1716), .Z(n1712) );
  XOR U1179 ( .A(n1717), .B(n1718), .Z(n1461) );
  XOR U1180 ( .A(n1719), .B(n1720), .Z(n1459) );
  XNOR U1181 ( .A(n1721), .B(n1716), .Z(n1720) );
  NOR U1182 ( .A(n1722), .B(n1717), .Z(n1721) );
  XOR U1183 ( .A(n1723), .B(n1724), .Z(n1719) );
  NOR U1184 ( .A(n1725), .B(n1718), .Z(n1724) );
  NOR U1185 ( .A(n1726), .B(n1463), .Z(n1723) );
  XOR U1186 ( .A(n1727), .B(n1728), .Z(n1457) );
  XNOR U1187 ( .A(n1452), .B(n1729), .Z(n1728) );
  XNOR U1188 ( .A(n1730), .B(n1456), .Z(n1729) );
  NOR U1189 ( .A(n1731), .B(n1732), .Z(n1730) );
  XNOR U1190 ( .A(n1732), .B(n1454), .Z(n1727) );
  XNOR U1191 ( .A(n1733), .B(n1734), .Z(n451) );
  NOR U1192 ( .A(n1735), .B(n1733), .Z(n1734) );
  XOR U1193 ( .A(n1736), .B(n1737), .Z(n442) );
  NOR U1194 ( .A(n1738), .B(n1736), .Z(n1737) );
  XOR U1195 ( .A(n1739), .B(n1740), .Z(n443) );
  NOR U1196 ( .A(n1741), .B(n1739), .Z(n1740) );
  XOR U1197 ( .A(n1742), .B(n1743), .Z(n440) );
  NOR U1198 ( .A(n1744), .B(n1742), .Z(n1743) );
  XOR U1199 ( .A(n1745), .B(n1746), .Z(n434) );
  NOR U1200 ( .A(n1747), .B(n1745), .Z(n1746) );
  XOR U1201 ( .A(n1748), .B(n1749), .Z(n431) );
  NOR U1202 ( .A(n1750), .B(n1748), .Z(n1749) );
  XOR U1203 ( .A(n1751), .B(n1752), .Z(n429) );
  NOR U1204 ( .A(n1753), .B(n1751), .Z(n1752) );
  XOR U1205 ( .A(n1754), .B(n1755), .Z(n430) );
  NOR U1206 ( .A(n1756), .B(n1754), .Z(n1755) );
  XOR U1207 ( .A(n1757), .B(n1758), .Z(n468) );
  NOR U1208 ( .A(n1759), .B(n1757), .Z(n1758) );
  XNOR U1209 ( .A(n1760), .B(n1761), .Z(n472) );
  NOR U1210 ( .A(n1762), .B(n1760), .Z(n1761) );
  XOR U1211 ( .A(n1763), .B(n1764), .Z(n419) );
  NOR U1212 ( .A(n1765), .B(n1763), .Z(n1764) );
  XOR U1213 ( .A(n1766), .B(n1767), .Z(n420) );
  NOR U1214 ( .A(n1768), .B(n1766), .Z(n1767) );
  XOR U1215 ( .A(n1769), .B(n1770), .Z(n480) );
  NOR U1216 ( .A(n1771), .B(n1769), .Z(n1770) );
  XOR U1217 ( .A(n1772), .B(n1773), .Z(n481) );
  NOR U1218 ( .A(n1774), .B(n1772), .Z(n1773) );
  XOR U1219 ( .A(n1775), .B(n1776), .Z(n482) );
  NOR U1220 ( .A(n1777), .B(n1775), .Z(n1776) );
  XOR U1221 ( .A(n1778), .B(n1779), .Z(n413) );
  NOR U1222 ( .A(n1780), .B(n1778), .Z(n1779) );
  XOR U1223 ( .A(n1781), .B(n1782), .Z(n407) );
  NOR U1224 ( .A(n1783), .B(n1781), .Z(n1782) );
  XOR U1225 ( .A(n1784), .B(n1785), .Z(n404) );
  NOR U1226 ( .A(n1786), .B(n1784), .Z(n1785) );
  XOR U1227 ( .A(n1787), .B(n1788), .Z(n402) );
  NOR U1228 ( .A(n1789), .B(n1787), .Z(n1788) );
  XOR U1229 ( .A(n1790), .B(n1791), .Z(n403) );
  NOR U1230 ( .A(n1792), .B(n1790), .Z(n1791) );
  XOR U1231 ( .A(n1793), .B(n1794), .Z(n501) );
  NOR U1232 ( .A(n1795), .B(n1793), .Z(n1794) );
  XNOR U1233 ( .A(n1796), .B(n1797), .Z(n505) );
  NOR U1234 ( .A(n1798), .B(n1796), .Z(n1797) );
  XOR U1235 ( .A(n1799), .B(n1800), .Z(n392) );
  NOR U1236 ( .A(n1801), .B(n1799), .Z(n1800) );
  XOR U1237 ( .A(n1802), .B(n1803), .Z(n393) );
  NOR U1238 ( .A(n1804), .B(n1802), .Z(n1803) );
  XOR U1239 ( .A(n1805), .B(n1806), .Z(n513) );
  NOR U1240 ( .A(n1807), .B(n1805), .Z(n1806) );
  XOR U1241 ( .A(n1808), .B(n1809), .Z(n514) );
  NOR U1242 ( .A(n1810), .B(n1808), .Z(n1809) );
  XOR U1243 ( .A(n1811), .B(n1812), .Z(n515) );
  NOR U1244 ( .A(n1813), .B(n1811), .Z(n1812) );
  XOR U1245 ( .A(n1814), .B(n1815), .Z(n386) );
  NOR U1246 ( .A(n1816), .B(n1814), .Z(n1815) );
  XOR U1247 ( .A(n1817), .B(n1818), .Z(n380) );
  NOR U1248 ( .A(n1819), .B(n1817), .Z(n1818) );
  XOR U1249 ( .A(n1820), .B(n1821), .Z(n377) );
  NOR U1250 ( .A(n1822), .B(n1820), .Z(n1821) );
  XOR U1251 ( .A(n1823), .B(n1824), .Z(n375) );
  NOR U1252 ( .A(n1825), .B(n1823), .Z(n1824) );
  XOR U1253 ( .A(n1826), .B(n1827), .Z(n376) );
  NOR U1254 ( .A(n1828), .B(n1826), .Z(n1827) );
  XOR U1255 ( .A(n1829), .B(n1830), .Z(n534) );
  NOR U1256 ( .A(n1831), .B(n1829), .Z(n1830) );
  XNOR U1257 ( .A(n1832), .B(n1833), .Z(n538) );
  NOR U1258 ( .A(n1834), .B(n1832), .Z(n1833) );
  XOR U1259 ( .A(n1835), .B(n1836), .Z(n365) );
  NOR U1260 ( .A(n1837), .B(n1835), .Z(n1836) );
  XOR U1261 ( .A(n1838), .B(n1839), .Z(n366) );
  NOR U1262 ( .A(n1840), .B(n1838), .Z(n1839) );
  XOR U1263 ( .A(n1841), .B(n1842), .Z(n546) );
  NOR U1264 ( .A(n1843), .B(n1841), .Z(n1842) );
  XOR U1265 ( .A(n1844), .B(n1845), .Z(n547) );
  NOR U1266 ( .A(n1846), .B(n1844), .Z(n1845) );
  XOR U1267 ( .A(n1847), .B(n1848), .Z(n548) );
  NOR U1268 ( .A(n1849), .B(n1847), .Z(n1848) );
  XOR U1269 ( .A(n1850), .B(n1851), .Z(n359) );
  NOR U1270 ( .A(n1852), .B(n1850), .Z(n1851) );
  XOR U1271 ( .A(n1853), .B(n1854), .Z(n353) );
  NOR U1272 ( .A(n1855), .B(n1853), .Z(n1854) );
  XOR U1273 ( .A(n1856), .B(n1857), .Z(n350) );
  NOR U1274 ( .A(n1858), .B(n1856), .Z(n1857) );
  XOR U1275 ( .A(n1859), .B(n1860), .Z(n348) );
  NOR U1276 ( .A(n1861), .B(n1859), .Z(n1860) );
  XOR U1277 ( .A(n1862), .B(n1863), .Z(n349) );
  NOR U1278 ( .A(n1864), .B(n1862), .Z(n1863) );
  XOR U1279 ( .A(n1865), .B(n1866), .Z(n567) );
  NOR U1280 ( .A(n1867), .B(n1865), .Z(n1866) );
  XNOR U1281 ( .A(n1868), .B(n1869), .Z(n571) );
  NOR U1282 ( .A(n1870), .B(n1868), .Z(n1869) );
  XOR U1283 ( .A(n1871), .B(n1872), .Z(n338) );
  NOR U1284 ( .A(n1873), .B(n1871), .Z(n1872) );
  XOR U1285 ( .A(n1874), .B(n1875), .Z(n339) );
  NOR U1286 ( .A(n1876), .B(n1874), .Z(n1875) );
  XOR U1287 ( .A(n1877), .B(n1878), .Z(n579) );
  NOR U1288 ( .A(n1879), .B(n1877), .Z(n1878) );
  XOR U1289 ( .A(n1880), .B(n1881), .Z(n580) );
  NOR U1290 ( .A(n1882), .B(n1880), .Z(n1881) );
  XOR U1291 ( .A(n1883), .B(n1884), .Z(n581) );
  NOR U1292 ( .A(n1885), .B(n1883), .Z(n1884) );
  XOR U1293 ( .A(n1886), .B(n1887), .Z(n332) );
  NOR U1294 ( .A(n1888), .B(n1886), .Z(n1887) );
  XOR U1295 ( .A(n1889), .B(n1890), .Z(n326) );
  NOR U1296 ( .A(n1891), .B(n1889), .Z(n1890) );
  XOR U1297 ( .A(n1892), .B(n1893), .Z(n323) );
  NOR U1298 ( .A(n1894), .B(n1892), .Z(n1893) );
  XOR U1299 ( .A(n1895), .B(n1896), .Z(n321) );
  NOR U1300 ( .A(n1897), .B(n1895), .Z(n1896) );
  XOR U1301 ( .A(n1898), .B(n1899), .Z(n322) );
  NOR U1302 ( .A(n1900), .B(n1898), .Z(n1899) );
  XOR U1303 ( .A(n1901), .B(n1902), .Z(n600) );
  NOR U1304 ( .A(n1903), .B(n1901), .Z(n1902) );
  XNOR U1305 ( .A(n1904), .B(n1905), .Z(n604) );
  NOR U1306 ( .A(n1906), .B(n1904), .Z(n1905) );
  XOR U1307 ( .A(n1907), .B(n1908), .Z(n311) );
  NOR U1308 ( .A(n1909), .B(n1907), .Z(n1908) );
  XOR U1309 ( .A(n1910), .B(n1911), .Z(n312) );
  NOR U1310 ( .A(n1912), .B(n1910), .Z(n1911) );
  XOR U1311 ( .A(n1913), .B(n1914), .Z(n612) );
  NOR U1312 ( .A(n1915), .B(n1913), .Z(n1914) );
  XOR U1313 ( .A(n1916), .B(n1917), .Z(n613) );
  NOR U1314 ( .A(n1918), .B(n1916), .Z(n1917) );
  XOR U1315 ( .A(n1919), .B(n1920), .Z(n614) );
  NOR U1316 ( .A(n1921), .B(n1919), .Z(n1920) );
  XOR U1317 ( .A(n1922), .B(n1923), .Z(n305) );
  NOR U1318 ( .A(n1924), .B(n1922), .Z(n1923) );
  XOR U1319 ( .A(n1925), .B(n1926), .Z(n299) );
  NOR U1320 ( .A(n1927), .B(n1925), .Z(n1926) );
  XOR U1321 ( .A(n1928), .B(n1929), .Z(n296) );
  NOR U1322 ( .A(n1930), .B(n1928), .Z(n1929) );
  XOR U1323 ( .A(n1931), .B(n1932), .Z(n294) );
  NOR U1324 ( .A(n1933), .B(n1931), .Z(n1932) );
  XOR U1325 ( .A(n1934), .B(n1935), .Z(n295) );
  NOR U1326 ( .A(n1936), .B(n1934), .Z(n1935) );
  XOR U1327 ( .A(n1937), .B(n1938), .Z(n633) );
  NOR U1328 ( .A(n1939), .B(n1937), .Z(n1938) );
  XNOR U1329 ( .A(n1940), .B(n1941), .Z(n637) );
  NOR U1330 ( .A(n1942), .B(n1940), .Z(n1941) );
  XOR U1331 ( .A(n1943), .B(n1944), .Z(n284) );
  NOR U1332 ( .A(n1945), .B(n1943), .Z(n1944) );
  XOR U1333 ( .A(n1946), .B(n1947), .Z(n285) );
  NOR U1334 ( .A(n1948), .B(n1946), .Z(n1947) );
  XOR U1335 ( .A(n1949), .B(n1950), .Z(n645) );
  NOR U1336 ( .A(n1951), .B(n1949), .Z(n1950) );
  XOR U1337 ( .A(n1952), .B(n1953), .Z(n646) );
  NOR U1338 ( .A(n1954), .B(n1952), .Z(n1953) );
  XOR U1339 ( .A(n1955), .B(n1956), .Z(n647) );
  NOR U1340 ( .A(n1957), .B(n1955), .Z(n1956) );
  XOR U1341 ( .A(n1958), .B(n1959), .Z(n278) );
  NOR U1342 ( .A(n1960), .B(n1958), .Z(n1959) );
  XOR U1343 ( .A(n1961), .B(n1962), .Z(n272) );
  NOR U1344 ( .A(n1963), .B(n1961), .Z(n1962) );
  XOR U1345 ( .A(n1964), .B(n1965), .Z(n269) );
  NOR U1346 ( .A(n1966), .B(n1964), .Z(n1965) );
  XOR U1347 ( .A(n1967), .B(n1968), .Z(n267) );
  NOR U1348 ( .A(n1969), .B(n1967), .Z(n1968) );
  XOR U1349 ( .A(n1970), .B(n1971), .Z(n268) );
  NOR U1350 ( .A(n1972), .B(n1970), .Z(n1971) );
  XOR U1351 ( .A(n1973), .B(n1974), .Z(n666) );
  NOR U1352 ( .A(n1975), .B(n1973), .Z(n1974) );
  XNOR U1353 ( .A(n1976), .B(n1977), .Z(n670) );
  NOR U1354 ( .A(n1978), .B(n1976), .Z(n1977) );
  XOR U1355 ( .A(n1979), .B(n1980), .Z(n257) );
  NOR U1356 ( .A(n1981), .B(n1979), .Z(n1980) );
  XOR U1357 ( .A(n1982), .B(n1983), .Z(n258) );
  NOR U1358 ( .A(n1984), .B(n1982), .Z(n1983) );
  XOR U1359 ( .A(n1985), .B(n1986), .Z(n678) );
  NOR U1360 ( .A(n1987), .B(n1985), .Z(n1986) );
  XOR U1361 ( .A(n1988), .B(n1989), .Z(n679) );
  NOR U1362 ( .A(n1990), .B(n1988), .Z(n1989) );
  XOR U1363 ( .A(n1991), .B(n1992), .Z(n680) );
  NOR U1364 ( .A(n1993), .B(n1991), .Z(n1992) );
  XOR U1365 ( .A(n1994), .B(n1995), .Z(n251) );
  NOR U1366 ( .A(n1996), .B(n1994), .Z(n1995) );
  XOR U1367 ( .A(n1997), .B(n1998), .Z(n245) );
  NOR U1368 ( .A(n1999), .B(n1997), .Z(n1998) );
  XOR U1369 ( .A(n2000), .B(n2001), .Z(n242) );
  NOR U1370 ( .A(n2002), .B(n2000), .Z(n2001) );
  XOR U1371 ( .A(n2003), .B(n2004), .Z(n240) );
  NOR U1372 ( .A(n2005), .B(n2003), .Z(n2004) );
  XOR U1373 ( .A(n2006), .B(n2007), .Z(n241) );
  NOR U1374 ( .A(n2008), .B(n2006), .Z(n2007) );
  XOR U1375 ( .A(n2009), .B(n2010), .Z(n699) );
  NOR U1376 ( .A(n2011), .B(n2009), .Z(n2010) );
  XNOR U1377 ( .A(n2012), .B(n2013), .Z(n703) );
  NOR U1378 ( .A(n2014), .B(n2012), .Z(n2013) );
  XOR U1379 ( .A(n2015), .B(n2016), .Z(n230) );
  NOR U1380 ( .A(n2017), .B(n2015), .Z(n2016) );
  XOR U1381 ( .A(n2018), .B(n2019), .Z(n231) );
  NOR U1382 ( .A(n2020), .B(n2018), .Z(n2019) );
  XOR U1383 ( .A(n2021), .B(n2022), .Z(n711) );
  NOR U1384 ( .A(n2023), .B(n2021), .Z(n2022) );
  XOR U1385 ( .A(n2024), .B(n2025), .Z(n712) );
  NOR U1386 ( .A(n2026), .B(n2024), .Z(n2025) );
  XOR U1387 ( .A(n2027), .B(n2028), .Z(n713) );
  NOR U1388 ( .A(n2029), .B(n2027), .Z(n2028) );
  XOR U1389 ( .A(n2030), .B(n2031), .Z(n224) );
  NOR U1390 ( .A(n2032), .B(n2030), .Z(n2031) );
  XOR U1391 ( .A(n2033), .B(n2034), .Z(n218) );
  NOR U1392 ( .A(n2035), .B(n2033), .Z(n2034) );
  XOR U1393 ( .A(n2036), .B(n2037), .Z(n215) );
  NOR U1394 ( .A(n2038), .B(n2036), .Z(n2037) );
  XOR U1395 ( .A(n2039), .B(n2040), .Z(n213) );
  NOR U1396 ( .A(n2041), .B(n2039), .Z(n2040) );
  XOR U1397 ( .A(n2042), .B(n2043), .Z(n214) );
  NOR U1398 ( .A(n2044), .B(n2042), .Z(n2043) );
  XOR U1399 ( .A(n2045), .B(n2046), .Z(n732) );
  NOR U1400 ( .A(n2047), .B(n2045), .Z(n2046) );
  XNOR U1401 ( .A(n2048), .B(n2049), .Z(n736) );
  NOR U1402 ( .A(n2050), .B(n2048), .Z(n2049) );
  XOR U1403 ( .A(n2051), .B(n2052), .Z(n203) );
  NOR U1404 ( .A(n2053), .B(n2051), .Z(n2052) );
  XOR U1405 ( .A(n2054), .B(n2055), .Z(n204) );
  NOR U1406 ( .A(n2056), .B(n2054), .Z(n2055) );
  XOR U1407 ( .A(n2057), .B(n2058), .Z(n744) );
  NOR U1408 ( .A(n2059), .B(n2057), .Z(n2058) );
  XOR U1409 ( .A(n2060), .B(n2061), .Z(n745) );
  NOR U1410 ( .A(n2062), .B(n2060), .Z(n2061) );
  XOR U1411 ( .A(n2063), .B(n2064), .Z(n746) );
  NOR U1412 ( .A(n2065), .B(n2063), .Z(n2064) );
  XOR U1413 ( .A(n2066), .B(n2067), .Z(n197) );
  NOR U1414 ( .A(n2068), .B(n2066), .Z(n2067) );
  XOR U1415 ( .A(n2069), .B(n2070), .Z(n191) );
  NOR U1416 ( .A(n2071), .B(n2069), .Z(n2070) );
  XOR U1417 ( .A(n2072), .B(n2073), .Z(n188) );
  NOR U1418 ( .A(n2074), .B(n2072), .Z(n2073) );
  XOR U1419 ( .A(n2075), .B(n2076), .Z(n186) );
  NOR U1420 ( .A(n2077), .B(n2075), .Z(n2076) );
  XOR U1421 ( .A(n2078), .B(n2079), .Z(n187) );
  NOR U1422 ( .A(n2080), .B(n2078), .Z(n2079) );
  XOR U1423 ( .A(n2081), .B(n2082), .Z(n765) );
  NOR U1424 ( .A(n2083), .B(n2081), .Z(n2082) );
  XNOR U1425 ( .A(n2084), .B(n2085), .Z(n769) );
  NOR U1426 ( .A(n2086), .B(n2084), .Z(n2085) );
  XOR U1427 ( .A(n2087), .B(n2088), .Z(n176) );
  NOR U1428 ( .A(n2089), .B(n2087), .Z(n2088) );
  XOR U1429 ( .A(n2090), .B(n2091), .Z(n177) );
  NOR U1430 ( .A(n2092), .B(n2090), .Z(n2091) );
  XOR U1431 ( .A(n2093), .B(n2094), .Z(n777) );
  NOR U1432 ( .A(n2095), .B(n2093), .Z(n2094) );
  XOR U1433 ( .A(n2096), .B(n2097), .Z(n778) );
  NOR U1434 ( .A(n2098), .B(n2096), .Z(n2097) );
  XOR U1435 ( .A(n2099), .B(n2100), .Z(n779) );
  NOR U1436 ( .A(n2101), .B(n2099), .Z(n2100) );
  XOR U1437 ( .A(n2102), .B(n2103), .Z(n170) );
  NOR U1438 ( .A(n2104), .B(n2102), .Z(n2103) );
  XOR U1439 ( .A(n2105), .B(n2106), .Z(n163) );
  NOR U1440 ( .A(n2107), .B(n2105), .Z(n2106) );
  XOR U1441 ( .A(n2108), .B(n2109), .Z(n159) );
  NOR U1442 ( .A(n2110), .B(n2108), .Z(n2109) );
  XOR U1443 ( .A(n2111), .B(n2112), .Z(n161) );
  NOR U1444 ( .A(n2113), .B(n2111), .Z(n2112) );
  IV U1445 ( .A(n793), .Z(n1444) );
  XOR U1446 ( .A(n2114), .B(n2115), .Z(n793) );
  AND U1447 ( .A(n2116), .B(n2114), .Z(n2115) );
  XNOR U1448 ( .A(n2117), .B(n2118), .Z(n794) );
  AND U1449 ( .A(n58), .B(n2117), .Z(n2118) );
  XOR U1450 ( .A(n1440), .B(n41), .Z(n1442) );
  XNOR U1451 ( .A(n1438), .B(n819), .Z(n41) );
  XOR U1452 ( .A(n818), .B(n807), .Z(n819) );
  XOR U1453 ( .A(n2119), .B(n805), .Z(n807) );
  XNOR U1454 ( .A(n806), .B(n802), .Z(n805) );
  XNOR U1455 ( .A(n801), .B(n828), .Z(n802) );
  XNOR U1456 ( .A(n827), .B(n1437), .Z(n828) );
  XNOR U1457 ( .A(n1428), .B(n1436), .Z(n1437) );
  XNOR U1458 ( .A(n1427), .B(n1433), .Z(n1436) );
  XNOR U1459 ( .A(n1432), .B(n837), .Z(n1433) );
  XNOR U1460 ( .A(n836), .B(n1426), .Z(n837) );
  XNOR U1461 ( .A(n1417), .B(n1425), .Z(n1426) );
  XNOR U1462 ( .A(n1416), .B(n1422), .Z(n1425) );
  XNOR U1463 ( .A(n1421), .B(n846), .Z(n1422) );
  XNOR U1464 ( .A(n845), .B(n1415), .Z(n846) );
  XNOR U1465 ( .A(n1406), .B(n1414), .Z(n1415) );
  XNOR U1466 ( .A(n1405), .B(n1411), .Z(n1414) );
  XNOR U1467 ( .A(n1410), .B(n855), .Z(n1411) );
  XNOR U1468 ( .A(n854), .B(n1404), .Z(n855) );
  XNOR U1469 ( .A(n1395), .B(n1403), .Z(n1404) );
  XNOR U1470 ( .A(n1394), .B(n1400), .Z(n1403) );
  XNOR U1471 ( .A(n1399), .B(n864), .Z(n1400) );
  XNOR U1472 ( .A(n863), .B(n1393), .Z(n864) );
  XNOR U1473 ( .A(n1384), .B(n1392), .Z(n1393) );
  XNOR U1474 ( .A(n1383), .B(n1389), .Z(n1392) );
  XNOR U1475 ( .A(n1388), .B(n873), .Z(n1389) );
  XNOR U1476 ( .A(n872), .B(n1382), .Z(n873) );
  XNOR U1477 ( .A(n1373), .B(n1381), .Z(n1382) );
  XNOR U1478 ( .A(n1372), .B(n1378), .Z(n1381) );
  XNOR U1479 ( .A(n1377), .B(n882), .Z(n1378) );
  XNOR U1480 ( .A(n881), .B(n1371), .Z(n882) );
  XNOR U1481 ( .A(n1362), .B(n1370), .Z(n1371) );
  XNOR U1482 ( .A(n1361), .B(n1367), .Z(n1370) );
  XNOR U1483 ( .A(n1366), .B(n891), .Z(n1367) );
  XNOR U1484 ( .A(n890), .B(n1360), .Z(n891) );
  XNOR U1485 ( .A(n1351), .B(n1359), .Z(n1360) );
  XNOR U1486 ( .A(n1350), .B(n1356), .Z(n1359) );
  XNOR U1487 ( .A(n1355), .B(n900), .Z(n1356) );
  XNOR U1488 ( .A(n899), .B(n1349), .Z(n900) );
  XNOR U1489 ( .A(n1340), .B(n1348), .Z(n1349) );
  XNOR U1490 ( .A(n1339), .B(n1345), .Z(n1348) );
  XNOR U1491 ( .A(n1344), .B(n909), .Z(n1345) );
  XNOR U1492 ( .A(n908), .B(n1338), .Z(n909) );
  XNOR U1493 ( .A(n1329), .B(n1337), .Z(n1338) );
  XNOR U1494 ( .A(n1328), .B(n1334), .Z(n1337) );
  XNOR U1495 ( .A(n1333), .B(n918), .Z(n1334) );
  XNOR U1496 ( .A(n917), .B(n1327), .Z(n918) );
  XNOR U1497 ( .A(n1318), .B(n1326), .Z(n1327) );
  XNOR U1498 ( .A(n1317), .B(n1323), .Z(n1326) );
  XNOR U1499 ( .A(n1322), .B(n927), .Z(n1323) );
  XNOR U1500 ( .A(n926), .B(n1316), .Z(n927) );
  XNOR U1501 ( .A(n1307), .B(n1315), .Z(n1316) );
  XNOR U1502 ( .A(n1306), .B(n1312), .Z(n1315) );
  XNOR U1503 ( .A(n1311), .B(n936), .Z(n1312) );
  XNOR U1504 ( .A(n935), .B(n1305), .Z(n936) );
  XNOR U1505 ( .A(n1296), .B(n1304), .Z(n1305) );
  XNOR U1506 ( .A(n1295), .B(n1301), .Z(n1304) );
  XNOR U1507 ( .A(n1300), .B(n945), .Z(n1301) );
  XNOR U1508 ( .A(n944), .B(n1294), .Z(n945) );
  XNOR U1509 ( .A(n1285), .B(n1293), .Z(n1294) );
  XNOR U1510 ( .A(n1284), .B(n1290), .Z(n1293) );
  XNOR U1511 ( .A(n1289), .B(n954), .Z(n1290) );
  XNOR U1512 ( .A(n953), .B(n1283), .Z(n954) );
  XNOR U1513 ( .A(n1274), .B(n1282), .Z(n1283) );
  XNOR U1514 ( .A(n1273), .B(n1279), .Z(n1282) );
  XNOR U1515 ( .A(n1278), .B(n963), .Z(n1279) );
  XNOR U1516 ( .A(n962), .B(n1272), .Z(n963) );
  XNOR U1517 ( .A(n1263), .B(n1271), .Z(n1272) );
  XNOR U1518 ( .A(n1262), .B(n1268), .Z(n1271) );
  XNOR U1519 ( .A(n1267), .B(n972), .Z(n1268) );
  XNOR U1520 ( .A(n971), .B(n1261), .Z(n972) );
  XNOR U1521 ( .A(n1252), .B(n1260), .Z(n1261) );
  XNOR U1522 ( .A(n1251), .B(n1257), .Z(n1260) );
  XNOR U1523 ( .A(n1256), .B(n981), .Z(n1257) );
  XNOR U1524 ( .A(n980), .B(n1250), .Z(n981) );
  XNOR U1525 ( .A(n1241), .B(n1249), .Z(n1250) );
  XNOR U1526 ( .A(n1240), .B(n1246), .Z(n1249) );
  XNOR U1527 ( .A(n1245), .B(n990), .Z(n1246) );
  XNOR U1528 ( .A(n989), .B(n1239), .Z(n990) );
  XNOR U1529 ( .A(n1230), .B(n1238), .Z(n1239) );
  XNOR U1530 ( .A(n1229), .B(n1235), .Z(n1238) );
  XNOR U1531 ( .A(n1234), .B(n999), .Z(n1235) );
  XNOR U1532 ( .A(n998), .B(n1228), .Z(n999) );
  XNOR U1533 ( .A(n1219), .B(n1227), .Z(n1228) );
  XNOR U1534 ( .A(n1218), .B(n1224), .Z(n1227) );
  XNOR U1535 ( .A(n1223), .B(n1008), .Z(n1224) );
  XNOR U1536 ( .A(n1007), .B(n1217), .Z(n1008) );
  XNOR U1537 ( .A(n1208), .B(n1216), .Z(n1217) );
  XNOR U1538 ( .A(n1207), .B(n1213), .Z(n1216) );
  XNOR U1539 ( .A(n1212), .B(n1017), .Z(n1213) );
  XNOR U1540 ( .A(n1016), .B(n1206), .Z(n1017) );
  XNOR U1541 ( .A(n1197), .B(n1205), .Z(n1206) );
  XNOR U1542 ( .A(n1196), .B(n1202), .Z(n1205) );
  XNOR U1543 ( .A(n1201), .B(n1026), .Z(n1202) );
  XNOR U1544 ( .A(n1025), .B(n1195), .Z(n1026) );
  XNOR U1545 ( .A(n1186), .B(n1194), .Z(n1195) );
  XNOR U1546 ( .A(n1185), .B(n1191), .Z(n1194) );
  XNOR U1547 ( .A(n1190), .B(n1035), .Z(n1191) );
  XNOR U1548 ( .A(n1034), .B(n1184), .Z(n1035) );
  XNOR U1549 ( .A(n1175), .B(n1183), .Z(n1184) );
  XNOR U1550 ( .A(n1174), .B(n1180), .Z(n1183) );
  XNOR U1551 ( .A(n1179), .B(n1044), .Z(n1180) );
  XNOR U1552 ( .A(n1043), .B(n1173), .Z(n1044) );
  XNOR U1553 ( .A(n1164), .B(n1172), .Z(n1173) );
  XNOR U1554 ( .A(n1163), .B(n1169), .Z(n1172) );
  XNOR U1555 ( .A(n1168), .B(n1053), .Z(n1169) );
  XNOR U1556 ( .A(n1052), .B(n1162), .Z(n1053) );
  XNOR U1557 ( .A(n1153), .B(n1161), .Z(n1162) );
  XNOR U1558 ( .A(n1152), .B(n1158), .Z(n1161) );
  XNOR U1559 ( .A(n1157), .B(n1062), .Z(n1158) );
  XNOR U1560 ( .A(n1061), .B(n1151), .Z(n1062) );
  XNOR U1561 ( .A(n1142), .B(n1150), .Z(n1151) );
  XNOR U1562 ( .A(n1141), .B(n1147), .Z(n1150) );
  XNOR U1563 ( .A(n1146), .B(n1071), .Z(n1147) );
  XNOR U1564 ( .A(n1070), .B(n1140), .Z(n1071) );
  XNOR U1565 ( .A(n1131), .B(n1139), .Z(n1140) );
  XNOR U1566 ( .A(n1130), .B(n1136), .Z(n1139) );
  XNOR U1567 ( .A(n1135), .B(n1118), .Z(n1136) );
  XNOR U1568 ( .A(n1077), .B(n1129), .Z(n1118) );
  XNOR U1569 ( .A(n1120), .B(n1128), .Z(n1129) );
  XNOR U1570 ( .A(n1119), .B(n1125), .Z(n1128) );
  XNOR U1571 ( .A(n1124), .B(n1108), .Z(n1125) );
  XNOR U1572 ( .A(n1080), .B(n1117), .Z(n1108) );
  XNOR U1573 ( .A(n1104), .B(n1114), .Z(n1117) );
  XNOR U1574 ( .A(n1107), .B(n1113), .Z(n1114) );
  XNOR U1575 ( .A(n1076), .B(n1103), .Z(n1113) );
  XNOR U1576 ( .A(n1086), .B(n1102), .Z(n1103) );
  XNOR U1577 ( .A(n1089), .B(n1099), .Z(n1102) );
  XOR U1578 ( .A(n1088), .B(n1096), .Z(n1099) );
  XOR U1579 ( .A(n1097), .B(n1095), .Z(n1096) );
  XOR U1580 ( .A(n2120), .B(n2121), .Z(n1095) );
  XOR U1581 ( .A(n2122), .B(n2123), .Z(n2121) );
  XNOR U1582 ( .A(n2124), .B(n2125), .Z(n2123) );
  NOR U1583 ( .A(n2126), .B(n2125), .Z(n2124) );
  XOR U1584 ( .A(n2127), .B(n2128), .Z(n2122) );
  NOR U1585 ( .A(n2129), .B(n2130), .Z(n2128) );
  NOR U1586 ( .A(n2131), .B(n2132), .Z(n2127) );
  XOR U1587 ( .A(n2133), .B(n2134), .Z(n2120) );
  XOR U1588 ( .A(n2135), .B(n2136), .Z(n2134) );
  XOR U1589 ( .A(n2137), .B(n2138), .Z(n2136) );
  XOR U1590 ( .A(n2139), .B(n2140), .Z(n2138) );
  XOR U1591 ( .A(n2141), .B(n2142), .Z(n2140) );
  AND U1592 ( .A(n2143), .B(n2142), .Z(n2141) );
  XOR U1593 ( .A(n2144), .B(n2145), .Z(n2139) );
  XOR U1594 ( .A(n2146), .B(n2147), .Z(n2145) );
  XOR U1595 ( .A(n2148), .B(n2149), .Z(n2147) );
  XNOR U1596 ( .A(n2150), .B(n2151), .Z(n2149) );
  NOR U1597 ( .A(n2152), .B(n2151), .Z(n2150) );
  XOR U1598 ( .A(n2153), .B(n2154), .Z(n2148) );
  XOR U1599 ( .A(n2155), .B(n2156), .Z(n2154) );
  XOR U1600 ( .A(n2157), .B(n2158), .Z(n2156) );
  XNOR U1601 ( .A(n2159), .B(n2160), .Z(n2158) );
  NOR U1602 ( .A(n2161), .B(n2160), .Z(n2159) );
  XOR U1603 ( .A(n2162), .B(n2163), .Z(n2157) );
  XOR U1604 ( .A(n2164), .B(n2165), .Z(n2163) );
  XOR U1605 ( .A(n2166), .B(n2167), .Z(n2165) );
  NOR U1606 ( .A(n2168), .B(n2169), .Z(n2166) );
  XOR U1607 ( .A(n2170), .B(n2171), .Z(n2164) );
  XOR U1608 ( .A(n2172), .B(n2173), .Z(n2171) );
  XOR U1609 ( .A(n2174), .B(n2175), .Z(n2173) );
  XOR U1610 ( .A(n2176), .B(n2177), .Z(n2175) );
  AND U1611 ( .A(n2177), .B(n2178), .Z(n2176) );
  XOR U1612 ( .A(n2179), .B(n2180), .Z(n2174) );
  XOR U1613 ( .A(n2181), .B(n2182), .Z(n2180) );
  XOR U1614 ( .A(n2183), .B(n2184), .Z(n2182) );
  XOR U1615 ( .A(n2185), .B(n2186), .Z(n2184) );
  XOR U1616 ( .A(n2187), .B(n2188), .Z(n2186) );
  XOR U1617 ( .A(n2189), .B(n2190), .Z(n2188) );
  XOR U1618 ( .A(n2191), .B(n2192), .Z(n2190) );
  XOR U1619 ( .A(n2193), .B(n2194), .Z(n2192) );
  XOR U1620 ( .A(n2195), .B(n2196), .Z(n2194) );
  AND U1621 ( .A(n2197), .B(n2198), .Z(n2196) );
  AND U1622 ( .A(n2199), .B(n2200), .Z(n2195) );
  XOR U1623 ( .A(n2201), .B(n2202), .Z(n2193) );
  AND U1624 ( .A(n2203), .B(n2204), .Z(n2202) );
  AND U1625 ( .A(n2205), .B(n2206), .Z(n2201) );
  AND U1626 ( .A(n2207), .B(n2208), .Z(n2206) );
  NOR U1627 ( .A(n2209), .B(n2210), .Z(n2208) );
  IV U1628 ( .A(n2211), .Z(n2209) );
  NOR U1629 ( .A(n2212), .B(n2213), .Z(n2211) );
  NOR U1630 ( .A(n2214), .B(n2215), .Z(n2207) );
  AND U1631 ( .A(n2216), .B(n2217), .Z(n2205) );
  NOR U1632 ( .A(n2218), .B(n2219), .Z(n2217) );
  NOR U1633 ( .A(n2220), .B(n2221), .Z(n2216) );
  XOR U1634 ( .A(n2222), .B(n2223), .Z(n2191) );
  XOR U1635 ( .A(n2224), .B(n2225), .Z(n2223) );
  NOR U1636 ( .A(n2226), .B(n2227), .Z(n2225) );
  NOR U1637 ( .A(n2228), .B(n2229), .Z(n2224) );
  AND U1638 ( .A(n2230), .B(n2231), .Z(n2229) );
  IV U1639 ( .A(n2232), .Z(n2228) );
  NOR U1640 ( .A(n2233), .B(n2234), .Z(n2232) );
  AND U1641 ( .A(n2226), .B(n2235), .Z(n2234) );
  AND U1642 ( .A(n2227), .B(n2236), .Z(n2233) );
  XOR U1643 ( .A(n2237), .B(n2238), .Z(n2222) );
  NOR U1644 ( .A(n2239), .B(n2240), .Z(n2238) );
  NOR U1645 ( .A(n2241), .B(n2242), .Z(n2237) );
  AND U1646 ( .A(n2243), .B(n2244), .Z(n2242) );
  IV U1647 ( .A(n2245), .Z(n2241) );
  NOR U1648 ( .A(n2246), .B(n2247), .Z(n2245) );
  AND U1649 ( .A(n2239), .B(n2248), .Z(n2247) );
  AND U1650 ( .A(n2240), .B(n2249), .Z(n2246) );
  AND U1651 ( .A(n2250), .B(n2251), .Z(n2189) );
  XOR U1652 ( .A(n2252), .B(n2253), .Z(n2187) );
  AND U1653 ( .A(n2254), .B(n2255), .Z(n2253) );
  NOR U1654 ( .A(n2256), .B(n2257), .Z(n2252) );
  XOR U1655 ( .A(n2258), .B(n2259), .Z(n2185) );
  XOR U1656 ( .A(n2260), .B(n2261), .Z(n2259) );
  NOR U1657 ( .A(n2262), .B(n2263), .Z(n2261) );
  AND U1658 ( .A(n2264), .B(n2265), .Z(n2263) );
  IV U1659 ( .A(n2266), .Z(n2262) );
  NOR U1660 ( .A(n2267), .B(n2268), .Z(n2266) );
  AND U1661 ( .A(n2256), .B(n2269), .Z(n2268) );
  AND U1662 ( .A(n2257), .B(n2270), .Z(n2267) );
  NOR U1663 ( .A(n2271), .B(n2272), .Z(n2260) );
  XOR U1664 ( .A(n2273), .B(n2274), .Z(n2258) );
  NOR U1665 ( .A(n2275), .B(n2276), .Z(n2274) );
  AND U1666 ( .A(n2277), .B(n2278), .Z(n2276) );
  IV U1667 ( .A(n2279), .Z(n2275) );
  NOR U1668 ( .A(n2280), .B(n2281), .Z(n2279) );
  AND U1669 ( .A(n2271), .B(n2282), .Z(n2281) );
  AND U1670 ( .A(n2272), .B(n2283), .Z(n2280) );
  NOR U1671 ( .A(n2284), .B(n2285), .Z(n2273) );
  AND U1672 ( .A(n2286), .B(n2287), .Z(n2183) );
  XOR U1673 ( .A(n2288), .B(n2289), .Z(n2181) );
  AND U1674 ( .A(n2290), .B(n2291), .Z(n2289) );
  NOR U1675 ( .A(n2292), .B(n2293), .Z(n2288) );
  AND U1676 ( .A(n2294), .B(n2295), .Z(n2293) );
  IV U1677 ( .A(n2296), .Z(n2292) );
  NOR U1678 ( .A(n2297), .B(n2298), .Z(n2296) );
  AND U1679 ( .A(n2284), .B(n2299), .Z(n2298) );
  AND U1680 ( .A(n2285), .B(n2300), .Z(n2297) );
  XOR U1681 ( .A(n2301), .B(n2302), .Z(n2179) );
  XOR U1682 ( .A(n2303), .B(n2304), .Z(n2302) );
  NOR U1683 ( .A(n2305), .B(n2306), .Z(n2304) );
  NOR U1684 ( .A(n2307), .B(n2308), .Z(n2303) );
  AND U1685 ( .A(n2309), .B(n2310), .Z(n2308) );
  IV U1686 ( .A(n2311), .Z(n2307) );
  NOR U1687 ( .A(n2312), .B(n2313), .Z(n2311) );
  AND U1688 ( .A(n2305), .B(n2314), .Z(n2313) );
  AND U1689 ( .A(n2306), .B(n2315), .Z(n2312) );
  XOR U1690 ( .A(n2316), .B(n2317), .Z(n2301) );
  NOR U1691 ( .A(n2318), .B(n2319), .Z(n2317) );
  NOR U1692 ( .A(n2320), .B(n2321), .Z(n2316) );
  AND U1693 ( .A(n2322), .B(n2323), .Z(n2321) );
  IV U1694 ( .A(n2324), .Z(n2320) );
  NOR U1695 ( .A(n2325), .B(n2326), .Z(n2324) );
  AND U1696 ( .A(n2318), .B(n2327), .Z(n2326) );
  AND U1697 ( .A(n2319), .B(n2328), .Z(n2325) );
  XOR U1698 ( .A(n2329), .B(n2330), .Z(n2172) );
  AND U1699 ( .A(n2331), .B(n2332), .Z(n2330) );
  AND U1700 ( .A(n2333), .B(n2334), .Z(n2329) );
  XOR U1701 ( .A(n2335), .B(n2336), .Z(n2170) );
  XOR U1702 ( .A(n2337), .B(n2338), .Z(n2336) );
  NOR U1703 ( .A(n2339), .B(n2340), .Z(n2338) );
  NOR U1704 ( .A(n2341), .B(n2342), .Z(n2337) );
  AND U1705 ( .A(n2343), .B(n2344), .Z(n2342) );
  IV U1706 ( .A(n2345), .Z(n2341) );
  NOR U1707 ( .A(n2346), .B(n2347), .Z(n2345) );
  AND U1708 ( .A(n2339), .B(n2348), .Z(n2347) );
  AND U1709 ( .A(n2340), .B(n2349), .Z(n2346) );
  XOR U1710 ( .A(n2350), .B(n2351), .Z(n2335) );
  NOR U1711 ( .A(n2352), .B(n2353), .Z(n2351) );
  NOR U1712 ( .A(n2354), .B(n2355), .Z(n2350) );
  AND U1713 ( .A(n2356), .B(n2357), .Z(n2355) );
  IV U1714 ( .A(n2358), .Z(n2354) );
  NOR U1715 ( .A(n2359), .B(n2360), .Z(n2358) );
  AND U1716 ( .A(n2352), .B(n2361), .Z(n2360) );
  AND U1717 ( .A(n2353), .B(n2362), .Z(n2359) );
  XOR U1718 ( .A(n2363), .B(n2364), .Z(n2162) );
  XOR U1719 ( .A(n2365), .B(n2366), .Z(n2364) );
  AND U1720 ( .A(n2367), .B(n2368), .Z(n2366) );
  AND U1721 ( .A(n2168), .B(n2369), .Z(n2365) );
  XOR U1722 ( .A(n2370), .B(n2371), .Z(n2363) );
  AND U1723 ( .A(n2169), .B(n2372), .Z(n2371) );
  AND U1724 ( .A(n2373), .B(n2167), .Z(n2370) );
  XNOR U1725 ( .A(n2374), .B(n2375), .Z(n2155) );
  XOR U1726 ( .A(n2376), .B(n2377), .Z(n2153) );
  XOR U1727 ( .A(n2378), .B(n2379), .Z(n2377) );
  AND U1728 ( .A(n2379), .B(n2380), .Z(n2378) );
  XOR U1729 ( .A(n2381), .B(n2382), .Z(n2376) );
  AND U1730 ( .A(n2383), .B(n2374), .Z(n2382) );
  AND U1731 ( .A(n2384), .B(n2385), .Z(n2381) );
  XOR U1732 ( .A(n2386), .B(n2387), .Z(n2146) );
  XOR U1733 ( .A(n2388), .B(n2389), .Z(n2144) );
  XOR U1734 ( .A(n2390), .B(n2391), .Z(n2389) );
  AND U1735 ( .A(n2392), .B(n2391), .Z(n2390) );
  XOR U1736 ( .A(n2393), .B(n2394), .Z(n2388) );
  NOR U1737 ( .A(n2395), .B(n2386), .Z(n2394) );
  NOR U1738 ( .A(n2396), .B(n2387), .Z(n2393) );
  XOR U1739 ( .A(n2397), .B(n2398), .Z(n2137) );
  XOR U1740 ( .A(n2399), .B(n2400), .Z(n2135) );
  XNOR U1741 ( .A(n2401), .B(n2402), .Z(n2400) );
  NOR U1742 ( .A(n2403), .B(n2402), .Z(n2401) );
  XOR U1743 ( .A(n2404), .B(n2405), .Z(n2399) );
  NOR U1744 ( .A(n2406), .B(n2397), .Z(n2405) );
  NOR U1745 ( .A(n2407), .B(n2398), .Z(n2404) );
  XNOR U1746 ( .A(n2132), .B(n2130), .Z(n2133) );
  XNOR U1747 ( .A(n2408), .B(n2409), .Z(n1097) );
  NOR U1748 ( .A(n2410), .B(n2408), .Z(n2409) );
  XOR U1749 ( .A(n2411), .B(n2412), .Z(n1088) );
  NOR U1750 ( .A(n2413), .B(n2411), .Z(n2412) );
  XOR U1751 ( .A(n2414), .B(n2415), .Z(n1089) );
  NOR U1752 ( .A(n2416), .B(n2414), .Z(n2415) );
  XOR U1753 ( .A(n2417), .B(n2418), .Z(n1086) );
  NOR U1754 ( .A(n2419), .B(n2417), .Z(n2418) );
  XOR U1755 ( .A(n2420), .B(n2421), .Z(n1076) );
  NOR U1756 ( .A(n2422), .B(n2420), .Z(n2421) );
  XOR U1757 ( .A(n2423), .B(n2424), .Z(n1107) );
  NOR U1758 ( .A(n2425), .B(n2423), .Z(n2424) );
  XOR U1759 ( .A(n2426), .B(n2427), .Z(n1104) );
  NOR U1760 ( .A(n2428), .B(n2426), .Z(n2427) );
  XOR U1761 ( .A(n2429), .B(n2430), .Z(n1080) );
  NOR U1762 ( .A(n2431), .B(n2429), .Z(n2430) );
  XOR U1763 ( .A(n2432), .B(n2433), .Z(n1124) );
  NOR U1764 ( .A(n2434), .B(n2432), .Z(n2433) );
  XOR U1765 ( .A(n2435), .B(n2436), .Z(n1119) );
  NOR U1766 ( .A(n2437), .B(n2435), .Z(n2436) );
  XOR U1767 ( .A(n2438), .B(n2439), .Z(n1120) );
  NOR U1768 ( .A(n2440), .B(n2438), .Z(n2439) );
  XOR U1769 ( .A(n2441), .B(n2442), .Z(n1077) );
  NOR U1770 ( .A(n2443), .B(n2441), .Z(n2442) );
  XOR U1771 ( .A(n2444), .B(n2445), .Z(n1135) );
  NOR U1772 ( .A(n2446), .B(n2444), .Z(n2445) );
  XOR U1773 ( .A(n2447), .B(n2448), .Z(n1130) );
  NOR U1774 ( .A(n2449), .B(n2447), .Z(n2448) );
  XOR U1775 ( .A(n2450), .B(n2451), .Z(n1131) );
  NOR U1776 ( .A(n2452), .B(n2450), .Z(n2451) );
  XOR U1777 ( .A(n2453), .B(n2454), .Z(n1070) );
  NOR U1778 ( .A(n2455), .B(n2453), .Z(n2454) );
  XOR U1779 ( .A(n2456), .B(n2457), .Z(n1146) );
  NOR U1780 ( .A(n2458), .B(n2456), .Z(n2457) );
  XOR U1781 ( .A(n2459), .B(n2460), .Z(n1141) );
  NOR U1782 ( .A(n2461), .B(n2459), .Z(n2460) );
  XOR U1783 ( .A(n2462), .B(n2463), .Z(n1142) );
  NOR U1784 ( .A(n2464), .B(n2462), .Z(n2463) );
  XOR U1785 ( .A(n2465), .B(n2466), .Z(n1061) );
  NOR U1786 ( .A(n2467), .B(n2465), .Z(n2466) );
  XOR U1787 ( .A(n2468), .B(n2469), .Z(n1157) );
  NOR U1788 ( .A(n2470), .B(n2468), .Z(n2469) );
  XOR U1789 ( .A(n2471), .B(n2472), .Z(n1152) );
  NOR U1790 ( .A(n2473), .B(n2471), .Z(n2472) );
  XOR U1791 ( .A(n2474), .B(n2475), .Z(n1153) );
  NOR U1792 ( .A(n2476), .B(n2474), .Z(n2475) );
  XOR U1793 ( .A(n2477), .B(n2478), .Z(n1052) );
  NOR U1794 ( .A(n2479), .B(n2477), .Z(n2478) );
  XOR U1795 ( .A(n2480), .B(n2481), .Z(n1168) );
  NOR U1796 ( .A(n2482), .B(n2480), .Z(n2481) );
  XOR U1797 ( .A(n2483), .B(n2484), .Z(n1163) );
  NOR U1798 ( .A(n2485), .B(n2483), .Z(n2484) );
  XOR U1799 ( .A(n2486), .B(n2487), .Z(n1164) );
  NOR U1800 ( .A(n2488), .B(n2486), .Z(n2487) );
  XOR U1801 ( .A(n2489), .B(n2490), .Z(n1043) );
  NOR U1802 ( .A(n2491), .B(n2489), .Z(n2490) );
  XOR U1803 ( .A(n2492), .B(n2493), .Z(n1179) );
  NOR U1804 ( .A(n2494), .B(n2492), .Z(n2493) );
  XOR U1805 ( .A(n2495), .B(n2496), .Z(n1174) );
  NOR U1806 ( .A(n2497), .B(n2495), .Z(n2496) );
  XOR U1807 ( .A(n2498), .B(n2499), .Z(n1175) );
  NOR U1808 ( .A(n2500), .B(n2498), .Z(n2499) );
  XOR U1809 ( .A(n2501), .B(n2502), .Z(n1034) );
  NOR U1810 ( .A(n2503), .B(n2501), .Z(n2502) );
  XOR U1811 ( .A(n2504), .B(n2505), .Z(n1190) );
  NOR U1812 ( .A(n2506), .B(n2504), .Z(n2505) );
  XOR U1813 ( .A(n2507), .B(n2508), .Z(n1185) );
  NOR U1814 ( .A(n2509), .B(n2507), .Z(n2508) );
  XOR U1815 ( .A(n2510), .B(n2511), .Z(n1186) );
  NOR U1816 ( .A(n2512), .B(n2510), .Z(n2511) );
  XOR U1817 ( .A(n2513), .B(n2514), .Z(n1025) );
  NOR U1818 ( .A(n2515), .B(n2513), .Z(n2514) );
  XOR U1819 ( .A(n2516), .B(n2517), .Z(n1201) );
  NOR U1820 ( .A(n2518), .B(n2516), .Z(n2517) );
  XOR U1821 ( .A(n2519), .B(n2520), .Z(n1196) );
  NOR U1822 ( .A(n2521), .B(n2519), .Z(n2520) );
  XOR U1823 ( .A(n2522), .B(n2523), .Z(n1197) );
  NOR U1824 ( .A(n2524), .B(n2522), .Z(n2523) );
  XOR U1825 ( .A(n2525), .B(n2526), .Z(n1016) );
  NOR U1826 ( .A(n2527), .B(n2525), .Z(n2526) );
  XOR U1827 ( .A(n2528), .B(n2529), .Z(n1212) );
  NOR U1828 ( .A(n2530), .B(n2528), .Z(n2529) );
  XOR U1829 ( .A(n2531), .B(n2532), .Z(n1207) );
  NOR U1830 ( .A(n2533), .B(n2531), .Z(n2532) );
  XOR U1831 ( .A(n2534), .B(n2535), .Z(n1208) );
  NOR U1832 ( .A(n2536), .B(n2534), .Z(n2535) );
  XOR U1833 ( .A(n2537), .B(n2538), .Z(n1007) );
  NOR U1834 ( .A(n2539), .B(n2537), .Z(n2538) );
  XOR U1835 ( .A(n2540), .B(n2541), .Z(n1223) );
  NOR U1836 ( .A(n2542), .B(n2540), .Z(n2541) );
  XOR U1837 ( .A(n2543), .B(n2544), .Z(n1218) );
  NOR U1838 ( .A(n2545), .B(n2543), .Z(n2544) );
  XOR U1839 ( .A(n2546), .B(n2547), .Z(n1219) );
  NOR U1840 ( .A(n2548), .B(n2546), .Z(n2547) );
  XOR U1841 ( .A(n2549), .B(n2550), .Z(n998) );
  NOR U1842 ( .A(n2551), .B(n2549), .Z(n2550) );
  XOR U1843 ( .A(n2552), .B(n2553), .Z(n1234) );
  NOR U1844 ( .A(n2554), .B(n2552), .Z(n2553) );
  XOR U1845 ( .A(n2555), .B(n2556), .Z(n1229) );
  NOR U1846 ( .A(n2557), .B(n2555), .Z(n2556) );
  XOR U1847 ( .A(n2558), .B(n2559), .Z(n1230) );
  NOR U1848 ( .A(n2560), .B(n2558), .Z(n2559) );
  XOR U1849 ( .A(n2561), .B(n2562), .Z(n989) );
  NOR U1850 ( .A(n2563), .B(n2561), .Z(n2562) );
  XOR U1851 ( .A(n2564), .B(n2565), .Z(n1245) );
  NOR U1852 ( .A(n2566), .B(n2564), .Z(n2565) );
  XOR U1853 ( .A(n2567), .B(n2568), .Z(n1240) );
  NOR U1854 ( .A(n2569), .B(n2567), .Z(n2568) );
  XOR U1855 ( .A(n2570), .B(n2571), .Z(n1241) );
  NOR U1856 ( .A(n2572), .B(n2570), .Z(n2571) );
  XOR U1857 ( .A(n2573), .B(n2574), .Z(n980) );
  NOR U1858 ( .A(n2575), .B(n2573), .Z(n2574) );
  XOR U1859 ( .A(n2576), .B(n2577), .Z(n1256) );
  NOR U1860 ( .A(n2578), .B(n2576), .Z(n2577) );
  XOR U1861 ( .A(n2579), .B(n2580), .Z(n1251) );
  NOR U1862 ( .A(n2581), .B(n2579), .Z(n2580) );
  XOR U1863 ( .A(n2582), .B(n2583), .Z(n1252) );
  NOR U1864 ( .A(n2584), .B(n2582), .Z(n2583) );
  XOR U1865 ( .A(n2585), .B(n2586), .Z(n971) );
  NOR U1866 ( .A(n2587), .B(n2585), .Z(n2586) );
  XOR U1867 ( .A(n2588), .B(n2589), .Z(n1267) );
  NOR U1868 ( .A(n2590), .B(n2588), .Z(n2589) );
  XOR U1869 ( .A(n2591), .B(n2592), .Z(n1262) );
  NOR U1870 ( .A(n2593), .B(n2591), .Z(n2592) );
  XOR U1871 ( .A(n2594), .B(n2595), .Z(n1263) );
  NOR U1872 ( .A(n2596), .B(n2594), .Z(n2595) );
  XOR U1873 ( .A(n2597), .B(n2598), .Z(n962) );
  NOR U1874 ( .A(n2599), .B(n2597), .Z(n2598) );
  XOR U1875 ( .A(n2600), .B(n2601), .Z(n1278) );
  NOR U1876 ( .A(n2602), .B(n2600), .Z(n2601) );
  XOR U1877 ( .A(n2603), .B(n2604), .Z(n1273) );
  NOR U1878 ( .A(n2605), .B(n2603), .Z(n2604) );
  XOR U1879 ( .A(n2606), .B(n2607), .Z(n1274) );
  NOR U1880 ( .A(n2608), .B(n2606), .Z(n2607) );
  XOR U1881 ( .A(n2609), .B(n2610), .Z(n953) );
  NOR U1882 ( .A(n2611), .B(n2609), .Z(n2610) );
  XOR U1883 ( .A(n2612), .B(n2613), .Z(n1289) );
  NOR U1884 ( .A(n2614), .B(n2612), .Z(n2613) );
  XOR U1885 ( .A(n2615), .B(n2616), .Z(n1284) );
  NOR U1886 ( .A(n2617), .B(n2615), .Z(n2616) );
  XOR U1887 ( .A(n2618), .B(n2619), .Z(n1285) );
  NOR U1888 ( .A(n2620), .B(n2618), .Z(n2619) );
  XOR U1889 ( .A(n2621), .B(n2622), .Z(n944) );
  NOR U1890 ( .A(n2623), .B(n2621), .Z(n2622) );
  XOR U1891 ( .A(n2624), .B(n2625), .Z(n1300) );
  NOR U1892 ( .A(n2626), .B(n2624), .Z(n2625) );
  XOR U1893 ( .A(n2627), .B(n2628), .Z(n1295) );
  NOR U1894 ( .A(n2629), .B(n2627), .Z(n2628) );
  XOR U1895 ( .A(n2630), .B(n2631), .Z(n1296) );
  NOR U1896 ( .A(n2632), .B(n2630), .Z(n2631) );
  XOR U1897 ( .A(n2633), .B(n2634), .Z(n935) );
  NOR U1898 ( .A(n2635), .B(n2633), .Z(n2634) );
  XOR U1899 ( .A(n2636), .B(n2637), .Z(n1311) );
  NOR U1900 ( .A(n2638), .B(n2636), .Z(n2637) );
  XOR U1901 ( .A(n2639), .B(n2640), .Z(n1306) );
  NOR U1902 ( .A(n2641), .B(n2639), .Z(n2640) );
  XOR U1903 ( .A(n2642), .B(n2643), .Z(n1307) );
  NOR U1904 ( .A(n2644), .B(n2642), .Z(n2643) );
  XOR U1905 ( .A(n2645), .B(n2646), .Z(n926) );
  NOR U1906 ( .A(n2647), .B(n2645), .Z(n2646) );
  XOR U1907 ( .A(n2648), .B(n2649), .Z(n1322) );
  NOR U1908 ( .A(n2650), .B(n2648), .Z(n2649) );
  XOR U1909 ( .A(n2651), .B(n2652), .Z(n1317) );
  NOR U1910 ( .A(n2653), .B(n2651), .Z(n2652) );
  XOR U1911 ( .A(n2654), .B(n2655), .Z(n1318) );
  NOR U1912 ( .A(n2656), .B(n2654), .Z(n2655) );
  XOR U1913 ( .A(n2657), .B(n2658), .Z(n917) );
  NOR U1914 ( .A(n2659), .B(n2657), .Z(n2658) );
  XOR U1915 ( .A(n2660), .B(n2661), .Z(n1333) );
  NOR U1916 ( .A(n2662), .B(n2660), .Z(n2661) );
  XOR U1917 ( .A(n2663), .B(n2664), .Z(n1328) );
  NOR U1918 ( .A(n2665), .B(n2663), .Z(n2664) );
  XOR U1919 ( .A(n2666), .B(n2667), .Z(n1329) );
  NOR U1920 ( .A(n2668), .B(n2666), .Z(n2667) );
  XOR U1921 ( .A(n2669), .B(n2670), .Z(n908) );
  NOR U1922 ( .A(n2671), .B(n2669), .Z(n2670) );
  XOR U1923 ( .A(n2672), .B(n2673), .Z(n1344) );
  NOR U1924 ( .A(n2674), .B(n2672), .Z(n2673) );
  XOR U1925 ( .A(n2675), .B(n2676), .Z(n1339) );
  NOR U1926 ( .A(n2677), .B(n2675), .Z(n2676) );
  XOR U1927 ( .A(n2678), .B(n2679), .Z(n1340) );
  NOR U1928 ( .A(n2680), .B(n2678), .Z(n2679) );
  XOR U1929 ( .A(n2681), .B(n2682), .Z(n899) );
  NOR U1930 ( .A(n2683), .B(n2681), .Z(n2682) );
  XOR U1931 ( .A(n2684), .B(n2685), .Z(n1355) );
  NOR U1932 ( .A(n2686), .B(n2684), .Z(n2685) );
  XOR U1933 ( .A(n2687), .B(n2688), .Z(n1350) );
  NOR U1934 ( .A(n2689), .B(n2687), .Z(n2688) );
  XOR U1935 ( .A(n2690), .B(n2691), .Z(n1351) );
  NOR U1936 ( .A(n2692), .B(n2690), .Z(n2691) );
  XOR U1937 ( .A(n2693), .B(n2694), .Z(n890) );
  NOR U1938 ( .A(n2695), .B(n2693), .Z(n2694) );
  XOR U1939 ( .A(n2696), .B(n2697), .Z(n1366) );
  NOR U1940 ( .A(n2698), .B(n2696), .Z(n2697) );
  XOR U1941 ( .A(n2699), .B(n2700), .Z(n1361) );
  NOR U1942 ( .A(n2701), .B(n2699), .Z(n2700) );
  XOR U1943 ( .A(n2702), .B(n2703), .Z(n1362) );
  NOR U1944 ( .A(n2704), .B(n2702), .Z(n2703) );
  XOR U1945 ( .A(n2705), .B(n2706), .Z(n881) );
  NOR U1946 ( .A(n2707), .B(n2705), .Z(n2706) );
  XOR U1947 ( .A(n2708), .B(n2709), .Z(n1377) );
  NOR U1948 ( .A(n2710), .B(n2708), .Z(n2709) );
  XOR U1949 ( .A(n2711), .B(n2712), .Z(n1372) );
  NOR U1950 ( .A(n2713), .B(n2711), .Z(n2712) );
  XOR U1951 ( .A(n2714), .B(n2715), .Z(n1373) );
  NOR U1952 ( .A(n2716), .B(n2714), .Z(n2715) );
  XOR U1953 ( .A(n2717), .B(n2718), .Z(n872) );
  NOR U1954 ( .A(n2719), .B(n2717), .Z(n2718) );
  XOR U1955 ( .A(n2720), .B(n2721), .Z(n1388) );
  NOR U1956 ( .A(n2722), .B(n2720), .Z(n2721) );
  XOR U1957 ( .A(n2723), .B(n2724), .Z(n1383) );
  NOR U1958 ( .A(n2725), .B(n2723), .Z(n2724) );
  XOR U1959 ( .A(n2726), .B(n2727), .Z(n1384) );
  NOR U1960 ( .A(n2728), .B(n2726), .Z(n2727) );
  XOR U1961 ( .A(n2729), .B(n2730), .Z(n863) );
  NOR U1962 ( .A(n2731), .B(n2729), .Z(n2730) );
  XOR U1963 ( .A(n2732), .B(n2733), .Z(n1399) );
  NOR U1964 ( .A(n2734), .B(n2732), .Z(n2733) );
  XOR U1965 ( .A(n2735), .B(n2736), .Z(n1394) );
  NOR U1966 ( .A(n2737), .B(n2735), .Z(n2736) );
  XOR U1967 ( .A(n2738), .B(n2739), .Z(n1395) );
  NOR U1968 ( .A(n2740), .B(n2738), .Z(n2739) );
  XOR U1969 ( .A(n2741), .B(n2742), .Z(n854) );
  NOR U1970 ( .A(n2743), .B(n2741), .Z(n2742) );
  XOR U1971 ( .A(n2744), .B(n2745), .Z(n1410) );
  NOR U1972 ( .A(n2746), .B(n2744), .Z(n2745) );
  XOR U1973 ( .A(n2747), .B(n2748), .Z(n1405) );
  NOR U1974 ( .A(n2749), .B(n2747), .Z(n2748) );
  XOR U1975 ( .A(n2750), .B(n2751), .Z(n1406) );
  NOR U1976 ( .A(n2752), .B(n2750), .Z(n2751) );
  XOR U1977 ( .A(n2753), .B(n2754), .Z(n845) );
  NOR U1978 ( .A(n2755), .B(n2753), .Z(n2754) );
  XOR U1979 ( .A(n2756), .B(n2757), .Z(n1421) );
  NOR U1980 ( .A(n2758), .B(n2756), .Z(n2757) );
  XOR U1981 ( .A(n2759), .B(n2760), .Z(n1416) );
  NOR U1982 ( .A(n2761), .B(n2759), .Z(n2760) );
  XOR U1983 ( .A(n2762), .B(n2763), .Z(n1417) );
  NOR U1984 ( .A(n2764), .B(n2762), .Z(n2763) );
  XOR U1985 ( .A(n2765), .B(n2766), .Z(n836) );
  NOR U1986 ( .A(n2767), .B(n2765), .Z(n2766) );
  XOR U1987 ( .A(n2768), .B(n2769), .Z(n1432) );
  NOR U1988 ( .A(n2770), .B(n2768), .Z(n2769) );
  XOR U1989 ( .A(n2771), .B(n2772), .Z(n1427) );
  NOR U1990 ( .A(n2773), .B(n2771), .Z(n2772) );
  XOR U1991 ( .A(n2774), .B(n2775), .Z(n1428) );
  NOR U1992 ( .A(n2776), .B(n2774), .Z(n2775) );
  XOR U1993 ( .A(n2777), .B(n2778), .Z(n827) );
  NOR U1994 ( .A(n2779), .B(n2777), .Z(n2778) );
  XOR U1995 ( .A(n2780), .B(n2781), .Z(n801) );
  NOR U1996 ( .A(n2782), .B(n2780), .Z(n2781) );
  XOR U1997 ( .A(n2783), .B(n2784), .Z(n806) );
  NOR U1998 ( .A(n2785), .B(n2783), .Z(n2784) );
  IV U1999 ( .A(n808), .Z(n2119) );
  XNOR U2000 ( .A(n2786), .B(n2787), .Z(n808) );
  NOR U2001 ( .A(n2788), .B(n2786), .Z(n2787) );
  XOR U2002 ( .A(n2789), .B(n2790), .Z(n818) );
  NOR U2003 ( .A(n2791), .B(n2789), .Z(n2790) );
  XNOR U2004 ( .A(n2792), .B(n2793), .Z(n1438) );
  NOR U2005 ( .A(n56), .B(n2794), .Z(n2793) );
  IV U2006 ( .A(n2792), .Z(n2794) );
  XOR U2007 ( .A(n2795), .B(n2796), .Z(n1440) );
  AND U2008 ( .A(n2797), .B(n2798), .Z(n2796) );
  XOR U2009 ( .A(n2795), .B(n58), .Z(n2798) );
  XOR U2010 ( .A(n2117), .B(n2116), .Z(n58) );
  XNOR U2011 ( .A(n2114), .B(n2113), .Z(n2116) );
  XNOR U2012 ( .A(n2111), .B(n2110), .Z(n2113) );
  XNOR U2013 ( .A(n2108), .B(n2107), .Z(n2110) );
  XNOR U2014 ( .A(n2105), .B(n2104), .Z(n2107) );
  XNOR U2015 ( .A(n2102), .B(n2101), .Z(n2104) );
  XNOR U2016 ( .A(n2099), .B(n2098), .Z(n2101) );
  XNOR U2017 ( .A(n2096), .B(n2095), .Z(n2098) );
  XNOR U2018 ( .A(n2093), .B(n2092), .Z(n2095) );
  XNOR U2019 ( .A(n2090), .B(n2089), .Z(n2092) );
  XNOR U2020 ( .A(n2087), .B(n2086), .Z(n2089) );
  XNOR U2021 ( .A(n2084), .B(n2083), .Z(n2086) );
  XNOR U2022 ( .A(n2081), .B(n2080), .Z(n2083) );
  XNOR U2023 ( .A(n2078), .B(n2077), .Z(n2080) );
  XNOR U2024 ( .A(n2075), .B(n2074), .Z(n2077) );
  XNOR U2025 ( .A(n2072), .B(n2071), .Z(n2074) );
  XNOR U2026 ( .A(n2069), .B(n2068), .Z(n2071) );
  XNOR U2027 ( .A(n2066), .B(n2065), .Z(n2068) );
  XNOR U2028 ( .A(n2063), .B(n2062), .Z(n2065) );
  XNOR U2029 ( .A(n2060), .B(n2059), .Z(n2062) );
  XNOR U2030 ( .A(n2057), .B(n2056), .Z(n2059) );
  XNOR U2031 ( .A(n2054), .B(n2053), .Z(n2056) );
  XNOR U2032 ( .A(n2051), .B(n2050), .Z(n2053) );
  XNOR U2033 ( .A(n2048), .B(n2047), .Z(n2050) );
  XNOR U2034 ( .A(n2045), .B(n2044), .Z(n2047) );
  XNOR U2035 ( .A(n2042), .B(n2041), .Z(n2044) );
  XNOR U2036 ( .A(n2039), .B(n2038), .Z(n2041) );
  XNOR U2037 ( .A(n2036), .B(n2035), .Z(n2038) );
  XNOR U2038 ( .A(n2033), .B(n2032), .Z(n2035) );
  XNOR U2039 ( .A(n2030), .B(n2029), .Z(n2032) );
  XNOR U2040 ( .A(n2027), .B(n2026), .Z(n2029) );
  XNOR U2041 ( .A(n2024), .B(n2023), .Z(n2026) );
  XNOR U2042 ( .A(n2021), .B(n2020), .Z(n2023) );
  XNOR U2043 ( .A(n2018), .B(n2017), .Z(n2020) );
  XNOR U2044 ( .A(n2015), .B(n2014), .Z(n2017) );
  XNOR U2045 ( .A(n2012), .B(n2011), .Z(n2014) );
  XNOR U2046 ( .A(n2009), .B(n2008), .Z(n2011) );
  XNOR U2047 ( .A(n2006), .B(n2005), .Z(n2008) );
  XNOR U2048 ( .A(n2003), .B(n2002), .Z(n2005) );
  XNOR U2049 ( .A(n2000), .B(n1999), .Z(n2002) );
  XNOR U2050 ( .A(n1997), .B(n1996), .Z(n1999) );
  XNOR U2051 ( .A(n1994), .B(n1993), .Z(n1996) );
  XNOR U2052 ( .A(n1991), .B(n1990), .Z(n1993) );
  XNOR U2053 ( .A(n1988), .B(n1987), .Z(n1990) );
  XNOR U2054 ( .A(n1985), .B(n1984), .Z(n1987) );
  XNOR U2055 ( .A(n1982), .B(n1981), .Z(n1984) );
  XNOR U2056 ( .A(n1979), .B(n1978), .Z(n1981) );
  XNOR U2057 ( .A(n1976), .B(n1975), .Z(n1978) );
  XNOR U2058 ( .A(n1973), .B(n1972), .Z(n1975) );
  XNOR U2059 ( .A(n1970), .B(n1969), .Z(n1972) );
  XNOR U2060 ( .A(n1967), .B(n1966), .Z(n1969) );
  XNOR U2061 ( .A(n1964), .B(n1963), .Z(n1966) );
  XNOR U2062 ( .A(n1961), .B(n1960), .Z(n1963) );
  XNOR U2063 ( .A(n1958), .B(n1957), .Z(n1960) );
  XNOR U2064 ( .A(n1955), .B(n1954), .Z(n1957) );
  XNOR U2065 ( .A(n1952), .B(n1951), .Z(n1954) );
  XNOR U2066 ( .A(n1949), .B(n1948), .Z(n1951) );
  XNOR U2067 ( .A(n1946), .B(n1945), .Z(n1948) );
  XNOR U2068 ( .A(n1943), .B(n1942), .Z(n1945) );
  XNOR U2069 ( .A(n1940), .B(n1939), .Z(n1942) );
  XNOR U2070 ( .A(n1937), .B(n1936), .Z(n1939) );
  XNOR U2071 ( .A(n1934), .B(n1933), .Z(n1936) );
  XNOR U2072 ( .A(n1931), .B(n1930), .Z(n1933) );
  XNOR U2073 ( .A(n1928), .B(n1927), .Z(n1930) );
  XNOR U2074 ( .A(n1925), .B(n1924), .Z(n1927) );
  XNOR U2075 ( .A(n1922), .B(n1921), .Z(n1924) );
  XNOR U2076 ( .A(n1919), .B(n1918), .Z(n1921) );
  XNOR U2077 ( .A(n1916), .B(n1915), .Z(n1918) );
  XNOR U2078 ( .A(n1913), .B(n1912), .Z(n1915) );
  XNOR U2079 ( .A(n1910), .B(n1909), .Z(n1912) );
  XNOR U2080 ( .A(n1907), .B(n1906), .Z(n1909) );
  XNOR U2081 ( .A(n1904), .B(n1903), .Z(n1906) );
  XNOR U2082 ( .A(n1901), .B(n1900), .Z(n1903) );
  XNOR U2083 ( .A(n1898), .B(n1897), .Z(n1900) );
  XNOR U2084 ( .A(n1895), .B(n1894), .Z(n1897) );
  XNOR U2085 ( .A(n1892), .B(n1891), .Z(n1894) );
  XNOR U2086 ( .A(n1889), .B(n1888), .Z(n1891) );
  XNOR U2087 ( .A(n1886), .B(n1885), .Z(n1888) );
  XNOR U2088 ( .A(n1883), .B(n1882), .Z(n1885) );
  XNOR U2089 ( .A(n1880), .B(n1879), .Z(n1882) );
  XNOR U2090 ( .A(n1877), .B(n1876), .Z(n1879) );
  XNOR U2091 ( .A(n1874), .B(n1873), .Z(n1876) );
  XNOR U2092 ( .A(n1871), .B(n1870), .Z(n1873) );
  XNOR U2093 ( .A(n1868), .B(n1867), .Z(n1870) );
  XNOR U2094 ( .A(n1865), .B(n1864), .Z(n1867) );
  XNOR U2095 ( .A(n1862), .B(n1861), .Z(n1864) );
  XNOR U2096 ( .A(n1859), .B(n1858), .Z(n1861) );
  XNOR U2097 ( .A(n1856), .B(n1855), .Z(n1858) );
  XNOR U2098 ( .A(n1853), .B(n1852), .Z(n1855) );
  XNOR U2099 ( .A(n1850), .B(n1849), .Z(n1852) );
  XNOR U2100 ( .A(n1847), .B(n1846), .Z(n1849) );
  XNOR U2101 ( .A(n1844), .B(n1843), .Z(n1846) );
  XNOR U2102 ( .A(n1841), .B(n1840), .Z(n1843) );
  XNOR U2103 ( .A(n1838), .B(n1837), .Z(n1840) );
  XNOR U2104 ( .A(n1835), .B(n1834), .Z(n1837) );
  XNOR U2105 ( .A(n1832), .B(n1831), .Z(n1834) );
  XNOR U2106 ( .A(n1829), .B(n1828), .Z(n1831) );
  XNOR U2107 ( .A(n1826), .B(n1825), .Z(n1828) );
  XNOR U2108 ( .A(n1823), .B(n1822), .Z(n1825) );
  XNOR U2109 ( .A(n1820), .B(n1819), .Z(n1822) );
  XNOR U2110 ( .A(n1817), .B(n1816), .Z(n1819) );
  XNOR U2111 ( .A(n1814), .B(n1813), .Z(n1816) );
  XNOR U2112 ( .A(n1811), .B(n1810), .Z(n1813) );
  XNOR U2113 ( .A(n1808), .B(n1807), .Z(n1810) );
  XNOR U2114 ( .A(n1805), .B(n1804), .Z(n1807) );
  XNOR U2115 ( .A(n1802), .B(n1801), .Z(n1804) );
  XNOR U2116 ( .A(n1799), .B(n1798), .Z(n1801) );
  XNOR U2117 ( .A(n1796), .B(n1795), .Z(n1798) );
  XNOR U2118 ( .A(n1793), .B(n1792), .Z(n1795) );
  XNOR U2119 ( .A(n1790), .B(n1789), .Z(n1792) );
  XNOR U2120 ( .A(n1787), .B(n1786), .Z(n1789) );
  XNOR U2121 ( .A(n1784), .B(n1783), .Z(n1786) );
  XNOR U2122 ( .A(n1781), .B(n1780), .Z(n1783) );
  XNOR U2123 ( .A(n1778), .B(n1777), .Z(n1780) );
  XNOR U2124 ( .A(n1775), .B(n1774), .Z(n1777) );
  XNOR U2125 ( .A(n1772), .B(n1771), .Z(n1774) );
  XNOR U2126 ( .A(n1769), .B(n1768), .Z(n1771) );
  XNOR U2127 ( .A(n1766), .B(n1765), .Z(n1768) );
  XNOR U2128 ( .A(n1763), .B(n1762), .Z(n1765) );
  XNOR U2129 ( .A(n1760), .B(n1759), .Z(n1762) );
  XNOR U2130 ( .A(n1757), .B(n1756), .Z(n1759) );
  XNOR U2131 ( .A(n1754), .B(n1753), .Z(n1756) );
  XNOR U2132 ( .A(n1751), .B(n1750), .Z(n1753) );
  XNOR U2133 ( .A(n1748), .B(n1747), .Z(n1750) );
  XNOR U2134 ( .A(n1745), .B(n1744), .Z(n1747) );
  XNOR U2135 ( .A(n1742), .B(n1741), .Z(n1744) );
  XNOR U2136 ( .A(n1739), .B(n1738), .Z(n1741) );
  XNOR U2137 ( .A(n1736), .B(n1735), .Z(n1738) );
  XNOR U2138 ( .A(n1733), .B(n1731), .Z(n1735) );
  XNOR U2139 ( .A(n1732), .B(n1453), .Z(n1731) );
  XNOR U2140 ( .A(n1454), .B(n1451), .Z(n1453) );
  XNOR U2141 ( .A(n1452), .B(n1455), .Z(n1451) );
  XNOR U2142 ( .A(n1456), .B(n1726), .Z(n1455) );
  XNOR U2143 ( .A(n1463), .B(n1725), .Z(n1726) );
  XNOR U2144 ( .A(n1718), .B(n1722), .Z(n1725) );
  XNOR U2145 ( .A(n1717), .B(n1715), .Z(n1722) );
  XNOR U2146 ( .A(n1716), .B(n1714), .Z(n1715) );
  XNOR U2147 ( .A(n1470), .B(n1709), .Z(n1714) );
  XOR U2148 ( .A(n1469), .B(n1707), .Z(n1709) );
  XNOR U2149 ( .A(n1708), .B(n1703), .Z(n1707) );
  XOR U2150 ( .A(n1704), .B(n1485), .Z(n1703) );
  XOR U2151 ( .A(n1486), .B(n1702), .Z(n1485) );
  XOR U2152 ( .A(n1479), .B(n1697), .Z(n1702) );
  XOR U2153 ( .A(n1481), .B(n1696), .Z(n1697) );
  XOR U2154 ( .A(n1693), .B(n1484), .Z(n1696) );
  AND U2155 ( .A(n2799), .B(n2800), .Z(n1484) );
  XOR U2156 ( .A(n1692), .B(n1683), .Z(n1693) );
  AND U2157 ( .A(n2801), .B(n2802), .Z(n1683) );
  XOR U2158 ( .A(n1689), .B(n1682), .Z(n1692) );
  AND U2159 ( .A(n2803), .B(n2804), .Z(n1682) );
  XOR U2160 ( .A(n1688), .B(n1681), .Z(n1689) );
  AND U2161 ( .A(n2805), .B(n2806), .Z(n1681) );
  XNOR U2162 ( .A(n1650), .B(n1680), .Z(n1688) );
  AND U2163 ( .A(n2807), .B(n2808), .Z(n1680) );
  XNOR U2164 ( .A(n1675), .B(n1651), .Z(n1650) );
  AND U2165 ( .A(n2809), .B(n2810), .Z(n1651) );
  XOR U2166 ( .A(n1674), .B(n1648), .Z(n1675) );
  AND U2167 ( .A(n2811), .B(n2812), .Z(n1648) );
  XOR U2168 ( .A(n1679), .B(n1655), .Z(n1674) );
  AND U2169 ( .A(n2813), .B(n2814), .Z(n1655) );
  XNOR U2170 ( .A(n1662), .B(n1654), .Z(n1679) );
  AND U2171 ( .A(n2815), .B(n2816), .Z(n1654) );
  XNOR U2172 ( .A(n1671), .B(n1663), .Z(n1662) );
  AND U2173 ( .A(n2817), .B(n2818), .Z(n1663) );
  XOR U2174 ( .A(n1670), .B(n1660), .Z(n1671) );
  AND U2175 ( .A(n2819), .B(n2820), .Z(n1660) );
  XOR U2176 ( .A(n1678), .B(n1659), .Z(n1670) );
  AND U2177 ( .A(n2821), .B(n2822), .Z(n1659) );
  XNOR U2178 ( .A(n1615), .B(n1658), .Z(n1678) );
  AND U2179 ( .A(n2823), .B(n2824), .Z(n1658) );
  XNOR U2180 ( .A(n1643), .B(n1616), .Z(n1615) );
  AND U2181 ( .A(n2825), .B(n2826), .Z(n1616) );
  XOR U2182 ( .A(n1642), .B(n1613), .Z(n1643) );
  AND U2183 ( .A(n2827), .B(n2828), .Z(n1613) );
  XOR U2184 ( .A(n1647), .B(n1612), .Z(n1642) );
  AND U2185 ( .A(n2829), .B(n2830), .Z(n1612) );
  XNOR U2186 ( .A(n1625), .B(n1611), .Z(n1647) );
  AND U2187 ( .A(n2831), .B(n2832), .Z(n1611) );
  XNOR U2188 ( .A(n1639), .B(n1626), .Z(n1625) );
  AND U2189 ( .A(n2833), .B(n2834), .Z(n1626) );
  XOR U2190 ( .A(n1638), .B(n1623), .Z(n1639) );
  AND U2191 ( .A(n2835), .B(n2836), .Z(n1623) );
  XOR U2192 ( .A(n1646), .B(n1622), .Z(n1638) );
  AND U2193 ( .A(n2837), .B(n2838), .Z(n1622) );
  XNOR U2194 ( .A(n1630), .B(n1621), .Z(n1646) );
  AND U2195 ( .A(n2839), .B(n2840), .Z(n1621) );
  XNOR U2196 ( .A(n1603), .B(n1631), .Z(n1630) );
  AND U2197 ( .A(n2841), .B(n2842), .Z(n1631) );
  XOR U2198 ( .A(n1601), .B(n1602), .Z(n1603) );
  AND U2199 ( .A(n2843), .B(n2844), .Z(n1602) );
  XOR U2200 ( .A(n1608), .B(n1600), .Z(n1601) );
  AND U2201 ( .A(n2845), .B(n2846), .Z(n1600) );
  XNOR U2202 ( .A(n1517), .B(n1607), .Z(n1608) );
  AND U2203 ( .A(n2847), .B(n2848), .Z(n1607) );
  XNOR U2204 ( .A(n1597), .B(n1518), .Z(n1517) );
  AND U2205 ( .A(n2849), .B(n2850), .Z(n1518) );
  XOR U2206 ( .A(n1596), .B(n1515), .Z(n1597) );
  AND U2207 ( .A(n2851), .B(n2852), .Z(n1515) );
  XOR U2208 ( .A(n1606), .B(n1514), .Z(n1596) );
  AND U2209 ( .A(n2853), .B(n2854), .Z(n1514) );
  XNOR U2210 ( .A(n1525), .B(n1513), .Z(n1606) );
  AND U2211 ( .A(n2855), .B(n2856), .Z(n1513) );
  XNOR U2212 ( .A(n1589), .B(n1526), .Z(n1525) );
  AND U2213 ( .A(n2857), .B(n2858), .Z(n1526) );
  XOR U2214 ( .A(n1588), .B(n1523), .Z(n1589) );
  AND U2215 ( .A(n2859), .B(n2860), .Z(n1523) );
  XOR U2216 ( .A(n1585), .B(n1522), .Z(n1588) );
  AND U2217 ( .A(n2861), .B(n2862), .Z(n1522) );
  XNOR U2218 ( .A(n1539), .B(n1521), .Z(n1585) );
  AND U2219 ( .A(n2863), .B(n2864), .Z(n1521) );
  XNOR U2220 ( .A(n1546), .B(n1540), .Z(n1539) );
  AND U2221 ( .A(n2865), .B(n2866), .Z(n1540) );
  XOR U2222 ( .A(n1545), .B(n1537), .Z(n1546) );
  AND U2223 ( .A(n2867), .B(n2868), .Z(n1537) );
  XOR U2224 ( .A(n1584), .B(n1536), .Z(n1545) );
  AND U2225 ( .A(n2869), .B(n2870), .Z(n1536) );
  XNOR U2226 ( .A(n1557), .B(n1535), .Z(n1584) );
  AND U2227 ( .A(n2871), .B(n2872), .Z(n1535) );
  XNOR U2228 ( .A(n1564), .B(n1558), .Z(n1557) );
  AND U2229 ( .A(n2873), .B(n2874), .Z(n1558) );
  XOR U2230 ( .A(n1563), .B(n1555), .Z(n1564) );
  AND U2231 ( .A(n2875), .B(n2876), .Z(n1555) );
  XOR U2232 ( .A(n1583), .B(n1554), .Z(n1563) );
  AND U2233 ( .A(n2877), .B(n2878), .Z(n1554) );
  XNOR U2234 ( .A(n2879), .B(n2880), .Z(n1583) );
  XOR U2235 ( .A(n2881), .B(n2882), .Z(n2880) );
  XOR U2236 ( .A(n2883), .B(n2884), .Z(n2882) );
  XNOR U2237 ( .A(n1581), .B(n1574), .Z(n2884) );
  XNOR U2238 ( .A(n2885), .B(n2886), .Z(n1574) );
  AND U2239 ( .A(n2887), .B(n2888), .Z(n2886) );
  NOR U2240 ( .A(n2889), .B(n2890), .Z(n2888) );
  NOR U2241 ( .A(n2891), .B(n2892), .Z(n2887) );
  AND U2242 ( .A(n2893), .B(n2894), .Z(n2892) );
  AND U2243 ( .A(n2895), .B(n2896), .Z(n2885) );
  NOR U2244 ( .A(n2897), .B(n2898), .Z(n2896) );
  AND U2245 ( .A(n2890), .B(n2899), .Z(n2898) );
  AND U2246 ( .A(n2891), .B(n2900), .Z(n2897) );
  NOR U2247 ( .A(n2901), .B(n2902), .Z(n2895) );
  XOR U2248 ( .A(n2903), .B(n2904), .Z(n2902) );
  AND U2249 ( .A(n2905), .B(n2906), .Z(n2904) );
  NOR U2250 ( .A(n2907), .B(n2908), .Z(n2906) );
  NOR U2251 ( .A(n2909), .B(n2910), .Z(n2905) );
  AND U2252 ( .A(n2911), .B(n2912), .Z(n2910) );
  AND U2253 ( .A(n2913), .B(n2914), .Z(n2903) );
  NOR U2254 ( .A(n2915), .B(n2916), .Z(n2914) );
  AND U2255 ( .A(n2908), .B(n2917), .Z(n2916) );
  AND U2256 ( .A(n2909), .B(n2918), .Z(n2915) );
  NOR U2257 ( .A(n2919), .B(n2920), .Z(n2913) );
  XOR U2258 ( .A(n2921), .B(n2922), .Z(n2920) );
  AND U2259 ( .A(n2923), .B(n2924), .Z(n2922) );
  NOR U2260 ( .A(n2925), .B(n2926), .Z(n2924) );
  NOR U2261 ( .A(n2927), .B(n2928), .Z(n2923) );
  AND U2262 ( .A(n2929), .B(n2930), .Z(n2928) );
  AND U2263 ( .A(n2931), .B(n2932), .Z(n2921) );
  NOR U2264 ( .A(n2933), .B(n2934), .Z(n2932) );
  AND U2265 ( .A(n2926), .B(n2935), .Z(n2934) );
  AND U2266 ( .A(n2927), .B(n2936), .Z(n2933) );
  NOR U2267 ( .A(n2937), .B(n2938), .Z(n2931) );
  XOR U2268 ( .A(n2939), .B(n2940), .Z(n2938) );
  AND U2269 ( .A(n2941), .B(n2942), .Z(n2940) );
  NOR U2270 ( .A(n2943), .B(n2944), .Z(n2942) );
  NOR U2271 ( .A(n2945), .B(n2946), .Z(n2941) );
  AND U2272 ( .A(n2947), .B(n2948), .Z(n2946) );
  AND U2273 ( .A(n2949), .B(n2950), .Z(n2939) );
  NOR U2274 ( .A(n2951), .B(n2952), .Z(n2950) );
  AND U2275 ( .A(n2944), .B(n2953), .Z(n2952) );
  AND U2276 ( .A(n2945), .B(n2954), .Z(n2951) );
  NOR U2277 ( .A(n2955), .B(n2956), .Z(n2949) );
  AND U2278 ( .A(n2957), .B(n2958), .Z(n2956) );
  AND U2279 ( .A(n2959), .B(n2960), .Z(n2958) );
  AND U2280 ( .A(n2961), .B(n2962), .Z(n2960) );
  AND U2281 ( .A(n2963), .B(n2964), .Z(n2962) );
  NOR U2282 ( .A(n2965), .B(n2966), .Z(n2963) );
  NOR U2283 ( .A(n2967), .B(n2968), .Z(n2961) );
  AND U2284 ( .A(n2969), .B(n2970), .Z(n2959) );
  NOR U2285 ( .A(n2971), .B(n2972), .Z(n2970) );
  NOR U2286 ( .A(n2973), .B(n2974), .Z(n2969) );
  AND U2287 ( .A(n2975), .B(n2976), .Z(n2957) );
  AND U2288 ( .A(n2977), .B(n2978), .Z(n2976) );
  NOR U2289 ( .A(n2979), .B(n2980), .Z(n2978) );
  NOR U2290 ( .A(n2981), .B(n2982), .Z(n2977) );
  AND U2291 ( .A(n2983), .B(n2984), .Z(n2975) );
  NOR U2292 ( .A(n2985), .B(n2986), .Z(n2984) );
  NOR U2293 ( .A(n2987), .B(n2988), .Z(n2983) );
  AND U2294 ( .A(n2943), .B(n2989), .Z(n2955) );
  AND U2295 ( .A(n2925), .B(n2990), .Z(n2937) );
  AND U2296 ( .A(n2907), .B(n2991), .Z(n2919) );
  AND U2297 ( .A(n2889), .B(n2992), .Z(n2901) );
  AND U2298 ( .A(n2993), .B(n2994), .Z(n1581) );
  XOR U2299 ( .A(n1579), .B(n1580), .Z(n2883) );
  AND U2300 ( .A(n2995), .B(n2996), .Z(n1580) );
  AND U2301 ( .A(n2997), .B(n2998), .Z(n1579) );
  XOR U2302 ( .A(n2999), .B(n3000), .Z(n2881) );
  XOR U2303 ( .A(n1575), .B(n1576), .Z(n3000) );
  AND U2304 ( .A(n3001), .B(n3002), .Z(n1576) );
  AND U2305 ( .A(n3003), .B(n3004), .Z(n1575) );
  XNOR U2306 ( .A(n1573), .B(n1572), .Z(n2999) );
  IV U2307 ( .A(n3005), .Z(n1572) );
  AND U2308 ( .A(n3006), .B(n3007), .Z(n3005) );
  AND U2309 ( .A(n3008), .B(n3009), .Z(n1573) );
  XNOR U2310 ( .A(n1582), .B(n1553), .Z(n2879) );
  AND U2311 ( .A(n3010), .B(n3011), .Z(n1553) );
  AND U2312 ( .A(n3012), .B(n3013), .Z(n1582) );
  XOR U2313 ( .A(n3014), .B(n3015), .Z(n1481) );
  AND U2314 ( .A(n3014), .B(n3016), .Z(n3015) );
  XOR U2315 ( .A(n3017), .B(n3018), .Z(n1479) );
  AND U2316 ( .A(n3017), .B(n3019), .Z(n3018) );
  IV U2317 ( .A(n1480), .Z(n1486) );
  XNOR U2318 ( .A(n3020), .B(n3021), .Z(n1480) );
  AND U2319 ( .A(n3020), .B(n3022), .Z(n3021) );
  XNOR U2320 ( .A(n3023), .B(n3024), .Z(n1704) );
  AND U2321 ( .A(n3023), .B(n3025), .Z(n3024) );
  XOR U2322 ( .A(n3026), .B(n3027), .Z(n1708) );
  AND U2323 ( .A(n3026), .B(n3028), .Z(n3027) );
  XNOR U2324 ( .A(n3029), .B(n3030), .Z(n1469) );
  AND U2325 ( .A(n3031), .B(n3029), .Z(n3030) );
  XOR U2326 ( .A(n3032), .B(n3033), .Z(n1470) );
  NOR U2327 ( .A(n3034), .B(n3032), .Z(n3033) );
  XOR U2328 ( .A(n3035), .B(n3036), .Z(n1716) );
  NOR U2329 ( .A(n3037), .B(n3035), .Z(n3036) );
  XOR U2330 ( .A(n3038), .B(n3039), .Z(n1717) );
  NOR U2331 ( .A(n3040), .B(n3038), .Z(n3039) );
  XOR U2332 ( .A(n3041), .B(n3042), .Z(n1718) );
  NOR U2333 ( .A(n3043), .B(n3041), .Z(n3042) );
  XOR U2334 ( .A(n3044), .B(n3045), .Z(n1463) );
  NOR U2335 ( .A(n3046), .B(n3044), .Z(n3045) );
  XOR U2336 ( .A(n3047), .B(n3048), .Z(n1456) );
  NOR U2337 ( .A(n3049), .B(n3047), .Z(n3048) );
  XOR U2338 ( .A(n3050), .B(n3051), .Z(n1452) );
  NOR U2339 ( .A(n3052), .B(n3050), .Z(n3051) );
  XOR U2340 ( .A(n3053), .B(n3054), .Z(n1454) );
  NOR U2341 ( .A(n3055), .B(n3053), .Z(n3054) );
  XOR U2342 ( .A(n3056), .B(n3057), .Z(n1732) );
  NOR U2343 ( .A(n3058), .B(n3056), .Z(n3057) );
  XOR U2344 ( .A(n3059), .B(n3060), .Z(n1733) );
  NOR U2345 ( .A(n3061), .B(n3059), .Z(n3060) );
  XOR U2346 ( .A(n3062), .B(n3063), .Z(n1736) );
  NOR U2347 ( .A(n3064), .B(n3062), .Z(n3063) );
  XOR U2348 ( .A(n3065), .B(n3066), .Z(n1739) );
  NOR U2349 ( .A(n3067), .B(n3065), .Z(n3066) );
  XOR U2350 ( .A(n3068), .B(n3069), .Z(n1742) );
  NOR U2351 ( .A(n3070), .B(n3068), .Z(n3069) );
  XOR U2352 ( .A(n3071), .B(n3072), .Z(n1745) );
  NOR U2353 ( .A(n3073), .B(n3071), .Z(n3072) );
  XOR U2354 ( .A(n3074), .B(n3075), .Z(n1748) );
  NOR U2355 ( .A(n3076), .B(n3074), .Z(n3075) );
  XOR U2356 ( .A(n3077), .B(n3078), .Z(n1751) );
  NOR U2357 ( .A(n3079), .B(n3077), .Z(n3078) );
  XOR U2358 ( .A(n3080), .B(n3081), .Z(n1754) );
  NOR U2359 ( .A(n3082), .B(n3080), .Z(n3081) );
  XOR U2360 ( .A(n3083), .B(n3084), .Z(n1757) );
  NOR U2361 ( .A(n3085), .B(n3083), .Z(n3084) );
  XOR U2362 ( .A(n3086), .B(n3087), .Z(n1760) );
  NOR U2363 ( .A(n3088), .B(n3086), .Z(n3087) );
  XOR U2364 ( .A(n3089), .B(n3090), .Z(n1763) );
  NOR U2365 ( .A(n3091), .B(n3089), .Z(n3090) );
  XOR U2366 ( .A(n3092), .B(n3093), .Z(n1766) );
  NOR U2367 ( .A(n3094), .B(n3092), .Z(n3093) );
  XOR U2368 ( .A(n3095), .B(n3096), .Z(n1769) );
  NOR U2369 ( .A(n3097), .B(n3095), .Z(n3096) );
  XOR U2370 ( .A(n3098), .B(n3099), .Z(n1772) );
  NOR U2371 ( .A(n3100), .B(n3098), .Z(n3099) );
  XOR U2372 ( .A(n3101), .B(n3102), .Z(n1775) );
  NOR U2373 ( .A(n3103), .B(n3101), .Z(n3102) );
  XOR U2374 ( .A(n3104), .B(n3105), .Z(n1778) );
  NOR U2375 ( .A(n3106), .B(n3104), .Z(n3105) );
  XOR U2376 ( .A(n3107), .B(n3108), .Z(n1781) );
  NOR U2377 ( .A(n3109), .B(n3107), .Z(n3108) );
  XOR U2378 ( .A(n3110), .B(n3111), .Z(n1784) );
  NOR U2379 ( .A(n3112), .B(n3110), .Z(n3111) );
  XOR U2380 ( .A(n3113), .B(n3114), .Z(n1787) );
  NOR U2381 ( .A(n3115), .B(n3113), .Z(n3114) );
  XOR U2382 ( .A(n3116), .B(n3117), .Z(n1790) );
  NOR U2383 ( .A(n3118), .B(n3116), .Z(n3117) );
  XOR U2384 ( .A(n3119), .B(n3120), .Z(n1793) );
  NOR U2385 ( .A(n3121), .B(n3119), .Z(n3120) );
  XOR U2386 ( .A(n3122), .B(n3123), .Z(n1796) );
  NOR U2387 ( .A(n3124), .B(n3122), .Z(n3123) );
  XOR U2388 ( .A(n3125), .B(n3126), .Z(n1799) );
  NOR U2389 ( .A(n3127), .B(n3125), .Z(n3126) );
  XOR U2390 ( .A(n3128), .B(n3129), .Z(n1802) );
  NOR U2391 ( .A(n3130), .B(n3128), .Z(n3129) );
  XOR U2392 ( .A(n3131), .B(n3132), .Z(n1805) );
  NOR U2393 ( .A(n3133), .B(n3131), .Z(n3132) );
  XOR U2394 ( .A(n3134), .B(n3135), .Z(n1808) );
  NOR U2395 ( .A(n3136), .B(n3134), .Z(n3135) );
  XOR U2396 ( .A(n3137), .B(n3138), .Z(n1811) );
  NOR U2397 ( .A(n3139), .B(n3137), .Z(n3138) );
  XOR U2398 ( .A(n3140), .B(n3141), .Z(n1814) );
  NOR U2399 ( .A(n3142), .B(n3140), .Z(n3141) );
  XOR U2400 ( .A(n3143), .B(n3144), .Z(n1817) );
  NOR U2401 ( .A(n3145), .B(n3143), .Z(n3144) );
  XOR U2402 ( .A(n3146), .B(n3147), .Z(n1820) );
  NOR U2403 ( .A(n3148), .B(n3146), .Z(n3147) );
  XOR U2404 ( .A(n3149), .B(n3150), .Z(n1823) );
  NOR U2405 ( .A(n3151), .B(n3149), .Z(n3150) );
  XOR U2406 ( .A(n3152), .B(n3153), .Z(n1826) );
  NOR U2407 ( .A(n3154), .B(n3152), .Z(n3153) );
  XOR U2408 ( .A(n3155), .B(n3156), .Z(n1829) );
  NOR U2409 ( .A(n3157), .B(n3155), .Z(n3156) );
  XOR U2410 ( .A(n3158), .B(n3159), .Z(n1832) );
  NOR U2411 ( .A(n3160), .B(n3158), .Z(n3159) );
  XOR U2412 ( .A(n3161), .B(n3162), .Z(n1835) );
  NOR U2413 ( .A(n3163), .B(n3161), .Z(n3162) );
  XOR U2414 ( .A(n3164), .B(n3165), .Z(n1838) );
  NOR U2415 ( .A(n3166), .B(n3164), .Z(n3165) );
  XOR U2416 ( .A(n3167), .B(n3168), .Z(n1841) );
  NOR U2417 ( .A(n3169), .B(n3167), .Z(n3168) );
  XOR U2418 ( .A(n3170), .B(n3171), .Z(n1844) );
  NOR U2419 ( .A(n3172), .B(n3170), .Z(n3171) );
  XOR U2420 ( .A(n3173), .B(n3174), .Z(n1847) );
  NOR U2421 ( .A(n3175), .B(n3173), .Z(n3174) );
  XOR U2422 ( .A(n3176), .B(n3177), .Z(n1850) );
  NOR U2423 ( .A(n3178), .B(n3176), .Z(n3177) );
  XOR U2424 ( .A(n3179), .B(n3180), .Z(n1853) );
  NOR U2425 ( .A(n3181), .B(n3179), .Z(n3180) );
  XOR U2426 ( .A(n3182), .B(n3183), .Z(n1856) );
  NOR U2427 ( .A(n3184), .B(n3182), .Z(n3183) );
  XOR U2428 ( .A(n3185), .B(n3186), .Z(n1859) );
  NOR U2429 ( .A(n3187), .B(n3185), .Z(n3186) );
  XOR U2430 ( .A(n3188), .B(n3189), .Z(n1862) );
  NOR U2431 ( .A(n3190), .B(n3188), .Z(n3189) );
  XOR U2432 ( .A(n3191), .B(n3192), .Z(n1865) );
  NOR U2433 ( .A(n3193), .B(n3191), .Z(n3192) );
  XOR U2434 ( .A(n3194), .B(n3195), .Z(n1868) );
  NOR U2435 ( .A(n3196), .B(n3194), .Z(n3195) );
  XOR U2436 ( .A(n3197), .B(n3198), .Z(n1871) );
  NOR U2437 ( .A(n3199), .B(n3197), .Z(n3198) );
  XOR U2438 ( .A(n3200), .B(n3201), .Z(n1874) );
  NOR U2439 ( .A(n3202), .B(n3200), .Z(n3201) );
  XOR U2440 ( .A(n3203), .B(n3204), .Z(n1877) );
  NOR U2441 ( .A(n3205), .B(n3203), .Z(n3204) );
  XOR U2442 ( .A(n3206), .B(n3207), .Z(n1880) );
  NOR U2443 ( .A(n3208), .B(n3206), .Z(n3207) );
  XOR U2444 ( .A(n3209), .B(n3210), .Z(n1883) );
  NOR U2445 ( .A(n3211), .B(n3209), .Z(n3210) );
  XOR U2446 ( .A(n3212), .B(n3213), .Z(n1886) );
  NOR U2447 ( .A(n3214), .B(n3212), .Z(n3213) );
  XOR U2448 ( .A(n3215), .B(n3216), .Z(n1889) );
  NOR U2449 ( .A(n3217), .B(n3215), .Z(n3216) );
  XOR U2450 ( .A(n3218), .B(n3219), .Z(n1892) );
  NOR U2451 ( .A(n3220), .B(n3218), .Z(n3219) );
  XOR U2452 ( .A(n3221), .B(n3222), .Z(n1895) );
  NOR U2453 ( .A(n3223), .B(n3221), .Z(n3222) );
  XOR U2454 ( .A(n3224), .B(n3225), .Z(n1898) );
  NOR U2455 ( .A(n3226), .B(n3224), .Z(n3225) );
  XOR U2456 ( .A(n3227), .B(n3228), .Z(n1901) );
  NOR U2457 ( .A(n3229), .B(n3227), .Z(n3228) );
  XOR U2458 ( .A(n3230), .B(n3231), .Z(n1904) );
  NOR U2459 ( .A(n3232), .B(n3230), .Z(n3231) );
  XOR U2460 ( .A(n3233), .B(n3234), .Z(n1907) );
  NOR U2461 ( .A(n3235), .B(n3233), .Z(n3234) );
  XOR U2462 ( .A(n3236), .B(n3237), .Z(n1910) );
  NOR U2463 ( .A(n3238), .B(n3236), .Z(n3237) );
  XOR U2464 ( .A(n3239), .B(n3240), .Z(n1913) );
  NOR U2465 ( .A(n3241), .B(n3239), .Z(n3240) );
  XOR U2466 ( .A(n3242), .B(n3243), .Z(n1916) );
  NOR U2467 ( .A(n3244), .B(n3242), .Z(n3243) );
  XOR U2468 ( .A(n3245), .B(n3246), .Z(n1919) );
  NOR U2469 ( .A(n3247), .B(n3245), .Z(n3246) );
  XOR U2470 ( .A(n3248), .B(n3249), .Z(n1922) );
  NOR U2471 ( .A(n3250), .B(n3248), .Z(n3249) );
  XOR U2472 ( .A(n3251), .B(n3252), .Z(n1925) );
  NOR U2473 ( .A(n3253), .B(n3251), .Z(n3252) );
  XOR U2474 ( .A(n3254), .B(n3255), .Z(n1928) );
  NOR U2475 ( .A(n3256), .B(n3254), .Z(n3255) );
  XOR U2476 ( .A(n3257), .B(n3258), .Z(n1931) );
  NOR U2477 ( .A(n3259), .B(n3257), .Z(n3258) );
  XOR U2478 ( .A(n3260), .B(n3261), .Z(n1934) );
  NOR U2479 ( .A(n3262), .B(n3260), .Z(n3261) );
  XOR U2480 ( .A(n3263), .B(n3264), .Z(n1937) );
  NOR U2481 ( .A(n3265), .B(n3263), .Z(n3264) );
  XOR U2482 ( .A(n3266), .B(n3267), .Z(n1940) );
  NOR U2483 ( .A(n3268), .B(n3266), .Z(n3267) );
  XOR U2484 ( .A(n3269), .B(n3270), .Z(n1943) );
  NOR U2485 ( .A(n3271), .B(n3269), .Z(n3270) );
  XOR U2486 ( .A(n3272), .B(n3273), .Z(n1946) );
  NOR U2487 ( .A(n3274), .B(n3272), .Z(n3273) );
  XOR U2488 ( .A(n3275), .B(n3276), .Z(n1949) );
  NOR U2489 ( .A(n3277), .B(n3275), .Z(n3276) );
  XOR U2490 ( .A(n3278), .B(n3279), .Z(n1952) );
  NOR U2491 ( .A(n3280), .B(n3278), .Z(n3279) );
  XOR U2492 ( .A(n3281), .B(n3282), .Z(n1955) );
  NOR U2493 ( .A(n3283), .B(n3281), .Z(n3282) );
  XOR U2494 ( .A(n3284), .B(n3285), .Z(n1958) );
  NOR U2495 ( .A(n3286), .B(n3284), .Z(n3285) );
  XOR U2496 ( .A(n3287), .B(n3288), .Z(n1961) );
  NOR U2497 ( .A(n3289), .B(n3287), .Z(n3288) );
  XOR U2498 ( .A(n3290), .B(n3291), .Z(n1964) );
  NOR U2499 ( .A(n3292), .B(n3290), .Z(n3291) );
  XOR U2500 ( .A(n3293), .B(n3294), .Z(n1967) );
  NOR U2501 ( .A(n3295), .B(n3293), .Z(n3294) );
  XOR U2502 ( .A(n3296), .B(n3297), .Z(n1970) );
  NOR U2503 ( .A(n3298), .B(n3296), .Z(n3297) );
  XOR U2504 ( .A(n3299), .B(n3300), .Z(n1973) );
  NOR U2505 ( .A(n3301), .B(n3299), .Z(n3300) );
  XOR U2506 ( .A(n3302), .B(n3303), .Z(n1976) );
  NOR U2507 ( .A(n3304), .B(n3302), .Z(n3303) );
  XOR U2508 ( .A(n3305), .B(n3306), .Z(n1979) );
  NOR U2509 ( .A(n3307), .B(n3305), .Z(n3306) );
  XOR U2510 ( .A(n3308), .B(n3309), .Z(n1982) );
  NOR U2511 ( .A(n3310), .B(n3308), .Z(n3309) );
  XOR U2512 ( .A(n3311), .B(n3312), .Z(n1985) );
  NOR U2513 ( .A(n3313), .B(n3311), .Z(n3312) );
  XOR U2514 ( .A(n3314), .B(n3315), .Z(n1988) );
  NOR U2515 ( .A(n3316), .B(n3314), .Z(n3315) );
  XOR U2516 ( .A(n3317), .B(n3318), .Z(n1991) );
  NOR U2517 ( .A(n3319), .B(n3317), .Z(n3318) );
  XOR U2518 ( .A(n3320), .B(n3321), .Z(n1994) );
  NOR U2519 ( .A(n3322), .B(n3320), .Z(n3321) );
  XOR U2520 ( .A(n3323), .B(n3324), .Z(n1997) );
  NOR U2521 ( .A(n3325), .B(n3323), .Z(n3324) );
  XOR U2522 ( .A(n3326), .B(n3327), .Z(n2000) );
  NOR U2523 ( .A(n3328), .B(n3326), .Z(n3327) );
  XOR U2524 ( .A(n3329), .B(n3330), .Z(n2003) );
  NOR U2525 ( .A(n3331), .B(n3329), .Z(n3330) );
  XOR U2526 ( .A(n3332), .B(n3333), .Z(n2006) );
  NOR U2527 ( .A(n3334), .B(n3332), .Z(n3333) );
  XOR U2528 ( .A(n3335), .B(n3336), .Z(n2009) );
  NOR U2529 ( .A(n3337), .B(n3335), .Z(n3336) );
  XOR U2530 ( .A(n3338), .B(n3339), .Z(n2012) );
  NOR U2531 ( .A(n3340), .B(n3338), .Z(n3339) );
  XOR U2532 ( .A(n3341), .B(n3342), .Z(n2015) );
  NOR U2533 ( .A(n3343), .B(n3341), .Z(n3342) );
  XOR U2534 ( .A(n3344), .B(n3345), .Z(n2018) );
  NOR U2535 ( .A(n3346), .B(n3344), .Z(n3345) );
  XOR U2536 ( .A(n3347), .B(n3348), .Z(n2021) );
  NOR U2537 ( .A(n3349), .B(n3347), .Z(n3348) );
  XOR U2538 ( .A(n3350), .B(n3351), .Z(n2024) );
  NOR U2539 ( .A(n3352), .B(n3350), .Z(n3351) );
  XOR U2540 ( .A(n3353), .B(n3354), .Z(n2027) );
  NOR U2541 ( .A(n3355), .B(n3353), .Z(n3354) );
  XOR U2542 ( .A(n3356), .B(n3357), .Z(n2030) );
  NOR U2543 ( .A(n3358), .B(n3356), .Z(n3357) );
  XOR U2544 ( .A(n3359), .B(n3360), .Z(n2033) );
  NOR U2545 ( .A(n3361), .B(n3359), .Z(n3360) );
  XOR U2546 ( .A(n3362), .B(n3363), .Z(n2036) );
  NOR U2547 ( .A(n3364), .B(n3362), .Z(n3363) );
  XOR U2548 ( .A(n3365), .B(n3366), .Z(n2039) );
  NOR U2549 ( .A(n3367), .B(n3365), .Z(n3366) );
  XOR U2550 ( .A(n3368), .B(n3369), .Z(n2042) );
  NOR U2551 ( .A(n3370), .B(n3368), .Z(n3369) );
  XOR U2552 ( .A(n3371), .B(n3372), .Z(n2045) );
  NOR U2553 ( .A(n3373), .B(n3371), .Z(n3372) );
  XOR U2554 ( .A(n3374), .B(n3375), .Z(n2048) );
  NOR U2555 ( .A(n3376), .B(n3374), .Z(n3375) );
  XOR U2556 ( .A(n3377), .B(n3378), .Z(n2051) );
  NOR U2557 ( .A(n3379), .B(n3377), .Z(n3378) );
  XOR U2558 ( .A(n3380), .B(n3381), .Z(n2054) );
  NOR U2559 ( .A(n3382), .B(n3380), .Z(n3381) );
  XOR U2560 ( .A(n3383), .B(n3384), .Z(n2057) );
  NOR U2561 ( .A(n3385), .B(n3383), .Z(n3384) );
  XOR U2562 ( .A(n3386), .B(n3387), .Z(n2060) );
  NOR U2563 ( .A(n3388), .B(n3386), .Z(n3387) );
  XOR U2564 ( .A(n3389), .B(n3390), .Z(n2063) );
  NOR U2565 ( .A(n3391), .B(n3389), .Z(n3390) );
  XOR U2566 ( .A(n3392), .B(n3393), .Z(n2066) );
  NOR U2567 ( .A(n3394), .B(n3392), .Z(n3393) );
  XOR U2568 ( .A(n3395), .B(n3396), .Z(n2069) );
  NOR U2569 ( .A(n3397), .B(n3395), .Z(n3396) );
  XOR U2570 ( .A(n3398), .B(n3399), .Z(n2072) );
  NOR U2571 ( .A(n3400), .B(n3398), .Z(n3399) );
  XOR U2572 ( .A(n3401), .B(n3402), .Z(n2075) );
  NOR U2573 ( .A(n3403), .B(n3401), .Z(n3402) );
  XOR U2574 ( .A(n3404), .B(n3405), .Z(n2078) );
  NOR U2575 ( .A(n3406), .B(n3404), .Z(n3405) );
  XOR U2576 ( .A(n3407), .B(n3408), .Z(n2081) );
  NOR U2577 ( .A(n3409), .B(n3407), .Z(n3408) );
  XOR U2578 ( .A(n3410), .B(n3411), .Z(n2084) );
  NOR U2579 ( .A(n3412), .B(n3410), .Z(n3411) );
  XOR U2580 ( .A(n3413), .B(n3414), .Z(n2087) );
  NOR U2581 ( .A(n3415), .B(n3413), .Z(n3414) );
  XOR U2582 ( .A(n3416), .B(n3417), .Z(n2090) );
  NOR U2583 ( .A(n3418), .B(n3416), .Z(n3417) );
  XOR U2584 ( .A(n3419), .B(n3420), .Z(n2093) );
  NOR U2585 ( .A(n3421), .B(n3419), .Z(n3420) );
  XOR U2586 ( .A(n3422), .B(n3423), .Z(n2096) );
  NOR U2587 ( .A(n3424), .B(n3422), .Z(n3423) );
  XOR U2588 ( .A(n3425), .B(n3426), .Z(n2099) );
  NOR U2589 ( .A(n3427), .B(n3425), .Z(n3426) );
  XOR U2590 ( .A(n3428), .B(n3429), .Z(n2102) );
  NOR U2591 ( .A(n3430), .B(n3428), .Z(n3429) );
  XOR U2592 ( .A(n3431), .B(n3432), .Z(n2105) );
  NOR U2593 ( .A(n3433), .B(n3431), .Z(n3432) );
  XOR U2594 ( .A(n3434), .B(n3435), .Z(n2108) );
  NOR U2595 ( .A(n3436), .B(n3434), .Z(n3435) );
  XOR U2596 ( .A(n3437), .B(n3438), .Z(n2111) );
  NOR U2597 ( .A(n3439), .B(n3437), .Z(n3438) );
  XOR U2598 ( .A(n3440), .B(n3441), .Z(n2114) );
  AND U2599 ( .A(n3442), .B(n3440), .Z(n3441) );
  XOR U2600 ( .A(n3443), .B(n3444), .Z(n2117) );
  AND U2601 ( .A(n73), .B(n3443), .Z(n3444) );
  XNOR U2602 ( .A(n3445), .B(n2795), .Z(n2797) );
  IV U2603 ( .A(n56), .Z(n3445) );
  XOR U2604 ( .A(n2792), .B(n2791), .Z(n56) );
  XNOR U2605 ( .A(n2789), .B(n2788), .Z(n2791) );
  XNOR U2606 ( .A(n2786), .B(n2785), .Z(n2788) );
  XNOR U2607 ( .A(n2783), .B(n2782), .Z(n2785) );
  XNOR U2608 ( .A(n2780), .B(n2779), .Z(n2782) );
  XNOR U2609 ( .A(n2777), .B(n2776), .Z(n2779) );
  XNOR U2610 ( .A(n2774), .B(n2773), .Z(n2776) );
  XNOR U2611 ( .A(n2771), .B(n2770), .Z(n2773) );
  XNOR U2612 ( .A(n2768), .B(n2767), .Z(n2770) );
  XNOR U2613 ( .A(n2765), .B(n2764), .Z(n2767) );
  XNOR U2614 ( .A(n2762), .B(n2761), .Z(n2764) );
  XNOR U2615 ( .A(n2759), .B(n2758), .Z(n2761) );
  XNOR U2616 ( .A(n2756), .B(n2755), .Z(n2758) );
  XNOR U2617 ( .A(n2753), .B(n2752), .Z(n2755) );
  XNOR U2618 ( .A(n2750), .B(n2749), .Z(n2752) );
  XNOR U2619 ( .A(n2747), .B(n2746), .Z(n2749) );
  XNOR U2620 ( .A(n2744), .B(n2743), .Z(n2746) );
  XNOR U2621 ( .A(n2741), .B(n2740), .Z(n2743) );
  XNOR U2622 ( .A(n2738), .B(n2737), .Z(n2740) );
  XNOR U2623 ( .A(n2735), .B(n2734), .Z(n2737) );
  XNOR U2624 ( .A(n2732), .B(n2731), .Z(n2734) );
  XNOR U2625 ( .A(n2729), .B(n2728), .Z(n2731) );
  XNOR U2626 ( .A(n2726), .B(n2725), .Z(n2728) );
  XNOR U2627 ( .A(n2723), .B(n2722), .Z(n2725) );
  XNOR U2628 ( .A(n2720), .B(n2719), .Z(n2722) );
  XNOR U2629 ( .A(n2717), .B(n2716), .Z(n2719) );
  XNOR U2630 ( .A(n2714), .B(n2713), .Z(n2716) );
  XNOR U2631 ( .A(n2711), .B(n2710), .Z(n2713) );
  XNOR U2632 ( .A(n2708), .B(n2707), .Z(n2710) );
  XNOR U2633 ( .A(n2705), .B(n2704), .Z(n2707) );
  XNOR U2634 ( .A(n2702), .B(n2701), .Z(n2704) );
  XNOR U2635 ( .A(n2699), .B(n2698), .Z(n2701) );
  XNOR U2636 ( .A(n2696), .B(n2695), .Z(n2698) );
  XNOR U2637 ( .A(n2693), .B(n2692), .Z(n2695) );
  XNOR U2638 ( .A(n2690), .B(n2689), .Z(n2692) );
  XNOR U2639 ( .A(n2687), .B(n2686), .Z(n2689) );
  XNOR U2640 ( .A(n2684), .B(n2683), .Z(n2686) );
  XNOR U2641 ( .A(n2681), .B(n2680), .Z(n2683) );
  XNOR U2642 ( .A(n2678), .B(n2677), .Z(n2680) );
  XNOR U2643 ( .A(n2675), .B(n2674), .Z(n2677) );
  XNOR U2644 ( .A(n2672), .B(n2671), .Z(n2674) );
  XNOR U2645 ( .A(n2669), .B(n2668), .Z(n2671) );
  XNOR U2646 ( .A(n2666), .B(n2665), .Z(n2668) );
  XNOR U2647 ( .A(n2663), .B(n2662), .Z(n2665) );
  XNOR U2648 ( .A(n2660), .B(n2659), .Z(n2662) );
  XNOR U2649 ( .A(n2657), .B(n2656), .Z(n2659) );
  XNOR U2650 ( .A(n2654), .B(n2653), .Z(n2656) );
  XNOR U2651 ( .A(n2651), .B(n2650), .Z(n2653) );
  XNOR U2652 ( .A(n2648), .B(n2647), .Z(n2650) );
  XNOR U2653 ( .A(n2645), .B(n2644), .Z(n2647) );
  XNOR U2654 ( .A(n2642), .B(n2641), .Z(n2644) );
  XNOR U2655 ( .A(n2639), .B(n2638), .Z(n2641) );
  XNOR U2656 ( .A(n2636), .B(n2635), .Z(n2638) );
  XNOR U2657 ( .A(n2633), .B(n2632), .Z(n2635) );
  XNOR U2658 ( .A(n2630), .B(n2629), .Z(n2632) );
  XNOR U2659 ( .A(n2627), .B(n2626), .Z(n2629) );
  XNOR U2660 ( .A(n2624), .B(n2623), .Z(n2626) );
  XNOR U2661 ( .A(n2621), .B(n2620), .Z(n2623) );
  XNOR U2662 ( .A(n2618), .B(n2617), .Z(n2620) );
  XNOR U2663 ( .A(n2615), .B(n2614), .Z(n2617) );
  XNOR U2664 ( .A(n2612), .B(n2611), .Z(n2614) );
  XNOR U2665 ( .A(n2609), .B(n2608), .Z(n2611) );
  XNOR U2666 ( .A(n2606), .B(n2605), .Z(n2608) );
  XNOR U2667 ( .A(n2603), .B(n2602), .Z(n2605) );
  XNOR U2668 ( .A(n2600), .B(n2599), .Z(n2602) );
  XNOR U2669 ( .A(n2597), .B(n2596), .Z(n2599) );
  XNOR U2670 ( .A(n2594), .B(n2593), .Z(n2596) );
  XNOR U2671 ( .A(n2591), .B(n2590), .Z(n2593) );
  XNOR U2672 ( .A(n2588), .B(n2587), .Z(n2590) );
  XNOR U2673 ( .A(n2585), .B(n2584), .Z(n2587) );
  XNOR U2674 ( .A(n2582), .B(n2581), .Z(n2584) );
  XNOR U2675 ( .A(n2579), .B(n2578), .Z(n2581) );
  XNOR U2676 ( .A(n2576), .B(n2575), .Z(n2578) );
  XNOR U2677 ( .A(n2573), .B(n2572), .Z(n2575) );
  XNOR U2678 ( .A(n2570), .B(n2569), .Z(n2572) );
  XNOR U2679 ( .A(n2567), .B(n2566), .Z(n2569) );
  XNOR U2680 ( .A(n2564), .B(n2563), .Z(n2566) );
  XNOR U2681 ( .A(n2561), .B(n2560), .Z(n2563) );
  XNOR U2682 ( .A(n2558), .B(n2557), .Z(n2560) );
  XNOR U2683 ( .A(n2555), .B(n2554), .Z(n2557) );
  XNOR U2684 ( .A(n2552), .B(n2551), .Z(n2554) );
  XNOR U2685 ( .A(n2549), .B(n2548), .Z(n2551) );
  XNOR U2686 ( .A(n2546), .B(n2545), .Z(n2548) );
  XNOR U2687 ( .A(n2543), .B(n2542), .Z(n2545) );
  XNOR U2688 ( .A(n2540), .B(n2539), .Z(n2542) );
  XNOR U2689 ( .A(n2537), .B(n2536), .Z(n2539) );
  XNOR U2690 ( .A(n2534), .B(n2533), .Z(n2536) );
  XNOR U2691 ( .A(n2531), .B(n2530), .Z(n2533) );
  XNOR U2692 ( .A(n2528), .B(n2527), .Z(n2530) );
  XNOR U2693 ( .A(n2525), .B(n2524), .Z(n2527) );
  XNOR U2694 ( .A(n2522), .B(n2521), .Z(n2524) );
  XNOR U2695 ( .A(n2519), .B(n2518), .Z(n2521) );
  XNOR U2696 ( .A(n2516), .B(n2515), .Z(n2518) );
  XNOR U2697 ( .A(n2513), .B(n2512), .Z(n2515) );
  XNOR U2698 ( .A(n2510), .B(n2509), .Z(n2512) );
  XNOR U2699 ( .A(n2507), .B(n2506), .Z(n2509) );
  XNOR U2700 ( .A(n2504), .B(n2503), .Z(n2506) );
  XNOR U2701 ( .A(n2501), .B(n2500), .Z(n2503) );
  XNOR U2702 ( .A(n2498), .B(n2497), .Z(n2500) );
  XNOR U2703 ( .A(n2495), .B(n2494), .Z(n2497) );
  XNOR U2704 ( .A(n2492), .B(n2491), .Z(n2494) );
  XNOR U2705 ( .A(n2489), .B(n2488), .Z(n2491) );
  XNOR U2706 ( .A(n2486), .B(n2485), .Z(n2488) );
  XNOR U2707 ( .A(n2483), .B(n2482), .Z(n2485) );
  XNOR U2708 ( .A(n2480), .B(n2479), .Z(n2482) );
  XNOR U2709 ( .A(n2477), .B(n2476), .Z(n2479) );
  XNOR U2710 ( .A(n2474), .B(n2473), .Z(n2476) );
  XNOR U2711 ( .A(n2471), .B(n2470), .Z(n2473) );
  XNOR U2712 ( .A(n2468), .B(n2467), .Z(n2470) );
  XNOR U2713 ( .A(n2465), .B(n2464), .Z(n2467) );
  XNOR U2714 ( .A(n2462), .B(n2461), .Z(n2464) );
  XNOR U2715 ( .A(n2459), .B(n2458), .Z(n2461) );
  XNOR U2716 ( .A(n2456), .B(n2455), .Z(n2458) );
  XNOR U2717 ( .A(n2453), .B(n2452), .Z(n2455) );
  XNOR U2718 ( .A(n2450), .B(n2449), .Z(n2452) );
  XNOR U2719 ( .A(n2447), .B(n2446), .Z(n2449) );
  XNOR U2720 ( .A(n2444), .B(n2443), .Z(n2446) );
  XNOR U2721 ( .A(n2441), .B(n2440), .Z(n2443) );
  XNOR U2722 ( .A(n2438), .B(n2437), .Z(n2440) );
  XNOR U2723 ( .A(n2435), .B(n2434), .Z(n2437) );
  XNOR U2724 ( .A(n2432), .B(n2431), .Z(n2434) );
  XNOR U2725 ( .A(n2429), .B(n2428), .Z(n2431) );
  XNOR U2726 ( .A(n2426), .B(n2425), .Z(n2428) );
  XNOR U2727 ( .A(n2423), .B(n2422), .Z(n2425) );
  XNOR U2728 ( .A(n2420), .B(n2419), .Z(n2422) );
  XNOR U2729 ( .A(n2417), .B(n2416), .Z(n2419) );
  XNOR U2730 ( .A(n2414), .B(n2413), .Z(n2416) );
  XNOR U2731 ( .A(n2411), .B(n2410), .Z(n2413) );
  XOR U2732 ( .A(n2408), .B(n2143), .Z(n2410) );
  XOR U2733 ( .A(n3446), .B(n2131), .Z(n2143) );
  XNOR U2734 ( .A(n2132), .B(n2129), .Z(n2131) );
  XNOR U2735 ( .A(n2130), .B(n2126), .Z(n2129) );
  XNOR U2736 ( .A(n2125), .B(n2152), .Z(n2126) );
  XNOR U2737 ( .A(n2151), .B(n2407), .Z(n2152) );
  XNOR U2738 ( .A(n2398), .B(n2406), .Z(n2407) );
  XNOR U2739 ( .A(n2397), .B(n2403), .Z(n2406) );
  XNOR U2740 ( .A(n2402), .B(n2161), .Z(n2403) );
  XNOR U2741 ( .A(n2160), .B(n2396), .Z(n2161) );
  XNOR U2742 ( .A(n2387), .B(n2395), .Z(n2396) );
  XOR U2743 ( .A(n2386), .B(n2392), .Z(n2395) );
  XOR U2744 ( .A(n2391), .B(n2373), .Z(n2392) );
  XOR U2745 ( .A(n2167), .B(n2384), .Z(n2373) );
  XOR U2746 ( .A(n2385), .B(n2383), .Z(n2384) );
  XOR U2747 ( .A(n2374), .B(n2380), .Z(n2383) );
  XOR U2748 ( .A(n2178), .B(n2379), .Z(n2380) );
  AND U2749 ( .A(n3447), .B(n3448), .Z(n2379) );
  XOR U2750 ( .A(n2372), .B(n2177), .Z(n2178) );
  AND U2751 ( .A(n3449), .B(n3450), .Z(n2177) );
  XOR U2752 ( .A(n2369), .B(n2169), .Z(n2372) );
  AND U2753 ( .A(n3451), .B(n3452), .Z(n2169) );
  XNOR U2754 ( .A(n2367), .B(n2168), .Z(n2369) );
  AND U2755 ( .A(n3453), .B(n3454), .Z(n2168) );
  XOR U2756 ( .A(n2331), .B(n2368), .Z(n2367) );
  AND U2757 ( .A(n3455), .B(n3456), .Z(n2368) );
  XNOR U2758 ( .A(n2362), .B(n2332), .Z(n2331) );
  AND U2759 ( .A(n3457), .B(n3458), .Z(n2332) );
  XOR U2760 ( .A(n2361), .B(n2353), .Z(n2362) );
  AND U2761 ( .A(n3459), .B(n3460), .Z(n2353) );
  XNOR U2762 ( .A(n2356), .B(n2352), .Z(n2361) );
  AND U2763 ( .A(n3461), .B(n3462), .Z(n2352) );
  XOR U2764 ( .A(n2333), .B(n2357), .Z(n2356) );
  AND U2765 ( .A(n3463), .B(n3464), .Z(n2357) );
  XNOR U2766 ( .A(n2349), .B(n2334), .Z(n2333) );
  AND U2767 ( .A(n3465), .B(n3466), .Z(n2334) );
  XOR U2768 ( .A(n2348), .B(n2340), .Z(n2349) );
  AND U2769 ( .A(n3467), .B(n3468), .Z(n2340) );
  XNOR U2770 ( .A(n2343), .B(n2339), .Z(n2348) );
  AND U2771 ( .A(n3469), .B(n3470), .Z(n2339) );
  XOR U2772 ( .A(n2286), .B(n2344), .Z(n2343) );
  AND U2773 ( .A(n3471), .B(n3472), .Z(n2344) );
  XNOR U2774 ( .A(n2328), .B(n2287), .Z(n2286) );
  AND U2775 ( .A(n3473), .B(n3474), .Z(n2287) );
  XOR U2776 ( .A(n2327), .B(n2319), .Z(n2328) );
  AND U2777 ( .A(n3475), .B(n3476), .Z(n2319) );
  XNOR U2778 ( .A(n2322), .B(n2318), .Z(n2327) );
  AND U2779 ( .A(n3477), .B(n3478), .Z(n2318) );
  XOR U2780 ( .A(n2290), .B(n2323), .Z(n2322) );
  AND U2781 ( .A(n3479), .B(n3480), .Z(n2323) );
  XNOR U2782 ( .A(n2315), .B(n2291), .Z(n2290) );
  AND U2783 ( .A(n3481), .B(n3482), .Z(n2291) );
  XOR U2784 ( .A(n2314), .B(n2306), .Z(n2315) );
  AND U2785 ( .A(n3483), .B(n3484), .Z(n2306) );
  XNOR U2786 ( .A(n2309), .B(n2305), .Z(n2314) );
  AND U2787 ( .A(n3485), .B(n3486), .Z(n2305) );
  XOR U2788 ( .A(n2250), .B(n2310), .Z(n2309) );
  AND U2789 ( .A(n3487), .B(n3488), .Z(n2310) );
  XNOR U2790 ( .A(n2300), .B(n2251), .Z(n2250) );
  AND U2791 ( .A(n3489), .B(n3490), .Z(n2251) );
  XOR U2792 ( .A(n2299), .B(n2285), .Z(n2300) );
  AND U2793 ( .A(n3491), .B(n3492), .Z(n2285) );
  XNOR U2794 ( .A(n2294), .B(n2284), .Z(n2299) );
  AND U2795 ( .A(n3493), .B(n3494), .Z(n2284) );
  XOR U2796 ( .A(n2254), .B(n2295), .Z(n2294) );
  AND U2797 ( .A(n3495), .B(n3496), .Z(n2295) );
  XNOR U2798 ( .A(n2283), .B(n2255), .Z(n2254) );
  AND U2799 ( .A(n3497), .B(n3498), .Z(n2255) );
  XOR U2800 ( .A(n2282), .B(n2272), .Z(n2283) );
  AND U2801 ( .A(n3499), .B(n3500), .Z(n2272) );
  XNOR U2802 ( .A(n2277), .B(n2271), .Z(n2282) );
  AND U2803 ( .A(n3501), .B(n3502), .Z(n2271) );
  XOR U2804 ( .A(n2197), .B(n2278), .Z(n2277) );
  AND U2805 ( .A(n3503), .B(n3504), .Z(n2278) );
  XNOR U2806 ( .A(n2270), .B(n2198), .Z(n2197) );
  AND U2807 ( .A(n3505), .B(n3506), .Z(n2198) );
  XOR U2808 ( .A(n2269), .B(n2257), .Z(n2270) );
  AND U2809 ( .A(n3507), .B(n3508), .Z(n2257) );
  XNOR U2810 ( .A(n2264), .B(n2256), .Z(n2269) );
  AND U2811 ( .A(n3509), .B(n3510), .Z(n2256) );
  XOR U2812 ( .A(n2199), .B(n2265), .Z(n2264) );
  AND U2813 ( .A(n3511), .B(n3512), .Z(n2265) );
  XNOR U2814 ( .A(n2249), .B(n2200), .Z(n2199) );
  AND U2815 ( .A(n3513), .B(n3514), .Z(n2200) );
  XOR U2816 ( .A(n2248), .B(n2240), .Z(n2249) );
  AND U2817 ( .A(n3515), .B(n3516), .Z(n2240) );
  XNOR U2818 ( .A(n2243), .B(n2239), .Z(n2248) );
  AND U2819 ( .A(n3517), .B(n3518), .Z(n2239) );
  XOR U2820 ( .A(n2203), .B(n2244), .Z(n2243) );
  AND U2821 ( .A(n3519), .B(n3520), .Z(n2244) );
  XNOR U2822 ( .A(n2236), .B(n2204), .Z(n2203) );
  AND U2823 ( .A(n3521), .B(n3522), .Z(n2204) );
  XOR U2824 ( .A(n2235), .B(n2227), .Z(n2236) );
  AND U2825 ( .A(n3523), .B(n3524), .Z(n2227) );
  XNOR U2826 ( .A(n2230), .B(n2226), .Z(n2235) );
  AND U2827 ( .A(n3525), .B(n3526), .Z(n2226) );
  XOR U2828 ( .A(n3527), .B(n3528), .Z(n2230) );
  XOR U2829 ( .A(n3529), .B(n3530), .Z(n3528) );
  XOR U2830 ( .A(n3531), .B(n3532), .Z(n3530) );
  XNOR U2831 ( .A(n2220), .B(n2213), .Z(n3532) );
  XOR U2832 ( .A(n3533), .B(n3534), .Z(n2213) );
  XOR U2833 ( .A(n3535), .B(n3536), .Z(n3534) );
  XOR U2834 ( .A(n3537), .B(n3538), .Z(n3536) );
  NOR U2835 ( .A(n3539), .B(n3540), .Z(n3538) );
  NOR U2836 ( .A(n3541), .B(n3542), .Z(n3537) );
  AND U2837 ( .A(n3543), .B(n3544), .Z(n3542) );
  IV U2838 ( .A(n3545), .Z(n3541) );
  NOR U2839 ( .A(n3546), .B(n3547), .Z(n3545) );
  AND U2840 ( .A(n3539), .B(n3548), .Z(n3547) );
  AND U2841 ( .A(n3540), .B(n3549), .Z(n3546) );
  NOR U2842 ( .A(n3550), .B(n3551), .Z(n3535) );
  AND U2843 ( .A(n3552), .B(n3553), .Z(n3551) );
  IV U2844 ( .A(n3554), .Z(n3550) );
  NOR U2845 ( .A(n3555), .B(n3556), .Z(n3554) );
  AND U2846 ( .A(n3557), .B(n3558), .Z(n3556) );
  AND U2847 ( .A(n3559), .B(n3560), .Z(n3555) );
  XOR U2848 ( .A(n3561), .B(n3562), .Z(n3533) );
  XOR U2849 ( .A(n3563), .B(n3564), .Z(n3562) );
  XOR U2850 ( .A(n3565), .B(n3566), .Z(n3564) );
  XOR U2851 ( .A(n3567), .B(n3568), .Z(n3566) );
  AND U2852 ( .A(n3569), .B(n3570), .Z(n3568) );
  AND U2853 ( .A(n3571), .B(n3572), .Z(n3567) );
  XOR U2854 ( .A(n3573), .B(n3574), .Z(n3565) );
  AND U2855 ( .A(n3575), .B(n3576), .Z(n3574) );
  AND U2856 ( .A(n3577), .B(n3578), .Z(n3573) );
  AND U2857 ( .A(n3579), .B(n3580), .Z(n3578) );
  AND U2858 ( .A(n3581), .B(n3582), .Z(n3580) );
  NOR U2859 ( .A(n3583), .B(n3584), .Z(n3582) );
  IV U2860 ( .A(n3585), .Z(n3583) );
  NOR U2861 ( .A(n3586), .B(n3587), .Z(n3585) );
  NOR U2862 ( .A(n3588), .B(n3589), .Z(n3581) );
  AND U2863 ( .A(n3590), .B(n3591), .Z(n3579) );
  NOR U2864 ( .A(n3592), .B(n3593), .Z(n3591) );
  NOR U2865 ( .A(n3594), .B(n3595), .Z(n3590) );
  AND U2866 ( .A(n3596), .B(n3597), .Z(n3577) );
  AND U2867 ( .A(n3598), .B(n3599), .Z(n3597) );
  NOR U2868 ( .A(n3600), .B(n3601), .Z(n3599) );
  NOR U2869 ( .A(n3602), .B(n3603), .Z(n3598) );
  AND U2870 ( .A(n3604), .B(n3605), .Z(n3596) );
  NOR U2871 ( .A(n3606), .B(n3607), .Z(n3605) );
  NOR U2872 ( .A(n3608), .B(n3609), .Z(n3604) );
  XOR U2873 ( .A(n3610), .B(n3611), .Z(n3563) );
  XOR U2874 ( .A(n3612), .B(n3613), .Z(n3611) );
  NOR U2875 ( .A(n3614), .B(n3615), .Z(n3613) );
  NOR U2876 ( .A(n3616), .B(n3617), .Z(n3612) );
  AND U2877 ( .A(n3618), .B(n3619), .Z(n3617) );
  IV U2878 ( .A(n3620), .Z(n3616) );
  NOR U2879 ( .A(n3621), .B(n3622), .Z(n3620) );
  AND U2880 ( .A(n3614), .B(n3623), .Z(n3622) );
  AND U2881 ( .A(n3615), .B(n3624), .Z(n3621) );
  XOR U2882 ( .A(n3625), .B(n3626), .Z(n3610) );
  NOR U2883 ( .A(n3627), .B(n3628), .Z(n3626) );
  NOR U2884 ( .A(n3629), .B(n3630), .Z(n3625) );
  AND U2885 ( .A(n3631), .B(n3632), .Z(n3630) );
  IV U2886 ( .A(n3633), .Z(n3629) );
  NOR U2887 ( .A(n3634), .B(n3635), .Z(n3633) );
  AND U2888 ( .A(n3627), .B(n3636), .Z(n3635) );
  AND U2889 ( .A(n3628), .B(n3637), .Z(n3634) );
  XNOR U2890 ( .A(n3638), .B(n3639), .Z(n3561) );
  AND U2891 ( .A(n3640), .B(n3641), .Z(n3639) );
  NOR U2892 ( .A(n3557), .B(n3559), .Z(n3638) );
  AND U2893 ( .A(n3642), .B(n3643), .Z(n2220) );
  XOR U2894 ( .A(n2218), .B(n2219), .Z(n3531) );
  AND U2895 ( .A(n3644), .B(n3645), .Z(n2219) );
  AND U2896 ( .A(n3646), .B(n3647), .Z(n2218) );
  XOR U2897 ( .A(n3648), .B(n3649), .Z(n3529) );
  XOR U2898 ( .A(n2214), .B(n2215), .Z(n3649) );
  AND U2899 ( .A(n3650), .B(n3651), .Z(n2215) );
  AND U2900 ( .A(n3652), .B(n3653), .Z(n2214) );
  XOR U2901 ( .A(n2212), .B(n2210), .Z(n3648) );
  AND U2902 ( .A(n3654), .B(n3655), .Z(n2210) );
  AND U2903 ( .A(n3656), .B(n3657), .Z(n2212) );
  XNOR U2904 ( .A(n2221), .B(n2231), .Z(n3527) );
  AND U2905 ( .A(n3658), .B(n3659), .Z(n2231) );
  AND U2906 ( .A(n3660), .B(n3661), .Z(n2221) );
  XOR U2907 ( .A(n3662), .B(n3663), .Z(n2374) );
  AND U2908 ( .A(n3662), .B(n3664), .Z(n3663) );
  IV U2909 ( .A(n2375), .Z(n2385) );
  XNOR U2910 ( .A(n3665), .B(n3666), .Z(n2375) );
  AND U2911 ( .A(n3665), .B(n3667), .Z(n3666) );
  XOR U2912 ( .A(n3668), .B(n3669), .Z(n2167) );
  AND U2913 ( .A(n3668), .B(n3670), .Z(n3669) );
  XOR U2914 ( .A(n3671), .B(n3672), .Z(n2391) );
  AND U2915 ( .A(n3671), .B(n3673), .Z(n3672) );
  XNOR U2916 ( .A(n3674), .B(n3675), .Z(n2386) );
  AND U2917 ( .A(n3674), .B(n3676), .Z(n3675) );
  XNOR U2918 ( .A(n3677), .B(n3678), .Z(n2387) );
  AND U2919 ( .A(n3679), .B(n3677), .Z(n3678) );
  XOR U2920 ( .A(n3680), .B(n3681), .Z(n2160) );
  NOR U2921 ( .A(n3682), .B(n3680), .Z(n3681) );
  XOR U2922 ( .A(n3683), .B(n3684), .Z(n2402) );
  NOR U2923 ( .A(n3685), .B(n3683), .Z(n3684) );
  XOR U2924 ( .A(n3686), .B(n3687), .Z(n2397) );
  NOR U2925 ( .A(n3688), .B(n3686), .Z(n3687) );
  XOR U2926 ( .A(n3689), .B(n3690), .Z(n2398) );
  NOR U2927 ( .A(n3691), .B(n3689), .Z(n3690) );
  XOR U2928 ( .A(n3692), .B(n3693), .Z(n2151) );
  NOR U2929 ( .A(n3694), .B(n3692), .Z(n3693) );
  XOR U2930 ( .A(n3695), .B(n3696), .Z(n2125) );
  NOR U2931 ( .A(n3697), .B(n3695), .Z(n3696) );
  XOR U2932 ( .A(n3698), .B(n3699), .Z(n2130) );
  NOR U2933 ( .A(n3700), .B(n3698), .Z(n3699) );
  XOR U2934 ( .A(n3701), .B(n3702), .Z(n2132) );
  NOR U2935 ( .A(n3703), .B(n3701), .Z(n3702) );
  IV U2936 ( .A(n2142), .Z(n3446) );
  XNOR U2937 ( .A(n3704), .B(n3705), .Z(n2142) );
  NOR U2938 ( .A(n3706), .B(n3704), .Z(n3705) );
  XOR U2939 ( .A(n3707), .B(n3708), .Z(n2408) );
  NOR U2940 ( .A(n3709), .B(n3707), .Z(n3708) );
  XOR U2941 ( .A(n3710), .B(n3711), .Z(n2411) );
  NOR U2942 ( .A(n3712), .B(n3710), .Z(n3711) );
  XOR U2943 ( .A(n3713), .B(n3714), .Z(n2414) );
  NOR U2944 ( .A(n3715), .B(n3713), .Z(n3714) );
  XOR U2945 ( .A(n3716), .B(n3717), .Z(n2417) );
  NOR U2946 ( .A(n3718), .B(n3716), .Z(n3717) );
  XOR U2947 ( .A(n3719), .B(n3720), .Z(n2420) );
  NOR U2948 ( .A(n3721), .B(n3719), .Z(n3720) );
  XOR U2949 ( .A(n3722), .B(n3723), .Z(n2423) );
  NOR U2950 ( .A(n3724), .B(n3722), .Z(n3723) );
  XOR U2951 ( .A(n3725), .B(n3726), .Z(n2426) );
  NOR U2952 ( .A(n3727), .B(n3725), .Z(n3726) );
  XOR U2953 ( .A(n3728), .B(n3729), .Z(n2429) );
  NOR U2954 ( .A(n3730), .B(n3728), .Z(n3729) );
  XOR U2955 ( .A(n3731), .B(n3732), .Z(n2432) );
  NOR U2956 ( .A(n3733), .B(n3731), .Z(n3732) );
  XOR U2957 ( .A(n3734), .B(n3735), .Z(n2435) );
  NOR U2958 ( .A(n3736), .B(n3734), .Z(n3735) );
  XOR U2959 ( .A(n3737), .B(n3738), .Z(n2438) );
  NOR U2960 ( .A(n3739), .B(n3737), .Z(n3738) );
  XOR U2961 ( .A(n3740), .B(n3741), .Z(n2441) );
  NOR U2962 ( .A(n3742), .B(n3740), .Z(n3741) );
  XOR U2963 ( .A(n3743), .B(n3744), .Z(n2444) );
  NOR U2964 ( .A(n3745), .B(n3743), .Z(n3744) );
  XOR U2965 ( .A(n3746), .B(n3747), .Z(n2447) );
  NOR U2966 ( .A(n3748), .B(n3746), .Z(n3747) );
  XOR U2967 ( .A(n3749), .B(n3750), .Z(n2450) );
  NOR U2968 ( .A(n3751), .B(n3749), .Z(n3750) );
  XOR U2969 ( .A(n3752), .B(n3753), .Z(n2453) );
  NOR U2970 ( .A(n3754), .B(n3752), .Z(n3753) );
  XOR U2971 ( .A(n3755), .B(n3756), .Z(n2456) );
  NOR U2972 ( .A(n3757), .B(n3755), .Z(n3756) );
  XOR U2973 ( .A(n3758), .B(n3759), .Z(n2459) );
  NOR U2974 ( .A(n3760), .B(n3758), .Z(n3759) );
  XOR U2975 ( .A(n3761), .B(n3762), .Z(n2462) );
  NOR U2976 ( .A(n3763), .B(n3761), .Z(n3762) );
  XOR U2977 ( .A(n3764), .B(n3765), .Z(n2465) );
  NOR U2978 ( .A(n3766), .B(n3764), .Z(n3765) );
  XOR U2979 ( .A(n3767), .B(n3768), .Z(n2468) );
  NOR U2980 ( .A(n3769), .B(n3767), .Z(n3768) );
  XOR U2981 ( .A(n3770), .B(n3771), .Z(n2471) );
  NOR U2982 ( .A(n3772), .B(n3770), .Z(n3771) );
  XOR U2983 ( .A(n3773), .B(n3774), .Z(n2474) );
  NOR U2984 ( .A(n3775), .B(n3773), .Z(n3774) );
  XOR U2985 ( .A(n3776), .B(n3777), .Z(n2477) );
  NOR U2986 ( .A(n3778), .B(n3776), .Z(n3777) );
  XOR U2987 ( .A(n3779), .B(n3780), .Z(n2480) );
  NOR U2988 ( .A(n3781), .B(n3779), .Z(n3780) );
  XOR U2989 ( .A(n3782), .B(n3783), .Z(n2483) );
  NOR U2990 ( .A(n3784), .B(n3782), .Z(n3783) );
  XOR U2991 ( .A(n3785), .B(n3786), .Z(n2486) );
  NOR U2992 ( .A(n3787), .B(n3785), .Z(n3786) );
  XOR U2993 ( .A(n3788), .B(n3789), .Z(n2489) );
  NOR U2994 ( .A(n3790), .B(n3788), .Z(n3789) );
  XOR U2995 ( .A(n3791), .B(n3792), .Z(n2492) );
  NOR U2996 ( .A(n3793), .B(n3791), .Z(n3792) );
  XOR U2997 ( .A(n3794), .B(n3795), .Z(n2495) );
  NOR U2998 ( .A(n3796), .B(n3794), .Z(n3795) );
  XOR U2999 ( .A(n3797), .B(n3798), .Z(n2498) );
  NOR U3000 ( .A(n3799), .B(n3797), .Z(n3798) );
  XOR U3001 ( .A(n3800), .B(n3801), .Z(n2501) );
  NOR U3002 ( .A(n3802), .B(n3800), .Z(n3801) );
  XOR U3003 ( .A(n3803), .B(n3804), .Z(n2504) );
  NOR U3004 ( .A(n3805), .B(n3803), .Z(n3804) );
  XOR U3005 ( .A(n3806), .B(n3807), .Z(n2507) );
  NOR U3006 ( .A(n3808), .B(n3806), .Z(n3807) );
  XOR U3007 ( .A(n3809), .B(n3810), .Z(n2510) );
  NOR U3008 ( .A(n3811), .B(n3809), .Z(n3810) );
  XOR U3009 ( .A(n3812), .B(n3813), .Z(n2513) );
  NOR U3010 ( .A(n3814), .B(n3812), .Z(n3813) );
  XOR U3011 ( .A(n3815), .B(n3816), .Z(n2516) );
  NOR U3012 ( .A(n3817), .B(n3815), .Z(n3816) );
  XOR U3013 ( .A(n3818), .B(n3819), .Z(n2519) );
  NOR U3014 ( .A(n3820), .B(n3818), .Z(n3819) );
  XOR U3015 ( .A(n3821), .B(n3822), .Z(n2522) );
  NOR U3016 ( .A(n3823), .B(n3821), .Z(n3822) );
  XOR U3017 ( .A(n3824), .B(n3825), .Z(n2525) );
  NOR U3018 ( .A(n3826), .B(n3824), .Z(n3825) );
  XOR U3019 ( .A(n3827), .B(n3828), .Z(n2528) );
  NOR U3020 ( .A(n3829), .B(n3827), .Z(n3828) );
  XOR U3021 ( .A(n3830), .B(n3831), .Z(n2531) );
  NOR U3022 ( .A(n3832), .B(n3830), .Z(n3831) );
  XOR U3023 ( .A(n3833), .B(n3834), .Z(n2534) );
  NOR U3024 ( .A(n3835), .B(n3833), .Z(n3834) );
  XOR U3025 ( .A(n3836), .B(n3837), .Z(n2537) );
  NOR U3026 ( .A(n3838), .B(n3836), .Z(n3837) );
  XOR U3027 ( .A(n3839), .B(n3840), .Z(n2540) );
  NOR U3028 ( .A(n3841), .B(n3839), .Z(n3840) );
  XOR U3029 ( .A(n3842), .B(n3843), .Z(n2543) );
  NOR U3030 ( .A(n3844), .B(n3842), .Z(n3843) );
  XOR U3031 ( .A(n3845), .B(n3846), .Z(n2546) );
  NOR U3032 ( .A(n3847), .B(n3845), .Z(n3846) );
  XOR U3033 ( .A(n3848), .B(n3849), .Z(n2549) );
  NOR U3034 ( .A(n3850), .B(n3848), .Z(n3849) );
  XOR U3035 ( .A(n3851), .B(n3852), .Z(n2552) );
  NOR U3036 ( .A(n3853), .B(n3851), .Z(n3852) );
  XOR U3037 ( .A(n3854), .B(n3855), .Z(n2555) );
  NOR U3038 ( .A(n3856), .B(n3854), .Z(n3855) );
  XOR U3039 ( .A(n3857), .B(n3858), .Z(n2558) );
  NOR U3040 ( .A(n3859), .B(n3857), .Z(n3858) );
  XOR U3041 ( .A(n3860), .B(n3861), .Z(n2561) );
  NOR U3042 ( .A(n3862), .B(n3860), .Z(n3861) );
  XOR U3043 ( .A(n3863), .B(n3864), .Z(n2564) );
  NOR U3044 ( .A(n3865), .B(n3863), .Z(n3864) );
  XOR U3045 ( .A(n3866), .B(n3867), .Z(n2567) );
  NOR U3046 ( .A(n3868), .B(n3866), .Z(n3867) );
  XOR U3047 ( .A(n3869), .B(n3870), .Z(n2570) );
  NOR U3048 ( .A(n3871), .B(n3869), .Z(n3870) );
  XOR U3049 ( .A(n3872), .B(n3873), .Z(n2573) );
  NOR U3050 ( .A(n3874), .B(n3872), .Z(n3873) );
  XOR U3051 ( .A(n3875), .B(n3876), .Z(n2576) );
  NOR U3052 ( .A(n3877), .B(n3875), .Z(n3876) );
  XOR U3053 ( .A(n3878), .B(n3879), .Z(n2579) );
  NOR U3054 ( .A(n3880), .B(n3878), .Z(n3879) );
  XOR U3055 ( .A(n3881), .B(n3882), .Z(n2582) );
  NOR U3056 ( .A(n3883), .B(n3881), .Z(n3882) );
  XOR U3057 ( .A(n3884), .B(n3885), .Z(n2585) );
  NOR U3058 ( .A(n3886), .B(n3884), .Z(n3885) );
  XOR U3059 ( .A(n3887), .B(n3888), .Z(n2588) );
  NOR U3060 ( .A(n3889), .B(n3887), .Z(n3888) );
  XOR U3061 ( .A(n3890), .B(n3891), .Z(n2591) );
  NOR U3062 ( .A(n3892), .B(n3890), .Z(n3891) );
  XOR U3063 ( .A(n3893), .B(n3894), .Z(n2594) );
  NOR U3064 ( .A(n3895), .B(n3893), .Z(n3894) );
  XOR U3065 ( .A(n3896), .B(n3897), .Z(n2597) );
  NOR U3066 ( .A(n3898), .B(n3896), .Z(n3897) );
  XOR U3067 ( .A(n3899), .B(n3900), .Z(n2600) );
  NOR U3068 ( .A(n3901), .B(n3899), .Z(n3900) );
  XOR U3069 ( .A(n3902), .B(n3903), .Z(n2603) );
  NOR U3070 ( .A(n3904), .B(n3902), .Z(n3903) );
  XOR U3071 ( .A(n3905), .B(n3906), .Z(n2606) );
  NOR U3072 ( .A(n3907), .B(n3905), .Z(n3906) );
  XOR U3073 ( .A(n3908), .B(n3909), .Z(n2609) );
  NOR U3074 ( .A(n3910), .B(n3908), .Z(n3909) );
  XOR U3075 ( .A(n3911), .B(n3912), .Z(n2612) );
  NOR U3076 ( .A(n3913), .B(n3911), .Z(n3912) );
  XOR U3077 ( .A(n3914), .B(n3915), .Z(n2615) );
  NOR U3078 ( .A(n3916), .B(n3914), .Z(n3915) );
  XOR U3079 ( .A(n3917), .B(n3918), .Z(n2618) );
  NOR U3080 ( .A(n3919), .B(n3917), .Z(n3918) );
  XOR U3081 ( .A(n3920), .B(n3921), .Z(n2621) );
  NOR U3082 ( .A(n3922), .B(n3920), .Z(n3921) );
  XOR U3083 ( .A(n3923), .B(n3924), .Z(n2624) );
  NOR U3084 ( .A(n3925), .B(n3923), .Z(n3924) );
  XOR U3085 ( .A(n3926), .B(n3927), .Z(n2627) );
  NOR U3086 ( .A(n3928), .B(n3926), .Z(n3927) );
  XOR U3087 ( .A(n3929), .B(n3930), .Z(n2630) );
  NOR U3088 ( .A(n3931), .B(n3929), .Z(n3930) );
  XOR U3089 ( .A(n3932), .B(n3933), .Z(n2633) );
  NOR U3090 ( .A(n3934), .B(n3932), .Z(n3933) );
  XOR U3091 ( .A(n3935), .B(n3936), .Z(n2636) );
  NOR U3092 ( .A(n3937), .B(n3935), .Z(n3936) );
  XOR U3093 ( .A(n3938), .B(n3939), .Z(n2639) );
  NOR U3094 ( .A(n3940), .B(n3938), .Z(n3939) );
  XOR U3095 ( .A(n3941), .B(n3942), .Z(n2642) );
  NOR U3096 ( .A(n3943), .B(n3941), .Z(n3942) );
  XOR U3097 ( .A(n3944), .B(n3945), .Z(n2645) );
  NOR U3098 ( .A(n3946), .B(n3944), .Z(n3945) );
  XOR U3099 ( .A(n3947), .B(n3948), .Z(n2648) );
  NOR U3100 ( .A(n3949), .B(n3947), .Z(n3948) );
  XOR U3101 ( .A(n3950), .B(n3951), .Z(n2651) );
  NOR U3102 ( .A(n3952), .B(n3950), .Z(n3951) );
  XOR U3103 ( .A(n3953), .B(n3954), .Z(n2654) );
  NOR U3104 ( .A(n3955), .B(n3953), .Z(n3954) );
  XOR U3105 ( .A(n3956), .B(n3957), .Z(n2657) );
  NOR U3106 ( .A(n3958), .B(n3956), .Z(n3957) );
  XOR U3107 ( .A(n3959), .B(n3960), .Z(n2660) );
  NOR U3108 ( .A(n3961), .B(n3959), .Z(n3960) );
  XOR U3109 ( .A(n3962), .B(n3963), .Z(n2663) );
  NOR U3110 ( .A(n3964), .B(n3962), .Z(n3963) );
  XOR U3111 ( .A(n3965), .B(n3966), .Z(n2666) );
  NOR U3112 ( .A(n3967), .B(n3965), .Z(n3966) );
  XOR U3113 ( .A(n3968), .B(n3969), .Z(n2669) );
  NOR U3114 ( .A(n3970), .B(n3968), .Z(n3969) );
  XOR U3115 ( .A(n3971), .B(n3972), .Z(n2672) );
  NOR U3116 ( .A(n3973), .B(n3971), .Z(n3972) );
  XOR U3117 ( .A(n3974), .B(n3975), .Z(n2675) );
  NOR U3118 ( .A(n3976), .B(n3974), .Z(n3975) );
  XOR U3119 ( .A(n3977), .B(n3978), .Z(n2678) );
  NOR U3120 ( .A(n3979), .B(n3977), .Z(n3978) );
  XOR U3121 ( .A(n3980), .B(n3981), .Z(n2681) );
  NOR U3122 ( .A(n3982), .B(n3980), .Z(n3981) );
  XOR U3123 ( .A(n3983), .B(n3984), .Z(n2684) );
  NOR U3124 ( .A(n3985), .B(n3983), .Z(n3984) );
  XOR U3125 ( .A(n3986), .B(n3987), .Z(n2687) );
  NOR U3126 ( .A(n3988), .B(n3986), .Z(n3987) );
  XOR U3127 ( .A(n3989), .B(n3990), .Z(n2690) );
  NOR U3128 ( .A(n3991), .B(n3989), .Z(n3990) );
  XOR U3129 ( .A(n3992), .B(n3993), .Z(n2693) );
  NOR U3130 ( .A(n3994), .B(n3992), .Z(n3993) );
  XOR U3131 ( .A(n3995), .B(n3996), .Z(n2696) );
  NOR U3132 ( .A(n3997), .B(n3995), .Z(n3996) );
  XOR U3133 ( .A(n3998), .B(n3999), .Z(n2699) );
  NOR U3134 ( .A(n4000), .B(n3998), .Z(n3999) );
  XOR U3135 ( .A(n4001), .B(n4002), .Z(n2702) );
  NOR U3136 ( .A(n4003), .B(n4001), .Z(n4002) );
  XOR U3137 ( .A(n4004), .B(n4005), .Z(n2705) );
  NOR U3138 ( .A(n4006), .B(n4004), .Z(n4005) );
  XOR U3139 ( .A(n4007), .B(n4008), .Z(n2708) );
  NOR U3140 ( .A(n4009), .B(n4007), .Z(n4008) );
  XOR U3141 ( .A(n4010), .B(n4011), .Z(n2711) );
  NOR U3142 ( .A(n4012), .B(n4010), .Z(n4011) );
  XOR U3143 ( .A(n4013), .B(n4014), .Z(n2714) );
  NOR U3144 ( .A(n4015), .B(n4013), .Z(n4014) );
  XOR U3145 ( .A(n4016), .B(n4017), .Z(n2717) );
  NOR U3146 ( .A(n4018), .B(n4016), .Z(n4017) );
  XOR U3147 ( .A(n4019), .B(n4020), .Z(n2720) );
  NOR U3148 ( .A(n4021), .B(n4019), .Z(n4020) );
  XOR U3149 ( .A(n4022), .B(n4023), .Z(n2723) );
  NOR U3150 ( .A(n4024), .B(n4022), .Z(n4023) );
  XOR U3151 ( .A(n4025), .B(n4026), .Z(n2726) );
  NOR U3152 ( .A(n4027), .B(n4025), .Z(n4026) );
  XOR U3153 ( .A(n4028), .B(n4029), .Z(n2729) );
  NOR U3154 ( .A(n4030), .B(n4028), .Z(n4029) );
  XOR U3155 ( .A(n4031), .B(n4032), .Z(n2732) );
  NOR U3156 ( .A(n4033), .B(n4031), .Z(n4032) );
  XOR U3157 ( .A(n4034), .B(n4035), .Z(n2735) );
  NOR U3158 ( .A(n4036), .B(n4034), .Z(n4035) );
  XOR U3159 ( .A(n4037), .B(n4038), .Z(n2738) );
  NOR U3160 ( .A(n4039), .B(n4037), .Z(n4038) );
  XOR U3161 ( .A(n4040), .B(n4041), .Z(n2741) );
  NOR U3162 ( .A(n4042), .B(n4040), .Z(n4041) );
  XOR U3163 ( .A(n4043), .B(n4044), .Z(n2744) );
  NOR U3164 ( .A(n4045), .B(n4043), .Z(n4044) );
  XOR U3165 ( .A(n4046), .B(n4047), .Z(n2747) );
  NOR U3166 ( .A(n4048), .B(n4046), .Z(n4047) );
  XOR U3167 ( .A(n4049), .B(n4050), .Z(n2750) );
  NOR U3168 ( .A(n4051), .B(n4049), .Z(n4050) );
  XOR U3169 ( .A(n4052), .B(n4053), .Z(n2753) );
  NOR U3170 ( .A(n4054), .B(n4052), .Z(n4053) );
  XOR U3171 ( .A(n4055), .B(n4056), .Z(n2756) );
  NOR U3172 ( .A(n4057), .B(n4055), .Z(n4056) );
  XOR U3173 ( .A(n4058), .B(n4059), .Z(n2759) );
  NOR U3174 ( .A(n4060), .B(n4058), .Z(n4059) );
  XOR U3175 ( .A(n4061), .B(n4062), .Z(n2762) );
  NOR U3176 ( .A(n4063), .B(n4061), .Z(n4062) );
  XOR U3177 ( .A(n4064), .B(n4065), .Z(n2765) );
  NOR U3178 ( .A(n4066), .B(n4064), .Z(n4065) );
  XOR U3179 ( .A(n4067), .B(n4068), .Z(n2768) );
  NOR U3180 ( .A(n4069), .B(n4067), .Z(n4068) );
  XOR U3181 ( .A(n4070), .B(n4071), .Z(n2771) );
  NOR U3182 ( .A(n4072), .B(n4070), .Z(n4071) );
  XOR U3183 ( .A(n4073), .B(n4074), .Z(n2774) );
  NOR U3184 ( .A(n4075), .B(n4073), .Z(n4074) );
  XOR U3185 ( .A(n4076), .B(n4077), .Z(n2777) );
  NOR U3186 ( .A(n4078), .B(n4076), .Z(n4077) );
  XOR U3187 ( .A(n4079), .B(n4080), .Z(n2780) );
  NOR U3188 ( .A(n4081), .B(n4079), .Z(n4080) );
  XOR U3189 ( .A(n4082), .B(n4083), .Z(n2783) );
  NOR U3190 ( .A(n4084), .B(n4082), .Z(n4083) );
  XOR U3191 ( .A(n4085), .B(n4086), .Z(n2786) );
  NOR U3192 ( .A(n4087), .B(n4085), .Z(n4086) );
  XOR U3193 ( .A(n4088), .B(n4089), .Z(n2789) );
  NOR U3194 ( .A(n4090), .B(n4088), .Z(n4089) );
  XOR U3195 ( .A(n4091), .B(n4092), .Z(n2792) );
  NOR U3196 ( .A(n71), .B(n4093), .Z(n4092) );
  IV U3197 ( .A(n4091), .Z(n4093) );
  XOR U3198 ( .A(n4094), .B(n4095), .Z(n2795) );
  AND U3199 ( .A(n4096), .B(n4097), .Z(n4095) );
  XOR U3200 ( .A(n4094), .B(n73), .Z(n4097) );
  XOR U3201 ( .A(n3443), .B(n3442), .Z(n73) );
  XNOR U3202 ( .A(n3440), .B(n3439), .Z(n3442) );
  XNOR U3203 ( .A(n3437), .B(n3436), .Z(n3439) );
  XNOR U3204 ( .A(n3434), .B(n3433), .Z(n3436) );
  XNOR U3205 ( .A(n3431), .B(n3430), .Z(n3433) );
  XNOR U3206 ( .A(n3428), .B(n3427), .Z(n3430) );
  XNOR U3207 ( .A(n3425), .B(n3424), .Z(n3427) );
  XNOR U3208 ( .A(n3422), .B(n3421), .Z(n3424) );
  XNOR U3209 ( .A(n3419), .B(n3418), .Z(n3421) );
  XNOR U3210 ( .A(n3416), .B(n3415), .Z(n3418) );
  XNOR U3211 ( .A(n3413), .B(n3412), .Z(n3415) );
  XNOR U3212 ( .A(n3410), .B(n3409), .Z(n3412) );
  XNOR U3213 ( .A(n3407), .B(n3406), .Z(n3409) );
  XNOR U3214 ( .A(n3404), .B(n3403), .Z(n3406) );
  XNOR U3215 ( .A(n3401), .B(n3400), .Z(n3403) );
  XNOR U3216 ( .A(n3398), .B(n3397), .Z(n3400) );
  XNOR U3217 ( .A(n3395), .B(n3394), .Z(n3397) );
  XNOR U3218 ( .A(n3392), .B(n3391), .Z(n3394) );
  XNOR U3219 ( .A(n3389), .B(n3388), .Z(n3391) );
  XNOR U3220 ( .A(n3386), .B(n3385), .Z(n3388) );
  XNOR U3221 ( .A(n3383), .B(n3382), .Z(n3385) );
  XNOR U3222 ( .A(n3380), .B(n3379), .Z(n3382) );
  XNOR U3223 ( .A(n3377), .B(n3376), .Z(n3379) );
  XNOR U3224 ( .A(n3374), .B(n3373), .Z(n3376) );
  XNOR U3225 ( .A(n3371), .B(n3370), .Z(n3373) );
  XNOR U3226 ( .A(n3368), .B(n3367), .Z(n3370) );
  XNOR U3227 ( .A(n3365), .B(n3364), .Z(n3367) );
  XNOR U3228 ( .A(n3362), .B(n3361), .Z(n3364) );
  XNOR U3229 ( .A(n3359), .B(n3358), .Z(n3361) );
  XNOR U3230 ( .A(n3356), .B(n3355), .Z(n3358) );
  XNOR U3231 ( .A(n3353), .B(n3352), .Z(n3355) );
  XNOR U3232 ( .A(n3350), .B(n3349), .Z(n3352) );
  XNOR U3233 ( .A(n3347), .B(n3346), .Z(n3349) );
  XNOR U3234 ( .A(n3344), .B(n3343), .Z(n3346) );
  XNOR U3235 ( .A(n3341), .B(n3340), .Z(n3343) );
  XNOR U3236 ( .A(n3338), .B(n3337), .Z(n3340) );
  XNOR U3237 ( .A(n3335), .B(n3334), .Z(n3337) );
  XNOR U3238 ( .A(n3332), .B(n3331), .Z(n3334) );
  XNOR U3239 ( .A(n3329), .B(n3328), .Z(n3331) );
  XNOR U3240 ( .A(n3326), .B(n3325), .Z(n3328) );
  XNOR U3241 ( .A(n3323), .B(n3322), .Z(n3325) );
  XNOR U3242 ( .A(n3320), .B(n3319), .Z(n3322) );
  XNOR U3243 ( .A(n3317), .B(n3316), .Z(n3319) );
  XNOR U3244 ( .A(n3314), .B(n3313), .Z(n3316) );
  XNOR U3245 ( .A(n3311), .B(n3310), .Z(n3313) );
  XNOR U3246 ( .A(n3308), .B(n3307), .Z(n3310) );
  XNOR U3247 ( .A(n3305), .B(n3304), .Z(n3307) );
  XNOR U3248 ( .A(n3302), .B(n3301), .Z(n3304) );
  XNOR U3249 ( .A(n3299), .B(n3298), .Z(n3301) );
  XNOR U3250 ( .A(n3296), .B(n3295), .Z(n3298) );
  XNOR U3251 ( .A(n3293), .B(n3292), .Z(n3295) );
  XNOR U3252 ( .A(n3290), .B(n3289), .Z(n3292) );
  XNOR U3253 ( .A(n3287), .B(n3286), .Z(n3289) );
  XNOR U3254 ( .A(n3284), .B(n3283), .Z(n3286) );
  XNOR U3255 ( .A(n3281), .B(n3280), .Z(n3283) );
  XNOR U3256 ( .A(n3278), .B(n3277), .Z(n3280) );
  XNOR U3257 ( .A(n3275), .B(n3274), .Z(n3277) );
  XNOR U3258 ( .A(n3272), .B(n3271), .Z(n3274) );
  XNOR U3259 ( .A(n3269), .B(n3268), .Z(n3271) );
  XNOR U3260 ( .A(n3266), .B(n3265), .Z(n3268) );
  XNOR U3261 ( .A(n3263), .B(n3262), .Z(n3265) );
  XNOR U3262 ( .A(n3260), .B(n3259), .Z(n3262) );
  XNOR U3263 ( .A(n3257), .B(n3256), .Z(n3259) );
  XNOR U3264 ( .A(n3254), .B(n3253), .Z(n3256) );
  XNOR U3265 ( .A(n3251), .B(n3250), .Z(n3253) );
  XNOR U3266 ( .A(n3248), .B(n3247), .Z(n3250) );
  XNOR U3267 ( .A(n3245), .B(n3244), .Z(n3247) );
  XNOR U3268 ( .A(n3242), .B(n3241), .Z(n3244) );
  XNOR U3269 ( .A(n3239), .B(n3238), .Z(n3241) );
  XNOR U3270 ( .A(n3236), .B(n3235), .Z(n3238) );
  XNOR U3271 ( .A(n3233), .B(n3232), .Z(n3235) );
  XNOR U3272 ( .A(n3230), .B(n3229), .Z(n3232) );
  XNOR U3273 ( .A(n3227), .B(n3226), .Z(n3229) );
  XNOR U3274 ( .A(n3224), .B(n3223), .Z(n3226) );
  XNOR U3275 ( .A(n3221), .B(n3220), .Z(n3223) );
  XNOR U3276 ( .A(n3218), .B(n3217), .Z(n3220) );
  XNOR U3277 ( .A(n3215), .B(n3214), .Z(n3217) );
  XNOR U3278 ( .A(n3212), .B(n3211), .Z(n3214) );
  XNOR U3279 ( .A(n3209), .B(n3208), .Z(n3211) );
  XNOR U3280 ( .A(n3206), .B(n3205), .Z(n3208) );
  XNOR U3281 ( .A(n3203), .B(n3202), .Z(n3205) );
  XNOR U3282 ( .A(n3200), .B(n3199), .Z(n3202) );
  XNOR U3283 ( .A(n3197), .B(n3196), .Z(n3199) );
  XNOR U3284 ( .A(n3194), .B(n3193), .Z(n3196) );
  XNOR U3285 ( .A(n3191), .B(n3190), .Z(n3193) );
  XNOR U3286 ( .A(n3188), .B(n3187), .Z(n3190) );
  XNOR U3287 ( .A(n3185), .B(n3184), .Z(n3187) );
  XNOR U3288 ( .A(n3182), .B(n3181), .Z(n3184) );
  XNOR U3289 ( .A(n3179), .B(n3178), .Z(n3181) );
  XNOR U3290 ( .A(n3176), .B(n3175), .Z(n3178) );
  XNOR U3291 ( .A(n3173), .B(n3172), .Z(n3175) );
  XNOR U3292 ( .A(n3170), .B(n3169), .Z(n3172) );
  XNOR U3293 ( .A(n3167), .B(n3166), .Z(n3169) );
  XNOR U3294 ( .A(n3164), .B(n3163), .Z(n3166) );
  XNOR U3295 ( .A(n3161), .B(n3160), .Z(n3163) );
  XNOR U3296 ( .A(n3158), .B(n3157), .Z(n3160) );
  XNOR U3297 ( .A(n3155), .B(n3154), .Z(n3157) );
  XNOR U3298 ( .A(n3152), .B(n3151), .Z(n3154) );
  XNOR U3299 ( .A(n3149), .B(n3148), .Z(n3151) );
  XNOR U3300 ( .A(n3146), .B(n3145), .Z(n3148) );
  XNOR U3301 ( .A(n3143), .B(n3142), .Z(n3145) );
  XNOR U3302 ( .A(n3140), .B(n3139), .Z(n3142) );
  XNOR U3303 ( .A(n3137), .B(n3136), .Z(n3139) );
  XNOR U3304 ( .A(n3134), .B(n3133), .Z(n3136) );
  XNOR U3305 ( .A(n3131), .B(n3130), .Z(n3133) );
  XNOR U3306 ( .A(n3128), .B(n3127), .Z(n3130) );
  XNOR U3307 ( .A(n3125), .B(n3124), .Z(n3127) );
  XNOR U3308 ( .A(n3122), .B(n3121), .Z(n3124) );
  XNOR U3309 ( .A(n3119), .B(n3118), .Z(n3121) );
  XNOR U3310 ( .A(n3116), .B(n3115), .Z(n3118) );
  XNOR U3311 ( .A(n3113), .B(n3112), .Z(n3115) );
  XNOR U3312 ( .A(n3110), .B(n3109), .Z(n3112) );
  XNOR U3313 ( .A(n3107), .B(n3106), .Z(n3109) );
  XNOR U3314 ( .A(n3104), .B(n3103), .Z(n3106) );
  XNOR U3315 ( .A(n3101), .B(n3100), .Z(n3103) );
  XNOR U3316 ( .A(n3098), .B(n3097), .Z(n3100) );
  XNOR U3317 ( .A(n3095), .B(n3094), .Z(n3097) );
  XNOR U3318 ( .A(n3092), .B(n3091), .Z(n3094) );
  XNOR U3319 ( .A(n3089), .B(n3088), .Z(n3091) );
  XNOR U3320 ( .A(n3086), .B(n3085), .Z(n3088) );
  XNOR U3321 ( .A(n3083), .B(n3082), .Z(n3085) );
  XNOR U3322 ( .A(n3080), .B(n3079), .Z(n3082) );
  XNOR U3323 ( .A(n3077), .B(n3076), .Z(n3079) );
  XNOR U3324 ( .A(n3074), .B(n3073), .Z(n3076) );
  XNOR U3325 ( .A(n3071), .B(n3070), .Z(n3073) );
  XNOR U3326 ( .A(n3068), .B(n3067), .Z(n3070) );
  XNOR U3327 ( .A(n3065), .B(n3064), .Z(n3067) );
  XNOR U3328 ( .A(n3062), .B(n3061), .Z(n3064) );
  XNOR U3329 ( .A(n3059), .B(n3058), .Z(n3061) );
  XNOR U3330 ( .A(n3056), .B(n3055), .Z(n3058) );
  XNOR U3331 ( .A(n3053), .B(n3052), .Z(n3055) );
  XNOR U3332 ( .A(n3050), .B(n3049), .Z(n3052) );
  XNOR U3333 ( .A(n3047), .B(n3046), .Z(n3049) );
  XNOR U3334 ( .A(n3044), .B(n3043), .Z(n3046) );
  XNOR U3335 ( .A(n3041), .B(n3040), .Z(n3043) );
  XNOR U3336 ( .A(n3038), .B(n3037), .Z(n3040) );
  XOR U3337 ( .A(n4098), .B(n3034), .Z(n3037) );
  XOR U3338 ( .A(n3032), .B(n3031), .Z(n3034) );
  XOR U3339 ( .A(n3029), .B(n3028), .Z(n3031) );
  XOR U3340 ( .A(n3025), .B(n3026), .Z(n3028) );
  AND U3341 ( .A(n4099), .B(n4100), .Z(n3026) );
  XOR U3342 ( .A(n3022), .B(n3023), .Z(n3025) );
  AND U3343 ( .A(n4101), .B(n4102), .Z(n3023) );
  XOR U3344 ( .A(n3019), .B(n3020), .Z(n3022) );
  AND U3345 ( .A(n4103), .B(n4104), .Z(n3020) );
  XOR U3346 ( .A(n3016), .B(n3017), .Z(n3019) );
  AND U3347 ( .A(n4105), .B(n4106), .Z(n3017) );
  XNOR U3348 ( .A(n2799), .B(n3014), .Z(n3016) );
  AND U3349 ( .A(n4107), .B(n4108), .Z(n3014) );
  XOR U3350 ( .A(n2801), .B(n2800), .Z(n2799) );
  AND U3351 ( .A(n4109), .B(n4110), .Z(n2800) );
  XOR U3352 ( .A(n2803), .B(n2802), .Z(n2801) );
  AND U3353 ( .A(n4111), .B(n4112), .Z(n2802) );
  XOR U3354 ( .A(n2805), .B(n2804), .Z(n2803) );
  AND U3355 ( .A(n4113), .B(n4114), .Z(n2804) );
  XOR U3356 ( .A(n2807), .B(n2806), .Z(n2805) );
  AND U3357 ( .A(n4115), .B(n4116), .Z(n2806) );
  XOR U3358 ( .A(n2809), .B(n2808), .Z(n2807) );
  AND U3359 ( .A(n4117), .B(n4118), .Z(n2808) );
  XOR U3360 ( .A(n2811), .B(n2810), .Z(n2809) );
  AND U3361 ( .A(n4119), .B(n4120), .Z(n2810) );
  XOR U3362 ( .A(n2813), .B(n2812), .Z(n2811) );
  AND U3363 ( .A(n4121), .B(n4122), .Z(n2812) );
  XOR U3364 ( .A(n2815), .B(n2814), .Z(n2813) );
  AND U3365 ( .A(n4123), .B(n4124), .Z(n2814) );
  XOR U3366 ( .A(n2817), .B(n2816), .Z(n2815) );
  AND U3367 ( .A(n4125), .B(n4126), .Z(n2816) );
  XOR U3368 ( .A(n2819), .B(n2818), .Z(n2817) );
  AND U3369 ( .A(n4127), .B(n4128), .Z(n2818) );
  XOR U3370 ( .A(n2821), .B(n2820), .Z(n2819) );
  AND U3371 ( .A(n4129), .B(n4130), .Z(n2820) );
  XOR U3372 ( .A(n2823), .B(n2822), .Z(n2821) );
  AND U3373 ( .A(n4131), .B(n4132), .Z(n2822) );
  XOR U3374 ( .A(n2825), .B(n2824), .Z(n2823) );
  AND U3375 ( .A(n4133), .B(n4134), .Z(n2824) );
  XOR U3376 ( .A(n2827), .B(n2826), .Z(n2825) );
  AND U3377 ( .A(n4135), .B(n4136), .Z(n2826) );
  XOR U3378 ( .A(n2829), .B(n2828), .Z(n2827) );
  AND U3379 ( .A(n4137), .B(n4138), .Z(n2828) );
  XOR U3380 ( .A(n2831), .B(n2830), .Z(n2829) );
  AND U3381 ( .A(n4139), .B(n4140), .Z(n2830) );
  XOR U3382 ( .A(n2833), .B(n2832), .Z(n2831) );
  AND U3383 ( .A(n4141), .B(n4142), .Z(n2832) );
  XOR U3384 ( .A(n2835), .B(n2834), .Z(n2833) );
  AND U3385 ( .A(n4143), .B(n4144), .Z(n2834) );
  XOR U3386 ( .A(n2837), .B(n2836), .Z(n2835) );
  AND U3387 ( .A(n4145), .B(n4146), .Z(n2836) );
  XOR U3388 ( .A(n2839), .B(n2838), .Z(n2837) );
  AND U3389 ( .A(n4147), .B(n4148), .Z(n2838) );
  XOR U3390 ( .A(n2841), .B(n2840), .Z(n2839) );
  AND U3391 ( .A(n4149), .B(n4150), .Z(n2840) );
  XOR U3392 ( .A(n2843), .B(n2842), .Z(n2841) );
  AND U3393 ( .A(n4151), .B(n4152), .Z(n2842) );
  XOR U3394 ( .A(n2845), .B(n2844), .Z(n2843) );
  AND U3395 ( .A(n4153), .B(n4154), .Z(n2844) );
  XOR U3396 ( .A(n2847), .B(n2846), .Z(n2845) );
  AND U3397 ( .A(n4155), .B(n4156), .Z(n2846) );
  XOR U3398 ( .A(n2849), .B(n2848), .Z(n2847) );
  AND U3399 ( .A(n4157), .B(n4158), .Z(n2848) );
  XOR U3400 ( .A(n2851), .B(n2850), .Z(n2849) );
  AND U3401 ( .A(n4159), .B(n4160), .Z(n2850) );
  XOR U3402 ( .A(n2853), .B(n2852), .Z(n2851) );
  AND U3403 ( .A(n4161), .B(n4162), .Z(n2852) );
  XOR U3404 ( .A(n2855), .B(n2854), .Z(n2853) );
  AND U3405 ( .A(n4163), .B(n4164), .Z(n2854) );
  XOR U3406 ( .A(n2857), .B(n2856), .Z(n2855) );
  AND U3407 ( .A(n4165), .B(n4166), .Z(n2856) );
  XOR U3408 ( .A(n2859), .B(n2858), .Z(n2857) );
  AND U3409 ( .A(n4167), .B(n4168), .Z(n2858) );
  XOR U3410 ( .A(n2861), .B(n2860), .Z(n2859) );
  AND U3411 ( .A(n4169), .B(n4170), .Z(n2860) );
  XOR U3412 ( .A(n2863), .B(n2862), .Z(n2861) );
  AND U3413 ( .A(n4171), .B(n4172), .Z(n2862) );
  XOR U3414 ( .A(n2865), .B(n2864), .Z(n2863) );
  AND U3415 ( .A(n4173), .B(n4174), .Z(n2864) );
  XOR U3416 ( .A(n2867), .B(n2866), .Z(n2865) );
  AND U3417 ( .A(n4175), .B(n4176), .Z(n2866) );
  XOR U3418 ( .A(n2869), .B(n2868), .Z(n2867) );
  AND U3419 ( .A(n4177), .B(n4178), .Z(n2868) );
  XOR U3420 ( .A(n2871), .B(n2870), .Z(n2869) );
  AND U3421 ( .A(n4179), .B(n4180), .Z(n2870) );
  XOR U3422 ( .A(n2873), .B(n2872), .Z(n2871) );
  AND U3423 ( .A(n4181), .B(n4182), .Z(n2872) );
  XOR U3424 ( .A(n2875), .B(n2874), .Z(n2873) );
  AND U3425 ( .A(n4183), .B(n4184), .Z(n2874) );
  XOR U3426 ( .A(n2877), .B(n2876), .Z(n2875) );
  AND U3427 ( .A(n4185), .B(n4186), .Z(n2876) );
  XOR U3428 ( .A(n3010), .B(n2878), .Z(n2877) );
  AND U3429 ( .A(n4187), .B(n4188), .Z(n2878) );
  XOR U3430 ( .A(n3012), .B(n3011), .Z(n3010) );
  AND U3431 ( .A(n4189), .B(n4190), .Z(n3011) );
  XOR U3432 ( .A(n2993), .B(n3013), .Z(n3012) );
  AND U3433 ( .A(n4191), .B(n4192), .Z(n3013) );
  XOR U3434 ( .A(n2995), .B(n2994), .Z(n2993) );
  AND U3435 ( .A(n4193), .B(n4194), .Z(n2994) );
  XOR U3436 ( .A(n2997), .B(n2996), .Z(n2995) );
  AND U3437 ( .A(n4195), .B(n4196), .Z(n2996) );
  XOR U3438 ( .A(n3001), .B(n2998), .Z(n2997) );
  AND U3439 ( .A(n4197), .B(n4198), .Z(n2998) );
  XOR U3440 ( .A(n3003), .B(n3002), .Z(n3001) );
  AND U3441 ( .A(n4199), .B(n4200), .Z(n3002) );
  XOR U3442 ( .A(n3006), .B(n3004), .Z(n3003) );
  AND U3443 ( .A(n4201), .B(n4202), .Z(n3004) );
  XOR U3444 ( .A(n3008), .B(n3007), .Z(n3006) );
  AND U3445 ( .A(n4203), .B(n4204), .Z(n3007) );
  XOR U3446 ( .A(n2893), .B(n3009), .Z(n3008) );
  AND U3447 ( .A(n4205), .B(n4206), .Z(n3009) );
  XNOR U3448 ( .A(n2900), .B(n2894), .Z(n2893) );
  AND U3449 ( .A(n4207), .B(n4208), .Z(n2894) );
  XOR U3450 ( .A(n2899), .B(n2891), .Z(n2900) );
  AND U3451 ( .A(n4209), .B(n4210), .Z(n2891) );
  XOR U3452 ( .A(n2992), .B(n2890), .Z(n2899) );
  AND U3453 ( .A(n4211), .B(n4212), .Z(n2890) );
  XNOR U3454 ( .A(n2911), .B(n2889), .Z(n2992) );
  AND U3455 ( .A(n4213), .B(n4214), .Z(n2889) );
  XNOR U3456 ( .A(n2918), .B(n2912), .Z(n2911) );
  AND U3457 ( .A(n4215), .B(n4216), .Z(n2912) );
  XOR U3458 ( .A(n2917), .B(n2909), .Z(n2918) );
  AND U3459 ( .A(n4217), .B(n4218), .Z(n2909) );
  XOR U3460 ( .A(n2991), .B(n2908), .Z(n2917) );
  AND U3461 ( .A(n4219), .B(n4220), .Z(n2908) );
  XNOR U3462 ( .A(n2929), .B(n2907), .Z(n2991) );
  AND U3463 ( .A(n4221), .B(n4222), .Z(n2907) );
  XNOR U3464 ( .A(n2936), .B(n2930), .Z(n2929) );
  AND U3465 ( .A(n4223), .B(n4224), .Z(n2930) );
  XOR U3466 ( .A(n2935), .B(n2927), .Z(n2936) );
  AND U3467 ( .A(n4225), .B(n4226), .Z(n2927) );
  XOR U3468 ( .A(n2990), .B(n2926), .Z(n2935) );
  AND U3469 ( .A(n4227), .B(n4228), .Z(n2926) );
  XNOR U3470 ( .A(n2947), .B(n2925), .Z(n2990) );
  AND U3471 ( .A(n4229), .B(n4230), .Z(n2925) );
  XNOR U3472 ( .A(n2954), .B(n2948), .Z(n2947) );
  AND U3473 ( .A(n4231), .B(n4232), .Z(n2948) );
  XOR U3474 ( .A(n2953), .B(n2945), .Z(n2954) );
  AND U3475 ( .A(n4233), .B(n4234), .Z(n2945) );
  XOR U3476 ( .A(n2989), .B(n2944), .Z(n2953) );
  AND U3477 ( .A(n4235), .B(n4236), .Z(n2944) );
  XNOR U3478 ( .A(n4237), .B(n4238), .Z(n2989) );
  XOR U3479 ( .A(n2987), .B(n2988), .Z(n4238) );
  AND U3480 ( .A(n4239), .B(n4240), .Z(n2988) );
  AND U3481 ( .A(n4241), .B(n4242), .Z(n2987) );
  XOR U3482 ( .A(n4243), .B(n2943), .Z(n4237) );
  AND U3483 ( .A(n4244), .B(n4245), .Z(n2943) );
  XOR U3484 ( .A(n4246), .B(n4247), .Z(n4243) );
  XOR U3485 ( .A(n4248), .B(n4249), .Z(n4247) );
  XOR U3486 ( .A(n2980), .B(n2981), .Z(n4249) );
  AND U3487 ( .A(n4250), .B(n4251), .Z(n2981) );
  AND U3488 ( .A(n4252), .B(n4253), .Z(n2980) );
  XOR U3489 ( .A(n2974), .B(n2979), .Z(n4248) );
  AND U3490 ( .A(n4254), .B(n4255), .Z(n2979) );
  AND U3491 ( .A(n4256), .B(n4257), .Z(n2974) );
  XOR U3492 ( .A(n4258), .B(n4259), .Z(n4246) );
  XOR U3493 ( .A(n2982), .B(n2985), .Z(n4259) );
  AND U3494 ( .A(n4260), .B(n4261), .Z(n2985) );
  AND U3495 ( .A(n4262), .B(n4263), .Z(n2982) );
  XOR U3496 ( .A(n4264), .B(n2986), .Z(n4258) );
  AND U3497 ( .A(n4265), .B(n4266), .Z(n2986) );
  XOR U3498 ( .A(n4267), .B(n4268), .Z(n4264) );
  XOR U3499 ( .A(n4269), .B(n4270), .Z(n4268) );
  XOR U3500 ( .A(n2967), .B(n2968), .Z(n4270) );
  AND U3501 ( .A(n4271), .B(n4272), .Z(n2968) );
  AND U3502 ( .A(n4273), .B(n4274), .Z(n2967) );
  XNOR U3503 ( .A(n2965), .B(n2964), .Z(n4269) );
  IV U3504 ( .A(n4275), .Z(n2964) );
  AND U3505 ( .A(n4276), .B(n4277), .Z(n4275) );
  AND U3506 ( .A(n4278), .B(n4279), .Z(n2965) );
  XOR U3507 ( .A(n4280), .B(n4281), .Z(n4267) );
  XOR U3508 ( .A(n2971), .B(n2972), .Z(n4281) );
  AND U3509 ( .A(n4282), .B(n4283), .Z(n2972) );
  AND U3510 ( .A(n4284), .B(n4285), .Z(n2971) );
  XOR U3511 ( .A(n2966), .B(n2973), .Z(n4280) );
  AND U3512 ( .A(n4286), .B(n4287), .Z(n2973) );
  XNOR U3513 ( .A(n4288), .B(n4289), .Z(n2966) );
  AND U3514 ( .A(n4290), .B(n4291), .Z(n4289) );
  NOR U3515 ( .A(n4292), .B(n4293), .Z(n4291) );
  NOR U3516 ( .A(n4294), .B(n4295), .Z(n4290) );
  AND U3517 ( .A(n4296), .B(n4297), .Z(n4295) );
  AND U3518 ( .A(n4298), .B(n4299), .Z(n4288) );
  NOR U3519 ( .A(n4300), .B(n4301), .Z(n4299) );
  AND U3520 ( .A(n4293), .B(n4302), .Z(n4301) );
  AND U3521 ( .A(n4294), .B(n4303), .Z(n4300) );
  NOR U3522 ( .A(n4304), .B(n4305), .Z(n4298) );
  XOR U3523 ( .A(n4306), .B(n4307), .Z(n4305) );
  AND U3524 ( .A(n4308), .B(n4309), .Z(n4307) );
  NOR U3525 ( .A(n4310), .B(n4311), .Z(n4309) );
  NOR U3526 ( .A(n4312), .B(n4313), .Z(n4308) );
  AND U3527 ( .A(n4314), .B(n4315), .Z(n4313) );
  AND U3528 ( .A(n4316), .B(n4317), .Z(n4306) );
  NOR U3529 ( .A(n4318), .B(n4319), .Z(n4317) );
  AND U3530 ( .A(n4311), .B(n4320), .Z(n4319) );
  AND U3531 ( .A(n4312), .B(n4321), .Z(n4318) );
  NOR U3532 ( .A(n4322), .B(n4323), .Z(n4316) );
  AND U3533 ( .A(n4324), .B(n4325), .Z(n4323) );
  AND U3534 ( .A(n4326), .B(n4327), .Z(n4325) );
  AND U3535 ( .A(n4328), .B(n4329), .Z(n4327) );
  NOR U3536 ( .A(n4330), .B(n4331), .Z(n4328) );
  NOR U3537 ( .A(n4332), .B(n4333), .Z(n4326) );
  AND U3538 ( .A(n4334), .B(n4335), .Z(n4324) );
  NOR U3539 ( .A(n4336), .B(n4337), .Z(n4335) );
  NOR U3540 ( .A(n4338), .B(n4339), .Z(n4334) );
  AND U3541 ( .A(n4310), .B(n4340), .Z(n4322) );
  AND U3542 ( .A(n4292), .B(n4341), .Z(n4304) );
  XOR U3543 ( .A(n4342), .B(n4343), .Z(n3029) );
  AND U3544 ( .A(n4342), .B(n4344), .Z(n4343) );
  XNOR U3545 ( .A(n4345), .B(n4346), .Z(n3032) );
  AND U3546 ( .A(n4345), .B(n4347), .Z(n4346) );
  IV U3547 ( .A(n3035), .Z(n4098) );
  XNOR U3548 ( .A(n4348), .B(n4349), .Z(n3035) );
  AND U3549 ( .A(n4348), .B(n4350), .Z(n4349) );
  XNOR U3550 ( .A(n4351), .B(n4352), .Z(n3038) );
  AND U3551 ( .A(n4351), .B(n4353), .Z(n4352) );
  XNOR U3552 ( .A(n4354), .B(n4355), .Z(n3041) );
  AND U3553 ( .A(n4356), .B(n4354), .Z(n4355) );
  XOR U3554 ( .A(n4357), .B(n4358), .Z(n3044) );
  NOR U3555 ( .A(n4359), .B(n4357), .Z(n4358) );
  XOR U3556 ( .A(n4360), .B(n4361), .Z(n3047) );
  NOR U3557 ( .A(n4362), .B(n4360), .Z(n4361) );
  XOR U3558 ( .A(n4363), .B(n4364), .Z(n3050) );
  NOR U3559 ( .A(n4365), .B(n4363), .Z(n4364) );
  XOR U3560 ( .A(n4366), .B(n4367), .Z(n3053) );
  NOR U3561 ( .A(n4368), .B(n4366), .Z(n4367) );
  XOR U3562 ( .A(n4369), .B(n4370), .Z(n3056) );
  NOR U3563 ( .A(n4371), .B(n4369), .Z(n4370) );
  XOR U3564 ( .A(n4372), .B(n4373), .Z(n3059) );
  NOR U3565 ( .A(n4374), .B(n4372), .Z(n4373) );
  XOR U3566 ( .A(n4375), .B(n4376), .Z(n3062) );
  NOR U3567 ( .A(n4377), .B(n4375), .Z(n4376) );
  XOR U3568 ( .A(n4378), .B(n4379), .Z(n3065) );
  NOR U3569 ( .A(n4380), .B(n4378), .Z(n4379) );
  XOR U3570 ( .A(n4381), .B(n4382), .Z(n3068) );
  NOR U3571 ( .A(n4383), .B(n4381), .Z(n4382) );
  XOR U3572 ( .A(n4384), .B(n4385), .Z(n3071) );
  NOR U3573 ( .A(n4386), .B(n4384), .Z(n4385) );
  XOR U3574 ( .A(n4387), .B(n4388), .Z(n3074) );
  NOR U3575 ( .A(n4389), .B(n4387), .Z(n4388) );
  XOR U3576 ( .A(n4390), .B(n4391), .Z(n3077) );
  NOR U3577 ( .A(n4392), .B(n4390), .Z(n4391) );
  XOR U3578 ( .A(n4393), .B(n4394), .Z(n3080) );
  NOR U3579 ( .A(n4395), .B(n4393), .Z(n4394) );
  XOR U3580 ( .A(n4396), .B(n4397), .Z(n3083) );
  NOR U3581 ( .A(n4398), .B(n4396), .Z(n4397) );
  XOR U3582 ( .A(n4399), .B(n4400), .Z(n3086) );
  NOR U3583 ( .A(n4401), .B(n4399), .Z(n4400) );
  XOR U3584 ( .A(n4402), .B(n4403), .Z(n3089) );
  NOR U3585 ( .A(n4404), .B(n4402), .Z(n4403) );
  XOR U3586 ( .A(n4405), .B(n4406), .Z(n3092) );
  NOR U3587 ( .A(n4407), .B(n4405), .Z(n4406) );
  XOR U3588 ( .A(n4408), .B(n4409), .Z(n3095) );
  NOR U3589 ( .A(n4410), .B(n4408), .Z(n4409) );
  XOR U3590 ( .A(n4411), .B(n4412), .Z(n3098) );
  NOR U3591 ( .A(n4413), .B(n4411), .Z(n4412) );
  XOR U3592 ( .A(n4414), .B(n4415), .Z(n3101) );
  NOR U3593 ( .A(n4416), .B(n4414), .Z(n4415) );
  XOR U3594 ( .A(n4417), .B(n4418), .Z(n3104) );
  NOR U3595 ( .A(n4419), .B(n4417), .Z(n4418) );
  XOR U3596 ( .A(n4420), .B(n4421), .Z(n3107) );
  NOR U3597 ( .A(n4422), .B(n4420), .Z(n4421) );
  XOR U3598 ( .A(n4423), .B(n4424), .Z(n3110) );
  NOR U3599 ( .A(n4425), .B(n4423), .Z(n4424) );
  XOR U3600 ( .A(n4426), .B(n4427), .Z(n3113) );
  NOR U3601 ( .A(n4428), .B(n4426), .Z(n4427) );
  XOR U3602 ( .A(n4429), .B(n4430), .Z(n3116) );
  NOR U3603 ( .A(n4431), .B(n4429), .Z(n4430) );
  XOR U3604 ( .A(n4432), .B(n4433), .Z(n3119) );
  NOR U3605 ( .A(n4434), .B(n4432), .Z(n4433) );
  XOR U3606 ( .A(n4435), .B(n4436), .Z(n3122) );
  NOR U3607 ( .A(n4437), .B(n4435), .Z(n4436) );
  XOR U3608 ( .A(n4438), .B(n4439), .Z(n3125) );
  NOR U3609 ( .A(n4440), .B(n4438), .Z(n4439) );
  XOR U3610 ( .A(n4441), .B(n4442), .Z(n3128) );
  NOR U3611 ( .A(n4443), .B(n4441), .Z(n4442) );
  XOR U3612 ( .A(n4444), .B(n4445), .Z(n3131) );
  NOR U3613 ( .A(n4446), .B(n4444), .Z(n4445) );
  XOR U3614 ( .A(n4447), .B(n4448), .Z(n3134) );
  NOR U3615 ( .A(n4449), .B(n4447), .Z(n4448) );
  XOR U3616 ( .A(n4450), .B(n4451), .Z(n3137) );
  NOR U3617 ( .A(n4452), .B(n4450), .Z(n4451) );
  XOR U3618 ( .A(n4453), .B(n4454), .Z(n3140) );
  NOR U3619 ( .A(n4455), .B(n4453), .Z(n4454) );
  XOR U3620 ( .A(n4456), .B(n4457), .Z(n3143) );
  NOR U3621 ( .A(n4458), .B(n4456), .Z(n4457) );
  XOR U3622 ( .A(n4459), .B(n4460), .Z(n3146) );
  NOR U3623 ( .A(n4461), .B(n4459), .Z(n4460) );
  XOR U3624 ( .A(n4462), .B(n4463), .Z(n3149) );
  NOR U3625 ( .A(n4464), .B(n4462), .Z(n4463) );
  XOR U3626 ( .A(n4465), .B(n4466), .Z(n3152) );
  NOR U3627 ( .A(n4467), .B(n4465), .Z(n4466) );
  XOR U3628 ( .A(n4468), .B(n4469), .Z(n3155) );
  NOR U3629 ( .A(n4470), .B(n4468), .Z(n4469) );
  XOR U3630 ( .A(n4471), .B(n4472), .Z(n3158) );
  NOR U3631 ( .A(n4473), .B(n4471), .Z(n4472) );
  XOR U3632 ( .A(n4474), .B(n4475), .Z(n3161) );
  NOR U3633 ( .A(n4476), .B(n4474), .Z(n4475) );
  XOR U3634 ( .A(n4477), .B(n4478), .Z(n3164) );
  NOR U3635 ( .A(n4479), .B(n4477), .Z(n4478) );
  XOR U3636 ( .A(n4480), .B(n4481), .Z(n3167) );
  NOR U3637 ( .A(n4482), .B(n4480), .Z(n4481) );
  XOR U3638 ( .A(n4483), .B(n4484), .Z(n3170) );
  NOR U3639 ( .A(n4485), .B(n4483), .Z(n4484) );
  XOR U3640 ( .A(n4486), .B(n4487), .Z(n3173) );
  NOR U3641 ( .A(n4488), .B(n4486), .Z(n4487) );
  XOR U3642 ( .A(n4489), .B(n4490), .Z(n3176) );
  NOR U3643 ( .A(n4491), .B(n4489), .Z(n4490) );
  XOR U3644 ( .A(n4492), .B(n4493), .Z(n3179) );
  NOR U3645 ( .A(n4494), .B(n4492), .Z(n4493) );
  XOR U3646 ( .A(n4495), .B(n4496), .Z(n3182) );
  NOR U3647 ( .A(n4497), .B(n4495), .Z(n4496) );
  XOR U3648 ( .A(n4498), .B(n4499), .Z(n3185) );
  NOR U3649 ( .A(n4500), .B(n4498), .Z(n4499) );
  XOR U3650 ( .A(n4501), .B(n4502), .Z(n3188) );
  NOR U3651 ( .A(n4503), .B(n4501), .Z(n4502) );
  XOR U3652 ( .A(n4504), .B(n4505), .Z(n3191) );
  NOR U3653 ( .A(n4506), .B(n4504), .Z(n4505) );
  XOR U3654 ( .A(n4507), .B(n4508), .Z(n3194) );
  NOR U3655 ( .A(n4509), .B(n4507), .Z(n4508) );
  XOR U3656 ( .A(n4510), .B(n4511), .Z(n3197) );
  NOR U3657 ( .A(n4512), .B(n4510), .Z(n4511) );
  XOR U3658 ( .A(n4513), .B(n4514), .Z(n3200) );
  NOR U3659 ( .A(n4515), .B(n4513), .Z(n4514) );
  XOR U3660 ( .A(n4516), .B(n4517), .Z(n3203) );
  NOR U3661 ( .A(n4518), .B(n4516), .Z(n4517) );
  XOR U3662 ( .A(n4519), .B(n4520), .Z(n3206) );
  NOR U3663 ( .A(n4521), .B(n4519), .Z(n4520) );
  XOR U3664 ( .A(n4522), .B(n4523), .Z(n3209) );
  NOR U3665 ( .A(n4524), .B(n4522), .Z(n4523) );
  XOR U3666 ( .A(n4525), .B(n4526), .Z(n3212) );
  NOR U3667 ( .A(n4527), .B(n4525), .Z(n4526) );
  XOR U3668 ( .A(n4528), .B(n4529), .Z(n3215) );
  NOR U3669 ( .A(n4530), .B(n4528), .Z(n4529) );
  XOR U3670 ( .A(n4531), .B(n4532), .Z(n3218) );
  NOR U3671 ( .A(n4533), .B(n4531), .Z(n4532) );
  XOR U3672 ( .A(n4534), .B(n4535), .Z(n3221) );
  NOR U3673 ( .A(n4536), .B(n4534), .Z(n4535) );
  XOR U3674 ( .A(n4537), .B(n4538), .Z(n3224) );
  NOR U3675 ( .A(n4539), .B(n4537), .Z(n4538) );
  XOR U3676 ( .A(n4540), .B(n4541), .Z(n3227) );
  NOR U3677 ( .A(n4542), .B(n4540), .Z(n4541) );
  XOR U3678 ( .A(n4543), .B(n4544), .Z(n3230) );
  NOR U3679 ( .A(n4545), .B(n4543), .Z(n4544) );
  XOR U3680 ( .A(n4546), .B(n4547), .Z(n3233) );
  NOR U3681 ( .A(n4548), .B(n4546), .Z(n4547) );
  XOR U3682 ( .A(n4549), .B(n4550), .Z(n3236) );
  NOR U3683 ( .A(n4551), .B(n4549), .Z(n4550) );
  XOR U3684 ( .A(n4552), .B(n4553), .Z(n3239) );
  NOR U3685 ( .A(n4554), .B(n4552), .Z(n4553) );
  XOR U3686 ( .A(n4555), .B(n4556), .Z(n3242) );
  NOR U3687 ( .A(n4557), .B(n4555), .Z(n4556) );
  XOR U3688 ( .A(n4558), .B(n4559), .Z(n3245) );
  NOR U3689 ( .A(n4560), .B(n4558), .Z(n4559) );
  XOR U3690 ( .A(n4561), .B(n4562), .Z(n3248) );
  NOR U3691 ( .A(n4563), .B(n4561), .Z(n4562) );
  XOR U3692 ( .A(n4564), .B(n4565), .Z(n3251) );
  NOR U3693 ( .A(n4566), .B(n4564), .Z(n4565) );
  XOR U3694 ( .A(n4567), .B(n4568), .Z(n3254) );
  NOR U3695 ( .A(n4569), .B(n4567), .Z(n4568) );
  XOR U3696 ( .A(n4570), .B(n4571), .Z(n3257) );
  NOR U3697 ( .A(n4572), .B(n4570), .Z(n4571) );
  XOR U3698 ( .A(n4573), .B(n4574), .Z(n3260) );
  NOR U3699 ( .A(n4575), .B(n4573), .Z(n4574) );
  XOR U3700 ( .A(n4576), .B(n4577), .Z(n3263) );
  NOR U3701 ( .A(n4578), .B(n4576), .Z(n4577) );
  XOR U3702 ( .A(n4579), .B(n4580), .Z(n3266) );
  NOR U3703 ( .A(n4581), .B(n4579), .Z(n4580) );
  XOR U3704 ( .A(n4582), .B(n4583), .Z(n3269) );
  NOR U3705 ( .A(n4584), .B(n4582), .Z(n4583) );
  XOR U3706 ( .A(n4585), .B(n4586), .Z(n3272) );
  NOR U3707 ( .A(n4587), .B(n4585), .Z(n4586) );
  XOR U3708 ( .A(n4588), .B(n4589), .Z(n3275) );
  NOR U3709 ( .A(n4590), .B(n4588), .Z(n4589) );
  XOR U3710 ( .A(n4591), .B(n4592), .Z(n3278) );
  NOR U3711 ( .A(n4593), .B(n4591), .Z(n4592) );
  XOR U3712 ( .A(n4594), .B(n4595), .Z(n3281) );
  NOR U3713 ( .A(n4596), .B(n4594), .Z(n4595) );
  XOR U3714 ( .A(n4597), .B(n4598), .Z(n3284) );
  NOR U3715 ( .A(n4599), .B(n4597), .Z(n4598) );
  XOR U3716 ( .A(n4600), .B(n4601), .Z(n3287) );
  NOR U3717 ( .A(n4602), .B(n4600), .Z(n4601) );
  XOR U3718 ( .A(n4603), .B(n4604), .Z(n3290) );
  NOR U3719 ( .A(n4605), .B(n4603), .Z(n4604) );
  XOR U3720 ( .A(n4606), .B(n4607), .Z(n3293) );
  NOR U3721 ( .A(n4608), .B(n4606), .Z(n4607) );
  XOR U3722 ( .A(n4609), .B(n4610), .Z(n3296) );
  NOR U3723 ( .A(n4611), .B(n4609), .Z(n4610) );
  XOR U3724 ( .A(n4612), .B(n4613), .Z(n3299) );
  NOR U3725 ( .A(n4614), .B(n4612), .Z(n4613) );
  XOR U3726 ( .A(n4615), .B(n4616), .Z(n3302) );
  NOR U3727 ( .A(n4617), .B(n4615), .Z(n4616) );
  XOR U3728 ( .A(n4618), .B(n4619), .Z(n3305) );
  NOR U3729 ( .A(n4620), .B(n4618), .Z(n4619) );
  XOR U3730 ( .A(n4621), .B(n4622), .Z(n3308) );
  NOR U3731 ( .A(n4623), .B(n4621), .Z(n4622) );
  XOR U3732 ( .A(n4624), .B(n4625), .Z(n3311) );
  NOR U3733 ( .A(n4626), .B(n4624), .Z(n4625) );
  XOR U3734 ( .A(n4627), .B(n4628), .Z(n3314) );
  NOR U3735 ( .A(n4629), .B(n4627), .Z(n4628) );
  XOR U3736 ( .A(n4630), .B(n4631), .Z(n3317) );
  NOR U3737 ( .A(n4632), .B(n4630), .Z(n4631) );
  XOR U3738 ( .A(n4633), .B(n4634), .Z(n3320) );
  NOR U3739 ( .A(n4635), .B(n4633), .Z(n4634) );
  XOR U3740 ( .A(n4636), .B(n4637), .Z(n3323) );
  NOR U3741 ( .A(n4638), .B(n4636), .Z(n4637) );
  XOR U3742 ( .A(n4639), .B(n4640), .Z(n3326) );
  NOR U3743 ( .A(n4641), .B(n4639), .Z(n4640) );
  XOR U3744 ( .A(n4642), .B(n4643), .Z(n3329) );
  NOR U3745 ( .A(n4644), .B(n4642), .Z(n4643) );
  XOR U3746 ( .A(n4645), .B(n4646), .Z(n3332) );
  NOR U3747 ( .A(n4647), .B(n4645), .Z(n4646) );
  XOR U3748 ( .A(n4648), .B(n4649), .Z(n3335) );
  NOR U3749 ( .A(n4650), .B(n4648), .Z(n4649) );
  XOR U3750 ( .A(n4651), .B(n4652), .Z(n3338) );
  NOR U3751 ( .A(n4653), .B(n4651), .Z(n4652) );
  XOR U3752 ( .A(n4654), .B(n4655), .Z(n3341) );
  NOR U3753 ( .A(n4656), .B(n4654), .Z(n4655) );
  XOR U3754 ( .A(n4657), .B(n4658), .Z(n3344) );
  NOR U3755 ( .A(n4659), .B(n4657), .Z(n4658) );
  XOR U3756 ( .A(n4660), .B(n4661), .Z(n3347) );
  NOR U3757 ( .A(n4662), .B(n4660), .Z(n4661) );
  XOR U3758 ( .A(n4663), .B(n4664), .Z(n3350) );
  NOR U3759 ( .A(n4665), .B(n4663), .Z(n4664) );
  XOR U3760 ( .A(n4666), .B(n4667), .Z(n3353) );
  NOR U3761 ( .A(n4668), .B(n4666), .Z(n4667) );
  XOR U3762 ( .A(n4669), .B(n4670), .Z(n3356) );
  NOR U3763 ( .A(n4671), .B(n4669), .Z(n4670) );
  XOR U3764 ( .A(n4672), .B(n4673), .Z(n3359) );
  NOR U3765 ( .A(n4674), .B(n4672), .Z(n4673) );
  XOR U3766 ( .A(n4675), .B(n4676), .Z(n3362) );
  NOR U3767 ( .A(n4677), .B(n4675), .Z(n4676) );
  XOR U3768 ( .A(n4678), .B(n4679), .Z(n3365) );
  NOR U3769 ( .A(n4680), .B(n4678), .Z(n4679) );
  XOR U3770 ( .A(n4681), .B(n4682), .Z(n3368) );
  NOR U3771 ( .A(n4683), .B(n4681), .Z(n4682) );
  XOR U3772 ( .A(n4684), .B(n4685), .Z(n3371) );
  NOR U3773 ( .A(n4686), .B(n4684), .Z(n4685) );
  XOR U3774 ( .A(n4687), .B(n4688), .Z(n3374) );
  NOR U3775 ( .A(n4689), .B(n4687), .Z(n4688) );
  XOR U3776 ( .A(n4690), .B(n4691), .Z(n3377) );
  NOR U3777 ( .A(n4692), .B(n4690), .Z(n4691) );
  XOR U3778 ( .A(n4693), .B(n4694), .Z(n3380) );
  NOR U3779 ( .A(n4695), .B(n4693), .Z(n4694) );
  XOR U3780 ( .A(n4696), .B(n4697), .Z(n3383) );
  NOR U3781 ( .A(n4698), .B(n4696), .Z(n4697) );
  XOR U3782 ( .A(n4699), .B(n4700), .Z(n3386) );
  NOR U3783 ( .A(n4701), .B(n4699), .Z(n4700) );
  XOR U3784 ( .A(n4702), .B(n4703), .Z(n3389) );
  NOR U3785 ( .A(n4704), .B(n4702), .Z(n4703) );
  XOR U3786 ( .A(n4705), .B(n4706), .Z(n3392) );
  NOR U3787 ( .A(n4707), .B(n4705), .Z(n4706) );
  XOR U3788 ( .A(n4708), .B(n4709), .Z(n3395) );
  NOR U3789 ( .A(n4710), .B(n4708), .Z(n4709) );
  XOR U3790 ( .A(n4711), .B(n4712), .Z(n3398) );
  NOR U3791 ( .A(n4713), .B(n4711), .Z(n4712) );
  XOR U3792 ( .A(n4714), .B(n4715), .Z(n3401) );
  NOR U3793 ( .A(n4716), .B(n4714), .Z(n4715) );
  XOR U3794 ( .A(n4717), .B(n4718), .Z(n3404) );
  NOR U3795 ( .A(n4719), .B(n4717), .Z(n4718) );
  XOR U3796 ( .A(n4720), .B(n4721), .Z(n3407) );
  NOR U3797 ( .A(n4722), .B(n4720), .Z(n4721) );
  XOR U3798 ( .A(n4723), .B(n4724), .Z(n3410) );
  NOR U3799 ( .A(n4725), .B(n4723), .Z(n4724) );
  XOR U3800 ( .A(n4726), .B(n4727), .Z(n3413) );
  NOR U3801 ( .A(n4728), .B(n4726), .Z(n4727) );
  XOR U3802 ( .A(n4729), .B(n4730), .Z(n3416) );
  NOR U3803 ( .A(n4731), .B(n4729), .Z(n4730) );
  XOR U3804 ( .A(n4732), .B(n4733), .Z(n3419) );
  NOR U3805 ( .A(n4734), .B(n4732), .Z(n4733) );
  XOR U3806 ( .A(n4735), .B(n4736), .Z(n3422) );
  NOR U3807 ( .A(n4737), .B(n4735), .Z(n4736) );
  XOR U3808 ( .A(n4738), .B(n4739), .Z(n3425) );
  NOR U3809 ( .A(n4740), .B(n4738), .Z(n4739) );
  XOR U3810 ( .A(n4741), .B(n4742), .Z(n3428) );
  NOR U3811 ( .A(n4743), .B(n4741), .Z(n4742) );
  XOR U3812 ( .A(n4744), .B(n4745), .Z(n3431) );
  NOR U3813 ( .A(n4746), .B(n4744), .Z(n4745) );
  XOR U3814 ( .A(n4747), .B(n4748), .Z(n3434) );
  NOR U3815 ( .A(n4749), .B(n4747), .Z(n4748) );
  XOR U3816 ( .A(n4750), .B(n4751), .Z(n3437) );
  NOR U3817 ( .A(n4752), .B(n4750), .Z(n4751) );
  XOR U3818 ( .A(n4753), .B(n4754), .Z(n3440) );
  AND U3819 ( .A(n4755), .B(n4753), .Z(n4754) );
  XOR U3820 ( .A(n4756), .B(n4757), .Z(n3443) );
  AND U3821 ( .A(n88), .B(n4756), .Z(n4757) );
  XNOR U3822 ( .A(n4758), .B(n4094), .Z(n4096) );
  IV U3823 ( .A(n71), .Z(n4758) );
  XOR U3824 ( .A(n4091), .B(n4090), .Z(n71) );
  XNOR U3825 ( .A(n4088), .B(n4087), .Z(n4090) );
  XNOR U3826 ( .A(n4085), .B(n4084), .Z(n4087) );
  XNOR U3827 ( .A(n4082), .B(n4081), .Z(n4084) );
  XNOR U3828 ( .A(n4079), .B(n4078), .Z(n4081) );
  XNOR U3829 ( .A(n4076), .B(n4075), .Z(n4078) );
  XNOR U3830 ( .A(n4073), .B(n4072), .Z(n4075) );
  XNOR U3831 ( .A(n4070), .B(n4069), .Z(n4072) );
  XNOR U3832 ( .A(n4067), .B(n4066), .Z(n4069) );
  XNOR U3833 ( .A(n4064), .B(n4063), .Z(n4066) );
  XNOR U3834 ( .A(n4061), .B(n4060), .Z(n4063) );
  XNOR U3835 ( .A(n4058), .B(n4057), .Z(n4060) );
  XNOR U3836 ( .A(n4055), .B(n4054), .Z(n4057) );
  XNOR U3837 ( .A(n4052), .B(n4051), .Z(n4054) );
  XNOR U3838 ( .A(n4049), .B(n4048), .Z(n4051) );
  XNOR U3839 ( .A(n4046), .B(n4045), .Z(n4048) );
  XNOR U3840 ( .A(n4043), .B(n4042), .Z(n4045) );
  XNOR U3841 ( .A(n4040), .B(n4039), .Z(n4042) );
  XNOR U3842 ( .A(n4037), .B(n4036), .Z(n4039) );
  XNOR U3843 ( .A(n4034), .B(n4033), .Z(n4036) );
  XNOR U3844 ( .A(n4031), .B(n4030), .Z(n4033) );
  XNOR U3845 ( .A(n4028), .B(n4027), .Z(n4030) );
  XNOR U3846 ( .A(n4025), .B(n4024), .Z(n4027) );
  XNOR U3847 ( .A(n4022), .B(n4021), .Z(n4024) );
  XNOR U3848 ( .A(n4019), .B(n4018), .Z(n4021) );
  XNOR U3849 ( .A(n4016), .B(n4015), .Z(n4018) );
  XNOR U3850 ( .A(n4013), .B(n4012), .Z(n4015) );
  XNOR U3851 ( .A(n4010), .B(n4009), .Z(n4012) );
  XNOR U3852 ( .A(n4007), .B(n4006), .Z(n4009) );
  XNOR U3853 ( .A(n4004), .B(n4003), .Z(n4006) );
  XNOR U3854 ( .A(n4001), .B(n4000), .Z(n4003) );
  XNOR U3855 ( .A(n3998), .B(n3997), .Z(n4000) );
  XNOR U3856 ( .A(n3995), .B(n3994), .Z(n3997) );
  XNOR U3857 ( .A(n3992), .B(n3991), .Z(n3994) );
  XNOR U3858 ( .A(n3989), .B(n3988), .Z(n3991) );
  XNOR U3859 ( .A(n3986), .B(n3985), .Z(n3988) );
  XNOR U3860 ( .A(n3983), .B(n3982), .Z(n3985) );
  XNOR U3861 ( .A(n3980), .B(n3979), .Z(n3982) );
  XNOR U3862 ( .A(n3977), .B(n3976), .Z(n3979) );
  XNOR U3863 ( .A(n3974), .B(n3973), .Z(n3976) );
  XNOR U3864 ( .A(n3971), .B(n3970), .Z(n3973) );
  XNOR U3865 ( .A(n3968), .B(n3967), .Z(n3970) );
  XNOR U3866 ( .A(n3965), .B(n3964), .Z(n3967) );
  XNOR U3867 ( .A(n3962), .B(n3961), .Z(n3964) );
  XNOR U3868 ( .A(n3959), .B(n3958), .Z(n3961) );
  XNOR U3869 ( .A(n3956), .B(n3955), .Z(n3958) );
  XNOR U3870 ( .A(n3953), .B(n3952), .Z(n3955) );
  XNOR U3871 ( .A(n3950), .B(n3949), .Z(n3952) );
  XNOR U3872 ( .A(n3947), .B(n3946), .Z(n3949) );
  XNOR U3873 ( .A(n3944), .B(n3943), .Z(n3946) );
  XNOR U3874 ( .A(n3941), .B(n3940), .Z(n3943) );
  XNOR U3875 ( .A(n3938), .B(n3937), .Z(n3940) );
  XNOR U3876 ( .A(n3935), .B(n3934), .Z(n3937) );
  XNOR U3877 ( .A(n3932), .B(n3931), .Z(n3934) );
  XNOR U3878 ( .A(n3929), .B(n3928), .Z(n3931) );
  XNOR U3879 ( .A(n3926), .B(n3925), .Z(n3928) );
  XNOR U3880 ( .A(n3923), .B(n3922), .Z(n3925) );
  XNOR U3881 ( .A(n3920), .B(n3919), .Z(n3922) );
  XNOR U3882 ( .A(n3917), .B(n3916), .Z(n3919) );
  XNOR U3883 ( .A(n3914), .B(n3913), .Z(n3916) );
  XNOR U3884 ( .A(n3911), .B(n3910), .Z(n3913) );
  XNOR U3885 ( .A(n3908), .B(n3907), .Z(n3910) );
  XNOR U3886 ( .A(n3905), .B(n3904), .Z(n3907) );
  XNOR U3887 ( .A(n3902), .B(n3901), .Z(n3904) );
  XNOR U3888 ( .A(n3899), .B(n3898), .Z(n3901) );
  XNOR U3889 ( .A(n3896), .B(n3895), .Z(n3898) );
  XNOR U3890 ( .A(n3893), .B(n3892), .Z(n3895) );
  XNOR U3891 ( .A(n3890), .B(n3889), .Z(n3892) );
  XNOR U3892 ( .A(n3887), .B(n3886), .Z(n3889) );
  XNOR U3893 ( .A(n3884), .B(n3883), .Z(n3886) );
  XNOR U3894 ( .A(n3881), .B(n3880), .Z(n3883) );
  XNOR U3895 ( .A(n3878), .B(n3877), .Z(n3880) );
  XNOR U3896 ( .A(n3875), .B(n3874), .Z(n3877) );
  XNOR U3897 ( .A(n3872), .B(n3871), .Z(n3874) );
  XNOR U3898 ( .A(n3869), .B(n3868), .Z(n3871) );
  XNOR U3899 ( .A(n3866), .B(n3865), .Z(n3868) );
  XNOR U3900 ( .A(n3863), .B(n3862), .Z(n3865) );
  XNOR U3901 ( .A(n3860), .B(n3859), .Z(n3862) );
  XNOR U3902 ( .A(n3857), .B(n3856), .Z(n3859) );
  XNOR U3903 ( .A(n3854), .B(n3853), .Z(n3856) );
  XNOR U3904 ( .A(n3851), .B(n3850), .Z(n3853) );
  XNOR U3905 ( .A(n3848), .B(n3847), .Z(n3850) );
  XNOR U3906 ( .A(n3845), .B(n3844), .Z(n3847) );
  XNOR U3907 ( .A(n3842), .B(n3841), .Z(n3844) );
  XNOR U3908 ( .A(n3839), .B(n3838), .Z(n3841) );
  XNOR U3909 ( .A(n3836), .B(n3835), .Z(n3838) );
  XNOR U3910 ( .A(n3833), .B(n3832), .Z(n3835) );
  XNOR U3911 ( .A(n3830), .B(n3829), .Z(n3832) );
  XNOR U3912 ( .A(n3827), .B(n3826), .Z(n3829) );
  XNOR U3913 ( .A(n3824), .B(n3823), .Z(n3826) );
  XNOR U3914 ( .A(n3821), .B(n3820), .Z(n3823) );
  XNOR U3915 ( .A(n3818), .B(n3817), .Z(n3820) );
  XNOR U3916 ( .A(n3815), .B(n3814), .Z(n3817) );
  XNOR U3917 ( .A(n3812), .B(n3811), .Z(n3814) );
  XNOR U3918 ( .A(n3809), .B(n3808), .Z(n3811) );
  XNOR U3919 ( .A(n3806), .B(n3805), .Z(n3808) );
  XNOR U3920 ( .A(n3803), .B(n3802), .Z(n3805) );
  XNOR U3921 ( .A(n3800), .B(n3799), .Z(n3802) );
  XNOR U3922 ( .A(n3797), .B(n3796), .Z(n3799) );
  XNOR U3923 ( .A(n3794), .B(n3793), .Z(n3796) );
  XNOR U3924 ( .A(n3791), .B(n3790), .Z(n3793) );
  XNOR U3925 ( .A(n3788), .B(n3787), .Z(n3790) );
  XNOR U3926 ( .A(n3785), .B(n3784), .Z(n3787) );
  XNOR U3927 ( .A(n3782), .B(n3781), .Z(n3784) );
  XNOR U3928 ( .A(n3779), .B(n3778), .Z(n3781) );
  XNOR U3929 ( .A(n3776), .B(n3775), .Z(n3778) );
  XNOR U3930 ( .A(n3773), .B(n3772), .Z(n3775) );
  XNOR U3931 ( .A(n3770), .B(n3769), .Z(n3772) );
  XNOR U3932 ( .A(n3767), .B(n3766), .Z(n3769) );
  XNOR U3933 ( .A(n3764), .B(n3763), .Z(n3766) );
  XNOR U3934 ( .A(n3761), .B(n3760), .Z(n3763) );
  XNOR U3935 ( .A(n3758), .B(n3757), .Z(n3760) );
  XNOR U3936 ( .A(n3755), .B(n3754), .Z(n3757) );
  XNOR U3937 ( .A(n3752), .B(n3751), .Z(n3754) );
  XNOR U3938 ( .A(n3749), .B(n3748), .Z(n3751) );
  XNOR U3939 ( .A(n3746), .B(n3745), .Z(n3748) );
  XNOR U3940 ( .A(n3743), .B(n3742), .Z(n3745) );
  XNOR U3941 ( .A(n3740), .B(n3739), .Z(n3742) );
  XNOR U3942 ( .A(n3737), .B(n3736), .Z(n3739) );
  XNOR U3943 ( .A(n3734), .B(n3733), .Z(n3736) );
  XNOR U3944 ( .A(n3731), .B(n3730), .Z(n3733) );
  XNOR U3945 ( .A(n3728), .B(n3727), .Z(n3730) );
  XNOR U3946 ( .A(n3725), .B(n3724), .Z(n3727) );
  XNOR U3947 ( .A(n3722), .B(n3721), .Z(n3724) );
  XNOR U3948 ( .A(n3719), .B(n3718), .Z(n3721) );
  XNOR U3949 ( .A(n3716), .B(n3715), .Z(n3718) );
  XNOR U3950 ( .A(n3713), .B(n3712), .Z(n3715) );
  XNOR U3951 ( .A(n3710), .B(n3709), .Z(n3712) );
  XNOR U3952 ( .A(n3707), .B(n3706), .Z(n3709) );
  XNOR U3953 ( .A(n3704), .B(n3703), .Z(n3706) );
  XNOR U3954 ( .A(n3701), .B(n3700), .Z(n3703) );
  XNOR U3955 ( .A(n3698), .B(n3697), .Z(n3700) );
  XNOR U3956 ( .A(n3695), .B(n3694), .Z(n3697) );
  XNOR U3957 ( .A(n3692), .B(n3691), .Z(n3694) );
  XNOR U3958 ( .A(n3689), .B(n3688), .Z(n3691) );
  XNOR U3959 ( .A(n3686), .B(n3685), .Z(n3688) );
  XOR U3960 ( .A(n4759), .B(n3682), .Z(n3685) );
  XOR U3961 ( .A(n3680), .B(n3679), .Z(n3682) );
  XOR U3962 ( .A(n3677), .B(n3676), .Z(n3679) );
  XOR U3963 ( .A(n3673), .B(n3674), .Z(n3676) );
  AND U3964 ( .A(n4760), .B(n4761), .Z(n3674) );
  XOR U3965 ( .A(n3670), .B(n3671), .Z(n3673) );
  AND U3966 ( .A(n4762), .B(n4763), .Z(n3671) );
  XOR U3967 ( .A(n3667), .B(n3668), .Z(n3670) );
  AND U3968 ( .A(n4764), .B(n4765), .Z(n3668) );
  XOR U3969 ( .A(n3664), .B(n3665), .Z(n3667) );
  AND U3970 ( .A(n4766), .B(n4767), .Z(n3665) );
  XNOR U3971 ( .A(n3447), .B(n3662), .Z(n3664) );
  AND U3972 ( .A(n4768), .B(n4769), .Z(n3662) );
  XOR U3973 ( .A(n3449), .B(n3448), .Z(n3447) );
  AND U3974 ( .A(n4770), .B(n4771), .Z(n3448) );
  XOR U3975 ( .A(n3451), .B(n3450), .Z(n3449) );
  AND U3976 ( .A(n4772), .B(n4773), .Z(n3450) );
  XOR U3977 ( .A(n3453), .B(n3452), .Z(n3451) );
  AND U3978 ( .A(n4774), .B(n4775), .Z(n3452) );
  XOR U3979 ( .A(n3455), .B(n3454), .Z(n3453) );
  AND U3980 ( .A(n4776), .B(n4777), .Z(n3454) );
  XOR U3981 ( .A(n3457), .B(n3456), .Z(n3455) );
  AND U3982 ( .A(n4778), .B(n4779), .Z(n3456) );
  XOR U3983 ( .A(n3459), .B(n3458), .Z(n3457) );
  AND U3984 ( .A(n4780), .B(n4781), .Z(n3458) );
  XOR U3985 ( .A(n3461), .B(n3460), .Z(n3459) );
  AND U3986 ( .A(n4782), .B(n4783), .Z(n3460) );
  XOR U3987 ( .A(n3463), .B(n3462), .Z(n3461) );
  AND U3988 ( .A(n4784), .B(n4785), .Z(n3462) );
  XOR U3989 ( .A(n3465), .B(n3464), .Z(n3463) );
  AND U3990 ( .A(n4786), .B(n4787), .Z(n3464) );
  XOR U3991 ( .A(n3467), .B(n3466), .Z(n3465) );
  AND U3992 ( .A(n4788), .B(n4789), .Z(n3466) );
  XOR U3993 ( .A(n3469), .B(n3468), .Z(n3467) );
  AND U3994 ( .A(n4790), .B(n4791), .Z(n3468) );
  XOR U3995 ( .A(n3471), .B(n3470), .Z(n3469) );
  AND U3996 ( .A(n4792), .B(n4793), .Z(n3470) );
  XOR U3997 ( .A(n3473), .B(n3472), .Z(n3471) );
  AND U3998 ( .A(n4794), .B(n4795), .Z(n3472) );
  XOR U3999 ( .A(n3475), .B(n3474), .Z(n3473) );
  AND U4000 ( .A(n4796), .B(n4797), .Z(n3474) );
  XOR U4001 ( .A(n3477), .B(n3476), .Z(n3475) );
  AND U4002 ( .A(n4798), .B(n4799), .Z(n3476) );
  XOR U4003 ( .A(n3479), .B(n3478), .Z(n3477) );
  AND U4004 ( .A(n4800), .B(n4801), .Z(n3478) );
  XOR U4005 ( .A(n3481), .B(n3480), .Z(n3479) );
  AND U4006 ( .A(n4802), .B(n4803), .Z(n3480) );
  XOR U4007 ( .A(n3483), .B(n3482), .Z(n3481) );
  AND U4008 ( .A(n4804), .B(n4805), .Z(n3482) );
  XOR U4009 ( .A(n3485), .B(n3484), .Z(n3483) );
  AND U4010 ( .A(n4806), .B(n4807), .Z(n3484) );
  XOR U4011 ( .A(n3487), .B(n3486), .Z(n3485) );
  AND U4012 ( .A(n4808), .B(n4809), .Z(n3486) );
  XOR U4013 ( .A(n3489), .B(n3488), .Z(n3487) );
  AND U4014 ( .A(n4810), .B(n4811), .Z(n3488) );
  XOR U4015 ( .A(n3491), .B(n3490), .Z(n3489) );
  AND U4016 ( .A(n4812), .B(n4813), .Z(n3490) );
  XOR U4017 ( .A(n3493), .B(n3492), .Z(n3491) );
  AND U4018 ( .A(n4814), .B(n4815), .Z(n3492) );
  XOR U4019 ( .A(n3495), .B(n3494), .Z(n3493) );
  AND U4020 ( .A(n4816), .B(n4817), .Z(n3494) );
  XOR U4021 ( .A(n3497), .B(n3496), .Z(n3495) );
  AND U4022 ( .A(n4818), .B(n4819), .Z(n3496) );
  XOR U4023 ( .A(n3499), .B(n3498), .Z(n3497) );
  AND U4024 ( .A(n4820), .B(n4821), .Z(n3498) );
  XOR U4025 ( .A(n3501), .B(n3500), .Z(n3499) );
  AND U4026 ( .A(n4822), .B(n4823), .Z(n3500) );
  XOR U4027 ( .A(n3503), .B(n3502), .Z(n3501) );
  AND U4028 ( .A(n4824), .B(n4825), .Z(n3502) );
  XOR U4029 ( .A(n3505), .B(n3504), .Z(n3503) );
  AND U4030 ( .A(n4826), .B(n4827), .Z(n3504) );
  XOR U4031 ( .A(n3507), .B(n3506), .Z(n3505) );
  AND U4032 ( .A(n4828), .B(n4829), .Z(n3506) );
  XOR U4033 ( .A(n3509), .B(n3508), .Z(n3507) );
  AND U4034 ( .A(n4830), .B(n4831), .Z(n3508) );
  XOR U4035 ( .A(n3511), .B(n3510), .Z(n3509) );
  AND U4036 ( .A(n4832), .B(n4833), .Z(n3510) );
  XOR U4037 ( .A(n3513), .B(n3512), .Z(n3511) );
  AND U4038 ( .A(n4834), .B(n4835), .Z(n3512) );
  XOR U4039 ( .A(n3515), .B(n3514), .Z(n3513) );
  AND U4040 ( .A(n4836), .B(n4837), .Z(n3514) );
  XOR U4041 ( .A(n3517), .B(n3516), .Z(n3515) );
  AND U4042 ( .A(n4838), .B(n4839), .Z(n3516) );
  XOR U4043 ( .A(n3519), .B(n3518), .Z(n3517) );
  AND U4044 ( .A(n4840), .B(n4841), .Z(n3518) );
  XOR U4045 ( .A(n3521), .B(n3520), .Z(n3519) );
  AND U4046 ( .A(n4842), .B(n4843), .Z(n3520) );
  XOR U4047 ( .A(n3523), .B(n3522), .Z(n3521) );
  AND U4048 ( .A(n4844), .B(n4845), .Z(n3522) );
  XOR U4049 ( .A(n3525), .B(n3524), .Z(n3523) );
  AND U4050 ( .A(n4846), .B(n4847), .Z(n3524) );
  XOR U4051 ( .A(n3658), .B(n3526), .Z(n3525) );
  AND U4052 ( .A(n4848), .B(n4849), .Z(n3526) );
  XOR U4053 ( .A(n3660), .B(n3659), .Z(n3658) );
  AND U4054 ( .A(n4850), .B(n4851), .Z(n3659) );
  XOR U4055 ( .A(n3642), .B(n3661), .Z(n3660) );
  AND U4056 ( .A(n4852), .B(n4853), .Z(n3661) );
  XOR U4057 ( .A(n3644), .B(n3643), .Z(n3642) );
  AND U4058 ( .A(n4854), .B(n4855), .Z(n3643) );
  XOR U4059 ( .A(n3646), .B(n3645), .Z(n3644) );
  AND U4060 ( .A(n4856), .B(n4857), .Z(n3645) );
  XOR U4061 ( .A(n3650), .B(n3647), .Z(n3646) );
  AND U4062 ( .A(n4858), .B(n4859), .Z(n3647) );
  XOR U4063 ( .A(n3652), .B(n3651), .Z(n3650) );
  AND U4064 ( .A(n4860), .B(n4861), .Z(n3651) );
  XOR U4065 ( .A(n3654), .B(n3653), .Z(n3652) );
  AND U4066 ( .A(n4862), .B(n4863), .Z(n3653) );
  XOR U4067 ( .A(n3656), .B(n3655), .Z(n3654) );
  AND U4068 ( .A(n4864), .B(n4865), .Z(n3655) );
  XOR U4069 ( .A(n3640), .B(n3657), .Z(n3656) );
  AND U4070 ( .A(n4866), .B(n4867), .Z(n3657) );
  XNOR U4071 ( .A(n3549), .B(n3641), .Z(n3640) );
  AND U4072 ( .A(n4868), .B(n4869), .Z(n3641) );
  XOR U4073 ( .A(n3548), .B(n3540), .Z(n3549) );
  AND U4074 ( .A(n4870), .B(n4871), .Z(n3540) );
  XNOR U4075 ( .A(n3543), .B(n3539), .Z(n3548) );
  AND U4076 ( .A(n4872), .B(n4873), .Z(n3539) );
  XOR U4077 ( .A(n3569), .B(n3544), .Z(n3543) );
  AND U4078 ( .A(n4874), .B(n4875), .Z(n3544) );
  XNOR U4079 ( .A(n3560), .B(n3570), .Z(n3569) );
  AND U4080 ( .A(n4876), .B(n4877), .Z(n3570) );
  XOR U4081 ( .A(n3558), .B(n3559), .Z(n3560) );
  AND U4082 ( .A(n4878), .B(n4879), .Z(n3559) );
  XNOR U4083 ( .A(n3552), .B(n3557), .Z(n3558) );
  AND U4084 ( .A(n4880), .B(n4881), .Z(n3557) );
  XOR U4085 ( .A(n3571), .B(n3553), .Z(n3552) );
  AND U4086 ( .A(n4882), .B(n4883), .Z(n3553) );
  XNOR U4087 ( .A(n3637), .B(n3572), .Z(n3571) );
  AND U4088 ( .A(n4884), .B(n4885), .Z(n3572) );
  XOR U4089 ( .A(n3636), .B(n3628), .Z(n3637) );
  AND U4090 ( .A(n4886), .B(n4887), .Z(n3628) );
  XNOR U4091 ( .A(n3631), .B(n3627), .Z(n3636) );
  AND U4092 ( .A(n4888), .B(n4889), .Z(n3627) );
  XOR U4093 ( .A(n3575), .B(n3632), .Z(n3631) );
  AND U4094 ( .A(n4890), .B(n4891), .Z(n3632) );
  XNOR U4095 ( .A(n3624), .B(n3576), .Z(n3575) );
  AND U4096 ( .A(n4892), .B(n4893), .Z(n3576) );
  XOR U4097 ( .A(n3623), .B(n3615), .Z(n3624) );
  AND U4098 ( .A(n4894), .B(n4895), .Z(n3615) );
  XNOR U4099 ( .A(n3618), .B(n3614), .Z(n3623) );
  AND U4100 ( .A(n4896), .B(n4897), .Z(n3614) );
  XOR U4101 ( .A(n4898), .B(n4899), .Z(n3618) );
  XOR U4102 ( .A(n3608), .B(n3609), .Z(n4899) );
  AND U4103 ( .A(n4900), .B(n4901), .Z(n3609) );
  AND U4104 ( .A(n4902), .B(n4903), .Z(n3608) );
  XOR U4105 ( .A(n4904), .B(n3619), .Z(n4898) );
  AND U4106 ( .A(n4905), .B(n4906), .Z(n3619) );
  XOR U4107 ( .A(n4907), .B(n4908), .Z(n4904) );
  XOR U4108 ( .A(n4909), .B(n4910), .Z(n4908) );
  XOR U4109 ( .A(n3601), .B(n3602), .Z(n4910) );
  AND U4110 ( .A(n4911), .B(n4912), .Z(n3602) );
  AND U4111 ( .A(n4913), .B(n4914), .Z(n3601) );
  XOR U4112 ( .A(n3595), .B(n3600), .Z(n4909) );
  AND U4113 ( .A(n4915), .B(n4916), .Z(n3600) );
  AND U4114 ( .A(n4917), .B(n4918), .Z(n3595) );
  XOR U4115 ( .A(n4919), .B(n4920), .Z(n4907) );
  XOR U4116 ( .A(n3603), .B(n3606), .Z(n4920) );
  AND U4117 ( .A(n4921), .B(n4922), .Z(n3606) );
  AND U4118 ( .A(n4923), .B(n4924), .Z(n3603) );
  XOR U4119 ( .A(n4925), .B(n3607), .Z(n4919) );
  AND U4120 ( .A(n4926), .B(n4927), .Z(n3607) );
  XOR U4121 ( .A(n4928), .B(n4929), .Z(n4925) );
  XOR U4122 ( .A(n4930), .B(n4931), .Z(n4929) );
  XOR U4123 ( .A(n3588), .B(n3589), .Z(n4931) );
  AND U4124 ( .A(n4932), .B(n4933), .Z(n3589) );
  AND U4125 ( .A(n4934), .B(n4935), .Z(n3588) );
  XOR U4126 ( .A(n3586), .B(n3584), .Z(n4930) );
  AND U4127 ( .A(n4936), .B(n4937), .Z(n3584) );
  AND U4128 ( .A(n4938), .B(n4939), .Z(n3586) );
  XOR U4129 ( .A(n4940), .B(n4941), .Z(n4928) );
  XOR U4130 ( .A(n3592), .B(n3593), .Z(n4941) );
  AND U4131 ( .A(n4942), .B(n4943), .Z(n3593) );
  AND U4132 ( .A(n4944), .B(n4945), .Z(n3592) );
  XOR U4133 ( .A(n3587), .B(n3594), .Z(n4940) );
  AND U4134 ( .A(n4946), .B(n4947), .Z(n3594) );
  XOR U4135 ( .A(n4948), .B(n4949), .Z(n3587) );
  XOR U4136 ( .A(n4950), .B(n4951), .Z(n4949) );
  XOR U4137 ( .A(n4952), .B(n4953), .Z(n4951) );
  NOR U4138 ( .A(n4954), .B(n4955), .Z(n4953) );
  NOR U4139 ( .A(n4956), .B(n4957), .Z(n4952) );
  AND U4140 ( .A(n4958), .B(n4959), .Z(n4957) );
  IV U4141 ( .A(n4960), .Z(n4956) );
  NOR U4142 ( .A(n4961), .B(n4962), .Z(n4960) );
  AND U4143 ( .A(n4954), .B(n4963), .Z(n4962) );
  AND U4144 ( .A(n4955), .B(n4964), .Z(n4961) );
  XOR U4145 ( .A(n4965), .B(n4966), .Z(n4950) );
  NOR U4146 ( .A(n4967), .B(n4968), .Z(n4966) );
  NOR U4147 ( .A(n4969), .B(n4970), .Z(n4965) );
  AND U4148 ( .A(n4971), .B(n4972), .Z(n4970) );
  IV U4149 ( .A(n4973), .Z(n4969) );
  NOR U4150 ( .A(n4974), .B(n4975), .Z(n4973) );
  AND U4151 ( .A(n4967), .B(n4976), .Z(n4975) );
  AND U4152 ( .A(n4968), .B(n4977), .Z(n4974) );
  XOR U4153 ( .A(n4978), .B(n4979), .Z(n4948) );
  AND U4154 ( .A(n4980), .B(n4981), .Z(n4979) );
  XNOR U4155 ( .A(n4982), .B(n4983), .Z(n4978) );
  AND U4156 ( .A(n4984), .B(n4985), .Z(n4983) );
  AND U4157 ( .A(n4986), .B(n4987), .Z(n4982) );
  AND U4158 ( .A(n4988), .B(n4989), .Z(n4987) );
  NOR U4159 ( .A(n4990), .B(n4991), .Z(n4989) );
  IV U4160 ( .A(n4992), .Z(n4990) );
  NOR U4161 ( .A(n4993), .B(n4994), .Z(n4992) );
  NOR U4162 ( .A(n4995), .B(n4996), .Z(n4988) );
  AND U4163 ( .A(n4997), .B(n4998), .Z(n4986) );
  NOR U4164 ( .A(n4999), .B(n5000), .Z(n4998) );
  NOR U4165 ( .A(n5001), .B(n5002), .Z(n4997) );
  XOR U4166 ( .A(n5003), .B(n5004), .Z(n3677) );
  AND U4167 ( .A(n5003), .B(n5005), .Z(n5004) );
  XNOR U4168 ( .A(n5006), .B(n5007), .Z(n3680) );
  AND U4169 ( .A(n5006), .B(n5008), .Z(n5007) );
  IV U4170 ( .A(n3683), .Z(n4759) );
  XNOR U4171 ( .A(n5009), .B(n5010), .Z(n3683) );
  AND U4172 ( .A(n5009), .B(n5011), .Z(n5010) );
  XNOR U4173 ( .A(n5012), .B(n5013), .Z(n3686) );
  AND U4174 ( .A(n5012), .B(n5014), .Z(n5013) );
  XNOR U4175 ( .A(n5015), .B(n5016), .Z(n3689) );
  AND U4176 ( .A(n5017), .B(n5015), .Z(n5016) );
  XOR U4177 ( .A(n5018), .B(n5019), .Z(n3692) );
  NOR U4178 ( .A(n5020), .B(n5018), .Z(n5019) );
  XOR U4179 ( .A(n5021), .B(n5022), .Z(n3695) );
  NOR U4180 ( .A(n5023), .B(n5021), .Z(n5022) );
  XOR U4181 ( .A(n5024), .B(n5025), .Z(n3698) );
  NOR U4182 ( .A(n5026), .B(n5024), .Z(n5025) );
  XOR U4183 ( .A(n5027), .B(n5028), .Z(n3701) );
  NOR U4184 ( .A(n5029), .B(n5027), .Z(n5028) );
  XOR U4185 ( .A(n5030), .B(n5031), .Z(n3704) );
  NOR U4186 ( .A(n5032), .B(n5030), .Z(n5031) );
  XOR U4187 ( .A(n5033), .B(n5034), .Z(n3707) );
  NOR U4188 ( .A(n5035), .B(n5033), .Z(n5034) );
  XOR U4189 ( .A(n5036), .B(n5037), .Z(n3710) );
  NOR U4190 ( .A(n5038), .B(n5036), .Z(n5037) );
  XOR U4191 ( .A(n5039), .B(n5040), .Z(n3713) );
  NOR U4192 ( .A(n5041), .B(n5039), .Z(n5040) );
  XOR U4193 ( .A(n5042), .B(n5043), .Z(n3716) );
  NOR U4194 ( .A(n5044), .B(n5042), .Z(n5043) );
  XOR U4195 ( .A(n5045), .B(n5046), .Z(n3719) );
  NOR U4196 ( .A(n5047), .B(n5045), .Z(n5046) );
  XOR U4197 ( .A(n5048), .B(n5049), .Z(n3722) );
  NOR U4198 ( .A(n5050), .B(n5048), .Z(n5049) );
  XOR U4199 ( .A(n5051), .B(n5052), .Z(n3725) );
  NOR U4200 ( .A(n5053), .B(n5051), .Z(n5052) );
  XOR U4201 ( .A(n5054), .B(n5055), .Z(n3728) );
  NOR U4202 ( .A(n5056), .B(n5054), .Z(n5055) );
  XOR U4203 ( .A(n5057), .B(n5058), .Z(n3731) );
  NOR U4204 ( .A(n5059), .B(n5057), .Z(n5058) );
  XOR U4205 ( .A(n5060), .B(n5061), .Z(n3734) );
  NOR U4206 ( .A(n5062), .B(n5060), .Z(n5061) );
  XOR U4207 ( .A(n5063), .B(n5064), .Z(n3737) );
  NOR U4208 ( .A(n5065), .B(n5063), .Z(n5064) );
  XOR U4209 ( .A(n5066), .B(n5067), .Z(n3740) );
  NOR U4210 ( .A(n5068), .B(n5066), .Z(n5067) );
  XOR U4211 ( .A(n5069), .B(n5070), .Z(n3743) );
  NOR U4212 ( .A(n5071), .B(n5069), .Z(n5070) );
  XOR U4213 ( .A(n5072), .B(n5073), .Z(n3746) );
  NOR U4214 ( .A(n5074), .B(n5072), .Z(n5073) );
  XOR U4215 ( .A(n5075), .B(n5076), .Z(n3749) );
  NOR U4216 ( .A(n5077), .B(n5075), .Z(n5076) );
  XOR U4217 ( .A(n5078), .B(n5079), .Z(n3752) );
  NOR U4218 ( .A(n5080), .B(n5078), .Z(n5079) );
  XOR U4219 ( .A(n5081), .B(n5082), .Z(n3755) );
  NOR U4220 ( .A(n5083), .B(n5081), .Z(n5082) );
  XOR U4221 ( .A(n5084), .B(n5085), .Z(n3758) );
  NOR U4222 ( .A(n5086), .B(n5084), .Z(n5085) );
  XOR U4223 ( .A(n5087), .B(n5088), .Z(n3761) );
  NOR U4224 ( .A(n5089), .B(n5087), .Z(n5088) );
  XOR U4225 ( .A(n5090), .B(n5091), .Z(n3764) );
  NOR U4226 ( .A(n5092), .B(n5090), .Z(n5091) );
  XOR U4227 ( .A(n5093), .B(n5094), .Z(n3767) );
  NOR U4228 ( .A(n5095), .B(n5093), .Z(n5094) );
  XOR U4229 ( .A(n5096), .B(n5097), .Z(n3770) );
  NOR U4230 ( .A(n5098), .B(n5096), .Z(n5097) );
  XOR U4231 ( .A(n5099), .B(n5100), .Z(n3773) );
  NOR U4232 ( .A(n5101), .B(n5099), .Z(n5100) );
  XOR U4233 ( .A(n5102), .B(n5103), .Z(n3776) );
  NOR U4234 ( .A(n5104), .B(n5102), .Z(n5103) );
  XOR U4235 ( .A(n5105), .B(n5106), .Z(n3779) );
  NOR U4236 ( .A(n5107), .B(n5105), .Z(n5106) );
  XOR U4237 ( .A(n5108), .B(n5109), .Z(n3782) );
  NOR U4238 ( .A(n5110), .B(n5108), .Z(n5109) );
  XOR U4239 ( .A(n5111), .B(n5112), .Z(n3785) );
  NOR U4240 ( .A(n5113), .B(n5111), .Z(n5112) );
  XOR U4241 ( .A(n5114), .B(n5115), .Z(n3788) );
  NOR U4242 ( .A(n5116), .B(n5114), .Z(n5115) );
  XOR U4243 ( .A(n5117), .B(n5118), .Z(n3791) );
  NOR U4244 ( .A(n5119), .B(n5117), .Z(n5118) );
  XOR U4245 ( .A(n5120), .B(n5121), .Z(n3794) );
  NOR U4246 ( .A(n5122), .B(n5120), .Z(n5121) );
  XOR U4247 ( .A(n5123), .B(n5124), .Z(n3797) );
  NOR U4248 ( .A(n5125), .B(n5123), .Z(n5124) );
  XOR U4249 ( .A(n5126), .B(n5127), .Z(n3800) );
  NOR U4250 ( .A(n5128), .B(n5126), .Z(n5127) );
  XOR U4251 ( .A(n5129), .B(n5130), .Z(n3803) );
  NOR U4252 ( .A(n5131), .B(n5129), .Z(n5130) );
  XOR U4253 ( .A(n5132), .B(n5133), .Z(n3806) );
  NOR U4254 ( .A(n5134), .B(n5132), .Z(n5133) );
  XOR U4255 ( .A(n5135), .B(n5136), .Z(n3809) );
  NOR U4256 ( .A(n5137), .B(n5135), .Z(n5136) );
  XOR U4257 ( .A(n5138), .B(n5139), .Z(n3812) );
  NOR U4258 ( .A(n5140), .B(n5138), .Z(n5139) );
  XOR U4259 ( .A(n5141), .B(n5142), .Z(n3815) );
  NOR U4260 ( .A(n5143), .B(n5141), .Z(n5142) );
  XOR U4261 ( .A(n5144), .B(n5145), .Z(n3818) );
  NOR U4262 ( .A(n5146), .B(n5144), .Z(n5145) );
  XOR U4263 ( .A(n5147), .B(n5148), .Z(n3821) );
  NOR U4264 ( .A(n5149), .B(n5147), .Z(n5148) );
  XOR U4265 ( .A(n5150), .B(n5151), .Z(n3824) );
  NOR U4266 ( .A(n5152), .B(n5150), .Z(n5151) );
  XOR U4267 ( .A(n5153), .B(n5154), .Z(n3827) );
  NOR U4268 ( .A(n5155), .B(n5153), .Z(n5154) );
  XOR U4269 ( .A(n5156), .B(n5157), .Z(n3830) );
  NOR U4270 ( .A(n5158), .B(n5156), .Z(n5157) );
  XOR U4271 ( .A(n5159), .B(n5160), .Z(n3833) );
  NOR U4272 ( .A(n5161), .B(n5159), .Z(n5160) );
  XOR U4273 ( .A(n5162), .B(n5163), .Z(n3836) );
  NOR U4274 ( .A(n5164), .B(n5162), .Z(n5163) );
  XOR U4275 ( .A(n5165), .B(n5166), .Z(n3839) );
  NOR U4276 ( .A(n5167), .B(n5165), .Z(n5166) );
  XOR U4277 ( .A(n5168), .B(n5169), .Z(n3842) );
  NOR U4278 ( .A(n5170), .B(n5168), .Z(n5169) );
  XOR U4279 ( .A(n5171), .B(n5172), .Z(n3845) );
  NOR U4280 ( .A(n5173), .B(n5171), .Z(n5172) );
  XOR U4281 ( .A(n5174), .B(n5175), .Z(n3848) );
  NOR U4282 ( .A(n5176), .B(n5174), .Z(n5175) );
  XOR U4283 ( .A(n5177), .B(n5178), .Z(n3851) );
  NOR U4284 ( .A(n5179), .B(n5177), .Z(n5178) );
  XOR U4285 ( .A(n5180), .B(n5181), .Z(n3854) );
  NOR U4286 ( .A(n5182), .B(n5180), .Z(n5181) );
  XOR U4287 ( .A(n5183), .B(n5184), .Z(n3857) );
  NOR U4288 ( .A(n5185), .B(n5183), .Z(n5184) );
  XOR U4289 ( .A(n5186), .B(n5187), .Z(n3860) );
  NOR U4290 ( .A(n5188), .B(n5186), .Z(n5187) );
  XOR U4291 ( .A(n5189), .B(n5190), .Z(n3863) );
  NOR U4292 ( .A(n5191), .B(n5189), .Z(n5190) );
  XOR U4293 ( .A(n5192), .B(n5193), .Z(n3866) );
  NOR U4294 ( .A(n5194), .B(n5192), .Z(n5193) );
  XOR U4295 ( .A(n5195), .B(n5196), .Z(n3869) );
  NOR U4296 ( .A(n5197), .B(n5195), .Z(n5196) );
  XOR U4297 ( .A(n5198), .B(n5199), .Z(n3872) );
  NOR U4298 ( .A(n5200), .B(n5198), .Z(n5199) );
  XOR U4299 ( .A(n5201), .B(n5202), .Z(n3875) );
  NOR U4300 ( .A(n5203), .B(n5201), .Z(n5202) );
  XOR U4301 ( .A(n5204), .B(n5205), .Z(n3878) );
  NOR U4302 ( .A(n5206), .B(n5204), .Z(n5205) );
  XOR U4303 ( .A(n5207), .B(n5208), .Z(n3881) );
  NOR U4304 ( .A(n5209), .B(n5207), .Z(n5208) );
  XOR U4305 ( .A(n5210), .B(n5211), .Z(n3884) );
  NOR U4306 ( .A(n5212), .B(n5210), .Z(n5211) );
  XOR U4307 ( .A(n5213), .B(n5214), .Z(n3887) );
  NOR U4308 ( .A(n5215), .B(n5213), .Z(n5214) );
  XOR U4309 ( .A(n5216), .B(n5217), .Z(n3890) );
  NOR U4310 ( .A(n5218), .B(n5216), .Z(n5217) );
  XOR U4311 ( .A(n5219), .B(n5220), .Z(n3893) );
  NOR U4312 ( .A(n5221), .B(n5219), .Z(n5220) );
  XOR U4313 ( .A(n5222), .B(n5223), .Z(n3896) );
  NOR U4314 ( .A(n5224), .B(n5222), .Z(n5223) );
  XOR U4315 ( .A(n5225), .B(n5226), .Z(n3899) );
  NOR U4316 ( .A(n5227), .B(n5225), .Z(n5226) );
  XOR U4317 ( .A(n5228), .B(n5229), .Z(n3902) );
  NOR U4318 ( .A(n5230), .B(n5228), .Z(n5229) );
  XOR U4319 ( .A(n5231), .B(n5232), .Z(n3905) );
  NOR U4320 ( .A(n5233), .B(n5231), .Z(n5232) );
  XOR U4321 ( .A(n5234), .B(n5235), .Z(n3908) );
  NOR U4322 ( .A(n5236), .B(n5234), .Z(n5235) );
  XOR U4323 ( .A(n5237), .B(n5238), .Z(n3911) );
  NOR U4324 ( .A(n5239), .B(n5237), .Z(n5238) );
  XOR U4325 ( .A(n5240), .B(n5241), .Z(n3914) );
  NOR U4326 ( .A(n5242), .B(n5240), .Z(n5241) );
  XOR U4327 ( .A(n5243), .B(n5244), .Z(n3917) );
  NOR U4328 ( .A(n5245), .B(n5243), .Z(n5244) );
  XOR U4329 ( .A(n5246), .B(n5247), .Z(n3920) );
  NOR U4330 ( .A(n5248), .B(n5246), .Z(n5247) );
  XOR U4331 ( .A(n5249), .B(n5250), .Z(n3923) );
  NOR U4332 ( .A(n5251), .B(n5249), .Z(n5250) );
  XOR U4333 ( .A(n5252), .B(n5253), .Z(n3926) );
  NOR U4334 ( .A(n5254), .B(n5252), .Z(n5253) );
  XOR U4335 ( .A(n5255), .B(n5256), .Z(n3929) );
  NOR U4336 ( .A(n5257), .B(n5255), .Z(n5256) );
  XOR U4337 ( .A(n5258), .B(n5259), .Z(n3932) );
  NOR U4338 ( .A(n5260), .B(n5258), .Z(n5259) );
  XOR U4339 ( .A(n5261), .B(n5262), .Z(n3935) );
  NOR U4340 ( .A(n5263), .B(n5261), .Z(n5262) );
  XOR U4341 ( .A(n5264), .B(n5265), .Z(n3938) );
  NOR U4342 ( .A(n5266), .B(n5264), .Z(n5265) );
  XOR U4343 ( .A(n5267), .B(n5268), .Z(n3941) );
  NOR U4344 ( .A(n5269), .B(n5267), .Z(n5268) );
  XOR U4345 ( .A(n5270), .B(n5271), .Z(n3944) );
  NOR U4346 ( .A(n5272), .B(n5270), .Z(n5271) );
  XOR U4347 ( .A(n5273), .B(n5274), .Z(n3947) );
  NOR U4348 ( .A(n5275), .B(n5273), .Z(n5274) );
  XOR U4349 ( .A(n5276), .B(n5277), .Z(n3950) );
  NOR U4350 ( .A(n5278), .B(n5276), .Z(n5277) );
  XOR U4351 ( .A(n5279), .B(n5280), .Z(n3953) );
  NOR U4352 ( .A(n5281), .B(n5279), .Z(n5280) );
  XOR U4353 ( .A(n5282), .B(n5283), .Z(n3956) );
  NOR U4354 ( .A(n5284), .B(n5282), .Z(n5283) );
  XOR U4355 ( .A(n5285), .B(n5286), .Z(n3959) );
  NOR U4356 ( .A(n5287), .B(n5285), .Z(n5286) );
  XOR U4357 ( .A(n5288), .B(n5289), .Z(n3962) );
  NOR U4358 ( .A(n5290), .B(n5288), .Z(n5289) );
  XOR U4359 ( .A(n5291), .B(n5292), .Z(n3965) );
  NOR U4360 ( .A(n5293), .B(n5291), .Z(n5292) );
  XOR U4361 ( .A(n5294), .B(n5295), .Z(n3968) );
  NOR U4362 ( .A(n5296), .B(n5294), .Z(n5295) );
  XOR U4363 ( .A(n5297), .B(n5298), .Z(n3971) );
  NOR U4364 ( .A(n5299), .B(n5297), .Z(n5298) );
  XOR U4365 ( .A(n5300), .B(n5301), .Z(n3974) );
  NOR U4366 ( .A(n5302), .B(n5300), .Z(n5301) );
  XOR U4367 ( .A(n5303), .B(n5304), .Z(n3977) );
  NOR U4368 ( .A(n5305), .B(n5303), .Z(n5304) );
  XOR U4369 ( .A(n5306), .B(n5307), .Z(n3980) );
  NOR U4370 ( .A(n5308), .B(n5306), .Z(n5307) );
  XOR U4371 ( .A(n5309), .B(n5310), .Z(n3983) );
  NOR U4372 ( .A(n5311), .B(n5309), .Z(n5310) );
  XOR U4373 ( .A(n5312), .B(n5313), .Z(n3986) );
  NOR U4374 ( .A(n5314), .B(n5312), .Z(n5313) );
  XOR U4375 ( .A(n5315), .B(n5316), .Z(n3989) );
  NOR U4376 ( .A(n5317), .B(n5315), .Z(n5316) );
  XOR U4377 ( .A(n5318), .B(n5319), .Z(n3992) );
  NOR U4378 ( .A(n5320), .B(n5318), .Z(n5319) );
  XOR U4379 ( .A(n5321), .B(n5322), .Z(n3995) );
  NOR U4380 ( .A(n5323), .B(n5321), .Z(n5322) );
  XOR U4381 ( .A(n5324), .B(n5325), .Z(n3998) );
  NOR U4382 ( .A(n5326), .B(n5324), .Z(n5325) );
  XOR U4383 ( .A(n5327), .B(n5328), .Z(n4001) );
  NOR U4384 ( .A(n5329), .B(n5327), .Z(n5328) );
  XOR U4385 ( .A(n5330), .B(n5331), .Z(n4004) );
  NOR U4386 ( .A(n5332), .B(n5330), .Z(n5331) );
  XOR U4387 ( .A(n5333), .B(n5334), .Z(n4007) );
  NOR U4388 ( .A(n5335), .B(n5333), .Z(n5334) );
  XOR U4389 ( .A(n5336), .B(n5337), .Z(n4010) );
  NOR U4390 ( .A(n5338), .B(n5336), .Z(n5337) );
  XOR U4391 ( .A(n5339), .B(n5340), .Z(n4013) );
  NOR U4392 ( .A(n5341), .B(n5339), .Z(n5340) );
  XOR U4393 ( .A(n5342), .B(n5343), .Z(n4016) );
  NOR U4394 ( .A(n5344), .B(n5342), .Z(n5343) );
  XOR U4395 ( .A(n5345), .B(n5346), .Z(n4019) );
  NOR U4396 ( .A(n5347), .B(n5345), .Z(n5346) );
  XOR U4397 ( .A(n5348), .B(n5349), .Z(n4022) );
  NOR U4398 ( .A(n5350), .B(n5348), .Z(n5349) );
  XOR U4399 ( .A(n5351), .B(n5352), .Z(n4025) );
  NOR U4400 ( .A(n5353), .B(n5351), .Z(n5352) );
  XOR U4401 ( .A(n5354), .B(n5355), .Z(n4028) );
  NOR U4402 ( .A(n5356), .B(n5354), .Z(n5355) );
  XOR U4403 ( .A(n5357), .B(n5358), .Z(n4031) );
  NOR U4404 ( .A(n5359), .B(n5357), .Z(n5358) );
  XOR U4405 ( .A(n5360), .B(n5361), .Z(n4034) );
  NOR U4406 ( .A(n5362), .B(n5360), .Z(n5361) );
  XOR U4407 ( .A(n5363), .B(n5364), .Z(n4037) );
  NOR U4408 ( .A(n5365), .B(n5363), .Z(n5364) );
  XOR U4409 ( .A(n5366), .B(n5367), .Z(n4040) );
  NOR U4410 ( .A(n5368), .B(n5366), .Z(n5367) );
  XOR U4411 ( .A(n5369), .B(n5370), .Z(n4043) );
  NOR U4412 ( .A(n5371), .B(n5369), .Z(n5370) );
  XOR U4413 ( .A(n5372), .B(n5373), .Z(n4046) );
  NOR U4414 ( .A(n5374), .B(n5372), .Z(n5373) );
  XOR U4415 ( .A(n5375), .B(n5376), .Z(n4049) );
  NOR U4416 ( .A(n5377), .B(n5375), .Z(n5376) );
  XOR U4417 ( .A(n5378), .B(n5379), .Z(n4052) );
  NOR U4418 ( .A(n5380), .B(n5378), .Z(n5379) );
  XOR U4419 ( .A(n5381), .B(n5382), .Z(n4055) );
  NOR U4420 ( .A(n5383), .B(n5381), .Z(n5382) );
  XOR U4421 ( .A(n5384), .B(n5385), .Z(n4058) );
  NOR U4422 ( .A(n5386), .B(n5384), .Z(n5385) );
  XOR U4423 ( .A(n5387), .B(n5388), .Z(n4061) );
  NOR U4424 ( .A(n5389), .B(n5387), .Z(n5388) );
  XOR U4425 ( .A(n5390), .B(n5391), .Z(n4064) );
  NOR U4426 ( .A(n5392), .B(n5390), .Z(n5391) );
  XOR U4427 ( .A(n5393), .B(n5394), .Z(n4067) );
  NOR U4428 ( .A(n5395), .B(n5393), .Z(n5394) );
  XOR U4429 ( .A(n5396), .B(n5397), .Z(n4070) );
  NOR U4430 ( .A(n5398), .B(n5396), .Z(n5397) );
  XOR U4431 ( .A(n5399), .B(n5400), .Z(n4073) );
  NOR U4432 ( .A(n5401), .B(n5399), .Z(n5400) );
  XOR U4433 ( .A(n5402), .B(n5403), .Z(n4076) );
  NOR U4434 ( .A(n5404), .B(n5402), .Z(n5403) );
  XOR U4435 ( .A(n5405), .B(n5406), .Z(n4079) );
  NOR U4436 ( .A(n5407), .B(n5405), .Z(n5406) );
  XOR U4437 ( .A(n5408), .B(n5409), .Z(n4082) );
  NOR U4438 ( .A(n5410), .B(n5408), .Z(n5409) );
  XOR U4439 ( .A(n5411), .B(n5412), .Z(n4085) );
  NOR U4440 ( .A(n5413), .B(n5411), .Z(n5412) );
  XOR U4441 ( .A(n5414), .B(n5415), .Z(n4088) );
  NOR U4442 ( .A(n5416), .B(n5414), .Z(n5415) );
  XOR U4443 ( .A(n5417), .B(n5418), .Z(n4091) );
  NOR U4444 ( .A(n86), .B(n5419), .Z(n5418) );
  IV U4445 ( .A(n5417), .Z(n5419) );
  XOR U4446 ( .A(n5420), .B(n5421), .Z(n4094) );
  AND U4447 ( .A(n5422), .B(n5423), .Z(n5421) );
  XOR U4448 ( .A(n5420), .B(n88), .Z(n5423) );
  XOR U4449 ( .A(n4756), .B(n4755), .Z(n88) );
  XNOR U4450 ( .A(n4753), .B(n4752), .Z(n4755) );
  XNOR U4451 ( .A(n4750), .B(n4749), .Z(n4752) );
  XNOR U4452 ( .A(n4747), .B(n4746), .Z(n4749) );
  XNOR U4453 ( .A(n4744), .B(n4743), .Z(n4746) );
  XNOR U4454 ( .A(n4741), .B(n4740), .Z(n4743) );
  XNOR U4455 ( .A(n4738), .B(n4737), .Z(n4740) );
  XNOR U4456 ( .A(n4735), .B(n4734), .Z(n4737) );
  XNOR U4457 ( .A(n4732), .B(n4731), .Z(n4734) );
  XNOR U4458 ( .A(n4729), .B(n4728), .Z(n4731) );
  XNOR U4459 ( .A(n4726), .B(n4725), .Z(n4728) );
  XNOR U4460 ( .A(n4723), .B(n4722), .Z(n4725) );
  XNOR U4461 ( .A(n4720), .B(n4719), .Z(n4722) );
  XNOR U4462 ( .A(n4717), .B(n4716), .Z(n4719) );
  XNOR U4463 ( .A(n4714), .B(n4713), .Z(n4716) );
  XNOR U4464 ( .A(n4711), .B(n4710), .Z(n4713) );
  XNOR U4465 ( .A(n4708), .B(n4707), .Z(n4710) );
  XNOR U4466 ( .A(n4705), .B(n4704), .Z(n4707) );
  XNOR U4467 ( .A(n4702), .B(n4701), .Z(n4704) );
  XNOR U4468 ( .A(n4699), .B(n4698), .Z(n4701) );
  XNOR U4469 ( .A(n4696), .B(n4695), .Z(n4698) );
  XNOR U4470 ( .A(n4693), .B(n4692), .Z(n4695) );
  XNOR U4471 ( .A(n4690), .B(n4689), .Z(n4692) );
  XNOR U4472 ( .A(n4687), .B(n4686), .Z(n4689) );
  XNOR U4473 ( .A(n4684), .B(n4683), .Z(n4686) );
  XNOR U4474 ( .A(n4681), .B(n4680), .Z(n4683) );
  XNOR U4475 ( .A(n4678), .B(n4677), .Z(n4680) );
  XNOR U4476 ( .A(n4675), .B(n4674), .Z(n4677) );
  XNOR U4477 ( .A(n4672), .B(n4671), .Z(n4674) );
  XNOR U4478 ( .A(n4669), .B(n4668), .Z(n4671) );
  XNOR U4479 ( .A(n4666), .B(n4665), .Z(n4668) );
  XNOR U4480 ( .A(n4663), .B(n4662), .Z(n4665) );
  XNOR U4481 ( .A(n4660), .B(n4659), .Z(n4662) );
  XNOR U4482 ( .A(n4657), .B(n4656), .Z(n4659) );
  XNOR U4483 ( .A(n4654), .B(n4653), .Z(n4656) );
  XNOR U4484 ( .A(n4651), .B(n4650), .Z(n4653) );
  XNOR U4485 ( .A(n4648), .B(n4647), .Z(n4650) );
  XNOR U4486 ( .A(n4645), .B(n4644), .Z(n4647) );
  XNOR U4487 ( .A(n4642), .B(n4641), .Z(n4644) );
  XNOR U4488 ( .A(n4639), .B(n4638), .Z(n4641) );
  XNOR U4489 ( .A(n4636), .B(n4635), .Z(n4638) );
  XNOR U4490 ( .A(n4633), .B(n4632), .Z(n4635) );
  XNOR U4491 ( .A(n4630), .B(n4629), .Z(n4632) );
  XNOR U4492 ( .A(n4627), .B(n4626), .Z(n4629) );
  XNOR U4493 ( .A(n4624), .B(n4623), .Z(n4626) );
  XNOR U4494 ( .A(n4621), .B(n4620), .Z(n4623) );
  XNOR U4495 ( .A(n4618), .B(n4617), .Z(n4620) );
  XNOR U4496 ( .A(n4615), .B(n4614), .Z(n4617) );
  XNOR U4497 ( .A(n4612), .B(n4611), .Z(n4614) );
  XNOR U4498 ( .A(n4609), .B(n4608), .Z(n4611) );
  XNOR U4499 ( .A(n4606), .B(n4605), .Z(n4608) );
  XNOR U4500 ( .A(n4603), .B(n4602), .Z(n4605) );
  XNOR U4501 ( .A(n4600), .B(n4599), .Z(n4602) );
  XNOR U4502 ( .A(n4597), .B(n4596), .Z(n4599) );
  XNOR U4503 ( .A(n4594), .B(n4593), .Z(n4596) );
  XNOR U4504 ( .A(n4591), .B(n4590), .Z(n4593) );
  XNOR U4505 ( .A(n4588), .B(n4587), .Z(n4590) );
  XNOR U4506 ( .A(n4585), .B(n4584), .Z(n4587) );
  XNOR U4507 ( .A(n4582), .B(n4581), .Z(n4584) );
  XNOR U4508 ( .A(n4579), .B(n4578), .Z(n4581) );
  XNOR U4509 ( .A(n4576), .B(n4575), .Z(n4578) );
  XNOR U4510 ( .A(n4573), .B(n4572), .Z(n4575) );
  XNOR U4511 ( .A(n4570), .B(n4569), .Z(n4572) );
  XNOR U4512 ( .A(n4567), .B(n4566), .Z(n4569) );
  XNOR U4513 ( .A(n4564), .B(n4563), .Z(n4566) );
  XNOR U4514 ( .A(n4561), .B(n4560), .Z(n4563) );
  XNOR U4515 ( .A(n4558), .B(n4557), .Z(n4560) );
  XNOR U4516 ( .A(n4555), .B(n4554), .Z(n4557) );
  XNOR U4517 ( .A(n4552), .B(n4551), .Z(n4554) );
  XNOR U4518 ( .A(n4549), .B(n4548), .Z(n4551) );
  XNOR U4519 ( .A(n4546), .B(n4545), .Z(n4548) );
  XNOR U4520 ( .A(n4543), .B(n4542), .Z(n4545) );
  XNOR U4521 ( .A(n4540), .B(n4539), .Z(n4542) );
  XNOR U4522 ( .A(n4537), .B(n4536), .Z(n4539) );
  XNOR U4523 ( .A(n4534), .B(n4533), .Z(n4536) );
  XNOR U4524 ( .A(n4531), .B(n4530), .Z(n4533) );
  XNOR U4525 ( .A(n4528), .B(n4527), .Z(n4530) );
  XNOR U4526 ( .A(n4525), .B(n4524), .Z(n4527) );
  XNOR U4527 ( .A(n4522), .B(n4521), .Z(n4524) );
  XNOR U4528 ( .A(n4519), .B(n4518), .Z(n4521) );
  XNOR U4529 ( .A(n4516), .B(n4515), .Z(n4518) );
  XNOR U4530 ( .A(n4513), .B(n4512), .Z(n4515) );
  XNOR U4531 ( .A(n4510), .B(n4509), .Z(n4512) );
  XNOR U4532 ( .A(n4507), .B(n4506), .Z(n4509) );
  XNOR U4533 ( .A(n4504), .B(n4503), .Z(n4506) );
  XNOR U4534 ( .A(n4501), .B(n4500), .Z(n4503) );
  XNOR U4535 ( .A(n4498), .B(n4497), .Z(n4500) );
  XNOR U4536 ( .A(n4495), .B(n4494), .Z(n4497) );
  XNOR U4537 ( .A(n4492), .B(n4491), .Z(n4494) );
  XNOR U4538 ( .A(n4489), .B(n4488), .Z(n4491) );
  XNOR U4539 ( .A(n4486), .B(n4485), .Z(n4488) );
  XNOR U4540 ( .A(n4483), .B(n4482), .Z(n4485) );
  XNOR U4541 ( .A(n4480), .B(n4479), .Z(n4482) );
  XNOR U4542 ( .A(n4477), .B(n4476), .Z(n4479) );
  XNOR U4543 ( .A(n4474), .B(n4473), .Z(n4476) );
  XNOR U4544 ( .A(n4471), .B(n4470), .Z(n4473) );
  XNOR U4545 ( .A(n4468), .B(n4467), .Z(n4470) );
  XNOR U4546 ( .A(n4465), .B(n4464), .Z(n4467) );
  XNOR U4547 ( .A(n4462), .B(n4461), .Z(n4464) );
  XNOR U4548 ( .A(n4459), .B(n4458), .Z(n4461) );
  XNOR U4549 ( .A(n4456), .B(n4455), .Z(n4458) );
  XNOR U4550 ( .A(n4453), .B(n4452), .Z(n4455) );
  XNOR U4551 ( .A(n4450), .B(n4449), .Z(n4452) );
  XNOR U4552 ( .A(n4447), .B(n4446), .Z(n4449) );
  XNOR U4553 ( .A(n4444), .B(n4443), .Z(n4446) );
  XNOR U4554 ( .A(n4441), .B(n4440), .Z(n4443) );
  XNOR U4555 ( .A(n4438), .B(n4437), .Z(n4440) );
  XNOR U4556 ( .A(n4435), .B(n4434), .Z(n4437) );
  XNOR U4557 ( .A(n4432), .B(n4431), .Z(n4434) );
  XNOR U4558 ( .A(n4429), .B(n4428), .Z(n4431) );
  XNOR U4559 ( .A(n4426), .B(n4425), .Z(n4428) );
  XNOR U4560 ( .A(n4423), .B(n4422), .Z(n4425) );
  XNOR U4561 ( .A(n4420), .B(n4419), .Z(n4422) );
  XNOR U4562 ( .A(n4417), .B(n4416), .Z(n4419) );
  XNOR U4563 ( .A(n4414), .B(n4413), .Z(n4416) );
  XNOR U4564 ( .A(n4411), .B(n4410), .Z(n4413) );
  XNOR U4565 ( .A(n4408), .B(n4407), .Z(n4410) );
  XNOR U4566 ( .A(n4405), .B(n4404), .Z(n4407) );
  XNOR U4567 ( .A(n4402), .B(n4401), .Z(n4404) );
  XNOR U4568 ( .A(n4399), .B(n4398), .Z(n4401) );
  XNOR U4569 ( .A(n4396), .B(n4395), .Z(n4398) );
  XNOR U4570 ( .A(n4393), .B(n4392), .Z(n4395) );
  XNOR U4571 ( .A(n4390), .B(n4389), .Z(n4392) );
  XNOR U4572 ( .A(n4387), .B(n4386), .Z(n4389) );
  XNOR U4573 ( .A(n4384), .B(n4383), .Z(n4386) );
  XNOR U4574 ( .A(n4381), .B(n4380), .Z(n4383) );
  XNOR U4575 ( .A(n4378), .B(n4377), .Z(n4380) );
  XNOR U4576 ( .A(n4375), .B(n4374), .Z(n4377) );
  XNOR U4577 ( .A(n4372), .B(n4371), .Z(n4374) );
  XNOR U4578 ( .A(n4369), .B(n4368), .Z(n4371) );
  XNOR U4579 ( .A(n4366), .B(n4365), .Z(n4368) );
  XNOR U4580 ( .A(n4363), .B(n4362), .Z(n4365) );
  XNOR U4581 ( .A(n4360), .B(n4359), .Z(n4362) );
  XOR U4582 ( .A(n4357), .B(n4356), .Z(n4359) );
  XOR U4583 ( .A(n4354), .B(n4353), .Z(n4356) );
  XOR U4584 ( .A(n4350), .B(n4351), .Z(n4353) );
  AND U4585 ( .A(n5424), .B(n5425), .Z(n4351) );
  XOR U4586 ( .A(n4347), .B(n4348), .Z(n4350) );
  AND U4587 ( .A(n5426), .B(n5427), .Z(n4348) );
  XOR U4588 ( .A(n4344), .B(n4345), .Z(n4347) );
  AND U4589 ( .A(n5428), .B(n5429), .Z(n4345) );
  XNOR U4590 ( .A(n4099), .B(n4342), .Z(n4344) );
  AND U4591 ( .A(n5430), .B(n5431), .Z(n4342) );
  XOR U4592 ( .A(n4101), .B(n4100), .Z(n4099) );
  AND U4593 ( .A(n5432), .B(n5433), .Z(n4100) );
  XOR U4594 ( .A(n4103), .B(n4102), .Z(n4101) );
  AND U4595 ( .A(n5434), .B(n5435), .Z(n4102) );
  XOR U4596 ( .A(n4105), .B(n4104), .Z(n4103) );
  AND U4597 ( .A(n5436), .B(n5437), .Z(n4104) );
  XOR U4598 ( .A(n4107), .B(n4106), .Z(n4105) );
  AND U4599 ( .A(n5438), .B(n5439), .Z(n4106) );
  XOR U4600 ( .A(n4109), .B(n4108), .Z(n4107) );
  AND U4601 ( .A(n5440), .B(n5441), .Z(n4108) );
  XOR U4602 ( .A(n4111), .B(n4110), .Z(n4109) );
  AND U4603 ( .A(n5442), .B(n5443), .Z(n4110) );
  XOR U4604 ( .A(n4113), .B(n4112), .Z(n4111) );
  AND U4605 ( .A(n5444), .B(n5445), .Z(n4112) );
  XOR U4606 ( .A(n4115), .B(n4114), .Z(n4113) );
  AND U4607 ( .A(n5446), .B(n5447), .Z(n4114) );
  XOR U4608 ( .A(n4117), .B(n4116), .Z(n4115) );
  AND U4609 ( .A(n5448), .B(n5449), .Z(n4116) );
  XOR U4610 ( .A(n4119), .B(n4118), .Z(n4117) );
  AND U4611 ( .A(n5450), .B(n5451), .Z(n4118) );
  XOR U4612 ( .A(n4121), .B(n4120), .Z(n4119) );
  AND U4613 ( .A(n5452), .B(n5453), .Z(n4120) );
  XOR U4614 ( .A(n4123), .B(n4122), .Z(n4121) );
  AND U4615 ( .A(n5454), .B(n5455), .Z(n4122) );
  XOR U4616 ( .A(n4125), .B(n4124), .Z(n4123) );
  AND U4617 ( .A(n5456), .B(n5457), .Z(n4124) );
  XOR U4618 ( .A(n4127), .B(n4126), .Z(n4125) );
  AND U4619 ( .A(n5458), .B(n5459), .Z(n4126) );
  XOR U4620 ( .A(n4129), .B(n4128), .Z(n4127) );
  AND U4621 ( .A(n5460), .B(n5461), .Z(n4128) );
  XOR U4622 ( .A(n4131), .B(n4130), .Z(n4129) );
  AND U4623 ( .A(n5462), .B(n5463), .Z(n4130) );
  XOR U4624 ( .A(n4133), .B(n4132), .Z(n4131) );
  AND U4625 ( .A(n5464), .B(n5465), .Z(n4132) );
  XOR U4626 ( .A(n4135), .B(n4134), .Z(n4133) );
  AND U4627 ( .A(n5466), .B(n5467), .Z(n4134) );
  XOR U4628 ( .A(n4137), .B(n4136), .Z(n4135) );
  AND U4629 ( .A(n5468), .B(n5469), .Z(n4136) );
  XOR U4630 ( .A(n4139), .B(n4138), .Z(n4137) );
  AND U4631 ( .A(n5470), .B(n5471), .Z(n4138) );
  XOR U4632 ( .A(n4141), .B(n4140), .Z(n4139) );
  AND U4633 ( .A(n5472), .B(n5473), .Z(n4140) );
  XOR U4634 ( .A(n4143), .B(n4142), .Z(n4141) );
  AND U4635 ( .A(n5474), .B(n5475), .Z(n4142) );
  XOR U4636 ( .A(n4145), .B(n4144), .Z(n4143) );
  AND U4637 ( .A(n5476), .B(n5477), .Z(n4144) );
  XOR U4638 ( .A(n4147), .B(n4146), .Z(n4145) );
  AND U4639 ( .A(n5478), .B(n5479), .Z(n4146) );
  XOR U4640 ( .A(n4149), .B(n4148), .Z(n4147) );
  AND U4641 ( .A(n5480), .B(n5481), .Z(n4148) );
  XOR U4642 ( .A(n4151), .B(n4150), .Z(n4149) );
  AND U4643 ( .A(n5482), .B(n5483), .Z(n4150) );
  XOR U4644 ( .A(n4153), .B(n4152), .Z(n4151) );
  AND U4645 ( .A(n5484), .B(n5485), .Z(n4152) );
  XOR U4646 ( .A(n4155), .B(n4154), .Z(n4153) );
  AND U4647 ( .A(n5486), .B(n5487), .Z(n4154) );
  XOR U4648 ( .A(n4157), .B(n4156), .Z(n4155) );
  AND U4649 ( .A(n5488), .B(n5489), .Z(n4156) );
  XOR U4650 ( .A(n4159), .B(n4158), .Z(n4157) );
  AND U4651 ( .A(n5490), .B(n5491), .Z(n4158) );
  XOR U4652 ( .A(n4161), .B(n4160), .Z(n4159) );
  AND U4653 ( .A(n5492), .B(n5493), .Z(n4160) );
  XOR U4654 ( .A(n4163), .B(n4162), .Z(n4161) );
  AND U4655 ( .A(n5494), .B(n5495), .Z(n4162) );
  XOR U4656 ( .A(n4165), .B(n4164), .Z(n4163) );
  AND U4657 ( .A(n5496), .B(n5497), .Z(n4164) );
  XOR U4658 ( .A(n4167), .B(n4166), .Z(n4165) );
  AND U4659 ( .A(n5498), .B(n5499), .Z(n4166) );
  XOR U4660 ( .A(n4169), .B(n4168), .Z(n4167) );
  AND U4661 ( .A(n5500), .B(n5501), .Z(n4168) );
  XOR U4662 ( .A(n4171), .B(n4170), .Z(n4169) );
  AND U4663 ( .A(n5502), .B(n5503), .Z(n4170) );
  XOR U4664 ( .A(n4173), .B(n4172), .Z(n4171) );
  AND U4665 ( .A(n5504), .B(n5505), .Z(n4172) );
  XOR U4666 ( .A(n4175), .B(n4174), .Z(n4173) );
  AND U4667 ( .A(n5506), .B(n5507), .Z(n4174) );
  XOR U4668 ( .A(n4177), .B(n4176), .Z(n4175) );
  AND U4669 ( .A(n5508), .B(n5509), .Z(n4176) );
  XOR U4670 ( .A(n4179), .B(n4178), .Z(n4177) );
  AND U4671 ( .A(n5510), .B(n5511), .Z(n4178) );
  XOR U4672 ( .A(n4181), .B(n4180), .Z(n4179) );
  AND U4673 ( .A(n5512), .B(n5513), .Z(n4180) );
  XOR U4674 ( .A(n4183), .B(n4182), .Z(n4181) );
  AND U4675 ( .A(n5514), .B(n5515), .Z(n4182) );
  XOR U4676 ( .A(n4185), .B(n4184), .Z(n4183) );
  AND U4677 ( .A(n5516), .B(n5517), .Z(n4184) );
  XOR U4678 ( .A(n4187), .B(n4186), .Z(n4185) );
  AND U4679 ( .A(n5518), .B(n5519), .Z(n4186) );
  XOR U4680 ( .A(n4189), .B(n4188), .Z(n4187) );
  AND U4681 ( .A(n5520), .B(n5521), .Z(n4188) );
  XOR U4682 ( .A(n4191), .B(n4190), .Z(n4189) );
  AND U4683 ( .A(n5522), .B(n5523), .Z(n4190) );
  XOR U4684 ( .A(n4193), .B(n4192), .Z(n4191) );
  AND U4685 ( .A(n5524), .B(n5525), .Z(n4192) );
  XOR U4686 ( .A(n4195), .B(n4194), .Z(n4193) );
  AND U4687 ( .A(n5526), .B(n5527), .Z(n4194) );
  XOR U4688 ( .A(n4197), .B(n4196), .Z(n4195) );
  AND U4689 ( .A(n5528), .B(n5529), .Z(n4196) );
  XOR U4690 ( .A(n4199), .B(n4198), .Z(n4197) );
  AND U4691 ( .A(n5530), .B(n5531), .Z(n4198) );
  XOR U4692 ( .A(n4201), .B(n4200), .Z(n4199) );
  AND U4693 ( .A(n5532), .B(n5533), .Z(n4200) );
  XOR U4694 ( .A(n4203), .B(n4202), .Z(n4201) );
  AND U4695 ( .A(n5534), .B(n5535), .Z(n4202) );
  XOR U4696 ( .A(n4205), .B(n4204), .Z(n4203) );
  AND U4697 ( .A(n5536), .B(n5537), .Z(n4204) );
  XOR U4698 ( .A(n4207), .B(n4206), .Z(n4205) );
  AND U4699 ( .A(n5538), .B(n5539), .Z(n4206) );
  XOR U4700 ( .A(n4209), .B(n4208), .Z(n4207) );
  AND U4701 ( .A(n5540), .B(n5541), .Z(n4208) );
  XOR U4702 ( .A(n4211), .B(n4210), .Z(n4209) );
  AND U4703 ( .A(n5542), .B(n5543), .Z(n4210) );
  XOR U4704 ( .A(n4213), .B(n4212), .Z(n4211) );
  AND U4705 ( .A(n5544), .B(n5545), .Z(n4212) );
  XOR U4706 ( .A(n4215), .B(n4214), .Z(n4213) );
  AND U4707 ( .A(n5546), .B(n5547), .Z(n4214) );
  XOR U4708 ( .A(n4217), .B(n4216), .Z(n4215) );
  AND U4709 ( .A(n5548), .B(n5549), .Z(n4216) );
  XOR U4710 ( .A(n4219), .B(n4218), .Z(n4217) );
  AND U4711 ( .A(n5550), .B(n5551), .Z(n4218) );
  XOR U4712 ( .A(n4221), .B(n4220), .Z(n4219) );
  AND U4713 ( .A(n5552), .B(n5553), .Z(n4220) );
  XOR U4714 ( .A(n4223), .B(n4222), .Z(n4221) );
  AND U4715 ( .A(n5554), .B(n5555), .Z(n4222) );
  XOR U4716 ( .A(n4225), .B(n4224), .Z(n4223) );
  AND U4717 ( .A(n5556), .B(n5557), .Z(n4224) );
  XOR U4718 ( .A(n4227), .B(n4226), .Z(n4225) );
  AND U4719 ( .A(n5558), .B(n5559), .Z(n4226) );
  XOR U4720 ( .A(n4229), .B(n4228), .Z(n4227) );
  AND U4721 ( .A(n5560), .B(n5561), .Z(n4228) );
  XOR U4722 ( .A(n4231), .B(n4230), .Z(n4229) );
  AND U4723 ( .A(n5562), .B(n5563), .Z(n4230) );
  XOR U4724 ( .A(n4233), .B(n4232), .Z(n4231) );
  AND U4725 ( .A(n5564), .B(n5565), .Z(n4232) );
  XOR U4726 ( .A(n4235), .B(n4234), .Z(n4233) );
  AND U4727 ( .A(n5566), .B(n5567), .Z(n4234) );
  XOR U4728 ( .A(n4244), .B(n4236), .Z(n4235) );
  AND U4729 ( .A(n5568), .B(n5569), .Z(n4236) );
  XOR U4730 ( .A(n4239), .B(n4245), .Z(n4244) );
  AND U4731 ( .A(n5570), .B(n5571), .Z(n4245) );
  XOR U4732 ( .A(n4241), .B(n4240), .Z(n4239) );
  AND U4733 ( .A(n5572), .B(n5573), .Z(n4240) );
  XOR U4734 ( .A(n4265), .B(n4242), .Z(n4241) );
  AND U4735 ( .A(n5574), .B(n5575), .Z(n4242) );
  XOR U4736 ( .A(n4260), .B(n4266), .Z(n4265) );
  AND U4737 ( .A(n5576), .B(n5577), .Z(n4266) );
  XOR U4738 ( .A(n4262), .B(n4261), .Z(n4260) );
  AND U4739 ( .A(n5578), .B(n5579), .Z(n4261) );
  XOR U4740 ( .A(n4250), .B(n4263), .Z(n4262) );
  AND U4741 ( .A(n5580), .B(n5581), .Z(n4263) );
  XOR U4742 ( .A(n4252), .B(n4251), .Z(n4250) );
  AND U4743 ( .A(n5582), .B(n5583), .Z(n4251) );
  XOR U4744 ( .A(n4254), .B(n4253), .Z(n4252) );
  AND U4745 ( .A(n5584), .B(n5585), .Z(n4253) );
  XOR U4746 ( .A(n4256), .B(n4255), .Z(n4254) );
  AND U4747 ( .A(n5586), .B(n5587), .Z(n4255) );
  XOR U4748 ( .A(n4286), .B(n4257), .Z(n4256) );
  AND U4749 ( .A(n5588), .B(n5589), .Z(n4257) );
  XOR U4750 ( .A(n4282), .B(n4287), .Z(n4286) );
  AND U4751 ( .A(n5590), .B(n5591), .Z(n4287) );
  XOR U4752 ( .A(n4284), .B(n4283), .Z(n4282) );
  AND U4753 ( .A(n5592), .B(n5593), .Z(n4283) );
  XOR U4754 ( .A(n4271), .B(n4285), .Z(n4284) );
  AND U4755 ( .A(n5594), .B(n5595), .Z(n4285) );
  XOR U4756 ( .A(n4273), .B(n4272), .Z(n4271) );
  AND U4757 ( .A(n5596), .B(n5597), .Z(n4272) );
  XOR U4758 ( .A(n4276), .B(n4274), .Z(n4273) );
  AND U4759 ( .A(n5598), .B(n5599), .Z(n4274) );
  XOR U4760 ( .A(n4278), .B(n4277), .Z(n4276) );
  AND U4761 ( .A(n5600), .B(n5601), .Z(n4277) );
  XOR U4762 ( .A(n4296), .B(n4279), .Z(n4278) );
  AND U4763 ( .A(n5602), .B(n5603), .Z(n4279) );
  XNOR U4764 ( .A(n4303), .B(n4297), .Z(n4296) );
  AND U4765 ( .A(n5604), .B(n5605), .Z(n4297) );
  XOR U4766 ( .A(n4302), .B(n4294), .Z(n4303) );
  AND U4767 ( .A(n5606), .B(n5607), .Z(n4294) );
  XOR U4768 ( .A(n4341), .B(n4293), .Z(n4302) );
  AND U4769 ( .A(n5608), .B(n5609), .Z(n4293) );
  XNOR U4770 ( .A(n4314), .B(n4292), .Z(n4341) );
  AND U4771 ( .A(n5610), .B(n5611), .Z(n4292) );
  XNOR U4772 ( .A(n4321), .B(n4315), .Z(n4314) );
  AND U4773 ( .A(n5612), .B(n5613), .Z(n4315) );
  XOR U4774 ( .A(n4320), .B(n4312), .Z(n4321) );
  AND U4775 ( .A(n5614), .B(n5615), .Z(n4312) );
  XOR U4776 ( .A(n4340), .B(n4311), .Z(n4320) );
  AND U4777 ( .A(n5616), .B(n5617), .Z(n4311) );
  XNOR U4778 ( .A(n5618), .B(n5619), .Z(n4340) );
  XOR U4779 ( .A(n5620), .B(n5621), .Z(n5619) );
  XOR U4780 ( .A(n5622), .B(n5623), .Z(n5621) );
  XNOR U4781 ( .A(n4338), .B(n4331), .Z(n5623) );
  XNOR U4782 ( .A(n5624), .B(n5625), .Z(n4331) );
  AND U4783 ( .A(n5626), .B(n5627), .Z(n5625) );
  NOR U4784 ( .A(n5628), .B(n5629), .Z(n5627) );
  NOR U4785 ( .A(n5630), .B(n5631), .Z(n5626) );
  AND U4786 ( .A(n5632), .B(n5633), .Z(n5631) );
  AND U4787 ( .A(n5634), .B(n5635), .Z(n5624) );
  NOR U4788 ( .A(n5636), .B(n5637), .Z(n5635) );
  AND U4789 ( .A(n5629), .B(n5638), .Z(n5637) );
  AND U4790 ( .A(n5630), .B(n5639), .Z(n5636) );
  NOR U4791 ( .A(n5640), .B(n5641), .Z(n5634) );
  AND U4792 ( .A(n5642), .B(n5643), .Z(n5641) );
  NOR U4793 ( .A(n5644), .B(n5645), .Z(n5643) );
  IV U4794 ( .A(n5646), .Z(n5644) );
  NOR U4795 ( .A(n5647), .B(n5648), .Z(n5646) );
  NOR U4796 ( .A(n5649), .B(n5650), .Z(n5642) );
  AND U4797 ( .A(n5628), .B(n5651), .Z(n5640) );
  AND U4798 ( .A(n5652), .B(n5653), .Z(n4338) );
  XOR U4799 ( .A(n4336), .B(n4337), .Z(n5622) );
  AND U4800 ( .A(n5654), .B(n5655), .Z(n4337) );
  AND U4801 ( .A(n5656), .B(n5657), .Z(n4336) );
  XOR U4802 ( .A(n5658), .B(n5659), .Z(n5620) );
  XOR U4803 ( .A(n4332), .B(n4333), .Z(n5659) );
  AND U4804 ( .A(n5660), .B(n5661), .Z(n4333) );
  AND U4805 ( .A(n5662), .B(n5663), .Z(n4332) );
  XNOR U4806 ( .A(n4330), .B(n4329), .Z(n5658) );
  IV U4807 ( .A(n5664), .Z(n4329) );
  AND U4808 ( .A(n5665), .B(n5666), .Z(n5664) );
  AND U4809 ( .A(n5667), .B(n5668), .Z(n4330) );
  XNOR U4810 ( .A(n4339), .B(n4310), .Z(n5618) );
  AND U4811 ( .A(n5669), .B(n5670), .Z(n4310) );
  AND U4812 ( .A(n5671), .B(n5672), .Z(n4339) );
  XOR U4813 ( .A(n5673), .B(n5674), .Z(n4354) );
  AND U4814 ( .A(n5673), .B(n5675), .Z(n5674) );
  XNOR U4815 ( .A(n5676), .B(n5677), .Z(n4357) );
  AND U4816 ( .A(n5676), .B(n5678), .Z(n5677) );
  XNOR U4817 ( .A(n5679), .B(n5680), .Z(n4360) );
  AND U4818 ( .A(n5679), .B(n5681), .Z(n5680) );
  XNOR U4819 ( .A(n5682), .B(n5683), .Z(n4363) );
  AND U4820 ( .A(n5682), .B(n5684), .Z(n5683) );
  XNOR U4821 ( .A(n5685), .B(n5686), .Z(n4366) );
  AND U4822 ( .A(n5687), .B(n5685), .Z(n5686) );
  XOR U4823 ( .A(n5688), .B(n5689), .Z(n4369) );
  NOR U4824 ( .A(n5690), .B(n5688), .Z(n5689) );
  XOR U4825 ( .A(n5691), .B(n5692), .Z(n4372) );
  NOR U4826 ( .A(n5693), .B(n5691), .Z(n5692) );
  XOR U4827 ( .A(n5694), .B(n5695), .Z(n4375) );
  NOR U4828 ( .A(n5696), .B(n5694), .Z(n5695) );
  XOR U4829 ( .A(n5697), .B(n5698), .Z(n4378) );
  NOR U4830 ( .A(n5699), .B(n5697), .Z(n5698) );
  XOR U4831 ( .A(n5700), .B(n5701), .Z(n4381) );
  NOR U4832 ( .A(n5702), .B(n5700), .Z(n5701) );
  XOR U4833 ( .A(n5703), .B(n5704), .Z(n4384) );
  NOR U4834 ( .A(n5705), .B(n5703), .Z(n5704) );
  XOR U4835 ( .A(n5706), .B(n5707), .Z(n4387) );
  NOR U4836 ( .A(n5708), .B(n5706), .Z(n5707) );
  XOR U4837 ( .A(n5709), .B(n5710), .Z(n4390) );
  NOR U4838 ( .A(n5711), .B(n5709), .Z(n5710) );
  XOR U4839 ( .A(n5712), .B(n5713), .Z(n4393) );
  NOR U4840 ( .A(n5714), .B(n5712), .Z(n5713) );
  XOR U4841 ( .A(n5715), .B(n5716), .Z(n4396) );
  NOR U4842 ( .A(n5717), .B(n5715), .Z(n5716) );
  XOR U4843 ( .A(n5718), .B(n5719), .Z(n4399) );
  NOR U4844 ( .A(n5720), .B(n5718), .Z(n5719) );
  XOR U4845 ( .A(n5721), .B(n5722), .Z(n4402) );
  NOR U4846 ( .A(n5723), .B(n5721), .Z(n5722) );
  XOR U4847 ( .A(n5724), .B(n5725), .Z(n4405) );
  NOR U4848 ( .A(n5726), .B(n5724), .Z(n5725) );
  XOR U4849 ( .A(n5727), .B(n5728), .Z(n4408) );
  NOR U4850 ( .A(n5729), .B(n5727), .Z(n5728) );
  XOR U4851 ( .A(n5730), .B(n5731), .Z(n4411) );
  NOR U4852 ( .A(n5732), .B(n5730), .Z(n5731) );
  XOR U4853 ( .A(n5733), .B(n5734), .Z(n4414) );
  NOR U4854 ( .A(n5735), .B(n5733), .Z(n5734) );
  XOR U4855 ( .A(n5736), .B(n5737), .Z(n4417) );
  NOR U4856 ( .A(n5738), .B(n5736), .Z(n5737) );
  XOR U4857 ( .A(n5739), .B(n5740), .Z(n4420) );
  NOR U4858 ( .A(n5741), .B(n5739), .Z(n5740) );
  XOR U4859 ( .A(n5742), .B(n5743), .Z(n4423) );
  NOR U4860 ( .A(n5744), .B(n5742), .Z(n5743) );
  XOR U4861 ( .A(n5745), .B(n5746), .Z(n4426) );
  NOR U4862 ( .A(n5747), .B(n5745), .Z(n5746) );
  XOR U4863 ( .A(n5748), .B(n5749), .Z(n4429) );
  NOR U4864 ( .A(n5750), .B(n5748), .Z(n5749) );
  XOR U4865 ( .A(n5751), .B(n5752), .Z(n4432) );
  NOR U4866 ( .A(n5753), .B(n5751), .Z(n5752) );
  XOR U4867 ( .A(n5754), .B(n5755), .Z(n4435) );
  NOR U4868 ( .A(n5756), .B(n5754), .Z(n5755) );
  XOR U4869 ( .A(n5757), .B(n5758), .Z(n4438) );
  NOR U4870 ( .A(n5759), .B(n5757), .Z(n5758) );
  XOR U4871 ( .A(n5760), .B(n5761), .Z(n4441) );
  NOR U4872 ( .A(n5762), .B(n5760), .Z(n5761) );
  XOR U4873 ( .A(n5763), .B(n5764), .Z(n4444) );
  NOR U4874 ( .A(n5765), .B(n5763), .Z(n5764) );
  XOR U4875 ( .A(n5766), .B(n5767), .Z(n4447) );
  NOR U4876 ( .A(n5768), .B(n5766), .Z(n5767) );
  XOR U4877 ( .A(n5769), .B(n5770), .Z(n4450) );
  NOR U4878 ( .A(n5771), .B(n5769), .Z(n5770) );
  XOR U4879 ( .A(n5772), .B(n5773), .Z(n4453) );
  NOR U4880 ( .A(n5774), .B(n5772), .Z(n5773) );
  XOR U4881 ( .A(n5775), .B(n5776), .Z(n4456) );
  NOR U4882 ( .A(n5777), .B(n5775), .Z(n5776) );
  XOR U4883 ( .A(n5778), .B(n5779), .Z(n4459) );
  NOR U4884 ( .A(n5780), .B(n5778), .Z(n5779) );
  XOR U4885 ( .A(n5781), .B(n5782), .Z(n4462) );
  NOR U4886 ( .A(n5783), .B(n5781), .Z(n5782) );
  XOR U4887 ( .A(n5784), .B(n5785), .Z(n4465) );
  NOR U4888 ( .A(n5786), .B(n5784), .Z(n5785) );
  XOR U4889 ( .A(n5787), .B(n5788), .Z(n4468) );
  NOR U4890 ( .A(n5789), .B(n5787), .Z(n5788) );
  XOR U4891 ( .A(n5790), .B(n5791), .Z(n4471) );
  NOR U4892 ( .A(n5792), .B(n5790), .Z(n5791) );
  XOR U4893 ( .A(n5793), .B(n5794), .Z(n4474) );
  NOR U4894 ( .A(n5795), .B(n5793), .Z(n5794) );
  XOR U4895 ( .A(n5796), .B(n5797), .Z(n4477) );
  NOR U4896 ( .A(n5798), .B(n5796), .Z(n5797) );
  XOR U4897 ( .A(n5799), .B(n5800), .Z(n4480) );
  NOR U4898 ( .A(n5801), .B(n5799), .Z(n5800) );
  XOR U4899 ( .A(n5802), .B(n5803), .Z(n4483) );
  NOR U4900 ( .A(n5804), .B(n5802), .Z(n5803) );
  XOR U4901 ( .A(n5805), .B(n5806), .Z(n4486) );
  NOR U4902 ( .A(n5807), .B(n5805), .Z(n5806) );
  XOR U4903 ( .A(n5808), .B(n5809), .Z(n4489) );
  NOR U4904 ( .A(n5810), .B(n5808), .Z(n5809) );
  XOR U4905 ( .A(n5811), .B(n5812), .Z(n4492) );
  NOR U4906 ( .A(n5813), .B(n5811), .Z(n5812) );
  XOR U4907 ( .A(n5814), .B(n5815), .Z(n4495) );
  NOR U4908 ( .A(n5816), .B(n5814), .Z(n5815) );
  XOR U4909 ( .A(n5817), .B(n5818), .Z(n4498) );
  NOR U4910 ( .A(n5819), .B(n5817), .Z(n5818) );
  XOR U4911 ( .A(n5820), .B(n5821), .Z(n4501) );
  NOR U4912 ( .A(n5822), .B(n5820), .Z(n5821) );
  XOR U4913 ( .A(n5823), .B(n5824), .Z(n4504) );
  NOR U4914 ( .A(n5825), .B(n5823), .Z(n5824) );
  XOR U4915 ( .A(n5826), .B(n5827), .Z(n4507) );
  NOR U4916 ( .A(n5828), .B(n5826), .Z(n5827) );
  XOR U4917 ( .A(n5829), .B(n5830), .Z(n4510) );
  NOR U4918 ( .A(n5831), .B(n5829), .Z(n5830) );
  XOR U4919 ( .A(n5832), .B(n5833), .Z(n4513) );
  NOR U4920 ( .A(n5834), .B(n5832), .Z(n5833) );
  XOR U4921 ( .A(n5835), .B(n5836), .Z(n4516) );
  NOR U4922 ( .A(n5837), .B(n5835), .Z(n5836) );
  XOR U4923 ( .A(n5838), .B(n5839), .Z(n4519) );
  NOR U4924 ( .A(n5840), .B(n5838), .Z(n5839) );
  XOR U4925 ( .A(n5841), .B(n5842), .Z(n4522) );
  NOR U4926 ( .A(n5843), .B(n5841), .Z(n5842) );
  XOR U4927 ( .A(n5844), .B(n5845), .Z(n4525) );
  NOR U4928 ( .A(n5846), .B(n5844), .Z(n5845) );
  XOR U4929 ( .A(n5847), .B(n5848), .Z(n4528) );
  NOR U4930 ( .A(n5849), .B(n5847), .Z(n5848) );
  XOR U4931 ( .A(n5850), .B(n5851), .Z(n4531) );
  NOR U4932 ( .A(n5852), .B(n5850), .Z(n5851) );
  XOR U4933 ( .A(n5853), .B(n5854), .Z(n4534) );
  NOR U4934 ( .A(n5855), .B(n5853), .Z(n5854) );
  XOR U4935 ( .A(n5856), .B(n5857), .Z(n4537) );
  NOR U4936 ( .A(n5858), .B(n5856), .Z(n5857) );
  XOR U4937 ( .A(n5859), .B(n5860), .Z(n4540) );
  NOR U4938 ( .A(n5861), .B(n5859), .Z(n5860) );
  XOR U4939 ( .A(n5862), .B(n5863), .Z(n4543) );
  NOR U4940 ( .A(n5864), .B(n5862), .Z(n5863) );
  XOR U4941 ( .A(n5865), .B(n5866), .Z(n4546) );
  NOR U4942 ( .A(n5867), .B(n5865), .Z(n5866) );
  XOR U4943 ( .A(n5868), .B(n5869), .Z(n4549) );
  NOR U4944 ( .A(n5870), .B(n5868), .Z(n5869) );
  XOR U4945 ( .A(n5871), .B(n5872), .Z(n4552) );
  NOR U4946 ( .A(n5873), .B(n5871), .Z(n5872) );
  XOR U4947 ( .A(n5874), .B(n5875), .Z(n4555) );
  NOR U4948 ( .A(n5876), .B(n5874), .Z(n5875) );
  XOR U4949 ( .A(n5877), .B(n5878), .Z(n4558) );
  NOR U4950 ( .A(n5879), .B(n5877), .Z(n5878) );
  XOR U4951 ( .A(n5880), .B(n5881), .Z(n4561) );
  NOR U4952 ( .A(n5882), .B(n5880), .Z(n5881) );
  XOR U4953 ( .A(n5883), .B(n5884), .Z(n4564) );
  NOR U4954 ( .A(n5885), .B(n5883), .Z(n5884) );
  XOR U4955 ( .A(n5886), .B(n5887), .Z(n4567) );
  NOR U4956 ( .A(n5888), .B(n5886), .Z(n5887) );
  XOR U4957 ( .A(n5889), .B(n5890), .Z(n4570) );
  NOR U4958 ( .A(n5891), .B(n5889), .Z(n5890) );
  XOR U4959 ( .A(n5892), .B(n5893), .Z(n4573) );
  NOR U4960 ( .A(n5894), .B(n5892), .Z(n5893) );
  XOR U4961 ( .A(n5895), .B(n5896), .Z(n4576) );
  NOR U4962 ( .A(n5897), .B(n5895), .Z(n5896) );
  XOR U4963 ( .A(n5898), .B(n5899), .Z(n4579) );
  NOR U4964 ( .A(n5900), .B(n5898), .Z(n5899) );
  XOR U4965 ( .A(n5901), .B(n5902), .Z(n4582) );
  NOR U4966 ( .A(n5903), .B(n5901), .Z(n5902) );
  XOR U4967 ( .A(n5904), .B(n5905), .Z(n4585) );
  NOR U4968 ( .A(n5906), .B(n5904), .Z(n5905) );
  XOR U4969 ( .A(n5907), .B(n5908), .Z(n4588) );
  NOR U4970 ( .A(n5909), .B(n5907), .Z(n5908) );
  XOR U4971 ( .A(n5910), .B(n5911), .Z(n4591) );
  NOR U4972 ( .A(n5912), .B(n5910), .Z(n5911) );
  XOR U4973 ( .A(n5913), .B(n5914), .Z(n4594) );
  NOR U4974 ( .A(n5915), .B(n5913), .Z(n5914) );
  XOR U4975 ( .A(n5916), .B(n5917), .Z(n4597) );
  NOR U4976 ( .A(n5918), .B(n5916), .Z(n5917) );
  XOR U4977 ( .A(n5919), .B(n5920), .Z(n4600) );
  NOR U4978 ( .A(n5921), .B(n5919), .Z(n5920) );
  XOR U4979 ( .A(n5922), .B(n5923), .Z(n4603) );
  NOR U4980 ( .A(n5924), .B(n5922), .Z(n5923) );
  XOR U4981 ( .A(n5925), .B(n5926), .Z(n4606) );
  NOR U4982 ( .A(n5927), .B(n5925), .Z(n5926) );
  XOR U4983 ( .A(n5928), .B(n5929), .Z(n4609) );
  NOR U4984 ( .A(n5930), .B(n5928), .Z(n5929) );
  XOR U4985 ( .A(n5931), .B(n5932), .Z(n4612) );
  NOR U4986 ( .A(n5933), .B(n5931), .Z(n5932) );
  XOR U4987 ( .A(n5934), .B(n5935), .Z(n4615) );
  NOR U4988 ( .A(n5936), .B(n5934), .Z(n5935) );
  XOR U4989 ( .A(n5937), .B(n5938), .Z(n4618) );
  NOR U4990 ( .A(n5939), .B(n5937), .Z(n5938) );
  XOR U4991 ( .A(n5940), .B(n5941), .Z(n4621) );
  NOR U4992 ( .A(n5942), .B(n5940), .Z(n5941) );
  XOR U4993 ( .A(n5943), .B(n5944), .Z(n4624) );
  NOR U4994 ( .A(n5945), .B(n5943), .Z(n5944) );
  XOR U4995 ( .A(n5946), .B(n5947), .Z(n4627) );
  NOR U4996 ( .A(n5948), .B(n5946), .Z(n5947) );
  XOR U4997 ( .A(n5949), .B(n5950), .Z(n4630) );
  NOR U4998 ( .A(n5951), .B(n5949), .Z(n5950) );
  XOR U4999 ( .A(n5952), .B(n5953), .Z(n4633) );
  NOR U5000 ( .A(n5954), .B(n5952), .Z(n5953) );
  XOR U5001 ( .A(n5955), .B(n5956), .Z(n4636) );
  NOR U5002 ( .A(n5957), .B(n5955), .Z(n5956) );
  XOR U5003 ( .A(n5958), .B(n5959), .Z(n4639) );
  NOR U5004 ( .A(n5960), .B(n5958), .Z(n5959) );
  XOR U5005 ( .A(n5961), .B(n5962), .Z(n4642) );
  NOR U5006 ( .A(n5963), .B(n5961), .Z(n5962) );
  XOR U5007 ( .A(n5964), .B(n5965), .Z(n4645) );
  NOR U5008 ( .A(n5966), .B(n5964), .Z(n5965) );
  XOR U5009 ( .A(n5967), .B(n5968), .Z(n4648) );
  NOR U5010 ( .A(n5969), .B(n5967), .Z(n5968) );
  XOR U5011 ( .A(n5970), .B(n5971), .Z(n4651) );
  NOR U5012 ( .A(n5972), .B(n5970), .Z(n5971) );
  XOR U5013 ( .A(n5973), .B(n5974), .Z(n4654) );
  NOR U5014 ( .A(n5975), .B(n5973), .Z(n5974) );
  XOR U5015 ( .A(n5976), .B(n5977), .Z(n4657) );
  NOR U5016 ( .A(n5978), .B(n5976), .Z(n5977) );
  XOR U5017 ( .A(n5979), .B(n5980), .Z(n4660) );
  NOR U5018 ( .A(n5981), .B(n5979), .Z(n5980) );
  XOR U5019 ( .A(n5982), .B(n5983), .Z(n4663) );
  NOR U5020 ( .A(n5984), .B(n5982), .Z(n5983) );
  XOR U5021 ( .A(n5985), .B(n5986), .Z(n4666) );
  NOR U5022 ( .A(n5987), .B(n5985), .Z(n5986) );
  XOR U5023 ( .A(n5988), .B(n5989), .Z(n4669) );
  NOR U5024 ( .A(n5990), .B(n5988), .Z(n5989) );
  XOR U5025 ( .A(n5991), .B(n5992), .Z(n4672) );
  NOR U5026 ( .A(n5993), .B(n5991), .Z(n5992) );
  XOR U5027 ( .A(n5994), .B(n5995), .Z(n4675) );
  NOR U5028 ( .A(n5996), .B(n5994), .Z(n5995) );
  XOR U5029 ( .A(n5997), .B(n5998), .Z(n4678) );
  NOR U5030 ( .A(n5999), .B(n5997), .Z(n5998) );
  XOR U5031 ( .A(n6000), .B(n6001), .Z(n4681) );
  NOR U5032 ( .A(n6002), .B(n6000), .Z(n6001) );
  XOR U5033 ( .A(n6003), .B(n6004), .Z(n4684) );
  NOR U5034 ( .A(n6005), .B(n6003), .Z(n6004) );
  XOR U5035 ( .A(n6006), .B(n6007), .Z(n4687) );
  NOR U5036 ( .A(n6008), .B(n6006), .Z(n6007) );
  XOR U5037 ( .A(n6009), .B(n6010), .Z(n4690) );
  NOR U5038 ( .A(n6011), .B(n6009), .Z(n6010) );
  XOR U5039 ( .A(n6012), .B(n6013), .Z(n4693) );
  NOR U5040 ( .A(n6014), .B(n6012), .Z(n6013) );
  XOR U5041 ( .A(n6015), .B(n6016), .Z(n4696) );
  NOR U5042 ( .A(n6017), .B(n6015), .Z(n6016) );
  XOR U5043 ( .A(n6018), .B(n6019), .Z(n4699) );
  NOR U5044 ( .A(n6020), .B(n6018), .Z(n6019) );
  XOR U5045 ( .A(n6021), .B(n6022), .Z(n4702) );
  NOR U5046 ( .A(n6023), .B(n6021), .Z(n6022) );
  XOR U5047 ( .A(n6024), .B(n6025), .Z(n4705) );
  NOR U5048 ( .A(n6026), .B(n6024), .Z(n6025) );
  XOR U5049 ( .A(n6027), .B(n6028), .Z(n4708) );
  NOR U5050 ( .A(n6029), .B(n6027), .Z(n6028) );
  XOR U5051 ( .A(n6030), .B(n6031), .Z(n4711) );
  NOR U5052 ( .A(n6032), .B(n6030), .Z(n6031) );
  XOR U5053 ( .A(n6033), .B(n6034), .Z(n4714) );
  NOR U5054 ( .A(n6035), .B(n6033), .Z(n6034) );
  XOR U5055 ( .A(n6036), .B(n6037), .Z(n4717) );
  NOR U5056 ( .A(n6038), .B(n6036), .Z(n6037) );
  XOR U5057 ( .A(n6039), .B(n6040), .Z(n4720) );
  NOR U5058 ( .A(n6041), .B(n6039), .Z(n6040) );
  XOR U5059 ( .A(n6042), .B(n6043), .Z(n4723) );
  NOR U5060 ( .A(n6044), .B(n6042), .Z(n6043) );
  XOR U5061 ( .A(n6045), .B(n6046), .Z(n4726) );
  NOR U5062 ( .A(n6047), .B(n6045), .Z(n6046) );
  XOR U5063 ( .A(n6048), .B(n6049), .Z(n4729) );
  NOR U5064 ( .A(n6050), .B(n6048), .Z(n6049) );
  XOR U5065 ( .A(n6051), .B(n6052), .Z(n4732) );
  NOR U5066 ( .A(n6053), .B(n6051), .Z(n6052) );
  XOR U5067 ( .A(n6054), .B(n6055), .Z(n4735) );
  NOR U5068 ( .A(n6056), .B(n6054), .Z(n6055) );
  XOR U5069 ( .A(n6057), .B(n6058), .Z(n4738) );
  NOR U5070 ( .A(n6059), .B(n6057), .Z(n6058) );
  XOR U5071 ( .A(n6060), .B(n6061), .Z(n4741) );
  NOR U5072 ( .A(n6062), .B(n6060), .Z(n6061) );
  XOR U5073 ( .A(n6063), .B(n6064), .Z(n4744) );
  NOR U5074 ( .A(n6065), .B(n6063), .Z(n6064) );
  XOR U5075 ( .A(n6066), .B(n6067), .Z(n4747) );
  NOR U5076 ( .A(n6068), .B(n6066), .Z(n6067) );
  XOR U5077 ( .A(n6069), .B(n6070), .Z(n4750) );
  NOR U5078 ( .A(n6071), .B(n6069), .Z(n6070) );
  XNOR U5079 ( .A(n6072), .B(n6073), .Z(n4753) );
  NOR U5080 ( .A(n6074), .B(n6072), .Z(n6073) );
  XOR U5081 ( .A(n6075), .B(n6076), .Z(n4756) );
  AND U5082 ( .A(n103), .B(n6075), .Z(n6076) );
  XNOR U5083 ( .A(n6077), .B(n5420), .Z(n5422) );
  IV U5084 ( .A(n86), .Z(n6077) );
  XOR U5085 ( .A(n5417), .B(n5416), .Z(n86) );
  XNOR U5086 ( .A(n5414), .B(n5413), .Z(n5416) );
  XNOR U5087 ( .A(n5411), .B(n5410), .Z(n5413) );
  XNOR U5088 ( .A(n5408), .B(n5407), .Z(n5410) );
  XNOR U5089 ( .A(n5405), .B(n5404), .Z(n5407) );
  XNOR U5090 ( .A(n5402), .B(n5401), .Z(n5404) );
  XNOR U5091 ( .A(n5399), .B(n5398), .Z(n5401) );
  XNOR U5092 ( .A(n5396), .B(n5395), .Z(n5398) );
  XNOR U5093 ( .A(n5393), .B(n5392), .Z(n5395) );
  XNOR U5094 ( .A(n5390), .B(n5389), .Z(n5392) );
  XNOR U5095 ( .A(n5387), .B(n5386), .Z(n5389) );
  XNOR U5096 ( .A(n5384), .B(n5383), .Z(n5386) );
  XNOR U5097 ( .A(n5381), .B(n5380), .Z(n5383) );
  XNOR U5098 ( .A(n5378), .B(n5377), .Z(n5380) );
  XNOR U5099 ( .A(n5375), .B(n5374), .Z(n5377) );
  XNOR U5100 ( .A(n5372), .B(n5371), .Z(n5374) );
  XNOR U5101 ( .A(n5369), .B(n5368), .Z(n5371) );
  XNOR U5102 ( .A(n5366), .B(n5365), .Z(n5368) );
  XNOR U5103 ( .A(n5363), .B(n5362), .Z(n5365) );
  XNOR U5104 ( .A(n5360), .B(n5359), .Z(n5362) );
  XNOR U5105 ( .A(n5357), .B(n5356), .Z(n5359) );
  XNOR U5106 ( .A(n5354), .B(n5353), .Z(n5356) );
  XNOR U5107 ( .A(n5351), .B(n5350), .Z(n5353) );
  XNOR U5108 ( .A(n5348), .B(n5347), .Z(n5350) );
  XNOR U5109 ( .A(n5345), .B(n5344), .Z(n5347) );
  XNOR U5110 ( .A(n5342), .B(n5341), .Z(n5344) );
  XNOR U5111 ( .A(n5339), .B(n5338), .Z(n5341) );
  XNOR U5112 ( .A(n5336), .B(n5335), .Z(n5338) );
  XNOR U5113 ( .A(n5333), .B(n5332), .Z(n5335) );
  XNOR U5114 ( .A(n5330), .B(n5329), .Z(n5332) );
  XNOR U5115 ( .A(n5327), .B(n5326), .Z(n5329) );
  XNOR U5116 ( .A(n5324), .B(n5323), .Z(n5326) );
  XNOR U5117 ( .A(n5321), .B(n5320), .Z(n5323) );
  XNOR U5118 ( .A(n5318), .B(n5317), .Z(n5320) );
  XNOR U5119 ( .A(n5315), .B(n5314), .Z(n5317) );
  XNOR U5120 ( .A(n5312), .B(n5311), .Z(n5314) );
  XNOR U5121 ( .A(n5309), .B(n5308), .Z(n5311) );
  XNOR U5122 ( .A(n5306), .B(n5305), .Z(n5308) );
  XNOR U5123 ( .A(n5303), .B(n5302), .Z(n5305) );
  XNOR U5124 ( .A(n5300), .B(n5299), .Z(n5302) );
  XNOR U5125 ( .A(n5297), .B(n5296), .Z(n5299) );
  XNOR U5126 ( .A(n5294), .B(n5293), .Z(n5296) );
  XNOR U5127 ( .A(n5291), .B(n5290), .Z(n5293) );
  XNOR U5128 ( .A(n5288), .B(n5287), .Z(n5290) );
  XNOR U5129 ( .A(n5285), .B(n5284), .Z(n5287) );
  XNOR U5130 ( .A(n5282), .B(n5281), .Z(n5284) );
  XNOR U5131 ( .A(n5279), .B(n5278), .Z(n5281) );
  XNOR U5132 ( .A(n5276), .B(n5275), .Z(n5278) );
  XNOR U5133 ( .A(n5273), .B(n5272), .Z(n5275) );
  XNOR U5134 ( .A(n5270), .B(n5269), .Z(n5272) );
  XNOR U5135 ( .A(n5267), .B(n5266), .Z(n5269) );
  XNOR U5136 ( .A(n5264), .B(n5263), .Z(n5266) );
  XNOR U5137 ( .A(n5261), .B(n5260), .Z(n5263) );
  XNOR U5138 ( .A(n5258), .B(n5257), .Z(n5260) );
  XNOR U5139 ( .A(n5255), .B(n5254), .Z(n5257) );
  XNOR U5140 ( .A(n5252), .B(n5251), .Z(n5254) );
  XNOR U5141 ( .A(n5249), .B(n5248), .Z(n5251) );
  XNOR U5142 ( .A(n5246), .B(n5245), .Z(n5248) );
  XNOR U5143 ( .A(n5243), .B(n5242), .Z(n5245) );
  XNOR U5144 ( .A(n5240), .B(n5239), .Z(n5242) );
  XNOR U5145 ( .A(n5237), .B(n5236), .Z(n5239) );
  XNOR U5146 ( .A(n5234), .B(n5233), .Z(n5236) );
  XNOR U5147 ( .A(n5231), .B(n5230), .Z(n5233) );
  XNOR U5148 ( .A(n5228), .B(n5227), .Z(n5230) );
  XNOR U5149 ( .A(n5225), .B(n5224), .Z(n5227) );
  XNOR U5150 ( .A(n5222), .B(n5221), .Z(n5224) );
  XNOR U5151 ( .A(n5219), .B(n5218), .Z(n5221) );
  XNOR U5152 ( .A(n5216), .B(n5215), .Z(n5218) );
  XNOR U5153 ( .A(n5213), .B(n5212), .Z(n5215) );
  XNOR U5154 ( .A(n5210), .B(n5209), .Z(n5212) );
  XNOR U5155 ( .A(n5207), .B(n5206), .Z(n5209) );
  XNOR U5156 ( .A(n5204), .B(n5203), .Z(n5206) );
  XNOR U5157 ( .A(n5201), .B(n5200), .Z(n5203) );
  XNOR U5158 ( .A(n5198), .B(n5197), .Z(n5200) );
  XNOR U5159 ( .A(n5195), .B(n5194), .Z(n5197) );
  XNOR U5160 ( .A(n5192), .B(n5191), .Z(n5194) );
  XNOR U5161 ( .A(n5189), .B(n5188), .Z(n5191) );
  XNOR U5162 ( .A(n5186), .B(n5185), .Z(n5188) );
  XNOR U5163 ( .A(n5183), .B(n5182), .Z(n5185) );
  XNOR U5164 ( .A(n5180), .B(n5179), .Z(n5182) );
  XNOR U5165 ( .A(n5177), .B(n5176), .Z(n5179) );
  XNOR U5166 ( .A(n5174), .B(n5173), .Z(n5176) );
  XNOR U5167 ( .A(n5171), .B(n5170), .Z(n5173) );
  XNOR U5168 ( .A(n5168), .B(n5167), .Z(n5170) );
  XNOR U5169 ( .A(n5165), .B(n5164), .Z(n5167) );
  XNOR U5170 ( .A(n5162), .B(n5161), .Z(n5164) );
  XNOR U5171 ( .A(n5159), .B(n5158), .Z(n5161) );
  XNOR U5172 ( .A(n5156), .B(n5155), .Z(n5158) );
  XNOR U5173 ( .A(n5153), .B(n5152), .Z(n5155) );
  XNOR U5174 ( .A(n5150), .B(n5149), .Z(n5152) );
  XNOR U5175 ( .A(n5147), .B(n5146), .Z(n5149) );
  XNOR U5176 ( .A(n5144), .B(n5143), .Z(n5146) );
  XNOR U5177 ( .A(n5141), .B(n5140), .Z(n5143) );
  XNOR U5178 ( .A(n5138), .B(n5137), .Z(n5140) );
  XNOR U5179 ( .A(n5135), .B(n5134), .Z(n5137) );
  XNOR U5180 ( .A(n5132), .B(n5131), .Z(n5134) );
  XNOR U5181 ( .A(n5129), .B(n5128), .Z(n5131) );
  XNOR U5182 ( .A(n5126), .B(n5125), .Z(n5128) );
  XNOR U5183 ( .A(n5123), .B(n5122), .Z(n5125) );
  XNOR U5184 ( .A(n5120), .B(n5119), .Z(n5122) );
  XNOR U5185 ( .A(n5117), .B(n5116), .Z(n5119) );
  XNOR U5186 ( .A(n5114), .B(n5113), .Z(n5116) );
  XNOR U5187 ( .A(n5111), .B(n5110), .Z(n5113) );
  XNOR U5188 ( .A(n5108), .B(n5107), .Z(n5110) );
  XNOR U5189 ( .A(n5105), .B(n5104), .Z(n5107) );
  XNOR U5190 ( .A(n5102), .B(n5101), .Z(n5104) );
  XNOR U5191 ( .A(n5099), .B(n5098), .Z(n5101) );
  XNOR U5192 ( .A(n5096), .B(n5095), .Z(n5098) );
  XNOR U5193 ( .A(n5093), .B(n5092), .Z(n5095) );
  XNOR U5194 ( .A(n5090), .B(n5089), .Z(n5092) );
  XNOR U5195 ( .A(n5087), .B(n5086), .Z(n5089) );
  XNOR U5196 ( .A(n5084), .B(n5083), .Z(n5086) );
  XNOR U5197 ( .A(n5081), .B(n5080), .Z(n5083) );
  XNOR U5198 ( .A(n5078), .B(n5077), .Z(n5080) );
  XNOR U5199 ( .A(n5075), .B(n5074), .Z(n5077) );
  XNOR U5200 ( .A(n5072), .B(n5071), .Z(n5074) );
  XNOR U5201 ( .A(n5069), .B(n5068), .Z(n5071) );
  XNOR U5202 ( .A(n5066), .B(n5065), .Z(n5068) );
  XNOR U5203 ( .A(n5063), .B(n5062), .Z(n5065) );
  XNOR U5204 ( .A(n5060), .B(n5059), .Z(n5062) );
  XNOR U5205 ( .A(n5057), .B(n5056), .Z(n5059) );
  XNOR U5206 ( .A(n5054), .B(n5053), .Z(n5056) );
  XNOR U5207 ( .A(n5051), .B(n5050), .Z(n5053) );
  XNOR U5208 ( .A(n5048), .B(n5047), .Z(n5050) );
  XNOR U5209 ( .A(n5045), .B(n5044), .Z(n5047) );
  XNOR U5210 ( .A(n5042), .B(n5041), .Z(n5044) );
  XNOR U5211 ( .A(n5039), .B(n5038), .Z(n5041) );
  XNOR U5212 ( .A(n5036), .B(n5035), .Z(n5038) );
  XNOR U5213 ( .A(n5033), .B(n5032), .Z(n5035) );
  XNOR U5214 ( .A(n5030), .B(n5029), .Z(n5032) );
  XNOR U5215 ( .A(n5027), .B(n5026), .Z(n5029) );
  XNOR U5216 ( .A(n5024), .B(n5023), .Z(n5026) );
  XNOR U5217 ( .A(n5021), .B(n5020), .Z(n5023) );
  XOR U5218 ( .A(n5018), .B(n5017), .Z(n5020) );
  XOR U5219 ( .A(n5015), .B(n5014), .Z(n5017) );
  XOR U5220 ( .A(n5011), .B(n5012), .Z(n5014) );
  AND U5221 ( .A(n6078), .B(n6079), .Z(n5012) );
  XOR U5222 ( .A(n5008), .B(n5009), .Z(n5011) );
  AND U5223 ( .A(n6080), .B(n6081), .Z(n5009) );
  XOR U5224 ( .A(n5005), .B(n5006), .Z(n5008) );
  AND U5225 ( .A(n6082), .B(n6083), .Z(n5006) );
  XNOR U5226 ( .A(n4760), .B(n5003), .Z(n5005) );
  AND U5227 ( .A(n6084), .B(n6085), .Z(n5003) );
  XOR U5228 ( .A(n4762), .B(n4761), .Z(n4760) );
  AND U5229 ( .A(n6086), .B(n6087), .Z(n4761) );
  XOR U5230 ( .A(n4764), .B(n4763), .Z(n4762) );
  AND U5231 ( .A(n6088), .B(n6089), .Z(n4763) );
  XOR U5232 ( .A(n4766), .B(n4765), .Z(n4764) );
  AND U5233 ( .A(n6090), .B(n6091), .Z(n4765) );
  XOR U5234 ( .A(n4768), .B(n4767), .Z(n4766) );
  AND U5235 ( .A(n6092), .B(n6093), .Z(n4767) );
  XOR U5236 ( .A(n4770), .B(n4769), .Z(n4768) );
  AND U5237 ( .A(n6094), .B(n6095), .Z(n4769) );
  XOR U5238 ( .A(n4772), .B(n4771), .Z(n4770) );
  AND U5239 ( .A(n6096), .B(n6097), .Z(n4771) );
  XOR U5240 ( .A(n4774), .B(n4773), .Z(n4772) );
  AND U5241 ( .A(n6098), .B(n6099), .Z(n4773) );
  XOR U5242 ( .A(n4776), .B(n4775), .Z(n4774) );
  AND U5243 ( .A(n6100), .B(n6101), .Z(n4775) );
  XOR U5244 ( .A(n4778), .B(n4777), .Z(n4776) );
  AND U5245 ( .A(n6102), .B(n6103), .Z(n4777) );
  XOR U5246 ( .A(n4780), .B(n4779), .Z(n4778) );
  AND U5247 ( .A(n6104), .B(n6105), .Z(n4779) );
  XOR U5248 ( .A(n4782), .B(n4781), .Z(n4780) );
  AND U5249 ( .A(n6106), .B(n6107), .Z(n4781) );
  XOR U5250 ( .A(n4784), .B(n4783), .Z(n4782) );
  AND U5251 ( .A(n6108), .B(n6109), .Z(n4783) );
  XOR U5252 ( .A(n4786), .B(n4785), .Z(n4784) );
  AND U5253 ( .A(n6110), .B(n6111), .Z(n4785) );
  XOR U5254 ( .A(n4788), .B(n4787), .Z(n4786) );
  AND U5255 ( .A(n6112), .B(n6113), .Z(n4787) );
  XOR U5256 ( .A(n4790), .B(n4789), .Z(n4788) );
  AND U5257 ( .A(n6114), .B(n6115), .Z(n4789) );
  XOR U5258 ( .A(n4792), .B(n4791), .Z(n4790) );
  AND U5259 ( .A(n6116), .B(n6117), .Z(n4791) );
  XOR U5260 ( .A(n4794), .B(n4793), .Z(n4792) );
  AND U5261 ( .A(n6118), .B(n6119), .Z(n4793) );
  XOR U5262 ( .A(n4796), .B(n4795), .Z(n4794) );
  AND U5263 ( .A(n6120), .B(n6121), .Z(n4795) );
  XOR U5264 ( .A(n4798), .B(n4797), .Z(n4796) );
  AND U5265 ( .A(n6122), .B(n6123), .Z(n4797) );
  XOR U5266 ( .A(n4800), .B(n4799), .Z(n4798) );
  AND U5267 ( .A(n6124), .B(n6125), .Z(n4799) );
  XOR U5268 ( .A(n4802), .B(n4801), .Z(n4800) );
  AND U5269 ( .A(n6126), .B(n6127), .Z(n4801) );
  XOR U5270 ( .A(n4804), .B(n4803), .Z(n4802) );
  AND U5271 ( .A(n6128), .B(n6129), .Z(n4803) );
  XOR U5272 ( .A(n4806), .B(n4805), .Z(n4804) );
  AND U5273 ( .A(n6130), .B(n6131), .Z(n4805) );
  XOR U5274 ( .A(n4808), .B(n4807), .Z(n4806) );
  AND U5275 ( .A(n6132), .B(n6133), .Z(n4807) );
  XOR U5276 ( .A(n4810), .B(n4809), .Z(n4808) );
  AND U5277 ( .A(n6134), .B(n6135), .Z(n4809) );
  XOR U5278 ( .A(n4812), .B(n4811), .Z(n4810) );
  AND U5279 ( .A(n6136), .B(n6137), .Z(n4811) );
  XOR U5280 ( .A(n4814), .B(n4813), .Z(n4812) );
  AND U5281 ( .A(n6138), .B(n6139), .Z(n4813) );
  XOR U5282 ( .A(n4816), .B(n4815), .Z(n4814) );
  AND U5283 ( .A(n6140), .B(n6141), .Z(n4815) );
  XOR U5284 ( .A(n4818), .B(n4817), .Z(n4816) );
  AND U5285 ( .A(n6142), .B(n6143), .Z(n4817) );
  XOR U5286 ( .A(n4820), .B(n4819), .Z(n4818) );
  AND U5287 ( .A(n6144), .B(n6145), .Z(n4819) );
  XOR U5288 ( .A(n4822), .B(n4821), .Z(n4820) );
  AND U5289 ( .A(n6146), .B(n6147), .Z(n4821) );
  XOR U5290 ( .A(n4824), .B(n4823), .Z(n4822) );
  AND U5291 ( .A(n6148), .B(n6149), .Z(n4823) );
  XOR U5292 ( .A(n4826), .B(n4825), .Z(n4824) );
  AND U5293 ( .A(n6150), .B(n6151), .Z(n4825) );
  XOR U5294 ( .A(n4828), .B(n4827), .Z(n4826) );
  AND U5295 ( .A(n6152), .B(n6153), .Z(n4827) );
  XOR U5296 ( .A(n4830), .B(n4829), .Z(n4828) );
  AND U5297 ( .A(n6154), .B(n6155), .Z(n4829) );
  XOR U5298 ( .A(n4832), .B(n4831), .Z(n4830) );
  AND U5299 ( .A(n6156), .B(n6157), .Z(n4831) );
  XOR U5300 ( .A(n4834), .B(n4833), .Z(n4832) );
  AND U5301 ( .A(n6158), .B(n6159), .Z(n4833) );
  XOR U5302 ( .A(n4836), .B(n4835), .Z(n4834) );
  AND U5303 ( .A(n6160), .B(n6161), .Z(n4835) );
  XOR U5304 ( .A(n4838), .B(n4837), .Z(n4836) );
  AND U5305 ( .A(n6162), .B(n6163), .Z(n4837) );
  XOR U5306 ( .A(n4840), .B(n4839), .Z(n4838) );
  AND U5307 ( .A(n6164), .B(n6165), .Z(n4839) );
  XOR U5308 ( .A(n4842), .B(n4841), .Z(n4840) );
  AND U5309 ( .A(n6166), .B(n6167), .Z(n4841) );
  XOR U5310 ( .A(n4844), .B(n4843), .Z(n4842) );
  AND U5311 ( .A(n6168), .B(n6169), .Z(n4843) );
  XOR U5312 ( .A(n4846), .B(n4845), .Z(n4844) );
  AND U5313 ( .A(n6170), .B(n6171), .Z(n4845) );
  XOR U5314 ( .A(n4848), .B(n4847), .Z(n4846) );
  AND U5315 ( .A(n6172), .B(n6173), .Z(n4847) );
  XOR U5316 ( .A(n4850), .B(n4849), .Z(n4848) );
  AND U5317 ( .A(n6174), .B(n6175), .Z(n4849) );
  XOR U5318 ( .A(n4852), .B(n4851), .Z(n4850) );
  AND U5319 ( .A(n6176), .B(n6177), .Z(n4851) );
  XOR U5320 ( .A(n4854), .B(n4853), .Z(n4852) );
  AND U5321 ( .A(n6178), .B(n6179), .Z(n4853) );
  XOR U5322 ( .A(n4856), .B(n4855), .Z(n4854) );
  AND U5323 ( .A(n6180), .B(n6181), .Z(n4855) );
  XOR U5324 ( .A(n4858), .B(n4857), .Z(n4856) );
  AND U5325 ( .A(n6182), .B(n6183), .Z(n4857) );
  XOR U5326 ( .A(n4860), .B(n4859), .Z(n4858) );
  AND U5327 ( .A(n6184), .B(n6185), .Z(n4859) );
  XOR U5328 ( .A(n4862), .B(n4861), .Z(n4860) );
  AND U5329 ( .A(n6186), .B(n6187), .Z(n4861) );
  XOR U5330 ( .A(n4864), .B(n4863), .Z(n4862) );
  AND U5331 ( .A(n6188), .B(n6189), .Z(n4863) );
  XOR U5332 ( .A(n4866), .B(n4865), .Z(n4864) );
  AND U5333 ( .A(n6190), .B(n6191), .Z(n4865) );
  XOR U5334 ( .A(n4868), .B(n4867), .Z(n4866) );
  AND U5335 ( .A(n6192), .B(n6193), .Z(n4867) );
  XOR U5336 ( .A(n4870), .B(n4869), .Z(n4868) );
  AND U5337 ( .A(n6194), .B(n6195), .Z(n4869) );
  XOR U5338 ( .A(n4872), .B(n4871), .Z(n4870) );
  AND U5339 ( .A(n6196), .B(n6197), .Z(n4871) );
  XOR U5340 ( .A(n4874), .B(n4873), .Z(n4872) );
  AND U5341 ( .A(n6198), .B(n6199), .Z(n4873) );
  XOR U5342 ( .A(n4876), .B(n4875), .Z(n4874) );
  AND U5343 ( .A(n6200), .B(n6201), .Z(n4875) );
  XOR U5344 ( .A(n4878), .B(n4877), .Z(n4876) );
  AND U5345 ( .A(n6202), .B(n6203), .Z(n4877) );
  XOR U5346 ( .A(n4880), .B(n4879), .Z(n4878) );
  AND U5347 ( .A(n6204), .B(n6205), .Z(n4879) );
  XOR U5348 ( .A(n4882), .B(n4881), .Z(n4880) );
  AND U5349 ( .A(n6206), .B(n6207), .Z(n4881) );
  XOR U5350 ( .A(n4884), .B(n4883), .Z(n4882) );
  AND U5351 ( .A(n6208), .B(n6209), .Z(n4883) );
  XOR U5352 ( .A(n4886), .B(n4885), .Z(n4884) );
  AND U5353 ( .A(n6210), .B(n6211), .Z(n4885) );
  XOR U5354 ( .A(n4888), .B(n4887), .Z(n4886) );
  AND U5355 ( .A(n6212), .B(n6213), .Z(n4887) );
  XOR U5356 ( .A(n4890), .B(n4889), .Z(n4888) );
  AND U5357 ( .A(n6214), .B(n6215), .Z(n4889) );
  XOR U5358 ( .A(n4892), .B(n4891), .Z(n4890) );
  AND U5359 ( .A(n6216), .B(n6217), .Z(n4891) );
  XOR U5360 ( .A(n4894), .B(n4893), .Z(n4892) );
  AND U5361 ( .A(n6218), .B(n6219), .Z(n4893) );
  XOR U5362 ( .A(n4896), .B(n4895), .Z(n4894) );
  AND U5363 ( .A(n6220), .B(n6221), .Z(n4895) );
  XOR U5364 ( .A(n4905), .B(n4897), .Z(n4896) );
  AND U5365 ( .A(n6222), .B(n6223), .Z(n4897) );
  XOR U5366 ( .A(n4900), .B(n4906), .Z(n4905) );
  AND U5367 ( .A(n6224), .B(n6225), .Z(n4906) );
  XOR U5368 ( .A(n4902), .B(n4901), .Z(n4900) );
  AND U5369 ( .A(n6226), .B(n6227), .Z(n4901) );
  XOR U5370 ( .A(n4926), .B(n4903), .Z(n4902) );
  AND U5371 ( .A(n6228), .B(n6229), .Z(n4903) );
  XOR U5372 ( .A(n4921), .B(n4927), .Z(n4926) );
  AND U5373 ( .A(n6230), .B(n6231), .Z(n4927) );
  XOR U5374 ( .A(n4923), .B(n4922), .Z(n4921) );
  AND U5375 ( .A(n6232), .B(n6233), .Z(n4922) );
  XOR U5376 ( .A(n4911), .B(n4924), .Z(n4923) );
  AND U5377 ( .A(n6234), .B(n6235), .Z(n4924) );
  XOR U5378 ( .A(n4913), .B(n4912), .Z(n4911) );
  AND U5379 ( .A(n6236), .B(n6237), .Z(n4912) );
  XOR U5380 ( .A(n4915), .B(n4914), .Z(n4913) );
  AND U5381 ( .A(n6238), .B(n6239), .Z(n4914) );
  XOR U5382 ( .A(n4917), .B(n4916), .Z(n4915) );
  AND U5383 ( .A(n6240), .B(n6241), .Z(n4916) );
  XOR U5384 ( .A(n4946), .B(n4918), .Z(n4917) );
  AND U5385 ( .A(n6242), .B(n6243), .Z(n4918) );
  XOR U5386 ( .A(n4942), .B(n4947), .Z(n4946) );
  AND U5387 ( .A(n6244), .B(n6245), .Z(n4947) );
  XOR U5388 ( .A(n4944), .B(n4943), .Z(n4942) );
  AND U5389 ( .A(n6246), .B(n6247), .Z(n4943) );
  XOR U5390 ( .A(n4932), .B(n4945), .Z(n4944) );
  AND U5391 ( .A(n6248), .B(n6249), .Z(n4945) );
  XOR U5392 ( .A(n4934), .B(n4933), .Z(n4932) );
  AND U5393 ( .A(n6250), .B(n6251), .Z(n4933) );
  XOR U5394 ( .A(n4936), .B(n4935), .Z(n4934) );
  AND U5395 ( .A(n6252), .B(n6253), .Z(n4935) );
  XOR U5396 ( .A(n4938), .B(n4937), .Z(n4936) );
  AND U5397 ( .A(n6254), .B(n6255), .Z(n4937) );
  XOR U5398 ( .A(n4980), .B(n4939), .Z(n4938) );
  AND U5399 ( .A(n6256), .B(n6257), .Z(n4939) );
  XNOR U5400 ( .A(n4977), .B(n4981), .Z(n4980) );
  AND U5401 ( .A(n6258), .B(n6259), .Z(n4981) );
  XOR U5402 ( .A(n4976), .B(n4968), .Z(n4977) );
  AND U5403 ( .A(n6260), .B(n6261), .Z(n4968) );
  XNOR U5404 ( .A(n4971), .B(n4967), .Z(n4976) );
  AND U5405 ( .A(n6262), .B(n6263), .Z(n4967) );
  XOR U5406 ( .A(n4984), .B(n4972), .Z(n4971) );
  AND U5407 ( .A(n6264), .B(n6265), .Z(n4972) );
  XNOR U5408 ( .A(n4964), .B(n4985), .Z(n4984) );
  AND U5409 ( .A(n6266), .B(n6267), .Z(n4985) );
  XOR U5410 ( .A(n4963), .B(n4955), .Z(n4964) );
  AND U5411 ( .A(n6268), .B(n6269), .Z(n4955) );
  XNOR U5412 ( .A(n4958), .B(n4954), .Z(n4963) );
  AND U5413 ( .A(n6270), .B(n6271), .Z(n4954) );
  XOR U5414 ( .A(n6272), .B(n6273), .Z(n4958) );
  XOR U5415 ( .A(n6274), .B(n6275), .Z(n6273) );
  XOR U5416 ( .A(n6276), .B(n6277), .Z(n6275) );
  XNOR U5417 ( .A(n5001), .B(n4994), .Z(n6277) );
  XOR U5418 ( .A(n6278), .B(n6279), .Z(n4994) );
  XOR U5419 ( .A(n6280), .B(n6281), .Z(n6279) );
  NOR U5420 ( .A(n6282), .B(n6283), .Z(n6281) );
  NOR U5421 ( .A(n6284), .B(n6285), .Z(n6280) );
  AND U5422 ( .A(n6286), .B(n6287), .Z(n6285) );
  IV U5423 ( .A(n6288), .Z(n6284) );
  NOR U5424 ( .A(n6289), .B(n6290), .Z(n6288) );
  AND U5425 ( .A(n6282), .B(n6291), .Z(n6290) );
  AND U5426 ( .A(n6283), .B(n6292), .Z(n6289) );
  XNOR U5427 ( .A(n6293), .B(n6294), .Z(n6278) );
  AND U5428 ( .A(n6295), .B(n6296), .Z(n6294) );
  AND U5429 ( .A(n6297), .B(n6298), .Z(n6293) );
  NOR U5430 ( .A(n6299), .B(n6300), .Z(n6298) );
  IV U5431 ( .A(n6301), .Z(n6299) );
  NOR U5432 ( .A(n6302), .B(n6303), .Z(n6301) );
  NOR U5433 ( .A(n6304), .B(n6305), .Z(n6297) );
  AND U5434 ( .A(n6306), .B(n6307), .Z(n5001) );
  XOR U5435 ( .A(n4999), .B(n5000), .Z(n6276) );
  AND U5436 ( .A(n6308), .B(n6309), .Z(n5000) );
  AND U5437 ( .A(n6310), .B(n6311), .Z(n4999) );
  XOR U5438 ( .A(n6312), .B(n6313), .Z(n6274) );
  XOR U5439 ( .A(n4995), .B(n4996), .Z(n6313) );
  AND U5440 ( .A(n6314), .B(n6315), .Z(n4996) );
  AND U5441 ( .A(n6316), .B(n6317), .Z(n4995) );
  XOR U5442 ( .A(n4993), .B(n4991), .Z(n6312) );
  AND U5443 ( .A(n6318), .B(n6319), .Z(n4991) );
  AND U5444 ( .A(n6320), .B(n6321), .Z(n4993) );
  XNOR U5445 ( .A(n5002), .B(n4959), .Z(n6272) );
  AND U5446 ( .A(n6322), .B(n6323), .Z(n4959) );
  AND U5447 ( .A(n6324), .B(n6325), .Z(n5002) );
  XOR U5448 ( .A(n6326), .B(n6327), .Z(n5015) );
  AND U5449 ( .A(n6326), .B(n6328), .Z(n6327) );
  XNOR U5450 ( .A(n6329), .B(n6330), .Z(n5018) );
  AND U5451 ( .A(n6329), .B(n6331), .Z(n6330) );
  XNOR U5452 ( .A(n6332), .B(n6333), .Z(n5021) );
  AND U5453 ( .A(n6332), .B(n6334), .Z(n6333) );
  XNOR U5454 ( .A(n6335), .B(n6336), .Z(n5024) );
  AND U5455 ( .A(n6335), .B(n6337), .Z(n6336) );
  XNOR U5456 ( .A(n6338), .B(n6339), .Z(n5027) );
  AND U5457 ( .A(n6340), .B(n6338), .Z(n6339) );
  XOR U5458 ( .A(n6341), .B(n6342), .Z(n5030) );
  NOR U5459 ( .A(n6343), .B(n6341), .Z(n6342) );
  XOR U5460 ( .A(n6344), .B(n6345), .Z(n5033) );
  NOR U5461 ( .A(n6346), .B(n6344), .Z(n6345) );
  XOR U5462 ( .A(n6347), .B(n6348), .Z(n5036) );
  NOR U5463 ( .A(n6349), .B(n6347), .Z(n6348) );
  XOR U5464 ( .A(n6350), .B(n6351), .Z(n5039) );
  NOR U5465 ( .A(n6352), .B(n6350), .Z(n6351) );
  XOR U5466 ( .A(n6353), .B(n6354), .Z(n5042) );
  NOR U5467 ( .A(n6355), .B(n6353), .Z(n6354) );
  XOR U5468 ( .A(n6356), .B(n6357), .Z(n5045) );
  NOR U5469 ( .A(n6358), .B(n6356), .Z(n6357) );
  XOR U5470 ( .A(n6359), .B(n6360), .Z(n5048) );
  NOR U5471 ( .A(n6361), .B(n6359), .Z(n6360) );
  XOR U5472 ( .A(n6362), .B(n6363), .Z(n5051) );
  NOR U5473 ( .A(n6364), .B(n6362), .Z(n6363) );
  XOR U5474 ( .A(n6365), .B(n6366), .Z(n5054) );
  NOR U5475 ( .A(n6367), .B(n6365), .Z(n6366) );
  XOR U5476 ( .A(n6368), .B(n6369), .Z(n5057) );
  NOR U5477 ( .A(n6370), .B(n6368), .Z(n6369) );
  XOR U5478 ( .A(n6371), .B(n6372), .Z(n5060) );
  NOR U5479 ( .A(n6373), .B(n6371), .Z(n6372) );
  XOR U5480 ( .A(n6374), .B(n6375), .Z(n5063) );
  NOR U5481 ( .A(n6376), .B(n6374), .Z(n6375) );
  XOR U5482 ( .A(n6377), .B(n6378), .Z(n5066) );
  NOR U5483 ( .A(n6379), .B(n6377), .Z(n6378) );
  XOR U5484 ( .A(n6380), .B(n6381), .Z(n5069) );
  NOR U5485 ( .A(n6382), .B(n6380), .Z(n6381) );
  XOR U5486 ( .A(n6383), .B(n6384), .Z(n5072) );
  NOR U5487 ( .A(n6385), .B(n6383), .Z(n6384) );
  XOR U5488 ( .A(n6386), .B(n6387), .Z(n5075) );
  NOR U5489 ( .A(n6388), .B(n6386), .Z(n6387) );
  XOR U5490 ( .A(n6389), .B(n6390), .Z(n5078) );
  NOR U5491 ( .A(n6391), .B(n6389), .Z(n6390) );
  XOR U5492 ( .A(n6392), .B(n6393), .Z(n5081) );
  NOR U5493 ( .A(n6394), .B(n6392), .Z(n6393) );
  XOR U5494 ( .A(n6395), .B(n6396), .Z(n5084) );
  NOR U5495 ( .A(n6397), .B(n6395), .Z(n6396) );
  XOR U5496 ( .A(n6398), .B(n6399), .Z(n5087) );
  NOR U5497 ( .A(n6400), .B(n6398), .Z(n6399) );
  XOR U5498 ( .A(n6401), .B(n6402), .Z(n5090) );
  NOR U5499 ( .A(n6403), .B(n6401), .Z(n6402) );
  XOR U5500 ( .A(n6404), .B(n6405), .Z(n5093) );
  NOR U5501 ( .A(n6406), .B(n6404), .Z(n6405) );
  XOR U5502 ( .A(n6407), .B(n6408), .Z(n5096) );
  NOR U5503 ( .A(n6409), .B(n6407), .Z(n6408) );
  XOR U5504 ( .A(n6410), .B(n6411), .Z(n5099) );
  NOR U5505 ( .A(n6412), .B(n6410), .Z(n6411) );
  XOR U5506 ( .A(n6413), .B(n6414), .Z(n5102) );
  NOR U5507 ( .A(n6415), .B(n6413), .Z(n6414) );
  XOR U5508 ( .A(n6416), .B(n6417), .Z(n5105) );
  NOR U5509 ( .A(n6418), .B(n6416), .Z(n6417) );
  XOR U5510 ( .A(n6419), .B(n6420), .Z(n5108) );
  NOR U5511 ( .A(n6421), .B(n6419), .Z(n6420) );
  XOR U5512 ( .A(n6422), .B(n6423), .Z(n5111) );
  NOR U5513 ( .A(n6424), .B(n6422), .Z(n6423) );
  XOR U5514 ( .A(n6425), .B(n6426), .Z(n5114) );
  NOR U5515 ( .A(n6427), .B(n6425), .Z(n6426) );
  XOR U5516 ( .A(n6428), .B(n6429), .Z(n5117) );
  NOR U5517 ( .A(n6430), .B(n6428), .Z(n6429) );
  XOR U5518 ( .A(n6431), .B(n6432), .Z(n5120) );
  NOR U5519 ( .A(n6433), .B(n6431), .Z(n6432) );
  XOR U5520 ( .A(n6434), .B(n6435), .Z(n5123) );
  NOR U5521 ( .A(n6436), .B(n6434), .Z(n6435) );
  XOR U5522 ( .A(n6437), .B(n6438), .Z(n5126) );
  NOR U5523 ( .A(n6439), .B(n6437), .Z(n6438) );
  XOR U5524 ( .A(n6440), .B(n6441), .Z(n5129) );
  NOR U5525 ( .A(n6442), .B(n6440), .Z(n6441) );
  XOR U5526 ( .A(n6443), .B(n6444), .Z(n5132) );
  NOR U5527 ( .A(n6445), .B(n6443), .Z(n6444) );
  XOR U5528 ( .A(n6446), .B(n6447), .Z(n5135) );
  NOR U5529 ( .A(n6448), .B(n6446), .Z(n6447) );
  XOR U5530 ( .A(n6449), .B(n6450), .Z(n5138) );
  NOR U5531 ( .A(n6451), .B(n6449), .Z(n6450) );
  XOR U5532 ( .A(n6452), .B(n6453), .Z(n5141) );
  NOR U5533 ( .A(n6454), .B(n6452), .Z(n6453) );
  XOR U5534 ( .A(n6455), .B(n6456), .Z(n5144) );
  NOR U5535 ( .A(n6457), .B(n6455), .Z(n6456) );
  XOR U5536 ( .A(n6458), .B(n6459), .Z(n5147) );
  NOR U5537 ( .A(n6460), .B(n6458), .Z(n6459) );
  XOR U5538 ( .A(n6461), .B(n6462), .Z(n5150) );
  NOR U5539 ( .A(n6463), .B(n6461), .Z(n6462) );
  XOR U5540 ( .A(n6464), .B(n6465), .Z(n5153) );
  NOR U5541 ( .A(n6466), .B(n6464), .Z(n6465) );
  XOR U5542 ( .A(n6467), .B(n6468), .Z(n5156) );
  NOR U5543 ( .A(n6469), .B(n6467), .Z(n6468) );
  XOR U5544 ( .A(n6470), .B(n6471), .Z(n5159) );
  NOR U5545 ( .A(n6472), .B(n6470), .Z(n6471) );
  XOR U5546 ( .A(n6473), .B(n6474), .Z(n5162) );
  NOR U5547 ( .A(n6475), .B(n6473), .Z(n6474) );
  XOR U5548 ( .A(n6476), .B(n6477), .Z(n5165) );
  NOR U5549 ( .A(n6478), .B(n6476), .Z(n6477) );
  XOR U5550 ( .A(n6479), .B(n6480), .Z(n5168) );
  NOR U5551 ( .A(n6481), .B(n6479), .Z(n6480) );
  XOR U5552 ( .A(n6482), .B(n6483), .Z(n5171) );
  NOR U5553 ( .A(n6484), .B(n6482), .Z(n6483) );
  XOR U5554 ( .A(n6485), .B(n6486), .Z(n5174) );
  NOR U5555 ( .A(n6487), .B(n6485), .Z(n6486) );
  XOR U5556 ( .A(n6488), .B(n6489), .Z(n5177) );
  NOR U5557 ( .A(n6490), .B(n6488), .Z(n6489) );
  XOR U5558 ( .A(n6491), .B(n6492), .Z(n5180) );
  NOR U5559 ( .A(n6493), .B(n6491), .Z(n6492) );
  XOR U5560 ( .A(n6494), .B(n6495), .Z(n5183) );
  NOR U5561 ( .A(n6496), .B(n6494), .Z(n6495) );
  XOR U5562 ( .A(n6497), .B(n6498), .Z(n5186) );
  NOR U5563 ( .A(n6499), .B(n6497), .Z(n6498) );
  XOR U5564 ( .A(n6500), .B(n6501), .Z(n5189) );
  NOR U5565 ( .A(n6502), .B(n6500), .Z(n6501) );
  XOR U5566 ( .A(n6503), .B(n6504), .Z(n5192) );
  NOR U5567 ( .A(n6505), .B(n6503), .Z(n6504) );
  XOR U5568 ( .A(n6506), .B(n6507), .Z(n5195) );
  NOR U5569 ( .A(n6508), .B(n6506), .Z(n6507) );
  XOR U5570 ( .A(n6509), .B(n6510), .Z(n5198) );
  NOR U5571 ( .A(n6511), .B(n6509), .Z(n6510) );
  XOR U5572 ( .A(n6512), .B(n6513), .Z(n5201) );
  NOR U5573 ( .A(n6514), .B(n6512), .Z(n6513) );
  XOR U5574 ( .A(n6515), .B(n6516), .Z(n5204) );
  NOR U5575 ( .A(n6517), .B(n6515), .Z(n6516) );
  XOR U5576 ( .A(n6518), .B(n6519), .Z(n5207) );
  NOR U5577 ( .A(n6520), .B(n6518), .Z(n6519) );
  XOR U5578 ( .A(n6521), .B(n6522), .Z(n5210) );
  NOR U5579 ( .A(n6523), .B(n6521), .Z(n6522) );
  XOR U5580 ( .A(n6524), .B(n6525), .Z(n5213) );
  NOR U5581 ( .A(n6526), .B(n6524), .Z(n6525) );
  XOR U5582 ( .A(n6527), .B(n6528), .Z(n5216) );
  NOR U5583 ( .A(n6529), .B(n6527), .Z(n6528) );
  XOR U5584 ( .A(n6530), .B(n6531), .Z(n5219) );
  NOR U5585 ( .A(n6532), .B(n6530), .Z(n6531) );
  XOR U5586 ( .A(n6533), .B(n6534), .Z(n5222) );
  NOR U5587 ( .A(n6535), .B(n6533), .Z(n6534) );
  XOR U5588 ( .A(n6536), .B(n6537), .Z(n5225) );
  NOR U5589 ( .A(n6538), .B(n6536), .Z(n6537) );
  XOR U5590 ( .A(n6539), .B(n6540), .Z(n5228) );
  NOR U5591 ( .A(n6541), .B(n6539), .Z(n6540) );
  XOR U5592 ( .A(n6542), .B(n6543), .Z(n5231) );
  NOR U5593 ( .A(n6544), .B(n6542), .Z(n6543) );
  XOR U5594 ( .A(n6545), .B(n6546), .Z(n5234) );
  NOR U5595 ( .A(n6547), .B(n6545), .Z(n6546) );
  XOR U5596 ( .A(n6548), .B(n6549), .Z(n5237) );
  NOR U5597 ( .A(n6550), .B(n6548), .Z(n6549) );
  XOR U5598 ( .A(n6551), .B(n6552), .Z(n5240) );
  NOR U5599 ( .A(n6553), .B(n6551), .Z(n6552) );
  XOR U5600 ( .A(n6554), .B(n6555), .Z(n5243) );
  NOR U5601 ( .A(n6556), .B(n6554), .Z(n6555) );
  XOR U5602 ( .A(n6557), .B(n6558), .Z(n5246) );
  NOR U5603 ( .A(n6559), .B(n6557), .Z(n6558) );
  XOR U5604 ( .A(n6560), .B(n6561), .Z(n5249) );
  NOR U5605 ( .A(n6562), .B(n6560), .Z(n6561) );
  XOR U5606 ( .A(n6563), .B(n6564), .Z(n5252) );
  NOR U5607 ( .A(n6565), .B(n6563), .Z(n6564) );
  XOR U5608 ( .A(n6566), .B(n6567), .Z(n5255) );
  NOR U5609 ( .A(n6568), .B(n6566), .Z(n6567) );
  XOR U5610 ( .A(n6569), .B(n6570), .Z(n5258) );
  NOR U5611 ( .A(n6571), .B(n6569), .Z(n6570) );
  XOR U5612 ( .A(n6572), .B(n6573), .Z(n5261) );
  NOR U5613 ( .A(n6574), .B(n6572), .Z(n6573) );
  XOR U5614 ( .A(n6575), .B(n6576), .Z(n5264) );
  NOR U5615 ( .A(n6577), .B(n6575), .Z(n6576) );
  XOR U5616 ( .A(n6578), .B(n6579), .Z(n5267) );
  NOR U5617 ( .A(n6580), .B(n6578), .Z(n6579) );
  XOR U5618 ( .A(n6581), .B(n6582), .Z(n5270) );
  NOR U5619 ( .A(n6583), .B(n6581), .Z(n6582) );
  XOR U5620 ( .A(n6584), .B(n6585), .Z(n5273) );
  NOR U5621 ( .A(n6586), .B(n6584), .Z(n6585) );
  XOR U5622 ( .A(n6587), .B(n6588), .Z(n5276) );
  NOR U5623 ( .A(n6589), .B(n6587), .Z(n6588) );
  XOR U5624 ( .A(n6590), .B(n6591), .Z(n5279) );
  NOR U5625 ( .A(n6592), .B(n6590), .Z(n6591) );
  XOR U5626 ( .A(n6593), .B(n6594), .Z(n5282) );
  NOR U5627 ( .A(n6595), .B(n6593), .Z(n6594) );
  XOR U5628 ( .A(n6596), .B(n6597), .Z(n5285) );
  NOR U5629 ( .A(n6598), .B(n6596), .Z(n6597) );
  XOR U5630 ( .A(n6599), .B(n6600), .Z(n5288) );
  NOR U5631 ( .A(n6601), .B(n6599), .Z(n6600) );
  XOR U5632 ( .A(n6602), .B(n6603), .Z(n5291) );
  NOR U5633 ( .A(n6604), .B(n6602), .Z(n6603) );
  XOR U5634 ( .A(n6605), .B(n6606), .Z(n5294) );
  NOR U5635 ( .A(n6607), .B(n6605), .Z(n6606) );
  XOR U5636 ( .A(n6608), .B(n6609), .Z(n5297) );
  NOR U5637 ( .A(n6610), .B(n6608), .Z(n6609) );
  XOR U5638 ( .A(n6611), .B(n6612), .Z(n5300) );
  NOR U5639 ( .A(n6613), .B(n6611), .Z(n6612) );
  XOR U5640 ( .A(n6614), .B(n6615), .Z(n5303) );
  NOR U5641 ( .A(n6616), .B(n6614), .Z(n6615) );
  XOR U5642 ( .A(n6617), .B(n6618), .Z(n5306) );
  NOR U5643 ( .A(n6619), .B(n6617), .Z(n6618) );
  XOR U5644 ( .A(n6620), .B(n6621), .Z(n5309) );
  NOR U5645 ( .A(n6622), .B(n6620), .Z(n6621) );
  XOR U5646 ( .A(n6623), .B(n6624), .Z(n5312) );
  NOR U5647 ( .A(n6625), .B(n6623), .Z(n6624) );
  XOR U5648 ( .A(n6626), .B(n6627), .Z(n5315) );
  NOR U5649 ( .A(n6628), .B(n6626), .Z(n6627) );
  XOR U5650 ( .A(n6629), .B(n6630), .Z(n5318) );
  NOR U5651 ( .A(n6631), .B(n6629), .Z(n6630) );
  XOR U5652 ( .A(n6632), .B(n6633), .Z(n5321) );
  NOR U5653 ( .A(n6634), .B(n6632), .Z(n6633) );
  XOR U5654 ( .A(n6635), .B(n6636), .Z(n5324) );
  NOR U5655 ( .A(n6637), .B(n6635), .Z(n6636) );
  XOR U5656 ( .A(n6638), .B(n6639), .Z(n5327) );
  NOR U5657 ( .A(n6640), .B(n6638), .Z(n6639) );
  XOR U5658 ( .A(n6641), .B(n6642), .Z(n5330) );
  NOR U5659 ( .A(n6643), .B(n6641), .Z(n6642) );
  XOR U5660 ( .A(n6644), .B(n6645), .Z(n5333) );
  NOR U5661 ( .A(n6646), .B(n6644), .Z(n6645) );
  XOR U5662 ( .A(n6647), .B(n6648), .Z(n5336) );
  NOR U5663 ( .A(n6649), .B(n6647), .Z(n6648) );
  XOR U5664 ( .A(n6650), .B(n6651), .Z(n5339) );
  NOR U5665 ( .A(n6652), .B(n6650), .Z(n6651) );
  XOR U5666 ( .A(n6653), .B(n6654), .Z(n5342) );
  NOR U5667 ( .A(n6655), .B(n6653), .Z(n6654) );
  XOR U5668 ( .A(n6656), .B(n6657), .Z(n5345) );
  NOR U5669 ( .A(n6658), .B(n6656), .Z(n6657) );
  XOR U5670 ( .A(n6659), .B(n6660), .Z(n5348) );
  NOR U5671 ( .A(n6661), .B(n6659), .Z(n6660) );
  XOR U5672 ( .A(n6662), .B(n6663), .Z(n5351) );
  NOR U5673 ( .A(n6664), .B(n6662), .Z(n6663) );
  XOR U5674 ( .A(n6665), .B(n6666), .Z(n5354) );
  NOR U5675 ( .A(n6667), .B(n6665), .Z(n6666) );
  XOR U5676 ( .A(n6668), .B(n6669), .Z(n5357) );
  NOR U5677 ( .A(n6670), .B(n6668), .Z(n6669) );
  XOR U5678 ( .A(n6671), .B(n6672), .Z(n5360) );
  NOR U5679 ( .A(n6673), .B(n6671), .Z(n6672) );
  XOR U5680 ( .A(n6674), .B(n6675), .Z(n5363) );
  NOR U5681 ( .A(n6676), .B(n6674), .Z(n6675) );
  XOR U5682 ( .A(n6677), .B(n6678), .Z(n5366) );
  NOR U5683 ( .A(n6679), .B(n6677), .Z(n6678) );
  XOR U5684 ( .A(n6680), .B(n6681), .Z(n5369) );
  NOR U5685 ( .A(n6682), .B(n6680), .Z(n6681) );
  XOR U5686 ( .A(n6683), .B(n6684), .Z(n5372) );
  NOR U5687 ( .A(n6685), .B(n6683), .Z(n6684) );
  XOR U5688 ( .A(n6686), .B(n6687), .Z(n5375) );
  NOR U5689 ( .A(n6688), .B(n6686), .Z(n6687) );
  XOR U5690 ( .A(n6689), .B(n6690), .Z(n5378) );
  NOR U5691 ( .A(n6691), .B(n6689), .Z(n6690) );
  XOR U5692 ( .A(n6692), .B(n6693), .Z(n5381) );
  NOR U5693 ( .A(n6694), .B(n6692), .Z(n6693) );
  XOR U5694 ( .A(n6695), .B(n6696), .Z(n5384) );
  NOR U5695 ( .A(n6697), .B(n6695), .Z(n6696) );
  XOR U5696 ( .A(n6698), .B(n6699), .Z(n5387) );
  NOR U5697 ( .A(n6700), .B(n6698), .Z(n6699) );
  XOR U5698 ( .A(n6701), .B(n6702), .Z(n5390) );
  NOR U5699 ( .A(n6703), .B(n6701), .Z(n6702) );
  XOR U5700 ( .A(n6704), .B(n6705), .Z(n5393) );
  NOR U5701 ( .A(n6706), .B(n6704), .Z(n6705) );
  XOR U5702 ( .A(n6707), .B(n6708), .Z(n5396) );
  NOR U5703 ( .A(n6709), .B(n6707), .Z(n6708) );
  XOR U5704 ( .A(n6710), .B(n6711), .Z(n5399) );
  NOR U5705 ( .A(n6712), .B(n6710), .Z(n6711) );
  XOR U5706 ( .A(n6713), .B(n6714), .Z(n5402) );
  NOR U5707 ( .A(n6715), .B(n6713), .Z(n6714) );
  XOR U5708 ( .A(n6716), .B(n6717), .Z(n5405) );
  NOR U5709 ( .A(n6718), .B(n6716), .Z(n6717) );
  XOR U5710 ( .A(n6719), .B(n6720), .Z(n5408) );
  NOR U5711 ( .A(n6721), .B(n6719), .Z(n6720) );
  XOR U5712 ( .A(n6722), .B(n6723), .Z(n5411) );
  NOR U5713 ( .A(n6724), .B(n6722), .Z(n6723) );
  XOR U5714 ( .A(n6725), .B(n6726), .Z(n5414) );
  NOR U5715 ( .A(n6727), .B(n6725), .Z(n6726) );
  XOR U5716 ( .A(n6728), .B(n6729), .Z(n5417) );
  NOR U5717 ( .A(n101), .B(n6730), .Z(n6729) );
  XOR U5718 ( .A(n6731), .B(n6732), .Z(n5420) );
  AND U5719 ( .A(n6733), .B(n6734), .Z(n6732) );
  XOR U5720 ( .A(n6731), .B(n103), .Z(n6734) );
  XNOR U5721 ( .A(n6075), .B(n6074), .Z(n103) );
  XNOR U5722 ( .A(n6072), .B(n6071), .Z(n6074) );
  XNOR U5723 ( .A(n6069), .B(n6068), .Z(n6071) );
  XNOR U5724 ( .A(n6066), .B(n6065), .Z(n6068) );
  XNOR U5725 ( .A(n6063), .B(n6062), .Z(n6065) );
  XNOR U5726 ( .A(n6060), .B(n6059), .Z(n6062) );
  XNOR U5727 ( .A(n6057), .B(n6056), .Z(n6059) );
  XNOR U5728 ( .A(n6054), .B(n6053), .Z(n6056) );
  XNOR U5729 ( .A(n6051), .B(n6050), .Z(n6053) );
  XNOR U5730 ( .A(n6048), .B(n6047), .Z(n6050) );
  XNOR U5731 ( .A(n6045), .B(n6044), .Z(n6047) );
  XNOR U5732 ( .A(n6042), .B(n6041), .Z(n6044) );
  XNOR U5733 ( .A(n6039), .B(n6038), .Z(n6041) );
  XNOR U5734 ( .A(n6036), .B(n6035), .Z(n6038) );
  XNOR U5735 ( .A(n6033), .B(n6032), .Z(n6035) );
  XNOR U5736 ( .A(n6030), .B(n6029), .Z(n6032) );
  XNOR U5737 ( .A(n6027), .B(n6026), .Z(n6029) );
  XNOR U5738 ( .A(n6024), .B(n6023), .Z(n6026) );
  XNOR U5739 ( .A(n6021), .B(n6020), .Z(n6023) );
  XNOR U5740 ( .A(n6018), .B(n6017), .Z(n6020) );
  XNOR U5741 ( .A(n6015), .B(n6014), .Z(n6017) );
  XNOR U5742 ( .A(n6012), .B(n6011), .Z(n6014) );
  XNOR U5743 ( .A(n6009), .B(n6008), .Z(n6011) );
  XNOR U5744 ( .A(n6006), .B(n6005), .Z(n6008) );
  XNOR U5745 ( .A(n6003), .B(n6002), .Z(n6005) );
  XNOR U5746 ( .A(n6000), .B(n5999), .Z(n6002) );
  XNOR U5747 ( .A(n5997), .B(n5996), .Z(n5999) );
  XNOR U5748 ( .A(n5994), .B(n5993), .Z(n5996) );
  XNOR U5749 ( .A(n5991), .B(n5990), .Z(n5993) );
  XNOR U5750 ( .A(n5988), .B(n5987), .Z(n5990) );
  XNOR U5751 ( .A(n5985), .B(n5984), .Z(n5987) );
  XNOR U5752 ( .A(n5982), .B(n5981), .Z(n5984) );
  XNOR U5753 ( .A(n5979), .B(n5978), .Z(n5981) );
  XNOR U5754 ( .A(n5976), .B(n5975), .Z(n5978) );
  XNOR U5755 ( .A(n5973), .B(n5972), .Z(n5975) );
  XNOR U5756 ( .A(n5970), .B(n5969), .Z(n5972) );
  XNOR U5757 ( .A(n5967), .B(n5966), .Z(n5969) );
  XNOR U5758 ( .A(n5964), .B(n5963), .Z(n5966) );
  XNOR U5759 ( .A(n5961), .B(n5960), .Z(n5963) );
  XNOR U5760 ( .A(n5958), .B(n5957), .Z(n5960) );
  XNOR U5761 ( .A(n5955), .B(n5954), .Z(n5957) );
  XNOR U5762 ( .A(n5952), .B(n5951), .Z(n5954) );
  XNOR U5763 ( .A(n5949), .B(n5948), .Z(n5951) );
  XNOR U5764 ( .A(n5946), .B(n5945), .Z(n5948) );
  XNOR U5765 ( .A(n5943), .B(n5942), .Z(n5945) );
  XNOR U5766 ( .A(n5940), .B(n5939), .Z(n5942) );
  XNOR U5767 ( .A(n5937), .B(n5936), .Z(n5939) );
  XNOR U5768 ( .A(n5934), .B(n5933), .Z(n5936) );
  XNOR U5769 ( .A(n5931), .B(n5930), .Z(n5933) );
  XNOR U5770 ( .A(n5928), .B(n5927), .Z(n5930) );
  XNOR U5771 ( .A(n5925), .B(n5924), .Z(n5927) );
  XNOR U5772 ( .A(n5922), .B(n5921), .Z(n5924) );
  XNOR U5773 ( .A(n5919), .B(n5918), .Z(n5921) );
  XNOR U5774 ( .A(n5916), .B(n5915), .Z(n5918) );
  XNOR U5775 ( .A(n5913), .B(n5912), .Z(n5915) );
  XNOR U5776 ( .A(n5910), .B(n5909), .Z(n5912) );
  XNOR U5777 ( .A(n5907), .B(n5906), .Z(n5909) );
  XNOR U5778 ( .A(n5904), .B(n5903), .Z(n5906) );
  XNOR U5779 ( .A(n5901), .B(n5900), .Z(n5903) );
  XNOR U5780 ( .A(n5898), .B(n5897), .Z(n5900) );
  XNOR U5781 ( .A(n5895), .B(n5894), .Z(n5897) );
  XNOR U5782 ( .A(n5892), .B(n5891), .Z(n5894) );
  XNOR U5783 ( .A(n5889), .B(n5888), .Z(n5891) );
  XNOR U5784 ( .A(n5886), .B(n5885), .Z(n5888) );
  XNOR U5785 ( .A(n5883), .B(n5882), .Z(n5885) );
  XNOR U5786 ( .A(n5880), .B(n5879), .Z(n5882) );
  XNOR U5787 ( .A(n5877), .B(n5876), .Z(n5879) );
  XNOR U5788 ( .A(n5874), .B(n5873), .Z(n5876) );
  XNOR U5789 ( .A(n5871), .B(n5870), .Z(n5873) );
  XNOR U5790 ( .A(n5868), .B(n5867), .Z(n5870) );
  XNOR U5791 ( .A(n5865), .B(n5864), .Z(n5867) );
  XNOR U5792 ( .A(n5862), .B(n5861), .Z(n5864) );
  XNOR U5793 ( .A(n5859), .B(n5858), .Z(n5861) );
  XNOR U5794 ( .A(n5856), .B(n5855), .Z(n5858) );
  XNOR U5795 ( .A(n5853), .B(n5852), .Z(n5855) );
  XNOR U5796 ( .A(n5850), .B(n5849), .Z(n5852) );
  XNOR U5797 ( .A(n5847), .B(n5846), .Z(n5849) );
  XNOR U5798 ( .A(n5844), .B(n5843), .Z(n5846) );
  XNOR U5799 ( .A(n5841), .B(n5840), .Z(n5843) );
  XNOR U5800 ( .A(n5838), .B(n5837), .Z(n5840) );
  XNOR U5801 ( .A(n5835), .B(n5834), .Z(n5837) );
  XNOR U5802 ( .A(n5832), .B(n5831), .Z(n5834) );
  XNOR U5803 ( .A(n5829), .B(n5828), .Z(n5831) );
  XNOR U5804 ( .A(n5826), .B(n5825), .Z(n5828) );
  XNOR U5805 ( .A(n5823), .B(n5822), .Z(n5825) );
  XNOR U5806 ( .A(n5820), .B(n5819), .Z(n5822) );
  XNOR U5807 ( .A(n5817), .B(n5816), .Z(n5819) );
  XNOR U5808 ( .A(n5814), .B(n5813), .Z(n5816) );
  XNOR U5809 ( .A(n5811), .B(n5810), .Z(n5813) );
  XNOR U5810 ( .A(n5808), .B(n5807), .Z(n5810) );
  XNOR U5811 ( .A(n5805), .B(n5804), .Z(n5807) );
  XNOR U5812 ( .A(n5802), .B(n5801), .Z(n5804) );
  XNOR U5813 ( .A(n5799), .B(n5798), .Z(n5801) );
  XNOR U5814 ( .A(n5796), .B(n5795), .Z(n5798) );
  XNOR U5815 ( .A(n5793), .B(n5792), .Z(n5795) );
  XNOR U5816 ( .A(n5790), .B(n5789), .Z(n5792) );
  XNOR U5817 ( .A(n5787), .B(n5786), .Z(n5789) );
  XNOR U5818 ( .A(n5784), .B(n5783), .Z(n5786) );
  XNOR U5819 ( .A(n5781), .B(n5780), .Z(n5783) );
  XNOR U5820 ( .A(n5778), .B(n5777), .Z(n5780) );
  XNOR U5821 ( .A(n5775), .B(n5774), .Z(n5777) );
  XNOR U5822 ( .A(n5772), .B(n5771), .Z(n5774) );
  XNOR U5823 ( .A(n5769), .B(n5768), .Z(n5771) );
  XNOR U5824 ( .A(n5766), .B(n5765), .Z(n5768) );
  XNOR U5825 ( .A(n5763), .B(n5762), .Z(n5765) );
  XNOR U5826 ( .A(n5760), .B(n5759), .Z(n5762) );
  XNOR U5827 ( .A(n5757), .B(n5756), .Z(n5759) );
  XNOR U5828 ( .A(n5754), .B(n5753), .Z(n5756) );
  XNOR U5829 ( .A(n5751), .B(n5750), .Z(n5753) );
  XNOR U5830 ( .A(n5748), .B(n5747), .Z(n5750) );
  XNOR U5831 ( .A(n5745), .B(n5744), .Z(n5747) );
  XNOR U5832 ( .A(n5742), .B(n5741), .Z(n5744) );
  XNOR U5833 ( .A(n5739), .B(n5738), .Z(n5741) );
  XNOR U5834 ( .A(n5736), .B(n5735), .Z(n5738) );
  XNOR U5835 ( .A(n5733), .B(n5732), .Z(n5735) );
  XNOR U5836 ( .A(n5730), .B(n5729), .Z(n5732) );
  XNOR U5837 ( .A(n5727), .B(n5726), .Z(n5729) );
  XNOR U5838 ( .A(n5724), .B(n5723), .Z(n5726) );
  XNOR U5839 ( .A(n5721), .B(n5720), .Z(n5723) );
  XNOR U5840 ( .A(n5718), .B(n5717), .Z(n5720) );
  XNOR U5841 ( .A(n5715), .B(n5714), .Z(n5717) );
  XNOR U5842 ( .A(n5712), .B(n5711), .Z(n5714) );
  XNOR U5843 ( .A(n5709), .B(n5708), .Z(n5711) );
  XNOR U5844 ( .A(n5706), .B(n5705), .Z(n5708) );
  XNOR U5845 ( .A(n5703), .B(n5702), .Z(n5705) );
  XNOR U5846 ( .A(n5700), .B(n5699), .Z(n5702) );
  XNOR U5847 ( .A(n5697), .B(n5696), .Z(n5699) );
  XNOR U5848 ( .A(n5694), .B(n5693), .Z(n5696) );
  XNOR U5849 ( .A(n5691), .B(n5690), .Z(n5693) );
  XOR U5850 ( .A(n5688), .B(n5687), .Z(n5690) );
  XOR U5851 ( .A(n5685), .B(n5684), .Z(n5687) );
  XOR U5852 ( .A(n5681), .B(n5682), .Z(n5684) );
  AND U5853 ( .A(n6735), .B(n6736), .Z(n5682) );
  XOR U5854 ( .A(n5678), .B(n5679), .Z(n5681) );
  AND U5855 ( .A(n6737), .B(n6738), .Z(n5679) );
  XOR U5856 ( .A(n5675), .B(n5676), .Z(n5678) );
  AND U5857 ( .A(n6739), .B(n6740), .Z(n5676) );
  XNOR U5858 ( .A(n5424), .B(n5673), .Z(n5675) );
  AND U5859 ( .A(n6741), .B(n6742), .Z(n5673) );
  XOR U5860 ( .A(n5426), .B(n5425), .Z(n5424) );
  AND U5861 ( .A(n6743), .B(n6744), .Z(n5425) );
  XOR U5862 ( .A(n5428), .B(n5427), .Z(n5426) );
  AND U5863 ( .A(n6745), .B(n6746), .Z(n5427) );
  XOR U5864 ( .A(n5430), .B(n5429), .Z(n5428) );
  AND U5865 ( .A(n6747), .B(n6748), .Z(n5429) );
  XOR U5866 ( .A(n5432), .B(n5431), .Z(n5430) );
  AND U5867 ( .A(n6749), .B(n6750), .Z(n5431) );
  XOR U5868 ( .A(n5434), .B(n5433), .Z(n5432) );
  AND U5869 ( .A(n6751), .B(n6752), .Z(n5433) );
  XOR U5870 ( .A(n5436), .B(n5435), .Z(n5434) );
  AND U5871 ( .A(n6753), .B(n6754), .Z(n5435) );
  XOR U5872 ( .A(n5438), .B(n5437), .Z(n5436) );
  AND U5873 ( .A(n6755), .B(n6756), .Z(n5437) );
  XOR U5874 ( .A(n5440), .B(n5439), .Z(n5438) );
  AND U5875 ( .A(n6757), .B(n6758), .Z(n5439) );
  XOR U5876 ( .A(n5442), .B(n5441), .Z(n5440) );
  AND U5877 ( .A(n6759), .B(n6760), .Z(n5441) );
  XOR U5878 ( .A(n5444), .B(n5443), .Z(n5442) );
  AND U5879 ( .A(n6761), .B(n6762), .Z(n5443) );
  XOR U5880 ( .A(n5446), .B(n5445), .Z(n5444) );
  AND U5881 ( .A(n6763), .B(n6764), .Z(n5445) );
  XOR U5882 ( .A(n5448), .B(n5447), .Z(n5446) );
  AND U5883 ( .A(n6765), .B(n6766), .Z(n5447) );
  XOR U5884 ( .A(n5450), .B(n5449), .Z(n5448) );
  AND U5885 ( .A(n6767), .B(n6768), .Z(n5449) );
  XOR U5886 ( .A(n5452), .B(n5451), .Z(n5450) );
  AND U5887 ( .A(n6769), .B(n6770), .Z(n5451) );
  XOR U5888 ( .A(n5454), .B(n5453), .Z(n5452) );
  AND U5889 ( .A(n6771), .B(n6772), .Z(n5453) );
  XOR U5890 ( .A(n5456), .B(n5455), .Z(n5454) );
  AND U5891 ( .A(n6773), .B(n6774), .Z(n5455) );
  XOR U5892 ( .A(n5458), .B(n5457), .Z(n5456) );
  AND U5893 ( .A(n6775), .B(n6776), .Z(n5457) );
  XOR U5894 ( .A(n5460), .B(n5459), .Z(n5458) );
  AND U5895 ( .A(n6777), .B(n6778), .Z(n5459) );
  XOR U5896 ( .A(n5462), .B(n5461), .Z(n5460) );
  AND U5897 ( .A(n6779), .B(n6780), .Z(n5461) );
  XOR U5898 ( .A(n5464), .B(n5463), .Z(n5462) );
  AND U5899 ( .A(n6781), .B(n6782), .Z(n5463) );
  XOR U5900 ( .A(n5466), .B(n5465), .Z(n5464) );
  AND U5901 ( .A(n6783), .B(n6784), .Z(n5465) );
  XOR U5902 ( .A(n5468), .B(n5467), .Z(n5466) );
  AND U5903 ( .A(n6785), .B(n6786), .Z(n5467) );
  XOR U5904 ( .A(n5470), .B(n5469), .Z(n5468) );
  AND U5905 ( .A(n6787), .B(n6788), .Z(n5469) );
  XOR U5906 ( .A(n5472), .B(n5471), .Z(n5470) );
  AND U5907 ( .A(n6789), .B(n6790), .Z(n5471) );
  XOR U5908 ( .A(n5474), .B(n5473), .Z(n5472) );
  AND U5909 ( .A(n6791), .B(n6792), .Z(n5473) );
  XOR U5910 ( .A(n5476), .B(n5475), .Z(n5474) );
  AND U5911 ( .A(n6793), .B(n6794), .Z(n5475) );
  XOR U5912 ( .A(n5478), .B(n5477), .Z(n5476) );
  AND U5913 ( .A(n6795), .B(n6796), .Z(n5477) );
  XOR U5914 ( .A(n5480), .B(n5479), .Z(n5478) );
  AND U5915 ( .A(n6797), .B(n6798), .Z(n5479) );
  XOR U5916 ( .A(n5482), .B(n5481), .Z(n5480) );
  AND U5917 ( .A(n6799), .B(n6800), .Z(n5481) );
  XOR U5918 ( .A(n5484), .B(n5483), .Z(n5482) );
  AND U5919 ( .A(n6801), .B(n6802), .Z(n5483) );
  XOR U5920 ( .A(n5486), .B(n5485), .Z(n5484) );
  AND U5921 ( .A(n6803), .B(n6804), .Z(n5485) );
  XOR U5922 ( .A(n5488), .B(n5487), .Z(n5486) );
  AND U5923 ( .A(n6805), .B(n6806), .Z(n5487) );
  XOR U5924 ( .A(n5490), .B(n5489), .Z(n5488) );
  AND U5925 ( .A(n6807), .B(n6808), .Z(n5489) );
  XOR U5926 ( .A(n5492), .B(n5491), .Z(n5490) );
  AND U5927 ( .A(n6809), .B(n6810), .Z(n5491) );
  XOR U5928 ( .A(n5494), .B(n5493), .Z(n5492) );
  AND U5929 ( .A(n6811), .B(n6812), .Z(n5493) );
  XOR U5930 ( .A(n5496), .B(n5495), .Z(n5494) );
  AND U5931 ( .A(n6813), .B(n6814), .Z(n5495) );
  XOR U5932 ( .A(n5498), .B(n5497), .Z(n5496) );
  AND U5933 ( .A(n6815), .B(n6816), .Z(n5497) );
  XOR U5934 ( .A(n5500), .B(n5499), .Z(n5498) );
  AND U5935 ( .A(n6817), .B(n6818), .Z(n5499) );
  XOR U5936 ( .A(n5502), .B(n5501), .Z(n5500) );
  AND U5937 ( .A(n6819), .B(n6820), .Z(n5501) );
  XOR U5938 ( .A(n5504), .B(n5503), .Z(n5502) );
  AND U5939 ( .A(n6821), .B(n6822), .Z(n5503) );
  XOR U5940 ( .A(n5506), .B(n5505), .Z(n5504) );
  AND U5941 ( .A(n6823), .B(n6824), .Z(n5505) );
  XOR U5942 ( .A(n5508), .B(n5507), .Z(n5506) );
  AND U5943 ( .A(n6825), .B(n6826), .Z(n5507) );
  XOR U5944 ( .A(n5510), .B(n5509), .Z(n5508) );
  AND U5945 ( .A(n6827), .B(n6828), .Z(n5509) );
  XOR U5946 ( .A(n5512), .B(n5511), .Z(n5510) );
  AND U5947 ( .A(n6829), .B(n6830), .Z(n5511) );
  XOR U5948 ( .A(n5514), .B(n5513), .Z(n5512) );
  AND U5949 ( .A(n6831), .B(n6832), .Z(n5513) );
  XOR U5950 ( .A(n5516), .B(n5515), .Z(n5514) );
  AND U5951 ( .A(n6833), .B(n6834), .Z(n5515) );
  XOR U5952 ( .A(n5518), .B(n5517), .Z(n5516) );
  AND U5953 ( .A(n6835), .B(n6836), .Z(n5517) );
  XOR U5954 ( .A(n5520), .B(n5519), .Z(n5518) );
  AND U5955 ( .A(n6837), .B(n6838), .Z(n5519) );
  XOR U5956 ( .A(n5522), .B(n5521), .Z(n5520) );
  AND U5957 ( .A(n6839), .B(n6840), .Z(n5521) );
  XOR U5958 ( .A(n5524), .B(n5523), .Z(n5522) );
  AND U5959 ( .A(n6841), .B(n6842), .Z(n5523) );
  XOR U5960 ( .A(n5526), .B(n5525), .Z(n5524) );
  AND U5961 ( .A(n6843), .B(n6844), .Z(n5525) );
  XOR U5962 ( .A(n5528), .B(n5527), .Z(n5526) );
  AND U5963 ( .A(n6845), .B(n6846), .Z(n5527) );
  XOR U5964 ( .A(n5530), .B(n5529), .Z(n5528) );
  AND U5965 ( .A(n6847), .B(n6848), .Z(n5529) );
  XOR U5966 ( .A(n5532), .B(n5531), .Z(n5530) );
  AND U5967 ( .A(n6849), .B(n6850), .Z(n5531) );
  XOR U5968 ( .A(n5534), .B(n5533), .Z(n5532) );
  AND U5969 ( .A(n6851), .B(n6852), .Z(n5533) );
  XOR U5970 ( .A(n5536), .B(n5535), .Z(n5534) );
  AND U5971 ( .A(n6853), .B(n6854), .Z(n5535) );
  XOR U5972 ( .A(n5538), .B(n5537), .Z(n5536) );
  AND U5973 ( .A(n6855), .B(n6856), .Z(n5537) );
  XOR U5974 ( .A(n5540), .B(n5539), .Z(n5538) );
  AND U5975 ( .A(n6857), .B(n6858), .Z(n5539) );
  XOR U5976 ( .A(n5542), .B(n5541), .Z(n5540) );
  AND U5977 ( .A(n6859), .B(n6860), .Z(n5541) );
  XOR U5978 ( .A(n5544), .B(n5543), .Z(n5542) );
  AND U5979 ( .A(n6861), .B(n6862), .Z(n5543) );
  XOR U5980 ( .A(n5546), .B(n5545), .Z(n5544) );
  AND U5981 ( .A(n6863), .B(n6864), .Z(n5545) );
  XOR U5982 ( .A(n5548), .B(n5547), .Z(n5546) );
  AND U5983 ( .A(n6865), .B(n6866), .Z(n5547) );
  XOR U5984 ( .A(n5550), .B(n5549), .Z(n5548) );
  AND U5985 ( .A(n6867), .B(n6868), .Z(n5549) );
  XOR U5986 ( .A(n5552), .B(n5551), .Z(n5550) );
  AND U5987 ( .A(n6869), .B(n6870), .Z(n5551) );
  XOR U5988 ( .A(n5554), .B(n5553), .Z(n5552) );
  AND U5989 ( .A(n6871), .B(n6872), .Z(n5553) );
  XOR U5990 ( .A(n5556), .B(n5555), .Z(n5554) );
  AND U5991 ( .A(n6873), .B(n6874), .Z(n5555) );
  XOR U5992 ( .A(n5558), .B(n5557), .Z(n5556) );
  AND U5993 ( .A(n6875), .B(n6876), .Z(n5557) );
  XOR U5994 ( .A(n5560), .B(n5559), .Z(n5558) );
  AND U5995 ( .A(n6877), .B(n6878), .Z(n5559) );
  XOR U5996 ( .A(n5562), .B(n5561), .Z(n5560) );
  AND U5997 ( .A(n6879), .B(n6880), .Z(n5561) );
  XOR U5998 ( .A(n5564), .B(n5563), .Z(n5562) );
  AND U5999 ( .A(n6881), .B(n6882), .Z(n5563) );
  XOR U6000 ( .A(n5566), .B(n5565), .Z(n5564) );
  AND U6001 ( .A(n6883), .B(n6884), .Z(n5565) );
  XOR U6002 ( .A(n5568), .B(n5567), .Z(n5566) );
  AND U6003 ( .A(n6885), .B(n6886), .Z(n5567) );
  XOR U6004 ( .A(n5570), .B(n5569), .Z(n5568) );
  AND U6005 ( .A(n6887), .B(n6888), .Z(n5569) );
  XOR U6006 ( .A(n5572), .B(n5571), .Z(n5570) );
  AND U6007 ( .A(n6889), .B(n6890), .Z(n5571) );
  XOR U6008 ( .A(n5574), .B(n5573), .Z(n5572) );
  AND U6009 ( .A(n6891), .B(n6892), .Z(n5573) );
  XOR U6010 ( .A(n5576), .B(n5575), .Z(n5574) );
  AND U6011 ( .A(n6893), .B(n6894), .Z(n5575) );
  XOR U6012 ( .A(n5578), .B(n5577), .Z(n5576) );
  AND U6013 ( .A(n6895), .B(n6896), .Z(n5577) );
  XOR U6014 ( .A(n5580), .B(n5579), .Z(n5578) );
  AND U6015 ( .A(n6897), .B(n6898), .Z(n5579) );
  XOR U6016 ( .A(n5582), .B(n5581), .Z(n5580) );
  AND U6017 ( .A(n6899), .B(n6900), .Z(n5581) );
  XOR U6018 ( .A(n5584), .B(n5583), .Z(n5582) );
  AND U6019 ( .A(n6901), .B(n6902), .Z(n5583) );
  XOR U6020 ( .A(n5586), .B(n5585), .Z(n5584) );
  AND U6021 ( .A(n6903), .B(n6904), .Z(n5585) );
  XOR U6022 ( .A(n5588), .B(n5587), .Z(n5586) );
  AND U6023 ( .A(n6905), .B(n6906), .Z(n5587) );
  XOR U6024 ( .A(n5590), .B(n5589), .Z(n5588) );
  AND U6025 ( .A(n6907), .B(n6908), .Z(n5589) );
  XOR U6026 ( .A(n5592), .B(n5591), .Z(n5590) );
  AND U6027 ( .A(n6909), .B(n6910), .Z(n5591) );
  XOR U6028 ( .A(n5594), .B(n5593), .Z(n5592) );
  AND U6029 ( .A(n6911), .B(n6912), .Z(n5593) );
  XOR U6030 ( .A(n5596), .B(n5595), .Z(n5594) );
  AND U6031 ( .A(n6913), .B(n6914), .Z(n5595) );
  XOR U6032 ( .A(n5598), .B(n5597), .Z(n5596) );
  AND U6033 ( .A(n6915), .B(n6916), .Z(n5597) );
  XOR U6034 ( .A(n5600), .B(n5599), .Z(n5598) );
  AND U6035 ( .A(n6917), .B(n6918), .Z(n5599) );
  XOR U6036 ( .A(n5602), .B(n5601), .Z(n5600) );
  AND U6037 ( .A(n6919), .B(n6920), .Z(n5601) );
  XOR U6038 ( .A(n5604), .B(n5603), .Z(n5602) );
  AND U6039 ( .A(n6921), .B(n6922), .Z(n5603) );
  XOR U6040 ( .A(n5606), .B(n5605), .Z(n5604) );
  AND U6041 ( .A(n6923), .B(n6924), .Z(n5605) );
  XOR U6042 ( .A(n5608), .B(n5607), .Z(n5606) );
  AND U6043 ( .A(n6925), .B(n6926), .Z(n5607) );
  XOR U6044 ( .A(n5610), .B(n5609), .Z(n5608) );
  AND U6045 ( .A(n6927), .B(n6928), .Z(n5609) );
  XOR U6046 ( .A(n5612), .B(n5611), .Z(n5610) );
  AND U6047 ( .A(n6929), .B(n6930), .Z(n5611) );
  XOR U6048 ( .A(n5614), .B(n5613), .Z(n5612) );
  AND U6049 ( .A(n6931), .B(n6932), .Z(n5613) );
  XOR U6050 ( .A(n5616), .B(n5615), .Z(n5614) );
  AND U6051 ( .A(n6933), .B(n6934), .Z(n5615) );
  XOR U6052 ( .A(n5669), .B(n5617), .Z(n5616) );
  AND U6053 ( .A(n6935), .B(n6936), .Z(n5617) );
  XOR U6054 ( .A(n5671), .B(n5670), .Z(n5669) );
  AND U6055 ( .A(n6937), .B(n6938), .Z(n5670) );
  XOR U6056 ( .A(n5652), .B(n5672), .Z(n5671) );
  AND U6057 ( .A(n6939), .B(n6940), .Z(n5672) );
  XOR U6058 ( .A(n5654), .B(n5653), .Z(n5652) );
  AND U6059 ( .A(n6941), .B(n6942), .Z(n5653) );
  XOR U6060 ( .A(n5656), .B(n5655), .Z(n5654) );
  AND U6061 ( .A(n6943), .B(n6944), .Z(n5655) );
  XOR U6062 ( .A(n5660), .B(n5657), .Z(n5656) );
  AND U6063 ( .A(n6945), .B(n6946), .Z(n5657) );
  XOR U6064 ( .A(n5662), .B(n5661), .Z(n5660) );
  AND U6065 ( .A(n6947), .B(n6948), .Z(n5661) );
  XOR U6066 ( .A(n5665), .B(n5663), .Z(n5662) );
  AND U6067 ( .A(n6949), .B(n6950), .Z(n5663) );
  XOR U6068 ( .A(n5667), .B(n5666), .Z(n5665) );
  AND U6069 ( .A(n6951), .B(n6952), .Z(n5666) );
  XOR U6070 ( .A(n5632), .B(n5668), .Z(n5667) );
  AND U6071 ( .A(n6953), .B(n6954), .Z(n5668) );
  XNOR U6072 ( .A(n5639), .B(n5633), .Z(n5632) );
  AND U6073 ( .A(n6955), .B(n6956), .Z(n5633) );
  XOR U6074 ( .A(n5638), .B(n5630), .Z(n5639) );
  AND U6075 ( .A(n6957), .B(n6958), .Z(n5630) );
  XOR U6076 ( .A(n5651), .B(n5629), .Z(n5638) );
  AND U6077 ( .A(n6959), .B(n6960), .Z(n5629) );
  XNOR U6078 ( .A(n6961), .B(n6962), .Z(n5651) );
  XOR U6079 ( .A(n5649), .B(n6963), .Z(n6962) );
  XOR U6080 ( .A(n5647), .B(n5645), .Z(n6963) );
  AND U6081 ( .A(n6964), .B(n6965), .Z(n5645) );
  AND U6082 ( .A(n6966), .B(n6967), .Z(n5647) );
  AND U6083 ( .A(n6968), .B(n6969), .Z(n5649) );
  XNOR U6084 ( .A(n6970), .B(n5648), .Z(n6961) );
  XOR U6085 ( .A(n6971), .B(n6972), .Z(n5648) );
  XOR U6086 ( .A(n6973), .B(n6974), .Z(n6972) );
  AND U6087 ( .A(n6975), .B(n6976), .Z(n6974) );
  XNOR U6088 ( .A(n6977), .B(n6978), .Z(n6971) );
  NOR U6089 ( .A(n6979), .B(n6980), .Z(n6978) );
  AND U6090 ( .A(n6981), .B(n6982), .Z(n6980) );
  IV U6091 ( .A(n6983), .Z(n6979) );
  NOR U6092 ( .A(n6973), .B(n6984), .Z(n6983) );
  AND U6093 ( .A(n6985), .B(n6986), .Z(n6984) );
  NOR U6094 ( .A(n6975), .B(n6985), .Z(n6977) );
  XNOR U6095 ( .A(n5650), .B(n5628), .Z(n6970) );
  AND U6096 ( .A(n6987), .B(n6988), .Z(n5628) );
  AND U6097 ( .A(n6989), .B(n6990), .Z(n5650) );
  XOR U6098 ( .A(n6991), .B(n6992), .Z(n5685) );
  NOR U6099 ( .A(n6993), .B(n6994), .Z(n6992) );
  IV U6100 ( .A(n6991), .Z(n6993) );
  XOR U6101 ( .A(n6995), .B(n6996), .Z(n5688) );
  NOR U6102 ( .A(n6995), .B(n6997), .Z(n6996) );
  XNOR U6103 ( .A(n6998), .B(n6999), .Z(n5691) );
  AND U6104 ( .A(n6998), .B(n7000), .Z(n6999) );
  XNOR U6105 ( .A(n7001), .B(n7002), .Z(n5694) );
  AND U6106 ( .A(n7001), .B(n7003), .Z(n7002) );
  XNOR U6107 ( .A(n7004), .B(n7005), .Z(n5697) );
  AND U6108 ( .A(n7004), .B(n7006), .Z(n7005) );
  XNOR U6109 ( .A(n7007), .B(n7008), .Z(n5700) );
  AND U6110 ( .A(n7007), .B(n7009), .Z(n7008) );
  XNOR U6111 ( .A(n7010), .B(n7011), .Z(n5703) );
  AND U6112 ( .A(n7010), .B(n7012), .Z(n7011) );
  XNOR U6113 ( .A(n7013), .B(n7014), .Z(n5706) );
  AND U6114 ( .A(n7013), .B(n7015), .Z(n7014) );
  XNOR U6115 ( .A(n7016), .B(n7017), .Z(n5709) );
  AND U6116 ( .A(n7016), .B(n7018), .Z(n7017) );
  XNOR U6117 ( .A(n7019), .B(n7020), .Z(n5712) );
  AND U6118 ( .A(n7019), .B(n7021), .Z(n7020) );
  XNOR U6119 ( .A(n7022), .B(n7023), .Z(n5715) );
  AND U6120 ( .A(n7022), .B(n7024), .Z(n7023) );
  XNOR U6121 ( .A(n7025), .B(n7026), .Z(n5718) );
  AND U6122 ( .A(n7025), .B(n7027), .Z(n7026) );
  XNOR U6123 ( .A(n7028), .B(n7029), .Z(n5721) );
  AND U6124 ( .A(n7028), .B(n7030), .Z(n7029) );
  XNOR U6125 ( .A(n7031), .B(n7032), .Z(n5724) );
  AND U6126 ( .A(n7031), .B(n7033), .Z(n7032) );
  XNOR U6127 ( .A(n7034), .B(n7035), .Z(n5727) );
  AND U6128 ( .A(n7034), .B(n7036), .Z(n7035) );
  XNOR U6129 ( .A(n7037), .B(n7038), .Z(n5730) );
  AND U6130 ( .A(n7037), .B(n7039), .Z(n7038) );
  XNOR U6131 ( .A(n7040), .B(n7041), .Z(n5733) );
  AND U6132 ( .A(n7040), .B(n7042), .Z(n7041) );
  XNOR U6133 ( .A(n7043), .B(n7044), .Z(n5736) );
  AND U6134 ( .A(n7043), .B(n7045), .Z(n7044) );
  XNOR U6135 ( .A(n7046), .B(n7047), .Z(n5739) );
  AND U6136 ( .A(n7046), .B(n7048), .Z(n7047) );
  XNOR U6137 ( .A(n7049), .B(n7050), .Z(n5742) );
  AND U6138 ( .A(n7049), .B(n7051), .Z(n7050) );
  XNOR U6139 ( .A(n7052), .B(n7053), .Z(n5745) );
  AND U6140 ( .A(n7052), .B(n7054), .Z(n7053) );
  XNOR U6141 ( .A(n7055), .B(n7056), .Z(n5748) );
  AND U6142 ( .A(n7055), .B(n7057), .Z(n7056) );
  XNOR U6143 ( .A(n7058), .B(n7059), .Z(n5751) );
  AND U6144 ( .A(n7058), .B(n7060), .Z(n7059) );
  XNOR U6145 ( .A(n7061), .B(n7062), .Z(n5754) );
  AND U6146 ( .A(n7061), .B(n7063), .Z(n7062) );
  XNOR U6147 ( .A(n7064), .B(n7065), .Z(n5757) );
  AND U6148 ( .A(n7064), .B(n7066), .Z(n7065) );
  XNOR U6149 ( .A(n7067), .B(n7068), .Z(n5760) );
  AND U6150 ( .A(n7067), .B(n7069), .Z(n7068) );
  XNOR U6151 ( .A(n7070), .B(n7071), .Z(n5763) );
  AND U6152 ( .A(n7070), .B(n7072), .Z(n7071) );
  XNOR U6153 ( .A(n7073), .B(n7074), .Z(n5766) );
  AND U6154 ( .A(n7073), .B(n7075), .Z(n7074) );
  XNOR U6155 ( .A(n7076), .B(n7077), .Z(n5769) );
  AND U6156 ( .A(n7076), .B(n7078), .Z(n7077) );
  XNOR U6157 ( .A(n7079), .B(n7080), .Z(n5772) );
  AND U6158 ( .A(n7079), .B(n7081), .Z(n7080) );
  XNOR U6159 ( .A(n7082), .B(n7083), .Z(n5775) );
  AND U6160 ( .A(n7082), .B(n7084), .Z(n7083) );
  XNOR U6161 ( .A(n7085), .B(n7086), .Z(n5778) );
  AND U6162 ( .A(n7085), .B(n7087), .Z(n7086) );
  XNOR U6163 ( .A(n7088), .B(n7089), .Z(n5781) );
  AND U6164 ( .A(n7088), .B(n7090), .Z(n7089) );
  XNOR U6165 ( .A(n7091), .B(n7092), .Z(n5784) );
  AND U6166 ( .A(n7091), .B(n7093), .Z(n7092) );
  XNOR U6167 ( .A(n7094), .B(n7095), .Z(n5787) );
  AND U6168 ( .A(n7094), .B(n7096), .Z(n7095) );
  XNOR U6169 ( .A(n7097), .B(n7098), .Z(n5790) );
  AND U6170 ( .A(n7097), .B(n7099), .Z(n7098) );
  XNOR U6171 ( .A(n7100), .B(n7101), .Z(n5793) );
  AND U6172 ( .A(n7100), .B(n7102), .Z(n7101) );
  XNOR U6173 ( .A(n7103), .B(n7104), .Z(n5796) );
  AND U6174 ( .A(n7103), .B(n7105), .Z(n7104) );
  XNOR U6175 ( .A(n7106), .B(n7107), .Z(n5799) );
  AND U6176 ( .A(n7106), .B(n7108), .Z(n7107) );
  XNOR U6177 ( .A(n7109), .B(n7110), .Z(n5802) );
  AND U6178 ( .A(n7109), .B(n7111), .Z(n7110) );
  XNOR U6179 ( .A(n7112), .B(n7113), .Z(n5805) );
  AND U6180 ( .A(n7112), .B(n7114), .Z(n7113) );
  XNOR U6181 ( .A(n7115), .B(n7116), .Z(n5808) );
  AND U6182 ( .A(n7115), .B(n7117), .Z(n7116) );
  XNOR U6183 ( .A(n7118), .B(n7119), .Z(n5811) );
  AND U6184 ( .A(n7118), .B(n7120), .Z(n7119) );
  XNOR U6185 ( .A(n7121), .B(n7122), .Z(n5814) );
  AND U6186 ( .A(n7121), .B(n7123), .Z(n7122) );
  XNOR U6187 ( .A(n7124), .B(n7125), .Z(n5817) );
  AND U6188 ( .A(n7124), .B(n7126), .Z(n7125) );
  XNOR U6189 ( .A(n7127), .B(n7128), .Z(n5820) );
  AND U6190 ( .A(n7127), .B(n7129), .Z(n7128) );
  XNOR U6191 ( .A(n7130), .B(n7131), .Z(n5823) );
  AND U6192 ( .A(n7130), .B(n7132), .Z(n7131) );
  XNOR U6193 ( .A(n7133), .B(n7134), .Z(n5826) );
  AND U6194 ( .A(n7133), .B(n7135), .Z(n7134) );
  XNOR U6195 ( .A(n7136), .B(n7137), .Z(n5829) );
  AND U6196 ( .A(n7136), .B(n7138), .Z(n7137) );
  XNOR U6197 ( .A(n7139), .B(n7140), .Z(n5832) );
  AND U6198 ( .A(n7139), .B(n7141), .Z(n7140) );
  XNOR U6199 ( .A(n7142), .B(n7143), .Z(n5835) );
  AND U6200 ( .A(n7142), .B(n7144), .Z(n7143) );
  XNOR U6201 ( .A(n7145), .B(n7146), .Z(n5838) );
  AND U6202 ( .A(n7145), .B(n7147), .Z(n7146) );
  XNOR U6203 ( .A(n7148), .B(n7149), .Z(n5841) );
  AND U6204 ( .A(n7148), .B(n7150), .Z(n7149) );
  XNOR U6205 ( .A(n7151), .B(n7152), .Z(n5844) );
  AND U6206 ( .A(n7151), .B(n7153), .Z(n7152) );
  XNOR U6207 ( .A(n7154), .B(n7155), .Z(n5847) );
  AND U6208 ( .A(n7154), .B(n7156), .Z(n7155) );
  XNOR U6209 ( .A(n7157), .B(n7158), .Z(n5850) );
  AND U6210 ( .A(n7157), .B(n7159), .Z(n7158) );
  XNOR U6211 ( .A(n7160), .B(n7161), .Z(n5853) );
  AND U6212 ( .A(n7160), .B(n7162), .Z(n7161) );
  XNOR U6213 ( .A(n7163), .B(n7164), .Z(n5856) );
  AND U6214 ( .A(n7163), .B(n7165), .Z(n7164) );
  XNOR U6215 ( .A(n7166), .B(n7167), .Z(n5859) );
  AND U6216 ( .A(n7166), .B(n7168), .Z(n7167) );
  XNOR U6217 ( .A(n7169), .B(n7170), .Z(n5862) );
  AND U6218 ( .A(n7169), .B(n7171), .Z(n7170) );
  XNOR U6219 ( .A(n7172), .B(n7173), .Z(n5865) );
  AND U6220 ( .A(n7172), .B(n7174), .Z(n7173) );
  XNOR U6221 ( .A(n7175), .B(n7176), .Z(n5868) );
  AND U6222 ( .A(n7175), .B(n7177), .Z(n7176) );
  XNOR U6223 ( .A(n7178), .B(n7179), .Z(n5871) );
  AND U6224 ( .A(n7178), .B(n7180), .Z(n7179) );
  XNOR U6225 ( .A(n7181), .B(n7182), .Z(n5874) );
  AND U6226 ( .A(n7181), .B(n7183), .Z(n7182) );
  XNOR U6227 ( .A(n7184), .B(n7185), .Z(n5877) );
  AND U6228 ( .A(n7184), .B(n7186), .Z(n7185) );
  XNOR U6229 ( .A(n7187), .B(n7188), .Z(n5880) );
  AND U6230 ( .A(n7187), .B(n7189), .Z(n7188) );
  XNOR U6231 ( .A(n7190), .B(n7191), .Z(n5883) );
  AND U6232 ( .A(n7190), .B(n7192), .Z(n7191) );
  XNOR U6233 ( .A(n7193), .B(n7194), .Z(n5886) );
  AND U6234 ( .A(n7193), .B(n7195), .Z(n7194) );
  XNOR U6235 ( .A(n7196), .B(n7197), .Z(n5889) );
  AND U6236 ( .A(n7196), .B(n7198), .Z(n7197) );
  XNOR U6237 ( .A(n7199), .B(n7200), .Z(n5892) );
  AND U6238 ( .A(n7199), .B(n7201), .Z(n7200) );
  XNOR U6239 ( .A(n7202), .B(n7203), .Z(n5895) );
  AND U6240 ( .A(n7202), .B(n7204), .Z(n7203) );
  XNOR U6241 ( .A(n7205), .B(n7206), .Z(n5898) );
  AND U6242 ( .A(n7205), .B(n7207), .Z(n7206) );
  XNOR U6243 ( .A(n7208), .B(n7209), .Z(n5901) );
  AND U6244 ( .A(n7208), .B(n7210), .Z(n7209) );
  XNOR U6245 ( .A(n7211), .B(n7212), .Z(n5904) );
  AND U6246 ( .A(n7211), .B(n7213), .Z(n7212) );
  XNOR U6247 ( .A(n7214), .B(n7215), .Z(n5907) );
  AND U6248 ( .A(n7214), .B(n7216), .Z(n7215) );
  XNOR U6249 ( .A(n7217), .B(n7218), .Z(n5910) );
  AND U6250 ( .A(n7217), .B(n7219), .Z(n7218) );
  XNOR U6251 ( .A(n7220), .B(n7221), .Z(n5913) );
  AND U6252 ( .A(n7220), .B(n7222), .Z(n7221) );
  XNOR U6253 ( .A(n7223), .B(n7224), .Z(n5916) );
  AND U6254 ( .A(n7223), .B(n7225), .Z(n7224) );
  XNOR U6255 ( .A(n7226), .B(n7227), .Z(n5919) );
  AND U6256 ( .A(n7226), .B(n7228), .Z(n7227) );
  XNOR U6257 ( .A(n7229), .B(n7230), .Z(n5922) );
  AND U6258 ( .A(n7229), .B(n7231), .Z(n7230) );
  XNOR U6259 ( .A(n7232), .B(n7233), .Z(n5925) );
  AND U6260 ( .A(n7232), .B(n7234), .Z(n7233) );
  XNOR U6261 ( .A(n7235), .B(n7236), .Z(n5928) );
  AND U6262 ( .A(n7235), .B(n7237), .Z(n7236) );
  XNOR U6263 ( .A(n7238), .B(n7239), .Z(n5931) );
  AND U6264 ( .A(n7238), .B(n7240), .Z(n7239) );
  XNOR U6265 ( .A(n7241), .B(n7242), .Z(n5934) );
  AND U6266 ( .A(n7241), .B(n7243), .Z(n7242) );
  XNOR U6267 ( .A(n7244), .B(n7245), .Z(n5937) );
  AND U6268 ( .A(n7244), .B(n7246), .Z(n7245) );
  XNOR U6269 ( .A(n7247), .B(n7248), .Z(n5940) );
  AND U6270 ( .A(n7247), .B(n7249), .Z(n7248) );
  XNOR U6271 ( .A(n7250), .B(n7251), .Z(n5943) );
  AND U6272 ( .A(n7250), .B(n7252), .Z(n7251) );
  XNOR U6273 ( .A(n7253), .B(n7254), .Z(n5946) );
  AND U6274 ( .A(n7253), .B(n7255), .Z(n7254) );
  XNOR U6275 ( .A(n7256), .B(n7257), .Z(n5949) );
  AND U6276 ( .A(n7256), .B(n7258), .Z(n7257) );
  XNOR U6277 ( .A(n7259), .B(n7260), .Z(n5952) );
  AND U6278 ( .A(n7259), .B(n7261), .Z(n7260) );
  XNOR U6279 ( .A(n7262), .B(n7263), .Z(n5955) );
  AND U6280 ( .A(n7262), .B(n7264), .Z(n7263) );
  XNOR U6281 ( .A(n7265), .B(n7266), .Z(n5958) );
  AND U6282 ( .A(n7265), .B(n7267), .Z(n7266) );
  XNOR U6283 ( .A(n7268), .B(n7269), .Z(n5961) );
  AND U6284 ( .A(n7268), .B(n7270), .Z(n7269) );
  XNOR U6285 ( .A(n7271), .B(n7272), .Z(n5964) );
  AND U6286 ( .A(n7271), .B(n7273), .Z(n7272) );
  XNOR U6287 ( .A(n7274), .B(n7275), .Z(n5967) );
  AND U6288 ( .A(n7274), .B(n7276), .Z(n7275) );
  XNOR U6289 ( .A(n7277), .B(n7278), .Z(n5970) );
  AND U6290 ( .A(n7277), .B(n7279), .Z(n7278) );
  XNOR U6291 ( .A(n7280), .B(n7281), .Z(n5973) );
  AND U6292 ( .A(n7280), .B(n7282), .Z(n7281) );
  XNOR U6293 ( .A(n7283), .B(n7284), .Z(n5976) );
  AND U6294 ( .A(n7283), .B(n7285), .Z(n7284) );
  XNOR U6295 ( .A(n7286), .B(n7287), .Z(n5979) );
  AND U6296 ( .A(n7286), .B(n7288), .Z(n7287) );
  XNOR U6297 ( .A(n7289), .B(n7290), .Z(n5982) );
  AND U6298 ( .A(n7289), .B(n7291), .Z(n7290) );
  XNOR U6299 ( .A(n7292), .B(n7293), .Z(n5985) );
  AND U6300 ( .A(n7292), .B(n7294), .Z(n7293) );
  XNOR U6301 ( .A(n7295), .B(n7296), .Z(n5988) );
  AND U6302 ( .A(n7295), .B(n7297), .Z(n7296) );
  XNOR U6303 ( .A(n7298), .B(n7299), .Z(n5991) );
  AND U6304 ( .A(n7298), .B(n7300), .Z(n7299) );
  XNOR U6305 ( .A(n7301), .B(n7302), .Z(n5994) );
  AND U6306 ( .A(n7301), .B(n7303), .Z(n7302) );
  XNOR U6307 ( .A(n7304), .B(n7305), .Z(n5997) );
  AND U6308 ( .A(n7304), .B(n7306), .Z(n7305) );
  XNOR U6309 ( .A(n7307), .B(n7308), .Z(n6000) );
  AND U6310 ( .A(n7307), .B(n7309), .Z(n7308) );
  XNOR U6311 ( .A(n7310), .B(n7311), .Z(n6003) );
  AND U6312 ( .A(n7310), .B(n7312), .Z(n7311) );
  XNOR U6313 ( .A(n7313), .B(n7314), .Z(n6006) );
  AND U6314 ( .A(n7313), .B(n7315), .Z(n7314) );
  XNOR U6315 ( .A(n7316), .B(n7317), .Z(n6009) );
  AND U6316 ( .A(n7316), .B(n7318), .Z(n7317) );
  XNOR U6317 ( .A(n7319), .B(n7320), .Z(n6012) );
  AND U6318 ( .A(n7319), .B(n7321), .Z(n7320) );
  XNOR U6319 ( .A(n7322), .B(n7323), .Z(n6015) );
  AND U6320 ( .A(n7322), .B(n7324), .Z(n7323) );
  XNOR U6321 ( .A(n7325), .B(n7326), .Z(n6018) );
  AND U6322 ( .A(n7325), .B(n7327), .Z(n7326) );
  XNOR U6323 ( .A(n7328), .B(n7329), .Z(n6021) );
  AND U6324 ( .A(n7328), .B(n7330), .Z(n7329) );
  XNOR U6325 ( .A(n7331), .B(n7332), .Z(n6024) );
  AND U6326 ( .A(n7331), .B(n7333), .Z(n7332) );
  XNOR U6327 ( .A(n7334), .B(n7335), .Z(n6027) );
  AND U6328 ( .A(n7334), .B(n7336), .Z(n7335) );
  XNOR U6329 ( .A(n7337), .B(n7338), .Z(n6030) );
  AND U6330 ( .A(n7337), .B(n7339), .Z(n7338) );
  XNOR U6331 ( .A(n7340), .B(n7341), .Z(n6033) );
  AND U6332 ( .A(n7340), .B(n7342), .Z(n7341) );
  XNOR U6333 ( .A(n7343), .B(n7344), .Z(n6036) );
  AND U6334 ( .A(n7343), .B(n7345), .Z(n7344) );
  XNOR U6335 ( .A(n7346), .B(n7347), .Z(n6039) );
  AND U6336 ( .A(n7346), .B(n7348), .Z(n7347) );
  XNOR U6337 ( .A(n7349), .B(n7350), .Z(n6042) );
  AND U6338 ( .A(n7349), .B(n7351), .Z(n7350) );
  XNOR U6339 ( .A(n7352), .B(n7353), .Z(n6045) );
  AND U6340 ( .A(n7352), .B(n7354), .Z(n7353) );
  XNOR U6341 ( .A(n7355), .B(n7356), .Z(n6048) );
  AND U6342 ( .A(n7355), .B(n7357), .Z(n7356) );
  XNOR U6343 ( .A(n7358), .B(n7359), .Z(n6051) );
  AND U6344 ( .A(n7358), .B(n7360), .Z(n7359) );
  XNOR U6345 ( .A(n7361), .B(n7362), .Z(n6054) );
  AND U6346 ( .A(n7361), .B(n7363), .Z(n7362) );
  XNOR U6347 ( .A(n7364), .B(n7365), .Z(n6057) );
  AND U6348 ( .A(n7364), .B(n7366), .Z(n7365) );
  XNOR U6349 ( .A(n7367), .B(n7368), .Z(n6060) );
  AND U6350 ( .A(n7367), .B(n7369), .Z(n7368) );
  XNOR U6351 ( .A(n7370), .B(n7371), .Z(n6063) );
  AND U6352 ( .A(n7370), .B(n7372), .Z(n7371) );
  XNOR U6353 ( .A(n7373), .B(n7374), .Z(n6066) );
  AND U6354 ( .A(n7373), .B(n7375), .Z(n7374) );
  XNOR U6355 ( .A(n7376), .B(n7377), .Z(n6069) );
  AND U6356 ( .A(n7376), .B(n7378), .Z(n7377) );
  XNOR U6357 ( .A(n7379), .B(n7380), .Z(n6072) );
  AND U6358 ( .A(n7379), .B(n7381), .Z(n7380) );
  XOR U6359 ( .A(n7382), .B(n7383), .Z(n6075) );
  AND U6360 ( .A(n7382), .B(n118), .Z(n7383) );
  XNOR U6361 ( .A(n7384), .B(n6731), .Z(n6733) );
  IV U6362 ( .A(n101), .Z(n7384) );
  XOR U6363 ( .A(n6728), .B(n6727), .Z(n101) );
  XNOR U6364 ( .A(n6725), .B(n6724), .Z(n6727) );
  XNOR U6365 ( .A(n6722), .B(n6721), .Z(n6724) );
  XNOR U6366 ( .A(n6719), .B(n6718), .Z(n6721) );
  XNOR U6367 ( .A(n6716), .B(n6715), .Z(n6718) );
  XNOR U6368 ( .A(n6713), .B(n6712), .Z(n6715) );
  XNOR U6369 ( .A(n6710), .B(n6709), .Z(n6712) );
  XNOR U6370 ( .A(n6707), .B(n6706), .Z(n6709) );
  XNOR U6371 ( .A(n6704), .B(n6703), .Z(n6706) );
  XNOR U6372 ( .A(n6701), .B(n6700), .Z(n6703) );
  XNOR U6373 ( .A(n6698), .B(n6697), .Z(n6700) );
  XNOR U6374 ( .A(n6695), .B(n6694), .Z(n6697) );
  XNOR U6375 ( .A(n6692), .B(n6691), .Z(n6694) );
  XNOR U6376 ( .A(n6689), .B(n6688), .Z(n6691) );
  XNOR U6377 ( .A(n6686), .B(n6685), .Z(n6688) );
  XNOR U6378 ( .A(n6683), .B(n6682), .Z(n6685) );
  XNOR U6379 ( .A(n6680), .B(n6679), .Z(n6682) );
  XNOR U6380 ( .A(n6677), .B(n6676), .Z(n6679) );
  XNOR U6381 ( .A(n6674), .B(n6673), .Z(n6676) );
  XNOR U6382 ( .A(n6671), .B(n6670), .Z(n6673) );
  XNOR U6383 ( .A(n6668), .B(n6667), .Z(n6670) );
  XNOR U6384 ( .A(n6665), .B(n6664), .Z(n6667) );
  XNOR U6385 ( .A(n6662), .B(n6661), .Z(n6664) );
  XNOR U6386 ( .A(n6659), .B(n6658), .Z(n6661) );
  XNOR U6387 ( .A(n6656), .B(n6655), .Z(n6658) );
  XNOR U6388 ( .A(n6653), .B(n6652), .Z(n6655) );
  XNOR U6389 ( .A(n6650), .B(n6649), .Z(n6652) );
  XNOR U6390 ( .A(n6647), .B(n6646), .Z(n6649) );
  XNOR U6391 ( .A(n6644), .B(n6643), .Z(n6646) );
  XNOR U6392 ( .A(n6641), .B(n6640), .Z(n6643) );
  XNOR U6393 ( .A(n6638), .B(n6637), .Z(n6640) );
  XNOR U6394 ( .A(n6635), .B(n6634), .Z(n6637) );
  XNOR U6395 ( .A(n6632), .B(n6631), .Z(n6634) );
  XNOR U6396 ( .A(n6629), .B(n6628), .Z(n6631) );
  XNOR U6397 ( .A(n6626), .B(n6625), .Z(n6628) );
  XNOR U6398 ( .A(n6623), .B(n6622), .Z(n6625) );
  XNOR U6399 ( .A(n6620), .B(n6619), .Z(n6622) );
  XNOR U6400 ( .A(n6617), .B(n6616), .Z(n6619) );
  XNOR U6401 ( .A(n6614), .B(n6613), .Z(n6616) );
  XNOR U6402 ( .A(n6611), .B(n6610), .Z(n6613) );
  XNOR U6403 ( .A(n6608), .B(n6607), .Z(n6610) );
  XNOR U6404 ( .A(n6605), .B(n6604), .Z(n6607) );
  XNOR U6405 ( .A(n6602), .B(n6601), .Z(n6604) );
  XNOR U6406 ( .A(n6599), .B(n6598), .Z(n6601) );
  XNOR U6407 ( .A(n6596), .B(n6595), .Z(n6598) );
  XNOR U6408 ( .A(n6593), .B(n6592), .Z(n6595) );
  XNOR U6409 ( .A(n6590), .B(n6589), .Z(n6592) );
  XNOR U6410 ( .A(n6587), .B(n6586), .Z(n6589) );
  XNOR U6411 ( .A(n6584), .B(n6583), .Z(n6586) );
  XNOR U6412 ( .A(n6581), .B(n6580), .Z(n6583) );
  XNOR U6413 ( .A(n6578), .B(n6577), .Z(n6580) );
  XNOR U6414 ( .A(n6575), .B(n6574), .Z(n6577) );
  XNOR U6415 ( .A(n6572), .B(n6571), .Z(n6574) );
  XNOR U6416 ( .A(n6569), .B(n6568), .Z(n6571) );
  XNOR U6417 ( .A(n6566), .B(n6565), .Z(n6568) );
  XNOR U6418 ( .A(n6563), .B(n6562), .Z(n6565) );
  XNOR U6419 ( .A(n6560), .B(n6559), .Z(n6562) );
  XNOR U6420 ( .A(n6557), .B(n6556), .Z(n6559) );
  XNOR U6421 ( .A(n6554), .B(n6553), .Z(n6556) );
  XNOR U6422 ( .A(n6551), .B(n6550), .Z(n6553) );
  XNOR U6423 ( .A(n6548), .B(n6547), .Z(n6550) );
  XNOR U6424 ( .A(n6545), .B(n6544), .Z(n6547) );
  XNOR U6425 ( .A(n6542), .B(n6541), .Z(n6544) );
  XNOR U6426 ( .A(n6539), .B(n6538), .Z(n6541) );
  XNOR U6427 ( .A(n6536), .B(n6535), .Z(n6538) );
  XNOR U6428 ( .A(n6533), .B(n6532), .Z(n6535) );
  XNOR U6429 ( .A(n6530), .B(n6529), .Z(n6532) );
  XNOR U6430 ( .A(n6527), .B(n6526), .Z(n6529) );
  XNOR U6431 ( .A(n6524), .B(n6523), .Z(n6526) );
  XNOR U6432 ( .A(n6521), .B(n6520), .Z(n6523) );
  XNOR U6433 ( .A(n6518), .B(n6517), .Z(n6520) );
  XNOR U6434 ( .A(n6515), .B(n6514), .Z(n6517) );
  XNOR U6435 ( .A(n6512), .B(n6511), .Z(n6514) );
  XNOR U6436 ( .A(n6509), .B(n6508), .Z(n6511) );
  XNOR U6437 ( .A(n6506), .B(n6505), .Z(n6508) );
  XNOR U6438 ( .A(n6503), .B(n6502), .Z(n6505) );
  XNOR U6439 ( .A(n6500), .B(n6499), .Z(n6502) );
  XNOR U6440 ( .A(n6497), .B(n6496), .Z(n6499) );
  XNOR U6441 ( .A(n6494), .B(n6493), .Z(n6496) );
  XNOR U6442 ( .A(n6491), .B(n6490), .Z(n6493) );
  XNOR U6443 ( .A(n6488), .B(n6487), .Z(n6490) );
  XNOR U6444 ( .A(n6485), .B(n6484), .Z(n6487) );
  XNOR U6445 ( .A(n6482), .B(n6481), .Z(n6484) );
  XNOR U6446 ( .A(n6479), .B(n6478), .Z(n6481) );
  XNOR U6447 ( .A(n6476), .B(n6475), .Z(n6478) );
  XNOR U6448 ( .A(n6473), .B(n6472), .Z(n6475) );
  XNOR U6449 ( .A(n6470), .B(n6469), .Z(n6472) );
  XNOR U6450 ( .A(n6467), .B(n6466), .Z(n6469) );
  XNOR U6451 ( .A(n6464), .B(n6463), .Z(n6466) );
  XNOR U6452 ( .A(n6461), .B(n6460), .Z(n6463) );
  XNOR U6453 ( .A(n6458), .B(n6457), .Z(n6460) );
  XNOR U6454 ( .A(n6455), .B(n6454), .Z(n6457) );
  XNOR U6455 ( .A(n6452), .B(n6451), .Z(n6454) );
  XNOR U6456 ( .A(n6449), .B(n6448), .Z(n6451) );
  XNOR U6457 ( .A(n6446), .B(n6445), .Z(n6448) );
  XNOR U6458 ( .A(n6443), .B(n6442), .Z(n6445) );
  XNOR U6459 ( .A(n6440), .B(n6439), .Z(n6442) );
  XNOR U6460 ( .A(n6437), .B(n6436), .Z(n6439) );
  XNOR U6461 ( .A(n6434), .B(n6433), .Z(n6436) );
  XNOR U6462 ( .A(n6431), .B(n6430), .Z(n6433) );
  XNOR U6463 ( .A(n6428), .B(n6427), .Z(n6430) );
  XNOR U6464 ( .A(n6425), .B(n6424), .Z(n6427) );
  XNOR U6465 ( .A(n6422), .B(n6421), .Z(n6424) );
  XNOR U6466 ( .A(n6419), .B(n6418), .Z(n6421) );
  XNOR U6467 ( .A(n6416), .B(n6415), .Z(n6418) );
  XNOR U6468 ( .A(n6413), .B(n6412), .Z(n6415) );
  XNOR U6469 ( .A(n6410), .B(n6409), .Z(n6412) );
  XNOR U6470 ( .A(n6407), .B(n6406), .Z(n6409) );
  XNOR U6471 ( .A(n6404), .B(n6403), .Z(n6406) );
  XNOR U6472 ( .A(n6401), .B(n6400), .Z(n6403) );
  XNOR U6473 ( .A(n6398), .B(n6397), .Z(n6400) );
  XNOR U6474 ( .A(n6395), .B(n6394), .Z(n6397) );
  XNOR U6475 ( .A(n6392), .B(n6391), .Z(n6394) );
  XNOR U6476 ( .A(n6389), .B(n6388), .Z(n6391) );
  XNOR U6477 ( .A(n6386), .B(n6385), .Z(n6388) );
  XNOR U6478 ( .A(n6383), .B(n6382), .Z(n6385) );
  XNOR U6479 ( .A(n6380), .B(n6379), .Z(n6382) );
  XNOR U6480 ( .A(n6377), .B(n6376), .Z(n6379) );
  XNOR U6481 ( .A(n6374), .B(n6373), .Z(n6376) );
  XNOR U6482 ( .A(n6371), .B(n6370), .Z(n6373) );
  XNOR U6483 ( .A(n6368), .B(n6367), .Z(n6370) );
  XNOR U6484 ( .A(n6365), .B(n6364), .Z(n6367) );
  XNOR U6485 ( .A(n6362), .B(n6361), .Z(n6364) );
  XNOR U6486 ( .A(n6359), .B(n6358), .Z(n6361) );
  XNOR U6487 ( .A(n6356), .B(n6355), .Z(n6358) );
  XNOR U6488 ( .A(n6353), .B(n6352), .Z(n6355) );
  XNOR U6489 ( .A(n6350), .B(n6349), .Z(n6352) );
  XNOR U6490 ( .A(n6347), .B(n6346), .Z(n6349) );
  XNOR U6491 ( .A(n6344), .B(n6343), .Z(n6346) );
  XOR U6492 ( .A(n6341), .B(n6340), .Z(n6343) );
  XOR U6493 ( .A(n6338), .B(n6337), .Z(n6340) );
  XOR U6494 ( .A(n6334), .B(n6335), .Z(n6337) );
  AND U6495 ( .A(n7385), .B(n7386), .Z(n6335) );
  XOR U6496 ( .A(n6331), .B(n6332), .Z(n6334) );
  AND U6497 ( .A(n7387), .B(n7388), .Z(n6332) );
  XOR U6498 ( .A(n6328), .B(n6329), .Z(n6331) );
  AND U6499 ( .A(n7389), .B(n7390), .Z(n6329) );
  XNOR U6500 ( .A(n6078), .B(n6326), .Z(n6328) );
  AND U6501 ( .A(n7391), .B(n7392), .Z(n6326) );
  XOR U6502 ( .A(n6080), .B(n6079), .Z(n6078) );
  AND U6503 ( .A(n7393), .B(n7394), .Z(n6079) );
  XOR U6504 ( .A(n6082), .B(n6081), .Z(n6080) );
  AND U6505 ( .A(n7395), .B(n7396), .Z(n6081) );
  XOR U6506 ( .A(n6084), .B(n6083), .Z(n6082) );
  AND U6507 ( .A(n7397), .B(n7398), .Z(n6083) );
  XOR U6508 ( .A(n6086), .B(n6085), .Z(n6084) );
  AND U6509 ( .A(n7399), .B(n7400), .Z(n6085) );
  XOR U6510 ( .A(n6088), .B(n6087), .Z(n6086) );
  AND U6511 ( .A(n7401), .B(n7402), .Z(n6087) );
  XOR U6512 ( .A(n6090), .B(n6089), .Z(n6088) );
  AND U6513 ( .A(n7403), .B(n7404), .Z(n6089) );
  XOR U6514 ( .A(n6092), .B(n6091), .Z(n6090) );
  AND U6515 ( .A(n7405), .B(n7406), .Z(n6091) );
  XOR U6516 ( .A(n6094), .B(n6093), .Z(n6092) );
  AND U6517 ( .A(n7407), .B(n7408), .Z(n6093) );
  XOR U6518 ( .A(n6096), .B(n6095), .Z(n6094) );
  AND U6519 ( .A(n7409), .B(n7410), .Z(n6095) );
  XOR U6520 ( .A(n6098), .B(n6097), .Z(n6096) );
  AND U6521 ( .A(n7411), .B(n7412), .Z(n6097) );
  XOR U6522 ( .A(n6100), .B(n6099), .Z(n6098) );
  AND U6523 ( .A(n7413), .B(n7414), .Z(n6099) );
  XOR U6524 ( .A(n6102), .B(n6101), .Z(n6100) );
  AND U6525 ( .A(n7415), .B(n7416), .Z(n6101) );
  XOR U6526 ( .A(n6104), .B(n6103), .Z(n6102) );
  AND U6527 ( .A(n7417), .B(n7418), .Z(n6103) );
  XOR U6528 ( .A(n6106), .B(n6105), .Z(n6104) );
  AND U6529 ( .A(n7419), .B(n7420), .Z(n6105) );
  XOR U6530 ( .A(n6108), .B(n6107), .Z(n6106) );
  AND U6531 ( .A(n7421), .B(n7422), .Z(n6107) );
  XOR U6532 ( .A(n6110), .B(n6109), .Z(n6108) );
  AND U6533 ( .A(n7423), .B(n7424), .Z(n6109) );
  XOR U6534 ( .A(n6112), .B(n6111), .Z(n6110) );
  AND U6535 ( .A(n7425), .B(n7426), .Z(n6111) );
  XOR U6536 ( .A(n6114), .B(n6113), .Z(n6112) );
  AND U6537 ( .A(n7427), .B(n7428), .Z(n6113) );
  XOR U6538 ( .A(n6116), .B(n6115), .Z(n6114) );
  AND U6539 ( .A(n7429), .B(n7430), .Z(n6115) );
  XOR U6540 ( .A(n6118), .B(n6117), .Z(n6116) );
  AND U6541 ( .A(n7431), .B(n7432), .Z(n6117) );
  XOR U6542 ( .A(n6120), .B(n6119), .Z(n6118) );
  AND U6543 ( .A(n7433), .B(n7434), .Z(n6119) );
  XOR U6544 ( .A(n6122), .B(n6121), .Z(n6120) );
  AND U6545 ( .A(n7435), .B(n7436), .Z(n6121) );
  XOR U6546 ( .A(n6124), .B(n6123), .Z(n6122) );
  AND U6547 ( .A(n7437), .B(n7438), .Z(n6123) );
  XOR U6548 ( .A(n6126), .B(n6125), .Z(n6124) );
  AND U6549 ( .A(n7439), .B(n7440), .Z(n6125) );
  XOR U6550 ( .A(n6128), .B(n6127), .Z(n6126) );
  AND U6551 ( .A(n7441), .B(n7442), .Z(n6127) );
  XOR U6552 ( .A(n6130), .B(n6129), .Z(n6128) );
  AND U6553 ( .A(n7443), .B(n7444), .Z(n6129) );
  XOR U6554 ( .A(n6132), .B(n6131), .Z(n6130) );
  AND U6555 ( .A(n7445), .B(n7446), .Z(n6131) );
  XOR U6556 ( .A(n6134), .B(n6133), .Z(n6132) );
  AND U6557 ( .A(n7447), .B(n7448), .Z(n6133) );
  XOR U6558 ( .A(n6136), .B(n6135), .Z(n6134) );
  AND U6559 ( .A(n7449), .B(n7450), .Z(n6135) );
  XOR U6560 ( .A(n6138), .B(n6137), .Z(n6136) );
  AND U6561 ( .A(n7451), .B(n7452), .Z(n6137) );
  XOR U6562 ( .A(n6140), .B(n6139), .Z(n6138) );
  AND U6563 ( .A(n7453), .B(n7454), .Z(n6139) );
  XOR U6564 ( .A(n6142), .B(n6141), .Z(n6140) );
  AND U6565 ( .A(n7455), .B(n7456), .Z(n6141) );
  XOR U6566 ( .A(n6144), .B(n6143), .Z(n6142) );
  AND U6567 ( .A(n7457), .B(n7458), .Z(n6143) );
  XOR U6568 ( .A(n6146), .B(n6145), .Z(n6144) );
  AND U6569 ( .A(n7459), .B(n7460), .Z(n6145) );
  XOR U6570 ( .A(n6148), .B(n6147), .Z(n6146) );
  AND U6571 ( .A(n7461), .B(n7462), .Z(n6147) );
  XOR U6572 ( .A(n6150), .B(n6149), .Z(n6148) );
  AND U6573 ( .A(n7463), .B(n7464), .Z(n6149) );
  XOR U6574 ( .A(n6152), .B(n6151), .Z(n6150) );
  AND U6575 ( .A(n7465), .B(n7466), .Z(n6151) );
  XOR U6576 ( .A(n6154), .B(n6153), .Z(n6152) );
  AND U6577 ( .A(n7467), .B(n7468), .Z(n6153) );
  XOR U6578 ( .A(n6156), .B(n6155), .Z(n6154) );
  AND U6579 ( .A(n7469), .B(n7470), .Z(n6155) );
  XOR U6580 ( .A(n6158), .B(n6157), .Z(n6156) );
  AND U6581 ( .A(n7471), .B(n7472), .Z(n6157) );
  XOR U6582 ( .A(n6160), .B(n6159), .Z(n6158) );
  AND U6583 ( .A(n7473), .B(n7474), .Z(n6159) );
  XOR U6584 ( .A(n6162), .B(n6161), .Z(n6160) );
  AND U6585 ( .A(n7475), .B(n7476), .Z(n6161) );
  XOR U6586 ( .A(n6164), .B(n6163), .Z(n6162) );
  AND U6587 ( .A(n7477), .B(n7478), .Z(n6163) );
  XOR U6588 ( .A(n6166), .B(n6165), .Z(n6164) );
  AND U6589 ( .A(n7479), .B(n7480), .Z(n6165) );
  XOR U6590 ( .A(n6168), .B(n6167), .Z(n6166) );
  AND U6591 ( .A(n7481), .B(n7482), .Z(n6167) );
  XOR U6592 ( .A(n6170), .B(n6169), .Z(n6168) );
  AND U6593 ( .A(n7483), .B(n7484), .Z(n6169) );
  XOR U6594 ( .A(n6172), .B(n6171), .Z(n6170) );
  AND U6595 ( .A(n7485), .B(n7486), .Z(n6171) );
  XOR U6596 ( .A(n6174), .B(n6173), .Z(n6172) );
  AND U6597 ( .A(n7487), .B(n7488), .Z(n6173) );
  XOR U6598 ( .A(n6176), .B(n6175), .Z(n6174) );
  AND U6599 ( .A(n7489), .B(n7490), .Z(n6175) );
  XOR U6600 ( .A(n6178), .B(n6177), .Z(n6176) );
  AND U6601 ( .A(n7491), .B(n7492), .Z(n6177) );
  XOR U6602 ( .A(n6180), .B(n6179), .Z(n6178) );
  AND U6603 ( .A(n7493), .B(n7494), .Z(n6179) );
  XOR U6604 ( .A(n6182), .B(n6181), .Z(n6180) );
  AND U6605 ( .A(n7495), .B(n7496), .Z(n6181) );
  XOR U6606 ( .A(n6184), .B(n6183), .Z(n6182) );
  AND U6607 ( .A(n7497), .B(n7498), .Z(n6183) );
  XOR U6608 ( .A(n6186), .B(n6185), .Z(n6184) );
  AND U6609 ( .A(n7499), .B(n7500), .Z(n6185) );
  XOR U6610 ( .A(n6188), .B(n6187), .Z(n6186) );
  AND U6611 ( .A(n7501), .B(n7502), .Z(n6187) );
  XOR U6612 ( .A(n6190), .B(n6189), .Z(n6188) );
  AND U6613 ( .A(n7503), .B(n7504), .Z(n6189) );
  XOR U6614 ( .A(n6192), .B(n6191), .Z(n6190) );
  AND U6615 ( .A(n7505), .B(n7506), .Z(n6191) );
  XOR U6616 ( .A(n6194), .B(n6193), .Z(n6192) );
  AND U6617 ( .A(n7507), .B(n7508), .Z(n6193) );
  XOR U6618 ( .A(n6196), .B(n6195), .Z(n6194) );
  AND U6619 ( .A(n7509), .B(n7510), .Z(n6195) );
  XOR U6620 ( .A(n6198), .B(n6197), .Z(n6196) );
  AND U6621 ( .A(n7511), .B(n7512), .Z(n6197) );
  XOR U6622 ( .A(n6200), .B(n6199), .Z(n6198) );
  AND U6623 ( .A(n7513), .B(n7514), .Z(n6199) );
  XOR U6624 ( .A(n6202), .B(n6201), .Z(n6200) );
  AND U6625 ( .A(n7515), .B(n7516), .Z(n6201) );
  XOR U6626 ( .A(n6204), .B(n6203), .Z(n6202) );
  AND U6627 ( .A(n7517), .B(n7518), .Z(n6203) );
  XOR U6628 ( .A(n6206), .B(n6205), .Z(n6204) );
  AND U6629 ( .A(n7519), .B(n7520), .Z(n6205) );
  XOR U6630 ( .A(n6208), .B(n6207), .Z(n6206) );
  AND U6631 ( .A(n7521), .B(n7522), .Z(n6207) );
  XOR U6632 ( .A(n6210), .B(n6209), .Z(n6208) );
  AND U6633 ( .A(n7523), .B(n7524), .Z(n6209) );
  XOR U6634 ( .A(n6212), .B(n6211), .Z(n6210) );
  AND U6635 ( .A(n7525), .B(n7526), .Z(n6211) );
  XOR U6636 ( .A(n6214), .B(n6213), .Z(n6212) );
  AND U6637 ( .A(n7527), .B(n7528), .Z(n6213) );
  XOR U6638 ( .A(n6216), .B(n6215), .Z(n6214) );
  AND U6639 ( .A(n7529), .B(n7530), .Z(n6215) );
  XOR U6640 ( .A(n6218), .B(n6217), .Z(n6216) );
  AND U6641 ( .A(n7531), .B(n7532), .Z(n6217) );
  XOR U6642 ( .A(n6220), .B(n6219), .Z(n6218) );
  AND U6643 ( .A(n7533), .B(n7534), .Z(n6219) );
  XOR U6644 ( .A(n6222), .B(n6221), .Z(n6220) );
  AND U6645 ( .A(n7535), .B(n7536), .Z(n6221) );
  XOR U6646 ( .A(n6224), .B(n6223), .Z(n6222) );
  AND U6647 ( .A(n7537), .B(n7538), .Z(n6223) );
  XOR U6648 ( .A(n6226), .B(n6225), .Z(n6224) );
  AND U6649 ( .A(n7539), .B(n7540), .Z(n6225) );
  XOR U6650 ( .A(n6228), .B(n6227), .Z(n6226) );
  AND U6651 ( .A(n7541), .B(n7542), .Z(n6227) );
  XOR U6652 ( .A(n6230), .B(n6229), .Z(n6228) );
  AND U6653 ( .A(n7543), .B(n7544), .Z(n6229) );
  XOR U6654 ( .A(n6232), .B(n6231), .Z(n6230) );
  AND U6655 ( .A(n7545), .B(n7546), .Z(n6231) );
  XOR U6656 ( .A(n6234), .B(n6233), .Z(n6232) );
  AND U6657 ( .A(n7547), .B(n7548), .Z(n6233) );
  XOR U6658 ( .A(n6236), .B(n6235), .Z(n6234) );
  AND U6659 ( .A(n7549), .B(n7550), .Z(n6235) );
  XOR U6660 ( .A(n6238), .B(n6237), .Z(n6236) );
  AND U6661 ( .A(n7551), .B(n7552), .Z(n6237) );
  XOR U6662 ( .A(n6240), .B(n6239), .Z(n6238) );
  AND U6663 ( .A(n7553), .B(n7554), .Z(n6239) );
  XOR U6664 ( .A(n6242), .B(n6241), .Z(n6240) );
  AND U6665 ( .A(n7555), .B(n7556), .Z(n6241) );
  XOR U6666 ( .A(n6244), .B(n6243), .Z(n6242) );
  AND U6667 ( .A(n7557), .B(n7558), .Z(n6243) );
  XOR U6668 ( .A(n6246), .B(n6245), .Z(n6244) );
  AND U6669 ( .A(n7559), .B(n7560), .Z(n6245) );
  XOR U6670 ( .A(n6248), .B(n6247), .Z(n6246) );
  AND U6671 ( .A(n7561), .B(n7562), .Z(n6247) );
  XOR U6672 ( .A(n6250), .B(n6249), .Z(n6248) );
  AND U6673 ( .A(n7563), .B(n7564), .Z(n6249) );
  XOR U6674 ( .A(n6252), .B(n6251), .Z(n6250) );
  AND U6675 ( .A(n7565), .B(n7566), .Z(n6251) );
  XOR U6676 ( .A(n6254), .B(n6253), .Z(n6252) );
  AND U6677 ( .A(n7567), .B(n7568), .Z(n6253) );
  XOR U6678 ( .A(n6256), .B(n6255), .Z(n6254) );
  AND U6679 ( .A(n7569), .B(n7570), .Z(n6255) );
  XOR U6680 ( .A(n6258), .B(n6257), .Z(n6256) );
  AND U6681 ( .A(n7571), .B(n7572), .Z(n6257) );
  XOR U6682 ( .A(n6260), .B(n6259), .Z(n6258) );
  AND U6683 ( .A(n7573), .B(n7574), .Z(n6259) );
  XOR U6684 ( .A(n6262), .B(n6261), .Z(n6260) );
  AND U6685 ( .A(n7575), .B(n7576), .Z(n6261) );
  XOR U6686 ( .A(n6264), .B(n6263), .Z(n6262) );
  AND U6687 ( .A(n7577), .B(n7578), .Z(n6263) );
  XOR U6688 ( .A(n6266), .B(n6265), .Z(n6264) );
  AND U6689 ( .A(n7579), .B(n7580), .Z(n6265) );
  XOR U6690 ( .A(n6268), .B(n6267), .Z(n6266) );
  AND U6691 ( .A(n7581), .B(n7582), .Z(n6267) );
  XOR U6692 ( .A(n6270), .B(n6269), .Z(n6268) );
  AND U6693 ( .A(n7583), .B(n7584), .Z(n6269) );
  XOR U6694 ( .A(n6322), .B(n6271), .Z(n6270) );
  AND U6695 ( .A(n7585), .B(n7586), .Z(n6271) );
  XOR U6696 ( .A(n6324), .B(n6323), .Z(n6322) );
  AND U6697 ( .A(n7587), .B(n7588), .Z(n6323) );
  XOR U6698 ( .A(n6306), .B(n6325), .Z(n6324) );
  AND U6699 ( .A(n7589), .B(n7590), .Z(n6325) );
  XOR U6700 ( .A(n6308), .B(n6307), .Z(n6306) );
  AND U6701 ( .A(n7591), .B(n7592), .Z(n6307) );
  XOR U6702 ( .A(n6310), .B(n6309), .Z(n6308) );
  AND U6703 ( .A(n7593), .B(n7594), .Z(n6309) );
  XOR U6704 ( .A(n6314), .B(n6311), .Z(n6310) );
  AND U6705 ( .A(n7595), .B(n7596), .Z(n6311) );
  XOR U6706 ( .A(n6316), .B(n6315), .Z(n6314) );
  AND U6707 ( .A(n7597), .B(n7598), .Z(n6315) );
  XOR U6708 ( .A(n6318), .B(n6317), .Z(n6316) );
  AND U6709 ( .A(n7599), .B(n7600), .Z(n6317) );
  XOR U6710 ( .A(n6320), .B(n6319), .Z(n6318) );
  AND U6711 ( .A(n7601), .B(n7602), .Z(n6319) );
  XOR U6712 ( .A(n6295), .B(n6321), .Z(n6320) );
  AND U6713 ( .A(n7603), .B(n7604), .Z(n6321) );
  XNOR U6714 ( .A(n6292), .B(n6296), .Z(n6295) );
  AND U6715 ( .A(n7605), .B(n7606), .Z(n6296) );
  XOR U6716 ( .A(n6291), .B(n6283), .Z(n6292) );
  AND U6717 ( .A(n7607), .B(n7608), .Z(n6283) );
  XNOR U6718 ( .A(n6286), .B(n6282), .Z(n6291) );
  AND U6719 ( .A(n7609), .B(n7610), .Z(n6282) );
  XOR U6720 ( .A(n7611), .B(n7612), .Z(n6286) );
  XOR U6721 ( .A(n6304), .B(n7613), .Z(n7612) );
  XOR U6722 ( .A(n6302), .B(n6300), .Z(n7613) );
  AND U6723 ( .A(n7614), .B(n7615), .Z(n6300) );
  AND U6724 ( .A(n7616), .B(n7617), .Z(n6302) );
  AND U6725 ( .A(n7618), .B(n7619), .Z(n6304) );
  XNOR U6726 ( .A(n7620), .B(n6303), .Z(n7611) );
  XOR U6727 ( .A(n7621), .B(n7622), .Z(n6303) );
  XOR U6728 ( .A(n7623), .B(n7624), .Z(n7622) );
  AND U6729 ( .A(n7625), .B(n7626), .Z(n7624) );
  XNOR U6730 ( .A(n7627), .B(n7628), .Z(n7621) );
  NOR U6731 ( .A(n7629), .B(n7630), .Z(n7628) );
  AND U6732 ( .A(n7631), .B(n7632), .Z(n7630) );
  IV U6733 ( .A(n7633), .Z(n7629) );
  NOR U6734 ( .A(n7623), .B(n7634), .Z(n7633) );
  AND U6735 ( .A(n7635), .B(n7636), .Z(n7634) );
  NOR U6736 ( .A(n7625), .B(n7635), .Z(n7627) );
  XNOR U6737 ( .A(n6305), .B(n6287), .Z(n7620) );
  AND U6738 ( .A(n7637), .B(n7638), .Z(n6287) );
  AND U6739 ( .A(n7639), .B(n7640), .Z(n6305) );
  XOR U6740 ( .A(n7641), .B(n7642), .Z(n6338) );
  NOR U6741 ( .A(n7643), .B(n7644), .Z(n7642) );
  IV U6742 ( .A(n7641), .Z(n7643) );
  XOR U6743 ( .A(n7645), .B(n7646), .Z(n6341) );
  NOR U6744 ( .A(n7645), .B(n7647), .Z(n7646) );
  XNOR U6745 ( .A(n7648), .B(n7649), .Z(n6344) );
  AND U6746 ( .A(n7648), .B(n7650), .Z(n7649) );
  XNOR U6747 ( .A(n7651), .B(n7652), .Z(n6347) );
  AND U6748 ( .A(n7651), .B(n7653), .Z(n7652) );
  XNOR U6749 ( .A(n7654), .B(n7655), .Z(n6350) );
  AND U6750 ( .A(n7654), .B(n7656), .Z(n7655) );
  XNOR U6751 ( .A(n7657), .B(n7658), .Z(n6353) );
  AND U6752 ( .A(n7657), .B(n7659), .Z(n7658) );
  XNOR U6753 ( .A(n7660), .B(n7661), .Z(n6356) );
  AND U6754 ( .A(n7660), .B(n7662), .Z(n7661) );
  XNOR U6755 ( .A(n7663), .B(n7664), .Z(n6359) );
  AND U6756 ( .A(n7663), .B(n7665), .Z(n7664) );
  XNOR U6757 ( .A(n7666), .B(n7667), .Z(n6362) );
  AND U6758 ( .A(n7666), .B(n7668), .Z(n7667) );
  XNOR U6759 ( .A(n7669), .B(n7670), .Z(n6365) );
  AND U6760 ( .A(n7669), .B(n7671), .Z(n7670) );
  XNOR U6761 ( .A(n7672), .B(n7673), .Z(n6368) );
  AND U6762 ( .A(n7672), .B(n7674), .Z(n7673) );
  XNOR U6763 ( .A(n7675), .B(n7676), .Z(n6371) );
  AND U6764 ( .A(n7675), .B(n7677), .Z(n7676) );
  XNOR U6765 ( .A(n7678), .B(n7679), .Z(n6374) );
  AND U6766 ( .A(n7678), .B(n7680), .Z(n7679) );
  XNOR U6767 ( .A(n7681), .B(n7682), .Z(n6377) );
  AND U6768 ( .A(n7681), .B(n7683), .Z(n7682) );
  XNOR U6769 ( .A(n7684), .B(n7685), .Z(n6380) );
  AND U6770 ( .A(n7684), .B(n7686), .Z(n7685) );
  XNOR U6771 ( .A(n7687), .B(n7688), .Z(n6383) );
  AND U6772 ( .A(n7687), .B(n7689), .Z(n7688) );
  XNOR U6773 ( .A(n7690), .B(n7691), .Z(n6386) );
  AND U6774 ( .A(n7690), .B(n7692), .Z(n7691) );
  XNOR U6775 ( .A(n7693), .B(n7694), .Z(n6389) );
  AND U6776 ( .A(n7693), .B(n7695), .Z(n7694) );
  XNOR U6777 ( .A(n7696), .B(n7697), .Z(n6392) );
  AND U6778 ( .A(n7696), .B(n7698), .Z(n7697) );
  XNOR U6779 ( .A(n7699), .B(n7700), .Z(n6395) );
  AND U6780 ( .A(n7699), .B(n7701), .Z(n7700) );
  XNOR U6781 ( .A(n7702), .B(n7703), .Z(n6398) );
  AND U6782 ( .A(n7702), .B(n7704), .Z(n7703) );
  XNOR U6783 ( .A(n7705), .B(n7706), .Z(n6401) );
  AND U6784 ( .A(n7705), .B(n7707), .Z(n7706) );
  XNOR U6785 ( .A(n7708), .B(n7709), .Z(n6404) );
  AND U6786 ( .A(n7708), .B(n7710), .Z(n7709) );
  XNOR U6787 ( .A(n7711), .B(n7712), .Z(n6407) );
  AND U6788 ( .A(n7711), .B(n7713), .Z(n7712) );
  XNOR U6789 ( .A(n7714), .B(n7715), .Z(n6410) );
  AND U6790 ( .A(n7714), .B(n7716), .Z(n7715) );
  XNOR U6791 ( .A(n7717), .B(n7718), .Z(n6413) );
  AND U6792 ( .A(n7717), .B(n7719), .Z(n7718) );
  XNOR U6793 ( .A(n7720), .B(n7721), .Z(n6416) );
  AND U6794 ( .A(n7720), .B(n7722), .Z(n7721) );
  XNOR U6795 ( .A(n7723), .B(n7724), .Z(n6419) );
  AND U6796 ( .A(n7723), .B(n7725), .Z(n7724) );
  XNOR U6797 ( .A(n7726), .B(n7727), .Z(n6422) );
  AND U6798 ( .A(n7726), .B(n7728), .Z(n7727) );
  XNOR U6799 ( .A(n7729), .B(n7730), .Z(n6425) );
  AND U6800 ( .A(n7729), .B(n7731), .Z(n7730) );
  XNOR U6801 ( .A(n7732), .B(n7733), .Z(n6428) );
  AND U6802 ( .A(n7732), .B(n7734), .Z(n7733) );
  XNOR U6803 ( .A(n7735), .B(n7736), .Z(n6431) );
  AND U6804 ( .A(n7735), .B(n7737), .Z(n7736) );
  XNOR U6805 ( .A(n7738), .B(n7739), .Z(n6434) );
  AND U6806 ( .A(n7738), .B(n7740), .Z(n7739) );
  XNOR U6807 ( .A(n7741), .B(n7742), .Z(n6437) );
  AND U6808 ( .A(n7741), .B(n7743), .Z(n7742) );
  XNOR U6809 ( .A(n7744), .B(n7745), .Z(n6440) );
  AND U6810 ( .A(n7744), .B(n7746), .Z(n7745) );
  XNOR U6811 ( .A(n7747), .B(n7748), .Z(n6443) );
  AND U6812 ( .A(n7747), .B(n7749), .Z(n7748) );
  XNOR U6813 ( .A(n7750), .B(n7751), .Z(n6446) );
  AND U6814 ( .A(n7750), .B(n7752), .Z(n7751) );
  XNOR U6815 ( .A(n7753), .B(n7754), .Z(n6449) );
  AND U6816 ( .A(n7753), .B(n7755), .Z(n7754) );
  XNOR U6817 ( .A(n7756), .B(n7757), .Z(n6452) );
  AND U6818 ( .A(n7756), .B(n7758), .Z(n7757) );
  XNOR U6819 ( .A(n7759), .B(n7760), .Z(n6455) );
  AND U6820 ( .A(n7759), .B(n7761), .Z(n7760) );
  XNOR U6821 ( .A(n7762), .B(n7763), .Z(n6458) );
  AND U6822 ( .A(n7762), .B(n7764), .Z(n7763) );
  XNOR U6823 ( .A(n7765), .B(n7766), .Z(n6461) );
  AND U6824 ( .A(n7765), .B(n7767), .Z(n7766) );
  XNOR U6825 ( .A(n7768), .B(n7769), .Z(n6464) );
  AND U6826 ( .A(n7768), .B(n7770), .Z(n7769) );
  XNOR U6827 ( .A(n7771), .B(n7772), .Z(n6467) );
  AND U6828 ( .A(n7771), .B(n7773), .Z(n7772) );
  XNOR U6829 ( .A(n7774), .B(n7775), .Z(n6470) );
  AND U6830 ( .A(n7774), .B(n7776), .Z(n7775) );
  XNOR U6831 ( .A(n7777), .B(n7778), .Z(n6473) );
  AND U6832 ( .A(n7777), .B(n7779), .Z(n7778) );
  XNOR U6833 ( .A(n7780), .B(n7781), .Z(n6476) );
  AND U6834 ( .A(n7780), .B(n7782), .Z(n7781) );
  XNOR U6835 ( .A(n7783), .B(n7784), .Z(n6479) );
  AND U6836 ( .A(n7783), .B(n7785), .Z(n7784) );
  XNOR U6837 ( .A(n7786), .B(n7787), .Z(n6482) );
  AND U6838 ( .A(n7786), .B(n7788), .Z(n7787) );
  XNOR U6839 ( .A(n7789), .B(n7790), .Z(n6485) );
  AND U6840 ( .A(n7789), .B(n7791), .Z(n7790) );
  XNOR U6841 ( .A(n7792), .B(n7793), .Z(n6488) );
  AND U6842 ( .A(n7792), .B(n7794), .Z(n7793) );
  XNOR U6843 ( .A(n7795), .B(n7796), .Z(n6491) );
  AND U6844 ( .A(n7795), .B(n7797), .Z(n7796) );
  XNOR U6845 ( .A(n7798), .B(n7799), .Z(n6494) );
  AND U6846 ( .A(n7798), .B(n7800), .Z(n7799) );
  XNOR U6847 ( .A(n7801), .B(n7802), .Z(n6497) );
  AND U6848 ( .A(n7801), .B(n7803), .Z(n7802) );
  XNOR U6849 ( .A(n7804), .B(n7805), .Z(n6500) );
  AND U6850 ( .A(n7804), .B(n7806), .Z(n7805) );
  XNOR U6851 ( .A(n7807), .B(n7808), .Z(n6503) );
  AND U6852 ( .A(n7807), .B(n7809), .Z(n7808) );
  XNOR U6853 ( .A(n7810), .B(n7811), .Z(n6506) );
  AND U6854 ( .A(n7810), .B(n7812), .Z(n7811) );
  XNOR U6855 ( .A(n7813), .B(n7814), .Z(n6509) );
  AND U6856 ( .A(n7813), .B(n7815), .Z(n7814) );
  XNOR U6857 ( .A(n7816), .B(n7817), .Z(n6512) );
  AND U6858 ( .A(n7816), .B(n7818), .Z(n7817) );
  XNOR U6859 ( .A(n7819), .B(n7820), .Z(n6515) );
  AND U6860 ( .A(n7819), .B(n7821), .Z(n7820) );
  XNOR U6861 ( .A(n7822), .B(n7823), .Z(n6518) );
  AND U6862 ( .A(n7822), .B(n7824), .Z(n7823) );
  XNOR U6863 ( .A(n7825), .B(n7826), .Z(n6521) );
  AND U6864 ( .A(n7825), .B(n7827), .Z(n7826) );
  XNOR U6865 ( .A(n7828), .B(n7829), .Z(n6524) );
  AND U6866 ( .A(n7828), .B(n7830), .Z(n7829) );
  XNOR U6867 ( .A(n7831), .B(n7832), .Z(n6527) );
  AND U6868 ( .A(n7831), .B(n7833), .Z(n7832) );
  XNOR U6869 ( .A(n7834), .B(n7835), .Z(n6530) );
  AND U6870 ( .A(n7834), .B(n7836), .Z(n7835) );
  XNOR U6871 ( .A(n7837), .B(n7838), .Z(n6533) );
  AND U6872 ( .A(n7837), .B(n7839), .Z(n7838) );
  XNOR U6873 ( .A(n7840), .B(n7841), .Z(n6536) );
  AND U6874 ( .A(n7840), .B(n7842), .Z(n7841) );
  XNOR U6875 ( .A(n7843), .B(n7844), .Z(n6539) );
  AND U6876 ( .A(n7843), .B(n7845), .Z(n7844) );
  XNOR U6877 ( .A(n7846), .B(n7847), .Z(n6542) );
  AND U6878 ( .A(n7846), .B(n7848), .Z(n7847) );
  XNOR U6879 ( .A(n7849), .B(n7850), .Z(n6545) );
  AND U6880 ( .A(n7849), .B(n7851), .Z(n7850) );
  XNOR U6881 ( .A(n7852), .B(n7853), .Z(n6548) );
  AND U6882 ( .A(n7852), .B(n7854), .Z(n7853) );
  XNOR U6883 ( .A(n7855), .B(n7856), .Z(n6551) );
  AND U6884 ( .A(n7855), .B(n7857), .Z(n7856) );
  XNOR U6885 ( .A(n7858), .B(n7859), .Z(n6554) );
  AND U6886 ( .A(n7858), .B(n7860), .Z(n7859) );
  XNOR U6887 ( .A(n7861), .B(n7862), .Z(n6557) );
  AND U6888 ( .A(n7861), .B(n7863), .Z(n7862) );
  XNOR U6889 ( .A(n7864), .B(n7865), .Z(n6560) );
  AND U6890 ( .A(n7864), .B(n7866), .Z(n7865) );
  XNOR U6891 ( .A(n7867), .B(n7868), .Z(n6563) );
  AND U6892 ( .A(n7867), .B(n7869), .Z(n7868) );
  XNOR U6893 ( .A(n7870), .B(n7871), .Z(n6566) );
  AND U6894 ( .A(n7870), .B(n7872), .Z(n7871) );
  XNOR U6895 ( .A(n7873), .B(n7874), .Z(n6569) );
  AND U6896 ( .A(n7873), .B(n7875), .Z(n7874) );
  XNOR U6897 ( .A(n7876), .B(n7877), .Z(n6572) );
  AND U6898 ( .A(n7876), .B(n7878), .Z(n7877) );
  XNOR U6899 ( .A(n7879), .B(n7880), .Z(n6575) );
  AND U6900 ( .A(n7879), .B(n7881), .Z(n7880) );
  XNOR U6901 ( .A(n7882), .B(n7883), .Z(n6578) );
  AND U6902 ( .A(n7882), .B(n7884), .Z(n7883) );
  XNOR U6903 ( .A(n7885), .B(n7886), .Z(n6581) );
  AND U6904 ( .A(n7885), .B(n7887), .Z(n7886) );
  XNOR U6905 ( .A(n7888), .B(n7889), .Z(n6584) );
  AND U6906 ( .A(n7888), .B(n7890), .Z(n7889) );
  XNOR U6907 ( .A(n7891), .B(n7892), .Z(n6587) );
  AND U6908 ( .A(n7891), .B(n7893), .Z(n7892) );
  XNOR U6909 ( .A(n7894), .B(n7895), .Z(n6590) );
  AND U6910 ( .A(n7894), .B(n7896), .Z(n7895) );
  XNOR U6911 ( .A(n7897), .B(n7898), .Z(n6593) );
  AND U6912 ( .A(n7897), .B(n7899), .Z(n7898) );
  XNOR U6913 ( .A(n7900), .B(n7901), .Z(n6596) );
  AND U6914 ( .A(n7900), .B(n7902), .Z(n7901) );
  XNOR U6915 ( .A(n7903), .B(n7904), .Z(n6599) );
  AND U6916 ( .A(n7903), .B(n7905), .Z(n7904) );
  XNOR U6917 ( .A(n7906), .B(n7907), .Z(n6602) );
  AND U6918 ( .A(n7906), .B(n7908), .Z(n7907) );
  XNOR U6919 ( .A(n7909), .B(n7910), .Z(n6605) );
  AND U6920 ( .A(n7909), .B(n7911), .Z(n7910) );
  XNOR U6921 ( .A(n7912), .B(n7913), .Z(n6608) );
  AND U6922 ( .A(n7912), .B(n7914), .Z(n7913) );
  XNOR U6923 ( .A(n7915), .B(n7916), .Z(n6611) );
  AND U6924 ( .A(n7915), .B(n7917), .Z(n7916) );
  XNOR U6925 ( .A(n7918), .B(n7919), .Z(n6614) );
  AND U6926 ( .A(n7918), .B(n7920), .Z(n7919) );
  XNOR U6927 ( .A(n7921), .B(n7922), .Z(n6617) );
  AND U6928 ( .A(n7921), .B(n7923), .Z(n7922) );
  XNOR U6929 ( .A(n7924), .B(n7925), .Z(n6620) );
  AND U6930 ( .A(n7924), .B(n7926), .Z(n7925) );
  XNOR U6931 ( .A(n7927), .B(n7928), .Z(n6623) );
  AND U6932 ( .A(n7927), .B(n7929), .Z(n7928) );
  XNOR U6933 ( .A(n7930), .B(n7931), .Z(n6626) );
  AND U6934 ( .A(n7930), .B(n7932), .Z(n7931) );
  XNOR U6935 ( .A(n7933), .B(n7934), .Z(n6629) );
  AND U6936 ( .A(n7933), .B(n7935), .Z(n7934) );
  XNOR U6937 ( .A(n7936), .B(n7937), .Z(n6632) );
  AND U6938 ( .A(n7936), .B(n7938), .Z(n7937) );
  XNOR U6939 ( .A(n7939), .B(n7940), .Z(n6635) );
  AND U6940 ( .A(n7939), .B(n7941), .Z(n7940) );
  XNOR U6941 ( .A(n7942), .B(n7943), .Z(n6638) );
  AND U6942 ( .A(n7942), .B(n7944), .Z(n7943) );
  XNOR U6943 ( .A(n7945), .B(n7946), .Z(n6641) );
  AND U6944 ( .A(n7945), .B(n7947), .Z(n7946) );
  XNOR U6945 ( .A(n7948), .B(n7949), .Z(n6644) );
  AND U6946 ( .A(n7948), .B(n7950), .Z(n7949) );
  XNOR U6947 ( .A(n7951), .B(n7952), .Z(n6647) );
  AND U6948 ( .A(n7951), .B(n7953), .Z(n7952) );
  XNOR U6949 ( .A(n7954), .B(n7955), .Z(n6650) );
  AND U6950 ( .A(n7954), .B(n7956), .Z(n7955) );
  XNOR U6951 ( .A(n7957), .B(n7958), .Z(n6653) );
  AND U6952 ( .A(n7957), .B(n7959), .Z(n7958) );
  XNOR U6953 ( .A(n7960), .B(n7961), .Z(n6656) );
  AND U6954 ( .A(n7960), .B(n7962), .Z(n7961) );
  XNOR U6955 ( .A(n7963), .B(n7964), .Z(n6659) );
  AND U6956 ( .A(n7963), .B(n7965), .Z(n7964) );
  XNOR U6957 ( .A(n7966), .B(n7967), .Z(n6662) );
  AND U6958 ( .A(n7966), .B(n7968), .Z(n7967) );
  XNOR U6959 ( .A(n7969), .B(n7970), .Z(n6665) );
  AND U6960 ( .A(n7969), .B(n7971), .Z(n7970) );
  XNOR U6961 ( .A(n7972), .B(n7973), .Z(n6668) );
  AND U6962 ( .A(n7972), .B(n7974), .Z(n7973) );
  XNOR U6963 ( .A(n7975), .B(n7976), .Z(n6671) );
  AND U6964 ( .A(n7975), .B(n7977), .Z(n7976) );
  XNOR U6965 ( .A(n7978), .B(n7979), .Z(n6674) );
  AND U6966 ( .A(n7978), .B(n7980), .Z(n7979) );
  XNOR U6967 ( .A(n7981), .B(n7982), .Z(n6677) );
  AND U6968 ( .A(n7981), .B(n7983), .Z(n7982) );
  XNOR U6969 ( .A(n7984), .B(n7985), .Z(n6680) );
  AND U6970 ( .A(n7984), .B(n7986), .Z(n7985) );
  XNOR U6971 ( .A(n7987), .B(n7988), .Z(n6683) );
  AND U6972 ( .A(n7987), .B(n7989), .Z(n7988) );
  XNOR U6973 ( .A(n7990), .B(n7991), .Z(n6686) );
  AND U6974 ( .A(n7990), .B(n7992), .Z(n7991) );
  XNOR U6975 ( .A(n7993), .B(n7994), .Z(n6689) );
  AND U6976 ( .A(n7993), .B(n7995), .Z(n7994) );
  XNOR U6977 ( .A(n7996), .B(n7997), .Z(n6692) );
  AND U6978 ( .A(n7996), .B(n7998), .Z(n7997) );
  XNOR U6979 ( .A(n7999), .B(n8000), .Z(n6695) );
  AND U6980 ( .A(n7999), .B(n8001), .Z(n8000) );
  XNOR U6981 ( .A(n8002), .B(n8003), .Z(n6698) );
  AND U6982 ( .A(n8002), .B(n8004), .Z(n8003) );
  XNOR U6983 ( .A(n8005), .B(n8006), .Z(n6701) );
  AND U6984 ( .A(n8005), .B(n8007), .Z(n8006) );
  XNOR U6985 ( .A(n8008), .B(n8009), .Z(n6704) );
  AND U6986 ( .A(n8008), .B(n8010), .Z(n8009) );
  XNOR U6987 ( .A(n8011), .B(n8012), .Z(n6707) );
  AND U6988 ( .A(n8011), .B(n8013), .Z(n8012) );
  XNOR U6989 ( .A(n8014), .B(n8015), .Z(n6710) );
  AND U6990 ( .A(n8014), .B(n8016), .Z(n8015) );
  XNOR U6991 ( .A(n8017), .B(n8018), .Z(n6713) );
  AND U6992 ( .A(n8017), .B(n8019), .Z(n8018) );
  XNOR U6993 ( .A(n8020), .B(n8021), .Z(n6716) );
  AND U6994 ( .A(n8020), .B(n8022), .Z(n8021) );
  XNOR U6995 ( .A(n8023), .B(n8024), .Z(n6719) );
  AND U6996 ( .A(n8023), .B(n8025), .Z(n8024) );
  XNOR U6997 ( .A(n8026), .B(n8027), .Z(n6722) );
  AND U6998 ( .A(n8026), .B(n8028), .Z(n8027) );
  XNOR U6999 ( .A(n8029), .B(n8030), .Z(n6725) );
  AND U7000 ( .A(n8029), .B(n8031), .Z(n8030) );
  IV U7001 ( .A(n6730), .Z(n6728) );
  XNOR U7002 ( .A(n8032), .B(n8033), .Z(n6730) );
  AND U7003 ( .A(n8032), .B(n114), .Z(n8033) );
  XOR U7004 ( .A(n8034), .B(n8035), .Z(n6731) );
  AND U7005 ( .A(n8036), .B(n8037), .Z(n8035) );
  XOR U7006 ( .A(n118), .B(n8034), .Z(n8037) );
  XOR U7007 ( .A(n7381), .B(n7382), .Z(n118) );
  AND U7008 ( .A(n8038), .B(n8039), .Z(n7382) );
  XOR U7009 ( .A(n7378), .B(n7379), .Z(n7381) );
  AND U7010 ( .A(n8040), .B(n8041), .Z(n7379) );
  XOR U7011 ( .A(n7375), .B(n7376), .Z(n7378) );
  AND U7012 ( .A(n8042), .B(n8043), .Z(n7376) );
  XOR U7013 ( .A(n7372), .B(n7373), .Z(n7375) );
  AND U7014 ( .A(n8044), .B(n8045), .Z(n7373) );
  XOR U7015 ( .A(n7369), .B(n7370), .Z(n7372) );
  AND U7016 ( .A(n8046), .B(n8047), .Z(n7370) );
  XOR U7017 ( .A(n7366), .B(n7367), .Z(n7369) );
  AND U7018 ( .A(n8048), .B(n8049), .Z(n7367) );
  XOR U7019 ( .A(n7363), .B(n7364), .Z(n7366) );
  AND U7020 ( .A(n8050), .B(n8051), .Z(n7364) );
  XOR U7021 ( .A(n7360), .B(n7361), .Z(n7363) );
  AND U7022 ( .A(n8052), .B(n8053), .Z(n7361) );
  XOR U7023 ( .A(n7357), .B(n7358), .Z(n7360) );
  AND U7024 ( .A(n8054), .B(n8055), .Z(n7358) );
  XOR U7025 ( .A(n7354), .B(n7355), .Z(n7357) );
  AND U7026 ( .A(n8056), .B(n8057), .Z(n7355) );
  XOR U7027 ( .A(n7351), .B(n7352), .Z(n7354) );
  AND U7028 ( .A(n8058), .B(n8059), .Z(n7352) );
  XOR U7029 ( .A(n7348), .B(n7349), .Z(n7351) );
  AND U7030 ( .A(n8060), .B(n8061), .Z(n7349) );
  XOR U7031 ( .A(n7345), .B(n7346), .Z(n7348) );
  AND U7032 ( .A(n8062), .B(n8063), .Z(n7346) );
  XOR U7033 ( .A(n7342), .B(n7343), .Z(n7345) );
  AND U7034 ( .A(n8064), .B(n8065), .Z(n7343) );
  XOR U7035 ( .A(n7339), .B(n7340), .Z(n7342) );
  AND U7036 ( .A(n8066), .B(n8067), .Z(n7340) );
  XOR U7037 ( .A(n7336), .B(n7337), .Z(n7339) );
  AND U7038 ( .A(n8068), .B(n8069), .Z(n7337) );
  XOR U7039 ( .A(n7333), .B(n7334), .Z(n7336) );
  AND U7040 ( .A(n8070), .B(n8071), .Z(n7334) );
  XOR U7041 ( .A(n7330), .B(n7331), .Z(n7333) );
  AND U7042 ( .A(n8072), .B(n8073), .Z(n7331) );
  XOR U7043 ( .A(n7327), .B(n7328), .Z(n7330) );
  AND U7044 ( .A(n8074), .B(n8075), .Z(n7328) );
  XOR U7045 ( .A(n7324), .B(n7325), .Z(n7327) );
  AND U7046 ( .A(n8076), .B(n8077), .Z(n7325) );
  XOR U7047 ( .A(n7321), .B(n7322), .Z(n7324) );
  AND U7048 ( .A(n8078), .B(n8079), .Z(n7322) );
  XOR U7049 ( .A(n7318), .B(n7319), .Z(n7321) );
  AND U7050 ( .A(n8080), .B(n8081), .Z(n7319) );
  XOR U7051 ( .A(n7315), .B(n7316), .Z(n7318) );
  AND U7052 ( .A(n8082), .B(n8083), .Z(n7316) );
  XOR U7053 ( .A(n7312), .B(n7313), .Z(n7315) );
  AND U7054 ( .A(n8084), .B(n8085), .Z(n7313) );
  XOR U7055 ( .A(n7309), .B(n7310), .Z(n7312) );
  AND U7056 ( .A(n8086), .B(n8087), .Z(n7310) );
  XOR U7057 ( .A(n7306), .B(n7307), .Z(n7309) );
  AND U7058 ( .A(n8088), .B(n8089), .Z(n7307) );
  XOR U7059 ( .A(n7303), .B(n7304), .Z(n7306) );
  AND U7060 ( .A(n8090), .B(n8091), .Z(n7304) );
  XOR U7061 ( .A(n7300), .B(n7301), .Z(n7303) );
  AND U7062 ( .A(n8092), .B(n8093), .Z(n7301) );
  XOR U7063 ( .A(n7297), .B(n7298), .Z(n7300) );
  AND U7064 ( .A(n8094), .B(n8095), .Z(n7298) );
  XOR U7065 ( .A(n7294), .B(n7295), .Z(n7297) );
  AND U7066 ( .A(n8096), .B(n8097), .Z(n7295) );
  XOR U7067 ( .A(n7291), .B(n7292), .Z(n7294) );
  AND U7068 ( .A(n8098), .B(n8099), .Z(n7292) );
  XOR U7069 ( .A(n7288), .B(n7289), .Z(n7291) );
  AND U7070 ( .A(n8100), .B(n8101), .Z(n7289) );
  XOR U7071 ( .A(n7285), .B(n7286), .Z(n7288) );
  AND U7072 ( .A(n8102), .B(n8103), .Z(n7286) );
  XOR U7073 ( .A(n7282), .B(n7283), .Z(n7285) );
  AND U7074 ( .A(n8104), .B(n8105), .Z(n7283) );
  XOR U7075 ( .A(n7279), .B(n7280), .Z(n7282) );
  AND U7076 ( .A(n8106), .B(n8107), .Z(n7280) );
  XOR U7077 ( .A(n7276), .B(n7277), .Z(n7279) );
  AND U7078 ( .A(n8108), .B(n8109), .Z(n7277) );
  XOR U7079 ( .A(n7273), .B(n7274), .Z(n7276) );
  AND U7080 ( .A(n8110), .B(n8111), .Z(n7274) );
  XOR U7081 ( .A(n7270), .B(n7271), .Z(n7273) );
  AND U7082 ( .A(n8112), .B(n8113), .Z(n7271) );
  XOR U7083 ( .A(n7267), .B(n7268), .Z(n7270) );
  AND U7084 ( .A(n8114), .B(n8115), .Z(n7268) );
  XOR U7085 ( .A(n7264), .B(n7265), .Z(n7267) );
  AND U7086 ( .A(n8116), .B(n8117), .Z(n7265) );
  XOR U7087 ( .A(n7261), .B(n7262), .Z(n7264) );
  AND U7088 ( .A(n8118), .B(n8119), .Z(n7262) );
  XOR U7089 ( .A(n7258), .B(n7259), .Z(n7261) );
  AND U7090 ( .A(n8120), .B(n8121), .Z(n7259) );
  XOR U7091 ( .A(n7255), .B(n7256), .Z(n7258) );
  AND U7092 ( .A(n8122), .B(n8123), .Z(n7256) );
  XOR U7093 ( .A(n7252), .B(n7253), .Z(n7255) );
  AND U7094 ( .A(n8124), .B(n8125), .Z(n7253) );
  XOR U7095 ( .A(n7249), .B(n7250), .Z(n7252) );
  AND U7096 ( .A(n8126), .B(n8127), .Z(n7250) );
  XOR U7097 ( .A(n7246), .B(n7247), .Z(n7249) );
  AND U7098 ( .A(n8128), .B(n8129), .Z(n7247) );
  XOR U7099 ( .A(n7243), .B(n7244), .Z(n7246) );
  AND U7100 ( .A(n8130), .B(n8131), .Z(n7244) );
  XOR U7101 ( .A(n7240), .B(n7241), .Z(n7243) );
  AND U7102 ( .A(n8132), .B(n8133), .Z(n7241) );
  XOR U7103 ( .A(n7237), .B(n7238), .Z(n7240) );
  AND U7104 ( .A(n8134), .B(n8135), .Z(n7238) );
  XOR U7105 ( .A(n7234), .B(n7235), .Z(n7237) );
  AND U7106 ( .A(n8136), .B(n8137), .Z(n7235) );
  XOR U7107 ( .A(n7231), .B(n7232), .Z(n7234) );
  AND U7108 ( .A(n8138), .B(n8139), .Z(n7232) );
  XOR U7109 ( .A(n7228), .B(n7229), .Z(n7231) );
  AND U7110 ( .A(n8140), .B(n8141), .Z(n7229) );
  XOR U7111 ( .A(n7225), .B(n7226), .Z(n7228) );
  AND U7112 ( .A(n8142), .B(n8143), .Z(n7226) );
  XOR U7113 ( .A(n7222), .B(n7223), .Z(n7225) );
  AND U7114 ( .A(n8144), .B(n8145), .Z(n7223) );
  XOR U7115 ( .A(n7219), .B(n7220), .Z(n7222) );
  AND U7116 ( .A(n8146), .B(n8147), .Z(n7220) );
  XOR U7117 ( .A(n7216), .B(n7217), .Z(n7219) );
  AND U7118 ( .A(n8148), .B(n8149), .Z(n7217) );
  XOR U7119 ( .A(n7213), .B(n7214), .Z(n7216) );
  AND U7120 ( .A(n8150), .B(n8151), .Z(n7214) );
  XOR U7121 ( .A(n7210), .B(n7211), .Z(n7213) );
  AND U7122 ( .A(n8152), .B(n8153), .Z(n7211) );
  XOR U7123 ( .A(n7207), .B(n7208), .Z(n7210) );
  AND U7124 ( .A(n8154), .B(n8155), .Z(n7208) );
  XOR U7125 ( .A(n7204), .B(n7205), .Z(n7207) );
  AND U7126 ( .A(n8156), .B(n8157), .Z(n7205) );
  XOR U7127 ( .A(n7201), .B(n7202), .Z(n7204) );
  AND U7128 ( .A(n8158), .B(n8159), .Z(n7202) );
  XOR U7129 ( .A(n7198), .B(n7199), .Z(n7201) );
  AND U7130 ( .A(n8160), .B(n8161), .Z(n7199) );
  XOR U7131 ( .A(n7195), .B(n7196), .Z(n7198) );
  AND U7132 ( .A(n8162), .B(n8163), .Z(n7196) );
  XOR U7133 ( .A(n7192), .B(n7193), .Z(n7195) );
  AND U7134 ( .A(n8164), .B(n8165), .Z(n7193) );
  XOR U7135 ( .A(n7189), .B(n7190), .Z(n7192) );
  AND U7136 ( .A(n8166), .B(n8167), .Z(n7190) );
  XOR U7137 ( .A(n7186), .B(n7187), .Z(n7189) );
  AND U7138 ( .A(n8168), .B(n8169), .Z(n7187) );
  XOR U7139 ( .A(n7183), .B(n7184), .Z(n7186) );
  AND U7140 ( .A(n8170), .B(n8171), .Z(n7184) );
  XOR U7141 ( .A(n7180), .B(n7181), .Z(n7183) );
  AND U7142 ( .A(n8172), .B(n8173), .Z(n7181) );
  XOR U7143 ( .A(n7177), .B(n7178), .Z(n7180) );
  AND U7144 ( .A(n8174), .B(n8175), .Z(n7178) );
  XOR U7145 ( .A(n7174), .B(n7175), .Z(n7177) );
  AND U7146 ( .A(n8176), .B(n8177), .Z(n7175) );
  XOR U7147 ( .A(n7171), .B(n7172), .Z(n7174) );
  AND U7148 ( .A(n8178), .B(n8179), .Z(n7172) );
  XOR U7149 ( .A(n7168), .B(n7169), .Z(n7171) );
  AND U7150 ( .A(n8180), .B(n8181), .Z(n7169) );
  XOR U7151 ( .A(n7165), .B(n7166), .Z(n7168) );
  AND U7152 ( .A(n8182), .B(n8183), .Z(n7166) );
  XOR U7153 ( .A(n7162), .B(n7163), .Z(n7165) );
  AND U7154 ( .A(n8184), .B(n8185), .Z(n7163) );
  XOR U7155 ( .A(n7159), .B(n7160), .Z(n7162) );
  AND U7156 ( .A(n8186), .B(n8187), .Z(n7160) );
  XOR U7157 ( .A(n7156), .B(n7157), .Z(n7159) );
  AND U7158 ( .A(n8188), .B(n8189), .Z(n7157) );
  XOR U7159 ( .A(n7153), .B(n7154), .Z(n7156) );
  AND U7160 ( .A(n8190), .B(n8191), .Z(n7154) );
  XOR U7161 ( .A(n7150), .B(n7151), .Z(n7153) );
  AND U7162 ( .A(n8192), .B(n8193), .Z(n7151) );
  XOR U7163 ( .A(n7147), .B(n7148), .Z(n7150) );
  AND U7164 ( .A(n8194), .B(n8195), .Z(n7148) );
  XOR U7165 ( .A(n7144), .B(n7145), .Z(n7147) );
  AND U7166 ( .A(n8196), .B(n8197), .Z(n7145) );
  XOR U7167 ( .A(n7141), .B(n7142), .Z(n7144) );
  AND U7168 ( .A(n8198), .B(n8199), .Z(n7142) );
  XOR U7169 ( .A(n7138), .B(n7139), .Z(n7141) );
  AND U7170 ( .A(n8200), .B(n8201), .Z(n7139) );
  XOR U7171 ( .A(n7135), .B(n7136), .Z(n7138) );
  AND U7172 ( .A(n8202), .B(n8203), .Z(n7136) );
  XOR U7173 ( .A(n7132), .B(n7133), .Z(n7135) );
  AND U7174 ( .A(n8204), .B(n8205), .Z(n7133) );
  XOR U7175 ( .A(n7129), .B(n7130), .Z(n7132) );
  AND U7176 ( .A(n8206), .B(n8207), .Z(n7130) );
  XOR U7177 ( .A(n7126), .B(n7127), .Z(n7129) );
  AND U7178 ( .A(n8208), .B(n8209), .Z(n7127) );
  XOR U7179 ( .A(n7123), .B(n7124), .Z(n7126) );
  AND U7180 ( .A(n8210), .B(n8211), .Z(n7124) );
  XOR U7181 ( .A(n7120), .B(n7121), .Z(n7123) );
  AND U7182 ( .A(n8212), .B(n8213), .Z(n7121) );
  XOR U7183 ( .A(n7117), .B(n7118), .Z(n7120) );
  AND U7184 ( .A(n8214), .B(n8215), .Z(n7118) );
  XOR U7185 ( .A(n7114), .B(n7115), .Z(n7117) );
  AND U7186 ( .A(n8216), .B(n8217), .Z(n7115) );
  XOR U7187 ( .A(n7111), .B(n7112), .Z(n7114) );
  AND U7188 ( .A(n8218), .B(n8219), .Z(n7112) );
  XOR U7189 ( .A(n7108), .B(n7109), .Z(n7111) );
  AND U7190 ( .A(n8220), .B(n8221), .Z(n7109) );
  XOR U7191 ( .A(n7105), .B(n7106), .Z(n7108) );
  AND U7192 ( .A(n8222), .B(n8223), .Z(n7106) );
  XOR U7193 ( .A(n7102), .B(n7103), .Z(n7105) );
  AND U7194 ( .A(n8224), .B(n8225), .Z(n7103) );
  XOR U7195 ( .A(n7099), .B(n7100), .Z(n7102) );
  AND U7196 ( .A(n8226), .B(n8227), .Z(n7100) );
  XOR U7197 ( .A(n7096), .B(n7097), .Z(n7099) );
  AND U7198 ( .A(n8228), .B(n8229), .Z(n7097) );
  XOR U7199 ( .A(n7093), .B(n7094), .Z(n7096) );
  AND U7200 ( .A(n8230), .B(n8231), .Z(n7094) );
  XOR U7201 ( .A(n7090), .B(n7091), .Z(n7093) );
  AND U7202 ( .A(n8232), .B(n8233), .Z(n7091) );
  XOR U7203 ( .A(n7087), .B(n7088), .Z(n7090) );
  AND U7204 ( .A(n8234), .B(n8235), .Z(n7088) );
  XOR U7205 ( .A(n7084), .B(n7085), .Z(n7087) );
  AND U7206 ( .A(n8236), .B(n8237), .Z(n7085) );
  XOR U7207 ( .A(n7081), .B(n7082), .Z(n7084) );
  AND U7208 ( .A(n8238), .B(n8239), .Z(n7082) );
  XOR U7209 ( .A(n7078), .B(n7079), .Z(n7081) );
  AND U7210 ( .A(n8240), .B(n8241), .Z(n7079) );
  XOR U7211 ( .A(n7075), .B(n7076), .Z(n7078) );
  AND U7212 ( .A(n8242), .B(n8243), .Z(n7076) );
  XOR U7213 ( .A(n7072), .B(n7073), .Z(n7075) );
  AND U7214 ( .A(n8244), .B(n8245), .Z(n7073) );
  XOR U7215 ( .A(n7069), .B(n7070), .Z(n7072) );
  AND U7216 ( .A(n8246), .B(n8247), .Z(n7070) );
  XOR U7217 ( .A(n7066), .B(n7067), .Z(n7069) );
  AND U7218 ( .A(n8248), .B(n8249), .Z(n7067) );
  XOR U7219 ( .A(n7063), .B(n7064), .Z(n7066) );
  AND U7220 ( .A(n8250), .B(n8251), .Z(n7064) );
  XOR U7221 ( .A(n7060), .B(n7061), .Z(n7063) );
  AND U7222 ( .A(n8252), .B(n8253), .Z(n7061) );
  XOR U7223 ( .A(n7057), .B(n7058), .Z(n7060) );
  AND U7224 ( .A(n8254), .B(n8255), .Z(n7058) );
  XOR U7225 ( .A(n7054), .B(n7055), .Z(n7057) );
  AND U7226 ( .A(n8256), .B(n8257), .Z(n7055) );
  XOR U7227 ( .A(n7051), .B(n7052), .Z(n7054) );
  AND U7228 ( .A(n8258), .B(n8259), .Z(n7052) );
  XOR U7229 ( .A(n7048), .B(n7049), .Z(n7051) );
  AND U7230 ( .A(n8260), .B(n8261), .Z(n7049) );
  XOR U7231 ( .A(n7045), .B(n7046), .Z(n7048) );
  AND U7232 ( .A(n8262), .B(n8263), .Z(n7046) );
  XOR U7233 ( .A(n7042), .B(n7043), .Z(n7045) );
  AND U7234 ( .A(n8264), .B(n8265), .Z(n7043) );
  XOR U7235 ( .A(n7039), .B(n7040), .Z(n7042) );
  AND U7236 ( .A(n8266), .B(n8267), .Z(n7040) );
  XOR U7237 ( .A(n7036), .B(n7037), .Z(n7039) );
  AND U7238 ( .A(n8268), .B(n8269), .Z(n7037) );
  XOR U7239 ( .A(n7033), .B(n7034), .Z(n7036) );
  AND U7240 ( .A(n8270), .B(n8271), .Z(n7034) );
  XOR U7241 ( .A(n7030), .B(n7031), .Z(n7033) );
  AND U7242 ( .A(n8272), .B(n8273), .Z(n7031) );
  XOR U7243 ( .A(n7027), .B(n7028), .Z(n7030) );
  AND U7244 ( .A(n8274), .B(n8275), .Z(n7028) );
  XOR U7245 ( .A(n7024), .B(n7025), .Z(n7027) );
  AND U7246 ( .A(n8276), .B(n8277), .Z(n7025) );
  XOR U7247 ( .A(n7021), .B(n7022), .Z(n7024) );
  AND U7248 ( .A(n8278), .B(n8279), .Z(n7022) );
  XOR U7249 ( .A(n7018), .B(n7019), .Z(n7021) );
  AND U7250 ( .A(n8280), .B(n8281), .Z(n7019) );
  XOR U7251 ( .A(n7015), .B(n7016), .Z(n7018) );
  AND U7252 ( .A(n8282), .B(n8283), .Z(n7016) );
  XOR U7253 ( .A(n7012), .B(n7013), .Z(n7015) );
  AND U7254 ( .A(n8284), .B(n8285), .Z(n7013) );
  XOR U7255 ( .A(n7009), .B(n7010), .Z(n7012) );
  AND U7256 ( .A(n8286), .B(n8287), .Z(n7010) );
  XOR U7257 ( .A(n7006), .B(n7007), .Z(n7009) );
  AND U7258 ( .A(n8288), .B(n8289), .Z(n7007) );
  XOR U7259 ( .A(n7003), .B(n7004), .Z(n7006) );
  AND U7260 ( .A(n8290), .B(n8291), .Z(n7004) );
  XOR U7261 ( .A(n7000), .B(n7001), .Z(n7003) );
  AND U7262 ( .A(n8292), .B(n8293), .Z(n7001) );
  XNOR U7263 ( .A(n6997), .B(n6998), .Z(n7000) );
  AND U7264 ( .A(n8294), .B(n8295), .Z(n6998) );
  XOR U7265 ( .A(n8296), .B(n6995), .Z(n6997) );
  IV U7266 ( .A(n8297), .Z(n6995) );
  AND U7267 ( .A(n8298), .B(n8299), .Z(n8297) );
  IV U7268 ( .A(n6994), .Z(n8296) );
  XOR U7269 ( .A(n6735), .B(n6991), .Z(n6994) );
  AND U7270 ( .A(n8300), .B(n8301), .Z(n6991) );
  XOR U7271 ( .A(n6737), .B(n6736), .Z(n6735) );
  AND U7272 ( .A(n8302), .B(n8303), .Z(n6736) );
  XOR U7273 ( .A(n6739), .B(n6738), .Z(n6737) );
  AND U7274 ( .A(n8304), .B(n8305), .Z(n6738) );
  XOR U7275 ( .A(n6741), .B(n6740), .Z(n6739) );
  AND U7276 ( .A(n8306), .B(n8307), .Z(n6740) );
  XOR U7277 ( .A(n6743), .B(n6742), .Z(n6741) );
  AND U7278 ( .A(n8308), .B(n8309), .Z(n6742) );
  XOR U7279 ( .A(n6745), .B(n6744), .Z(n6743) );
  AND U7280 ( .A(n8310), .B(n8311), .Z(n6744) );
  XOR U7281 ( .A(n6747), .B(n6746), .Z(n6745) );
  AND U7282 ( .A(n8312), .B(n8313), .Z(n6746) );
  XOR U7283 ( .A(n6749), .B(n6748), .Z(n6747) );
  AND U7284 ( .A(n8314), .B(n8315), .Z(n6748) );
  XOR U7285 ( .A(n6751), .B(n6750), .Z(n6749) );
  AND U7286 ( .A(n8316), .B(n8317), .Z(n6750) );
  XOR U7287 ( .A(n6753), .B(n6752), .Z(n6751) );
  AND U7288 ( .A(n8318), .B(n8319), .Z(n6752) );
  XOR U7289 ( .A(n6755), .B(n6754), .Z(n6753) );
  AND U7290 ( .A(n8320), .B(n8321), .Z(n6754) );
  XOR U7291 ( .A(n6757), .B(n6756), .Z(n6755) );
  AND U7292 ( .A(n8322), .B(n8323), .Z(n6756) );
  XOR U7293 ( .A(n6759), .B(n6758), .Z(n6757) );
  AND U7294 ( .A(n8324), .B(n8325), .Z(n6758) );
  XOR U7295 ( .A(n6761), .B(n6760), .Z(n6759) );
  AND U7296 ( .A(n8326), .B(n8327), .Z(n6760) );
  XOR U7297 ( .A(n6763), .B(n6762), .Z(n6761) );
  AND U7298 ( .A(n8328), .B(n8329), .Z(n6762) );
  XOR U7299 ( .A(n6765), .B(n6764), .Z(n6763) );
  AND U7300 ( .A(n8330), .B(n8331), .Z(n6764) );
  XOR U7301 ( .A(n6767), .B(n6766), .Z(n6765) );
  AND U7302 ( .A(n8332), .B(n8333), .Z(n6766) );
  XOR U7303 ( .A(n6769), .B(n6768), .Z(n6767) );
  AND U7304 ( .A(n8334), .B(n8335), .Z(n6768) );
  XOR U7305 ( .A(n6771), .B(n6770), .Z(n6769) );
  AND U7306 ( .A(n8336), .B(n8337), .Z(n6770) );
  XOR U7307 ( .A(n6773), .B(n6772), .Z(n6771) );
  AND U7308 ( .A(n8338), .B(n8339), .Z(n6772) );
  XOR U7309 ( .A(n6775), .B(n6774), .Z(n6773) );
  AND U7310 ( .A(n8340), .B(n8341), .Z(n6774) );
  XOR U7311 ( .A(n6777), .B(n6776), .Z(n6775) );
  AND U7312 ( .A(n8342), .B(n8343), .Z(n6776) );
  XOR U7313 ( .A(n6779), .B(n6778), .Z(n6777) );
  AND U7314 ( .A(n8344), .B(n8345), .Z(n6778) );
  XOR U7315 ( .A(n6781), .B(n6780), .Z(n6779) );
  AND U7316 ( .A(n8346), .B(n8347), .Z(n6780) );
  XOR U7317 ( .A(n6783), .B(n6782), .Z(n6781) );
  AND U7318 ( .A(n8348), .B(n8349), .Z(n6782) );
  XOR U7319 ( .A(n6785), .B(n6784), .Z(n6783) );
  AND U7320 ( .A(n8350), .B(n8351), .Z(n6784) );
  XOR U7321 ( .A(n6787), .B(n6786), .Z(n6785) );
  AND U7322 ( .A(n8352), .B(n8353), .Z(n6786) );
  XOR U7323 ( .A(n6789), .B(n6788), .Z(n6787) );
  AND U7324 ( .A(n8354), .B(n8355), .Z(n6788) );
  XOR U7325 ( .A(n6791), .B(n6790), .Z(n6789) );
  AND U7326 ( .A(n8356), .B(n8357), .Z(n6790) );
  XOR U7327 ( .A(n6793), .B(n6792), .Z(n6791) );
  AND U7328 ( .A(n8358), .B(n8359), .Z(n6792) );
  XOR U7329 ( .A(n6795), .B(n6794), .Z(n6793) );
  AND U7330 ( .A(n8360), .B(n8361), .Z(n6794) );
  XOR U7331 ( .A(n6797), .B(n6796), .Z(n6795) );
  AND U7332 ( .A(n8362), .B(n8363), .Z(n6796) );
  XOR U7333 ( .A(n6799), .B(n6798), .Z(n6797) );
  AND U7334 ( .A(n8364), .B(n8365), .Z(n6798) );
  XOR U7335 ( .A(n6801), .B(n6800), .Z(n6799) );
  AND U7336 ( .A(n8366), .B(n8367), .Z(n6800) );
  XOR U7337 ( .A(n6803), .B(n6802), .Z(n6801) );
  AND U7338 ( .A(n8368), .B(n8369), .Z(n6802) );
  XOR U7339 ( .A(n6805), .B(n6804), .Z(n6803) );
  AND U7340 ( .A(n8370), .B(n8371), .Z(n6804) );
  XOR U7341 ( .A(n6807), .B(n6806), .Z(n6805) );
  AND U7342 ( .A(n8372), .B(n8373), .Z(n6806) );
  XOR U7343 ( .A(n6809), .B(n6808), .Z(n6807) );
  AND U7344 ( .A(n8374), .B(n8375), .Z(n6808) );
  XOR U7345 ( .A(n6811), .B(n6810), .Z(n6809) );
  AND U7346 ( .A(n8376), .B(n8377), .Z(n6810) );
  XOR U7347 ( .A(n6813), .B(n6812), .Z(n6811) );
  AND U7348 ( .A(n8378), .B(n8379), .Z(n6812) );
  XOR U7349 ( .A(n6815), .B(n6814), .Z(n6813) );
  AND U7350 ( .A(n8380), .B(n8381), .Z(n6814) );
  XOR U7351 ( .A(n6817), .B(n6816), .Z(n6815) );
  AND U7352 ( .A(n8382), .B(n8383), .Z(n6816) );
  XOR U7353 ( .A(n6819), .B(n6818), .Z(n6817) );
  AND U7354 ( .A(n8384), .B(n8385), .Z(n6818) );
  XOR U7355 ( .A(n6821), .B(n6820), .Z(n6819) );
  AND U7356 ( .A(n8386), .B(n8387), .Z(n6820) );
  XOR U7357 ( .A(n6823), .B(n6822), .Z(n6821) );
  AND U7358 ( .A(n8388), .B(n8389), .Z(n6822) );
  XOR U7359 ( .A(n6825), .B(n6824), .Z(n6823) );
  AND U7360 ( .A(n8390), .B(n8391), .Z(n6824) );
  XOR U7361 ( .A(n6827), .B(n6826), .Z(n6825) );
  AND U7362 ( .A(n8392), .B(n8393), .Z(n6826) );
  XOR U7363 ( .A(n6829), .B(n6828), .Z(n6827) );
  AND U7364 ( .A(n8394), .B(n8395), .Z(n6828) );
  XOR U7365 ( .A(n6831), .B(n6830), .Z(n6829) );
  AND U7366 ( .A(n8396), .B(n8397), .Z(n6830) );
  XOR U7367 ( .A(n6833), .B(n6832), .Z(n6831) );
  AND U7368 ( .A(n8398), .B(n8399), .Z(n6832) );
  XOR U7369 ( .A(n6835), .B(n6834), .Z(n6833) );
  AND U7370 ( .A(n8400), .B(n8401), .Z(n6834) );
  XOR U7371 ( .A(n6837), .B(n6836), .Z(n6835) );
  AND U7372 ( .A(n8402), .B(n8403), .Z(n6836) );
  XOR U7373 ( .A(n6839), .B(n6838), .Z(n6837) );
  AND U7374 ( .A(n8404), .B(n8405), .Z(n6838) );
  XOR U7375 ( .A(n6841), .B(n6840), .Z(n6839) );
  AND U7376 ( .A(n8406), .B(n8407), .Z(n6840) );
  XOR U7377 ( .A(n6843), .B(n6842), .Z(n6841) );
  AND U7378 ( .A(n8408), .B(n8409), .Z(n6842) );
  XOR U7379 ( .A(n6845), .B(n6844), .Z(n6843) );
  AND U7380 ( .A(n8410), .B(n8411), .Z(n6844) );
  XOR U7381 ( .A(n6847), .B(n6846), .Z(n6845) );
  AND U7382 ( .A(n8412), .B(n8413), .Z(n6846) );
  XOR U7383 ( .A(n6849), .B(n6848), .Z(n6847) );
  AND U7384 ( .A(n8414), .B(n8415), .Z(n6848) );
  XOR U7385 ( .A(n6851), .B(n6850), .Z(n6849) );
  AND U7386 ( .A(n8416), .B(n8417), .Z(n6850) );
  XOR U7387 ( .A(n6853), .B(n6852), .Z(n6851) );
  AND U7388 ( .A(n8418), .B(n8419), .Z(n6852) );
  XOR U7389 ( .A(n6855), .B(n6854), .Z(n6853) );
  AND U7390 ( .A(n8420), .B(n8421), .Z(n6854) );
  XOR U7391 ( .A(n6857), .B(n6856), .Z(n6855) );
  AND U7392 ( .A(n8422), .B(n8423), .Z(n6856) );
  XOR U7393 ( .A(n6859), .B(n6858), .Z(n6857) );
  AND U7394 ( .A(n8424), .B(n8425), .Z(n6858) );
  XOR U7395 ( .A(n6861), .B(n6860), .Z(n6859) );
  AND U7396 ( .A(n8426), .B(n8427), .Z(n6860) );
  XOR U7397 ( .A(n6863), .B(n6862), .Z(n6861) );
  AND U7398 ( .A(n8428), .B(n8429), .Z(n6862) );
  XOR U7399 ( .A(n6865), .B(n6864), .Z(n6863) );
  AND U7400 ( .A(n8430), .B(n8431), .Z(n6864) );
  XOR U7401 ( .A(n6867), .B(n6866), .Z(n6865) );
  AND U7402 ( .A(n8432), .B(n8433), .Z(n6866) );
  XOR U7403 ( .A(n6869), .B(n6868), .Z(n6867) );
  AND U7404 ( .A(n8434), .B(n8435), .Z(n6868) );
  XOR U7405 ( .A(n6871), .B(n6870), .Z(n6869) );
  AND U7406 ( .A(n8436), .B(n8437), .Z(n6870) );
  XOR U7407 ( .A(n6873), .B(n6872), .Z(n6871) );
  AND U7408 ( .A(n8438), .B(n8439), .Z(n6872) );
  XOR U7409 ( .A(n6875), .B(n6874), .Z(n6873) );
  AND U7410 ( .A(n8440), .B(n8441), .Z(n6874) );
  XOR U7411 ( .A(n6877), .B(n6876), .Z(n6875) );
  AND U7412 ( .A(n8442), .B(n8443), .Z(n6876) );
  XOR U7413 ( .A(n6879), .B(n6878), .Z(n6877) );
  AND U7414 ( .A(n8444), .B(n8445), .Z(n6878) );
  XOR U7415 ( .A(n6881), .B(n6880), .Z(n6879) );
  AND U7416 ( .A(n8446), .B(n8447), .Z(n6880) );
  XOR U7417 ( .A(n6883), .B(n6882), .Z(n6881) );
  AND U7418 ( .A(n8448), .B(n8449), .Z(n6882) );
  XOR U7419 ( .A(n6885), .B(n6884), .Z(n6883) );
  AND U7420 ( .A(n8450), .B(n8451), .Z(n6884) );
  XOR U7421 ( .A(n6887), .B(n6886), .Z(n6885) );
  AND U7422 ( .A(n8452), .B(n8453), .Z(n6886) );
  XOR U7423 ( .A(n6889), .B(n6888), .Z(n6887) );
  AND U7424 ( .A(n8454), .B(n8455), .Z(n6888) );
  XOR U7425 ( .A(n6891), .B(n6890), .Z(n6889) );
  AND U7426 ( .A(n8456), .B(n8457), .Z(n6890) );
  XOR U7427 ( .A(n6893), .B(n6892), .Z(n6891) );
  AND U7428 ( .A(n8458), .B(n8459), .Z(n6892) );
  XOR U7429 ( .A(n6895), .B(n6894), .Z(n6893) );
  AND U7430 ( .A(n8460), .B(n8461), .Z(n6894) );
  XOR U7431 ( .A(n6897), .B(n6896), .Z(n6895) );
  AND U7432 ( .A(n8462), .B(n8463), .Z(n6896) );
  XOR U7433 ( .A(n6899), .B(n6898), .Z(n6897) );
  AND U7434 ( .A(n8464), .B(n8465), .Z(n6898) );
  XOR U7435 ( .A(n6901), .B(n6900), .Z(n6899) );
  AND U7436 ( .A(n8466), .B(n8467), .Z(n6900) );
  XOR U7437 ( .A(n6903), .B(n6902), .Z(n6901) );
  AND U7438 ( .A(n8468), .B(n8469), .Z(n6902) );
  XOR U7439 ( .A(n6905), .B(n6904), .Z(n6903) );
  AND U7440 ( .A(n8470), .B(n8471), .Z(n6904) );
  XOR U7441 ( .A(n6907), .B(n6906), .Z(n6905) );
  AND U7442 ( .A(n8472), .B(n8473), .Z(n6906) );
  XOR U7443 ( .A(n6909), .B(n6908), .Z(n6907) );
  AND U7444 ( .A(n8474), .B(n8475), .Z(n6908) );
  XOR U7445 ( .A(n6911), .B(n6910), .Z(n6909) );
  AND U7446 ( .A(n8476), .B(n8477), .Z(n6910) );
  XOR U7447 ( .A(n6913), .B(n6912), .Z(n6911) );
  AND U7448 ( .A(n8478), .B(n8479), .Z(n6912) );
  XOR U7449 ( .A(n6915), .B(n6914), .Z(n6913) );
  AND U7450 ( .A(n8480), .B(n8481), .Z(n6914) );
  XOR U7451 ( .A(n6917), .B(n6916), .Z(n6915) );
  AND U7452 ( .A(n8482), .B(n8483), .Z(n6916) );
  XOR U7453 ( .A(n6919), .B(n6918), .Z(n6917) );
  AND U7454 ( .A(n8484), .B(n8485), .Z(n6918) );
  XOR U7455 ( .A(n6921), .B(n6920), .Z(n6919) );
  AND U7456 ( .A(n8486), .B(n8487), .Z(n6920) );
  XOR U7457 ( .A(n6923), .B(n6922), .Z(n6921) );
  AND U7458 ( .A(n8488), .B(n8489), .Z(n6922) );
  XOR U7459 ( .A(n6925), .B(n6924), .Z(n6923) );
  AND U7460 ( .A(n8490), .B(n8491), .Z(n6924) );
  XOR U7461 ( .A(n6927), .B(n6926), .Z(n6925) );
  AND U7462 ( .A(n8492), .B(n8493), .Z(n6926) );
  XOR U7463 ( .A(n6929), .B(n6928), .Z(n6927) );
  AND U7464 ( .A(n8494), .B(n8495), .Z(n6928) );
  XOR U7465 ( .A(n6931), .B(n6930), .Z(n6929) );
  AND U7466 ( .A(n8496), .B(n8497), .Z(n6930) );
  XOR U7467 ( .A(n6933), .B(n6932), .Z(n6931) );
  AND U7468 ( .A(n8498), .B(n8499), .Z(n6932) );
  XOR U7469 ( .A(n6935), .B(n6934), .Z(n6933) );
  AND U7470 ( .A(n8500), .B(n8501), .Z(n6934) );
  XOR U7471 ( .A(n6937), .B(n6936), .Z(n6935) );
  AND U7472 ( .A(n8502), .B(n8503), .Z(n6936) );
  XOR U7473 ( .A(n6939), .B(n6938), .Z(n6937) );
  AND U7474 ( .A(n8504), .B(n8505), .Z(n6938) );
  XOR U7475 ( .A(n6941), .B(n6940), .Z(n6939) );
  AND U7476 ( .A(n8506), .B(n8507), .Z(n6940) );
  XOR U7477 ( .A(n6943), .B(n6942), .Z(n6941) );
  AND U7478 ( .A(n8508), .B(n8509), .Z(n6942) );
  XOR U7479 ( .A(n6945), .B(n6944), .Z(n6943) );
  AND U7480 ( .A(n8510), .B(n8511), .Z(n6944) );
  XOR U7481 ( .A(n6947), .B(n6946), .Z(n6945) );
  AND U7482 ( .A(n8512), .B(n8513), .Z(n6946) );
  XOR U7483 ( .A(n6949), .B(n6948), .Z(n6947) );
  AND U7484 ( .A(n8514), .B(n8515), .Z(n6948) );
  XOR U7485 ( .A(n6951), .B(n6950), .Z(n6949) );
  AND U7486 ( .A(n8516), .B(n8517), .Z(n6950) );
  XOR U7487 ( .A(n6953), .B(n6952), .Z(n6951) );
  AND U7488 ( .A(n8518), .B(n8519), .Z(n6952) );
  XOR U7489 ( .A(n6955), .B(n6954), .Z(n6953) );
  AND U7490 ( .A(n8520), .B(n8521), .Z(n6954) );
  XOR U7491 ( .A(n6957), .B(n6956), .Z(n6955) );
  AND U7492 ( .A(n8522), .B(n8523), .Z(n6956) );
  XOR U7493 ( .A(n6959), .B(n6958), .Z(n6957) );
  AND U7494 ( .A(n8524), .B(n8525), .Z(n6958) );
  XOR U7495 ( .A(n6987), .B(n6960), .Z(n6959) );
  AND U7496 ( .A(n8526), .B(n8527), .Z(n6960) );
  XOR U7497 ( .A(n6989), .B(n6988), .Z(n6987) );
  AND U7498 ( .A(n8528), .B(n8529), .Z(n6988) );
  XOR U7499 ( .A(n6968), .B(n6990), .Z(n6989) );
  AND U7500 ( .A(n8530), .B(n8531), .Z(n6990) );
  XOR U7501 ( .A(n6964), .B(n6969), .Z(n6968) );
  AND U7502 ( .A(n8532), .B(n8533), .Z(n6969) );
  XOR U7503 ( .A(n6966), .B(n6965), .Z(n6964) );
  AND U7504 ( .A(n8534), .B(n8535), .Z(n6965) );
  XNOR U7505 ( .A(n6976), .B(n6967), .Z(n6966) );
  AND U7506 ( .A(n8536), .B(n8537), .Z(n6967) );
  XOR U7507 ( .A(n6986), .B(n6975), .Z(n6976) );
  AND U7508 ( .A(n8538), .B(n8539), .Z(n6975) );
  XNOR U7509 ( .A(n8540), .B(n6981), .Z(n6986) );
  XOR U7510 ( .A(n6982), .B(n8541), .Z(n6981) );
  AND U7511 ( .A(n8542), .B(n8543), .Z(n8541) );
  XOR U7512 ( .A(n8544), .B(n8545), .Z(n6982) );
  NOR U7513 ( .A(n8546), .B(n8547), .Z(n8545) );
  AND U7514 ( .A(n8548), .B(n8549), .Z(n8547) );
  AND U7515 ( .A(n8550), .B(n8551), .Z(n8546) );
  XNOR U7516 ( .A(n8548), .B(n8549), .Z(n8544) );
  XNOR U7517 ( .A(n6973), .B(n6985), .Z(n8540) );
  AND U7518 ( .A(n8552), .B(n8553), .Z(n6985) );
  AND U7519 ( .A(n8554), .B(n8555), .Z(n6973) );
  XNOR U7520 ( .A(n8034), .B(n114), .Z(n8036) );
  XOR U7521 ( .A(n8031), .B(n8032), .Z(n114) );
  AND U7522 ( .A(n8556), .B(n8557), .Z(n8032) );
  XOR U7523 ( .A(n8028), .B(n8029), .Z(n8031) );
  AND U7524 ( .A(n8558), .B(n8559), .Z(n8029) );
  XOR U7525 ( .A(n8025), .B(n8026), .Z(n8028) );
  AND U7526 ( .A(n8560), .B(n8561), .Z(n8026) );
  XOR U7527 ( .A(n8022), .B(n8023), .Z(n8025) );
  AND U7528 ( .A(n8562), .B(n8563), .Z(n8023) );
  XOR U7529 ( .A(n8019), .B(n8020), .Z(n8022) );
  AND U7530 ( .A(n8564), .B(n8565), .Z(n8020) );
  XOR U7531 ( .A(n8016), .B(n8017), .Z(n8019) );
  AND U7532 ( .A(n8566), .B(n8567), .Z(n8017) );
  XOR U7533 ( .A(n8013), .B(n8014), .Z(n8016) );
  AND U7534 ( .A(n8568), .B(n8569), .Z(n8014) );
  XOR U7535 ( .A(n8010), .B(n8011), .Z(n8013) );
  AND U7536 ( .A(n8570), .B(n8571), .Z(n8011) );
  XOR U7537 ( .A(n8007), .B(n8008), .Z(n8010) );
  AND U7538 ( .A(n8572), .B(n8573), .Z(n8008) );
  XOR U7539 ( .A(n8004), .B(n8005), .Z(n8007) );
  AND U7540 ( .A(n8574), .B(n8575), .Z(n8005) );
  XOR U7541 ( .A(n8001), .B(n8002), .Z(n8004) );
  AND U7542 ( .A(n8576), .B(n8577), .Z(n8002) );
  XOR U7543 ( .A(n7998), .B(n7999), .Z(n8001) );
  AND U7544 ( .A(n8578), .B(n8579), .Z(n7999) );
  XOR U7545 ( .A(n7995), .B(n7996), .Z(n7998) );
  AND U7546 ( .A(n8580), .B(n8581), .Z(n7996) );
  XOR U7547 ( .A(n7992), .B(n7993), .Z(n7995) );
  AND U7548 ( .A(n8582), .B(n8583), .Z(n7993) );
  XOR U7549 ( .A(n7989), .B(n7990), .Z(n7992) );
  AND U7550 ( .A(n8584), .B(n8585), .Z(n7990) );
  XOR U7551 ( .A(n7986), .B(n7987), .Z(n7989) );
  AND U7552 ( .A(n8586), .B(n8587), .Z(n7987) );
  XOR U7553 ( .A(n7983), .B(n7984), .Z(n7986) );
  AND U7554 ( .A(n8588), .B(n8589), .Z(n7984) );
  XOR U7555 ( .A(n7980), .B(n7981), .Z(n7983) );
  AND U7556 ( .A(n8590), .B(n8591), .Z(n7981) );
  XOR U7557 ( .A(n7977), .B(n7978), .Z(n7980) );
  AND U7558 ( .A(n8592), .B(n8593), .Z(n7978) );
  XOR U7559 ( .A(n7974), .B(n7975), .Z(n7977) );
  AND U7560 ( .A(n8594), .B(n8595), .Z(n7975) );
  XOR U7561 ( .A(n7971), .B(n7972), .Z(n7974) );
  AND U7562 ( .A(n8596), .B(n8597), .Z(n7972) );
  XOR U7563 ( .A(n7968), .B(n7969), .Z(n7971) );
  AND U7564 ( .A(n8598), .B(n8599), .Z(n7969) );
  XOR U7565 ( .A(n7965), .B(n7966), .Z(n7968) );
  AND U7566 ( .A(n8600), .B(n8601), .Z(n7966) );
  XOR U7567 ( .A(n7962), .B(n7963), .Z(n7965) );
  AND U7568 ( .A(n8602), .B(n8603), .Z(n7963) );
  XOR U7569 ( .A(n7959), .B(n7960), .Z(n7962) );
  AND U7570 ( .A(n8604), .B(n8605), .Z(n7960) );
  XOR U7571 ( .A(n7956), .B(n7957), .Z(n7959) );
  AND U7572 ( .A(n8606), .B(n8607), .Z(n7957) );
  XOR U7573 ( .A(n7953), .B(n7954), .Z(n7956) );
  AND U7574 ( .A(n8608), .B(n8609), .Z(n7954) );
  XOR U7575 ( .A(n7950), .B(n7951), .Z(n7953) );
  AND U7576 ( .A(n8610), .B(n8611), .Z(n7951) );
  XOR U7577 ( .A(n7947), .B(n7948), .Z(n7950) );
  AND U7578 ( .A(n8612), .B(n8613), .Z(n7948) );
  XOR U7579 ( .A(n7944), .B(n7945), .Z(n7947) );
  AND U7580 ( .A(n8614), .B(n8615), .Z(n7945) );
  XOR U7581 ( .A(n7941), .B(n7942), .Z(n7944) );
  AND U7582 ( .A(n8616), .B(n8617), .Z(n7942) );
  XOR U7583 ( .A(n7938), .B(n7939), .Z(n7941) );
  AND U7584 ( .A(n8618), .B(n8619), .Z(n7939) );
  XOR U7585 ( .A(n7935), .B(n7936), .Z(n7938) );
  AND U7586 ( .A(n8620), .B(n8621), .Z(n7936) );
  XOR U7587 ( .A(n7932), .B(n7933), .Z(n7935) );
  AND U7588 ( .A(n8622), .B(n8623), .Z(n7933) );
  XOR U7589 ( .A(n7929), .B(n7930), .Z(n7932) );
  AND U7590 ( .A(n8624), .B(n8625), .Z(n7930) );
  XOR U7591 ( .A(n7926), .B(n7927), .Z(n7929) );
  AND U7592 ( .A(n8626), .B(n8627), .Z(n7927) );
  XOR U7593 ( .A(n7923), .B(n7924), .Z(n7926) );
  AND U7594 ( .A(n8628), .B(n8629), .Z(n7924) );
  XOR U7595 ( .A(n7920), .B(n7921), .Z(n7923) );
  AND U7596 ( .A(n8630), .B(n8631), .Z(n7921) );
  XOR U7597 ( .A(n7917), .B(n7918), .Z(n7920) );
  AND U7598 ( .A(n8632), .B(n8633), .Z(n7918) );
  XOR U7599 ( .A(n7914), .B(n7915), .Z(n7917) );
  AND U7600 ( .A(n8634), .B(n8635), .Z(n7915) );
  XOR U7601 ( .A(n7911), .B(n7912), .Z(n7914) );
  AND U7602 ( .A(n8636), .B(n8637), .Z(n7912) );
  XOR U7603 ( .A(n7908), .B(n7909), .Z(n7911) );
  AND U7604 ( .A(n8638), .B(n8639), .Z(n7909) );
  XOR U7605 ( .A(n7905), .B(n7906), .Z(n7908) );
  AND U7606 ( .A(n8640), .B(n8641), .Z(n7906) );
  XOR U7607 ( .A(n7902), .B(n7903), .Z(n7905) );
  AND U7608 ( .A(n8642), .B(n8643), .Z(n7903) );
  XOR U7609 ( .A(n7899), .B(n7900), .Z(n7902) );
  AND U7610 ( .A(n8644), .B(n8645), .Z(n7900) );
  XOR U7611 ( .A(n7896), .B(n7897), .Z(n7899) );
  AND U7612 ( .A(n8646), .B(n8647), .Z(n7897) );
  XOR U7613 ( .A(n7893), .B(n7894), .Z(n7896) );
  AND U7614 ( .A(n8648), .B(n8649), .Z(n7894) );
  XOR U7615 ( .A(n7890), .B(n7891), .Z(n7893) );
  AND U7616 ( .A(n8650), .B(n8651), .Z(n7891) );
  XOR U7617 ( .A(n7887), .B(n7888), .Z(n7890) );
  AND U7618 ( .A(n8652), .B(n8653), .Z(n7888) );
  XOR U7619 ( .A(n7884), .B(n7885), .Z(n7887) );
  AND U7620 ( .A(n8654), .B(n8655), .Z(n7885) );
  XOR U7621 ( .A(n7881), .B(n7882), .Z(n7884) );
  AND U7622 ( .A(n8656), .B(n8657), .Z(n7882) );
  XOR U7623 ( .A(n7878), .B(n7879), .Z(n7881) );
  AND U7624 ( .A(n8658), .B(n8659), .Z(n7879) );
  XOR U7625 ( .A(n7875), .B(n7876), .Z(n7878) );
  AND U7626 ( .A(n8660), .B(n8661), .Z(n7876) );
  XOR U7627 ( .A(n7872), .B(n7873), .Z(n7875) );
  AND U7628 ( .A(n8662), .B(n8663), .Z(n7873) );
  XOR U7629 ( .A(n7869), .B(n7870), .Z(n7872) );
  AND U7630 ( .A(n8664), .B(n8665), .Z(n7870) );
  XOR U7631 ( .A(n7866), .B(n7867), .Z(n7869) );
  AND U7632 ( .A(n8666), .B(n8667), .Z(n7867) );
  XOR U7633 ( .A(n7863), .B(n7864), .Z(n7866) );
  AND U7634 ( .A(n8668), .B(n8669), .Z(n7864) );
  XOR U7635 ( .A(n7860), .B(n7861), .Z(n7863) );
  AND U7636 ( .A(n8670), .B(n8671), .Z(n7861) );
  XOR U7637 ( .A(n7857), .B(n7858), .Z(n7860) );
  AND U7638 ( .A(n8672), .B(n8673), .Z(n7858) );
  XOR U7639 ( .A(n7854), .B(n7855), .Z(n7857) );
  AND U7640 ( .A(n8674), .B(n8675), .Z(n7855) );
  XOR U7641 ( .A(n7851), .B(n7852), .Z(n7854) );
  AND U7642 ( .A(n8676), .B(n8677), .Z(n7852) );
  XOR U7643 ( .A(n7848), .B(n7849), .Z(n7851) );
  AND U7644 ( .A(n8678), .B(n8679), .Z(n7849) );
  XOR U7645 ( .A(n7845), .B(n7846), .Z(n7848) );
  AND U7646 ( .A(n8680), .B(n8681), .Z(n7846) );
  XOR U7647 ( .A(n7842), .B(n7843), .Z(n7845) );
  AND U7648 ( .A(n8682), .B(n8683), .Z(n7843) );
  XOR U7649 ( .A(n7839), .B(n7840), .Z(n7842) );
  AND U7650 ( .A(n8684), .B(n8685), .Z(n7840) );
  XOR U7651 ( .A(n7836), .B(n7837), .Z(n7839) );
  AND U7652 ( .A(n8686), .B(n8687), .Z(n7837) );
  XOR U7653 ( .A(n7833), .B(n7834), .Z(n7836) );
  AND U7654 ( .A(n8688), .B(n8689), .Z(n7834) );
  XOR U7655 ( .A(n7830), .B(n7831), .Z(n7833) );
  AND U7656 ( .A(n8690), .B(n8691), .Z(n7831) );
  XOR U7657 ( .A(n7827), .B(n7828), .Z(n7830) );
  AND U7658 ( .A(n8692), .B(n8693), .Z(n7828) );
  XOR U7659 ( .A(n7824), .B(n7825), .Z(n7827) );
  AND U7660 ( .A(n8694), .B(n8695), .Z(n7825) );
  XOR U7661 ( .A(n7821), .B(n7822), .Z(n7824) );
  AND U7662 ( .A(n8696), .B(n8697), .Z(n7822) );
  XOR U7663 ( .A(n7818), .B(n7819), .Z(n7821) );
  AND U7664 ( .A(n8698), .B(n8699), .Z(n7819) );
  XOR U7665 ( .A(n7815), .B(n7816), .Z(n7818) );
  AND U7666 ( .A(n8700), .B(n8701), .Z(n7816) );
  XOR U7667 ( .A(n7812), .B(n7813), .Z(n7815) );
  AND U7668 ( .A(n8702), .B(n8703), .Z(n7813) );
  XOR U7669 ( .A(n7809), .B(n7810), .Z(n7812) );
  AND U7670 ( .A(n8704), .B(n8705), .Z(n7810) );
  XOR U7671 ( .A(n7806), .B(n7807), .Z(n7809) );
  AND U7672 ( .A(n8706), .B(n8707), .Z(n7807) );
  XOR U7673 ( .A(n7803), .B(n7804), .Z(n7806) );
  AND U7674 ( .A(n8708), .B(n8709), .Z(n7804) );
  XOR U7675 ( .A(n7800), .B(n7801), .Z(n7803) );
  AND U7676 ( .A(n8710), .B(n8711), .Z(n7801) );
  XOR U7677 ( .A(n7797), .B(n7798), .Z(n7800) );
  AND U7678 ( .A(n8712), .B(n8713), .Z(n7798) );
  XOR U7679 ( .A(n7794), .B(n7795), .Z(n7797) );
  AND U7680 ( .A(n8714), .B(n8715), .Z(n7795) );
  XOR U7681 ( .A(n7791), .B(n7792), .Z(n7794) );
  AND U7682 ( .A(n8716), .B(n8717), .Z(n7792) );
  XOR U7683 ( .A(n7788), .B(n7789), .Z(n7791) );
  AND U7684 ( .A(n8718), .B(n8719), .Z(n7789) );
  XOR U7685 ( .A(n7785), .B(n7786), .Z(n7788) );
  AND U7686 ( .A(n8720), .B(n8721), .Z(n7786) );
  XOR U7687 ( .A(n7782), .B(n7783), .Z(n7785) );
  AND U7688 ( .A(n8722), .B(n8723), .Z(n7783) );
  XOR U7689 ( .A(n7779), .B(n7780), .Z(n7782) );
  AND U7690 ( .A(n8724), .B(n8725), .Z(n7780) );
  XOR U7691 ( .A(n7776), .B(n7777), .Z(n7779) );
  AND U7692 ( .A(n8726), .B(n8727), .Z(n7777) );
  XOR U7693 ( .A(n7773), .B(n7774), .Z(n7776) );
  AND U7694 ( .A(n8728), .B(n8729), .Z(n7774) );
  XOR U7695 ( .A(n7770), .B(n7771), .Z(n7773) );
  AND U7696 ( .A(n8730), .B(n8731), .Z(n7771) );
  XOR U7697 ( .A(n7767), .B(n7768), .Z(n7770) );
  AND U7698 ( .A(n8732), .B(n8733), .Z(n7768) );
  XOR U7699 ( .A(n7764), .B(n7765), .Z(n7767) );
  AND U7700 ( .A(n8734), .B(n8735), .Z(n7765) );
  XOR U7701 ( .A(n7761), .B(n7762), .Z(n7764) );
  AND U7702 ( .A(n8736), .B(n8737), .Z(n7762) );
  XOR U7703 ( .A(n7758), .B(n7759), .Z(n7761) );
  AND U7704 ( .A(n8738), .B(n8739), .Z(n7759) );
  XOR U7705 ( .A(n7755), .B(n7756), .Z(n7758) );
  AND U7706 ( .A(n8740), .B(n8741), .Z(n7756) );
  XOR U7707 ( .A(n7752), .B(n7753), .Z(n7755) );
  AND U7708 ( .A(n8742), .B(n8743), .Z(n7753) );
  XOR U7709 ( .A(n7749), .B(n7750), .Z(n7752) );
  AND U7710 ( .A(n8744), .B(n8745), .Z(n7750) );
  XOR U7711 ( .A(n7746), .B(n7747), .Z(n7749) );
  AND U7712 ( .A(n8746), .B(n8747), .Z(n7747) );
  XOR U7713 ( .A(n7743), .B(n7744), .Z(n7746) );
  AND U7714 ( .A(n8748), .B(n8749), .Z(n7744) );
  XOR U7715 ( .A(n7740), .B(n7741), .Z(n7743) );
  AND U7716 ( .A(n8750), .B(n8751), .Z(n7741) );
  XOR U7717 ( .A(n7737), .B(n7738), .Z(n7740) );
  AND U7718 ( .A(n8752), .B(n8753), .Z(n7738) );
  XOR U7719 ( .A(n7734), .B(n7735), .Z(n7737) );
  AND U7720 ( .A(n8754), .B(n8755), .Z(n7735) );
  XOR U7721 ( .A(n7731), .B(n7732), .Z(n7734) );
  AND U7722 ( .A(n8756), .B(n8757), .Z(n7732) );
  XOR U7723 ( .A(n7728), .B(n7729), .Z(n7731) );
  AND U7724 ( .A(n8758), .B(n8759), .Z(n7729) );
  XOR U7725 ( .A(n7725), .B(n7726), .Z(n7728) );
  AND U7726 ( .A(n8760), .B(n8761), .Z(n7726) );
  XOR U7727 ( .A(n7722), .B(n7723), .Z(n7725) );
  AND U7728 ( .A(n8762), .B(n8763), .Z(n7723) );
  XOR U7729 ( .A(n7719), .B(n7720), .Z(n7722) );
  AND U7730 ( .A(n8764), .B(n8765), .Z(n7720) );
  XOR U7731 ( .A(n7716), .B(n7717), .Z(n7719) );
  AND U7732 ( .A(n8766), .B(n8767), .Z(n7717) );
  XOR U7733 ( .A(n7713), .B(n7714), .Z(n7716) );
  AND U7734 ( .A(n8768), .B(n8769), .Z(n7714) );
  XOR U7735 ( .A(n7710), .B(n7711), .Z(n7713) );
  AND U7736 ( .A(n8770), .B(n8771), .Z(n7711) );
  XOR U7737 ( .A(n7707), .B(n7708), .Z(n7710) );
  AND U7738 ( .A(n8772), .B(n8773), .Z(n7708) );
  XOR U7739 ( .A(n7704), .B(n7705), .Z(n7707) );
  AND U7740 ( .A(n8774), .B(n8775), .Z(n7705) );
  XOR U7741 ( .A(n7701), .B(n7702), .Z(n7704) );
  AND U7742 ( .A(n8776), .B(n8777), .Z(n7702) );
  XOR U7743 ( .A(n7698), .B(n7699), .Z(n7701) );
  AND U7744 ( .A(n8778), .B(n8779), .Z(n7699) );
  XOR U7745 ( .A(n7695), .B(n7696), .Z(n7698) );
  AND U7746 ( .A(n8780), .B(n8781), .Z(n7696) );
  XOR U7747 ( .A(n7692), .B(n7693), .Z(n7695) );
  AND U7748 ( .A(n8782), .B(n8783), .Z(n7693) );
  XOR U7749 ( .A(n7689), .B(n7690), .Z(n7692) );
  AND U7750 ( .A(n8784), .B(n8785), .Z(n7690) );
  XOR U7751 ( .A(n7686), .B(n7687), .Z(n7689) );
  AND U7752 ( .A(n8786), .B(n8787), .Z(n7687) );
  XOR U7753 ( .A(n7683), .B(n7684), .Z(n7686) );
  AND U7754 ( .A(n8788), .B(n8789), .Z(n7684) );
  XOR U7755 ( .A(n7680), .B(n7681), .Z(n7683) );
  AND U7756 ( .A(n8790), .B(n8791), .Z(n7681) );
  XOR U7757 ( .A(n7677), .B(n7678), .Z(n7680) );
  AND U7758 ( .A(n8792), .B(n8793), .Z(n7678) );
  XOR U7759 ( .A(n7674), .B(n7675), .Z(n7677) );
  AND U7760 ( .A(n8794), .B(n8795), .Z(n7675) );
  XOR U7761 ( .A(n7671), .B(n7672), .Z(n7674) );
  AND U7762 ( .A(n8796), .B(n8797), .Z(n7672) );
  XOR U7763 ( .A(n7668), .B(n7669), .Z(n7671) );
  AND U7764 ( .A(n8798), .B(n8799), .Z(n7669) );
  XOR U7765 ( .A(n7665), .B(n7666), .Z(n7668) );
  AND U7766 ( .A(n8800), .B(n8801), .Z(n7666) );
  XOR U7767 ( .A(n7662), .B(n7663), .Z(n7665) );
  AND U7768 ( .A(n8802), .B(n8803), .Z(n7663) );
  XOR U7769 ( .A(n7659), .B(n7660), .Z(n7662) );
  AND U7770 ( .A(n8804), .B(n8805), .Z(n7660) );
  XOR U7771 ( .A(n7656), .B(n7657), .Z(n7659) );
  AND U7772 ( .A(n8806), .B(n8807), .Z(n7657) );
  XOR U7773 ( .A(n7653), .B(n7654), .Z(n7656) );
  AND U7774 ( .A(n8808), .B(n8809), .Z(n7654) );
  XOR U7775 ( .A(n7650), .B(n7651), .Z(n7653) );
  AND U7776 ( .A(n8810), .B(n8811), .Z(n7651) );
  XNOR U7777 ( .A(n7647), .B(n7648), .Z(n7650) );
  AND U7778 ( .A(n8812), .B(n8813), .Z(n7648) );
  XOR U7779 ( .A(n8814), .B(n7645), .Z(n7647) );
  IV U7780 ( .A(n8815), .Z(n7645) );
  AND U7781 ( .A(n8816), .B(n8817), .Z(n8815) );
  IV U7782 ( .A(n7644), .Z(n8814) );
  XOR U7783 ( .A(n7385), .B(n7641), .Z(n7644) );
  AND U7784 ( .A(n8818), .B(n8819), .Z(n7641) );
  XOR U7785 ( .A(n7387), .B(n7386), .Z(n7385) );
  AND U7786 ( .A(n8820), .B(n8821), .Z(n7386) );
  XOR U7787 ( .A(n7389), .B(n7388), .Z(n7387) );
  AND U7788 ( .A(n8822), .B(n8823), .Z(n7388) );
  XOR U7789 ( .A(n7391), .B(n7390), .Z(n7389) );
  AND U7790 ( .A(n8824), .B(n8825), .Z(n7390) );
  XOR U7791 ( .A(n7393), .B(n7392), .Z(n7391) );
  AND U7792 ( .A(n8826), .B(n8827), .Z(n7392) );
  XOR U7793 ( .A(n7395), .B(n7394), .Z(n7393) );
  AND U7794 ( .A(n8828), .B(n8829), .Z(n7394) );
  XOR U7795 ( .A(n7397), .B(n7396), .Z(n7395) );
  AND U7796 ( .A(n8830), .B(n8831), .Z(n7396) );
  XOR U7797 ( .A(n7399), .B(n7398), .Z(n7397) );
  AND U7798 ( .A(n8832), .B(n8833), .Z(n7398) );
  XOR U7799 ( .A(n7401), .B(n7400), .Z(n7399) );
  AND U7800 ( .A(n8834), .B(n8835), .Z(n7400) );
  XOR U7801 ( .A(n7403), .B(n7402), .Z(n7401) );
  AND U7802 ( .A(n8836), .B(n8837), .Z(n7402) );
  XOR U7803 ( .A(n7405), .B(n7404), .Z(n7403) );
  AND U7804 ( .A(n8838), .B(n8839), .Z(n7404) );
  XOR U7805 ( .A(n7407), .B(n7406), .Z(n7405) );
  AND U7806 ( .A(n8840), .B(n8841), .Z(n7406) );
  XOR U7807 ( .A(n7409), .B(n7408), .Z(n7407) );
  AND U7808 ( .A(n8842), .B(n8843), .Z(n7408) );
  XOR U7809 ( .A(n7411), .B(n7410), .Z(n7409) );
  AND U7810 ( .A(n8844), .B(n8845), .Z(n7410) );
  XOR U7811 ( .A(n7413), .B(n7412), .Z(n7411) );
  AND U7812 ( .A(n8846), .B(n8847), .Z(n7412) );
  XOR U7813 ( .A(n7415), .B(n7414), .Z(n7413) );
  AND U7814 ( .A(n8848), .B(n8849), .Z(n7414) );
  XOR U7815 ( .A(n7417), .B(n7416), .Z(n7415) );
  AND U7816 ( .A(n8850), .B(n8851), .Z(n7416) );
  XOR U7817 ( .A(n7419), .B(n7418), .Z(n7417) );
  AND U7818 ( .A(n8852), .B(n8853), .Z(n7418) );
  XOR U7819 ( .A(n7421), .B(n7420), .Z(n7419) );
  AND U7820 ( .A(n8854), .B(n8855), .Z(n7420) );
  XOR U7821 ( .A(n7423), .B(n7422), .Z(n7421) );
  AND U7822 ( .A(n8856), .B(n8857), .Z(n7422) );
  XOR U7823 ( .A(n7425), .B(n7424), .Z(n7423) );
  AND U7824 ( .A(n8858), .B(n8859), .Z(n7424) );
  XOR U7825 ( .A(n7427), .B(n7426), .Z(n7425) );
  AND U7826 ( .A(n8860), .B(n8861), .Z(n7426) );
  XOR U7827 ( .A(n7429), .B(n7428), .Z(n7427) );
  AND U7828 ( .A(n8862), .B(n8863), .Z(n7428) );
  XOR U7829 ( .A(n7431), .B(n7430), .Z(n7429) );
  AND U7830 ( .A(n8864), .B(n8865), .Z(n7430) );
  XOR U7831 ( .A(n7433), .B(n7432), .Z(n7431) );
  AND U7832 ( .A(n8866), .B(n8867), .Z(n7432) );
  XOR U7833 ( .A(n7435), .B(n7434), .Z(n7433) );
  AND U7834 ( .A(n8868), .B(n8869), .Z(n7434) );
  XOR U7835 ( .A(n7437), .B(n7436), .Z(n7435) );
  AND U7836 ( .A(n8870), .B(n8871), .Z(n7436) );
  XOR U7837 ( .A(n7439), .B(n7438), .Z(n7437) );
  AND U7838 ( .A(n8872), .B(n8873), .Z(n7438) );
  XOR U7839 ( .A(n7441), .B(n7440), .Z(n7439) );
  AND U7840 ( .A(n8874), .B(n8875), .Z(n7440) );
  XOR U7841 ( .A(n7443), .B(n7442), .Z(n7441) );
  AND U7842 ( .A(n8876), .B(n8877), .Z(n7442) );
  XOR U7843 ( .A(n7445), .B(n7444), .Z(n7443) );
  AND U7844 ( .A(n8878), .B(n8879), .Z(n7444) );
  XOR U7845 ( .A(n7447), .B(n7446), .Z(n7445) );
  AND U7846 ( .A(n8880), .B(n8881), .Z(n7446) );
  XOR U7847 ( .A(n7449), .B(n7448), .Z(n7447) );
  AND U7848 ( .A(n8882), .B(n8883), .Z(n7448) );
  XOR U7849 ( .A(n7451), .B(n7450), .Z(n7449) );
  AND U7850 ( .A(n8884), .B(n8885), .Z(n7450) );
  XOR U7851 ( .A(n7453), .B(n7452), .Z(n7451) );
  AND U7852 ( .A(n8886), .B(n8887), .Z(n7452) );
  XOR U7853 ( .A(n7455), .B(n7454), .Z(n7453) );
  AND U7854 ( .A(n8888), .B(n8889), .Z(n7454) );
  XOR U7855 ( .A(n7457), .B(n7456), .Z(n7455) );
  AND U7856 ( .A(n8890), .B(n8891), .Z(n7456) );
  XOR U7857 ( .A(n7459), .B(n7458), .Z(n7457) );
  AND U7858 ( .A(n8892), .B(n8893), .Z(n7458) );
  XOR U7859 ( .A(n7461), .B(n7460), .Z(n7459) );
  AND U7860 ( .A(n8894), .B(n8895), .Z(n7460) );
  XOR U7861 ( .A(n7463), .B(n7462), .Z(n7461) );
  AND U7862 ( .A(n8896), .B(n8897), .Z(n7462) );
  XOR U7863 ( .A(n7465), .B(n7464), .Z(n7463) );
  AND U7864 ( .A(n8898), .B(n8899), .Z(n7464) );
  XOR U7865 ( .A(n7467), .B(n7466), .Z(n7465) );
  AND U7866 ( .A(n8900), .B(n8901), .Z(n7466) );
  XOR U7867 ( .A(n7469), .B(n7468), .Z(n7467) );
  AND U7868 ( .A(n8902), .B(n8903), .Z(n7468) );
  XOR U7869 ( .A(n7471), .B(n7470), .Z(n7469) );
  AND U7870 ( .A(n8904), .B(n8905), .Z(n7470) );
  XOR U7871 ( .A(n7473), .B(n7472), .Z(n7471) );
  AND U7872 ( .A(n8906), .B(n8907), .Z(n7472) );
  XOR U7873 ( .A(n7475), .B(n7474), .Z(n7473) );
  AND U7874 ( .A(n8908), .B(n8909), .Z(n7474) );
  XOR U7875 ( .A(n7477), .B(n7476), .Z(n7475) );
  AND U7876 ( .A(n8910), .B(n8911), .Z(n7476) );
  XOR U7877 ( .A(n7479), .B(n7478), .Z(n7477) );
  AND U7878 ( .A(n8912), .B(n8913), .Z(n7478) );
  XOR U7879 ( .A(n7481), .B(n7480), .Z(n7479) );
  AND U7880 ( .A(n8914), .B(n8915), .Z(n7480) );
  XOR U7881 ( .A(n7483), .B(n7482), .Z(n7481) );
  AND U7882 ( .A(n8916), .B(n8917), .Z(n7482) );
  XOR U7883 ( .A(n7485), .B(n7484), .Z(n7483) );
  AND U7884 ( .A(n8918), .B(n8919), .Z(n7484) );
  XOR U7885 ( .A(n7487), .B(n7486), .Z(n7485) );
  AND U7886 ( .A(n8920), .B(n8921), .Z(n7486) );
  XOR U7887 ( .A(n7489), .B(n7488), .Z(n7487) );
  AND U7888 ( .A(n8922), .B(n8923), .Z(n7488) );
  XOR U7889 ( .A(n7491), .B(n7490), .Z(n7489) );
  AND U7890 ( .A(n8924), .B(n8925), .Z(n7490) );
  XOR U7891 ( .A(n7493), .B(n7492), .Z(n7491) );
  AND U7892 ( .A(n8926), .B(n8927), .Z(n7492) );
  XOR U7893 ( .A(n7495), .B(n7494), .Z(n7493) );
  AND U7894 ( .A(n8928), .B(n8929), .Z(n7494) );
  XOR U7895 ( .A(n7497), .B(n7496), .Z(n7495) );
  AND U7896 ( .A(n8930), .B(n8931), .Z(n7496) );
  XOR U7897 ( .A(n7499), .B(n7498), .Z(n7497) );
  AND U7898 ( .A(n8932), .B(n8933), .Z(n7498) );
  XOR U7899 ( .A(n7501), .B(n7500), .Z(n7499) );
  AND U7900 ( .A(n8934), .B(n8935), .Z(n7500) );
  XOR U7901 ( .A(n7503), .B(n7502), .Z(n7501) );
  AND U7902 ( .A(n8936), .B(n8937), .Z(n7502) );
  XOR U7903 ( .A(n7505), .B(n7504), .Z(n7503) );
  AND U7904 ( .A(n8938), .B(n8939), .Z(n7504) );
  XOR U7905 ( .A(n7507), .B(n7506), .Z(n7505) );
  AND U7906 ( .A(n8940), .B(n8941), .Z(n7506) );
  XOR U7907 ( .A(n7509), .B(n7508), .Z(n7507) );
  AND U7908 ( .A(n8942), .B(n8943), .Z(n7508) );
  XOR U7909 ( .A(n7511), .B(n7510), .Z(n7509) );
  AND U7910 ( .A(n8944), .B(n8945), .Z(n7510) );
  XOR U7911 ( .A(n7513), .B(n7512), .Z(n7511) );
  AND U7912 ( .A(n8946), .B(n8947), .Z(n7512) );
  XOR U7913 ( .A(n7515), .B(n7514), .Z(n7513) );
  AND U7914 ( .A(n8948), .B(n8949), .Z(n7514) );
  XOR U7915 ( .A(n7517), .B(n7516), .Z(n7515) );
  AND U7916 ( .A(n8950), .B(n8951), .Z(n7516) );
  XOR U7917 ( .A(n7519), .B(n7518), .Z(n7517) );
  AND U7918 ( .A(n8952), .B(n8953), .Z(n7518) );
  XOR U7919 ( .A(n7521), .B(n7520), .Z(n7519) );
  AND U7920 ( .A(n8954), .B(n8955), .Z(n7520) );
  XOR U7921 ( .A(n7523), .B(n7522), .Z(n7521) );
  AND U7922 ( .A(n8956), .B(n8957), .Z(n7522) );
  XOR U7923 ( .A(n7525), .B(n7524), .Z(n7523) );
  AND U7924 ( .A(n8958), .B(n8959), .Z(n7524) );
  XOR U7925 ( .A(n7527), .B(n7526), .Z(n7525) );
  AND U7926 ( .A(n8960), .B(n8961), .Z(n7526) );
  XOR U7927 ( .A(n7529), .B(n7528), .Z(n7527) );
  AND U7928 ( .A(n8962), .B(n8963), .Z(n7528) );
  XOR U7929 ( .A(n7531), .B(n7530), .Z(n7529) );
  AND U7930 ( .A(n8964), .B(n8965), .Z(n7530) );
  XOR U7931 ( .A(n7533), .B(n7532), .Z(n7531) );
  AND U7932 ( .A(n8966), .B(n8967), .Z(n7532) );
  XOR U7933 ( .A(n7535), .B(n7534), .Z(n7533) );
  AND U7934 ( .A(n8968), .B(n8969), .Z(n7534) );
  XOR U7935 ( .A(n7537), .B(n7536), .Z(n7535) );
  AND U7936 ( .A(n8970), .B(n8971), .Z(n7536) );
  XOR U7937 ( .A(n7539), .B(n7538), .Z(n7537) );
  AND U7938 ( .A(n8972), .B(n8973), .Z(n7538) );
  XOR U7939 ( .A(n7541), .B(n7540), .Z(n7539) );
  AND U7940 ( .A(n8974), .B(n8975), .Z(n7540) );
  XOR U7941 ( .A(n7543), .B(n7542), .Z(n7541) );
  AND U7942 ( .A(n8976), .B(n8977), .Z(n7542) );
  XOR U7943 ( .A(n7545), .B(n7544), .Z(n7543) );
  AND U7944 ( .A(n8978), .B(n8979), .Z(n7544) );
  XOR U7945 ( .A(n7547), .B(n7546), .Z(n7545) );
  AND U7946 ( .A(n8980), .B(n8981), .Z(n7546) );
  XOR U7947 ( .A(n7549), .B(n7548), .Z(n7547) );
  AND U7948 ( .A(n8982), .B(n8983), .Z(n7548) );
  XOR U7949 ( .A(n7551), .B(n7550), .Z(n7549) );
  AND U7950 ( .A(n8984), .B(n8985), .Z(n7550) );
  XOR U7951 ( .A(n7553), .B(n7552), .Z(n7551) );
  AND U7952 ( .A(n8986), .B(n8987), .Z(n7552) );
  XOR U7953 ( .A(n7555), .B(n7554), .Z(n7553) );
  AND U7954 ( .A(n8988), .B(n8989), .Z(n7554) );
  XOR U7955 ( .A(n7557), .B(n7556), .Z(n7555) );
  AND U7956 ( .A(n8990), .B(n8991), .Z(n7556) );
  XOR U7957 ( .A(n7559), .B(n7558), .Z(n7557) );
  AND U7958 ( .A(n8992), .B(n8993), .Z(n7558) );
  XOR U7959 ( .A(n7561), .B(n7560), .Z(n7559) );
  AND U7960 ( .A(n8994), .B(n8995), .Z(n7560) );
  XOR U7961 ( .A(n7563), .B(n7562), .Z(n7561) );
  AND U7962 ( .A(n8996), .B(n8997), .Z(n7562) );
  XOR U7963 ( .A(n7565), .B(n7564), .Z(n7563) );
  AND U7964 ( .A(n8998), .B(n8999), .Z(n7564) );
  XOR U7965 ( .A(n7567), .B(n7566), .Z(n7565) );
  AND U7966 ( .A(n9000), .B(n9001), .Z(n7566) );
  XOR U7967 ( .A(n7569), .B(n7568), .Z(n7567) );
  AND U7968 ( .A(n9002), .B(n9003), .Z(n7568) );
  XOR U7969 ( .A(n7571), .B(n7570), .Z(n7569) );
  AND U7970 ( .A(n9004), .B(n9005), .Z(n7570) );
  XOR U7971 ( .A(n7573), .B(n7572), .Z(n7571) );
  AND U7972 ( .A(n9006), .B(n9007), .Z(n7572) );
  XOR U7973 ( .A(n7575), .B(n7574), .Z(n7573) );
  AND U7974 ( .A(n9008), .B(n9009), .Z(n7574) );
  XOR U7975 ( .A(n7577), .B(n7576), .Z(n7575) );
  AND U7976 ( .A(n9010), .B(n9011), .Z(n7576) );
  XOR U7977 ( .A(n7579), .B(n7578), .Z(n7577) );
  AND U7978 ( .A(n9012), .B(n9013), .Z(n7578) );
  XOR U7979 ( .A(n7581), .B(n7580), .Z(n7579) );
  AND U7980 ( .A(n9014), .B(n9015), .Z(n7580) );
  XOR U7981 ( .A(n7583), .B(n7582), .Z(n7581) );
  AND U7982 ( .A(n9016), .B(n9017), .Z(n7582) );
  XOR U7983 ( .A(n7585), .B(n7584), .Z(n7583) );
  AND U7984 ( .A(n9018), .B(n9019), .Z(n7584) );
  XOR U7985 ( .A(n7587), .B(n7586), .Z(n7585) );
  AND U7986 ( .A(n9020), .B(n9021), .Z(n7586) );
  XOR U7987 ( .A(n7589), .B(n7588), .Z(n7587) );
  AND U7988 ( .A(n9022), .B(n9023), .Z(n7588) );
  XOR U7989 ( .A(n7591), .B(n7590), .Z(n7589) );
  AND U7990 ( .A(n9024), .B(n9025), .Z(n7590) );
  XOR U7991 ( .A(n7593), .B(n7592), .Z(n7591) );
  AND U7992 ( .A(n9026), .B(n9027), .Z(n7592) );
  XOR U7993 ( .A(n7595), .B(n7594), .Z(n7593) );
  AND U7994 ( .A(n9028), .B(n9029), .Z(n7594) );
  XOR U7995 ( .A(n7597), .B(n7596), .Z(n7595) );
  AND U7996 ( .A(n9030), .B(n9031), .Z(n7596) );
  XOR U7997 ( .A(n7599), .B(n7598), .Z(n7597) );
  AND U7998 ( .A(n9032), .B(n9033), .Z(n7598) );
  XOR U7999 ( .A(n7601), .B(n7600), .Z(n7599) );
  AND U8000 ( .A(n9034), .B(n9035), .Z(n7600) );
  XOR U8001 ( .A(n7603), .B(n7602), .Z(n7601) );
  AND U8002 ( .A(n9036), .B(n9037), .Z(n7602) );
  XOR U8003 ( .A(n7605), .B(n7604), .Z(n7603) );
  AND U8004 ( .A(n9038), .B(n9039), .Z(n7604) );
  XOR U8005 ( .A(n7607), .B(n7606), .Z(n7605) );
  AND U8006 ( .A(n9040), .B(n9041), .Z(n7606) );
  XOR U8007 ( .A(n7609), .B(n7608), .Z(n7607) );
  AND U8008 ( .A(n9042), .B(n9043), .Z(n7608) );
  XOR U8009 ( .A(n7637), .B(n7610), .Z(n7609) );
  AND U8010 ( .A(n9044), .B(n9045), .Z(n7610) );
  XOR U8011 ( .A(n7639), .B(n7638), .Z(n7637) );
  AND U8012 ( .A(n9046), .B(n9047), .Z(n7638) );
  XOR U8013 ( .A(n7618), .B(n7640), .Z(n7639) );
  AND U8014 ( .A(n9048), .B(n9049), .Z(n7640) );
  XOR U8015 ( .A(n7614), .B(n7619), .Z(n7618) );
  AND U8016 ( .A(n9050), .B(n9051), .Z(n7619) );
  XOR U8017 ( .A(n7616), .B(n7615), .Z(n7614) );
  AND U8018 ( .A(n9052), .B(n9053), .Z(n7615) );
  XNOR U8019 ( .A(n7626), .B(n7617), .Z(n7616) );
  AND U8020 ( .A(n9054), .B(n9055), .Z(n7617) );
  XOR U8021 ( .A(n7636), .B(n7625), .Z(n7626) );
  AND U8022 ( .A(n9056), .B(n9057), .Z(n7625) );
  XNOR U8023 ( .A(n9058), .B(n7631), .Z(n7636) );
  XOR U8024 ( .A(n7632), .B(n9059), .Z(n7631) );
  AND U8025 ( .A(n9060), .B(n9061), .Z(n9059) );
  XOR U8026 ( .A(n9062), .B(n9063), .Z(n7632) );
  NOR U8027 ( .A(n9064), .B(n9065), .Z(n9063) );
  AND U8028 ( .A(n9066), .B(n9067), .Z(n9065) );
  AND U8029 ( .A(n9068), .B(n9069), .Z(n9064) );
  XNOR U8030 ( .A(n9066), .B(n9067), .Z(n9062) );
  XNOR U8031 ( .A(n7623), .B(n7635), .Z(n9058) );
  AND U8032 ( .A(n9070), .B(n9071), .Z(n7635) );
  AND U8033 ( .A(n9072), .B(n9073), .Z(n7623) );
  AND U8034 ( .A(n127), .B(n129), .Z(n8034) );
  XOR U8035 ( .A(n8039), .B(n8038), .Z(n129) );
  NOR U8036 ( .A(n9074), .B(n9075), .Z(n8038) );
  XOR U8037 ( .A(n8041), .B(n8040), .Z(n8039) );
  NOR U8038 ( .A(n9076), .B(n9077), .Z(n8040) );
  XOR U8039 ( .A(n8043), .B(n8042), .Z(n8041) );
  NOR U8040 ( .A(n9078), .B(n9079), .Z(n8042) );
  XOR U8041 ( .A(n8045), .B(n8044), .Z(n8043) );
  NOR U8042 ( .A(n9080), .B(n9081), .Z(n8044) );
  XOR U8043 ( .A(n8047), .B(n8046), .Z(n8045) );
  NOR U8044 ( .A(n9082), .B(n9083), .Z(n8046) );
  XOR U8045 ( .A(n8049), .B(n8048), .Z(n8047) );
  NOR U8046 ( .A(n9084), .B(n9085), .Z(n8048) );
  XOR U8047 ( .A(n8051), .B(n8050), .Z(n8049) );
  NOR U8048 ( .A(n9086), .B(n9087), .Z(n8050) );
  XOR U8049 ( .A(n8053), .B(n8052), .Z(n8051) );
  NOR U8050 ( .A(n9088), .B(n9089), .Z(n8052) );
  XOR U8051 ( .A(n8055), .B(n8054), .Z(n8053) );
  NOR U8052 ( .A(n9090), .B(n9091), .Z(n8054) );
  XOR U8053 ( .A(n8057), .B(n8056), .Z(n8055) );
  NOR U8054 ( .A(n9092), .B(n9093), .Z(n8056) );
  XOR U8055 ( .A(n8059), .B(n8058), .Z(n8057) );
  NOR U8056 ( .A(n9094), .B(n9095), .Z(n8058) );
  XOR U8057 ( .A(n8061), .B(n8060), .Z(n8059) );
  NOR U8058 ( .A(n9096), .B(n9097), .Z(n8060) );
  XOR U8059 ( .A(n8063), .B(n8062), .Z(n8061) );
  NOR U8060 ( .A(n9098), .B(n9099), .Z(n8062) );
  XOR U8061 ( .A(n8065), .B(n8064), .Z(n8063) );
  NOR U8062 ( .A(n9100), .B(n9101), .Z(n8064) );
  XOR U8063 ( .A(n8067), .B(n8066), .Z(n8065) );
  NOR U8064 ( .A(n9102), .B(n9103), .Z(n8066) );
  XOR U8065 ( .A(n8069), .B(n8068), .Z(n8067) );
  NOR U8066 ( .A(n9104), .B(n9105), .Z(n8068) );
  XOR U8067 ( .A(n8071), .B(n8070), .Z(n8069) );
  NOR U8068 ( .A(n9106), .B(n9107), .Z(n8070) );
  XOR U8069 ( .A(n8073), .B(n8072), .Z(n8071) );
  NOR U8070 ( .A(n9108), .B(n9109), .Z(n8072) );
  XOR U8071 ( .A(n8075), .B(n8074), .Z(n8073) );
  NOR U8072 ( .A(n9110), .B(n9111), .Z(n8074) );
  XOR U8073 ( .A(n8077), .B(n8076), .Z(n8075) );
  NOR U8074 ( .A(n9112), .B(n9113), .Z(n8076) );
  XOR U8075 ( .A(n8079), .B(n8078), .Z(n8077) );
  NOR U8076 ( .A(n9114), .B(n9115), .Z(n8078) );
  XOR U8077 ( .A(n8081), .B(n8080), .Z(n8079) );
  NOR U8078 ( .A(n9116), .B(n9117), .Z(n8080) );
  XOR U8079 ( .A(n8083), .B(n8082), .Z(n8081) );
  NOR U8080 ( .A(n9118), .B(n9119), .Z(n8082) );
  XOR U8081 ( .A(n8085), .B(n8084), .Z(n8083) );
  NOR U8082 ( .A(n9120), .B(n9121), .Z(n8084) );
  XOR U8083 ( .A(n8087), .B(n8086), .Z(n8085) );
  NOR U8084 ( .A(n9122), .B(n9123), .Z(n8086) );
  XOR U8085 ( .A(n8089), .B(n8088), .Z(n8087) );
  NOR U8086 ( .A(n9124), .B(n9125), .Z(n8088) );
  XOR U8087 ( .A(n8091), .B(n8090), .Z(n8089) );
  NOR U8088 ( .A(n9126), .B(n9127), .Z(n8090) );
  XOR U8089 ( .A(n8093), .B(n8092), .Z(n8091) );
  NOR U8090 ( .A(n9128), .B(n9129), .Z(n8092) );
  XOR U8091 ( .A(n8095), .B(n8094), .Z(n8093) );
  NOR U8092 ( .A(n9130), .B(n9131), .Z(n8094) );
  XOR U8093 ( .A(n8097), .B(n8096), .Z(n8095) );
  NOR U8094 ( .A(n9132), .B(n9133), .Z(n8096) );
  XOR U8095 ( .A(n8099), .B(n8098), .Z(n8097) );
  NOR U8096 ( .A(n9134), .B(n9135), .Z(n8098) );
  XOR U8097 ( .A(n8101), .B(n8100), .Z(n8099) );
  NOR U8098 ( .A(n9136), .B(n9137), .Z(n8100) );
  XOR U8099 ( .A(n8103), .B(n8102), .Z(n8101) );
  NOR U8100 ( .A(n9138), .B(n9139), .Z(n8102) );
  XOR U8101 ( .A(n8105), .B(n8104), .Z(n8103) );
  NOR U8102 ( .A(n9140), .B(n9141), .Z(n8104) );
  XOR U8103 ( .A(n8107), .B(n8106), .Z(n8105) );
  NOR U8104 ( .A(n9142), .B(n9143), .Z(n8106) );
  XOR U8105 ( .A(n8109), .B(n8108), .Z(n8107) );
  NOR U8106 ( .A(n9144), .B(n9145), .Z(n8108) );
  XOR U8107 ( .A(n8111), .B(n8110), .Z(n8109) );
  NOR U8108 ( .A(n9146), .B(n9147), .Z(n8110) );
  XOR U8109 ( .A(n8113), .B(n8112), .Z(n8111) );
  NOR U8110 ( .A(n9148), .B(n9149), .Z(n8112) );
  XOR U8111 ( .A(n8115), .B(n8114), .Z(n8113) );
  NOR U8112 ( .A(n9150), .B(n9151), .Z(n8114) );
  XOR U8113 ( .A(n8117), .B(n8116), .Z(n8115) );
  NOR U8114 ( .A(n9152), .B(n9153), .Z(n8116) );
  XOR U8115 ( .A(n8119), .B(n8118), .Z(n8117) );
  NOR U8116 ( .A(n9154), .B(n9155), .Z(n8118) );
  XOR U8117 ( .A(n8121), .B(n8120), .Z(n8119) );
  NOR U8118 ( .A(n9156), .B(n9157), .Z(n8120) );
  XOR U8119 ( .A(n8123), .B(n8122), .Z(n8121) );
  NOR U8120 ( .A(n9158), .B(n9159), .Z(n8122) );
  XOR U8121 ( .A(n8125), .B(n8124), .Z(n8123) );
  NOR U8122 ( .A(n9160), .B(n9161), .Z(n8124) );
  XOR U8123 ( .A(n8127), .B(n8126), .Z(n8125) );
  NOR U8124 ( .A(n9162), .B(n9163), .Z(n8126) );
  XOR U8125 ( .A(n8129), .B(n8128), .Z(n8127) );
  NOR U8126 ( .A(n9164), .B(n9165), .Z(n8128) );
  XOR U8127 ( .A(n8131), .B(n8130), .Z(n8129) );
  NOR U8128 ( .A(n9166), .B(n9167), .Z(n8130) );
  XOR U8129 ( .A(n8133), .B(n8132), .Z(n8131) );
  NOR U8130 ( .A(n9168), .B(n9169), .Z(n8132) );
  XOR U8131 ( .A(n8135), .B(n8134), .Z(n8133) );
  NOR U8132 ( .A(n9170), .B(n9171), .Z(n8134) );
  XOR U8133 ( .A(n8137), .B(n8136), .Z(n8135) );
  NOR U8134 ( .A(n9172), .B(n9173), .Z(n8136) );
  XOR U8135 ( .A(n8139), .B(n8138), .Z(n8137) );
  NOR U8136 ( .A(n9174), .B(n9175), .Z(n8138) );
  XOR U8137 ( .A(n8141), .B(n8140), .Z(n8139) );
  NOR U8138 ( .A(n9176), .B(n9177), .Z(n8140) );
  XOR U8139 ( .A(n8143), .B(n8142), .Z(n8141) );
  NOR U8140 ( .A(n9178), .B(n9179), .Z(n8142) );
  XOR U8141 ( .A(n8145), .B(n8144), .Z(n8143) );
  NOR U8142 ( .A(n9180), .B(n9181), .Z(n8144) );
  XOR U8143 ( .A(n8147), .B(n8146), .Z(n8145) );
  NOR U8144 ( .A(n9182), .B(n9183), .Z(n8146) );
  XOR U8145 ( .A(n8149), .B(n8148), .Z(n8147) );
  NOR U8146 ( .A(n9184), .B(n9185), .Z(n8148) );
  XOR U8147 ( .A(n8151), .B(n8150), .Z(n8149) );
  NOR U8148 ( .A(n9186), .B(n9187), .Z(n8150) );
  XOR U8149 ( .A(n8153), .B(n8152), .Z(n8151) );
  NOR U8150 ( .A(n9188), .B(n9189), .Z(n8152) );
  XOR U8151 ( .A(n8155), .B(n8154), .Z(n8153) );
  NOR U8152 ( .A(n9190), .B(n9191), .Z(n8154) );
  XOR U8153 ( .A(n8157), .B(n8156), .Z(n8155) );
  NOR U8154 ( .A(n9192), .B(n9193), .Z(n8156) );
  XOR U8155 ( .A(n8159), .B(n8158), .Z(n8157) );
  NOR U8156 ( .A(n9194), .B(n9195), .Z(n8158) );
  XOR U8157 ( .A(n8161), .B(n8160), .Z(n8159) );
  NOR U8158 ( .A(n9196), .B(n9197), .Z(n8160) );
  XOR U8159 ( .A(n8163), .B(n8162), .Z(n8161) );
  NOR U8160 ( .A(n9198), .B(n9199), .Z(n8162) );
  XOR U8161 ( .A(n8165), .B(n8164), .Z(n8163) );
  NOR U8162 ( .A(n9200), .B(n9201), .Z(n8164) );
  XOR U8163 ( .A(n8167), .B(n8166), .Z(n8165) );
  NOR U8164 ( .A(n9202), .B(n9203), .Z(n8166) );
  XOR U8165 ( .A(n8169), .B(n8168), .Z(n8167) );
  NOR U8166 ( .A(n9204), .B(n9205), .Z(n8168) );
  XOR U8167 ( .A(n8171), .B(n8170), .Z(n8169) );
  NOR U8168 ( .A(n9206), .B(n9207), .Z(n8170) );
  XOR U8169 ( .A(n8173), .B(n8172), .Z(n8171) );
  NOR U8170 ( .A(n9208), .B(n9209), .Z(n8172) );
  XOR U8171 ( .A(n8175), .B(n8174), .Z(n8173) );
  NOR U8172 ( .A(n9210), .B(n9211), .Z(n8174) );
  XOR U8173 ( .A(n8177), .B(n8176), .Z(n8175) );
  NOR U8174 ( .A(n9212), .B(n9213), .Z(n8176) );
  XOR U8175 ( .A(n8179), .B(n8178), .Z(n8177) );
  NOR U8176 ( .A(n9214), .B(n9215), .Z(n8178) );
  XOR U8177 ( .A(n8181), .B(n8180), .Z(n8179) );
  NOR U8178 ( .A(n9216), .B(n9217), .Z(n8180) );
  XOR U8179 ( .A(n8183), .B(n8182), .Z(n8181) );
  NOR U8180 ( .A(n9218), .B(n9219), .Z(n8182) );
  XOR U8181 ( .A(n8185), .B(n8184), .Z(n8183) );
  NOR U8182 ( .A(n9220), .B(n9221), .Z(n8184) );
  XOR U8183 ( .A(n8187), .B(n8186), .Z(n8185) );
  NOR U8184 ( .A(n9222), .B(n9223), .Z(n8186) );
  XOR U8185 ( .A(n8189), .B(n8188), .Z(n8187) );
  NOR U8186 ( .A(n9224), .B(n9225), .Z(n8188) );
  XOR U8187 ( .A(n8191), .B(n8190), .Z(n8189) );
  NOR U8188 ( .A(n9226), .B(n9227), .Z(n8190) );
  XOR U8189 ( .A(n8193), .B(n8192), .Z(n8191) );
  NOR U8190 ( .A(n9228), .B(n9229), .Z(n8192) );
  XOR U8191 ( .A(n8195), .B(n8194), .Z(n8193) );
  NOR U8192 ( .A(n9230), .B(n9231), .Z(n8194) );
  XOR U8193 ( .A(n8197), .B(n8196), .Z(n8195) );
  NOR U8194 ( .A(n9232), .B(n9233), .Z(n8196) );
  XOR U8195 ( .A(n8199), .B(n8198), .Z(n8197) );
  NOR U8196 ( .A(n9234), .B(n9235), .Z(n8198) );
  XOR U8197 ( .A(n8201), .B(n8200), .Z(n8199) );
  NOR U8198 ( .A(n9236), .B(n9237), .Z(n8200) );
  XOR U8199 ( .A(n8203), .B(n8202), .Z(n8201) );
  NOR U8200 ( .A(n9238), .B(n9239), .Z(n8202) );
  XOR U8201 ( .A(n8205), .B(n8204), .Z(n8203) );
  NOR U8202 ( .A(n9240), .B(n9241), .Z(n8204) );
  XOR U8203 ( .A(n8207), .B(n8206), .Z(n8205) );
  NOR U8204 ( .A(n9242), .B(n9243), .Z(n8206) );
  XOR U8205 ( .A(n8209), .B(n8208), .Z(n8207) );
  NOR U8206 ( .A(n9244), .B(n9245), .Z(n8208) );
  XOR U8207 ( .A(n8211), .B(n8210), .Z(n8209) );
  NOR U8208 ( .A(n9246), .B(n9247), .Z(n8210) );
  XOR U8209 ( .A(n8213), .B(n8212), .Z(n8211) );
  NOR U8210 ( .A(n9248), .B(n9249), .Z(n8212) );
  XOR U8211 ( .A(n8215), .B(n8214), .Z(n8213) );
  NOR U8212 ( .A(n9250), .B(n9251), .Z(n8214) );
  XOR U8213 ( .A(n8217), .B(n8216), .Z(n8215) );
  NOR U8214 ( .A(n9252), .B(n9253), .Z(n8216) );
  XOR U8215 ( .A(n8219), .B(n8218), .Z(n8217) );
  NOR U8216 ( .A(n9254), .B(n9255), .Z(n8218) );
  XOR U8217 ( .A(n8221), .B(n8220), .Z(n8219) );
  NOR U8218 ( .A(n9256), .B(n9257), .Z(n8220) );
  XOR U8219 ( .A(n8223), .B(n8222), .Z(n8221) );
  NOR U8220 ( .A(n9258), .B(n9259), .Z(n8222) );
  XOR U8221 ( .A(n8225), .B(n8224), .Z(n8223) );
  NOR U8222 ( .A(n9260), .B(n9261), .Z(n8224) );
  XOR U8223 ( .A(n8227), .B(n8226), .Z(n8225) );
  NOR U8224 ( .A(n9262), .B(n9263), .Z(n8226) );
  XOR U8225 ( .A(n8229), .B(n8228), .Z(n8227) );
  NOR U8226 ( .A(n9264), .B(n9265), .Z(n8228) );
  XOR U8227 ( .A(n8231), .B(n8230), .Z(n8229) );
  NOR U8228 ( .A(n9266), .B(n9267), .Z(n8230) );
  XOR U8229 ( .A(n8233), .B(n8232), .Z(n8231) );
  NOR U8230 ( .A(n9268), .B(n9269), .Z(n8232) );
  XOR U8231 ( .A(n8235), .B(n8234), .Z(n8233) );
  NOR U8232 ( .A(n9270), .B(n9271), .Z(n8234) );
  XOR U8233 ( .A(n8237), .B(n8236), .Z(n8235) );
  NOR U8234 ( .A(n9272), .B(n9273), .Z(n8236) );
  XOR U8235 ( .A(n8239), .B(n8238), .Z(n8237) );
  NOR U8236 ( .A(n9274), .B(n9275), .Z(n8238) );
  XOR U8237 ( .A(n8241), .B(n8240), .Z(n8239) );
  NOR U8238 ( .A(n9276), .B(n9277), .Z(n8240) );
  XOR U8239 ( .A(n8243), .B(n8242), .Z(n8241) );
  NOR U8240 ( .A(n9278), .B(n9279), .Z(n8242) );
  XOR U8241 ( .A(n8245), .B(n8244), .Z(n8243) );
  NOR U8242 ( .A(n9280), .B(n9281), .Z(n8244) );
  XOR U8243 ( .A(n8247), .B(n8246), .Z(n8245) );
  NOR U8244 ( .A(n9282), .B(n9283), .Z(n8246) );
  XOR U8245 ( .A(n8249), .B(n8248), .Z(n8247) );
  NOR U8246 ( .A(n9284), .B(n9285), .Z(n8248) );
  XOR U8247 ( .A(n8251), .B(n8250), .Z(n8249) );
  NOR U8248 ( .A(n9286), .B(n9287), .Z(n8250) );
  XOR U8249 ( .A(n8253), .B(n8252), .Z(n8251) );
  NOR U8250 ( .A(n9288), .B(n9289), .Z(n8252) );
  XOR U8251 ( .A(n8255), .B(n8254), .Z(n8253) );
  NOR U8252 ( .A(n9290), .B(n9291), .Z(n8254) );
  XOR U8253 ( .A(n8257), .B(n8256), .Z(n8255) );
  NOR U8254 ( .A(n9292), .B(n9293), .Z(n8256) );
  XOR U8255 ( .A(n8259), .B(n8258), .Z(n8257) );
  NOR U8256 ( .A(n9294), .B(n9295), .Z(n8258) );
  XOR U8257 ( .A(n8261), .B(n8260), .Z(n8259) );
  NOR U8258 ( .A(n9296), .B(n9297), .Z(n8260) );
  XOR U8259 ( .A(n8263), .B(n8262), .Z(n8261) );
  NOR U8260 ( .A(n9298), .B(n9299), .Z(n8262) );
  XOR U8261 ( .A(n8265), .B(n8264), .Z(n8263) );
  NOR U8262 ( .A(n9300), .B(n9301), .Z(n8264) );
  XOR U8263 ( .A(n8267), .B(n8266), .Z(n8265) );
  NOR U8264 ( .A(n9302), .B(n9303), .Z(n8266) );
  XOR U8265 ( .A(n8269), .B(n8268), .Z(n8267) );
  NOR U8266 ( .A(n9304), .B(n9305), .Z(n8268) );
  XOR U8267 ( .A(n8271), .B(n8270), .Z(n8269) );
  NOR U8268 ( .A(n9306), .B(n9307), .Z(n8270) );
  XOR U8269 ( .A(n8273), .B(n8272), .Z(n8271) );
  NOR U8270 ( .A(n9308), .B(n9309), .Z(n8272) );
  XOR U8271 ( .A(n8275), .B(n8274), .Z(n8273) );
  NOR U8272 ( .A(n9310), .B(n9311), .Z(n8274) );
  XOR U8273 ( .A(n8277), .B(n8276), .Z(n8275) );
  NOR U8274 ( .A(n9312), .B(n9313), .Z(n8276) );
  XOR U8275 ( .A(n8279), .B(n8278), .Z(n8277) );
  NOR U8276 ( .A(n9314), .B(n9315), .Z(n8278) );
  XOR U8277 ( .A(n8281), .B(n8280), .Z(n8279) );
  NOR U8278 ( .A(n9316), .B(n9317), .Z(n8280) );
  XOR U8279 ( .A(n8283), .B(n8282), .Z(n8281) );
  NOR U8280 ( .A(n9318), .B(n9319), .Z(n8282) );
  XOR U8281 ( .A(n8285), .B(n8284), .Z(n8283) );
  NOR U8282 ( .A(n9320), .B(n9321), .Z(n8284) );
  XOR U8283 ( .A(n8287), .B(n8286), .Z(n8285) );
  NOR U8284 ( .A(n9322), .B(n9323), .Z(n8286) );
  XOR U8285 ( .A(n8289), .B(n8288), .Z(n8287) );
  NOR U8286 ( .A(n9324), .B(n9325), .Z(n8288) );
  XOR U8287 ( .A(n8291), .B(n8290), .Z(n8289) );
  NOR U8288 ( .A(n9326), .B(n9327), .Z(n8290) );
  XOR U8289 ( .A(n8293), .B(n8292), .Z(n8291) );
  NOR U8290 ( .A(n9328), .B(n9329), .Z(n8292) );
  XOR U8291 ( .A(n8295), .B(n8294), .Z(n8293) );
  NOR U8292 ( .A(n9330), .B(n9331), .Z(n8294) );
  XOR U8293 ( .A(n8299), .B(n8298), .Z(n8295) );
  NOR U8294 ( .A(n9332), .B(n9333), .Z(n8298) );
  XOR U8295 ( .A(n8301), .B(n8300), .Z(n8299) );
  NOR U8296 ( .A(n9334), .B(n9335), .Z(n8300) );
  XOR U8297 ( .A(n8303), .B(n8302), .Z(n8301) );
  NOR U8298 ( .A(n9336), .B(n9337), .Z(n8302) );
  XOR U8299 ( .A(n8305), .B(n8304), .Z(n8303) );
  NOR U8300 ( .A(n9338), .B(n9339), .Z(n8304) );
  XOR U8301 ( .A(n8307), .B(n8306), .Z(n8305) );
  NOR U8302 ( .A(n9340), .B(n9341), .Z(n8306) );
  XOR U8303 ( .A(n8309), .B(n8308), .Z(n8307) );
  NOR U8304 ( .A(n9342), .B(n9343), .Z(n8308) );
  XOR U8305 ( .A(n8311), .B(n8310), .Z(n8309) );
  NOR U8306 ( .A(n9344), .B(n9345), .Z(n8310) );
  XOR U8307 ( .A(n8313), .B(n8312), .Z(n8311) );
  NOR U8308 ( .A(n9346), .B(n9347), .Z(n8312) );
  XOR U8309 ( .A(n8315), .B(n8314), .Z(n8313) );
  NOR U8310 ( .A(n9348), .B(n9349), .Z(n8314) );
  XOR U8311 ( .A(n8317), .B(n8316), .Z(n8315) );
  NOR U8312 ( .A(n9350), .B(n9351), .Z(n8316) );
  XOR U8313 ( .A(n8319), .B(n8318), .Z(n8317) );
  NOR U8314 ( .A(n9352), .B(n9353), .Z(n8318) );
  XOR U8315 ( .A(n8321), .B(n8320), .Z(n8319) );
  NOR U8316 ( .A(n9354), .B(n9355), .Z(n8320) );
  XOR U8317 ( .A(n8323), .B(n8322), .Z(n8321) );
  NOR U8318 ( .A(n9356), .B(n9357), .Z(n8322) );
  XOR U8319 ( .A(n8325), .B(n8324), .Z(n8323) );
  NOR U8320 ( .A(n9358), .B(n9359), .Z(n8324) );
  XOR U8321 ( .A(n8327), .B(n8326), .Z(n8325) );
  NOR U8322 ( .A(n9360), .B(n9361), .Z(n8326) );
  XOR U8323 ( .A(n8329), .B(n8328), .Z(n8327) );
  NOR U8324 ( .A(n9362), .B(n9363), .Z(n8328) );
  XOR U8325 ( .A(n8331), .B(n8330), .Z(n8329) );
  NOR U8326 ( .A(n9364), .B(n9365), .Z(n8330) );
  XOR U8327 ( .A(n8333), .B(n8332), .Z(n8331) );
  NOR U8328 ( .A(n9366), .B(n9367), .Z(n8332) );
  XOR U8329 ( .A(n8335), .B(n8334), .Z(n8333) );
  NOR U8330 ( .A(n9368), .B(n9369), .Z(n8334) );
  XOR U8331 ( .A(n8337), .B(n8336), .Z(n8335) );
  NOR U8332 ( .A(n9370), .B(n9371), .Z(n8336) );
  XOR U8333 ( .A(n8339), .B(n8338), .Z(n8337) );
  NOR U8334 ( .A(n9372), .B(n9373), .Z(n8338) );
  XOR U8335 ( .A(n8341), .B(n8340), .Z(n8339) );
  NOR U8336 ( .A(n9374), .B(n9375), .Z(n8340) );
  XOR U8337 ( .A(n8343), .B(n8342), .Z(n8341) );
  NOR U8338 ( .A(n9376), .B(n9377), .Z(n8342) );
  XOR U8339 ( .A(n8345), .B(n8344), .Z(n8343) );
  NOR U8340 ( .A(n9378), .B(n9379), .Z(n8344) );
  XOR U8341 ( .A(n8347), .B(n8346), .Z(n8345) );
  NOR U8342 ( .A(n9380), .B(n9381), .Z(n8346) );
  XOR U8343 ( .A(n8349), .B(n8348), .Z(n8347) );
  NOR U8344 ( .A(n9382), .B(n9383), .Z(n8348) );
  XOR U8345 ( .A(n8351), .B(n8350), .Z(n8349) );
  NOR U8346 ( .A(n9384), .B(n9385), .Z(n8350) );
  XOR U8347 ( .A(n8353), .B(n8352), .Z(n8351) );
  NOR U8348 ( .A(n9386), .B(n9387), .Z(n8352) );
  XOR U8349 ( .A(n8355), .B(n8354), .Z(n8353) );
  NOR U8350 ( .A(n9388), .B(n9389), .Z(n8354) );
  XOR U8351 ( .A(n8357), .B(n8356), .Z(n8355) );
  NOR U8352 ( .A(n9390), .B(n9391), .Z(n8356) );
  XOR U8353 ( .A(n8359), .B(n8358), .Z(n8357) );
  NOR U8354 ( .A(n9392), .B(n9393), .Z(n8358) );
  XOR U8355 ( .A(n8361), .B(n8360), .Z(n8359) );
  NOR U8356 ( .A(n9394), .B(n9395), .Z(n8360) );
  XOR U8357 ( .A(n8363), .B(n8362), .Z(n8361) );
  NOR U8358 ( .A(n9396), .B(n9397), .Z(n8362) );
  XOR U8359 ( .A(n8365), .B(n8364), .Z(n8363) );
  NOR U8360 ( .A(n9398), .B(n9399), .Z(n8364) );
  XOR U8361 ( .A(n8367), .B(n8366), .Z(n8365) );
  NOR U8362 ( .A(n9400), .B(n9401), .Z(n8366) );
  XOR U8363 ( .A(n8369), .B(n8368), .Z(n8367) );
  NOR U8364 ( .A(n9402), .B(n9403), .Z(n8368) );
  XOR U8365 ( .A(n8371), .B(n8370), .Z(n8369) );
  NOR U8366 ( .A(n9404), .B(n9405), .Z(n8370) );
  XOR U8367 ( .A(n8373), .B(n8372), .Z(n8371) );
  NOR U8368 ( .A(n9406), .B(n9407), .Z(n8372) );
  XOR U8369 ( .A(n8375), .B(n8374), .Z(n8373) );
  NOR U8370 ( .A(n9408), .B(n9409), .Z(n8374) );
  XOR U8371 ( .A(n8377), .B(n8376), .Z(n8375) );
  NOR U8372 ( .A(n9410), .B(n9411), .Z(n8376) );
  XOR U8373 ( .A(n8379), .B(n8378), .Z(n8377) );
  NOR U8374 ( .A(n9412), .B(n9413), .Z(n8378) );
  XOR U8375 ( .A(n8381), .B(n8380), .Z(n8379) );
  NOR U8376 ( .A(n9414), .B(n9415), .Z(n8380) );
  XOR U8377 ( .A(n8383), .B(n8382), .Z(n8381) );
  NOR U8378 ( .A(n9416), .B(n9417), .Z(n8382) );
  XOR U8379 ( .A(n8385), .B(n8384), .Z(n8383) );
  NOR U8380 ( .A(n9418), .B(n9419), .Z(n8384) );
  XOR U8381 ( .A(n8387), .B(n8386), .Z(n8385) );
  NOR U8382 ( .A(n9420), .B(n9421), .Z(n8386) );
  XOR U8383 ( .A(n8389), .B(n8388), .Z(n8387) );
  NOR U8384 ( .A(n9422), .B(n9423), .Z(n8388) );
  XOR U8385 ( .A(n8391), .B(n8390), .Z(n8389) );
  NOR U8386 ( .A(n9424), .B(n9425), .Z(n8390) );
  XOR U8387 ( .A(n8393), .B(n8392), .Z(n8391) );
  NOR U8388 ( .A(n9426), .B(n9427), .Z(n8392) );
  XOR U8389 ( .A(n8395), .B(n8394), .Z(n8393) );
  NOR U8390 ( .A(n9428), .B(n9429), .Z(n8394) );
  XOR U8391 ( .A(n8397), .B(n8396), .Z(n8395) );
  NOR U8392 ( .A(n9430), .B(n9431), .Z(n8396) );
  XOR U8393 ( .A(n8399), .B(n8398), .Z(n8397) );
  NOR U8394 ( .A(n9432), .B(n9433), .Z(n8398) );
  XOR U8395 ( .A(n8401), .B(n8400), .Z(n8399) );
  NOR U8396 ( .A(n9434), .B(n9435), .Z(n8400) );
  XOR U8397 ( .A(n8403), .B(n8402), .Z(n8401) );
  NOR U8398 ( .A(n9436), .B(n9437), .Z(n8402) );
  XOR U8399 ( .A(n8405), .B(n8404), .Z(n8403) );
  NOR U8400 ( .A(n9438), .B(n9439), .Z(n8404) );
  XOR U8401 ( .A(n8407), .B(n8406), .Z(n8405) );
  NOR U8402 ( .A(n9440), .B(n9441), .Z(n8406) );
  XOR U8403 ( .A(n8409), .B(n8408), .Z(n8407) );
  NOR U8404 ( .A(n9442), .B(n9443), .Z(n8408) );
  XOR U8405 ( .A(n8411), .B(n8410), .Z(n8409) );
  NOR U8406 ( .A(n9444), .B(n9445), .Z(n8410) );
  XOR U8407 ( .A(n8413), .B(n8412), .Z(n8411) );
  NOR U8408 ( .A(n9446), .B(n9447), .Z(n8412) );
  XOR U8409 ( .A(n8415), .B(n8414), .Z(n8413) );
  NOR U8410 ( .A(n9448), .B(n9449), .Z(n8414) );
  XOR U8411 ( .A(n8417), .B(n8416), .Z(n8415) );
  NOR U8412 ( .A(n9450), .B(n9451), .Z(n8416) );
  XOR U8413 ( .A(n8419), .B(n8418), .Z(n8417) );
  NOR U8414 ( .A(n9452), .B(n9453), .Z(n8418) );
  XOR U8415 ( .A(n8421), .B(n8420), .Z(n8419) );
  NOR U8416 ( .A(n9454), .B(n9455), .Z(n8420) );
  XOR U8417 ( .A(n8423), .B(n8422), .Z(n8421) );
  NOR U8418 ( .A(n9456), .B(n9457), .Z(n8422) );
  XOR U8419 ( .A(n8425), .B(n8424), .Z(n8423) );
  NOR U8420 ( .A(n9458), .B(n9459), .Z(n8424) );
  XOR U8421 ( .A(n8427), .B(n8426), .Z(n8425) );
  NOR U8422 ( .A(n9460), .B(n9461), .Z(n8426) );
  XOR U8423 ( .A(n8429), .B(n8428), .Z(n8427) );
  NOR U8424 ( .A(n9462), .B(n9463), .Z(n8428) );
  XOR U8425 ( .A(n8431), .B(n8430), .Z(n8429) );
  NOR U8426 ( .A(n9464), .B(n9465), .Z(n8430) );
  XOR U8427 ( .A(n8433), .B(n8432), .Z(n8431) );
  NOR U8428 ( .A(n9466), .B(n9467), .Z(n8432) );
  XOR U8429 ( .A(n8435), .B(n8434), .Z(n8433) );
  NOR U8430 ( .A(n9468), .B(n9469), .Z(n8434) );
  XOR U8431 ( .A(n8437), .B(n8436), .Z(n8435) );
  NOR U8432 ( .A(n9470), .B(n9471), .Z(n8436) );
  XOR U8433 ( .A(n8439), .B(n8438), .Z(n8437) );
  NOR U8434 ( .A(n9472), .B(n9473), .Z(n8438) );
  XOR U8435 ( .A(n8441), .B(n8440), .Z(n8439) );
  NOR U8436 ( .A(n9474), .B(n9475), .Z(n8440) );
  XOR U8437 ( .A(n8443), .B(n8442), .Z(n8441) );
  NOR U8438 ( .A(n9476), .B(n9477), .Z(n8442) );
  XOR U8439 ( .A(n8445), .B(n8444), .Z(n8443) );
  NOR U8440 ( .A(n9478), .B(n9479), .Z(n8444) );
  XOR U8441 ( .A(n8447), .B(n8446), .Z(n8445) );
  NOR U8442 ( .A(n9480), .B(n9481), .Z(n8446) );
  XOR U8443 ( .A(n8449), .B(n8448), .Z(n8447) );
  NOR U8444 ( .A(n9482), .B(n9483), .Z(n8448) );
  XOR U8445 ( .A(n8451), .B(n8450), .Z(n8449) );
  NOR U8446 ( .A(n9484), .B(n9485), .Z(n8450) );
  XOR U8447 ( .A(n8453), .B(n8452), .Z(n8451) );
  NOR U8448 ( .A(n9486), .B(n9487), .Z(n8452) );
  XOR U8449 ( .A(n8455), .B(n8454), .Z(n8453) );
  NOR U8450 ( .A(n9488), .B(n9489), .Z(n8454) );
  XOR U8451 ( .A(n8457), .B(n8456), .Z(n8455) );
  NOR U8452 ( .A(n9490), .B(n9491), .Z(n8456) );
  XOR U8453 ( .A(n8459), .B(n8458), .Z(n8457) );
  NOR U8454 ( .A(n9492), .B(n9493), .Z(n8458) );
  XOR U8455 ( .A(n8461), .B(n8460), .Z(n8459) );
  NOR U8456 ( .A(n9494), .B(n9495), .Z(n8460) );
  XOR U8457 ( .A(n8463), .B(n8462), .Z(n8461) );
  NOR U8458 ( .A(n9496), .B(n9497), .Z(n8462) );
  XOR U8459 ( .A(n8465), .B(n8464), .Z(n8463) );
  NOR U8460 ( .A(n9498), .B(n9499), .Z(n8464) );
  XOR U8461 ( .A(n8467), .B(n8466), .Z(n8465) );
  NOR U8462 ( .A(n9500), .B(n9501), .Z(n8466) );
  XOR U8463 ( .A(n8469), .B(n8468), .Z(n8467) );
  NOR U8464 ( .A(n9502), .B(n9503), .Z(n8468) );
  XOR U8465 ( .A(n8471), .B(n8470), .Z(n8469) );
  NOR U8466 ( .A(n9504), .B(n9505), .Z(n8470) );
  XOR U8467 ( .A(n8473), .B(n8472), .Z(n8471) );
  NOR U8468 ( .A(n9506), .B(n9507), .Z(n8472) );
  XOR U8469 ( .A(n8475), .B(n8474), .Z(n8473) );
  NOR U8470 ( .A(n9508), .B(n9509), .Z(n8474) );
  XOR U8471 ( .A(n8477), .B(n8476), .Z(n8475) );
  NOR U8472 ( .A(n9510), .B(n9511), .Z(n8476) );
  XOR U8473 ( .A(n8479), .B(n8478), .Z(n8477) );
  NOR U8474 ( .A(n9512), .B(n9513), .Z(n8478) );
  XOR U8475 ( .A(n8481), .B(n8480), .Z(n8479) );
  NOR U8476 ( .A(n9514), .B(n9515), .Z(n8480) );
  XOR U8477 ( .A(n8483), .B(n8482), .Z(n8481) );
  NOR U8478 ( .A(n9516), .B(n9517), .Z(n8482) );
  XOR U8479 ( .A(n8485), .B(n8484), .Z(n8483) );
  NOR U8480 ( .A(n9518), .B(n9519), .Z(n8484) );
  XOR U8481 ( .A(n8487), .B(n8486), .Z(n8485) );
  NOR U8482 ( .A(n9520), .B(n9521), .Z(n8486) );
  XOR U8483 ( .A(n8489), .B(n8488), .Z(n8487) );
  NOR U8484 ( .A(n9522), .B(n9523), .Z(n8488) );
  XOR U8485 ( .A(n8491), .B(n8490), .Z(n8489) );
  NOR U8486 ( .A(n9524), .B(n9525), .Z(n8490) );
  XOR U8487 ( .A(n8493), .B(n8492), .Z(n8491) );
  NOR U8488 ( .A(n9526), .B(n9527), .Z(n8492) );
  XOR U8489 ( .A(n8495), .B(n8494), .Z(n8493) );
  NOR U8490 ( .A(n9528), .B(n9529), .Z(n8494) );
  XOR U8491 ( .A(n8497), .B(n8496), .Z(n8495) );
  NOR U8492 ( .A(n9530), .B(n9531), .Z(n8496) );
  XOR U8493 ( .A(n8499), .B(n8498), .Z(n8497) );
  NOR U8494 ( .A(n9532), .B(n9533), .Z(n8498) );
  XOR U8495 ( .A(n8501), .B(n8500), .Z(n8499) );
  NOR U8496 ( .A(n9534), .B(n9535), .Z(n8500) );
  XOR U8497 ( .A(n8503), .B(n8502), .Z(n8501) );
  NOR U8498 ( .A(n9536), .B(n9537), .Z(n8502) );
  XOR U8499 ( .A(n8505), .B(n8504), .Z(n8503) );
  NOR U8500 ( .A(n9538), .B(n9539), .Z(n8504) );
  XOR U8501 ( .A(n8507), .B(n8506), .Z(n8505) );
  NOR U8502 ( .A(n9540), .B(n9541), .Z(n8506) );
  XOR U8503 ( .A(n8509), .B(n8508), .Z(n8507) );
  NOR U8504 ( .A(n9542), .B(n9543), .Z(n8508) );
  XOR U8505 ( .A(n8511), .B(n8510), .Z(n8509) );
  NOR U8506 ( .A(n9544), .B(n9545), .Z(n8510) );
  XOR U8507 ( .A(n8513), .B(n8512), .Z(n8511) );
  NOR U8508 ( .A(n9546), .B(n9547), .Z(n8512) );
  XOR U8509 ( .A(n8515), .B(n8514), .Z(n8513) );
  NOR U8510 ( .A(n9548), .B(n9549), .Z(n8514) );
  XOR U8511 ( .A(n8517), .B(n8516), .Z(n8515) );
  NOR U8512 ( .A(n9550), .B(n9551), .Z(n8516) );
  XOR U8513 ( .A(n8519), .B(n8518), .Z(n8517) );
  NOR U8514 ( .A(n9552), .B(n9553), .Z(n8518) );
  XOR U8515 ( .A(n8521), .B(n8520), .Z(n8519) );
  NOR U8516 ( .A(n9554), .B(n9555), .Z(n8520) );
  XOR U8517 ( .A(n8523), .B(n8522), .Z(n8521) );
  NOR U8518 ( .A(n9556), .B(n9557), .Z(n8522) );
  XOR U8519 ( .A(n8525), .B(n8524), .Z(n8523) );
  NOR U8520 ( .A(n9558), .B(n9559), .Z(n8524) );
  XOR U8521 ( .A(n8527), .B(n8526), .Z(n8525) );
  NOR U8522 ( .A(n9560), .B(n9561), .Z(n8526) );
  XOR U8523 ( .A(n8529), .B(n8528), .Z(n8527) );
  NOR U8524 ( .A(n9562), .B(n9563), .Z(n8528) );
  XOR U8525 ( .A(n8531), .B(n8530), .Z(n8529) );
  NOR U8526 ( .A(n9564), .B(n9565), .Z(n8530) );
  XOR U8527 ( .A(n8533), .B(n8532), .Z(n8531) );
  NOR U8528 ( .A(n9566), .B(n9567), .Z(n8532) );
  XOR U8529 ( .A(n8535), .B(n8534), .Z(n8533) );
  NOR U8530 ( .A(n9568), .B(n9569), .Z(n8534) );
  XOR U8531 ( .A(n8537), .B(n8536), .Z(n8535) );
  NOR U8532 ( .A(n9570), .B(n9571), .Z(n8536) );
  XOR U8533 ( .A(n8539), .B(n8538), .Z(n8537) );
  NOR U8534 ( .A(n9572), .B(n9573), .Z(n8538) );
  XOR U8535 ( .A(n8553), .B(n8552), .Z(n8539) );
  NOR U8536 ( .A(n9574), .B(n9575), .Z(n8552) );
  XOR U8537 ( .A(n8555), .B(n8554), .Z(n8553) );
  NOR U8538 ( .A(n9576), .B(n9577), .Z(n8554) );
  XOR U8539 ( .A(n8543), .B(n8542), .Z(n8555) );
  NOR U8540 ( .A(n9578), .B(n9579), .Z(n8542) );
  XOR U8541 ( .A(n8550), .B(n8551), .Z(n8543) );
  XOR U8542 ( .A(n8548), .B(n8549), .Z(n8551) );
  NOR U8543 ( .A(n9580), .B(n9581), .Z(n8549) );
  NOR U8544 ( .A(n9582), .B(n9583), .Z(n8548) );
  NOR U8545 ( .A(n9584), .B(n9585), .Z(n8550) );
  XNOR U8546 ( .A(n8557), .B(n8556), .Z(n127) );
  NOR U8547 ( .A(n9074), .B(p_input[510]), .Z(n8556) );
  XOR U8548 ( .A(n8559), .B(n8558), .Z(n8557) );
  NOR U8549 ( .A(n9076), .B(p_input[508]), .Z(n8558) );
  XOR U8550 ( .A(n8561), .B(n8560), .Z(n8559) );
  NOR U8551 ( .A(n9078), .B(p_input[506]), .Z(n8560) );
  XOR U8552 ( .A(n8563), .B(n8562), .Z(n8561) );
  NOR U8553 ( .A(n9080), .B(p_input[504]), .Z(n8562) );
  XOR U8554 ( .A(n8565), .B(n8564), .Z(n8563) );
  NOR U8555 ( .A(n9082), .B(p_input[502]), .Z(n8564) );
  XOR U8556 ( .A(n8567), .B(n8566), .Z(n8565) );
  NOR U8557 ( .A(n9084), .B(p_input[500]), .Z(n8566) );
  XOR U8558 ( .A(n8569), .B(n8568), .Z(n8567) );
  NOR U8559 ( .A(n9086), .B(p_input[498]), .Z(n8568) );
  XOR U8560 ( .A(n8571), .B(n8570), .Z(n8569) );
  NOR U8561 ( .A(n9088), .B(p_input[496]), .Z(n8570) );
  XOR U8562 ( .A(n8573), .B(n8572), .Z(n8571) );
  NOR U8563 ( .A(n9090), .B(p_input[494]), .Z(n8572) );
  XOR U8564 ( .A(n8575), .B(n8574), .Z(n8573) );
  NOR U8565 ( .A(n9092), .B(p_input[492]), .Z(n8574) );
  XOR U8566 ( .A(n8577), .B(n8576), .Z(n8575) );
  NOR U8567 ( .A(n9094), .B(p_input[490]), .Z(n8576) );
  XOR U8568 ( .A(n8579), .B(n8578), .Z(n8577) );
  NOR U8569 ( .A(n9096), .B(p_input[488]), .Z(n8578) );
  XOR U8570 ( .A(n8581), .B(n8580), .Z(n8579) );
  NOR U8571 ( .A(n9098), .B(p_input[486]), .Z(n8580) );
  XOR U8572 ( .A(n8583), .B(n8582), .Z(n8581) );
  NOR U8573 ( .A(n9100), .B(p_input[484]), .Z(n8582) );
  XOR U8574 ( .A(n8585), .B(n8584), .Z(n8583) );
  NOR U8575 ( .A(n9102), .B(p_input[482]), .Z(n8584) );
  XOR U8576 ( .A(n8587), .B(n8586), .Z(n8585) );
  NOR U8577 ( .A(n9104), .B(p_input[480]), .Z(n8586) );
  XOR U8578 ( .A(n8589), .B(n8588), .Z(n8587) );
  NOR U8579 ( .A(n9106), .B(p_input[478]), .Z(n8588) );
  XOR U8580 ( .A(n8591), .B(n8590), .Z(n8589) );
  NOR U8581 ( .A(n9108), .B(p_input[476]), .Z(n8590) );
  XOR U8582 ( .A(n8593), .B(n8592), .Z(n8591) );
  NOR U8583 ( .A(n9110), .B(p_input[474]), .Z(n8592) );
  XOR U8584 ( .A(n8595), .B(n8594), .Z(n8593) );
  NOR U8585 ( .A(n9112), .B(p_input[472]), .Z(n8594) );
  XOR U8586 ( .A(n8597), .B(n8596), .Z(n8595) );
  NOR U8587 ( .A(n9114), .B(p_input[470]), .Z(n8596) );
  XOR U8588 ( .A(n8599), .B(n8598), .Z(n8597) );
  NOR U8589 ( .A(n9116), .B(p_input[468]), .Z(n8598) );
  XOR U8590 ( .A(n8601), .B(n8600), .Z(n8599) );
  NOR U8591 ( .A(n9118), .B(p_input[466]), .Z(n8600) );
  XOR U8592 ( .A(n8603), .B(n8602), .Z(n8601) );
  NOR U8593 ( .A(n9120), .B(p_input[464]), .Z(n8602) );
  XOR U8594 ( .A(n8605), .B(n8604), .Z(n8603) );
  NOR U8595 ( .A(n9122), .B(p_input[462]), .Z(n8604) );
  XOR U8596 ( .A(n8607), .B(n8606), .Z(n8605) );
  NOR U8597 ( .A(n9124), .B(p_input[460]), .Z(n8606) );
  XOR U8598 ( .A(n8609), .B(n8608), .Z(n8607) );
  NOR U8599 ( .A(n9126), .B(p_input[458]), .Z(n8608) );
  XOR U8600 ( .A(n8611), .B(n8610), .Z(n8609) );
  NOR U8601 ( .A(n9128), .B(p_input[456]), .Z(n8610) );
  XOR U8602 ( .A(n8613), .B(n8612), .Z(n8611) );
  NOR U8603 ( .A(n9130), .B(p_input[454]), .Z(n8612) );
  XOR U8604 ( .A(n8615), .B(n8614), .Z(n8613) );
  NOR U8605 ( .A(n9132), .B(p_input[452]), .Z(n8614) );
  XOR U8606 ( .A(n8617), .B(n8616), .Z(n8615) );
  NOR U8607 ( .A(n9134), .B(p_input[450]), .Z(n8616) );
  XOR U8608 ( .A(n8619), .B(n8618), .Z(n8617) );
  NOR U8609 ( .A(n9136), .B(p_input[448]), .Z(n8618) );
  XOR U8610 ( .A(n8621), .B(n8620), .Z(n8619) );
  NOR U8611 ( .A(n9138), .B(p_input[446]), .Z(n8620) );
  XOR U8612 ( .A(n8623), .B(n8622), .Z(n8621) );
  NOR U8613 ( .A(n9140), .B(p_input[444]), .Z(n8622) );
  XOR U8614 ( .A(n8625), .B(n8624), .Z(n8623) );
  NOR U8615 ( .A(n9142), .B(p_input[442]), .Z(n8624) );
  XOR U8616 ( .A(n8627), .B(n8626), .Z(n8625) );
  NOR U8617 ( .A(n9144), .B(p_input[440]), .Z(n8626) );
  XOR U8618 ( .A(n8629), .B(n8628), .Z(n8627) );
  NOR U8619 ( .A(n9146), .B(p_input[438]), .Z(n8628) );
  XOR U8620 ( .A(n8631), .B(n8630), .Z(n8629) );
  NOR U8621 ( .A(n9148), .B(p_input[436]), .Z(n8630) );
  XOR U8622 ( .A(n8633), .B(n8632), .Z(n8631) );
  NOR U8623 ( .A(n9150), .B(p_input[434]), .Z(n8632) );
  XOR U8624 ( .A(n8635), .B(n8634), .Z(n8633) );
  NOR U8625 ( .A(n9152), .B(p_input[432]), .Z(n8634) );
  XOR U8626 ( .A(n8637), .B(n8636), .Z(n8635) );
  NOR U8627 ( .A(n9154), .B(p_input[430]), .Z(n8636) );
  XOR U8628 ( .A(n8639), .B(n8638), .Z(n8637) );
  NOR U8629 ( .A(n9156), .B(p_input[428]), .Z(n8638) );
  XOR U8630 ( .A(n8641), .B(n8640), .Z(n8639) );
  NOR U8631 ( .A(n9158), .B(p_input[426]), .Z(n8640) );
  XOR U8632 ( .A(n8643), .B(n8642), .Z(n8641) );
  NOR U8633 ( .A(n9160), .B(p_input[424]), .Z(n8642) );
  XOR U8634 ( .A(n8645), .B(n8644), .Z(n8643) );
  NOR U8635 ( .A(n9162), .B(p_input[422]), .Z(n8644) );
  XOR U8636 ( .A(n8647), .B(n8646), .Z(n8645) );
  NOR U8637 ( .A(n9164), .B(p_input[420]), .Z(n8646) );
  XOR U8638 ( .A(n8649), .B(n8648), .Z(n8647) );
  NOR U8639 ( .A(n9166), .B(p_input[418]), .Z(n8648) );
  XOR U8640 ( .A(n8651), .B(n8650), .Z(n8649) );
  NOR U8641 ( .A(n9168), .B(p_input[416]), .Z(n8650) );
  XOR U8642 ( .A(n8653), .B(n8652), .Z(n8651) );
  NOR U8643 ( .A(n9170), .B(p_input[414]), .Z(n8652) );
  XOR U8644 ( .A(n8655), .B(n8654), .Z(n8653) );
  NOR U8645 ( .A(n9172), .B(p_input[412]), .Z(n8654) );
  XOR U8646 ( .A(n8657), .B(n8656), .Z(n8655) );
  NOR U8647 ( .A(n9174), .B(p_input[410]), .Z(n8656) );
  XOR U8648 ( .A(n8659), .B(n8658), .Z(n8657) );
  NOR U8649 ( .A(n9176), .B(p_input[408]), .Z(n8658) );
  XOR U8650 ( .A(n8661), .B(n8660), .Z(n8659) );
  NOR U8651 ( .A(n9178), .B(p_input[406]), .Z(n8660) );
  XOR U8652 ( .A(n8663), .B(n8662), .Z(n8661) );
  NOR U8653 ( .A(n9180), .B(p_input[404]), .Z(n8662) );
  XOR U8654 ( .A(n8665), .B(n8664), .Z(n8663) );
  NOR U8655 ( .A(n9182), .B(p_input[402]), .Z(n8664) );
  XOR U8656 ( .A(n8667), .B(n8666), .Z(n8665) );
  NOR U8657 ( .A(n9184), .B(p_input[400]), .Z(n8666) );
  XOR U8658 ( .A(n8669), .B(n8668), .Z(n8667) );
  NOR U8659 ( .A(n9186), .B(p_input[398]), .Z(n8668) );
  XOR U8660 ( .A(n8671), .B(n8670), .Z(n8669) );
  NOR U8661 ( .A(n9188), .B(p_input[396]), .Z(n8670) );
  XOR U8662 ( .A(n8673), .B(n8672), .Z(n8671) );
  NOR U8663 ( .A(n9190), .B(p_input[394]), .Z(n8672) );
  XOR U8664 ( .A(n8675), .B(n8674), .Z(n8673) );
  NOR U8665 ( .A(n9192), .B(p_input[392]), .Z(n8674) );
  XOR U8666 ( .A(n8677), .B(n8676), .Z(n8675) );
  NOR U8667 ( .A(n9194), .B(p_input[390]), .Z(n8676) );
  XOR U8668 ( .A(n8679), .B(n8678), .Z(n8677) );
  NOR U8669 ( .A(n9196), .B(p_input[388]), .Z(n8678) );
  XOR U8670 ( .A(n8681), .B(n8680), .Z(n8679) );
  NOR U8671 ( .A(n9198), .B(p_input[386]), .Z(n8680) );
  XOR U8672 ( .A(n8683), .B(n8682), .Z(n8681) );
  NOR U8673 ( .A(n9200), .B(p_input[384]), .Z(n8682) );
  XOR U8674 ( .A(n8685), .B(n8684), .Z(n8683) );
  NOR U8675 ( .A(n9202), .B(p_input[382]), .Z(n8684) );
  XOR U8676 ( .A(n8687), .B(n8686), .Z(n8685) );
  NOR U8677 ( .A(n9204), .B(p_input[380]), .Z(n8686) );
  XOR U8678 ( .A(n8689), .B(n8688), .Z(n8687) );
  NOR U8679 ( .A(n9206), .B(p_input[378]), .Z(n8688) );
  XOR U8680 ( .A(n8691), .B(n8690), .Z(n8689) );
  NOR U8681 ( .A(n9208), .B(p_input[376]), .Z(n8690) );
  XOR U8682 ( .A(n8693), .B(n8692), .Z(n8691) );
  NOR U8683 ( .A(n9210), .B(p_input[374]), .Z(n8692) );
  XOR U8684 ( .A(n8695), .B(n8694), .Z(n8693) );
  NOR U8685 ( .A(n9212), .B(p_input[372]), .Z(n8694) );
  XOR U8686 ( .A(n8697), .B(n8696), .Z(n8695) );
  NOR U8687 ( .A(n9214), .B(p_input[370]), .Z(n8696) );
  XOR U8688 ( .A(n8699), .B(n8698), .Z(n8697) );
  NOR U8689 ( .A(n9216), .B(p_input[368]), .Z(n8698) );
  XOR U8690 ( .A(n8701), .B(n8700), .Z(n8699) );
  NOR U8691 ( .A(n9218), .B(p_input[366]), .Z(n8700) );
  XOR U8692 ( .A(n8703), .B(n8702), .Z(n8701) );
  NOR U8693 ( .A(n9220), .B(p_input[364]), .Z(n8702) );
  XOR U8694 ( .A(n8705), .B(n8704), .Z(n8703) );
  NOR U8695 ( .A(n9222), .B(p_input[362]), .Z(n8704) );
  XOR U8696 ( .A(n8707), .B(n8706), .Z(n8705) );
  NOR U8697 ( .A(n9224), .B(p_input[360]), .Z(n8706) );
  XOR U8698 ( .A(n8709), .B(n8708), .Z(n8707) );
  NOR U8699 ( .A(n9226), .B(p_input[358]), .Z(n8708) );
  XOR U8700 ( .A(n8711), .B(n8710), .Z(n8709) );
  NOR U8701 ( .A(n9228), .B(p_input[356]), .Z(n8710) );
  XOR U8702 ( .A(n8713), .B(n8712), .Z(n8711) );
  NOR U8703 ( .A(n9230), .B(p_input[354]), .Z(n8712) );
  XOR U8704 ( .A(n8715), .B(n8714), .Z(n8713) );
  NOR U8705 ( .A(n9232), .B(p_input[352]), .Z(n8714) );
  XOR U8706 ( .A(n8717), .B(n8716), .Z(n8715) );
  NOR U8707 ( .A(n9234), .B(p_input[350]), .Z(n8716) );
  XOR U8708 ( .A(n8719), .B(n8718), .Z(n8717) );
  NOR U8709 ( .A(n9236), .B(p_input[348]), .Z(n8718) );
  XOR U8710 ( .A(n8721), .B(n8720), .Z(n8719) );
  NOR U8711 ( .A(n9238), .B(p_input[346]), .Z(n8720) );
  XOR U8712 ( .A(n8723), .B(n8722), .Z(n8721) );
  NOR U8713 ( .A(n9240), .B(p_input[344]), .Z(n8722) );
  XOR U8714 ( .A(n8725), .B(n8724), .Z(n8723) );
  NOR U8715 ( .A(n9242), .B(p_input[342]), .Z(n8724) );
  XOR U8716 ( .A(n8727), .B(n8726), .Z(n8725) );
  NOR U8717 ( .A(n9244), .B(p_input[340]), .Z(n8726) );
  XOR U8718 ( .A(n8729), .B(n8728), .Z(n8727) );
  NOR U8719 ( .A(n9246), .B(p_input[338]), .Z(n8728) );
  XOR U8720 ( .A(n8731), .B(n8730), .Z(n8729) );
  NOR U8721 ( .A(n9248), .B(p_input[336]), .Z(n8730) );
  XOR U8722 ( .A(n8733), .B(n8732), .Z(n8731) );
  NOR U8723 ( .A(n9250), .B(p_input[334]), .Z(n8732) );
  XOR U8724 ( .A(n8735), .B(n8734), .Z(n8733) );
  NOR U8725 ( .A(n9252), .B(p_input[332]), .Z(n8734) );
  XOR U8726 ( .A(n8737), .B(n8736), .Z(n8735) );
  NOR U8727 ( .A(n9254), .B(p_input[330]), .Z(n8736) );
  XOR U8728 ( .A(n8739), .B(n8738), .Z(n8737) );
  NOR U8729 ( .A(n9256), .B(p_input[328]), .Z(n8738) );
  XOR U8730 ( .A(n8741), .B(n8740), .Z(n8739) );
  NOR U8731 ( .A(n9258), .B(p_input[326]), .Z(n8740) );
  XOR U8732 ( .A(n8743), .B(n8742), .Z(n8741) );
  NOR U8733 ( .A(n9260), .B(p_input[324]), .Z(n8742) );
  XOR U8734 ( .A(n8745), .B(n8744), .Z(n8743) );
  NOR U8735 ( .A(n9262), .B(p_input[322]), .Z(n8744) );
  XOR U8736 ( .A(n8747), .B(n8746), .Z(n8745) );
  NOR U8737 ( .A(n9264), .B(p_input[320]), .Z(n8746) );
  XOR U8738 ( .A(n8749), .B(n8748), .Z(n8747) );
  NOR U8739 ( .A(n9266), .B(p_input[318]), .Z(n8748) );
  XOR U8740 ( .A(n8751), .B(n8750), .Z(n8749) );
  NOR U8741 ( .A(n9268), .B(p_input[316]), .Z(n8750) );
  XOR U8742 ( .A(n8753), .B(n8752), .Z(n8751) );
  NOR U8743 ( .A(n9270), .B(p_input[314]), .Z(n8752) );
  XOR U8744 ( .A(n8755), .B(n8754), .Z(n8753) );
  NOR U8745 ( .A(n9272), .B(p_input[312]), .Z(n8754) );
  XOR U8746 ( .A(n8757), .B(n8756), .Z(n8755) );
  NOR U8747 ( .A(n9274), .B(p_input[310]), .Z(n8756) );
  XOR U8748 ( .A(n8759), .B(n8758), .Z(n8757) );
  NOR U8749 ( .A(n9276), .B(p_input[308]), .Z(n8758) );
  XOR U8750 ( .A(n8761), .B(n8760), .Z(n8759) );
  NOR U8751 ( .A(n9278), .B(p_input[306]), .Z(n8760) );
  XOR U8752 ( .A(n8763), .B(n8762), .Z(n8761) );
  NOR U8753 ( .A(n9280), .B(p_input[304]), .Z(n8762) );
  XOR U8754 ( .A(n8765), .B(n8764), .Z(n8763) );
  NOR U8755 ( .A(n9282), .B(p_input[302]), .Z(n8764) );
  XOR U8756 ( .A(n8767), .B(n8766), .Z(n8765) );
  NOR U8757 ( .A(n9284), .B(p_input[300]), .Z(n8766) );
  XOR U8758 ( .A(n8769), .B(n8768), .Z(n8767) );
  NOR U8759 ( .A(n9286), .B(p_input[298]), .Z(n8768) );
  XOR U8760 ( .A(n8771), .B(n8770), .Z(n8769) );
  NOR U8761 ( .A(n9288), .B(p_input[296]), .Z(n8770) );
  XOR U8762 ( .A(n8773), .B(n8772), .Z(n8771) );
  NOR U8763 ( .A(n9290), .B(p_input[294]), .Z(n8772) );
  XOR U8764 ( .A(n8775), .B(n8774), .Z(n8773) );
  NOR U8765 ( .A(n9292), .B(p_input[292]), .Z(n8774) );
  XOR U8766 ( .A(n8777), .B(n8776), .Z(n8775) );
  NOR U8767 ( .A(n9294), .B(p_input[290]), .Z(n8776) );
  XOR U8768 ( .A(n8779), .B(n8778), .Z(n8777) );
  NOR U8769 ( .A(n9296), .B(p_input[288]), .Z(n8778) );
  XOR U8770 ( .A(n8781), .B(n8780), .Z(n8779) );
  NOR U8771 ( .A(n9298), .B(p_input[286]), .Z(n8780) );
  XOR U8772 ( .A(n8783), .B(n8782), .Z(n8781) );
  NOR U8773 ( .A(n9300), .B(p_input[284]), .Z(n8782) );
  XOR U8774 ( .A(n8785), .B(n8784), .Z(n8783) );
  NOR U8775 ( .A(n9302), .B(p_input[282]), .Z(n8784) );
  XOR U8776 ( .A(n8787), .B(n8786), .Z(n8785) );
  NOR U8777 ( .A(n9304), .B(p_input[280]), .Z(n8786) );
  XOR U8778 ( .A(n8789), .B(n8788), .Z(n8787) );
  NOR U8779 ( .A(n9306), .B(p_input[278]), .Z(n8788) );
  XOR U8780 ( .A(n8791), .B(n8790), .Z(n8789) );
  NOR U8781 ( .A(n9308), .B(p_input[276]), .Z(n8790) );
  XOR U8782 ( .A(n8793), .B(n8792), .Z(n8791) );
  NOR U8783 ( .A(n9310), .B(p_input[274]), .Z(n8792) );
  XOR U8784 ( .A(n8795), .B(n8794), .Z(n8793) );
  NOR U8785 ( .A(n9312), .B(p_input[272]), .Z(n8794) );
  XOR U8786 ( .A(n8797), .B(n8796), .Z(n8795) );
  NOR U8787 ( .A(n9314), .B(p_input[270]), .Z(n8796) );
  XOR U8788 ( .A(n8799), .B(n8798), .Z(n8797) );
  NOR U8789 ( .A(n9316), .B(p_input[268]), .Z(n8798) );
  XOR U8790 ( .A(n8801), .B(n8800), .Z(n8799) );
  NOR U8791 ( .A(n9318), .B(p_input[266]), .Z(n8800) );
  XOR U8792 ( .A(n8803), .B(n8802), .Z(n8801) );
  NOR U8793 ( .A(n9320), .B(p_input[264]), .Z(n8802) );
  XOR U8794 ( .A(n8805), .B(n8804), .Z(n8803) );
  NOR U8795 ( .A(n9322), .B(p_input[262]), .Z(n8804) );
  XOR U8796 ( .A(n8807), .B(n8806), .Z(n8805) );
  NOR U8797 ( .A(n9324), .B(p_input[260]), .Z(n8806) );
  XOR U8798 ( .A(n8809), .B(n8808), .Z(n8807) );
  NOR U8799 ( .A(n9326), .B(p_input[258]), .Z(n8808) );
  XOR U8800 ( .A(n8811), .B(n8810), .Z(n8809) );
  NOR U8801 ( .A(n9328), .B(p_input[256]), .Z(n8810) );
  XOR U8802 ( .A(n8813), .B(n8812), .Z(n8811) );
  NOR U8803 ( .A(n9330), .B(p_input[254]), .Z(n8812) );
  XOR U8804 ( .A(n8817), .B(n8816), .Z(n8813) );
  NOR U8805 ( .A(n9332), .B(p_input[252]), .Z(n8816) );
  XOR U8806 ( .A(n8819), .B(n8818), .Z(n8817) );
  NOR U8807 ( .A(n9334), .B(p_input[250]), .Z(n8818) );
  XOR U8808 ( .A(n8821), .B(n8820), .Z(n8819) );
  NOR U8809 ( .A(n9336), .B(p_input[248]), .Z(n8820) );
  XOR U8810 ( .A(n8823), .B(n8822), .Z(n8821) );
  NOR U8811 ( .A(n9338), .B(p_input[246]), .Z(n8822) );
  XOR U8812 ( .A(n8825), .B(n8824), .Z(n8823) );
  NOR U8813 ( .A(n9340), .B(p_input[244]), .Z(n8824) );
  XOR U8814 ( .A(n8827), .B(n8826), .Z(n8825) );
  NOR U8815 ( .A(n9342), .B(p_input[242]), .Z(n8826) );
  XOR U8816 ( .A(n8829), .B(n8828), .Z(n8827) );
  NOR U8817 ( .A(n9344), .B(p_input[240]), .Z(n8828) );
  XOR U8818 ( .A(n8831), .B(n8830), .Z(n8829) );
  NOR U8819 ( .A(n9346), .B(p_input[238]), .Z(n8830) );
  XOR U8820 ( .A(n8833), .B(n8832), .Z(n8831) );
  NOR U8821 ( .A(n9348), .B(p_input[236]), .Z(n8832) );
  XOR U8822 ( .A(n8835), .B(n8834), .Z(n8833) );
  NOR U8823 ( .A(n9350), .B(p_input[234]), .Z(n8834) );
  XOR U8824 ( .A(n8837), .B(n8836), .Z(n8835) );
  NOR U8825 ( .A(n9352), .B(p_input[232]), .Z(n8836) );
  XOR U8826 ( .A(n8839), .B(n8838), .Z(n8837) );
  NOR U8827 ( .A(n9354), .B(p_input[230]), .Z(n8838) );
  XOR U8828 ( .A(n8841), .B(n8840), .Z(n8839) );
  NOR U8829 ( .A(n9356), .B(p_input[228]), .Z(n8840) );
  XOR U8830 ( .A(n8843), .B(n8842), .Z(n8841) );
  NOR U8831 ( .A(n9358), .B(p_input[226]), .Z(n8842) );
  XOR U8832 ( .A(n8845), .B(n8844), .Z(n8843) );
  NOR U8833 ( .A(n9360), .B(p_input[224]), .Z(n8844) );
  XOR U8834 ( .A(n8847), .B(n8846), .Z(n8845) );
  NOR U8835 ( .A(n9362), .B(p_input[222]), .Z(n8846) );
  XOR U8836 ( .A(n8849), .B(n8848), .Z(n8847) );
  NOR U8837 ( .A(n9364), .B(p_input[220]), .Z(n8848) );
  XOR U8838 ( .A(n8851), .B(n8850), .Z(n8849) );
  NOR U8839 ( .A(n9366), .B(p_input[218]), .Z(n8850) );
  XOR U8840 ( .A(n8853), .B(n8852), .Z(n8851) );
  NOR U8841 ( .A(n9368), .B(p_input[216]), .Z(n8852) );
  XOR U8842 ( .A(n8855), .B(n8854), .Z(n8853) );
  NOR U8843 ( .A(n9370), .B(p_input[214]), .Z(n8854) );
  XOR U8844 ( .A(n8857), .B(n8856), .Z(n8855) );
  NOR U8845 ( .A(n9372), .B(p_input[212]), .Z(n8856) );
  XOR U8846 ( .A(n8859), .B(n8858), .Z(n8857) );
  NOR U8847 ( .A(n9374), .B(p_input[210]), .Z(n8858) );
  XOR U8848 ( .A(n8861), .B(n8860), .Z(n8859) );
  NOR U8849 ( .A(n9376), .B(p_input[208]), .Z(n8860) );
  XOR U8850 ( .A(n8863), .B(n8862), .Z(n8861) );
  NOR U8851 ( .A(n9378), .B(p_input[206]), .Z(n8862) );
  XOR U8852 ( .A(n8865), .B(n8864), .Z(n8863) );
  NOR U8853 ( .A(n9380), .B(p_input[204]), .Z(n8864) );
  XOR U8854 ( .A(n8867), .B(n8866), .Z(n8865) );
  NOR U8855 ( .A(n9382), .B(p_input[202]), .Z(n8866) );
  XOR U8856 ( .A(n8869), .B(n8868), .Z(n8867) );
  NOR U8857 ( .A(n9384), .B(p_input[200]), .Z(n8868) );
  XOR U8858 ( .A(n8871), .B(n8870), .Z(n8869) );
  NOR U8859 ( .A(n9386), .B(p_input[198]), .Z(n8870) );
  XOR U8860 ( .A(n8873), .B(n8872), .Z(n8871) );
  NOR U8861 ( .A(n9388), .B(p_input[196]), .Z(n8872) );
  XOR U8862 ( .A(n8875), .B(n8874), .Z(n8873) );
  NOR U8863 ( .A(n9390), .B(p_input[194]), .Z(n8874) );
  XOR U8864 ( .A(n8877), .B(n8876), .Z(n8875) );
  NOR U8865 ( .A(n9392), .B(p_input[192]), .Z(n8876) );
  XOR U8866 ( .A(n8879), .B(n8878), .Z(n8877) );
  NOR U8867 ( .A(n9394), .B(p_input[190]), .Z(n8878) );
  XOR U8868 ( .A(n8881), .B(n8880), .Z(n8879) );
  NOR U8869 ( .A(n9396), .B(p_input[188]), .Z(n8880) );
  XOR U8870 ( .A(n8883), .B(n8882), .Z(n8881) );
  NOR U8871 ( .A(n9398), .B(p_input[186]), .Z(n8882) );
  XOR U8872 ( .A(n8885), .B(n8884), .Z(n8883) );
  NOR U8873 ( .A(n9400), .B(p_input[184]), .Z(n8884) );
  XOR U8874 ( .A(n8887), .B(n8886), .Z(n8885) );
  NOR U8875 ( .A(n9402), .B(p_input[182]), .Z(n8886) );
  XOR U8876 ( .A(n8889), .B(n8888), .Z(n8887) );
  NOR U8877 ( .A(n9404), .B(p_input[180]), .Z(n8888) );
  XOR U8878 ( .A(n8891), .B(n8890), .Z(n8889) );
  NOR U8879 ( .A(n9406), .B(p_input[178]), .Z(n8890) );
  XOR U8880 ( .A(n8893), .B(n8892), .Z(n8891) );
  NOR U8881 ( .A(n9408), .B(p_input[176]), .Z(n8892) );
  XOR U8882 ( .A(n8895), .B(n8894), .Z(n8893) );
  NOR U8883 ( .A(n9410), .B(p_input[174]), .Z(n8894) );
  XOR U8884 ( .A(n8897), .B(n8896), .Z(n8895) );
  NOR U8885 ( .A(n9412), .B(p_input[172]), .Z(n8896) );
  XOR U8886 ( .A(n8899), .B(n8898), .Z(n8897) );
  NOR U8887 ( .A(n9414), .B(p_input[170]), .Z(n8898) );
  XOR U8888 ( .A(n8901), .B(n8900), .Z(n8899) );
  NOR U8889 ( .A(n9416), .B(p_input[168]), .Z(n8900) );
  XOR U8890 ( .A(n8903), .B(n8902), .Z(n8901) );
  NOR U8891 ( .A(n9418), .B(p_input[166]), .Z(n8902) );
  XOR U8892 ( .A(n8905), .B(n8904), .Z(n8903) );
  NOR U8893 ( .A(n9420), .B(p_input[164]), .Z(n8904) );
  XOR U8894 ( .A(n8907), .B(n8906), .Z(n8905) );
  NOR U8895 ( .A(n9422), .B(p_input[162]), .Z(n8906) );
  XOR U8896 ( .A(n8909), .B(n8908), .Z(n8907) );
  NOR U8897 ( .A(n9424), .B(p_input[160]), .Z(n8908) );
  XOR U8898 ( .A(n8911), .B(n8910), .Z(n8909) );
  NOR U8899 ( .A(n9426), .B(p_input[158]), .Z(n8910) );
  XOR U8900 ( .A(n8913), .B(n8912), .Z(n8911) );
  NOR U8901 ( .A(n9428), .B(p_input[156]), .Z(n8912) );
  XOR U8902 ( .A(n8915), .B(n8914), .Z(n8913) );
  NOR U8903 ( .A(n9430), .B(p_input[154]), .Z(n8914) );
  XOR U8904 ( .A(n8917), .B(n8916), .Z(n8915) );
  NOR U8905 ( .A(n9432), .B(p_input[152]), .Z(n8916) );
  XOR U8906 ( .A(n8919), .B(n8918), .Z(n8917) );
  NOR U8907 ( .A(n9434), .B(p_input[150]), .Z(n8918) );
  XOR U8908 ( .A(n8921), .B(n8920), .Z(n8919) );
  NOR U8909 ( .A(n9436), .B(p_input[148]), .Z(n8920) );
  XOR U8910 ( .A(n8923), .B(n8922), .Z(n8921) );
  NOR U8911 ( .A(n9438), .B(p_input[146]), .Z(n8922) );
  XOR U8912 ( .A(n8925), .B(n8924), .Z(n8923) );
  NOR U8913 ( .A(n9440), .B(p_input[144]), .Z(n8924) );
  XOR U8914 ( .A(n8927), .B(n8926), .Z(n8925) );
  NOR U8915 ( .A(n9442), .B(p_input[142]), .Z(n8926) );
  XOR U8916 ( .A(n8929), .B(n8928), .Z(n8927) );
  NOR U8917 ( .A(n9444), .B(p_input[140]), .Z(n8928) );
  XOR U8918 ( .A(n8931), .B(n8930), .Z(n8929) );
  NOR U8919 ( .A(n9446), .B(p_input[138]), .Z(n8930) );
  XOR U8920 ( .A(n8933), .B(n8932), .Z(n8931) );
  NOR U8921 ( .A(n9448), .B(p_input[136]), .Z(n8932) );
  XOR U8922 ( .A(n8935), .B(n8934), .Z(n8933) );
  NOR U8923 ( .A(n9450), .B(p_input[134]), .Z(n8934) );
  XOR U8924 ( .A(n8937), .B(n8936), .Z(n8935) );
  NOR U8925 ( .A(n9452), .B(p_input[132]), .Z(n8936) );
  XOR U8926 ( .A(n8939), .B(n8938), .Z(n8937) );
  NOR U8927 ( .A(n9454), .B(p_input[130]), .Z(n8938) );
  XOR U8928 ( .A(n8941), .B(n8940), .Z(n8939) );
  NOR U8929 ( .A(n9456), .B(p_input[128]), .Z(n8940) );
  XOR U8930 ( .A(n8943), .B(n8942), .Z(n8941) );
  NOR U8931 ( .A(n9458), .B(p_input[126]), .Z(n8942) );
  XOR U8932 ( .A(n8945), .B(n8944), .Z(n8943) );
  NOR U8933 ( .A(n9460), .B(p_input[124]), .Z(n8944) );
  XOR U8934 ( .A(n8947), .B(n8946), .Z(n8945) );
  NOR U8935 ( .A(n9462), .B(p_input[122]), .Z(n8946) );
  XOR U8936 ( .A(n8949), .B(n8948), .Z(n8947) );
  NOR U8937 ( .A(n9464), .B(p_input[120]), .Z(n8948) );
  XOR U8938 ( .A(n8951), .B(n8950), .Z(n8949) );
  NOR U8939 ( .A(n9466), .B(p_input[118]), .Z(n8950) );
  XOR U8940 ( .A(n8953), .B(n8952), .Z(n8951) );
  NOR U8941 ( .A(n9468), .B(p_input[116]), .Z(n8952) );
  XOR U8942 ( .A(n8955), .B(n8954), .Z(n8953) );
  NOR U8943 ( .A(n9470), .B(p_input[114]), .Z(n8954) );
  XOR U8944 ( .A(n8957), .B(n8956), .Z(n8955) );
  NOR U8945 ( .A(n9472), .B(p_input[112]), .Z(n8956) );
  XOR U8946 ( .A(n8959), .B(n8958), .Z(n8957) );
  NOR U8947 ( .A(n9474), .B(p_input[110]), .Z(n8958) );
  XOR U8948 ( .A(n8961), .B(n8960), .Z(n8959) );
  NOR U8949 ( .A(n9476), .B(p_input[108]), .Z(n8960) );
  XOR U8950 ( .A(n8963), .B(n8962), .Z(n8961) );
  NOR U8951 ( .A(n9478), .B(p_input[106]), .Z(n8962) );
  XOR U8952 ( .A(n8965), .B(n8964), .Z(n8963) );
  NOR U8953 ( .A(n9480), .B(p_input[104]), .Z(n8964) );
  XOR U8954 ( .A(n8967), .B(n8966), .Z(n8965) );
  NOR U8955 ( .A(n9482), .B(p_input[102]), .Z(n8966) );
  XOR U8956 ( .A(n8969), .B(n8968), .Z(n8967) );
  NOR U8957 ( .A(n9484), .B(p_input[100]), .Z(n8968) );
  XOR U8958 ( .A(n8971), .B(n8970), .Z(n8969) );
  NOR U8959 ( .A(n9486), .B(p_input[98]), .Z(n8970) );
  XOR U8960 ( .A(n8973), .B(n8972), .Z(n8971) );
  NOR U8961 ( .A(n9488), .B(p_input[96]), .Z(n8972) );
  XOR U8962 ( .A(n8975), .B(n8974), .Z(n8973) );
  NOR U8963 ( .A(n9490), .B(p_input[94]), .Z(n8974) );
  XOR U8964 ( .A(n8977), .B(n8976), .Z(n8975) );
  NOR U8965 ( .A(n9492), .B(p_input[92]), .Z(n8976) );
  XOR U8966 ( .A(n8979), .B(n8978), .Z(n8977) );
  NOR U8967 ( .A(n9494), .B(p_input[90]), .Z(n8978) );
  XOR U8968 ( .A(n8981), .B(n8980), .Z(n8979) );
  NOR U8969 ( .A(n9496), .B(p_input[88]), .Z(n8980) );
  XOR U8970 ( .A(n8983), .B(n8982), .Z(n8981) );
  NOR U8971 ( .A(n9498), .B(p_input[86]), .Z(n8982) );
  XOR U8972 ( .A(n8985), .B(n8984), .Z(n8983) );
  NOR U8973 ( .A(n9500), .B(p_input[84]), .Z(n8984) );
  XOR U8974 ( .A(n8987), .B(n8986), .Z(n8985) );
  NOR U8975 ( .A(n9502), .B(p_input[82]), .Z(n8986) );
  XOR U8976 ( .A(n8989), .B(n8988), .Z(n8987) );
  NOR U8977 ( .A(n9504), .B(p_input[80]), .Z(n8988) );
  XOR U8978 ( .A(n8991), .B(n8990), .Z(n8989) );
  NOR U8979 ( .A(n9506), .B(p_input[78]), .Z(n8990) );
  XOR U8980 ( .A(n8993), .B(n8992), .Z(n8991) );
  NOR U8981 ( .A(n9508), .B(p_input[76]), .Z(n8992) );
  XOR U8982 ( .A(n8995), .B(n8994), .Z(n8993) );
  NOR U8983 ( .A(n9510), .B(p_input[74]), .Z(n8994) );
  XOR U8984 ( .A(n8997), .B(n8996), .Z(n8995) );
  NOR U8985 ( .A(n9512), .B(p_input[72]), .Z(n8996) );
  XOR U8986 ( .A(n8999), .B(n8998), .Z(n8997) );
  NOR U8987 ( .A(n9514), .B(p_input[70]), .Z(n8998) );
  XOR U8988 ( .A(n9001), .B(n9000), .Z(n8999) );
  NOR U8989 ( .A(n9516), .B(p_input[68]), .Z(n9000) );
  XOR U8990 ( .A(n9003), .B(n9002), .Z(n9001) );
  NOR U8991 ( .A(n9518), .B(p_input[66]), .Z(n9002) );
  XOR U8992 ( .A(n9005), .B(n9004), .Z(n9003) );
  NOR U8993 ( .A(n9520), .B(p_input[64]), .Z(n9004) );
  XOR U8994 ( .A(n9007), .B(n9006), .Z(n9005) );
  NOR U8995 ( .A(n9522), .B(p_input[62]), .Z(n9006) );
  XOR U8996 ( .A(n9009), .B(n9008), .Z(n9007) );
  NOR U8997 ( .A(n9524), .B(p_input[60]), .Z(n9008) );
  XOR U8998 ( .A(n9011), .B(n9010), .Z(n9009) );
  NOR U8999 ( .A(n9526), .B(p_input[58]), .Z(n9010) );
  XOR U9000 ( .A(n9013), .B(n9012), .Z(n9011) );
  NOR U9001 ( .A(n9528), .B(p_input[56]), .Z(n9012) );
  XOR U9002 ( .A(n9015), .B(n9014), .Z(n9013) );
  NOR U9003 ( .A(n9530), .B(p_input[54]), .Z(n9014) );
  XOR U9004 ( .A(n9017), .B(n9016), .Z(n9015) );
  NOR U9005 ( .A(n9532), .B(p_input[52]), .Z(n9016) );
  XOR U9006 ( .A(n9019), .B(n9018), .Z(n9017) );
  NOR U9007 ( .A(n9534), .B(p_input[50]), .Z(n9018) );
  XOR U9008 ( .A(n9021), .B(n9020), .Z(n9019) );
  NOR U9009 ( .A(n9536), .B(p_input[48]), .Z(n9020) );
  XOR U9010 ( .A(n9023), .B(n9022), .Z(n9021) );
  NOR U9011 ( .A(n9538), .B(p_input[46]), .Z(n9022) );
  XOR U9012 ( .A(n9025), .B(n9024), .Z(n9023) );
  NOR U9013 ( .A(n9540), .B(p_input[44]), .Z(n9024) );
  XOR U9014 ( .A(n9027), .B(n9026), .Z(n9025) );
  NOR U9015 ( .A(n9542), .B(p_input[42]), .Z(n9026) );
  XOR U9016 ( .A(n9029), .B(n9028), .Z(n9027) );
  NOR U9017 ( .A(n9544), .B(p_input[40]), .Z(n9028) );
  XOR U9018 ( .A(n9031), .B(n9030), .Z(n9029) );
  NOR U9019 ( .A(n9546), .B(p_input[38]), .Z(n9030) );
  XOR U9020 ( .A(n9033), .B(n9032), .Z(n9031) );
  NOR U9021 ( .A(n9548), .B(p_input[36]), .Z(n9032) );
  XOR U9022 ( .A(n9035), .B(n9034), .Z(n9033) );
  NOR U9023 ( .A(n9550), .B(p_input[34]), .Z(n9034) );
  XOR U9024 ( .A(n9037), .B(n9036), .Z(n9035) );
  NOR U9025 ( .A(n9552), .B(p_input[32]), .Z(n9036) );
  XOR U9026 ( .A(n9039), .B(n9038), .Z(n9037) );
  NOR U9027 ( .A(n9554), .B(p_input[30]), .Z(n9038) );
  XOR U9028 ( .A(n9041), .B(n9040), .Z(n9039) );
  NOR U9029 ( .A(n9556), .B(p_input[28]), .Z(n9040) );
  XOR U9030 ( .A(n9043), .B(n9042), .Z(n9041) );
  NOR U9031 ( .A(n9558), .B(p_input[26]), .Z(n9042) );
  XOR U9032 ( .A(n9045), .B(n9044), .Z(n9043) );
  NOR U9033 ( .A(n9560), .B(p_input[24]), .Z(n9044) );
  XOR U9034 ( .A(n9047), .B(n9046), .Z(n9045) );
  NOR U9035 ( .A(n9562), .B(p_input[22]), .Z(n9046) );
  XOR U9036 ( .A(n9049), .B(n9048), .Z(n9047) );
  NOR U9037 ( .A(n9564), .B(p_input[20]), .Z(n9048) );
  XOR U9038 ( .A(n9051), .B(n9050), .Z(n9049) );
  NOR U9039 ( .A(n9566), .B(p_input[18]), .Z(n9050) );
  XOR U9040 ( .A(n9053), .B(n9052), .Z(n9051) );
  NOR U9041 ( .A(n9568), .B(p_input[16]), .Z(n9052) );
  XOR U9042 ( .A(n9055), .B(n9054), .Z(n9053) );
  NOR U9043 ( .A(n9570), .B(p_input[14]), .Z(n9054) );
  XOR U9044 ( .A(n9057), .B(n9056), .Z(n9055) );
  NOR U9045 ( .A(n9572), .B(p_input[12]), .Z(n9056) );
  XOR U9046 ( .A(n9071), .B(n9070), .Z(n9057) );
  NOR U9047 ( .A(n9574), .B(p_input[10]), .Z(n9070) );
  XOR U9048 ( .A(n9073), .B(n9072), .Z(n9071) );
  NOR U9049 ( .A(n9576), .B(p_input[8]), .Z(n9072) );
  XOR U9050 ( .A(n9061), .B(n9060), .Z(n9073) );
  NOR U9051 ( .A(n9578), .B(p_input[6]), .Z(n9060) );
  XOR U9052 ( .A(n9068), .B(n9069), .Z(n9061) );
  XOR U9053 ( .A(n9066), .B(n9067), .Z(n9069) );
  NOR U9054 ( .A(n9580), .B(p_input[2]), .Z(n9067) );
  NOR U9055 ( .A(n9582), .B(p_input[0]), .Z(n9066) );
  NOR U9056 ( .A(n9584), .B(p_input[4]), .Z(n9068) );
  XNOR U9057 ( .A(n9586), .B(n9587), .Z(n124) );
  AND U9058 ( .A(n1), .B(n9588), .Z(n9587) );
  XNOR U9059 ( .A(n9586), .B(n9589), .Z(n9588) );
  XNOR U9060 ( .A(n9590), .B(n9591), .Z(n1) );
  AND U9061 ( .A(n9592), .B(n9593), .Z(n9591) );
  XNOR U9062 ( .A(n9590), .B(n19), .Z(n9593) );
  XOR U9063 ( .A(n9594), .B(n9595), .Z(n19) );
  AND U9064 ( .A(n9596), .B(n9597), .Z(n9595) );
  XNOR U9065 ( .A(n34), .B(n9594), .Z(n9596) );
  XNOR U9066 ( .A(n9598), .B(n9599), .Z(n9594) );
  AND U9067 ( .A(n34), .B(n9598), .Z(n9599) );
  XOR U9068 ( .A(n16), .B(n9590), .Z(n9592) );
  IV U9069 ( .A(n20), .Z(n16) );
  XOR U9070 ( .A(n9600), .B(n9601), .Z(n20) );
  AND U9071 ( .A(n9602), .B(n9603), .Z(n9601) );
  XOR U9072 ( .A(n35), .B(n9600), .Z(n9602) );
  XOR U9073 ( .A(n9604), .B(n9605), .Z(n9600) );
  NOR U9074 ( .A(n31), .B(n9606), .Z(n9605) );
  IV U9075 ( .A(n9604), .Z(n9606) );
  XOR U9076 ( .A(n9607), .B(n9608), .Z(n9590) );
  AND U9077 ( .A(n9609), .B(n9610), .Z(n9608) );
  XOR U9078 ( .A(n9607), .B(n34), .Z(n9610) );
  XOR U9079 ( .A(n9598), .B(n9597), .Z(n34) );
  XNOR U9080 ( .A(n9611), .B(n9612), .Z(n9597) );
  XOR U9081 ( .A(n9613), .B(n9614), .Z(n9612) );
  XOR U9082 ( .A(n9615), .B(n9616), .Z(n9614) );
  NOR U9083 ( .A(n9617), .B(n9618), .Z(n9616) );
  NOR U9084 ( .A(n9619), .B(n9620), .Z(n9615) );
  NOR U9085 ( .A(n9621), .B(n9622), .Z(n9613) );
  XOR U9086 ( .A(n9623), .B(n9624), .Z(n9611) );
  XOR U9087 ( .A(n9625), .B(n9626), .Z(n9624) );
  XOR U9088 ( .A(n9627), .B(n9628), .Z(n9626) );
  XNOR U9089 ( .A(n9629), .B(n9630), .Z(n9628) );
  XOR U9090 ( .A(n9631), .B(n9632), .Z(n9630) );
  XOR U9091 ( .A(n9633), .B(n9634), .Z(n9632) );
  XOR U9092 ( .A(n9635), .B(n9636), .Z(n9634) );
  XOR U9093 ( .A(n9637), .B(n9638), .Z(n9633) );
  XOR U9094 ( .A(n9639), .B(n9640), .Z(n9638) );
  XOR U9095 ( .A(n9641), .B(n9642), .Z(n9640) );
  XOR U9096 ( .A(n9643), .B(n9644), .Z(n9642) );
  XOR U9097 ( .A(n9645), .B(n9646), .Z(n9644) );
  XNOR U9098 ( .A(n9647), .B(n9648), .Z(n9643) );
  XNOR U9099 ( .A(n9649), .B(n9650), .Z(n9648) );
  NOR U9100 ( .A(n9651), .B(n9646), .Z(n9649) );
  XOR U9101 ( .A(n9652), .B(n9653), .Z(n9641) );
  XOR U9102 ( .A(n9654), .B(n9655), .Z(n9653) );
  XNOR U9103 ( .A(n9656), .B(n9657), .Z(n9655) );
  XOR U9104 ( .A(n9658), .B(n9659), .Z(n9657) );
  XOR U9105 ( .A(n9660), .B(n9661), .Z(n9659) );
  XOR U9106 ( .A(n9662), .B(n9663), .Z(n9661) );
  XOR U9107 ( .A(n9664), .B(n9665), .Z(n9660) );
  XOR U9108 ( .A(n9666), .B(n9667), .Z(n9665) );
  XOR U9109 ( .A(n9668), .B(n9669), .Z(n9667) );
  XOR U9110 ( .A(n9670), .B(n9671), .Z(n9669) );
  XOR U9111 ( .A(n9672), .B(n9673), .Z(n9671) );
  XNOR U9112 ( .A(n9674), .B(n9675), .Z(n9670) );
  XNOR U9113 ( .A(n9676), .B(n9677), .Z(n9675) );
  NOR U9114 ( .A(n9678), .B(n9673), .Z(n9676) );
  XOR U9115 ( .A(n9679), .B(n9680), .Z(n9668) );
  XOR U9116 ( .A(n9681), .B(n9682), .Z(n9680) );
  XNOR U9117 ( .A(n9683), .B(n9684), .Z(n9682) );
  XOR U9118 ( .A(n9685), .B(n9686), .Z(n9684) );
  XOR U9119 ( .A(n9687), .B(n9688), .Z(n9686) );
  XOR U9120 ( .A(n9689), .B(n9690), .Z(n9688) );
  XOR U9121 ( .A(n9691), .B(n9692), .Z(n9687) );
  XOR U9122 ( .A(n9693), .B(n9694), .Z(n9692) );
  XOR U9123 ( .A(n9695), .B(n9696), .Z(n9694) );
  XOR U9124 ( .A(n9697), .B(n9698), .Z(n9696) );
  XOR U9125 ( .A(n9699), .B(n9700), .Z(n9698) );
  XNOR U9126 ( .A(n9701), .B(n9702), .Z(n9697) );
  XNOR U9127 ( .A(n9703), .B(n9704), .Z(n9702) );
  NOR U9128 ( .A(n9705), .B(n9700), .Z(n9703) );
  XOR U9129 ( .A(n9706), .B(n9707), .Z(n9695) );
  XOR U9130 ( .A(n9708), .B(n9709), .Z(n9707) );
  XNOR U9131 ( .A(n9710), .B(n9711), .Z(n9709) );
  XOR U9132 ( .A(n9712), .B(n9713), .Z(n9711) );
  XOR U9133 ( .A(n9714), .B(n9715), .Z(n9713) );
  XOR U9134 ( .A(n9716), .B(n9717), .Z(n9715) );
  XOR U9135 ( .A(n9718), .B(n9719), .Z(n9714) );
  XOR U9136 ( .A(n9720), .B(n9721), .Z(n9719) );
  XOR U9137 ( .A(n9722), .B(n9723), .Z(n9721) );
  XOR U9138 ( .A(n9724), .B(n9725), .Z(n9723) );
  XOR U9139 ( .A(n9726), .B(n9727), .Z(n9725) );
  XNOR U9140 ( .A(n9728), .B(n9729), .Z(n9724) );
  XNOR U9141 ( .A(n9730), .B(n9731), .Z(n9729) );
  NOR U9142 ( .A(n9732), .B(n9727), .Z(n9730) );
  XOR U9143 ( .A(n9733), .B(n9734), .Z(n9722) );
  XOR U9144 ( .A(n9735), .B(n9736), .Z(n9734) );
  XNOR U9145 ( .A(n9737), .B(n9738), .Z(n9736) );
  XOR U9146 ( .A(n9739), .B(n9740), .Z(n9738) );
  XOR U9147 ( .A(n9741), .B(n9742), .Z(n9740) );
  XOR U9148 ( .A(n9743), .B(n9744), .Z(n9742) );
  XOR U9149 ( .A(n9745), .B(n9746), .Z(n9741) );
  XOR U9150 ( .A(n9747), .B(n9748), .Z(n9746) );
  XOR U9151 ( .A(n9749), .B(n9750), .Z(n9748) );
  XOR U9152 ( .A(n9751), .B(n9752), .Z(n9750) );
  XOR U9153 ( .A(n9753), .B(n9754), .Z(n9752) );
  XNOR U9154 ( .A(n9755), .B(n9756), .Z(n9751) );
  XNOR U9155 ( .A(n9757), .B(n9758), .Z(n9756) );
  NOR U9156 ( .A(n9759), .B(n9754), .Z(n9757) );
  XOR U9157 ( .A(n9760), .B(n9761), .Z(n9749) );
  XOR U9158 ( .A(n9762), .B(n9763), .Z(n9761) );
  XNOR U9159 ( .A(n9764), .B(n9765), .Z(n9763) );
  XOR U9160 ( .A(n9766), .B(n9767), .Z(n9765) );
  XOR U9161 ( .A(n9768), .B(n9769), .Z(n9767) );
  XOR U9162 ( .A(n9770), .B(n9771), .Z(n9769) );
  XOR U9163 ( .A(n9772), .B(n9773), .Z(n9768) );
  XOR U9164 ( .A(n9774), .B(n9775), .Z(n9773) );
  XOR U9165 ( .A(n9776), .B(n9777), .Z(n9775) );
  XOR U9166 ( .A(n9778), .B(n9779), .Z(n9777) );
  XOR U9167 ( .A(n9780), .B(n9781), .Z(n9779) );
  XNOR U9168 ( .A(n9782), .B(n9783), .Z(n9778) );
  XNOR U9169 ( .A(n9784), .B(n9785), .Z(n9783) );
  NOR U9170 ( .A(n9786), .B(n9781), .Z(n9784) );
  XOR U9171 ( .A(n9787), .B(n9788), .Z(n9776) );
  XOR U9172 ( .A(n9789), .B(n9790), .Z(n9788) );
  XNOR U9173 ( .A(n9791), .B(n9792), .Z(n9790) );
  XOR U9174 ( .A(n9793), .B(n9794), .Z(n9792) );
  XOR U9175 ( .A(n9795), .B(n9796), .Z(n9794) );
  XOR U9176 ( .A(n9797), .B(n9798), .Z(n9796) );
  XOR U9177 ( .A(n9799), .B(n9800), .Z(n9795) );
  XOR U9178 ( .A(n9801), .B(n9802), .Z(n9800) );
  XOR U9179 ( .A(n9803), .B(n9804), .Z(n9802) );
  XOR U9180 ( .A(n9805), .B(n9806), .Z(n9804) );
  XOR U9181 ( .A(n9807), .B(n9808), .Z(n9806) );
  XNOR U9182 ( .A(n9809), .B(n9810), .Z(n9805) );
  XNOR U9183 ( .A(n9811), .B(n9812), .Z(n9810) );
  NOR U9184 ( .A(n9813), .B(n9808), .Z(n9811) );
  XOR U9185 ( .A(n9814), .B(n9815), .Z(n9803) );
  XOR U9186 ( .A(n9816), .B(n9817), .Z(n9815) );
  XNOR U9187 ( .A(n9818), .B(n9819), .Z(n9817) );
  XOR U9188 ( .A(n9820), .B(n9821), .Z(n9819) );
  XOR U9189 ( .A(n9822), .B(n9823), .Z(n9821) );
  XOR U9190 ( .A(n9824), .B(n9825), .Z(n9823) );
  XOR U9191 ( .A(n9826), .B(n9827), .Z(n9822) );
  XOR U9192 ( .A(n9828), .B(n9829), .Z(n9827) );
  XOR U9193 ( .A(n9830), .B(n9831), .Z(n9829) );
  XOR U9194 ( .A(n9832), .B(n9833), .Z(n9831) );
  XOR U9195 ( .A(n9834), .B(n9835), .Z(n9833) );
  XNOR U9196 ( .A(n9836), .B(n9837), .Z(n9832) );
  XNOR U9197 ( .A(n9838), .B(n9839), .Z(n9837) );
  NOR U9198 ( .A(n9840), .B(n9835), .Z(n9838) );
  XOR U9199 ( .A(n9841), .B(n9842), .Z(n9830) );
  XOR U9200 ( .A(n9843), .B(n9844), .Z(n9842) );
  XNOR U9201 ( .A(n9845), .B(n9846), .Z(n9844) );
  XOR U9202 ( .A(n9847), .B(n9848), .Z(n9846) );
  XOR U9203 ( .A(n9849), .B(n9850), .Z(n9848) );
  XOR U9204 ( .A(n9851), .B(n9852), .Z(n9850) );
  XOR U9205 ( .A(n9853), .B(n9854), .Z(n9849) );
  XOR U9206 ( .A(n9855), .B(n9856), .Z(n9854) );
  XOR U9207 ( .A(n9857), .B(n9858), .Z(n9856) );
  XOR U9208 ( .A(n9859), .B(n9860), .Z(n9858) );
  XOR U9209 ( .A(n9861), .B(n9862), .Z(n9860) );
  XNOR U9210 ( .A(n9863), .B(n9864), .Z(n9859) );
  XNOR U9211 ( .A(n9865), .B(n9866), .Z(n9864) );
  NOR U9212 ( .A(n9867), .B(n9862), .Z(n9865) );
  XOR U9213 ( .A(n9868), .B(n9869), .Z(n9857) );
  XOR U9214 ( .A(n9870), .B(n9871), .Z(n9869) );
  XNOR U9215 ( .A(n9872), .B(n9873), .Z(n9871) );
  XOR U9216 ( .A(n9874), .B(n9875), .Z(n9873) );
  XOR U9217 ( .A(n9876), .B(n9877), .Z(n9875) );
  XOR U9218 ( .A(n9878), .B(n9879), .Z(n9877) );
  XOR U9219 ( .A(n9880), .B(n9881), .Z(n9876) );
  XOR U9220 ( .A(n9882), .B(n9883), .Z(n9881) );
  XOR U9221 ( .A(n9884), .B(n9885), .Z(n9883) );
  XOR U9222 ( .A(n9886), .B(n9887), .Z(n9885) );
  XOR U9223 ( .A(n9888), .B(n9889), .Z(n9887) );
  XNOR U9224 ( .A(n9890), .B(n9891), .Z(n9886) );
  XNOR U9225 ( .A(n9892), .B(n9893), .Z(n9891) );
  NOR U9226 ( .A(n9894), .B(n9889), .Z(n9892) );
  XOR U9227 ( .A(n9895), .B(n9896), .Z(n9884) );
  XOR U9228 ( .A(n9897), .B(n9898), .Z(n9896) );
  XNOR U9229 ( .A(n9899), .B(n9900), .Z(n9898) );
  XOR U9230 ( .A(n9901), .B(n9902), .Z(n9897) );
  XOR U9231 ( .A(n9903), .B(n9904), .Z(n9895) );
  XOR U9232 ( .A(n9905), .B(n9906), .Z(n9904) );
  AND U9233 ( .A(n9907), .B(n9908), .Z(n9906) );
  XOR U9234 ( .A(n9900), .B(n9909), .Z(n9907) );
  XOR U9235 ( .A(n9910), .B(n9911), .Z(n9900) );
  AND U9236 ( .A(n9909), .B(n9910), .Z(n9911) );
  NOR U9237 ( .A(n9912), .B(n9901), .Z(n9905) );
  XOR U9238 ( .A(n9913), .B(n9914), .Z(n9903) );
  NOR U9239 ( .A(n9915), .B(n9902), .Z(n9914) );
  NOR U9240 ( .A(n9916), .B(n9899), .Z(n9913) );
  XOR U9241 ( .A(n9917), .B(n9918), .Z(n9882) );
  NOR U9242 ( .A(n9919), .B(n9893), .Z(n9918) );
  NOR U9243 ( .A(n9920), .B(n9890), .Z(n9917) );
  XOR U9244 ( .A(n9921), .B(n9922), .Z(n9880) );
  XOR U9245 ( .A(n9923), .B(n9924), .Z(n9922) );
  NOR U9246 ( .A(n9925), .B(n9888), .Z(n9924) );
  NOR U9247 ( .A(n9926), .B(n9927), .Z(n9923) );
  XOR U9248 ( .A(n9928), .B(n9929), .Z(n9921) );
  AND U9249 ( .A(n9930), .B(n9931), .Z(n9929) );
  NOR U9250 ( .A(n9932), .B(n9878), .Z(n9928) );
  XOR U9251 ( .A(n9933), .B(n9934), .Z(n9874) );
  XNOR U9252 ( .A(n9927), .B(n9931), .Z(n9934) );
  XOR U9253 ( .A(n9935), .B(n9936), .Z(n9933) );
  NOR U9254 ( .A(n9937), .B(n9879), .Z(n9936) );
  NOR U9255 ( .A(n9938), .B(n9939), .Z(n9935) );
  XOR U9256 ( .A(n9940), .B(n9941), .Z(n9870) );
  XOR U9257 ( .A(n9942), .B(n9943), .Z(n9868) );
  XNOR U9258 ( .A(n9944), .B(n9939), .Z(n9943) );
  NOR U9259 ( .A(n9945), .B(n9940), .Z(n9944) );
  XOR U9260 ( .A(n9946), .B(n9947), .Z(n9942) );
  NOR U9261 ( .A(n9948), .B(n9941), .Z(n9947) );
  NOR U9262 ( .A(n9949), .B(n9872), .Z(n9946) );
  XOR U9263 ( .A(n9950), .B(n9951), .Z(n9855) );
  NOR U9264 ( .A(n9952), .B(n9866), .Z(n9951) );
  NOR U9265 ( .A(n9953), .B(n9863), .Z(n9950) );
  XOR U9266 ( .A(n9954), .B(n9955), .Z(n9853) );
  XOR U9267 ( .A(n9956), .B(n9957), .Z(n9955) );
  NOR U9268 ( .A(n9958), .B(n9861), .Z(n9957) );
  NOR U9269 ( .A(n9959), .B(n9960), .Z(n9956) );
  XOR U9270 ( .A(n9961), .B(n9962), .Z(n9954) );
  AND U9271 ( .A(n9963), .B(n9964), .Z(n9962) );
  NOR U9272 ( .A(n9965), .B(n9851), .Z(n9961) );
  XOR U9273 ( .A(n9966), .B(n9967), .Z(n9847) );
  XNOR U9274 ( .A(n9960), .B(n9964), .Z(n9967) );
  XOR U9275 ( .A(n9968), .B(n9969), .Z(n9966) );
  NOR U9276 ( .A(n9970), .B(n9852), .Z(n9969) );
  NOR U9277 ( .A(n9971), .B(n9972), .Z(n9968) );
  XOR U9278 ( .A(n9973), .B(n9974), .Z(n9843) );
  XOR U9279 ( .A(n9975), .B(n9976), .Z(n9841) );
  XNOR U9280 ( .A(n9977), .B(n9972), .Z(n9976) );
  NOR U9281 ( .A(n9978), .B(n9973), .Z(n9977) );
  XOR U9282 ( .A(n9979), .B(n9980), .Z(n9975) );
  NOR U9283 ( .A(n9981), .B(n9974), .Z(n9980) );
  NOR U9284 ( .A(n9982), .B(n9845), .Z(n9979) );
  XOR U9285 ( .A(n9983), .B(n9984), .Z(n9828) );
  NOR U9286 ( .A(n9985), .B(n9839), .Z(n9984) );
  NOR U9287 ( .A(n9986), .B(n9836), .Z(n9983) );
  XOR U9288 ( .A(n9987), .B(n9988), .Z(n9826) );
  XOR U9289 ( .A(n9989), .B(n9990), .Z(n9988) );
  NOR U9290 ( .A(n9991), .B(n9834), .Z(n9990) );
  NOR U9291 ( .A(n9992), .B(n9993), .Z(n9989) );
  XOR U9292 ( .A(n9994), .B(n9995), .Z(n9987) );
  AND U9293 ( .A(n9996), .B(n9997), .Z(n9995) );
  NOR U9294 ( .A(n9998), .B(n9824), .Z(n9994) );
  XOR U9295 ( .A(n9999), .B(n10000), .Z(n9820) );
  XNOR U9296 ( .A(n9993), .B(n9997), .Z(n10000) );
  XOR U9297 ( .A(n10001), .B(n10002), .Z(n9999) );
  NOR U9298 ( .A(n10003), .B(n9825), .Z(n10002) );
  NOR U9299 ( .A(n10004), .B(n10005), .Z(n10001) );
  XOR U9300 ( .A(n10006), .B(n10007), .Z(n9816) );
  XOR U9301 ( .A(n10008), .B(n10009), .Z(n9814) );
  XNOR U9302 ( .A(n10010), .B(n10005), .Z(n10009) );
  NOR U9303 ( .A(n10011), .B(n10006), .Z(n10010) );
  XOR U9304 ( .A(n10012), .B(n10013), .Z(n10008) );
  NOR U9305 ( .A(n10014), .B(n10007), .Z(n10013) );
  NOR U9306 ( .A(n10015), .B(n9818), .Z(n10012) );
  XOR U9307 ( .A(n10016), .B(n10017), .Z(n9801) );
  NOR U9308 ( .A(n10018), .B(n9812), .Z(n10017) );
  NOR U9309 ( .A(n10019), .B(n9809), .Z(n10016) );
  XOR U9310 ( .A(n10020), .B(n10021), .Z(n9799) );
  XOR U9311 ( .A(n10022), .B(n10023), .Z(n10021) );
  NOR U9312 ( .A(n10024), .B(n9807), .Z(n10023) );
  NOR U9313 ( .A(n10025), .B(n10026), .Z(n10022) );
  XOR U9314 ( .A(n10027), .B(n10028), .Z(n10020) );
  AND U9315 ( .A(n10029), .B(n10030), .Z(n10028) );
  NOR U9316 ( .A(n10031), .B(n9797), .Z(n10027) );
  XOR U9317 ( .A(n10032), .B(n10033), .Z(n9793) );
  XNOR U9318 ( .A(n10026), .B(n10030), .Z(n10033) );
  XOR U9319 ( .A(n10034), .B(n10035), .Z(n10032) );
  NOR U9320 ( .A(n10036), .B(n9798), .Z(n10035) );
  NOR U9321 ( .A(n10037), .B(n10038), .Z(n10034) );
  XOR U9322 ( .A(n10039), .B(n10040), .Z(n9789) );
  XOR U9323 ( .A(n10041), .B(n10042), .Z(n9787) );
  XNOR U9324 ( .A(n10043), .B(n10038), .Z(n10042) );
  NOR U9325 ( .A(n10044), .B(n10039), .Z(n10043) );
  XOR U9326 ( .A(n10045), .B(n10046), .Z(n10041) );
  NOR U9327 ( .A(n10047), .B(n10040), .Z(n10046) );
  NOR U9328 ( .A(n10048), .B(n9791), .Z(n10045) );
  XOR U9329 ( .A(n10049), .B(n10050), .Z(n9774) );
  NOR U9330 ( .A(n10051), .B(n9785), .Z(n10050) );
  NOR U9331 ( .A(n10052), .B(n9782), .Z(n10049) );
  XOR U9332 ( .A(n10053), .B(n10054), .Z(n9772) );
  XOR U9333 ( .A(n10055), .B(n10056), .Z(n10054) );
  NOR U9334 ( .A(n10057), .B(n9780), .Z(n10056) );
  NOR U9335 ( .A(n10058), .B(n10059), .Z(n10055) );
  XOR U9336 ( .A(n10060), .B(n10061), .Z(n10053) );
  AND U9337 ( .A(n10062), .B(n10063), .Z(n10061) );
  NOR U9338 ( .A(n10064), .B(n9770), .Z(n10060) );
  XOR U9339 ( .A(n10065), .B(n10066), .Z(n9766) );
  XNOR U9340 ( .A(n10059), .B(n10063), .Z(n10066) );
  XOR U9341 ( .A(n10067), .B(n10068), .Z(n10065) );
  NOR U9342 ( .A(n10069), .B(n9771), .Z(n10068) );
  NOR U9343 ( .A(n10070), .B(n10071), .Z(n10067) );
  XOR U9344 ( .A(n10072), .B(n10073), .Z(n9762) );
  XOR U9345 ( .A(n10074), .B(n10075), .Z(n9760) );
  XNOR U9346 ( .A(n10076), .B(n10071), .Z(n10075) );
  NOR U9347 ( .A(n10077), .B(n10072), .Z(n10076) );
  XOR U9348 ( .A(n10078), .B(n10079), .Z(n10074) );
  NOR U9349 ( .A(n10080), .B(n10073), .Z(n10079) );
  NOR U9350 ( .A(n10081), .B(n9764), .Z(n10078) );
  XOR U9351 ( .A(n10082), .B(n10083), .Z(n9747) );
  NOR U9352 ( .A(n10084), .B(n9758), .Z(n10083) );
  NOR U9353 ( .A(n10085), .B(n9755), .Z(n10082) );
  XOR U9354 ( .A(n10086), .B(n10087), .Z(n9745) );
  XOR U9355 ( .A(n10088), .B(n10089), .Z(n10087) );
  NOR U9356 ( .A(n10090), .B(n9753), .Z(n10089) );
  NOR U9357 ( .A(n10091), .B(n10092), .Z(n10088) );
  XOR U9358 ( .A(n10093), .B(n10094), .Z(n10086) );
  AND U9359 ( .A(n10095), .B(n10096), .Z(n10094) );
  NOR U9360 ( .A(n10097), .B(n9743), .Z(n10093) );
  XOR U9361 ( .A(n10098), .B(n10099), .Z(n9739) );
  XNOR U9362 ( .A(n10092), .B(n10096), .Z(n10099) );
  XOR U9363 ( .A(n10100), .B(n10101), .Z(n10098) );
  NOR U9364 ( .A(n10102), .B(n9744), .Z(n10101) );
  NOR U9365 ( .A(n10103), .B(n10104), .Z(n10100) );
  XOR U9366 ( .A(n10105), .B(n10106), .Z(n9735) );
  XOR U9367 ( .A(n10107), .B(n10108), .Z(n9733) );
  XNOR U9368 ( .A(n10109), .B(n10104), .Z(n10108) );
  NOR U9369 ( .A(n10110), .B(n10105), .Z(n10109) );
  XOR U9370 ( .A(n10111), .B(n10112), .Z(n10107) );
  NOR U9371 ( .A(n10113), .B(n10106), .Z(n10112) );
  NOR U9372 ( .A(n10114), .B(n9737), .Z(n10111) );
  XOR U9373 ( .A(n10115), .B(n10116), .Z(n9720) );
  NOR U9374 ( .A(n10117), .B(n9731), .Z(n10116) );
  NOR U9375 ( .A(n10118), .B(n9728), .Z(n10115) );
  XOR U9376 ( .A(n10119), .B(n10120), .Z(n9718) );
  XOR U9377 ( .A(n10121), .B(n10122), .Z(n10120) );
  NOR U9378 ( .A(n10123), .B(n9726), .Z(n10122) );
  NOR U9379 ( .A(n10124), .B(n10125), .Z(n10121) );
  XOR U9380 ( .A(n10126), .B(n10127), .Z(n10119) );
  AND U9381 ( .A(n10128), .B(n10129), .Z(n10127) );
  NOR U9382 ( .A(n10130), .B(n9716), .Z(n10126) );
  XOR U9383 ( .A(n10131), .B(n10132), .Z(n9712) );
  XNOR U9384 ( .A(n10125), .B(n10129), .Z(n10132) );
  XOR U9385 ( .A(n10133), .B(n10134), .Z(n10131) );
  NOR U9386 ( .A(n10135), .B(n9717), .Z(n10134) );
  NOR U9387 ( .A(n10136), .B(n10137), .Z(n10133) );
  XOR U9388 ( .A(n10138), .B(n10139), .Z(n9708) );
  XOR U9389 ( .A(n10140), .B(n10141), .Z(n9706) );
  XNOR U9390 ( .A(n10142), .B(n10137), .Z(n10141) );
  NOR U9391 ( .A(n10143), .B(n10138), .Z(n10142) );
  XOR U9392 ( .A(n10144), .B(n10145), .Z(n10140) );
  NOR U9393 ( .A(n10146), .B(n10139), .Z(n10145) );
  NOR U9394 ( .A(n10147), .B(n9710), .Z(n10144) );
  XOR U9395 ( .A(n10148), .B(n10149), .Z(n9693) );
  NOR U9396 ( .A(n10150), .B(n9704), .Z(n10149) );
  NOR U9397 ( .A(n10151), .B(n9701), .Z(n10148) );
  XOR U9398 ( .A(n10152), .B(n10153), .Z(n9691) );
  XOR U9399 ( .A(n10154), .B(n10155), .Z(n10153) );
  NOR U9400 ( .A(n10156), .B(n9699), .Z(n10155) );
  NOR U9401 ( .A(n10157), .B(n10158), .Z(n10154) );
  XOR U9402 ( .A(n10159), .B(n10160), .Z(n10152) );
  AND U9403 ( .A(n10161), .B(n10162), .Z(n10160) );
  NOR U9404 ( .A(n10163), .B(n9689), .Z(n10159) );
  XOR U9405 ( .A(n10164), .B(n10165), .Z(n9685) );
  XNOR U9406 ( .A(n10158), .B(n10162), .Z(n10165) );
  XOR U9407 ( .A(n10166), .B(n10167), .Z(n10164) );
  NOR U9408 ( .A(n10168), .B(n9690), .Z(n10167) );
  NOR U9409 ( .A(n10169), .B(n10170), .Z(n10166) );
  XOR U9410 ( .A(n10171), .B(n10172), .Z(n9681) );
  XOR U9411 ( .A(n10173), .B(n10174), .Z(n9679) );
  XNOR U9412 ( .A(n10175), .B(n10170), .Z(n10174) );
  NOR U9413 ( .A(n10176), .B(n10171), .Z(n10175) );
  XOR U9414 ( .A(n10177), .B(n10178), .Z(n10173) );
  NOR U9415 ( .A(n10179), .B(n10172), .Z(n10178) );
  NOR U9416 ( .A(n10180), .B(n9683), .Z(n10177) );
  XOR U9417 ( .A(n10181), .B(n10182), .Z(n9666) );
  NOR U9418 ( .A(n10183), .B(n9677), .Z(n10182) );
  NOR U9419 ( .A(n10184), .B(n9674), .Z(n10181) );
  XOR U9420 ( .A(n10185), .B(n10186), .Z(n9664) );
  XOR U9421 ( .A(n10187), .B(n10188), .Z(n10186) );
  NOR U9422 ( .A(n10189), .B(n9672), .Z(n10188) );
  NOR U9423 ( .A(n10190), .B(n10191), .Z(n10187) );
  XOR U9424 ( .A(n10192), .B(n10193), .Z(n10185) );
  AND U9425 ( .A(n10194), .B(n10195), .Z(n10193) );
  NOR U9426 ( .A(n10196), .B(n9662), .Z(n10192) );
  XOR U9427 ( .A(n10197), .B(n10198), .Z(n9658) );
  XNOR U9428 ( .A(n10191), .B(n10195), .Z(n10198) );
  XOR U9429 ( .A(n10199), .B(n10200), .Z(n10197) );
  NOR U9430 ( .A(n10201), .B(n9663), .Z(n10200) );
  NOR U9431 ( .A(n10202), .B(n10203), .Z(n10199) );
  XOR U9432 ( .A(n10204), .B(n10205), .Z(n9654) );
  XOR U9433 ( .A(n10206), .B(n10207), .Z(n9652) );
  XNOR U9434 ( .A(n10208), .B(n10203), .Z(n10207) );
  NOR U9435 ( .A(n10209), .B(n10204), .Z(n10208) );
  XOR U9436 ( .A(n10210), .B(n10211), .Z(n10206) );
  NOR U9437 ( .A(n10212), .B(n10205), .Z(n10211) );
  NOR U9438 ( .A(n10213), .B(n9656), .Z(n10210) );
  XOR U9439 ( .A(n10214), .B(n10215), .Z(n9639) );
  NOR U9440 ( .A(n10216), .B(n9650), .Z(n10215) );
  NOR U9441 ( .A(n10217), .B(n9647), .Z(n10214) );
  XOR U9442 ( .A(n10218), .B(n10219), .Z(n9637) );
  XOR U9443 ( .A(n10220), .B(n10221), .Z(n10219) );
  NOR U9444 ( .A(n10222), .B(n9645), .Z(n10221) );
  NOR U9445 ( .A(n10223), .B(n10224), .Z(n10220) );
  XOR U9446 ( .A(n10225), .B(n10226), .Z(n10218) );
  AND U9447 ( .A(n10227), .B(n10228), .Z(n10226) );
  NOR U9448 ( .A(n10229), .B(n9635), .Z(n10225) );
  XOR U9449 ( .A(n10230), .B(n10231), .Z(n9631) );
  XNOR U9450 ( .A(n10224), .B(n10228), .Z(n10231) );
  XOR U9451 ( .A(n10232), .B(n10233), .Z(n10230) );
  NOR U9452 ( .A(n10234), .B(n9636), .Z(n10233) );
  NOR U9453 ( .A(n10235), .B(n10236), .Z(n10232) );
  XOR U9454 ( .A(n10237), .B(n10238), .Z(n9627) );
  XOR U9455 ( .A(n10239), .B(n10240), .Z(n9625) );
  XNOR U9456 ( .A(n10241), .B(n10236), .Z(n10240) );
  NOR U9457 ( .A(n10242), .B(n10237), .Z(n10241) );
  XOR U9458 ( .A(n10243), .B(n10244), .Z(n10239) );
  NOR U9459 ( .A(n10245), .B(n10238), .Z(n10244) );
  NOR U9460 ( .A(n10246), .B(n9629), .Z(n10243) );
  XOR U9461 ( .A(n10247), .B(n10248), .Z(n9623) );
  XNOR U9462 ( .A(n9618), .B(n10249), .Z(n10248) );
  XNOR U9463 ( .A(n10250), .B(n9622), .Z(n10249) );
  AND U9464 ( .A(n10251), .B(n10252), .Z(n10250) );
  XOR U9465 ( .A(n10252), .B(n9620), .Z(n10247) );
  XNOR U9466 ( .A(n10253), .B(n10254), .Z(n9598) );
  NOR U9467 ( .A(n49), .B(n10253), .Z(n10254) );
  XOR U9468 ( .A(n31), .B(n9607), .Z(n9609) );
  IV U9469 ( .A(n35), .Z(n31) );
  XOR U9470 ( .A(n9604), .B(n9603), .Z(n35) );
  XNOR U9471 ( .A(n10255), .B(n10256), .Z(n9603) );
  XOR U9472 ( .A(n10257), .B(n10258), .Z(n10256) );
  XNOR U9473 ( .A(n10259), .B(n10260), .Z(n10258) );
  NOR U9474 ( .A(n10261), .B(n10260), .Z(n10259) );
  XOR U9475 ( .A(n10262), .B(n10263), .Z(n10257) );
  NOR U9476 ( .A(n10264), .B(n10265), .Z(n10263) );
  AND U9477 ( .A(n10266), .B(n10267), .Z(n10262) );
  XOR U9478 ( .A(n10268), .B(n10269), .Z(n10255) );
  XOR U9479 ( .A(n10270), .B(n10271), .Z(n10269) );
  XOR U9480 ( .A(n10272), .B(n10273), .Z(n10271) );
  XOR U9481 ( .A(n10274), .B(n10275), .Z(n10273) );
  XNOR U9482 ( .A(n10276), .B(n10277), .Z(n10275) );
  NOR U9483 ( .A(n10278), .B(n10277), .Z(n10276) );
  XOR U9484 ( .A(n10279), .B(n10280), .Z(n10274) );
  XOR U9485 ( .A(n10281), .B(n10282), .Z(n10280) );
  XOR U9486 ( .A(n10283), .B(n10284), .Z(n10282) );
  XNOR U9487 ( .A(n10285), .B(n10286), .Z(n10284) );
  NOR U9488 ( .A(n10287), .B(n10286), .Z(n10285) );
  XOR U9489 ( .A(n10288), .B(n10289), .Z(n10283) );
  XOR U9490 ( .A(n10290), .B(n10291), .Z(n10289) );
  XOR U9491 ( .A(n10292), .B(n10293), .Z(n10291) );
  XNOR U9492 ( .A(n10294), .B(n10295), .Z(n10293) );
  NOR U9493 ( .A(n10296), .B(n10295), .Z(n10294) );
  XOR U9494 ( .A(n10297), .B(n10298), .Z(n10292) );
  XOR U9495 ( .A(n10299), .B(n10300), .Z(n10298) );
  XOR U9496 ( .A(n10301), .B(n10302), .Z(n10300) );
  XNOR U9497 ( .A(n10303), .B(n10304), .Z(n10302) );
  NOR U9498 ( .A(n10305), .B(n10304), .Z(n10303) );
  XOR U9499 ( .A(n10306), .B(n10307), .Z(n10301) );
  XOR U9500 ( .A(n10308), .B(n10309), .Z(n10307) );
  XOR U9501 ( .A(n10310), .B(n10311), .Z(n10309) );
  XNOR U9502 ( .A(n10312), .B(n10313), .Z(n10311) );
  NOR U9503 ( .A(n10314), .B(n10313), .Z(n10312) );
  XOR U9504 ( .A(n10315), .B(n10316), .Z(n10310) );
  XOR U9505 ( .A(n10317), .B(n10318), .Z(n10316) );
  XOR U9506 ( .A(n10319), .B(n10320), .Z(n10318) );
  XNOR U9507 ( .A(n10321), .B(n10322), .Z(n10320) );
  NOR U9508 ( .A(n10323), .B(n10322), .Z(n10321) );
  XOR U9509 ( .A(n10324), .B(n10325), .Z(n10319) );
  XOR U9510 ( .A(n10326), .B(n10327), .Z(n10325) );
  XOR U9511 ( .A(n10328), .B(n10329), .Z(n10327) );
  XNOR U9512 ( .A(n10330), .B(n10331), .Z(n10329) );
  NOR U9513 ( .A(n10332), .B(n10331), .Z(n10330) );
  XOR U9514 ( .A(n10333), .B(n10334), .Z(n10328) );
  XOR U9515 ( .A(n10335), .B(n10336), .Z(n10334) );
  XOR U9516 ( .A(n10337), .B(n10338), .Z(n10336) );
  XNOR U9517 ( .A(n10339), .B(n10340), .Z(n10338) );
  NOR U9518 ( .A(n10341), .B(n10340), .Z(n10339) );
  XOR U9519 ( .A(n10342), .B(n10343), .Z(n10337) );
  XOR U9520 ( .A(n10344), .B(n10345), .Z(n10343) );
  XOR U9521 ( .A(n10346), .B(n10347), .Z(n10345) );
  XNOR U9522 ( .A(n10348), .B(n10349), .Z(n10347) );
  NOR U9523 ( .A(n10350), .B(n10349), .Z(n10348) );
  XOR U9524 ( .A(n10351), .B(n10352), .Z(n10346) );
  XOR U9525 ( .A(n10353), .B(n10354), .Z(n10352) );
  XOR U9526 ( .A(n10355), .B(n10356), .Z(n10354) );
  XNOR U9527 ( .A(n10357), .B(n10358), .Z(n10356) );
  NOR U9528 ( .A(n10359), .B(n10358), .Z(n10357) );
  XOR U9529 ( .A(n10360), .B(n10361), .Z(n10355) );
  XOR U9530 ( .A(n10362), .B(n10363), .Z(n10361) );
  XOR U9531 ( .A(n10364), .B(n10365), .Z(n10363) );
  XNOR U9532 ( .A(n10366), .B(n10367), .Z(n10365) );
  NOR U9533 ( .A(n10368), .B(n10367), .Z(n10366) );
  XOR U9534 ( .A(n10369), .B(n10370), .Z(n10364) );
  XOR U9535 ( .A(n10371), .B(n10372), .Z(n10370) );
  XOR U9536 ( .A(n10373), .B(n10374), .Z(n10372) );
  XNOR U9537 ( .A(n10375), .B(n10376), .Z(n10374) );
  NOR U9538 ( .A(n10377), .B(n10376), .Z(n10375) );
  XOR U9539 ( .A(n10378), .B(n10379), .Z(n10373) );
  XOR U9540 ( .A(n10380), .B(n10381), .Z(n10379) );
  XOR U9541 ( .A(n10382), .B(n10383), .Z(n10381) );
  XNOR U9542 ( .A(n10384), .B(n10385), .Z(n10383) );
  NOR U9543 ( .A(n10386), .B(n10385), .Z(n10384) );
  XOR U9544 ( .A(n10387), .B(n10388), .Z(n10382) );
  XOR U9545 ( .A(n10389), .B(n10390), .Z(n10388) );
  XOR U9546 ( .A(n10391), .B(n10392), .Z(n10390) );
  XNOR U9547 ( .A(n10393), .B(n10394), .Z(n10392) );
  NOR U9548 ( .A(n10395), .B(n10394), .Z(n10393) );
  XOR U9549 ( .A(n10396), .B(n10397), .Z(n10391) );
  XOR U9550 ( .A(n10398), .B(n10399), .Z(n10397) );
  XOR U9551 ( .A(n10400), .B(n10401), .Z(n10399) );
  XNOR U9552 ( .A(n10402), .B(n10403), .Z(n10401) );
  NOR U9553 ( .A(n10404), .B(n10403), .Z(n10402) );
  XOR U9554 ( .A(n10405), .B(n10406), .Z(n10400) );
  XOR U9555 ( .A(n10407), .B(n10408), .Z(n10406) );
  XOR U9556 ( .A(n10409), .B(n10410), .Z(n10408) );
  XNOR U9557 ( .A(n10411), .B(n10412), .Z(n10410) );
  NOR U9558 ( .A(n10413), .B(n10412), .Z(n10411) );
  XOR U9559 ( .A(n10414), .B(n10415), .Z(n10409) );
  XOR U9560 ( .A(n10416), .B(n10417), .Z(n10415) );
  XOR U9561 ( .A(n10418), .B(n10419), .Z(n10417) );
  XNOR U9562 ( .A(n10420), .B(n10421), .Z(n10419) );
  NOR U9563 ( .A(n10422), .B(n10421), .Z(n10420) );
  XOR U9564 ( .A(n10423), .B(n10424), .Z(n10418) );
  XOR U9565 ( .A(n10425), .B(n10426), .Z(n10424) );
  XOR U9566 ( .A(n10427), .B(n10428), .Z(n10426) );
  XNOR U9567 ( .A(n10429), .B(n10430), .Z(n10428) );
  NOR U9568 ( .A(n10431), .B(n10430), .Z(n10429) );
  XOR U9569 ( .A(n10432), .B(n10433), .Z(n10427) );
  XOR U9570 ( .A(n10434), .B(n10435), .Z(n10433) );
  XOR U9571 ( .A(n10436), .B(n10437), .Z(n10435) );
  XNOR U9572 ( .A(n10438), .B(n10439), .Z(n10437) );
  NOR U9573 ( .A(n10440), .B(n10439), .Z(n10438) );
  XOR U9574 ( .A(n10441), .B(n10442), .Z(n10436) );
  XOR U9575 ( .A(n10443), .B(n10444), .Z(n10442) );
  XOR U9576 ( .A(n10445), .B(n10446), .Z(n10444) );
  XNOR U9577 ( .A(n10447), .B(n10448), .Z(n10446) );
  NOR U9578 ( .A(n10449), .B(n10448), .Z(n10447) );
  XOR U9579 ( .A(n10450), .B(n10451), .Z(n10445) );
  XOR U9580 ( .A(n10452), .B(n10453), .Z(n10451) );
  XOR U9581 ( .A(n10454), .B(n10455), .Z(n10453) );
  XNOR U9582 ( .A(n10456), .B(n10457), .Z(n10455) );
  NOR U9583 ( .A(n10458), .B(n10457), .Z(n10456) );
  XOR U9584 ( .A(n10459), .B(n10460), .Z(n10454) );
  XOR U9585 ( .A(n10461), .B(n10462), .Z(n10460) );
  XOR U9586 ( .A(n10463), .B(n10464), .Z(n10462) );
  XNOR U9587 ( .A(n10465), .B(n10466), .Z(n10464) );
  NOR U9588 ( .A(n10467), .B(n10466), .Z(n10465) );
  XOR U9589 ( .A(n10468), .B(n10469), .Z(n10463) );
  XOR U9590 ( .A(n10470), .B(n10471), .Z(n10469) );
  XOR U9591 ( .A(n10472), .B(n10473), .Z(n10471) );
  XNOR U9592 ( .A(n10474), .B(n10475), .Z(n10473) );
  NOR U9593 ( .A(n10476), .B(n10475), .Z(n10474) );
  XOR U9594 ( .A(n10477), .B(n10478), .Z(n10472) );
  XOR U9595 ( .A(n10479), .B(n10480), .Z(n10478) );
  XOR U9596 ( .A(n10481), .B(n10482), .Z(n10480) );
  XNOR U9597 ( .A(n10483), .B(n10484), .Z(n10482) );
  NOR U9598 ( .A(n10485), .B(n10484), .Z(n10483) );
  XOR U9599 ( .A(n10486), .B(n10487), .Z(n10481) );
  XOR U9600 ( .A(n10488), .B(n10489), .Z(n10487) );
  XOR U9601 ( .A(n10490), .B(n10491), .Z(n10489) );
  XNOR U9602 ( .A(n10492), .B(n10493), .Z(n10491) );
  NOR U9603 ( .A(n10494), .B(n10493), .Z(n10492) );
  XOR U9604 ( .A(n10495), .B(n10496), .Z(n10490) );
  XOR U9605 ( .A(n10497), .B(n10498), .Z(n10496) );
  XOR U9606 ( .A(n10499), .B(n10500), .Z(n10498) );
  XNOR U9607 ( .A(n10501), .B(n10502), .Z(n10500) );
  NOR U9608 ( .A(n10503), .B(n10502), .Z(n10501) );
  XOR U9609 ( .A(n10504), .B(n10505), .Z(n10499) );
  XOR U9610 ( .A(n10506), .B(n10507), .Z(n10505) );
  XOR U9611 ( .A(n10508), .B(n10509), .Z(n10507) );
  XNOR U9612 ( .A(n10510), .B(n10511), .Z(n10509) );
  NOR U9613 ( .A(n10512), .B(n10511), .Z(n10510) );
  XOR U9614 ( .A(n10513), .B(n10514), .Z(n10508) );
  XOR U9615 ( .A(n10515), .B(n10516), .Z(n10514) );
  XOR U9616 ( .A(n10517), .B(n10518), .Z(n10516) );
  XNOR U9617 ( .A(n10519), .B(n10520), .Z(n10518) );
  NOR U9618 ( .A(n10521), .B(n10520), .Z(n10519) );
  XOR U9619 ( .A(n10522), .B(n10523), .Z(n10517) );
  XOR U9620 ( .A(n10524), .B(n10525), .Z(n10523) );
  XOR U9621 ( .A(n10526), .B(n10527), .Z(n10525) );
  XNOR U9622 ( .A(n10528), .B(n10529), .Z(n10527) );
  NOR U9623 ( .A(n10530), .B(n10529), .Z(n10528) );
  XOR U9624 ( .A(n10531), .B(n10532), .Z(n10526) );
  XOR U9625 ( .A(n10533), .B(n10534), .Z(n10532) );
  XOR U9626 ( .A(n10535), .B(n10536), .Z(n10534) );
  XOR U9627 ( .A(n10537), .B(n10538), .Z(n10533) );
  XNOR U9628 ( .A(n10539), .B(n10540), .Z(n10538) );
  XOR U9629 ( .A(n10541), .B(n10542), .Z(n10540) );
  XOR U9630 ( .A(n10543), .B(n10544), .Z(n10542) );
  XNOR U9631 ( .A(n10545), .B(n10546), .Z(n10544) );
  XOR U9632 ( .A(n10547), .B(n10548), .Z(n10543) );
  XOR U9633 ( .A(n10549), .B(n10550), .Z(n10541) );
  XOR U9634 ( .A(n10551), .B(n10552), .Z(n10550) );
  AND U9635 ( .A(n10553), .B(n10554), .Z(n10552) );
  XOR U9636 ( .A(n10546), .B(n10555), .Z(n10553) );
  XOR U9637 ( .A(n10556), .B(n10557), .Z(n10546) );
  AND U9638 ( .A(n10555), .B(n10556), .Z(n10557) );
  NOR U9639 ( .A(n10558), .B(n10547), .Z(n10551) );
  XOR U9640 ( .A(n10559), .B(n10560), .Z(n10549) );
  NOR U9641 ( .A(n10561), .B(n10548), .Z(n10560) );
  NOR U9642 ( .A(n10562), .B(n10545), .Z(n10559) );
  XNOR U9643 ( .A(n10563), .B(n10564), .Z(n10537) );
  XNOR U9644 ( .A(n10565), .B(n10566), .Z(n10564) );
  NOR U9645 ( .A(n10567), .B(n10539), .Z(n10565) );
  XOR U9646 ( .A(n10568), .B(n10569), .Z(n10531) );
  XOR U9647 ( .A(n10570), .B(n10571), .Z(n10569) );
  NOR U9648 ( .A(n10572), .B(n10535), .Z(n10571) );
  NOR U9649 ( .A(n10573), .B(n10566), .Z(n10570) );
  XOR U9650 ( .A(n10574), .B(n10575), .Z(n10568) );
  NOR U9651 ( .A(n10576), .B(n10563), .Z(n10575) );
  NOR U9652 ( .A(n10577), .B(n10536), .Z(n10574) );
  XOR U9653 ( .A(n10578), .B(n10579), .Z(n10524) );
  XOR U9654 ( .A(n10580), .B(n10581), .Z(n10522) );
  XNOR U9655 ( .A(n10582), .B(n10583), .Z(n10581) );
  NOR U9656 ( .A(n10584), .B(n10583), .Z(n10582) );
  XOR U9657 ( .A(n10585), .B(n10586), .Z(n10580) );
  NOR U9658 ( .A(n10587), .B(n10578), .Z(n10586) );
  NOR U9659 ( .A(n10588), .B(n10579), .Z(n10585) );
  XOR U9660 ( .A(n10589), .B(n10590), .Z(n10515) );
  XOR U9661 ( .A(n10591), .B(n10592), .Z(n10513) );
  XNOR U9662 ( .A(n10593), .B(n10594), .Z(n10592) );
  NOR U9663 ( .A(n10595), .B(n10594), .Z(n10593) );
  XOR U9664 ( .A(n10596), .B(n10597), .Z(n10591) );
  NOR U9665 ( .A(n10598), .B(n10589), .Z(n10597) );
  NOR U9666 ( .A(n10599), .B(n10590), .Z(n10596) );
  XOR U9667 ( .A(n10600), .B(n10601), .Z(n10506) );
  XOR U9668 ( .A(n10602), .B(n10603), .Z(n10504) );
  XNOR U9669 ( .A(n10604), .B(n10605), .Z(n10603) );
  NOR U9670 ( .A(n10606), .B(n10605), .Z(n10604) );
  XOR U9671 ( .A(n10607), .B(n10608), .Z(n10602) );
  NOR U9672 ( .A(n10609), .B(n10600), .Z(n10608) );
  NOR U9673 ( .A(n10610), .B(n10601), .Z(n10607) );
  XOR U9674 ( .A(n10611), .B(n10612), .Z(n10497) );
  XOR U9675 ( .A(n10613), .B(n10614), .Z(n10495) );
  XNOR U9676 ( .A(n10615), .B(n10616), .Z(n10614) );
  NOR U9677 ( .A(n10617), .B(n10616), .Z(n10615) );
  XOR U9678 ( .A(n10618), .B(n10619), .Z(n10613) );
  NOR U9679 ( .A(n10620), .B(n10611), .Z(n10619) );
  NOR U9680 ( .A(n10621), .B(n10612), .Z(n10618) );
  XOR U9681 ( .A(n10622), .B(n10623), .Z(n10488) );
  XOR U9682 ( .A(n10624), .B(n10625), .Z(n10486) );
  XNOR U9683 ( .A(n10626), .B(n10627), .Z(n10625) );
  NOR U9684 ( .A(n10628), .B(n10627), .Z(n10626) );
  XOR U9685 ( .A(n10629), .B(n10630), .Z(n10624) );
  NOR U9686 ( .A(n10631), .B(n10622), .Z(n10630) );
  NOR U9687 ( .A(n10632), .B(n10623), .Z(n10629) );
  XOR U9688 ( .A(n10633), .B(n10634), .Z(n10479) );
  XOR U9689 ( .A(n10635), .B(n10636), .Z(n10477) );
  XNOR U9690 ( .A(n10637), .B(n10638), .Z(n10636) );
  NOR U9691 ( .A(n10639), .B(n10638), .Z(n10637) );
  XOR U9692 ( .A(n10640), .B(n10641), .Z(n10635) );
  NOR U9693 ( .A(n10642), .B(n10633), .Z(n10641) );
  NOR U9694 ( .A(n10643), .B(n10634), .Z(n10640) );
  XOR U9695 ( .A(n10644), .B(n10645), .Z(n10470) );
  XOR U9696 ( .A(n10646), .B(n10647), .Z(n10468) );
  XNOR U9697 ( .A(n10648), .B(n10649), .Z(n10647) );
  NOR U9698 ( .A(n10650), .B(n10649), .Z(n10648) );
  XOR U9699 ( .A(n10651), .B(n10652), .Z(n10646) );
  NOR U9700 ( .A(n10653), .B(n10644), .Z(n10652) );
  NOR U9701 ( .A(n10654), .B(n10645), .Z(n10651) );
  XOR U9702 ( .A(n10655), .B(n10656), .Z(n10461) );
  XOR U9703 ( .A(n10657), .B(n10658), .Z(n10459) );
  XNOR U9704 ( .A(n10659), .B(n10660), .Z(n10658) );
  NOR U9705 ( .A(n10661), .B(n10660), .Z(n10659) );
  XOR U9706 ( .A(n10662), .B(n10663), .Z(n10657) );
  NOR U9707 ( .A(n10664), .B(n10655), .Z(n10663) );
  NOR U9708 ( .A(n10665), .B(n10656), .Z(n10662) );
  XOR U9709 ( .A(n10666), .B(n10667), .Z(n10452) );
  XOR U9710 ( .A(n10668), .B(n10669), .Z(n10450) );
  XNOR U9711 ( .A(n10670), .B(n10671), .Z(n10669) );
  NOR U9712 ( .A(n10672), .B(n10671), .Z(n10670) );
  XOR U9713 ( .A(n10673), .B(n10674), .Z(n10668) );
  NOR U9714 ( .A(n10675), .B(n10666), .Z(n10674) );
  NOR U9715 ( .A(n10676), .B(n10667), .Z(n10673) );
  XOR U9716 ( .A(n10677), .B(n10678), .Z(n10443) );
  XOR U9717 ( .A(n10679), .B(n10680), .Z(n10441) );
  XNOR U9718 ( .A(n10681), .B(n10682), .Z(n10680) );
  NOR U9719 ( .A(n10683), .B(n10682), .Z(n10681) );
  XOR U9720 ( .A(n10684), .B(n10685), .Z(n10679) );
  NOR U9721 ( .A(n10686), .B(n10677), .Z(n10685) );
  NOR U9722 ( .A(n10687), .B(n10678), .Z(n10684) );
  XOR U9723 ( .A(n10688), .B(n10689), .Z(n10434) );
  XOR U9724 ( .A(n10690), .B(n10691), .Z(n10432) );
  XNOR U9725 ( .A(n10692), .B(n10693), .Z(n10691) );
  NOR U9726 ( .A(n10694), .B(n10693), .Z(n10692) );
  XOR U9727 ( .A(n10695), .B(n10696), .Z(n10690) );
  NOR U9728 ( .A(n10697), .B(n10688), .Z(n10696) );
  NOR U9729 ( .A(n10698), .B(n10689), .Z(n10695) );
  XOR U9730 ( .A(n10699), .B(n10700), .Z(n10425) );
  XOR U9731 ( .A(n10701), .B(n10702), .Z(n10423) );
  XNOR U9732 ( .A(n10703), .B(n10704), .Z(n10702) );
  NOR U9733 ( .A(n10705), .B(n10704), .Z(n10703) );
  XOR U9734 ( .A(n10706), .B(n10707), .Z(n10701) );
  NOR U9735 ( .A(n10708), .B(n10699), .Z(n10707) );
  NOR U9736 ( .A(n10709), .B(n10700), .Z(n10706) );
  XOR U9737 ( .A(n10710), .B(n10711), .Z(n10416) );
  XOR U9738 ( .A(n10712), .B(n10713), .Z(n10414) );
  XNOR U9739 ( .A(n10714), .B(n10715), .Z(n10713) );
  NOR U9740 ( .A(n10716), .B(n10715), .Z(n10714) );
  XOR U9741 ( .A(n10717), .B(n10718), .Z(n10712) );
  NOR U9742 ( .A(n10719), .B(n10710), .Z(n10718) );
  NOR U9743 ( .A(n10720), .B(n10711), .Z(n10717) );
  XOR U9744 ( .A(n10721), .B(n10722), .Z(n10407) );
  XOR U9745 ( .A(n10723), .B(n10724), .Z(n10405) );
  XNOR U9746 ( .A(n10725), .B(n10726), .Z(n10724) );
  NOR U9747 ( .A(n10727), .B(n10726), .Z(n10725) );
  XOR U9748 ( .A(n10728), .B(n10729), .Z(n10723) );
  NOR U9749 ( .A(n10730), .B(n10721), .Z(n10729) );
  NOR U9750 ( .A(n10731), .B(n10722), .Z(n10728) );
  XOR U9751 ( .A(n10732), .B(n10733), .Z(n10398) );
  XOR U9752 ( .A(n10734), .B(n10735), .Z(n10396) );
  XNOR U9753 ( .A(n10736), .B(n10737), .Z(n10735) );
  NOR U9754 ( .A(n10738), .B(n10737), .Z(n10736) );
  XOR U9755 ( .A(n10739), .B(n10740), .Z(n10734) );
  NOR U9756 ( .A(n10741), .B(n10732), .Z(n10740) );
  NOR U9757 ( .A(n10742), .B(n10733), .Z(n10739) );
  XOR U9758 ( .A(n10743), .B(n10744), .Z(n10389) );
  XOR U9759 ( .A(n10745), .B(n10746), .Z(n10387) );
  XNOR U9760 ( .A(n10747), .B(n10748), .Z(n10746) );
  NOR U9761 ( .A(n10749), .B(n10748), .Z(n10747) );
  XOR U9762 ( .A(n10750), .B(n10751), .Z(n10745) );
  NOR U9763 ( .A(n10752), .B(n10743), .Z(n10751) );
  NOR U9764 ( .A(n10753), .B(n10744), .Z(n10750) );
  XOR U9765 ( .A(n10754), .B(n10755), .Z(n10380) );
  XOR U9766 ( .A(n10756), .B(n10757), .Z(n10378) );
  XNOR U9767 ( .A(n10758), .B(n10759), .Z(n10757) );
  NOR U9768 ( .A(n10760), .B(n10759), .Z(n10758) );
  XOR U9769 ( .A(n10761), .B(n10762), .Z(n10756) );
  NOR U9770 ( .A(n10763), .B(n10754), .Z(n10762) );
  NOR U9771 ( .A(n10764), .B(n10755), .Z(n10761) );
  XOR U9772 ( .A(n10765), .B(n10766), .Z(n10371) );
  XOR U9773 ( .A(n10767), .B(n10768), .Z(n10369) );
  XNOR U9774 ( .A(n10769), .B(n10770), .Z(n10768) );
  NOR U9775 ( .A(n10771), .B(n10770), .Z(n10769) );
  XOR U9776 ( .A(n10772), .B(n10773), .Z(n10767) );
  NOR U9777 ( .A(n10774), .B(n10765), .Z(n10773) );
  NOR U9778 ( .A(n10775), .B(n10766), .Z(n10772) );
  XOR U9779 ( .A(n10776), .B(n10777), .Z(n10362) );
  XOR U9780 ( .A(n10778), .B(n10779), .Z(n10360) );
  XNOR U9781 ( .A(n10780), .B(n10781), .Z(n10779) );
  NOR U9782 ( .A(n10782), .B(n10781), .Z(n10780) );
  XOR U9783 ( .A(n10783), .B(n10784), .Z(n10778) );
  NOR U9784 ( .A(n10785), .B(n10776), .Z(n10784) );
  NOR U9785 ( .A(n10786), .B(n10777), .Z(n10783) );
  XOR U9786 ( .A(n10787), .B(n10788), .Z(n10353) );
  XOR U9787 ( .A(n10789), .B(n10790), .Z(n10351) );
  XNOR U9788 ( .A(n10791), .B(n10792), .Z(n10790) );
  NOR U9789 ( .A(n10793), .B(n10792), .Z(n10791) );
  XOR U9790 ( .A(n10794), .B(n10795), .Z(n10789) );
  NOR U9791 ( .A(n10796), .B(n10787), .Z(n10795) );
  NOR U9792 ( .A(n10797), .B(n10788), .Z(n10794) );
  XOR U9793 ( .A(n10798), .B(n10799), .Z(n10344) );
  XOR U9794 ( .A(n10800), .B(n10801), .Z(n10342) );
  XNOR U9795 ( .A(n10802), .B(n10803), .Z(n10801) );
  NOR U9796 ( .A(n10804), .B(n10803), .Z(n10802) );
  XOR U9797 ( .A(n10805), .B(n10806), .Z(n10800) );
  NOR U9798 ( .A(n10807), .B(n10798), .Z(n10806) );
  NOR U9799 ( .A(n10808), .B(n10799), .Z(n10805) );
  XOR U9800 ( .A(n10809), .B(n10810), .Z(n10335) );
  XOR U9801 ( .A(n10811), .B(n10812), .Z(n10333) );
  XNOR U9802 ( .A(n10813), .B(n10814), .Z(n10812) );
  NOR U9803 ( .A(n10815), .B(n10814), .Z(n10813) );
  XOR U9804 ( .A(n10816), .B(n10817), .Z(n10811) );
  NOR U9805 ( .A(n10818), .B(n10809), .Z(n10817) );
  NOR U9806 ( .A(n10819), .B(n10810), .Z(n10816) );
  XOR U9807 ( .A(n10820), .B(n10821), .Z(n10326) );
  XOR U9808 ( .A(n10822), .B(n10823), .Z(n10324) );
  XNOR U9809 ( .A(n10824), .B(n10825), .Z(n10823) );
  NOR U9810 ( .A(n10826), .B(n10825), .Z(n10824) );
  XOR U9811 ( .A(n10827), .B(n10828), .Z(n10822) );
  NOR U9812 ( .A(n10829), .B(n10820), .Z(n10828) );
  NOR U9813 ( .A(n10830), .B(n10821), .Z(n10827) );
  XOR U9814 ( .A(n10831), .B(n10832), .Z(n10317) );
  XOR U9815 ( .A(n10833), .B(n10834), .Z(n10315) );
  XNOR U9816 ( .A(n10835), .B(n10836), .Z(n10834) );
  NOR U9817 ( .A(n10837), .B(n10836), .Z(n10835) );
  XOR U9818 ( .A(n10838), .B(n10839), .Z(n10833) );
  NOR U9819 ( .A(n10840), .B(n10831), .Z(n10839) );
  NOR U9820 ( .A(n10841), .B(n10832), .Z(n10838) );
  XOR U9821 ( .A(n10842), .B(n10843), .Z(n10308) );
  XOR U9822 ( .A(n10844), .B(n10845), .Z(n10306) );
  XNOR U9823 ( .A(n10846), .B(n10847), .Z(n10845) );
  NOR U9824 ( .A(n10848), .B(n10847), .Z(n10846) );
  XOR U9825 ( .A(n10849), .B(n10850), .Z(n10844) );
  NOR U9826 ( .A(n10851), .B(n10842), .Z(n10850) );
  NOR U9827 ( .A(n10852), .B(n10843), .Z(n10849) );
  XOR U9828 ( .A(n10853), .B(n10854), .Z(n10299) );
  XOR U9829 ( .A(n10855), .B(n10856), .Z(n10297) );
  XNOR U9830 ( .A(n10857), .B(n10858), .Z(n10856) );
  NOR U9831 ( .A(n10859), .B(n10858), .Z(n10857) );
  XOR U9832 ( .A(n10860), .B(n10861), .Z(n10855) );
  NOR U9833 ( .A(n10862), .B(n10853), .Z(n10861) );
  NOR U9834 ( .A(n10863), .B(n10854), .Z(n10860) );
  XOR U9835 ( .A(n10864), .B(n10865), .Z(n10290) );
  XOR U9836 ( .A(n10866), .B(n10867), .Z(n10288) );
  XNOR U9837 ( .A(n10868), .B(n10869), .Z(n10867) );
  NOR U9838 ( .A(n10870), .B(n10869), .Z(n10868) );
  XOR U9839 ( .A(n10871), .B(n10872), .Z(n10866) );
  NOR U9840 ( .A(n10873), .B(n10864), .Z(n10872) );
  NOR U9841 ( .A(n10874), .B(n10865), .Z(n10871) );
  XOR U9842 ( .A(n10875), .B(n10876), .Z(n10281) );
  XOR U9843 ( .A(n10877), .B(n10878), .Z(n10279) );
  XNOR U9844 ( .A(n10879), .B(n10880), .Z(n10878) );
  NOR U9845 ( .A(n10881), .B(n10880), .Z(n10879) );
  XOR U9846 ( .A(n10882), .B(n10883), .Z(n10877) );
  NOR U9847 ( .A(n10884), .B(n10875), .Z(n10883) );
  NOR U9848 ( .A(n10885), .B(n10876), .Z(n10882) );
  XOR U9849 ( .A(n10886), .B(n10887), .Z(n10272) );
  XOR U9850 ( .A(n10888), .B(n10889), .Z(n10270) );
  XNOR U9851 ( .A(n10890), .B(n10891), .Z(n10889) );
  NOR U9852 ( .A(n10892), .B(n10891), .Z(n10890) );
  XOR U9853 ( .A(n10893), .B(n10894), .Z(n10888) );
  NOR U9854 ( .A(n10895), .B(n10886), .Z(n10894) );
  NOR U9855 ( .A(n10896), .B(n10887), .Z(n10893) );
  XOR U9856 ( .A(n10267), .B(n10265), .Z(n10268) );
  XOR U9857 ( .A(n10897), .B(n10898), .Z(n9604) );
  AND U9858 ( .A(n47), .B(n10897), .Z(n10898) );
  XOR U9859 ( .A(n10899), .B(n10900), .Z(n9607) );
  AND U9860 ( .A(n10901), .B(n10902), .Z(n10900) );
  XNOR U9861 ( .A(n49), .B(n10899), .Z(n10902) );
  XOR U9862 ( .A(n10253), .B(n10251), .Z(n49) );
  XOR U9863 ( .A(n10903), .B(n9619), .Z(n10251) );
  XNOR U9864 ( .A(n9620), .B(n9617), .Z(n9619) );
  XNOR U9865 ( .A(n9618), .B(n9621), .Z(n9617) );
  XNOR U9866 ( .A(n9622), .B(n10246), .Z(n9621) );
  XNOR U9867 ( .A(n9629), .B(n10245), .Z(n10246) );
  XNOR U9868 ( .A(n10238), .B(n10242), .Z(n10245) );
  XNOR U9869 ( .A(n10237), .B(n10235), .Z(n10242) );
  XNOR U9870 ( .A(n10236), .B(n10234), .Z(n10235) );
  XNOR U9871 ( .A(n9636), .B(n10229), .Z(n10234) );
  XOR U9872 ( .A(n9635), .B(n10227), .Z(n10229) );
  XNOR U9873 ( .A(n10228), .B(n10223), .Z(n10227) );
  XNOR U9874 ( .A(n10224), .B(n9651), .Z(n10223) );
  XNOR U9875 ( .A(n9646), .B(n10222), .Z(n9651) );
  XNOR U9876 ( .A(n9645), .B(n10217), .Z(n10222) );
  XNOR U9877 ( .A(n9647), .B(n10216), .Z(n10217) );
  XNOR U9878 ( .A(n9650), .B(n10213), .Z(n10216) );
  XNOR U9879 ( .A(n9656), .B(n10212), .Z(n10213) );
  XNOR U9880 ( .A(n10205), .B(n10209), .Z(n10212) );
  XNOR U9881 ( .A(n10204), .B(n10202), .Z(n10209) );
  XNOR U9882 ( .A(n10203), .B(n10201), .Z(n10202) );
  XNOR U9883 ( .A(n9663), .B(n10196), .Z(n10201) );
  XOR U9884 ( .A(n9662), .B(n10194), .Z(n10196) );
  XNOR U9885 ( .A(n10195), .B(n10190), .Z(n10194) );
  XNOR U9886 ( .A(n10191), .B(n9678), .Z(n10190) );
  XNOR U9887 ( .A(n9673), .B(n10189), .Z(n9678) );
  XNOR U9888 ( .A(n9672), .B(n10184), .Z(n10189) );
  XNOR U9889 ( .A(n9674), .B(n10183), .Z(n10184) );
  XNOR U9890 ( .A(n9677), .B(n10180), .Z(n10183) );
  XNOR U9891 ( .A(n9683), .B(n10179), .Z(n10180) );
  XNOR U9892 ( .A(n10172), .B(n10176), .Z(n10179) );
  XNOR U9893 ( .A(n10171), .B(n10169), .Z(n10176) );
  XNOR U9894 ( .A(n10170), .B(n10168), .Z(n10169) );
  XNOR U9895 ( .A(n9690), .B(n10163), .Z(n10168) );
  XOR U9896 ( .A(n9689), .B(n10161), .Z(n10163) );
  XNOR U9897 ( .A(n10162), .B(n10157), .Z(n10161) );
  XNOR U9898 ( .A(n10158), .B(n9705), .Z(n10157) );
  XNOR U9899 ( .A(n9700), .B(n10156), .Z(n9705) );
  XNOR U9900 ( .A(n9699), .B(n10151), .Z(n10156) );
  XNOR U9901 ( .A(n9701), .B(n10150), .Z(n10151) );
  XNOR U9902 ( .A(n9704), .B(n10147), .Z(n10150) );
  XNOR U9903 ( .A(n9710), .B(n10146), .Z(n10147) );
  XNOR U9904 ( .A(n10139), .B(n10143), .Z(n10146) );
  XNOR U9905 ( .A(n10138), .B(n10136), .Z(n10143) );
  XNOR U9906 ( .A(n10137), .B(n10135), .Z(n10136) );
  XNOR U9907 ( .A(n9717), .B(n10130), .Z(n10135) );
  XOR U9908 ( .A(n9716), .B(n10128), .Z(n10130) );
  XNOR U9909 ( .A(n10129), .B(n10124), .Z(n10128) );
  XNOR U9910 ( .A(n10125), .B(n9732), .Z(n10124) );
  XNOR U9911 ( .A(n9727), .B(n10123), .Z(n9732) );
  XNOR U9912 ( .A(n9726), .B(n10118), .Z(n10123) );
  XNOR U9913 ( .A(n9728), .B(n10117), .Z(n10118) );
  XNOR U9914 ( .A(n9731), .B(n10114), .Z(n10117) );
  XNOR U9915 ( .A(n9737), .B(n10113), .Z(n10114) );
  XNOR U9916 ( .A(n10106), .B(n10110), .Z(n10113) );
  XNOR U9917 ( .A(n10105), .B(n10103), .Z(n10110) );
  XNOR U9918 ( .A(n10104), .B(n10102), .Z(n10103) );
  XNOR U9919 ( .A(n9744), .B(n10097), .Z(n10102) );
  XOR U9920 ( .A(n9743), .B(n10095), .Z(n10097) );
  XNOR U9921 ( .A(n10096), .B(n10091), .Z(n10095) );
  XNOR U9922 ( .A(n10092), .B(n9759), .Z(n10091) );
  XNOR U9923 ( .A(n9754), .B(n10090), .Z(n9759) );
  XNOR U9924 ( .A(n9753), .B(n10085), .Z(n10090) );
  XNOR U9925 ( .A(n9755), .B(n10084), .Z(n10085) );
  XNOR U9926 ( .A(n9758), .B(n10081), .Z(n10084) );
  XNOR U9927 ( .A(n9764), .B(n10080), .Z(n10081) );
  XNOR U9928 ( .A(n10073), .B(n10077), .Z(n10080) );
  XNOR U9929 ( .A(n10072), .B(n10070), .Z(n10077) );
  XNOR U9930 ( .A(n10071), .B(n10069), .Z(n10070) );
  XNOR U9931 ( .A(n9771), .B(n10064), .Z(n10069) );
  XOR U9932 ( .A(n9770), .B(n10062), .Z(n10064) );
  XNOR U9933 ( .A(n10063), .B(n10058), .Z(n10062) );
  XNOR U9934 ( .A(n10059), .B(n9786), .Z(n10058) );
  XNOR U9935 ( .A(n9781), .B(n10057), .Z(n9786) );
  XNOR U9936 ( .A(n9780), .B(n10052), .Z(n10057) );
  XNOR U9937 ( .A(n9782), .B(n10051), .Z(n10052) );
  XNOR U9938 ( .A(n9785), .B(n10048), .Z(n10051) );
  XNOR U9939 ( .A(n9791), .B(n10047), .Z(n10048) );
  XNOR U9940 ( .A(n10040), .B(n10044), .Z(n10047) );
  XNOR U9941 ( .A(n10039), .B(n10037), .Z(n10044) );
  XNOR U9942 ( .A(n10038), .B(n10036), .Z(n10037) );
  XNOR U9943 ( .A(n9798), .B(n10031), .Z(n10036) );
  XOR U9944 ( .A(n9797), .B(n10029), .Z(n10031) );
  XNOR U9945 ( .A(n10030), .B(n10025), .Z(n10029) );
  XNOR U9946 ( .A(n10026), .B(n9813), .Z(n10025) );
  XNOR U9947 ( .A(n9808), .B(n10024), .Z(n9813) );
  XNOR U9948 ( .A(n9807), .B(n10019), .Z(n10024) );
  XNOR U9949 ( .A(n9809), .B(n10018), .Z(n10019) );
  XNOR U9950 ( .A(n9812), .B(n10015), .Z(n10018) );
  XNOR U9951 ( .A(n9818), .B(n10014), .Z(n10015) );
  XNOR U9952 ( .A(n10007), .B(n10011), .Z(n10014) );
  XNOR U9953 ( .A(n10006), .B(n10004), .Z(n10011) );
  XNOR U9954 ( .A(n10005), .B(n10003), .Z(n10004) );
  XNOR U9955 ( .A(n9825), .B(n9998), .Z(n10003) );
  XOR U9956 ( .A(n9824), .B(n9996), .Z(n9998) );
  XNOR U9957 ( .A(n9997), .B(n9992), .Z(n9996) );
  XNOR U9958 ( .A(n9993), .B(n9840), .Z(n9992) );
  XNOR U9959 ( .A(n9835), .B(n9991), .Z(n9840) );
  XNOR U9960 ( .A(n9834), .B(n9986), .Z(n9991) );
  XNOR U9961 ( .A(n9836), .B(n9985), .Z(n9986) );
  XNOR U9962 ( .A(n9839), .B(n9982), .Z(n9985) );
  XNOR U9963 ( .A(n9845), .B(n9981), .Z(n9982) );
  XNOR U9964 ( .A(n9974), .B(n9978), .Z(n9981) );
  XNOR U9965 ( .A(n9973), .B(n9971), .Z(n9978) );
  XNOR U9966 ( .A(n9972), .B(n9970), .Z(n9971) );
  XNOR U9967 ( .A(n9852), .B(n9965), .Z(n9970) );
  XOR U9968 ( .A(n9851), .B(n9963), .Z(n9965) );
  XNOR U9969 ( .A(n9964), .B(n9959), .Z(n9963) );
  XNOR U9970 ( .A(n9960), .B(n9867), .Z(n9959) );
  XNOR U9971 ( .A(n9862), .B(n9958), .Z(n9867) );
  XNOR U9972 ( .A(n9861), .B(n9953), .Z(n9958) );
  XNOR U9973 ( .A(n9863), .B(n9952), .Z(n9953) );
  XNOR U9974 ( .A(n9866), .B(n9949), .Z(n9952) );
  XNOR U9975 ( .A(n9872), .B(n9948), .Z(n9949) );
  XNOR U9976 ( .A(n9941), .B(n9945), .Z(n9948) );
  XNOR U9977 ( .A(n9940), .B(n9938), .Z(n9945) );
  XNOR U9978 ( .A(n9939), .B(n9937), .Z(n9938) );
  XNOR U9979 ( .A(n9879), .B(n9932), .Z(n9937) );
  XOR U9980 ( .A(n9878), .B(n9930), .Z(n9932) );
  XNOR U9981 ( .A(n9931), .B(n9926), .Z(n9930) );
  XNOR U9982 ( .A(n9927), .B(n9894), .Z(n9926) );
  XNOR U9983 ( .A(n9889), .B(n9925), .Z(n9894) );
  XNOR U9984 ( .A(n9888), .B(n9920), .Z(n9925) );
  XNOR U9985 ( .A(n9890), .B(n9919), .Z(n9920) );
  XNOR U9986 ( .A(n9893), .B(n9916), .Z(n9919) );
  XNOR U9987 ( .A(n9899), .B(n9915), .Z(n9916) );
  XNOR U9988 ( .A(n9902), .B(n9912), .Z(n9915) );
  XOR U9989 ( .A(n9901), .B(n9909), .Z(n9912) );
  XOR U9990 ( .A(n9910), .B(n9908), .Z(n9909) );
  XOR U9991 ( .A(n10904), .B(n10905), .Z(n9908) );
  XOR U9992 ( .A(n10906), .B(n10907), .Z(n10905) );
  XOR U9993 ( .A(n10908), .B(n10909), .Z(n10907) );
  NOR U9994 ( .A(n10910), .B(n10911), .Z(n10909) );
  NOR U9995 ( .A(n10912), .B(n10913), .Z(n10908) );
  NOR U9996 ( .A(n10914), .B(n10915), .Z(n10906) );
  XOR U9997 ( .A(n10916), .B(n10917), .Z(n10904) );
  XOR U9998 ( .A(n10918), .B(n10919), .Z(n10917) );
  XOR U9999 ( .A(n10920), .B(n10921), .Z(n10919) );
  XNOR U10000 ( .A(n10922), .B(n10923), .Z(n10921) );
  XOR U10001 ( .A(n10924), .B(n10925), .Z(n10923) );
  XOR U10002 ( .A(n10926), .B(n10927), .Z(n10925) );
  XOR U10003 ( .A(n10928), .B(n10929), .Z(n10927) );
  XOR U10004 ( .A(n10930), .B(n10931), .Z(n10926) );
  XOR U10005 ( .A(n10932), .B(n10933), .Z(n10931) );
  XOR U10006 ( .A(n10934), .B(n10935), .Z(n10933) );
  XOR U10007 ( .A(n10936), .B(n10937), .Z(n10935) );
  XNOR U10008 ( .A(n10938), .B(n10939), .Z(n10937) );
  XOR U10009 ( .A(n10940), .B(n10941), .Z(n10936) );
  XOR U10010 ( .A(n10942), .B(n10943), .Z(n10941) );
  AND U10011 ( .A(n10944), .B(n10945), .Z(n10942) );
  XOR U10012 ( .A(n10946), .B(n10947), .Z(n10934) );
  XOR U10013 ( .A(n10948), .B(n10949), .Z(n10947) );
  XOR U10014 ( .A(n10950), .B(n10951), .Z(n10949) );
  XOR U10015 ( .A(n10952), .B(n10953), .Z(n10951) );
  XOR U10016 ( .A(n10954), .B(n10955), .Z(n10953) );
  XOR U10017 ( .A(n10956), .B(n10957), .Z(n10955) );
  XOR U10018 ( .A(n10958), .B(n10959), .Z(n10957) );
  XOR U10019 ( .A(n10960), .B(n10961), .Z(n10959) );
  XOR U10020 ( .A(n10962), .B(n10963), .Z(n10961) );
  XOR U10021 ( .A(n10964), .B(n10965), .Z(n10963) );
  XOR U10022 ( .A(n10966), .B(n10967), .Z(n10965) );
  XOR U10023 ( .A(n10968), .B(n10969), .Z(n10967) );
  AND U10024 ( .A(n10970), .B(n10971), .Z(n10969) );
  NOR U10025 ( .A(n10972), .B(n10973), .Z(n10971) );
  NOR U10026 ( .A(n10974), .B(n10975), .Z(n10970) );
  AND U10027 ( .A(n10976), .B(n10977), .Z(n10975) );
  AND U10028 ( .A(n10978), .B(n10979), .Z(n10968) );
  NOR U10029 ( .A(n10980), .B(n10981), .Z(n10979) );
  NOR U10030 ( .A(n10982), .B(n10983), .Z(n10978) );
  AND U10031 ( .A(n10984), .B(n10985), .Z(n10983) );
  XOR U10032 ( .A(n10986), .B(n10987), .Z(n10966) );
  NOR U10033 ( .A(n10988), .B(n10989), .Z(n10987) );
  XOR U10034 ( .A(n10990), .B(n10991), .Z(n10989) );
  AND U10035 ( .A(n10992), .B(n10993), .Z(n10991) );
  NOR U10036 ( .A(n10994), .B(n10995), .Z(n10993) );
  NOR U10037 ( .A(n10996), .B(n10997), .Z(n10992) );
  AND U10038 ( .A(n10998), .B(n10999), .Z(n10997) );
  AND U10039 ( .A(n11000), .B(n11001), .Z(n10990) );
  NOR U10040 ( .A(n11002), .B(n11003), .Z(n11001) );
  AND U10041 ( .A(n10995), .B(n11004), .Z(n11003) );
  AND U10042 ( .A(n10996), .B(n11005), .Z(n11002) );
  NOR U10043 ( .A(n11006), .B(n11007), .Z(n11000) );
  XOR U10044 ( .A(n11008), .B(n11009), .Z(n11007) );
  AND U10045 ( .A(n11010), .B(n11011), .Z(n11009) );
  NOR U10046 ( .A(n11012), .B(n11013), .Z(n11011) );
  NOR U10047 ( .A(n11014), .B(n11015), .Z(n11010) );
  AND U10048 ( .A(n11016), .B(n11017), .Z(n11015) );
  AND U10049 ( .A(n11018), .B(n11019), .Z(n11008) );
  NOR U10050 ( .A(n11020), .B(n11021), .Z(n11019) );
  AND U10051 ( .A(n11013), .B(n11022), .Z(n11021) );
  AND U10052 ( .A(n11014), .B(n11023), .Z(n11020) );
  NOR U10053 ( .A(n11024), .B(n11025), .Z(n11018) );
  AND U10054 ( .A(n11026), .B(n11027), .Z(n11025) );
  AND U10055 ( .A(n11028), .B(n11029), .Z(n11027) );
  AND U10056 ( .A(n11030), .B(n11031), .Z(n11029) );
  NOR U10057 ( .A(n11032), .B(n11033), .Z(n11030) );
  NOR U10058 ( .A(n11034), .B(n11035), .Z(n11028) );
  AND U10059 ( .A(n11036), .B(n11037), .Z(n11026) );
  NOR U10060 ( .A(n11038), .B(n11039), .Z(n11037) );
  NOR U10061 ( .A(n11040), .B(n11041), .Z(n11036) );
  AND U10062 ( .A(n11012), .B(n11042), .Z(n11024) );
  AND U10063 ( .A(n10994), .B(n11043), .Z(n11006) );
  AND U10064 ( .A(n10980), .B(n11044), .Z(n10988) );
  NOR U10065 ( .A(n11045), .B(n11046), .Z(n10986) );
  AND U10066 ( .A(n10981), .B(n11047), .Z(n11046) );
  AND U10067 ( .A(n10982), .B(n11048), .Z(n11045) );
  XOR U10068 ( .A(n11049), .B(n11050), .Z(n10964) );
  XOR U10069 ( .A(n11051), .B(n11052), .Z(n11050) );
  NOR U10070 ( .A(n11053), .B(n11054), .Z(n11052) );
  AND U10071 ( .A(n10973), .B(n11055), .Z(n11054) );
  AND U10072 ( .A(n10974), .B(n11056), .Z(n11053) );
  NOR U10073 ( .A(n11057), .B(n11058), .Z(n11051) );
  AND U10074 ( .A(n11059), .B(n11060), .Z(n11058) );
  AND U10075 ( .A(n11061), .B(n11062), .Z(n11057) );
  XOR U10076 ( .A(n11063), .B(n11064), .Z(n11049) );
  AND U10077 ( .A(n10972), .B(n11065), .Z(n11064) );
  AND U10078 ( .A(n11066), .B(n11067), .Z(n11063) );
  AND U10079 ( .A(n11068), .B(n11069), .Z(n10962) );
  NOR U10080 ( .A(n11070), .B(n11071), .Z(n11069) );
  NOR U10081 ( .A(n11072), .B(n11073), .Z(n11068) );
  AND U10082 ( .A(n11074), .B(n11075), .Z(n11073) );
  XOR U10083 ( .A(n11076), .B(n11077), .Z(n10960) );
  AND U10084 ( .A(n11078), .B(n11079), .Z(n11077) );
  NOR U10085 ( .A(n11080), .B(n11081), .Z(n11079) );
  NOR U10086 ( .A(n11082), .B(n11083), .Z(n11078) );
  AND U10087 ( .A(n11084), .B(n11085), .Z(n11083) );
  AND U10088 ( .A(n11086), .B(n11087), .Z(n11076) );
  NOR U10089 ( .A(n11066), .B(n11059), .Z(n11087) );
  NOR U10090 ( .A(n11061), .B(n11088), .Z(n11086) );
  AND U10091 ( .A(n11089), .B(n11090), .Z(n11088) );
  XOR U10092 ( .A(n11091), .B(n11092), .Z(n10958) );
  XOR U10093 ( .A(n11093), .B(n11094), .Z(n11092) );
  NOR U10094 ( .A(n11095), .B(n11096), .Z(n11094) );
  AND U10095 ( .A(n11081), .B(n11097), .Z(n11096) );
  AND U10096 ( .A(n11082), .B(n11098), .Z(n11095) );
  NOR U10097 ( .A(n11099), .B(n11100), .Z(n11093) );
  AND U10098 ( .A(n11071), .B(n11101), .Z(n11100) );
  AND U10099 ( .A(n11072), .B(n11102), .Z(n11099) );
  XOR U10100 ( .A(n11103), .B(n11104), .Z(n11091) );
  AND U10101 ( .A(n11080), .B(n11105), .Z(n11104) );
  AND U10102 ( .A(n11070), .B(n11106), .Z(n11103) );
  NOR U10103 ( .A(n11107), .B(n11108), .Z(n10956) );
  AND U10104 ( .A(n11109), .B(n11110), .Z(n11108) );
  XOR U10105 ( .A(n11111), .B(n11112), .Z(n10954) );
  NOR U10106 ( .A(n11113), .B(n11114), .Z(n11112) );
  AND U10107 ( .A(n11115), .B(n11116), .Z(n11111) );
  NOR U10108 ( .A(n11117), .B(n11118), .Z(n11116) );
  NOR U10109 ( .A(n11119), .B(n11120), .Z(n11115) );
  AND U10110 ( .A(n11121), .B(n11122), .Z(n11120) );
  XOR U10111 ( .A(n11123), .B(n11124), .Z(n10952) );
  XOR U10112 ( .A(n11125), .B(n11126), .Z(n11124) );
  NOR U10113 ( .A(n11127), .B(n11128), .Z(n11126) );
  AND U10114 ( .A(n11118), .B(n11129), .Z(n11128) );
  AND U10115 ( .A(n11119), .B(n11130), .Z(n11127) );
  NOR U10116 ( .A(n11131), .B(n11132), .Z(n11125) );
  AND U10117 ( .A(n11114), .B(n11133), .Z(n11132) );
  AND U10118 ( .A(n11107), .B(n11134), .Z(n11131) );
  XOR U10119 ( .A(n11135), .B(n11136), .Z(n11123) );
  AND U10120 ( .A(n11117), .B(n11137), .Z(n11136) );
  AND U10121 ( .A(n11113), .B(n11138), .Z(n11135) );
  NOR U10122 ( .A(n11139), .B(n11140), .Z(n10950) );
  XOR U10123 ( .A(n11141), .B(n11142), .Z(n10948) );
  XOR U10124 ( .A(n11143), .B(n11144), .Z(n10946) );
  XOR U10125 ( .A(n11145), .B(n11146), .Z(n11144) );
  AND U10126 ( .A(n11139), .B(n11147), .Z(n11146) );
  AND U10127 ( .A(n11140), .B(n11148), .Z(n11145) );
  XOR U10128 ( .A(n11149), .B(n11150), .Z(n11143) );
  AND U10129 ( .A(n11141), .B(n11151), .Z(n11150) );
  AND U10130 ( .A(n11142), .B(n11152), .Z(n11149) );
  XOR U10131 ( .A(n11153), .B(n11154), .Z(n10932) );
  AND U10132 ( .A(n10943), .B(n11155), .Z(n11154) );
  AND U10133 ( .A(n11156), .B(n10940), .Z(n11153) );
  XOR U10134 ( .A(n11157), .B(n11158), .Z(n10930) );
  XOR U10135 ( .A(n11159), .B(n11160), .Z(n11158) );
  AND U10136 ( .A(n11161), .B(n10938), .Z(n11160) );
  NOR U10137 ( .A(n11162), .B(n11163), .Z(n11159) );
  XOR U10138 ( .A(n11164), .B(n11165), .Z(n11157) );
  AND U10139 ( .A(n11166), .B(n11167), .Z(n11165) );
  NOR U10140 ( .A(n11168), .B(n10928), .Z(n11164) );
  XOR U10141 ( .A(n11169), .B(n11170), .Z(n10924) );
  XNOR U10142 ( .A(n11163), .B(n11167), .Z(n11170) );
  XOR U10143 ( .A(n11171), .B(n11172), .Z(n11169) );
  NOR U10144 ( .A(n11173), .B(n10929), .Z(n11172) );
  NOR U10145 ( .A(n11174), .B(n11175), .Z(n11171) );
  XOR U10146 ( .A(n11176), .B(n11177), .Z(n10920) );
  XOR U10147 ( .A(n11178), .B(n11179), .Z(n10918) );
  XNOR U10148 ( .A(n11180), .B(n11175), .Z(n11179) );
  NOR U10149 ( .A(n11181), .B(n11176), .Z(n11180) );
  XOR U10150 ( .A(n11182), .B(n11183), .Z(n11178) );
  NOR U10151 ( .A(n11184), .B(n11177), .Z(n11183) );
  NOR U10152 ( .A(n11185), .B(n10922), .Z(n11182) );
  XOR U10153 ( .A(n11186), .B(n11187), .Z(n10916) );
  XNOR U10154 ( .A(n10911), .B(n11188), .Z(n11187) );
  XNOR U10155 ( .A(n11189), .B(n10915), .Z(n11188) );
  NOR U10156 ( .A(n11190), .B(n11191), .Z(n11189) );
  XNOR U10157 ( .A(n11191), .B(n10913), .Z(n11186) );
  XNOR U10158 ( .A(n11192), .B(n11193), .Z(n9910) );
  NOR U10159 ( .A(n11194), .B(n11192), .Z(n11193) );
  XOR U10160 ( .A(n11195), .B(n11196), .Z(n9901) );
  NOR U10161 ( .A(n11197), .B(n11195), .Z(n11196) );
  XOR U10162 ( .A(n11198), .B(n11199), .Z(n9902) );
  NOR U10163 ( .A(n11200), .B(n11198), .Z(n11199) );
  XOR U10164 ( .A(n11201), .B(n11202), .Z(n9899) );
  NOR U10165 ( .A(n11203), .B(n11201), .Z(n11202) );
  XOR U10166 ( .A(n11204), .B(n11205), .Z(n9893) );
  NOR U10167 ( .A(n11206), .B(n11204), .Z(n11205) );
  XOR U10168 ( .A(n11207), .B(n11208), .Z(n9890) );
  NOR U10169 ( .A(n11209), .B(n11207), .Z(n11208) );
  XOR U10170 ( .A(n11210), .B(n11211), .Z(n9888) );
  NOR U10171 ( .A(n11212), .B(n11210), .Z(n11211) );
  XOR U10172 ( .A(n11213), .B(n11214), .Z(n9889) );
  NOR U10173 ( .A(n11215), .B(n11213), .Z(n11214) );
  XOR U10174 ( .A(n11216), .B(n11217), .Z(n9927) );
  NOR U10175 ( .A(n11218), .B(n11216), .Z(n11217) );
  XNOR U10176 ( .A(n11219), .B(n11220), .Z(n9931) );
  NOR U10177 ( .A(n11221), .B(n11219), .Z(n11220) );
  XOR U10178 ( .A(n11222), .B(n11223), .Z(n9878) );
  NOR U10179 ( .A(n11224), .B(n11222), .Z(n11223) );
  XOR U10180 ( .A(n11225), .B(n11226), .Z(n9879) );
  NOR U10181 ( .A(n11227), .B(n11225), .Z(n11226) );
  XOR U10182 ( .A(n11228), .B(n11229), .Z(n9939) );
  NOR U10183 ( .A(n11230), .B(n11228), .Z(n11229) );
  XOR U10184 ( .A(n11231), .B(n11232), .Z(n9940) );
  NOR U10185 ( .A(n11233), .B(n11231), .Z(n11232) );
  XOR U10186 ( .A(n11234), .B(n11235), .Z(n9941) );
  NOR U10187 ( .A(n11236), .B(n11234), .Z(n11235) );
  XOR U10188 ( .A(n11237), .B(n11238), .Z(n9872) );
  NOR U10189 ( .A(n11239), .B(n11237), .Z(n11238) );
  XOR U10190 ( .A(n11240), .B(n11241), .Z(n9866) );
  NOR U10191 ( .A(n11242), .B(n11240), .Z(n11241) );
  XOR U10192 ( .A(n11243), .B(n11244), .Z(n9863) );
  NOR U10193 ( .A(n11245), .B(n11243), .Z(n11244) );
  XOR U10194 ( .A(n11246), .B(n11247), .Z(n9861) );
  NOR U10195 ( .A(n11248), .B(n11246), .Z(n11247) );
  XOR U10196 ( .A(n11249), .B(n11250), .Z(n9862) );
  NOR U10197 ( .A(n11251), .B(n11249), .Z(n11250) );
  XOR U10198 ( .A(n11252), .B(n11253), .Z(n9960) );
  NOR U10199 ( .A(n11254), .B(n11252), .Z(n11253) );
  XNOR U10200 ( .A(n11255), .B(n11256), .Z(n9964) );
  NOR U10201 ( .A(n11257), .B(n11255), .Z(n11256) );
  XOR U10202 ( .A(n11258), .B(n11259), .Z(n9851) );
  NOR U10203 ( .A(n11260), .B(n11258), .Z(n11259) );
  XOR U10204 ( .A(n11261), .B(n11262), .Z(n9852) );
  NOR U10205 ( .A(n11263), .B(n11261), .Z(n11262) );
  XOR U10206 ( .A(n11264), .B(n11265), .Z(n9972) );
  NOR U10207 ( .A(n11266), .B(n11264), .Z(n11265) );
  XOR U10208 ( .A(n11267), .B(n11268), .Z(n9973) );
  NOR U10209 ( .A(n11269), .B(n11267), .Z(n11268) );
  XOR U10210 ( .A(n11270), .B(n11271), .Z(n9974) );
  NOR U10211 ( .A(n11272), .B(n11270), .Z(n11271) );
  XOR U10212 ( .A(n11273), .B(n11274), .Z(n9845) );
  NOR U10213 ( .A(n11275), .B(n11273), .Z(n11274) );
  XOR U10214 ( .A(n11276), .B(n11277), .Z(n9839) );
  NOR U10215 ( .A(n11278), .B(n11276), .Z(n11277) );
  XOR U10216 ( .A(n11279), .B(n11280), .Z(n9836) );
  NOR U10217 ( .A(n11281), .B(n11279), .Z(n11280) );
  XOR U10218 ( .A(n11282), .B(n11283), .Z(n9834) );
  NOR U10219 ( .A(n11284), .B(n11282), .Z(n11283) );
  XOR U10220 ( .A(n11285), .B(n11286), .Z(n9835) );
  NOR U10221 ( .A(n11287), .B(n11285), .Z(n11286) );
  XOR U10222 ( .A(n11288), .B(n11289), .Z(n9993) );
  NOR U10223 ( .A(n11290), .B(n11288), .Z(n11289) );
  XNOR U10224 ( .A(n11291), .B(n11292), .Z(n9997) );
  NOR U10225 ( .A(n11293), .B(n11291), .Z(n11292) );
  XOR U10226 ( .A(n11294), .B(n11295), .Z(n9824) );
  NOR U10227 ( .A(n11296), .B(n11294), .Z(n11295) );
  XOR U10228 ( .A(n11297), .B(n11298), .Z(n9825) );
  NOR U10229 ( .A(n11299), .B(n11297), .Z(n11298) );
  XOR U10230 ( .A(n11300), .B(n11301), .Z(n10005) );
  NOR U10231 ( .A(n11302), .B(n11300), .Z(n11301) );
  XOR U10232 ( .A(n11303), .B(n11304), .Z(n10006) );
  NOR U10233 ( .A(n11305), .B(n11303), .Z(n11304) );
  XOR U10234 ( .A(n11306), .B(n11307), .Z(n10007) );
  NOR U10235 ( .A(n11308), .B(n11306), .Z(n11307) );
  XOR U10236 ( .A(n11309), .B(n11310), .Z(n9818) );
  NOR U10237 ( .A(n11311), .B(n11309), .Z(n11310) );
  XOR U10238 ( .A(n11312), .B(n11313), .Z(n9812) );
  NOR U10239 ( .A(n11314), .B(n11312), .Z(n11313) );
  XOR U10240 ( .A(n11315), .B(n11316), .Z(n9809) );
  NOR U10241 ( .A(n11317), .B(n11315), .Z(n11316) );
  XOR U10242 ( .A(n11318), .B(n11319), .Z(n9807) );
  NOR U10243 ( .A(n11320), .B(n11318), .Z(n11319) );
  XOR U10244 ( .A(n11321), .B(n11322), .Z(n9808) );
  NOR U10245 ( .A(n11323), .B(n11321), .Z(n11322) );
  XOR U10246 ( .A(n11324), .B(n11325), .Z(n10026) );
  NOR U10247 ( .A(n11326), .B(n11324), .Z(n11325) );
  XNOR U10248 ( .A(n11327), .B(n11328), .Z(n10030) );
  NOR U10249 ( .A(n11329), .B(n11327), .Z(n11328) );
  XOR U10250 ( .A(n11330), .B(n11331), .Z(n9797) );
  NOR U10251 ( .A(n11332), .B(n11330), .Z(n11331) );
  XOR U10252 ( .A(n11333), .B(n11334), .Z(n9798) );
  NOR U10253 ( .A(n11335), .B(n11333), .Z(n11334) );
  XOR U10254 ( .A(n11336), .B(n11337), .Z(n10038) );
  NOR U10255 ( .A(n11338), .B(n11336), .Z(n11337) );
  XOR U10256 ( .A(n11339), .B(n11340), .Z(n10039) );
  NOR U10257 ( .A(n11341), .B(n11339), .Z(n11340) );
  XOR U10258 ( .A(n11342), .B(n11343), .Z(n10040) );
  NOR U10259 ( .A(n11344), .B(n11342), .Z(n11343) );
  XOR U10260 ( .A(n11345), .B(n11346), .Z(n9791) );
  NOR U10261 ( .A(n11347), .B(n11345), .Z(n11346) );
  XOR U10262 ( .A(n11348), .B(n11349), .Z(n9785) );
  NOR U10263 ( .A(n11350), .B(n11348), .Z(n11349) );
  XOR U10264 ( .A(n11351), .B(n11352), .Z(n9782) );
  NOR U10265 ( .A(n11353), .B(n11351), .Z(n11352) );
  XOR U10266 ( .A(n11354), .B(n11355), .Z(n9780) );
  NOR U10267 ( .A(n11356), .B(n11354), .Z(n11355) );
  XOR U10268 ( .A(n11357), .B(n11358), .Z(n9781) );
  NOR U10269 ( .A(n11359), .B(n11357), .Z(n11358) );
  XOR U10270 ( .A(n11360), .B(n11361), .Z(n10059) );
  NOR U10271 ( .A(n11362), .B(n11360), .Z(n11361) );
  XNOR U10272 ( .A(n11363), .B(n11364), .Z(n10063) );
  NOR U10273 ( .A(n11365), .B(n11363), .Z(n11364) );
  XOR U10274 ( .A(n11366), .B(n11367), .Z(n9770) );
  NOR U10275 ( .A(n11368), .B(n11366), .Z(n11367) );
  XOR U10276 ( .A(n11369), .B(n11370), .Z(n9771) );
  NOR U10277 ( .A(n11371), .B(n11369), .Z(n11370) );
  XOR U10278 ( .A(n11372), .B(n11373), .Z(n10071) );
  NOR U10279 ( .A(n11374), .B(n11372), .Z(n11373) );
  XOR U10280 ( .A(n11375), .B(n11376), .Z(n10072) );
  NOR U10281 ( .A(n11377), .B(n11375), .Z(n11376) );
  XOR U10282 ( .A(n11378), .B(n11379), .Z(n10073) );
  NOR U10283 ( .A(n11380), .B(n11378), .Z(n11379) );
  XOR U10284 ( .A(n11381), .B(n11382), .Z(n9764) );
  NOR U10285 ( .A(n11383), .B(n11381), .Z(n11382) );
  XOR U10286 ( .A(n11384), .B(n11385), .Z(n9758) );
  NOR U10287 ( .A(n11386), .B(n11384), .Z(n11385) );
  XOR U10288 ( .A(n11387), .B(n11388), .Z(n9755) );
  NOR U10289 ( .A(n11389), .B(n11387), .Z(n11388) );
  XOR U10290 ( .A(n11390), .B(n11391), .Z(n9753) );
  NOR U10291 ( .A(n11392), .B(n11390), .Z(n11391) );
  XOR U10292 ( .A(n11393), .B(n11394), .Z(n9754) );
  NOR U10293 ( .A(n11395), .B(n11393), .Z(n11394) );
  XOR U10294 ( .A(n11396), .B(n11397), .Z(n10092) );
  NOR U10295 ( .A(n11398), .B(n11396), .Z(n11397) );
  XNOR U10296 ( .A(n11399), .B(n11400), .Z(n10096) );
  NOR U10297 ( .A(n11401), .B(n11399), .Z(n11400) );
  XOR U10298 ( .A(n11402), .B(n11403), .Z(n9743) );
  NOR U10299 ( .A(n11404), .B(n11402), .Z(n11403) );
  XOR U10300 ( .A(n11405), .B(n11406), .Z(n9744) );
  NOR U10301 ( .A(n11407), .B(n11405), .Z(n11406) );
  XOR U10302 ( .A(n11408), .B(n11409), .Z(n10104) );
  NOR U10303 ( .A(n11410), .B(n11408), .Z(n11409) );
  XOR U10304 ( .A(n11411), .B(n11412), .Z(n10105) );
  NOR U10305 ( .A(n11413), .B(n11411), .Z(n11412) );
  XOR U10306 ( .A(n11414), .B(n11415), .Z(n10106) );
  NOR U10307 ( .A(n11416), .B(n11414), .Z(n11415) );
  XOR U10308 ( .A(n11417), .B(n11418), .Z(n9737) );
  NOR U10309 ( .A(n11419), .B(n11417), .Z(n11418) );
  XOR U10310 ( .A(n11420), .B(n11421), .Z(n9731) );
  NOR U10311 ( .A(n11422), .B(n11420), .Z(n11421) );
  XOR U10312 ( .A(n11423), .B(n11424), .Z(n9728) );
  NOR U10313 ( .A(n11425), .B(n11423), .Z(n11424) );
  XOR U10314 ( .A(n11426), .B(n11427), .Z(n9726) );
  NOR U10315 ( .A(n11428), .B(n11426), .Z(n11427) );
  XOR U10316 ( .A(n11429), .B(n11430), .Z(n9727) );
  NOR U10317 ( .A(n11431), .B(n11429), .Z(n11430) );
  XOR U10318 ( .A(n11432), .B(n11433), .Z(n10125) );
  NOR U10319 ( .A(n11434), .B(n11432), .Z(n11433) );
  XNOR U10320 ( .A(n11435), .B(n11436), .Z(n10129) );
  NOR U10321 ( .A(n11437), .B(n11435), .Z(n11436) );
  XOR U10322 ( .A(n11438), .B(n11439), .Z(n9716) );
  NOR U10323 ( .A(n11440), .B(n11438), .Z(n11439) );
  XOR U10324 ( .A(n11441), .B(n11442), .Z(n9717) );
  NOR U10325 ( .A(n11443), .B(n11441), .Z(n11442) );
  XOR U10326 ( .A(n11444), .B(n11445), .Z(n10137) );
  NOR U10327 ( .A(n11446), .B(n11444), .Z(n11445) );
  XOR U10328 ( .A(n11447), .B(n11448), .Z(n10138) );
  NOR U10329 ( .A(n11449), .B(n11447), .Z(n11448) );
  XOR U10330 ( .A(n11450), .B(n11451), .Z(n10139) );
  NOR U10331 ( .A(n11452), .B(n11450), .Z(n11451) );
  XOR U10332 ( .A(n11453), .B(n11454), .Z(n9710) );
  NOR U10333 ( .A(n11455), .B(n11453), .Z(n11454) );
  XOR U10334 ( .A(n11456), .B(n11457), .Z(n9704) );
  NOR U10335 ( .A(n11458), .B(n11456), .Z(n11457) );
  XOR U10336 ( .A(n11459), .B(n11460), .Z(n9701) );
  NOR U10337 ( .A(n11461), .B(n11459), .Z(n11460) );
  XOR U10338 ( .A(n11462), .B(n11463), .Z(n9699) );
  NOR U10339 ( .A(n11464), .B(n11462), .Z(n11463) );
  XOR U10340 ( .A(n11465), .B(n11466), .Z(n9700) );
  NOR U10341 ( .A(n11467), .B(n11465), .Z(n11466) );
  XOR U10342 ( .A(n11468), .B(n11469), .Z(n10158) );
  NOR U10343 ( .A(n11470), .B(n11468), .Z(n11469) );
  XNOR U10344 ( .A(n11471), .B(n11472), .Z(n10162) );
  NOR U10345 ( .A(n11473), .B(n11471), .Z(n11472) );
  XOR U10346 ( .A(n11474), .B(n11475), .Z(n9689) );
  NOR U10347 ( .A(n11476), .B(n11474), .Z(n11475) );
  XOR U10348 ( .A(n11477), .B(n11478), .Z(n9690) );
  NOR U10349 ( .A(n11479), .B(n11477), .Z(n11478) );
  XOR U10350 ( .A(n11480), .B(n11481), .Z(n10170) );
  NOR U10351 ( .A(n11482), .B(n11480), .Z(n11481) );
  XOR U10352 ( .A(n11483), .B(n11484), .Z(n10171) );
  NOR U10353 ( .A(n11485), .B(n11483), .Z(n11484) );
  XOR U10354 ( .A(n11486), .B(n11487), .Z(n10172) );
  NOR U10355 ( .A(n11488), .B(n11486), .Z(n11487) );
  XOR U10356 ( .A(n11489), .B(n11490), .Z(n9683) );
  NOR U10357 ( .A(n11491), .B(n11489), .Z(n11490) );
  XOR U10358 ( .A(n11492), .B(n11493), .Z(n9677) );
  NOR U10359 ( .A(n11494), .B(n11492), .Z(n11493) );
  XOR U10360 ( .A(n11495), .B(n11496), .Z(n9674) );
  NOR U10361 ( .A(n11497), .B(n11495), .Z(n11496) );
  XOR U10362 ( .A(n11498), .B(n11499), .Z(n9672) );
  NOR U10363 ( .A(n11500), .B(n11498), .Z(n11499) );
  XOR U10364 ( .A(n11501), .B(n11502), .Z(n9673) );
  NOR U10365 ( .A(n11503), .B(n11501), .Z(n11502) );
  XOR U10366 ( .A(n11504), .B(n11505), .Z(n10191) );
  NOR U10367 ( .A(n11506), .B(n11504), .Z(n11505) );
  XNOR U10368 ( .A(n11507), .B(n11508), .Z(n10195) );
  NOR U10369 ( .A(n11509), .B(n11507), .Z(n11508) );
  XOR U10370 ( .A(n11510), .B(n11511), .Z(n9662) );
  NOR U10371 ( .A(n11512), .B(n11510), .Z(n11511) );
  XOR U10372 ( .A(n11513), .B(n11514), .Z(n9663) );
  NOR U10373 ( .A(n11515), .B(n11513), .Z(n11514) );
  XOR U10374 ( .A(n11516), .B(n11517), .Z(n10203) );
  NOR U10375 ( .A(n11518), .B(n11516), .Z(n11517) );
  XOR U10376 ( .A(n11519), .B(n11520), .Z(n10204) );
  NOR U10377 ( .A(n11521), .B(n11519), .Z(n11520) );
  XOR U10378 ( .A(n11522), .B(n11523), .Z(n10205) );
  NOR U10379 ( .A(n11524), .B(n11522), .Z(n11523) );
  XOR U10380 ( .A(n11525), .B(n11526), .Z(n9656) );
  NOR U10381 ( .A(n11527), .B(n11525), .Z(n11526) );
  XOR U10382 ( .A(n11528), .B(n11529), .Z(n9650) );
  NOR U10383 ( .A(n11530), .B(n11528), .Z(n11529) );
  XOR U10384 ( .A(n11531), .B(n11532), .Z(n9647) );
  NOR U10385 ( .A(n11533), .B(n11531), .Z(n11532) );
  XOR U10386 ( .A(n11534), .B(n11535), .Z(n9645) );
  NOR U10387 ( .A(n11536), .B(n11534), .Z(n11535) );
  XOR U10388 ( .A(n11537), .B(n11538), .Z(n9646) );
  NOR U10389 ( .A(n11539), .B(n11537), .Z(n11538) );
  XOR U10390 ( .A(n11540), .B(n11541), .Z(n10224) );
  NOR U10391 ( .A(n11542), .B(n11540), .Z(n11541) );
  XNOR U10392 ( .A(n11543), .B(n11544), .Z(n10228) );
  NOR U10393 ( .A(n11545), .B(n11543), .Z(n11544) );
  XOR U10394 ( .A(n11546), .B(n11547), .Z(n9635) );
  NOR U10395 ( .A(n11548), .B(n11546), .Z(n11547) );
  XOR U10396 ( .A(n11549), .B(n11550), .Z(n9636) );
  NOR U10397 ( .A(n11551), .B(n11549), .Z(n11550) );
  XOR U10398 ( .A(n11552), .B(n11553), .Z(n10236) );
  NOR U10399 ( .A(n11554), .B(n11552), .Z(n11553) );
  XOR U10400 ( .A(n11555), .B(n11556), .Z(n10237) );
  NOR U10401 ( .A(n11557), .B(n11555), .Z(n11556) );
  XOR U10402 ( .A(n11558), .B(n11559), .Z(n10238) );
  NOR U10403 ( .A(n11560), .B(n11558), .Z(n11559) );
  XOR U10404 ( .A(n11561), .B(n11562), .Z(n9629) );
  NOR U10405 ( .A(n11563), .B(n11561), .Z(n11562) );
  XOR U10406 ( .A(n11564), .B(n11565), .Z(n9622) );
  NOR U10407 ( .A(n11566), .B(n11564), .Z(n11565) );
  XOR U10408 ( .A(n11567), .B(n11568), .Z(n9618) );
  NOR U10409 ( .A(n11569), .B(n11567), .Z(n11568) );
  XOR U10410 ( .A(n11570), .B(n11571), .Z(n9620) );
  NOR U10411 ( .A(n11572), .B(n11570), .Z(n11571) );
  IV U10412 ( .A(n10252), .Z(n10903) );
  XOR U10413 ( .A(n11573), .B(n11574), .Z(n10252) );
  AND U10414 ( .A(n11575), .B(n11573), .Z(n11574) );
  XNOR U10415 ( .A(n11576), .B(n11577), .Z(n10253) );
  AND U10416 ( .A(n63), .B(n11576), .Z(n11577) );
  XNOR U10417 ( .A(n10899), .B(n47), .Z(n10901) );
  XOR U10418 ( .A(n11578), .B(n10278), .Z(n47) );
  XOR U10419 ( .A(n10277), .B(n10266), .Z(n10278) );
  XOR U10420 ( .A(n11579), .B(n10264), .Z(n10266) );
  XNOR U10421 ( .A(n10265), .B(n10261), .Z(n10264) );
  XNOR U10422 ( .A(n10260), .B(n10287), .Z(n10261) );
  XNOR U10423 ( .A(n10286), .B(n10896), .Z(n10287) );
  XNOR U10424 ( .A(n10887), .B(n10895), .Z(n10896) );
  XNOR U10425 ( .A(n10886), .B(n10892), .Z(n10895) );
  XNOR U10426 ( .A(n10891), .B(n10296), .Z(n10892) );
  XNOR U10427 ( .A(n10295), .B(n10885), .Z(n10296) );
  XNOR U10428 ( .A(n10876), .B(n10884), .Z(n10885) );
  XNOR U10429 ( .A(n10875), .B(n10881), .Z(n10884) );
  XNOR U10430 ( .A(n10880), .B(n10305), .Z(n10881) );
  XNOR U10431 ( .A(n10304), .B(n10874), .Z(n10305) );
  XNOR U10432 ( .A(n10865), .B(n10873), .Z(n10874) );
  XNOR U10433 ( .A(n10864), .B(n10870), .Z(n10873) );
  XNOR U10434 ( .A(n10869), .B(n10314), .Z(n10870) );
  XNOR U10435 ( .A(n10313), .B(n10863), .Z(n10314) );
  XNOR U10436 ( .A(n10854), .B(n10862), .Z(n10863) );
  XNOR U10437 ( .A(n10853), .B(n10859), .Z(n10862) );
  XNOR U10438 ( .A(n10858), .B(n10323), .Z(n10859) );
  XNOR U10439 ( .A(n10322), .B(n10852), .Z(n10323) );
  XNOR U10440 ( .A(n10843), .B(n10851), .Z(n10852) );
  XNOR U10441 ( .A(n10842), .B(n10848), .Z(n10851) );
  XNOR U10442 ( .A(n10847), .B(n10332), .Z(n10848) );
  XNOR U10443 ( .A(n10331), .B(n10841), .Z(n10332) );
  XNOR U10444 ( .A(n10832), .B(n10840), .Z(n10841) );
  XNOR U10445 ( .A(n10831), .B(n10837), .Z(n10840) );
  XNOR U10446 ( .A(n10836), .B(n10341), .Z(n10837) );
  XNOR U10447 ( .A(n10340), .B(n10830), .Z(n10341) );
  XNOR U10448 ( .A(n10821), .B(n10829), .Z(n10830) );
  XNOR U10449 ( .A(n10820), .B(n10826), .Z(n10829) );
  XNOR U10450 ( .A(n10825), .B(n10350), .Z(n10826) );
  XNOR U10451 ( .A(n10349), .B(n10819), .Z(n10350) );
  XNOR U10452 ( .A(n10810), .B(n10818), .Z(n10819) );
  XNOR U10453 ( .A(n10809), .B(n10815), .Z(n10818) );
  XNOR U10454 ( .A(n10814), .B(n10359), .Z(n10815) );
  XNOR U10455 ( .A(n10358), .B(n10808), .Z(n10359) );
  XNOR U10456 ( .A(n10799), .B(n10807), .Z(n10808) );
  XNOR U10457 ( .A(n10798), .B(n10804), .Z(n10807) );
  XNOR U10458 ( .A(n10803), .B(n10368), .Z(n10804) );
  XNOR U10459 ( .A(n10367), .B(n10797), .Z(n10368) );
  XNOR U10460 ( .A(n10788), .B(n10796), .Z(n10797) );
  XNOR U10461 ( .A(n10787), .B(n10793), .Z(n10796) );
  XNOR U10462 ( .A(n10792), .B(n10377), .Z(n10793) );
  XNOR U10463 ( .A(n10376), .B(n10786), .Z(n10377) );
  XNOR U10464 ( .A(n10777), .B(n10785), .Z(n10786) );
  XNOR U10465 ( .A(n10776), .B(n10782), .Z(n10785) );
  XNOR U10466 ( .A(n10781), .B(n10386), .Z(n10782) );
  XNOR U10467 ( .A(n10385), .B(n10775), .Z(n10386) );
  XNOR U10468 ( .A(n10766), .B(n10774), .Z(n10775) );
  XNOR U10469 ( .A(n10765), .B(n10771), .Z(n10774) );
  XNOR U10470 ( .A(n10770), .B(n10395), .Z(n10771) );
  XNOR U10471 ( .A(n10394), .B(n10764), .Z(n10395) );
  XNOR U10472 ( .A(n10755), .B(n10763), .Z(n10764) );
  XNOR U10473 ( .A(n10754), .B(n10760), .Z(n10763) );
  XNOR U10474 ( .A(n10759), .B(n10404), .Z(n10760) );
  XNOR U10475 ( .A(n10403), .B(n10753), .Z(n10404) );
  XNOR U10476 ( .A(n10744), .B(n10752), .Z(n10753) );
  XNOR U10477 ( .A(n10743), .B(n10749), .Z(n10752) );
  XNOR U10478 ( .A(n10748), .B(n10413), .Z(n10749) );
  XNOR U10479 ( .A(n10412), .B(n10742), .Z(n10413) );
  XNOR U10480 ( .A(n10733), .B(n10741), .Z(n10742) );
  XNOR U10481 ( .A(n10732), .B(n10738), .Z(n10741) );
  XNOR U10482 ( .A(n10737), .B(n10422), .Z(n10738) );
  XNOR U10483 ( .A(n10421), .B(n10731), .Z(n10422) );
  XNOR U10484 ( .A(n10722), .B(n10730), .Z(n10731) );
  XNOR U10485 ( .A(n10721), .B(n10727), .Z(n10730) );
  XNOR U10486 ( .A(n10726), .B(n10431), .Z(n10727) );
  XNOR U10487 ( .A(n10430), .B(n10720), .Z(n10431) );
  XNOR U10488 ( .A(n10711), .B(n10719), .Z(n10720) );
  XNOR U10489 ( .A(n10710), .B(n10716), .Z(n10719) );
  XNOR U10490 ( .A(n10715), .B(n10440), .Z(n10716) );
  XNOR U10491 ( .A(n10439), .B(n10709), .Z(n10440) );
  XNOR U10492 ( .A(n10700), .B(n10708), .Z(n10709) );
  XNOR U10493 ( .A(n10699), .B(n10705), .Z(n10708) );
  XNOR U10494 ( .A(n10704), .B(n10449), .Z(n10705) );
  XNOR U10495 ( .A(n10448), .B(n10698), .Z(n10449) );
  XNOR U10496 ( .A(n10689), .B(n10697), .Z(n10698) );
  XNOR U10497 ( .A(n10688), .B(n10694), .Z(n10697) );
  XNOR U10498 ( .A(n10693), .B(n10458), .Z(n10694) );
  XNOR U10499 ( .A(n10457), .B(n10687), .Z(n10458) );
  XNOR U10500 ( .A(n10678), .B(n10686), .Z(n10687) );
  XNOR U10501 ( .A(n10677), .B(n10683), .Z(n10686) );
  XNOR U10502 ( .A(n10682), .B(n10467), .Z(n10683) );
  XNOR U10503 ( .A(n10466), .B(n10676), .Z(n10467) );
  XNOR U10504 ( .A(n10667), .B(n10675), .Z(n10676) );
  XNOR U10505 ( .A(n10666), .B(n10672), .Z(n10675) );
  XNOR U10506 ( .A(n10671), .B(n10476), .Z(n10672) );
  XNOR U10507 ( .A(n10475), .B(n10665), .Z(n10476) );
  XNOR U10508 ( .A(n10656), .B(n10664), .Z(n10665) );
  XNOR U10509 ( .A(n10655), .B(n10661), .Z(n10664) );
  XNOR U10510 ( .A(n10660), .B(n10485), .Z(n10661) );
  XNOR U10511 ( .A(n10484), .B(n10654), .Z(n10485) );
  XNOR U10512 ( .A(n10645), .B(n10653), .Z(n10654) );
  XNOR U10513 ( .A(n10644), .B(n10650), .Z(n10653) );
  XNOR U10514 ( .A(n10649), .B(n10494), .Z(n10650) );
  XNOR U10515 ( .A(n10493), .B(n10643), .Z(n10494) );
  XNOR U10516 ( .A(n10634), .B(n10642), .Z(n10643) );
  XNOR U10517 ( .A(n10633), .B(n10639), .Z(n10642) );
  XNOR U10518 ( .A(n10638), .B(n10503), .Z(n10639) );
  XNOR U10519 ( .A(n10502), .B(n10632), .Z(n10503) );
  XNOR U10520 ( .A(n10623), .B(n10631), .Z(n10632) );
  XNOR U10521 ( .A(n10622), .B(n10628), .Z(n10631) );
  XNOR U10522 ( .A(n10627), .B(n10512), .Z(n10628) );
  XNOR U10523 ( .A(n10511), .B(n10621), .Z(n10512) );
  XNOR U10524 ( .A(n10612), .B(n10620), .Z(n10621) );
  XNOR U10525 ( .A(n10611), .B(n10617), .Z(n10620) );
  XNOR U10526 ( .A(n10616), .B(n10521), .Z(n10617) );
  XNOR U10527 ( .A(n10520), .B(n10610), .Z(n10521) );
  XNOR U10528 ( .A(n10601), .B(n10609), .Z(n10610) );
  XNOR U10529 ( .A(n10600), .B(n10606), .Z(n10609) );
  XNOR U10530 ( .A(n10605), .B(n10530), .Z(n10606) );
  XNOR U10531 ( .A(n10529), .B(n10599), .Z(n10530) );
  XNOR U10532 ( .A(n10590), .B(n10598), .Z(n10599) );
  XNOR U10533 ( .A(n10589), .B(n10595), .Z(n10598) );
  XNOR U10534 ( .A(n10594), .B(n10577), .Z(n10595) );
  XNOR U10535 ( .A(n10536), .B(n10588), .Z(n10577) );
  XNOR U10536 ( .A(n10579), .B(n10587), .Z(n10588) );
  XNOR U10537 ( .A(n10578), .B(n10584), .Z(n10587) );
  XNOR U10538 ( .A(n10583), .B(n10567), .Z(n10584) );
  XNOR U10539 ( .A(n10539), .B(n10576), .Z(n10567) );
  XNOR U10540 ( .A(n10563), .B(n10573), .Z(n10576) );
  XNOR U10541 ( .A(n10566), .B(n10572), .Z(n10573) );
  XNOR U10542 ( .A(n10535), .B(n10562), .Z(n10572) );
  XNOR U10543 ( .A(n10545), .B(n10561), .Z(n10562) );
  XNOR U10544 ( .A(n10548), .B(n10558), .Z(n10561) );
  XOR U10545 ( .A(n10547), .B(n10555), .Z(n10558) );
  XOR U10546 ( .A(n10556), .B(n10554), .Z(n10555) );
  XOR U10547 ( .A(n11580), .B(n11581), .Z(n10554) );
  XOR U10548 ( .A(n11582), .B(n11583), .Z(n11581) );
  XNOR U10549 ( .A(n11584), .B(n11585), .Z(n11583) );
  NOR U10550 ( .A(n11586), .B(n11585), .Z(n11584) );
  XOR U10551 ( .A(n11587), .B(n11588), .Z(n11582) );
  NOR U10552 ( .A(n11589), .B(n11590), .Z(n11588) );
  NOR U10553 ( .A(n11591), .B(n11592), .Z(n11587) );
  XOR U10554 ( .A(n11593), .B(n11594), .Z(n11580) );
  XOR U10555 ( .A(n11595), .B(n11596), .Z(n11594) );
  XOR U10556 ( .A(n11597), .B(n11598), .Z(n11596) );
  XOR U10557 ( .A(n11599), .B(n11600), .Z(n11598) );
  XOR U10558 ( .A(n11601), .B(n11602), .Z(n11600) );
  AND U10559 ( .A(n11603), .B(n11602), .Z(n11601) );
  XOR U10560 ( .A(n11604), .B(n11605), .Z(n11599) );
  XOR U10561 ( .A(n11606), .B(n11607), .Z(n11605) );
  XOR U10562 ( .A(n11608), .B(n11609), .Z(n11607) );
  XNOR U10563 ( .A(n11610), .B(n11611), .Z(n11609) );
  NOR U10564 ( .A(n11612), .B(n11611), .Z(n11610) );
  XOR U10565 ( .A(n11613), .B(n11614), .Z(n11608) );
  XOR U10566 ( .A(n11615), .B(n11616), .Z(n11614) );
  XOR U10567 ( .A(n11617), .B(n11618), .Z(n11616) );
  XNOR U10568 ( .A(n11619), .B(n11620), .Z(n11618) );
  NOR U10569 ( .A(n11621), .B(n11620), .Z(n11619) );
  XOR U10570 ( .A(n11622), .B(n11623), .Z(n11617) );
  XOR U10571 ( .A(n11624), .B(n11625), .Z(n11623) );
  XOR U10572 ( .A(n11626), .B(n11627), .Z(n11625) );
  NOR U10573 ( .A(n11628), .B(n11629), .Z(n11626) );
  XOR U10574 ( .A(n11630), .B(n11631), .Z(n11624) );
  XOR U10575 ( .A(n11632), .B(n11633), .Z(n11631) );
  XOR U10576 ( .A(n11634), .B(n11635), .Z(n11633) );
  XOR U10577 ( .A(n11636), .B(n11637), .Z(n11635) );
  AND U10578 ( .A(n11637), .B(n11638), .Z(n11636) );
  XOR U10579 ( .A(n11639), .B(n11640), .Z(n11634) );
  XOR U10580 ( .A(n11641), .B(n11642), .Z(n11640) );
  XOR U10581 ( .A(n11643), .B(n11644), .Z(n11642) );
  XOR U10582 ( .A(n11645), .B(n11646), .Z(n11644) );
  XOR U10583 ( .A(n11647), .B(n11648), .Z(n11646) );
  XOR U10584 ( .A(n11649), .B(n11650), .Z(n11648) );
  XOR U10585 ( .A(n11651), .B(n11652), .Z(n11650) );
  XOR U10586 ( .A(n11653), .B(n11654), .Z(n11652) );
  XOR U10587 ( .A(n11655), .B(n11656), .Z(n11654) );
  AND U10588 ( .A(n11657), .B(n11658), .Z(n11656) );
  AND U10589 ( .A(n11659), .B(n11660), .Z(n11655) );
  XOR U10590 ( .A(n11661), .B(n11662), .Z(n11653) );
  AND U10591 ( .A(n11663), .B(n11664), .Z(n11662) );
  AND U10592 ( .A(n11665), .B(n11666), .Z(n11661) );
  AND U10593 ( .A(n11667), .B(n11668), .Z(n11666) );
  NOR U10594 ( .A(n11669), .B(n11670), .Z(n11668) );
  IV U10595 ( .A(n11671), .Z(n11669) );
  NOR U10596 ( .A(n11672), .B(n11673), .Z(n11671) );
  NOR U10597 ( .A(n11674), .B(n11675), .Z(n11667) );
  AND U10598 ( .A(n11676), .B(n11677), .Z(n11665) );
  NOR U10599 ( .A(n11678), .B(n11679), .Z(n11677) );
  NOR U10600 ( .A(n11680), .B(n11681), .Z(n11676) );
  XOR U10601 ( .A(n11682), .B(n11683), .Z(n11651) );
  XOR U10602 ( .A(n11684), .B(n11685), .Z(n11683) );
  NOR U10603 ( .A(n11686), .B(n11687), .Z(n11685) );
  NOR U10604 ( .A(n11688), .B(n11689), .Z(n11684) );
  AND U10605 ( .A(n11690), .B(n11691), .Z(n11689) );
  IV U10606 ( .A(n11692), .Z(n11688) );
  NOR U10607 ( .A(n11693), .B(n11694), .Z(n11692) );
  AND U10608 ( .A(n11686), .B(n11695), .Z(n11694) );
  AND U10609 ( .A(n11687), .B(n11696), .Z(n11693) );
  XOR U10610 ( .A(n11697), .B(n11698), .Z(n11682) );
  NOR U10611 ( .A(n11699), .B(n11700), .Z(n11698) );
  NOR U10612 ( .A(n11701), .B(n11702), .Z(n11697) );
  AND U10613 ( .A(n11703), .B(n11704), .Z(n11702) );
  IV U10614 ( .A(n11705), .Z(n11701) );
  NOR U10615 ( .A(n11706), .B(n11707), .Z(n11705) );
  AND U10616 ( .A(n11699), .B(n11708), .Z(n11707) );
  AND U10617 ( .A(n11700), .B(n11709), .Z(n11706) );
  AND U10618 ( .A(n11710), .B(n11711), .Z(n11649) );
  XOR U10619 ( .A(n11712), .B(n11713), .Z(n11647) );
  AND U10620 ( .A(n11714), .B(n11715), .Z(n11713) );
  NOR U10621 ( .A(n11716), .B(n11717), .Z(n11712) );
  XOR U10622 ( .A(n11718), .B(n11719), .Z(n11645) );
  XOR U10623 ( .A(n11720), .B(n11721), .Z(n11719) );
  NOR U10624 ( .A(n11722), .B(n11723), .Z(n11721) );
  AND U10625 ( .A(n11724), .B(n11725), .Z(n11723) );
  IV U10626 ( .A(n11726), .Z(n11722) );
  NOR U10627 ( .A(n11727), .B(n11728), .Z(n11726) );
  AND U10628 ( .A(n11716), .B(n11729), .Z(n11728) );
  AND U10629 ( .A(n11717), .B(n11730), .Z(n11727) );
  NOR U10630 ( .A(n11731), .B(n11732), .Z(n11720) );
  XOR U10631 ( .A(n11733), .B(n11734), .Z(n11718) );
  NOR U10632 ( .A(n11735), .B(n11736), .Z(n11734) );
  AND U10633 ( .A(n11737), .B(n11738), .Z(n11736) );
  IV U10634 ( .A(n11739), .Z(n11735) );
  NOR U10635 ( .A(n11740), .B(n11741), .Z(n11739) );
  AND U10636 ( .A(n11731), .B(n11742), .Z(n11741) );
  AND U10637 ( .A(n11732), .B(n11743), .Z(n11740) );
  NOR U10638 ( .A(n11744), .B(n11745), .Z(n11733) );
  AND U10639 ( .A(n11746), .B(n11747), .Z(n11643) );
  XOR U10640 ( .A(n11748), .B(n11749), .Z(n11641) );
  AND U10641 ( .A(n11750), .B(n11751), .Z(n11749) );
  NOR U10642 ( .A(n11752), .B(n11753), .Z(n11748) );
  AND U10643 ( .A(n11754), .B(n11755), .Z(n11753) );
  IV U10644 ( .A(n11756), .Z(n11752) );
  NOR U10645 ( .A(n11757), .B(n11758), .Z(n11756) );
  AND U10646 ( .A(n11744), .B(n11759), .Z(n11758) );
  AND U10647 ( .A(n11745), .B(n11760), .Z(n11757) );
  XOR U10648 ( .A(n11761), .B(n11762), .Z(n11639) );
  XOR U10649 ( .A(n11763), .B(n11764), .Z(n11762) );
  NOR U10650 ( .A(n11765), .B(n11766), .Z(n11764) );
  NOR U10651 ( .A(n11767), .B(n11768), .Z(n11763) );
  AND U10652 ( .A(n11769), .B(n11770), .Z(n11768) );
  IV U10653 ( .A(n11771), .Z(n11767) );
  NOR U10654 ( .A(n11772), .B(n11773), .Z(n11771) );
  AND U10655 ( .A(n11765), .B(n11774), .Z(n11773) );
  AND U10656 ( .A(n11766), .B(n11775), .Z(n11772) );
  XOR U10657 ( .A(n11776), .B(n11777), .Z(n11761) );
  NOR U10658 ( .A(n11778), .B(n11779), .Z(n11777) );
  NOR U10659 ( .A(n11780), .B(n11781), .Z(n11776) );
  AND U10660 ( .A(n11782), .B(n11783), .Z(n11781) );
  IV U10661 ( .A(n11784), .Z(n11780) );
  NOR U10662 ( .A(n11785), .B(n11786), .Z(n11784) );
  AND U10663 ( .A(n11778), .B(n11787), .Z(n11786) );
  AND U10664 ( .A(n11779), .B(n11788), .Z(n11785) );
  XOR U10665 ( .A(n11789), .B(n11790), .Z(n11632) );
  AND U10666 ( .A(n11791), .B(n11792), .Z(n11790) );
  AND U10667 ( .A(n11793), .B(n11794), .Z(n11789) );
  XOR U10668 ( .A(n11795), .B(n11796), .Z(n11630) );
  XOR U10669 ( .A(n11797), .B(n11798), .Z(n11796) );
  NOR U10670 ( .A(n11799), .B(n11800), .Z(n11798) );
  NOR U10671 ( .A(n11801), .B(n11802), .Z(n11797) );
  AND U10672 ( .A(n11803), .B(n11804), .Z(n11802) );
  IV U10673 ( .A(n11805), .Z(n11801) );
  NOR U10674 ( .A(n11806), .B(n11807), .Z(n11805) );
  AND U10675 ( .A(n11799), .B(n11808), .Z(n11807) );
  AND U10676 ( .A(n11800), .B(n11809), .Z(n11806) );
  XOR U10677 ( .A(n11810), .B(n11811), .Z(n11795) );
  NOR U10678 ( .A(n11812), .B(n11813), .Z(n11811) );
  NOR U10679 ( .A(n11814), .B(n11815), .Z(n11810) );
  AND U10680 ( .A(n11816), .B(n11817), .Z(n11815) );
  IV U10681 ( .A(n11818), .Z(n11814) );
  NOR U10682 ( .A(n11819), .B(n11820), .Z(n11818) );
  AND U10683 ( .A(n11812), .B(n11821), .Z(n11820) );
  AND U10684 ( .A(n11813), .B(n11822), .Z(n11819) );
  XOR U10685 ( .A(n11823), .B(n11824), .Z(n11622) );
  XOR U10686 ( .A(n11825), .B(n11826), .Z(n11824) );
  AND U10687 ( .A(n11827), .B(n11828), .Z(n11826) );
  AND U10688 ( .A(n11628), .B(n11829), .Z(n11825) );
  XOR U10689 ( .A(n11830), .B(n11831), .Z(n11823) );
  AND U10690 ( .A(n11629), .B(n11832), .Z(n11831) );
  AND U10691 ( .A(n11833), .B(n11627), .Z(n11830) );
  XNOR U10692 ( .A(n11834), .B(n11835), .Z(n11615) );
  XOR U10693 ( .A(n11836), .B(n11837), .Z(n11613) );
  XOR U10694 ( .A(n11838), .B(n11839), .Z(n11837) );
  AND U10695 ( .A(n11839), .B(n11840), .Z(n11838) );
  XOR U10696 ( .A(n11841), .B(n11842), .Z(n11836) );
  AND U10697 ( .A(n11843), .B(n11834), .Z(n11842) );
  AND U10698 ( .A(n11844), .B(n11845), .Z(n11841) );
  XOR U10699 ( .A(n11846), .B(n11847), .Z(n11606) );
  XOR U10700 ( .A(n11848), .B(n11849), .Z(n11604) );
  XOR U10701 ( .A(n11850), .B(n11851), .Z(n11849) );
  AND U10702 ( .A(n11852), .B(n11851), .Z(n11850) );
  XOR U10703 ( .A(n11853), .B(n11854), .Z(n11848) );
  NOR U10704 ( .A(n11855), .B(n11846), .Z(n11854) );
  NOR U10705 ( .A(n11856), .B(n11847), .Z(n11853) );
  XOR U10706 ( .A(n11857), .B(n11858), .Z(n11597) );
  XOR U10707 ( .A(n11859), .B(n11860), .Z(n11595) );
  XNOR U10708 ( .A(n11861), .B(n11862), .Z(n11860) );
  NOR U10709 ( .A(n11863), .B(n11862), .Z(n11861) );
  XOR U10710 ( .A(n11864), .B(n11865), .Z(n11859) );
  NOR U10711 ( .A(n11866), .B(n11857), .Z(n11865) );
  NOR U10712 ( .A(n11867), .B(n11858), .Z(n11864) );
  XNOR U10713 ( .A(n11592), .B(n11590), .Z(n11593) );
  XNOR U10714 ( .A(n11868), .B(n11869), .Z(n10556) );
  NOR U10715 ( .A(n11870), .B(n11868), .Z(n11869) );
  XOR U10716 ( .A(n11871), .B(n11872), .Z(n10547) );
  NOR U10717 ( .A(n11873), .B(n11871), .Z(n11872) );
  XOR U10718 ( .A(n11874), .B(n11875), .Z(n10548) );
  NOR U10719 ( .A(n11876), .B(n11874), .Z(n11875) );
  XOR U10720 ( .A(n11877), .B(n11878), .Z(n10545) );
  NOR U10721 ( .A(n11879), .B(n11877), .Z(n11878) );
  XOR U10722 ( .A(n11880), .B(n11881), .Z(n10535) );
  NOR U10723 ( .A(n11882), .B(n11880), .Z(n11881) );
  XOR U10724 ( .A(n11883), .B(n11884), .Z(n10566) );
  NOR U10725 ( .A(n11885), .B(n11883), .Z(n11884) );
  XOR U10726 ( .A(n11886), .B(n11887), .Z(n10563) );
  NOR U10727 ( .A(n11888), .B(n11886), .Z(n11887) );
  XOR U10728 ( .A(n11889), .B(n11890), .Z(n10539) );
  NOR U10729 ( .A(n11891), .B(n11889), .Z(n11890) );
  XOR U10730 ( .A(n11892), .B(n11893), .Z(n10583) );
  NOR U10731 ( .A(n11894), .B(n11892), .Z(n11893) );
  XOR U10732 ( .A(n11895), .B(n11896), .Z(n10578) );
  NOR U10733 ( .A(n11897), .B(n11895), .Z(n11896) );
  XOR U10734 ( .A(n11898), .B(n11899), .Z(n10579) );
  NOR U10735 ( .A(n11900), .B(n11898), .Z(n11899) );
  XOR U10736 ( .A(n11901), .B(n11902), .Z(n10536) );
  NOR U10737 ( .A(n11903), .B(n11901), .Z(n11902) );
  XOR U10738 ( .A(n11904), .B(n11905), .Z(n10594) );
  NOR U10739 ( .A(n11906), .B(n11904), .Z(n11905) );
  XOR U10740 ( .A(n11907), .B(n11908), .Z(n10589) );
  NOR U10741 ( .A(n11909), .B(n11907), .Z(n11908) );
  XOR U10742 ( .A(n11910), .B(n11911), .Z(n10590) );
  NOR U10743 ( .A(n11912), .B(n11910), .Z(n11911) );
  XOR U10744 ( .A(n11913), .B(n11914), .Z(n10529) );
  NOR U10745 ( .A(n11915), .B(n11913), .Z(n11914) );
  XOR U10746 ( .A(n11916), .B(n11917), .Z(n10605) );
  NOR U10747 ( .A(n11918), .B(n11916), .Z(n11917) );
  XOR U10748 ( .A(n11919), .B(n11920), .Z(n10600) );
  NOR U10749 ( .A(n11921), .B(n11919), .Z(n11920) );
  XOR U10750 ( .A(n11922), .B(n11923), .Z(n10601) );
  NOR U10751 ( .A(n11924), .B(n11922), .Z(n11923) );
  XOR U10752 ( .A(n11925), .B(n11926), .Z(n10520) );
  NOR U10753 ( .A(n11927), .B(n11925), .Z(n11926) );
  XOR U10754 ( .A(n11928), .B(n11929), .Z(n10616) );
  NOR U10755 ( .A(n11930), .B(n11928), .Z(n11929) );
  XOR U10756 ( .A(n11931), .B(n11932), .Z(n10611) );
  NOR U10757 ( .A(n11933), .B(n11931), .Z(n11932) );
  XOR U10758 ( .A(n11934), .B(n11935), .Z(n10612) );
  NOR U10759 ( .A(n11936), .B(n11934), .Z(n11935) );
  XOR U10760 ( .A(n11937), .B(n11938), .Z(n10511) );
  NOR U10761 ( .A(n11939), .B(n11937), .Z(n11938) );
  XOR U10762 ( .A(n11940), .B(n11941), .Z(n10627) );
  NOR U10763 ( .A(n11942), .B(n11940), .Z(n11941) );
  XOR U10764 ( .A(n11943), .B(n11944), .Z(n10622) );
  NOR U10765 ( .A(n11945), .B(n11943), .Z(n11944) );
  XOR U10766 ( .A(n11946), .B(n11947), .Z(n10623) );
  NOR U10767 ( .A(n11948), .B(n11946), .Z(n11947) );
  XOR U10768 ( .A(n11949), .B(n11950), .Z(n10502) );
  NOR U10769 ( .A(n11951), .B(n11949), .Z(n11950) );
  XOR U10770 ( .A(n11952), .B(n11953), .Z(n10638) );
  NOR U10771 ( .A(n11954), .B(n11952), .Z(n11953) );
  XOR U10772 ( .A(n11955), .B(n11956), .Z(n10633) );
  NOR U10773 ( .A(n11957), .B(n11955), .Z(n11956) );
  XOR U10774 ( .A(n11958), .B(n11959), .Z(n10634) );
  NOR U10775 ( .A(n11960), .B(n11958), .Z(n11959) );
  XOR U10776 ( .A(n11961), .B(n11962), .Z(n10493) );
  NOR U10777 ( .A(n11963), .B(n11961), .Z(n11962) );
  XOR U10778 ( .A(n11964), .B(n11965), .Z(n10649) );
  NOR U10779 ( .A(n11966), .B(n11964), .Z(n11965) );
  XOR U10780 ( .A(n11967), .B(n11968), .Z(n10644) );
  NOR U10781 ( .A(n11969), .B(n11967), .Z(n11968) );
  XOR U10782 ( .A(n11970), .B(n11971), .Z(n10645) );
  NOR U10783 ( .A(n11972), .B(n11970), .Z(n11971) );
  XOR U10784 ( .A(n11973), .B(n11974), .Z(n10484) );
  NOR U10785 ( .A(n11975), .B(n11973), .Z(n11974) );
  XOR U10786 ( .A(n11976), .B(n11977), .Z(n10660) );
  NOR U10787 ( .A(n11978), .B(n11976), .Z(n11977) );
  XOR U10788 ( .A(n11979), .B(n11980), .Z(n10655) );
  NOR U10789 ( .A(n11981), .B(n11979), .Z(n11980) );
  XOR U10790 ( .A(n11982), .B(n11983), .Z(n10656) );
  NOR U10791 ( .A(n11984), .B(n11982), .Z(n11983) );
  XOR U10792 ( .A(n11985), .B(n11986), .Z(n10475) );
  NOR U10793 ( .A(n11987), .B(n11985), .Z(n11986) );
  XOR U10794 ( .A(n11988), .B(n11989), .Z(n10671) );
  NOR U10795 ( .A(n11990), .B(n11988), .Z(n11989) );
  XOR U10796 ( .A(n11991), .B(n11992), .Z(n10666) );
  NOR U10797 ( .A(n11993), .B(n11991), .Z(n11992) );
  XOR U10798 ( .A(n11994), .B(n11995), .Z(n10667) );
  NOR U10799 ( .A(n11996), .B(n11994), .Z(n11995) );
  XOR U10800 ( .A(n11997), .B(n11998), .Z(n10466) );
  NOR U10801 ( .A(n11999), .B(n11997), .Z(n11998) );
  XOR U10802 ( .A(n12000), .B(n12001), .Z(n10682) );
  NOR U10803 ( .A(n12002), .B(n12000), .Z(n12001) );
  XOR U10804 ( .A(n12003), .B(n12004), .Z(n10677) );
  NOR U10805 ( .A(n12005), .B(n12003), .Z(n12004) );
  XOR U10806 ( .A(n12006), .B(n12007), .Z(n10678) );
  NOR U10807 ( .A(n12008), .B(n12006), .Z(n12007) );
  XOR U10808 ( .A(n12009), .B(n12010), .Z(n10457) );
  NOR U10809 ( .A(n12011), .B(n12009), .Z(n12010) );
  XOR U10810 ( .A(n12012), .B(n12013), .Z(n10693) );
  NOR U10811 ( .A(n12014), .B(n12012), .Z(n12013) );
  XOR U10812 ( .A(n12015), .B(n12016), .Z(n10688) );
  NOR U10813 ( .A(n12017), .B(n12015), .Z(n12016) );
  XOR U10814 ( .A(n12018), .B(n12019), .Z(n10689) );
  NOR U10815 ( .A(n12020), .B(n12018), .Z(n12019) );
  XOR U10816 ( .A(n12021), .B(n12022), .Z(n10448) );
  NOR U10817 ( .A(n12023), .B(n12021), .Z(n12022) );
  XOR U10818 ( .A(n12024), .B(n12025), .Z(n10704) );
  NOR U10819 ( .A(n12026), .B(n12024), .Z(n12025) );
  XOR U10820 ( .A(n12027), .B(n12028), .Z(n10699) );
  NOR U10821 ( .A(n12029), .B(n12027), .Z(n12028) );
  XOR U10822 ( .A(n12030), .B(n12031), .Z(n10700) );
  NOR U10823 ( .A(n12032), .B(n12030), .Z(n12031) );
  XOR U10824 ( .A(n12033), .B(n12034), .Z(n10439) );
  NOR U10825 ( .A(n12035), .B(n12033), .Z(n12034) );
  XOR U10826 ( .A(n12036), .B(n12037), .Z(n10715) );
  NOR U10827 ( .A(n12038), .B(n12036), .Z(n12037) );
  XOR U10828 ( .A(n12039), .B(n12040), .Z(n10710) );
  NOR U10829 ( .A(n12041), .B(n12039), .Z(n12040) );
  XOR U10830 ( .A(n12042), .B(n12043), .Z(n10711) );
  NOR U10831 ( .A(n12044), .B(n12042), .Z(n12043) );
  XOR U10832 ( .A(n12045), .B(n12046), .Z(n10430) );
  NOR U10833 ( .A(n12047), .B(n12045), .Z(n12046) );
  XOR U10834 ( .A(n12048), .B(n12049), .Z(n10726) );
  NOR U10835 ( .A(n12050), .B(n12048), .Z(n12049) );
  XOR U10836 ( .A(n12051), .B(n12052), .Z(n10721) );
  NOR U10837 ( .A(n12053), .B(n12051), .Z(n12052) );
  XOR U10838 ( .A(n12054), .B(n12055), .Z(n10722) );
  NOR U10839 ( .A(n12056), .B(n12054), .Z(n12055) );
  XOR U10840 ( .A(n12057), .B(n12058), .Z(n10421) );
  NOR U10841 ( .A(n12059), .B(n12057), .Z(n12058) );
  XOR U10842 ( .A(n12060), .B(n12061), .Z(n10737) );
  NOR U10843 ( .A(n12062), .B(n12060), .Z(n12061) );
  XOR U10844 ( .A(n12063), .B(n12064), .Z(n10732) );
  NOR U10845 ( .A(n12065), .B(n12063), .Z(n12064) );
  XOR U10846 ( .A(n12066), .B(n12067), .Z(n10733) );
  NOR U10847 ( .A(n12068), .B(n12066), .Z(n12067) );
  XOR U10848 ( .A(n12069), .B(n12070), .Z(n10412) );
  NOR U10849 ( .A(n12071), .B(n12069), .Z(n12070) );
  XOR U10850 ( .A(n12072), .B(n12073), .Z(n10748) );
  NOR U10851 ( .A(n12074), .B(n12072), .Z(n12073) );
  XOR U10852 ( .A(n12075), .B(n12076), .Z(n10743) );
  NOR U10853 ( .A(n12077), .B(n12075), .Z(n12076) );
  XOR U10854 ( .A(n12078), .B(n12079), .Z(n10744) );
  NOR U10855 ( .A(n12080), .B(n12078), .Z(n12079) );
  XOR U10856 ( .A(n12081), .B(n12082), .Z(n10403) );
  NOR U10857 ( .A(n12083), .B(n12081), .Z(n12082) );
  XOR U10858 ( .A(n12084), .B(n12085), .Z(n10759) );
  NOR U10859 ( .A(n12086), .B(n12084), .Z(n12085) );
  XOR U10860 ( .A(n12087), .B(n12088), .Z(n10754) );
  NOR U10861 ( .A(n12089), .B(n12087), .Z(n12088) );
  XOR U10862 ( .A(n12090), .B(n12091), .Z(n10755) );
  NOR U10863 ( .A(n12092), .B(n12090), .Z(n12091) );
  XOR U10864 ( .A(n12093), .B(n12094), .Z(n10394) );
  NOR U10865 ( .A(n12095), .B(n12093), .Z(n12094) );
  XOR U10866 ( .A(n12096), .B(n12097), .Z(n10770) );
  NOR U10867 ( .A(n12098), .B(n12096), .Z(n12097) );
  XOR U10868 ( .A(n12099), .B(n12100), .Z(n10765) );
  NOR U10869 ( .A(n12101), .B(n12099), .Z(n12100) );
  XOR U10870 ( .A(n12102), .B(n12103), .Z(n10766) );
  NOR U10871 ( .A(n12104), .B(n12102), .Z(n12103) );
  XOR U10872 ( .A(n12105), .B(n12106), .Z(n10385) );
  NOR U10873 ( .A(n12107), .B(n12105), .Z(n12106) );
  XOR U10874 ( .A(n12108), .B(n12109), .Z(n10781) );
  NOR U10875 ( .A(n12110), .B(n12108), .Z(n12109) );
  XOR U10876 ( .A(n12111), .B(n12112), .Z(n10776) );
  NOR U10877 ( .A(n12113), .B(n12111), .Z(n12112) );
  XOR U10878 ( .A(n12114), .B(n12115), .Z(n10777) );
  NOR U10879 ( .A(n12116), .B(n12114), .Z(n12115) );
  XOR U10880 ( .A(n12117), .B(n12118), .Z(n10376) );
  NOR U10881 ( .A(n12119), .B(n12117), .Z(n12118) );
  XOR U10882 ( .A(n12120), .B(n12121), .Z(n10792) );
  NOR U10883 ( .A(n12122), .B(n12120), .Z(n12121) );
  XOR U10884 ( .A(n12123), .B(n12124), .Z(n10787) );
  NOR U10885 ( .A(n12125), .B(n12123), .Z(n12124) );
  XOR U10886 ( .A(n12126), .B(n12127), .Z(n10788) );
  NOR U10887 ( .A(n12128), .B(n12126), .Z(n12127) );
  XOR U10888 ( .A(n12129), .B(n12130), .Z(n10367) );
  NOR U10889 ( .A(n12131), .B(n12129), .Z(n12130) );
  XOR U10890 ( .A(n12132), .B(n12133), .Z(n10803) );
  NOR U10891 ( .A(n12134), .B(n12132), .Z(n12133) );
  XOR U10892 ( .A(n12135), .B(n12136), .Z(n10798) );
  NOR U10893 ( .A(n12137), .B(n12135), .Z(n12136) );
  XOR U10894 ( .A(n12138), .B(n12139), .Z(n10799) );
  NOR U10895 ( .A(n12140), .B(n12138), .Z(n12139) );
  XOR U10896 ( .A(n12141), .B(n12142), .Z(n10358) );
  NOR U10897 ( .A(n12143), .B(n12141), .Z(n12142) );
  XOR U10898 ( .A(n12144), .B(n12145), .Z(n10814) );
  NOR U10899 ( .A(n12146), .B(n12144), .Z(n12145) );
  XOR U10900 ( .A(n12147), .B(n12148), .Z(n10809) );
  NOR U10901 ( .A(n12149), .B(n12147), .Z(n12148) );
  XOR U10902 ( .A(n12150), .B(n12151), .Z(n10810) );
  NOR U10903 ( .A(n12152), .B(n12150), .Z(n12151) );
  XOR U10904 ( .A(n12153), .B(n12154), .Z(n10349) );
  NOR U10905 ( .A(n12155), .B(n12153), .Z(n12154) );
  XOR U10906 ( .A(n12156), .B(n12157), .Z(n10825) );
  NOR U10907 ( .A(n12158), .B(n12156), .Z(n12157) );
  XOR U10908 ( .A(n12159), .B(n12160), .Z(n10820) );
  NOR U10909 ( .A(n12161), .B(n12159), .Z(n12160) );
  XOR U10910 ( .A(n12162), .B(n12163), .Z(n10821) );
  NOR U10911 ( .A(n12164), .B(n12162), .Z(n12163) );
  XOR U10912 ( .A(n12165), .B(n12166), .Z(n10340) );
  NOR U10913 ( .A(n12167), .B(n12165), .Z(n12166) );
  XOR U10914 ( .A(n12168), .B(n12169), .Z(n10836) );
  NOR U10915 ( .A(n12170), .B(n12168), .Z(n12169) );
  XOR U10916 ( .A(n12171), .B(n12172), .Z(n10831) );
  NOR U10917 ( .A(n12173), .B(n12171), .Z(n12172) );
  XOR U10918 ( .A(n12174), .B(n12175), .Z(n10832) );
  NOR U10919 ( .A(n12176), .B(n12174), .Z(n12175) );
  XOR U10920 ( .A(n12177), .B(n12178), .Z(n10331) );
  NOR U10921 ( .A(n12179), .B(n12177), .Z(n12178) );
  XOR U10922 ( .A(n12180), .B(n12181), .Z(n10847) );
  NOR U10923 ( .A(n12182), .B(n12180), .Z(n12181) );
  XOR U10924 ( .A(n12183), .B(n12184), .Z(n10842) );
  NOR U10925 ( .A(n12185), .B(n12183), .Z(n12184) );
  XOR U10926 ( .A(n12186), .B(n12187), .Z(n10843) );
  NOR U10927 ( .A(n12188), .B(n12186), .Z(n12187) );
  XOR U10928 ( .A(n12189), .B(n12190), .Z(n10322) );
  NOR U10929 ( .A(n12191), .B(n12189), .Z(n12190) );
  XOR U10930 ( .A(n12192), .B(n12193), .Z(n10858) );
  NOR U10931 ( .A(n12194), .B(n12192), .Z(n12193) );
  XOR U10932 ( .A(n12195), .B(n12196), .Z(n10853) );
  NOR U10933 ( .A(n12197), .B(n12195), .Z(n12196) );
  XOR U10934 ( .A(n12198), .B(n12199), .Z(n10854) );
  NOR U10935 ( .A(n12200), .B(n12198), .Z(n12199) );
  XOR U10936 ( .A(n12201), .B(n12202), .Z(n10313) );
  NOR U10937 ( .A(n12203), .B(n12201), .Z(n12202) );
  XOR U10938 ( .A(n12204), .B(n12205), .Z(n10869) );
  NOR U10939 ( .A(n12206), .B(n12204), .Z(n12205) );
  XOR U10940 ( .A(n12207), .B(n12208), .Z(n10864) );
  NOR U10941 ( .A(n12209), .B(n12207), .Z(n12208) );
  XOR U10942 ( .A(n12210), .B(n12211), .Z(n10865) );
  NOR U10943 ( .A(n12212), .B(n12210), .Z(n12211) );
  XOR U10944 ( .A(n12213), .B(n12214), .Z(n10304) );
  NOR U10945 ( .A(n12215), .B(n12213), .Z(n12214) );
  XOR U10946 ( .A(n12216), .B(n12217), .Z(n10880) );
  NOR U10947 ( .A(n12218), .B(n12216), .Z(n12217) );
  XOR U10948 ( .A(n12219), .B(n12220), .Z(n10875) );
  NOR U10949 ( .A(n12221), .B(n12219), .Z(n12220) );
  XOR U10950 ( .A(n12222), .B(n12223), .Z(n10876) );
  NOR U10951 ( .A(n12224), .B(n12222), .Z(n12223) );
  XOR U10952 ( .A(n12225), .B(n12226), .Z(n10295) );
  NOR U10953 ( .A(n12227), .B(n12225), .Z(n12226) );
  XOR U10954 ( .A(n12228), .B(n12229), .Z(n10891) );
  NOR U10955 ( .A(n12230), .B(n12228), .Z(n12229) );
  XOR U10956 ( .A(n12231), .B(n12232), .Z(n10886) );
  NOR U10957 ( .A(n12233), .B(n12231), .Z(n12232) );
  XOR U10958 ( .A(n12234), .B(n12235), .Z(n10887) );
  NOR U10959 ( .A(n12236), .B(n12234), .Z(n12235) );
  XOR U10960 ( .A(n12237), .B(n12238), .Z(n10286) );
  NOR U10961 ( .A(n12239), .B(n12237), .Z(n12238) );
  XOR U10962 ( .A(n12240), .B(n12241), .Z(n10260) );
  NOR U10963 ( .A(n12242), .B(n12240), .Z(n12241) );
  XOR U10964 ( .A(n12243), .B(n12244), .Z(n10265) );
  NOR U10965 ( .A(n12245), .B(n12243), .Z(n12244) );
  IV U10966 ( .A(n10267), .Z(n11579) );
  XNOR U10967 ( .A(n12246), .B(n12247), .Z(n10267) );
  NOR U10968 ( .A(n12248), .B(n12246), .Z(n12247) );
  XOR U10969 ( .A(n12249), .B(n12250), .Z(n10277) );
  NOR U10970 ( .A(n12251), .B(n12249), .Z(n12250) );
  IV U10971 ( .A(n10897), .Z(n11578) );
  XOR U10972 ( .A(n12252), .B(n12253), .Z(n10897) );
  NOR U10973 ( .A(n60), .B(n12254), .Z(n12253) );
  IV U10974 ( .A(n12252), .Z(n12254) );
  XOR U10975 ( .A(n12255), .B(n12256), .Z(n10899) );
  AND U10976 ( .A(n12257), .B(n12258), .Z(n12256) );
  XOR U10977 ( .A(n12255), .B(n63), .Z(n12258) );
  XOR U10978 ( .A(n11576), .B(n11575), .Z(n63) );
  XNOR U10979 ( .A(n11573), .B(n11572), .Z(n11575) );
  XNOR U10980 ( .A(n11570), .B(n11569), .Z(n11572) );
  XNOR U10981 ( .A(n11567), .B(n11566), .Z(n11569) );
  XNOR U10982 ( .A(n11564), .B(n11563), .Z(n11566) );
  XNOR U10983 ( .A(n11561), .B(n11560), .Z(n11563) );
  XNOR U10984 ( .A(n11558), .B(n11557), .Z(n11560) );
  XNOR U10985 ( .A(n11555), .B(n11554), .Z(n11557) );
  XNOR U10986 ( .A(n11552), .B(n11551), .Z(n11554) );
  XNOR U10987 ( .A(n11549), .B(n11548), .Z(n11551) );
  XNOR U10988 ( .A(n11546), .B(n11545), .Z(n11548) );
  XNOR U10989 ( .A(n11543), .B(n11542), .Z(n11545) );
  XNOR U10990 ( .A(n11540), .B(n11539), .Z(n11542) );
  XNOR U10991 ( .A(n11537), .B(n11536), .Z(n11539) );
  XNOR U10992 ( .A(n11534), .B(n11533), .Z(n11536) );
  XNOR U10993 ( .A(n11531), .B(n11530), .Z(n11533) );
  XNOR U10994 ( .A(n11528), .B(n11527), .Z(n11530) );
  XNOR U10995 ( .A(n11525), .B(n11524), .Z(n11527) );
  XNOR U10996 ( .A(n11522), .B(n11521), .Z(n11524) );
  XNOR U10997 ( .A(n11519), .B(n11518), .Z(n11521) );
  XNOR U10998 ( .A(n11516), .B(n11515), .Z(n11518) );
  XNOR U10999 ( .A(n11513), .B(n11512), .Z(n11515) );
  XNOR U11000 ( .A(n11510), .B(n11509), .Z(n11512) );
  XNOR U11001 ( .A(n11507), .B(n11506), .Z(n11509) );
  XNOR U11002 ( .A(n11504), .B(n11503), .Z(n11506) );
  XNOR U11003 ( .A(n11501), .B(n11500), .Z(n11503) );
  XNOR U11004 ( .A(n11498), .B(n11497), .Z(n11500) );
  XNOR U11005 ( .A(n11495), .B(n11494), .Z(n11497) );
  XNOR U11006 ( .A(n11492), .B(n11491), .Z(n11494) );
  XNOR U11007 ( .A(n11489), .B(n11488), .Z(n11491) );
  XNOR U11008 ( .A(n11486), .B(n11485), .Z(n11488) );
  XNOR U11009 ( .A(n11483), .B(n11482), .Z(n11485) );
  XNOR U11010 ( .A(n11480), .B(n11479), .Z(n11482) );
  XNOR U11011 ( .A(n11477), .B(n11476), .Z(n11479) );
  XNOR U11012 ( .A(n11474), .B(n11473), .Z(n11476) );
  XNOR U11013 ( .A(n11471), .B(n11470), .Z(n11473) );
  XNOR U11014 ( .A(n11468), .B(n11467), .Z(n11470) );
  XNOR U11015 ( .A(n11465), .B(n11464), .Z(n11467) );
  XNOR U11016 ( .A(n11462), .B(n11461), .Z(n11464) );
  XNOR U11017 ( .A(n11459), .B(n11458), .Z(n11461) );
  XNOR U11018 ( .A(n11456), .B(n11455), .Z(n11458) );
  XNOR U11019 ( .A(n11453), .B(n11452), .Z(n11455) );
  XNOR U11020 ( .A(n11450), .B(n11449), .Z(n11452) );
  XNOR U11021 ( .A(n11447), .B(n11446), .Z(n11449) );
  XNOR U11022 ( .A(n11444), .B(n11443), .Z(n11446) );
  XNOR U11023 ( .A(n11441), .B(n11440), .Z(n11443) );
  XNOR U11024 ( .A(n11438), .B(n11437), .Z(n11440) );
  XNOR U11025 ( .A(n11435), .B(n11434), .Z(n11437) );
  XNOR U11026 ( .A(n11432), .B(n11431), .Z(n11434) );
  XNOR U11027 ( .A(n11429), .B(n11428), .Z(n11431) );
  XNOR U11028 ( .A(n11426), .B(n11425), .Z(n11428) );
  XNOR U11029 ( .A(n11423), .B(n11422), .Z(n11425) );
  XNOR U11030 ( .A(n11420), .B(n11419), .Z(n11422) );
  XNOR U11031 ( .A(n11417), .B(n11416), .Z(n11419) );
  XNOR U11032 ( .A(n11414), .B(n11413), .Z(n11416) );
  XNOR U11033 ( .A(n11411), .B(n11410), .Z(n11413) );
  XNOR U11034 ( .A(n11408), .B(n11407), .Z(n11410) );
  XNOR U11035 ( .A(n11405), .B(n11404), .Z(n11407) );
  XNOR U11036 ( .A(n11402), .B(n11401), .Z(n11404) );
  XNOR U11037 ( .A(n11399), .B(n11398), .Z(n11401) );
  XNOR U11038 ( .A(n11396), .B(n11395), .Z(n11398) );
  XNOR U11039 ( .A(n11393), .B(n11392), .Z(n11395) );
  XNOR U11040 ( .A(n11390), .B(n11389), .Z(n11392) );
  XNOR U11041 ( .A(n11387), .B(n11386), .Z(n11389) );
  XNOR U11042 ( .A(n11384), .B(n11383), .Z(n11386) );
  XNOR U11043 ( .A(n11381), .B(n11380), .Z(n11383) );
  XNOR U11044 ( .A(n11378), .B(n11377), .Z(n11380) );
  XNOR U11045 ( .A(n11375), .B(n11374), .Z(n11377) );
  XNOR U11046 ( .A(n11372), .B(n11371), .Z(n11374) );
  XNOR U11047 ( .A(n11369), .B(n11368), .Z(n11371) );
  XNOR U11048 ( .A(n11366), .B(n11365), .Z(n11368) );
  XNOR U11049 ( .A(n11363), .B(n11362), .Z(n11365) );
  XNOR U11050 ( .A(n11360), .B(n11359), .Z(n11362) );
  XNOR U11051 ( .A(n11357), .B(n11356), .Z(n11359) );
  XNOR U11052 ( .A(n11354), .B(n11353), .Z(n11356) );
  XNOR U11053 ( .A(n11351), .B(n11350), .Z(n11353) );
  XNOR U11054 ( .A(n11348), .B(n11347), .Z(n11350) );
  XNOR U11055 ( .A(n11345), .B(n11344), .Z(n11347) );
  XNOR U11056 ( .A(n11342), .B(n11341), .Z(n11344) );
  XNOR U11057 ( .A(n11339), .B(n11338), .Z(n11341) );
  XNOR U11058 ( .A(n11336), .B(n11335), .Z(n11338) );
  XNOR U11059 ( .A(n11333), .B(n11332), .Z(n11335) );
  XNOR U11060 ( .A(n11330), .B(n11329), .Z(n11332) );
  XNOR U11061 ( .A(n11327), .B(n11326), .Z(n11329) );
  XNOR U11062 ( .A(n11324), .B(n11323), .Z(n11326) );
  XNOR U11063 ( .A(n11321), .B(n11320), .Z(n11323) );
  XNOR U11064 ( .A(n11318), .B(n11317), .Z(n11320) );
  XNOR U11065 ( .A(n11315), .B(n11314), .Z(n11317) );
  XNOR U11066 ( .A(n11312), .B(n11311), .Z(n11314) );
  XNOR U11067 ( .A(n11309), .B(n11308), .Z(n11311) );
  XNOR U11068 ( .A(n11306), .B(n11305), .Z(n11308) );
  XNOR U11069 ( .A(n11303), .B(n11302), .Z(n11305) );
  XNOR U11070 ( .A(n11300), .B(n11299), .Z(n11302) );
  XNOR U11071 ( .A(n11297), .B(n11296), .Z(n11299) );
  XNOR U11072 ( .A(n11294), .B(n11293), .Z(n11296) );
  XNOR U11073 ( .A(n11291), .B(n11290), .Z(n11293) );
  XNOR U11074 ( .A(n11288), .B(n11287), .Z(n11290) );
  XNOR U11075 ( .A(n11285), .B(n11284), .Z(n11287) );
  XNOR U11076 ( .A(n11282), .B(n11281), .Z(n11284) );
  XNOR U11077 ( .A(n11279), .B(n11278), .Z(n11281) );
  XNOR U11078 ( .A(n11276), .B(n11275), .Z(n11278) );
  XNOR U11079 ( .A(n11273), .B(n11272), .Z(n11275) );
  XNOR U11080 ( .A(n11270), .B(n11269), .Z(n11272) );
  XNOR U11081 ( .A(n11267), .B(n11266), .Z(n11269) );
  XNOR U11082 ( .A(n11264), .B(n11263), .Z(n11266) );
  XNOR U11083 ( .A(n11261), .B(n11260), .Z(n11263) );
  XNOR U11084 ( .A(n11258), .B(n11257), .Z(n11260) );
  XNOR U11085 ( .A(n11255), .B(n11254), .Z(n11257) );
  XNOR U11086 ( .A(n11252), .B(n11251), .Z(n11254) );
  XNOR U11087 ( .A(n11249), .B(n11248), .Z(n11251) );
  XNOR U11088 ( .A(n11246), .B(n11245), .Z(n11248) );
  XNOR U11089 ( .A(n11243), .B(n11242), .Z(n11245) );
  XNOR U11090 ( .A(n11240), .B(n11239), .Z(n11242) );
  XNOR U11091 ( .A(n11237), .B(n11236), .Z(n11239) );
  XNOR U11092 ( .A(n11234), .B(n11233), .Z(n11236) );
  XNOR U11093 ( .A(n11231), .B(n11230), .Z(n11233) );
  XNOR U11094 ( .A(n11228), .B(n11227), .Z(n11230) );
  XNOR U11095 ( .A(n11225), .B(n11224), .Z(n11227) );
  XNOR U11096 ( .A(n11222), .B(n11221), .Z(n11224) );
  XNOR U11097 ( .A(n11219), .B(n11218), .Z(n11221) );
  XNOR U11098 ( .A(n11216), .B(n11215), .Z(n11218) );
  XNOR U11099 ( .A(n11213), .B(n11212), .Z(n11215) );
  XNOR U11100 ( .A(n11210), .B(n11209), .Z(n11212) );
  XNOR U11101 ( .A(n11207), .B(n11206), .Z(n11209) );
  XNOR U11102 ( .A(n11204), .B(n11203), .Z(n11206) );
  XNOR U11103 ( .A(n11201), .B(n11200), .Z(n11203) );
  XNOR U11104 ( .A(n11198), .B(n11197), .Z(n11200) );
  XNOR U11105 ( .A(n11195), .B(n11194), .Z(n11197) );
  XNOR U11106 ( .A(n11192), .B(n11190), .Z(n11194) );
  XNOR U11107 ( .A(n11191), .B(n10912), .Z(n11190) );
  XNOR U11108 ( .A(n10913), .B(n10910), .Z(n10912) );
  XNOR U11109 ( .A(n10911), .B(n10914), .Z(n10910) );
  XNOR U11110 ( .A(n10915), .B(n11185), .Z(n10914) );
  XNOR U11111 ( .A(n10922), .B(n11184), .Z(n11185) );
  XNOR U11112 ( .A(n11177), .B(n11181), .Z(n11184) );
  XNOR U11113 ( .A(n11176), .B(n11174), .Z(n11181) );
  XNOR U11114 ( .A(n11175), .B(n11173), .Z(n11174) );
  XNOR U11115 ( .A(n10929), .B(n11168), .Z(n11173) );
  XOR U11116 ( .A(n10928), .B(n11166), .Z(n11168) );
  XNOR U11117 ( .A(n11167), .B(n11162), .Z(n11166) );
  XOR U11118 ( .A(n11163), .B(n10944), .Z(n11162) );
  XOR U11119 ( .A(n10945), .B(n11161), .Z(n10944) );
  XOR U11120 ( .A(n10938), .B(n11156), .Z(n11161) );
  XOR U11121 ( .A(n10940), .B(n11155), .Z(n11156) );
  XOR U11122 ( .A(n11152), .B(n10943), .Z(n11155) );
  AND U11123 ( .A(n12259), .B(n12260), .Z(n10943) );
  XOR U11124 ( .A(n11151), .B(n11142), .Z(n11152) );
  AND U11125 ( .A(n12261), .B(n12262), .Z(n11142) );
  XOR U11126 ( .A(n11148), .B(n11141), .Z(n11151) );
  AND U11127 ( .A(n12263), .B(n12264), .Z(n11141) );
  XOR U11128 ( .A(n11147), .B(n11140), .Z(n11148) );
  AND U11129 ( .A(n12265), .B(n12266), .Z(n11140) );
  XNOR U11130 ( .A(n11109), .B(n11139), .Z(n11147) );
  AND U11131 ( .A(n12267), .B(n12268), .Z(n11139) );
  XNOR U11132 ( .A(n11134), .B(n11110), .Z(n11109) );
  AND U11133 ( .A(n12269), .B(n12270), .Z(n11110) );
  XOR U11134 ( .A(n11133), .B(n11107), .Z(n11134) );
  AND U11135 ( .A(n12271), .B(n12272), .Z(n11107) );
  XOR U11136 ( .A(n11138), .B(n11114), .Z(n11133) );
  AND U11137 ( .A(n12273), .B(n12274), .Z(n11114) );
  XNOR U11138 ( .A(n11121), .B(n11113), .Z(n11138) );
  AND U11139 ( .A(n12275), .B(n12276), .Z(n11113) );
  XNOR U11140 ( .A(n11130), .B(n11122), .Z(n11121) );
  AND U11141 ( .A(n12277), .B(n12278), .Z(n11122) );
  XOR U11142 ( .A(n11129), .B(n11119), .Z(n11130) );
  AND U11143 ( .A(n12279), .B(n12280), .Z(n11119) );
  XOR U11144 ( .A(n11137), .B(n11118), .Z(n11129) );
  AND U11145 ( .A(n12281), .B(n12282), .Z(n11118) );
  XNOR U11146 ( .A(n11074), .B(n11117), .Z(n11137) );
  AND U11147 ( .A(n12283), .B(n12284), .Z(n11117) );
  XNOR U11148 ( .A(n11102), .B(n11075), .Z(n11074) );
  AND U11149 ( .A(n12285), .B(n12286), .Z(n11075) );
  XOR U11150 ( .A(n11101), .B(n11072), .Z(n11102) );
  AND U11151 ( .A(n12287), .B(n12288), .Z(n11072) );
  XOR U11152 ( .A(n11106), .B(n11071), .Z(n11101) );
  AND U11153 ( .A(n12289), .B(n12290), .Z(n11071) );
  XNOR U11154 ( .A(n11084), .B(n11070), .Z(n11106) );
  AND U11155 ( .A(n12291), .B(n12292), .Z(n11070) );
  XNOR U11156 ( .A(n11098), .B(n11085), .Z(n11084) );
  AND U11157 ( .A(n12293), .B(n12294), .Z(n11085) );
  XOR U11158 ( .A(n11097), .B(n11082), .Z(n11098) );
  AND U11159 ( .A(n12295), .B(n12296), .Z(n11082) );
  XOR U11160 ( .A(n11105), .B(n11081), .Z(n11097) );
  AND U11161 ( .A(n12297), .B(n12298), .Z(n11081) );
  XNOR U11162 ( .A(n11089), .B(n11080), .Z(n11105) );
  AND U11163 ( .A(n12299), .B(n12300), .Z(n11080) );
  XNOR U11164 ( .A(n11062), .B(n11090), .Z(n11089) );
  AND U11165 ( .A(n12301), .B(n12302), .Z(n11090) );
  XOR U11166 ( .A(n11060), .B(n11061), .Z(n11062) );
  AND U11167 ( .A(n12303), .B(n12304), .Z(n11061) );
  XOR U11168 ( .A(n11067), .B(n11059), .Z(n11060) );
  AND U11169 ( .A(n12305), .B(n12306), .Z(n11059) );
  XNOR U11170 ( .A(n10976), .B(n11066), .Z(n11067) );
  AND U11171 ( .A(n12307), .B(n12308), .Z(n11066) );
  XNOR U11172 ( .A(n11056), .B(n10977), .Z(n10976) );
  AND U11173 ( .A(n12309), .B(n12310), .Z(n10977) );
  XOR U11174 ( .A(n11055), .B(n10974), .Z(n11056) );
  AND U11175 ( .A(n12311), .B(n12312), .Z(n10974) );
  XOR U11176 ( .A(n11065), .B(n10973), .Z(n11055) );
  AND U11177 ( .A(n12313), .B(n12314), .Z(n10973) );
  XNOR U11178 ( .A(n10984), .B(n10972), .Z(n11065) );
  AND U11179 ( .A(n12315), .B(n12316), .Z(n10972) );
  XNOR U11180 ( .A(n11048), .B(n10985), .Z(n10984) );
  AND U11181 ( .A(n12317), .B(n12318), .Z(n10985) );
  XOR U11182 ( .A(n11047), .B(n10982), .Z(n11048) );
  AND U11183 ( .A(n12319), .B(n12320), .Z(n10982) );
  XOR U11184 ( .A(n11044), .B(n10981), .Z(n11047) );
  AND U11185 ( .A(n12321), .B(n12322), .Z(n10981) );
  XNOR U11186 ( .A(n10998), .B(n10980), .Z(n11044) );
  AND U11187 ( .A(n12323), .B(n12324), .Z(n10980) );
  XNOR U11188 ( .A(n11005), .B(n10999), .Z(n10998) );
  AND U11189 ( .A(n12325), .B(n12326), .Z(n10999) );
  XOR U11190 ( .A(n11004), .B(n10996), .Z(n11005) );
  AND U11191 ( .A(n12327), .B(n12328), .Z(n10996) );
  XOR U11192 ( .A(n11043), .B(n10995), .Z(n11004) );
  AND U11193 ( .A(n12329), .B(n12330), .Z(n10995) );
  XNOR U11194 ( .A(n11016), .B(n10994), .Z(n11043) );
  AND U11195 ( .A(n12331), .B(n12332), .Z(n10994) );
  XNOR U11196 ( .A(n11023), .B(n11017), .Z(n11016) );
  AND U11197 ( .A(n12333), .B(n12334), .Z(n11017) );
  XOR U11198 ( .A(n11022), .B(n11014), .Z(n11023) );
  AND U11199 ( .A(n12335), .B(n12336), .Z(n11014) );
  XOR U11200 ( .A(n11042), .B(n11013), .Z(n11022) );
  AND U11201 ( .A(n12337), .B(n12338), .Z(n11013) );
  XNOR U11202 ( .A(n12339), .B(n12340), .Z(n11042) );
  XOR U11203 ( .A(n12341), .B(n12342), .Z(n12340) );
  XOR U11204 ( .A(n12343), .B(n12344), .Z(n12342) );
  XNOR U11205 ( .A(n11040), .B(n11033), .Z(n12344) );
  XNOR U11206 ( .A(n12345), .B(n12346), .Z(n11033) );
  AND U11207 ( .A(n12347), .B(n12348), .Z(n12346) );
  NOR U11208 ( .A(n12349), .B(n12350), .Z(n12348) );
  NOR U11209 ( .A(n12351), .B(n12352), .Z(n12347) );
  AND U11210 ( .A(n12353), .B(n12354), .Z(n12352) );
  AND U11211 ( .A(n12355), .B(n12356), .Z(n12345) );
  NOR U11212 ( .A(n12357), .B(n12358), .Z(n12356) );
  AND U11213 ( .A(n12350), .B(n12359), .Z(n12358) );
  AND U11214 ( .A(n12351), .B(n12360), .Z(n12357) );
  NOR U11215 ( .A(n12361), .B(n12362), .Z(n12355) );
  XOR U11216 ( .A(n12363), .B(n12364), .Z(n12362) );
  AND U11217 ( .A(n12365), .B(n12366), .Z(n12364) );
  NOR U11218 ( .A(n12367), .B(n12368), .Z(n12366) );
  NOR U11219 ( .A(n12369), .B(n12370), .Z(n12365) );
  AND U11220 ( .A(n12371), .B(n12372), .Z(n12370) );
  AND U11221 ( .A(n12373), .B(n12374), .Z(n12363) );
  NOR U11222 ( .A(n12375), .B(n12376), .Z(n12374) );
  AND U11223 ( .A(n12368), .B(n12377), .Z(n12376) );
  AND U11224 ( .A(n12369), .B(n12378), .Z(n12375) );
  NOR U11225 ( .A(n12379), .B(n12380), .Z(n12373) );
  XOR U11226 ( .A(n12381), .B(n12382), .Z(n12380) );
  AND U11227 ( .A(n12383), .B(n12384), .Z(n12382) );
  NOR U11228 ( .A(n12385), .B(n12386), .Z(n12384) );
  NOR U11229 ( .A(n12387), .B(n12388), .Z(n12383) );
  AND U11230 ( .A(n12389), .B(n12390), .Z(n12388) );
  AND U11231 ( .A(n12391), .B(n12392), .Z(n12381) );
  NOR U11232 ( .A(n12393), .B(n12394), .Z(n12392) );
  AND U11233 ( .A(n12386), .B(n12395), .Z(n12394) );
  AND U11234 ( .A(n12387), .B(n12396), .Z(n12393) );
  NOR U11235 ( .A(n12397), .B(n12398), .Z(n12391) );
  XOR U11236 ( .A(n12399), .B(n12400), .Z(n12398) );
  AND U11237 ( .A(n12401), .B(n12402), .Z(n12400) );
  NOR U11238 ( .A(n12403), .B(n12404), .Z(n12402) );
  NOR U11239 ( .A(n12405), .B(n12406), .Z(n12401) );
  AND U11240 ( .A(n12407), .B(n12408), .Z(n12406) );
  AND U11241 ( .A(n12409), .B(n12410), .Z(n12399) );
  NOR U11242 ( .A(n12411), .B(n12412), .Z(n12410) );
  AND U11243 ( .A(n12404), .B(n12413), .Z(n12412) );
  AND U11244 ( .A(n12405), .B(n12414), .Z(n12411) );
  NOR U11245 ( .A(n12415), .B(n12416), .Z(n12409) );
  AND U11246 ( .A(n12417), .B(n12418), .Z(n12416) );
  AND U11247 ( .A(n12419), .B(n12420), .Z(n12418) );
  AND U11248 ( .A(n12421), .B(n12422), .Z(n12420) );
  AND U11249 ( .A(n12423), .B(n12424), .Z(n12422) );
  NOR U11250 ( .A(n12425), .B(n12426), .Z(n12423) );
  NOR U11251 ( .A(n12427), .B(n12428), .Z(n12421) );
  AND U11252 ( .A(n12429), .B(n12430), .Z(n12419) );
  NOR U11253 ( .A(n12431), .B(n12432), .Z(n12430) );
  NOR U11254 ( .A(n12433), .B(n12434), .Z(n12429) );
  AND U11255 ( .A(n12435), .B(n12436), .Z(n12417) );
  AND U11256 ( .A(n12437), .B(n12438), .Z(n12436) );
  NOR U11257 ( .A(n12439), .B(n12440), .Z(n12438) );
  NOR U11258 ( .A(n12441), .B(n12442), .Z(n12437) );
  AND U11259 ( .A(n12443), .B(n12444), .Z(n12435) );
  NOR U11260 ( .A(n12445), .B(n12446), .Z(n12444) );
  NOR U11261 ( .A(n12447), .B(n12448), .Z(n12443) );
  AND U11262 ( .A(n12403), .B(n12449), .Z(n12415) );
  AND U11263 ( .A(n12385), .B(n12450), .Z(n12397) );
  AND U11264 ( .A(n12367), .B(n12451), .Z(n12379) );
  AND U11265 ( .A(n12349), .B(n12452), .Z(n12361) );
  AND U11266 ( .A(n12453), .B(n12454), .Z(n11040) );
  XOR U11267 ( .A(n11038), .B(n11039), .Z(n12343) );
  AND U11268 ( .A(n12455), .B(n12456), .Z(n11039) );
  AND U11269 ( .A(n12457), .B(n12458), .Z(n11038) );
  XOR U11270 ( .A(n12459), .B(n12460), .Z(n12341) );
  XOR U11271 ( .A(n11034), .B(n11035), .Z(n12460) );
  AND U11272 ( .A(n12461), .B(n12462), .Z(n11035) );
  AND U11273 ( .A(n12463), .B(n12464), .Z(n11034) );
  XNOR U11274 ( .A(n11032), .B(n11031), .Z(n12459) );
  IV U11275 ( .A(n12465), .Z(n11031) );
  AND U11276 ( .A(n12466), .B(n12467), .Z(n12465) );
  AND U11277 ( .A(n12468), .B(n12469), .Z(n11032) );
  XNOR U11278 ( .A(n11041), .B(n11012), .Z(n12339) );
  AND U11279 ( .A(n12470), .B(n12471), .Z(n11012) );
  AND U11280 ( .A(n12472), .B(n12473), .Z(n11041) );
  XOR U11281 ( .A(n12474), .B(n12475), .Z(n10940) );
  AND U11282 ( .A(n12474), .B(n12476), .Z(n12475) );
  XOR U11283 ( .A(n12477), .B(n12478), .Z(n10938) );
  AND U11284 ( .A(n12477), .B(n12479), .Z(n12478) );
  IV U11285 ( .A(n10939), .Z(n10945) );
  XNOR U11286 ( .A(n12480), .B(n12481), .Z(n10939) );
  AND U11287 ( .A(n12480), .B(n12482), .Z(n12481) );
  XNOR U11288 ( .A(n12483), .B(n12484), .Z(n11163) );
  AND U11289 ( .A(n12483), .B(n12485), .Z(n12484) );
  XOR U11290 ( .A(n12486), .B(n12487), .Z(n11167) );
  AND U11291 ( .A(n12486), .B(n12488), .Z(n12487) );
  XNOR U11292 ( .A(n12489), .B(n12490), .Z(n10928) );
  AND U11293 ( .A(n12491), .B(n12489), .Z(n12490) );
  XOR U11294 ( .A(n12492), .B(n12493), .Z(n10929) );
  NOR U11295 ( .A(n12494), .B(n12492), .Z(n12493) );
  XOR U11296 ( .A(n12495), .B(n12496), .Z(n11175) );
  NOR U11297 ( .A(n12497), .B(n12495), .Z(n12496) );
  XOR U11298 ( .A(n12498), .B(n12499), .Z(n11176) );
  NOR U11299 ( .A(n12500), .B(n12498), .Z(n12499) );
  XOR U11300 ( .A(n12501), .B(n12502), .Z(n11177) );
  NOR U11301 ( .A(n12503), .B(n12501), .Z(n12502) );
  XOR U11302 ( .A(n12504), .B(n12505), .Z(n10922) );
  NOR U11303 ( .A(n12506), .B(n12504), .Z(n12505) );
  XOR U11304 ( .A(n12507), .B(n12508), .Z(n10915) );
  NOR U11305 ( .A(n12509), .B(n12507), .Z(n12508) );
  XOR U11306 ( .A(n12510), .B(n12511), .Z(n10911) );
  NOR U11307 ( .A(n12512), .B(n12510), .Z(n12511) );
  XOR U11308 ( .A(n12513), .B(n12514), .Z(n10913) );
  NOR U11309 ( .A(n12515), .B(n12513), .Z(n12514) );
  XOR U11310 ( .A(n12516), .B(n12517), .Z(n11191) );
  NOR U11311 ( .A(n12518), .B(n12516), .Z(n12517) );
  XOR U11312 ( .A(n12519), .B(n12520), .Z(n11192) );
  NOR U11313 ( .A(n12521), .B(n12519), .Z(n12520) );
  XOR U11314 ( .A(n12522), .B(n12523), .Z(n11195) );
  NOR U11315 ( .A(n12524), .B(n12522), .Z(n12523) );
  XOR U11316 ( .A(n12525), .B(n12526), .Z(n11198) );
  NOR U11317 ( .A(n12527), .B(n12525), .Z(n12526) );
  XOR U11318 ( .A(n12528), .B(n12529), .Z(n11201) );
  NOR U11319 ( .A(n12530), .B(n12528), .Z(n12529) );
  XOR U11320 ( .A(n12531), .B(n12532), .Z(n11204) );
  NOR U11321 ( .A(n12533), .B(n12531), .Z(n12532) );
  XOR U11322 ( .A(n12534), .B(n12535), .Z(n11207) );
  NOR U11323 ( .A(n12536), .B(n12534), .Z(n12535) );
  XOR U11324 ( .A(n12537), .B(n12538), .Z(n11210) );
  NOR U11325 ( .A(n12539), .B(n12537), .Z(n12538) );
  XOR U11326 ( .A(n12540), .B(n12541), .Z(n11213) );
  NOR U11327 ( .A(n12542), .B(n12540), .Z(n12541) );
  XOR U11328 ( .A(n12543), .B(n12544), .Z(n11216) );
  NOR U11329 ( .A(n12545), .B(n12543), .Z(n12544) );
  XOR U11330 ( .A(n12546), .B(n12547), .Z(n11219) );
  NOR U11331 ( .A(n12548), .B(n12546), .Z(n12547) );
  XOR U11332 ( .A(n12549), .B(n12550), .Z(n11222) );
  NOR U11333 ( .A(n12551), .B(n12549), .Z(n12550) );
  XOR U11334 ( .A(n12552), .B(n12553), .Z(n11225) );
  NOR U11335 ( .A(n12554), .B(n12552), .Z(n12553) );
  XOR U11336 ( .A(n12555), .B(n12556), .Z(n11228) );
  NOR U11337 ( .A(n12557), .B(n12555), .Z(n12556) );
  XOR U11338 ( .A(n12558), .B(n12559), .Z(n11231) );
  NOR U11339 ( .A(n12560), .B(n12558), .Z(n12559) );
  XOR U11340 ( .A(n12561), .B(n12562), .Z(n11234) );
  NOR U11341 ( .A(n12563), .B(n12561), .Z(n12562) );
  XOR U11342 ( .A(n12564), .B(n12565), .Z(n11237) );
  NOR U11343 ( .A(n12566), .B(n12564), .Z(n12565) );
  XOR U11344 ( .A(n12567), .B(n12568), .Z(n11240) );
  NOR U11345 ( .A(n12569), .B(n12567), .Z(n12568) );
  XOR U11346 ( .A(n12570), .B(n12571), .Z(n11243) );
  NOR U11347 ( .A(n12572), .B(n12570), .Z(n12571) );
  XOR U11348 ( .A(n12573), .B(n12574), .Z(n11246) );
  NOR U11349 ( .A(n12575), .B(n12573), .Z(n12574) );
  XOR U11350 ( .A(n12576), .B(n12577), .Z(n11249) );
  NOR U11351 ( .A(n12578), .B(n12576), .Z(n12577) );
  XOR U11352 ( .A(n12579), .B(n12580), .Z(n11252) );
  NOR U11353 ( .A(n12581), .B(n12579), .Z(n12580) );
  XOR U11354 ( .A(n12582), .B(n12583), .Z(n11255) );
  NOR U11355 ( .A(n12584), .B(n12582), .Z(n12583) );
  XOR U11356 ( .A(n12585), .B(n12586), .Z(n11258) );
  NOR U11357 ( .A(n12587), .B(n12585), .Z(n12586) );
  XOR U11358 ( .A(n12588), .B(n12589), .Z(n11261) );
  NOR U11359 ( .A(n12590), .B(n12588), .Z(n12589) );
  XOR U11360 ( .A(n12591), .B(n12592), .Z(n11264) );
  NOR U11361 ( .A(n12593), .B(n12591), .Z(n12592) );
  XOR U11362 ( .A(n12594), .B(n12595), .Z(n11267) );
  NOR U11363 ( .A(n12596), .B(n12594), .Z(n12595) );
  XOR U11364 ( .A(n12597), .B(n12598), .Z(n11270) );
  NOR U11365 ( .A(n12599), .B(n12597), .Z(n12598) );
  XOR U11366 ( .A(n12600), .B(n12601), .Z(n11273) );
  NOR U11367 ( .A(n12602), .B(n12600), .Z(n12601) );
  XOR U11368 ( .A(n12603), .B(n12604), .Z(n11276) );
  NOR U11369 ( .A(n12605), .B(n12603), .Z(n12604) );
  XOR U11370 ( .A(n12606), .B(n12607), .Z(n11279) );
  NOR U11371 ( .A(n12608), .B(n12606), .Z(n12607) );
  XOR U11372 ( .A(n12609), .B(n12610), .Z(n11282) );
  NOR U11373 ( .A(n12611), .B(n12609), .Z(n12610) );
  XOR U11374 ( .A(n12612), .B(n12613), .Z(n11285) );
  NOR U11375 ( .A(n12614), .B(n12612), .Z(n12613) );
  XOR U11376 ( .A(n12615), .B(n12616), .Z(n11288) );
  NOR U11377 ( .A(n12617), .B(n12615), .Z(n12616) );
  XOR U11378 ( .A(n12618), .B(n12619), .Z(n11291) );
  NOR U11379 ( .A(n12620), .B(n12618), .Z(n12619) );
  XOR U11380 ( .A(n12621), .B(n12622), .Z(n11294) );
  NOR U11381 ( .A(n12623), .B(n12621), .Z(n12622) );
  XOR U11382 ( .A(n12624), .B(n12625), .Z(n11297) );
  NOR U11383 ( .A(n12626), .B(n12624), .Z(n12625) );
  XOR U11384 ( .A(n12627), .B(n12628), .Z(n11300) );
  NOR U11385 ( .A(n12629), .B(n12627), .Z(n12628) );
  XOR U11386 ( .A(n12630), .B(n12631), .Z(n11303) );
  NOR U11387 ( .A(n12632), .B(n12630), .Z(n12631) );
  XOR U11388 ( .A(n12633), .B(n12634), .Z(n11306) );
  NOR U11389 ( .A(n12635), .B(n12633), .Z(n12634) );
  XOR U11390 ( .A(n12636), .B(n12637), .Z(n11309) );
  NOR U11391 ( .A(n12638), .B(n12636), .Z(n12637) );
  XOR U11392 ( .A(n12639), .B(n12640), .Z(n11312) );
  NOR U11393 ( .A(n12641), .B(n12639), .Z(n12640) );
  XOR U11394 ( .A(n12642), .B(n12643), .Z(n11315) );
  NOR U11395 ( .A(n12644), .B(n12642), .Z(n12643) );
  XOR U11396 ( .A(n12645), .B(n12646), .Z(n11318) );
  NOR U11397 ( .A(n12647), .B(n12645), .Z(n12646) );
  XOR U11398 ( .A(n12648), .B(n12649), .Z(n11321) );
  NOR U11399 ( .A(n12650), .B(n12648), .Z(n12649) );
  XOR U11400 ( .A(n12651), .B(n12652), .Z(n11324) );
  NOR U11401 ( .A(n12653), .B(n12651), .Z(n12652) );
  XOR U11402 ( .A(n12654), .B(n12655), .Z(n11327) );
  NOR U11403 ( .A(n12656), .B(n12654), .Z(n12655) );
  XOR U11404 ( .A(n12657), .B(n12658), .Z(n11330) );
  NOR U11405 ( .A(n12659), .B(n12657), .Z(n12658) );
  XOR U11406 ( .A(n12660), .B(n12661), .Z(n11333) );
  NOR U11407 ( .A(n12662), .B(n12660), .Z(n12661) );
  XOR U11408 ( .A(n12663), .B(n12664), .Z(n11336) );
  NOR U11409 ( .A(n12665), .B(n12663), .Z(n12664) );
  XOR U11410 ( .A(n12666), .B(n12667), .Z(n11339) );
  NOR U11411 ( .A(n12668), .B(n12666), .Z(n12667) );
  XOR U11412 ( .A(n12669), .B(n12670), .Z(n11342) );
  NOR U11413 ( .A(n12671), .B(n12669), .Z(n12670) );
  XOR U11414 ( .A(n12672), .B(n12673), .Z(n11345) );
  NOR U11415 ( .A(n12674), .B(n12672), .Z(n12673) );
  XOR U11416 ( .A(n12675), .B(n12676), .Z(n11348) );
  NOR U11417 ( .A(n12677), .B(n12675), .Z(n12676) );
  XOR U11418 ( .A(n12678), .B(n12679), .Z(n11351) );
  NOR U11419 ( .A(n12680), .B(n12678), .Z(n12679) );
  XOR U11420 ( .A(n12681), .B(n12682), .Z(n11354) );
  NOR U11421 ( .A(n12683), .B(n12681), .Z(n12682) );
  XOR U11422 ( .A(n12684), .B(n12685), .Z(n11357) );
  NOR U11423 ( .A(n12686), .B(n12684), .Z(n12685) );
  XOR U11424 ( .A(n12687), .B(n12688), .Z(n11360) );
  NOR U11425 ( .A(n12689), .B(n12687), .Z(n12688) );
  XOR U11426 ( .A(n12690), .B(n12691), .Z(n11363) );
  NOR U11427 ( .A(n12692), .B(n12690), .Z(n12691) );
  XOR U11428 ( .A(n12693), .B(n12694), .Z(n11366) );
  NOR U11429 ( .A(n12695), .B(n12693), .Z(n12694) );
  XOR U11430 ( .A(n12696), .B(n12697), .Z(n11369) );
  NOR U11431 ( .A(n12698), .B(n12696), .Z(n12697) );
  XOR U11432 ( .A(n12699), .B(n12700), .Z(n11372) );
  NOR U11433 ( .A(n12701), .B(n12699), .Z(n12700) );
  XOR U11434 ( .A(n12702), .B(n12703), .Z(n11375) );
  NOR U11435 ( .A(n12704), .B(n12702), .Z(n12703) );
  XOR U11436 ( .A(n12705), .B(n12706), .Z(n11378) );
  NOR U11437 ( .A(n12707), .B(n12705), .Z(n12706) );
  XOR U11438 ( .A(n12708), .B(n12709), .Z(n11381) );
  NOR U11439 ( .A(n12710), .B(n12708), .Z(n12709) );
  XOR U11440 ( .A(n12711), .B(n12712), .Z(n11384) );
  NOR U11441 ( .A(n12713), .B(n12711), .Z(n12712) );
  XOR U11442 ( .A(n12714), .B(n12715), .Z(n11387) );
  NOR U11443 ( .A(n12716), .B(n12714), .Z(n12715) );
  XOR U11444 ( .A(n12717), .B(n12718), .Z(n11390) );
  NOR U11445 ( .A(n12719), .B(n12717), .Z(n12718) );
  XOR U11446 ( .A(n12720), .B(n12721), .Z(n11393) );
  NOR U11447 ( .A(n12722), .B(n12720), .Z(n12721) );
  XOR U11448 ( .A(n12723), .B(n12724), .Z(n11396) );
  NOR U11449 ( .A(n12725), .B(n12723), .Z(n12724) );
  XOR U11450 ( .A(n12726), .B(n12727), .Z(n11399) );
  NOR U11451 ( .A(n12728), .B(n12726), .Z(n12727) );
  XOR U11452 ( .A(n12729), .B(n12730), .Z(n11402) );
  NOR U11453 ( .A(n12731), .B(n12729), .Z(n12730) );
  XOR U11454 ( .A(n12732), .B(n12733), .Z(n11405) );
  NOR U11455 ( .A(n12734), .B(n12732), .Z(n12733) );
  XOR U11456 ( .A(n12735), .B(n12736), .Z(n11408) );
  NOR U11457 ( .A(n12737), .B(n12735), .Z(n12736) );
  XOR U11458 ( .A(n12738), .B(n12739), .Z(n11411) );
  NOR U11459 ( .A(n12740), .B(n12738), .Z(n12739) );
  XOR U11460 ( .A(n12741), .B(n12742), .Z(n11414) );
  NOR U11461 ( .A(n12743), .B(n12741), .Z(n12742) );
  XOR U11462 ( .A(n12744), .B(n12745), .Z(n11417) );
  NOR U11463 ( .A(n12746), .B(n12744), .Z(n12745) );
  XOR U11464 ( .A(n12747), .B(n12748), .Z(n11420) );
  NOR U11465 ( .A(n12749), .B(n12747), .Z(n12748) );
  XOR U11466 ( .A(n12750), .B(n12751), .Z(n11423) );
  NOR U11467 ( .A(n12752), .B(n12750), .Z(n12751) );
  XOR U11468 ( .A(n12753), .B(n12754), .Z(n11426) );
  NOR U11469 ( .A(n12755), .B(n12753), .Z(n12754) );
  XOR U11470 ( .A(n12756), .B(n12757), .Z(n11429) );
  NOR U11471 ( .A(n12758), .B(n12756), .Z(n12757) );
  XOR U11472 ( .A(n12759), .B(n12760), .Z(n11432) );
  NOR U11473 ( .A(n12761), .B(n12759), .Z(n12760) );
  XOR U11474 ( .A(n12762), .B(n12763), .Z(n11435) );
  NOR U11475 ( .A(n12764), .B(n12762), .Z(n12763) );
  XOR U11476 ( .A(n12765), .B(n12766), .Z(n11438) );
  NOR U11477 ( .A(n12767), .B(n12765), .Z(n12766) );
  XOR U11478 ( .A(n12768), .B(n12769), .Z(n11441) );
  NOR U11479 ( .A(n12770), .B(n12768), .Z(n12769) );
  XOR U11480 ( .A(n12771), .B(n12772), .Z(n11444) );
  NOR U11481 ( .A(n12773), .B(n12771), .Z(n12772) );
  XOR U11482 ( .A(n12774), .B(n12775), .Z(n11447) );
  NOR U11483 ( .A(n12776), .B(n12774), .Z(n12775) );
  XOR U11484 ( .A(n12777), .B(n12778), .Z(n11450) );
  NOR U11485 ( .A(n12779), .B(n12777), .Z(n12778) );
  XOR U11486 ( .A(n12780), .B(n12781), .Z(n11453) );
  NOR U11487 ( .A(n12782), .B(n12780), .Z(n12781) );
  XOR U11488 ( .A(n12783), .B(n12784), .Z(n11456) );
  NOR U11489 ( .A(n12785), .B(n12783), .Z(n12784) );
  XOR U11490 ( .A(n12786), .B(n12787), .Z(n11459) );
  NOR U11491 ( .A(n12788), .B(n12786), .Z(n12787) );
  XOR U11492 ( .A(n12789), .B(n12790), .Z(n11462) );
  NOR U11493 ( .A(n12791), .B(n12789), .Z(n12790) );
  XOR U11494 ( .A(n12792), .B(n12793), .Z(n11465) );
  NOR U11495 ( .A(n12794), .B(n12792), .Z(n12793) );
  XOR U11496 ( .A(n12795), .B(n12796), .Z(n11468) );
  NOR U11497 ( .A(n12797), .B(n12795), .Z(n12796) );
  XOR U11498 ( .A(n12798), .B(n12799), .Z(n11471) );
  NOR U11499 ( .A(n12800), .B(n12798), .Z(n12799) );
  XOR U11500 ( .A(n12801), .B(n12802), .Z(n11474) );
  NOR U11501 ( .A(n12803), .B(n12801), .Z(n12802) );
  XOR U11502 ( .A(n12804), .B(n12805), .Z(n11477) );
  NOR U11503 ( .A(n12806), .B(n12804), .Z(n12805) );
  XOR U11504 ( .A(n12807), .B(n12808), .Z(n11480) );
  NOR U11505 ( .A(n12809), .B(n12807), .Z(n12808) );
  XOR U11506 ( .A(n12810), .B(n12811), .Z(n11483) );
  NOR U11507 ( .A(n12812), .B(n12810), .Z(n12811) );
  XOR U11508 ( .A(n12813), .B(n12814), .Z(n11486) );
  NOR U11509 ( .A(n12815), .B(n12813), .Z(n12814) );
  XOR U11510 ( .A(n12816), .B(n12817), .Z(n11489) );
  NOR U11511 ( .A(n12818), .B(n12816), .Z(n12817) );
  XOR U11512 ( .A(n12819), .B(n12820), .Z(n11492) );
  NOR U11513 ( .A(n12821), .B(n12819), .Z(n12820) );
  XOR U11514 ( .A(n12822), .B(n12823), .Z(n11495) );
  NOR U11515 ( .A(n12824), .B(n12822), .Z(n12823) );
  XOR U11516 ( .A(n12825), .B(n12826), .Z(n11498) );
  NOR U11517 ( .A(n12827), .B(n12825), .Z(n12826) );
  XOR U11518 ( .A(n12828), .B(n12829), .Z(n11501) );
  NOR U11519 ( .A(n12830), .B(n12828), .Z(n12829) );
  XOR U11520 ( .A(n12831), .B(n12832), .Z(n11504) );
  NOR U11521 ( .A(n12833), .B(n12831), .Z(n12832) );
  XOR U11522 ( .A(n12834), .B(n12835), .Z(n11507) );
  NOR U11523 ( .A(n12836), .B(n12834), .Z(n12835) );
  XOR U11524 ( .A(n12837), .B(n12838), .Z(n11510) );
  NOR U11525 ( .A(n12839), .B(n12837), .Z(n12838) );
  XOR U11526 ( .A(n12840), .B(n12841), .Z(n11513) );
  NOR U11527 ( .A(n12842), .B(n12840), .Z(n12841) );
  XOR U11528 ( .A(n12843), .B(n12844), .Z(n11516) );
  NOR U11529 ( .A(n12845), .B(n12843), .Z(n12844) );
  XOR U11530 ( .A(n12846), .B(n12847), .Z(n11519) );
  NOR U11531 ( .A(n12848), .B(n12846), .Z(n12847) );
  XOR U11532 ( .A(n12849), .B(n12850), .Z(n11522) );
  NOR U11533 ( .A(n12851), .B(n12849), .Z(n12850) );
  XOR U11534 ( .A(n12852), .B(n12853), .Z(n11525) );
  NOR U11535 ( .A(n12854), .B(n12852), .Z(n12853) );
  XOR U11536 ( .A(n12855), .B(n12856), .Z(n11528) );
  NOR U11537 ( .A(n12857), .B(n12855), .Z(n12856) );
  XOR U11538 ( .A(n12858), .B(n12859), .Z(n11531) );
  NOR U11539 ( .A(n12860), .B(n12858), .Z(n12859) );
  XOR U11540 ( .A(n12861), .B(n12862), .Z(n11534) );
  NOR U11541 ( .A(n12863), .B(n12861), .Z(n12862) );
  XOR U11542 ( .A(n12864), .B(n12865), .Z(n11537) );
  NOR U11543 ( .A(n12866), .B(n12864), .Z(n12865) );
  XOR U11544 ( .A(n12867), .B(n12868), .Z(n11540) );
  NOR U11545 ( .A(n12869), .B(n12867), .Z(n12868) );
  XOR U11546 ( .A(n12870), .B(n12871), .Z(n11543) );
  NOR U11547 ( .A(n12872), .B(n12870), .Z(n12871) );
  XOR U11548 ( .A(n12873), .B(n12874), .Z(n11546) );
  NOR U11549 ( .A(n12875), .B(n12873), .Z(n12874) );
  XOR U11550 ( .A(n12876), .B(n12877), .Z(n11549) );
  NOR U11551 ( .A(n12878), .B(n12876), .Z(n12877) );
  XOR U11552 ( .A(n12879), .B(n12880), .Z(n11552) );
  NOR U11553 ( .A(n12881), .B(n12879), .Z(n12880) );
  XOR U11554 ( .A(n12882), .B(n12883), .Z(n11555) );
  NOR U11555 ( .A(n12884), .B(n12882), .Z(n12883) );
  XOR U11556 ( .A(n12885), .B(n12886), .Z(n11558) );
  NOR U11557 ( .A(n12887), .B(n12885), .Z(n12886) );
  XOR U11558 ( .A(n12888), .B(n12889), .Z(n11561) );
  NOR U11559 ( .A(n12890), .B(n12888), .Z(n12889) );
  XOR U11560 ( .A(n12891), .B(n12892), .Z(n11564) );
  NOR U11561 ( .A(n12893), .B(n12891), .Z(n12892) );
  XOR U11562 ( .A(n12894), .B(n12895), .Z(n11567) );
  NOR U11563 ( .A(n12896), .B(n12894), .Z(n12895) );
  XOR U11564 ( .A(n12897), .B(n12898), .Z(n11570) );
  NOR U11565 ( .A(n12899), .B(n12897), .Z(n12898) );
  XOR U11566 ( .A(n12900), .B(n12901), .Z(n11573) );
  AND U11567 ( .A(n12902), .B(n12900), .Z(n12901) );
  XOR U11568 ( .A(n12903), .B(n12904), .Z(n11576) );
  AND U11569 ( .A(n78), .B(n12903), .Z(n12904) );
  XOR U11570 ( .A(n60), .B(n12255), .Z(n12257) );
  XOR U11571 ( .A(n12252), .B(n12251), .Z(n60) );
  XNOR U11572 ( .A(n12249), .B(n12248), .Z(n12251) );
  XNOR U11573 ( .A(n12246), .B(n12245), .Z(n12248) );
  XNOR U11574 ( .A(n12243), .B(n12242), .Z(n12245) );
  XNOR U11575 ( .A(n12240), .B(n12239), .Z(n12242) );
  XNOR U11576 ( .A(n12237), .B(n12236), .Z(n12239) );
  XNOR U11577 ( .A(n12234), .B(n12233), .Z(n12236) );
  XNOR U11578 ( .A(n12231), .B(n12230), .Z(n12233) );
  XNOR U11579 ( .A(n12228), .B(n12227), .Z(n12230) );
  XNOR U11580 ( .A(n12225), .B(n12224), .Z(n12227) );
  XNOR U11581 ( .A(n12222), .B(n12221), .Z(n12224) );
  XNOR U11582 ( .A(n12219), .B(n12218), .Z(n12221) );
  XNOR U11583 ( .A(n12216), .B(n12215), .Z(n12218) );
  XNOR U11584 ( .A(n12213), .B(n12212), .Z(n12215) );
  XNOR U11585 ( .A(n12210), .B(n12209), .Z(n12212) );
  XNOR U11586 ( .A(n12207), .B(n12206), .Z(n12209) );
  XNOR U11587 ( .A(n12204), .B(n12203), .Z(n12206) );
  XNOR U11588 ( .A(n12201), .B(n12200), .Z(n12203) );
  XNOR U11589 ( .A(n12198), .B(n12197), .Z(n12200) );
  XNOR U11590 ( .A(n12195), .B(n12194), .Z(n12197) );
  XNOR U11591 ( .A(n12192), .B(n12191), .Z(n12194) );
  XNOR U11592 ( .A(n12189), .B(n12188), .Z(n12191) );
  XNOR U11593 ( .A(n12186), .B(n12185), .Z(n12188) );
  XNOR U11594 ( .A(n12183), .B(n12182), .Z(n12185) );
  XNOR U11595 ( .A(n12180), .B(n12179), .Z(n12182) );
  XNOR U11596 ( .A(n12177), .B(n12176), .Z(n12179) );
  XNOR U11597 ( .A(n12174), .B(n12173), .Z(n12176) );
  XNOR U11598 ( .A(n12171), .B(n12170), .Z(n12173) );
  XNOR U11599 ( .A(n12168), .B(n12167), .Z(n12170) );
  XNOR U11600 ( .A(n12165), .B(n12164), .Z(n12167) );
  XNOR U11601 ( .A(n12162), .B(n12161), .Z(n12164) );
  XNOR U11602 ( .A(n12159), .B(n12158), .Z(n12161) );
  XNOR U11603 ( .A(n12156), .B(n12155), .Z(n12158) );
  XNOR U11604 ( .A(n12153), .B(n12152), .Z(n12155) );
  XNOR U11605 ( .A(n12150), .B(n12149), .Z(n12152) );
  XNOR U11606 ( .A(n12147), .B(n12146), .Z(n12149) );
  XNOR U11607 ( .A(n12144), .B(n12143), .Z(n12146) );
  XNOR U11608 ( .A(n12141), .B(n12140), .Z(n12143) );
  XNOR U11609 ( .A(n12138), .B(n12137), .Z(n12140) );
  XNOR U11610 ( .A(n12135), .B(n12134), .Z(n12137) );
  XNOR U11611 ( .A(n12132), .B(n12131), .Z(n12134) );
  XNOR U11612 ( .A(n12129), .B(n12128), .Z(n12131) );
  XNOR U11613 ( .A(n12126), .B(n12125), .Z(n12128) );
  XNOR U11614 ( .A(n12123), .B(n12122), .Z(n12125) );
  XNOR U11615 ( .A(n12120), .B(n12119), .Z(n12122) );
  XNOR U11616 ( .A(n12117), .B(n12116), .Z(n12119) );
  XNOR U11617 ( .A(n12114), .B(n12113), .Z(n12116) );
  XNOR U11618 ( .A(n12111), .B(n12110), .Z(n12113) );
  XNOR U11619 ( .A(n12108), .B(n12107), .Z(n12110) );
  XNOR U11620 ( .A(n12105), .B(n12104), .Z(n12107) );
  XNOR U11621 ( .A(n12102), .B(n12101), .Z(n12104) );
  XNOR U11622 ( .A(n12099), .B(n12098), .Z(n12101) );
  XNOR U11623 ( .A(n12096), .B(n12095), .Z(n12098) );
  XNOR U11624 ( .A(n12093), .B(n12092), .Z(n12095) );
  XNOR U11625 ( .A(n12090), .B(n12089), .Z(n12092) );
  XNOR U11626 ( .A(n12087), .B(n12086), .Z(n12089) );
  XNOR U11627 ( .A(n12084), .B(n12083), .Z(n12086) );
  XNOR U11628 ( .A(n12081), .B(n12080), .Z(n12083) );
  XNOR U11629 ( .A(n12078), .B(n12077), .Z(n12080) );
  XNOR U11630 ( .A(n12075), .B(n12074), .Z(n12077) );
  XNOR U11631 ( .A(n12072), .B(n12071), .Z(n12074) );
  XNOR U11632 ( .A(n12069), .B(n12068), .Z(n12071) );
  XNOR U11633 ( .A(n12066), .B(n12065), .Z(n12068) );
  XNOR U11634 ( .A(n12063), .B(n12062), .Z(n12065) );
  XNOR U11635 ( .A(n12060), .B(n12059), .Z(n12062) );
  XNOR U11636 ( .A(n12057), .B(n12056), .Z(n12059) );
  XNOR U11637 ( .A(n12054), .B(n12053), .Z(n12056) );
  XNOR U11638 ( .A(n12051), .B(n12050), .Z(n12053) );
  XNOR U11639 ( .A(n12048), .B(n12047), .Z(n12050) );
  XNOR U11640 ( .A(n12045), .B(n12044), .Z(n12047) );
  XNOR U11641 ( .A(n12042), .B(n12041), .Z(n12044) );
  XNOR U11642 ( .A(n12039), .B(n12038), .Z(n12041) );
  XNOR U11643 ( .A(n12036), .B(n12035), .Z(n12038) );
  XNOR U11644 ( .A(n12033), .B(n12032), .Z(n12035) );
  XNOR U11645 ( .A(n12030), .B(n12029), .Z(n12032) );
  XNOR U11646 ( .A(n12027), .B(n12026), .Z(n12029) );
  XNOR U11647 ( .A(n12024), .B(n12023), .Z(n12026) );
  XNOR U11648 ( .A(n12021), .B(n12020), .Z(n12023) );
  XNOR U11649 ( .A(n12018), .B(n12017), .Z(n12020) );
  XNOR U11650 ( .A(n12015), .B(n12014), .Z(n12017) );
  XNOR U11651 ( .A(n12012), .B(n12011), .Z(n12014) );
  XNOR U11652 ( .A(n12009), .B(n12008), .Z(n12011) );
  XNOR U11653 ( .A(n12006), .B(n12005), .Z(n12008) );
  XNOR U11654 ( .A(n12003), .B(n12002), .Z(n12005) );
  XNOR U11655 ( .A(n12000), .B(n11999), .Z(n12002) );
  XNOR U11656 ( .A(n11997), .B(n11996), .Z(n11999) );
  XNOR U11657 ( .A(n11994), .B(n11993), .Z(n11996) );
  XNOR U11658 ( .A(n11991), .B(n11990), .Z(n11993) );
  XNOR U11659 ( .A(n11988), .B(n11987), .Z(n11990) );
  XNOR U11660 ( .A(n11985), .B(n11984), .Z(n11987) );
  XNOR U11661 ( .A(n11982), .B(n11981), .Z(n11984) );
  XNOR U11662 ( .A(n11979), .B(n11978), .Z(n11981) );
  XNOR U11663 ( .A(n11976), .B(n11975), .Z(n11978) );
  XNOR U11664 ( .A(n11973), .B(n11972), .Z(n11975) );
  XNOR U11665 ( .A(n11970), .B(n11969), .Z(n11972) );
  XNOR U11666 ( .A(n11967), .B(n11966), .Z(n11969) );
  XNOR U11667 ( .A(n11964), .B(n11963), .Z(n11966) );
  XNOR U11668 ( .A(n11961), .B(n11960), .Z(n11963) );
  XNOR U11669 ( .A(n11958), .B(n11957), .Z(n11960) );
  XNOR U11670 ( .A(n11955), .B(n11954), .Z(n11957) );
  XNOR U11671 ( .A(n11952), .B(n11951), .Z(n11954) );
  XNOR U11672 ( .A(n11949), .B(n11948), .Z(n11951) );
  XNOR U11673 ( .A(n11946), .B(n11945), .Z(n11948) );
  XNOR U11674 ( .A(n11943), .B(n11942), .Z(n11945) );
  XNOR U11675 ( .A(n11940), .B(n11939), .Z(n11942) );
  XNOR U11676 ( .A(n11937), .B(n11936), .Z(n11939) );
  XNOR U11677 ( .A(n11934), .B(n11933), .Z(n11936) );
  XNOR U11678 ( .A(n11931), .B(n11930), .Z(n11933) );
  XNOR U11679 ( .A(n11928), .B(n11927), .Z(n11930) );
  XNOR U11680 ( .A(n11925), .B(n11924), .Z(n11927) );
  XNOR U11681 ( .A(n11922), .B(n11921), .Z(n11924) );
  XNOR U11682 ( .A(n11919), .B(n11918), .Z(n11921) );
  XNOR U11683 ( .A(n11916), .B(n11915), .Z(n11918) );
  XNOR U11684 ( .A(n11913), .B(n11912), .Z(n11915) );
  XNOR U11685 ( .A(n11910), .B(n11909), .Z(n11912) );
  XNOR U11686 ( .A(n11907), .B(n11906), .Z(n11909) );
  XNOR U11687 ( .A(n11904), .B(n11903), .Z(n11906) );
  XNOR U11688 ( .A(n11901), .B(n11900), .Z(n11903) );
  XNOR U11689 ( .A(n11898), .B(n11897), .Z(n11900) );
  XNOR U11690 ( .A(n11895), .B(n11894), .Z(n11897) );
  XNOR U11691 ( .A(n11892), .B(n11891), .Z(n11894) );
  XNOR U11692 ( .A(n11889), .B(n11888), .Z(n11891) );
  XNOR U11693 ( .A(n11886), .B(n11885), .Z(n11888) );
  XNOR U11694 ( .A(n11883), .B(n11882), .Z(n11885) );
  XNOR U11695 ( .A(n11880), .B(n11879), .Z(n11882) );
  XNOR U11696 ( .A(n11877), .B(n11876), .Z(n11879) );
  XNOR U11697 ( .A(n11874), .B(n11873), .Z(n11876) );
  XNOR U11698 ( .A(n11871), .B(n11870), .Z(n11873) );
  XOR U11699 ( .A(n11868), .B(n11603), .Z(n11870) );
  XOR U11700 ( .A(n12905), .B(n11591), .Z(n11603) );
  XNOR U11701 ( .A(n11592), .B(n11589), .Z(n11591) );
  XNOR U11702 ( .A(n11590), .B(n11586), .Z(n11589) );
  XNOR U11703 ( .A(n11585), .B(n11612), .Z(n11586) );
  XNOR U11704 ( .A(n11611), .B(n11867), .Z(n11612) );
  XNOR U11705 ( .A(n11858), .B(n11866), .Z(n11867) );
  XNOR U11706 ( .A(n11857), .B(n11863), .Z(n11866) );
  XNOR U11707 ( .A(n11862), .B(n11621), .Z(n11863) );
  XNOR U11708 ( .A(n11620), .B(n11856), .Z(n11621) );
  XNOR U11709 ( .A(n11847), .B(n11855), .Z(n11856) );
  XOR U11710 ( .A(n11846), .B(n11852), .Z(n11855) );
  XOR U11711 ( .A(n11851), .B(n11833), .Z(n11852) );
  XOR U11712 ( .A(n11627), .B(n11844), .Z(n11833) );
  XOR U11713 ( .A(n11845), .B(n11843), .Z(n11844) );
  XOR U11714 ( .A(n11834), .B(n11840), .Z(n11843) );
  XOR U11715 ( .A(n11638), .B(n11839), .Z(n11840) );
  AND U11716 ( .A(n12906), .B(n12907), .Z(n11839) );
  XOR U11717 ( .A(n11832), .B(n11637), .Z(n11638) );
  AND U11718 ( .A(n12908), .B(n12909), .Z(n11637) );
  XOR U11719 ( .A(n11829), .B(n11629), .Z(n11832) );
  AND U11720 ( .A(n12910), .B(n12911), .Z(n11629) );
  XNOR U11721 ( .A(n11827), .B(n11628), .Z(n11829) );
  AND U11722 ( .A(n12912), .B(n12913), .Z(n11628) );
  XOR U11723 ( .A(n11791), .B(n11828), .Z(n11827) );
  AND U11724 ( .A(n12914), .B(n12915), .Z(n11828) );
  XNOR U11725 ( .A(n11822), .B(n11792), .Z(n11791) );
  AND U11726 ( .A(n12916), .B(n12917), .Z(n11792) );
  XOR U11727 ( .A(n11821), .B(n11813), .Z(n11822) );
  AND U11728 ( .A(n12918), .B(n12919), .Z(n11813) );
  XNOR U11729 ( .A(n11816), .B(n11812), .Z(n11821) );
  AND U11730 ( .A(n12920), .B(n12921), .Z(n11812) );
  XOR U11731 ( .A(n11793), .B(n11817), .Z(n11816) );
  AND U11732 ( .A(n12922), .B(n12923), .Z(n11817) );
  XNOR U11733 ( .A(n11809), .B(n11794), .Z(n11793) );
  AND U11734 ( .A(n12924), .B(n12925), .Z(n11794) );
  XOR U11735 ( .A(n11808), .B(n11800), .Z(n11809) );
  AND U11736 ( .A(n12926), .B(n12927), .Z(n11800) );
  XNOR U11737 ( .A(n11803), .B(n11799), .Z(n11808) );
  AND U11738 ( .A(n12928), .B(n12929), .Z(n11799) );
  XOR U11739 ( .A(n11746), .B(n11804), .Z(n11803) );
  AND U11740 ( .A(n12930), .B(n12931), .Z(n11804) );
  XNOR U11741 ( .A(n11788), .B(n11747), .Z(n11746) );
  AND U11742 ( .A(n12932), .B(n12933), .Z(n11747) );
  XOR U11743 ( .A(n11787), .B(n11779), .Z(n11788) );
  AND U11744 ( .A(n12934), .B(n12935), .Z(n11779) );
  XNOR U11745 ( .A(n11782), .B(n11778), .Z(n11787) );
  AND U11746 ( .A(n12936), .B(n12937), .Z(n11778) );
  XOR U11747 ( .A(n11750), .B(n11783), .Z(n11782) );
  AND U11748 ( .A(n12938), .B(n12939), .Z(n11783) );
  XNOR U11749 ( .A(n11775), .B(n11751), .Z(n11750) );
  AND U11750 ( .A(n12940), .B(n12941), .Z(n11751) );
  XOR U11751 ( .A(n11774), .B(n11766), .Z(n11775) );
  AND U11752 ( .A(n12942), .B(n12943), .Z(n11766) );
  XNOR U11753 ( .A(n11769), .B(n11765), .Z(n11774) );
  AND U11754 ( .A(n12944), .B(n12945), .Z(n11765) );
  XOR U11755 ( .A(n11710), .B(n11770), .Z(n11769) );
  AND U11756 ( .A(n12946), .B(n12947), .Z(n11770) );
  XNOR U11757 ( .A(n11760), .B(n11711), .Z(n11710) );
  AND U11758 ( .A(n12948), .B(n12949), .Z(n11711) );
  XOR U11759 ( .A(n11759), .B(n11745), .Z(n11760) );
  AND U11760 ( .A(n12950), .B(n12951), .Z(n11745) );
  XNOR U11761 ( .A(n11754), .B(n11744), .Z(n11759) );
  AND U11762 ( .A(n12952), .B(n12953), .Z(n11744) );
  XOR U11763 ( .A(n11714), .B(n11755), .Z(n11754) );
  AND U11764 ( .A(n12954), .B(n12955), .Z(n11755) );
  XNOR U11765 ( .A(n11743), .B(n11715), .Z(n11714) );
  AND U11766 ( .A(n12956), .B(n12957), .Z(n11715) );
  XOR U11767 ( .A(n11742), .B(n11732), .Z(n11743) );
  AND U11768 ( .A(n12958), .B(n12959), .Z(n11732) );
  XNOR U11769 ( .A(n11737), .B(n11731), .Z(n11742) );
  AND U11770 ( .A(n12960), .B(n12961), .Z(n11731) );
  XOR U11771 ( .A(n11657), .B(n11738), .Z(n11737) );
  AND U11772 ( .A(n12962), .B(n12963), .Z(n11738) );
  XNOR U11773 ( .A(n11730), .B(n11658), .Z(n11657) );
  AND U11774 ( .A(n12964), .B(n12965), .Z(n11658) );
  XOR U11775 ( .A(n11729), .B(n11717), .Z(n11730) );
  AND U11776 ( .A(n12966), .B(n12967), .Z(n11717) );
  XNOR U11777 ( .A(n11724), .B(n11716), .Z(n11729) );
  AND U11778 ( .A(n12968), .B(n12969), .Z(n11716) );
  XOR U11779 ( .A(n11659), .B(n11725), .Z(n11724) );
  AND U11780 ( .A(n12970), .B(n12971), .Z(n11725) );
  XNOR U11781 ( .A(n11709), .B(n11660), .Z(n11659) );
  AND U11782 ( .A(n12972), .B(n12973), .Z(n11660) );
  XOR U11783 ( .A(n11708), .B(n11700), .Z(n11709) );
  AND U11784 ( .A(n12974), .B(n12975), .Z(n11700) );
  XNOR U11785 ( .A(n11703), .B(n11699), .Z(n11708) );
  AND U11786 ( .A(n12976), .B(n12977), .Z(n11699) );
  XOR U11787 ( .A(n11663), .B(n11704), .Z(n11703) );
  AND U11788 ( .A(n12978), .B(n12979), .Z(n11704) );
  XNOR U11789 ( .A(n11696), .B(n11664), .Z(n11663) );
  AND U11790 ( .A(n12980), .B(n12981), .Z(n11664) );
  XOR U11791 ( .A(n11695), .B(n11687), .Z(n11696) );
  AND U11792 ( .A(n12982), .B(n12983), .Z(n11687) );
  XNOR U11793 ( .A(n11690), .B(n11686), .Z(n11695) );
  AND U11794 ( .A(n12984), .B(n12985), .Z(n11686) );
  XOR U11795 ( .A(n12986), .B(n12987), .Z(n11690) );
  XOR U11796 ( .A(n12988), .B(n12989), .Z(n12987) );
  XOR U11797 ( .A(n12990), .B(n12991), .Z(n12989) );
  XNOR U11798 ( .A(n11680), .B(n11673), .Z(n12991) );
  XOR U11799 ( .A(n12992), .B(n12993), .Z(n11673) );
  XOR U11800 ( .A(n12994), .B(n12995), .Z(n12993) );
  XOR U11801 ( .A(n12996), .B(n12997), .Z(n12995) );
  NOR U11802 ( .A(n12998), .B(n12999), .Z(n12997) );
  NOR U11803 ( .A(n13000), .B(n13001), .Z(n12996) );
  AND U11804 ( .A(n13002), .B(n13003), .Z(n13001) );
  IV U11805 ( .A(n13004), .Z(n13000) );
  NOR U11806 ( .A(n13005), .B(n13006), .Z(n13004) );
  AND U11807 ( .A(n12998), .B(n13007), .Z(n13006) );
  AND U11808 ( .A(n12999), .B(n13008), .Z(n13005) );
  NOR U11809 ( .A(n13009), .B(n13010), .Z(n12994) );
  AND U11810 ( .A(n13011), .B(n13012), .Z(n13010) );
  IV U11811 ( .A(n13013), .Z(n13009) );
  NOR U11812 ( .A(n13014), .B(n13015), .Z(n13013) );
  AND U11813 ( .A(n13016), .B(n13017), .Z(n13015) );
  AND U11814 ( .A(n13018), .B(n13019), .Z(n13014) );
  XOR U11815 ( .A(n13020), .B(n13021), .Z(n12992) );
  XOR U11816 ( .A(n13022), .B(n13023), .Z(n13021) );
  XOR U11817 ( .A(n13024), .B(n13025), .Z(n13023) );
  XOR U11818 ( .A(n13026), .B(n13027), .Z(n13025) );
  AND U11819 ( .A(n13028), .B(n13029), .Z(n13027) );
  AND U11820 ( .A(n13030), .B(n13031), .Z(n13026) );
  XOR U11821 ( .A(n13032), .B(n13033), .Z(n13024) );
  AND U11822 ( .A(n13034), .B(n13035), .Z(n13033) );
  AND U11823 ( .A(n13036), .B(n13037), .Z(n13032) );
  AND U11824 ( .A(n13038), .B(n13039), .Z(n13037) );
  AND U11825 ( .A(n13040), .B(n13041), .Z(n13039) );
  NOR U11826 ( .A(n13042), .B(n13043), .Z(n13041) );
  IV U11827 ( .A(n13044), .Z(n13042) );
  NOR U11828 ( .A(n13045), .B(n13046), .Z(n13044) );
  NOR U11829 ( .A(n13047), .B(n13048), .Z(n13040) );
  AND U11830 ( .A(n13049), .B(n13050), .Z(n13038) );
  NOR U11831 ( .A(n13051), .B(n13052), .Z(n13050) );
  NOR U11832 ( .A(n13053), .B(n13054), .Z(n13049) );
  AND U11833 ( .A(n13055), .B(n13056), .Z(n13036) );
  AND U11834 ( .A(n13057), .B(n13058), .Z(n13056) );
  NOR U11835 ( .A(n13059), .B(n13060), .Z(n13058) );
  NOR U11836 ( .A(n13061), .B(n13062), .Z(n13057) );
  AND U11837 ( .A(n13063), .B(n13064), .Z(n13055) );
  NOR U11838 ( .A(n13065), .B(n13066), .Z(n13064) );
  NOR U11839 ( .A(n13067), .B(n13068), .Z(n13063) );
  XOR U11840 ( .A(n13069), .B(n13070), .Z(n13022) );
  XOR U11841 ( .A(n13071), .B(n13072), .Z(n13070) );
  NOR U11842 ( .A(n13073), .B(n13074), .Z(n13072) );
  NOR U11843 ( .A(n13075), .B(n13076), .Z(n13071) );
  AND U11844 ( .A(n13077), .B(n13078), .Z(n13076) );
  IV U11845 ( .A(n13079), .Z(n13075) );
  NOR U11846 ( .A(n13080), .B(n13081), .Z(n13079) );
  AND U11847 ( .A(n13073), .B(n13082), .Z(n13081) );
  AND U11848 ( .A(n13074), .B(n13083), .Z(n13080) );
  XOR U11849 ( .A(n13084), .B(n13085), .Z(n13069) );
  NOR U11850 ( .A(n13086), .B(n13087), .Z(n13085) );
  NOR U11851 ( .A(n13088), .B(n13089), .Z(n13084) );
  AND U11852 ( .A(n13090), .B(n13091), .Z(n13089) );
  IV U11853 ( .A(n13092), .Z(n13088) );
  NOR U11854 ( .A(n13093), .B(n13094), .Z(n13092) );
  AND U11855 ( .A(n13086), .B(n13095), .Z(n13094) );
  AND U11856 ( .A(n13087), .B(n13096), .Z(n13093) );
  XNOR U11857 ( .A(n13097), .B(n13098), .Z(n13020) );
  AND U11858 ( .A(n13099), .B(n13100), .Z(n13098) );
  NOR U11859 ( .A(n13016), .B(n13018), .Z(n13097) );
  AND U11860 ( .A(n13101), .B(n13102), .Z(n11680) );
  XOR U11861 ( .A(n11678), .B(n11679), .Z(n12990) );
  AND U11862 ( .A(n13103), .B(n13104), .Z(n11679) );
  AND U11863 ( .A(n13105), .B(n13106), .Z(n11678) );
  XOR U11864 ( .A(n13107), .B(n13108), .Z(n12988) );
  XOR U11865 ( .A(n11674), .B(n11675), .Z(n13108) );
  AND U11866 ( .A(n13109), .B(n13110), .Z(n11675) );
  AND U11867 ( .A(n13111), .B(n13112), .Z(n11674) );
  XOR U11868 ( .A(n11672), .B(n11670), .Z(n13107) );
  AND U11869 ( .A(n13113), .B(n13114), .Z(n11670) );
  AND U11870 ( .A(n13115), .B(n13116), .Z(n11672) );
  XNOR U11871 ( .A(n11681), .B(n11691), .Z(n12986) );
  AND U11872 ( .A(n13117), .B(n13118), .Z(n11691) );
  AND U11873 ( .A(n13119), .B(n13120), .Z(n11681) );
  XOR U11874 ( .A(n13121), .B(n13122), .Z(n11834) );
  AND U11875 ( .A(n13121), .B(n13123), .Z(n13122) );
  IV U11876 ( .A(n11835), .Z(n11845) );
  XNOR U11877 ( .A(n13124), .B(n13125), .Z(n11835) );
  AND U11878 ( .A(n13124), .B(n13126), .Z(n13125) );
  XOR U11879 ( .A(n13127), .B(n13128), .Z(n11627) );
  AND U11880 ( .A(n13127), .B(n13129), .Z(n13128) );
  XOR U11881 ( .A(n13130), .B(n13131), .Z(n11851) );
  AND U11882 ( .A(n13130), .B(n13132), .Z(n13131) );
  XNOR U11883 ( .A(n13133), .B(n13134), .Z(n11846) );
  AND U11884 ( .A(n13133), .B(n13135), .Z(n13134) );
  XNOR U11885 ( .A(n13136), .B(n13137), .Z(n11847) );
  AND U11886 ( .A(n13138), .B(n13136), .Z(n13137) );
  XOR U11887 ( .A(n13139), .B(n13140), .Z(n11620) );
  NOR U11888 ( .A(n13141), .B(n13139), .Z(n13140) );
  XOR U11889 ( .A(n13142), .B(n13143), .Z(n11862) );
  NOR U11890 ( .A(n13144), .B(n13142), .Z(n13143) );
  XOR U11891 ( .A(n13145), .B(n13146), .Z(n11857) );
  NOR U11892 ( .A(n13147), .B(n13145), .Z(n13146) );
  XOR U11893 ( .A(n13148), .B(n13149), .Z(n11858) );
  NOR U11894 ( .A(n13150), .B(n13148), .Z(n13149) );
  XOR U11895 ( .A(n13151), .B(n13152), .Z(n11611) );
  NOR U11896 ( .A(n13153), .B(n13151), .Z(n13152) );
  XOR U11897 ( .A(n13154), .B(n13155), .Z(n11585) );
  NOR U11898 ( .A(n13156), .B(n13154), .Z(n13155) );
  XOR U11899 ( .A(n13157), .B(n13158), .Z(n11590) );
  NOR U11900 ( .A(n13159), .B(n13157), .Z(n13158) );
  XOR U11901 ( .A(n13160), .B(n13161), .Z(n11592) );
  NOR U11902 ( .A(n13162), .B(n13160), .Z(n13161) );
  IV U11903 ( .A(n11602), .Z(n12905) );
  XNOR U11904 ( .A(n13163), .B(n13164), .Z(n11602) );
  NOR U11905 ( .A(n13165), .B(n13163), .Z(n13164) );
  XOR U11906 ( .A(n13166), .B(n13167), .Z(n11868) );
  NOR U11907 ( .A(n13168), .B(n13166), .Z(n13167) );
  XOR U11908 ( .A(n13169), .B(n13170), .Z(n11871) );
  NOR U11909 ( .A(n13171), .B(n13169), .Z(n13170) );
  XOR U11910 ( .A(n13172), .B(n13173), .Z(n11874) );
  NOR U11911 ( .A(n13174), .B(n13172), .Z(n13173) );
  XOR U11912 ( .A(n13175), .B(n13176), .Z(n11877) );
  NOR U11913 ( .A(n13177), .B(n13175), .Z(n13176) );
  XOR U11914 ( .A(n13178), .B(n13179), .Z(n11880) );
  NOR U11915 ( .A(n13180), .B(n13178), .Z(n13179) );
  XOR U11916 ( .A(n13181), .B(n13182), .Z(n11883) );
  NOR U11917 ( .A(n13183), .B(n13181), .Z(n13182) );
  XOR U11918 ( .A(n13184), .B(n13185), .Z(n11886) );
  NOR U11919 ( .A(n13186), .B(n13184), .Z(n13185) );
  XOR U11920 ( .A(n13187), .B(n13188), .Z(n11889) );
  NOR U11921 ( .A(n13189), .B(n13187), .Z(n13188) );
  XOR U11922 ( .A(n13190), .B(n13191), .Z(n11892) );
  NOR U11923 ( .A(n13192), .B(n13190), .Z(n13191) );
  XOR U11924 ( .A(n13193), .B(n13194), .Z(n11895) );
  NOR U11925 ( .A(n13195), .B(n13193), .Z(n13194) );
  XOR U11926 ( .A(n13196), .B(n13197), .Z(n11898) );
  NOR U11927 ( .A(n13198), .B(n13196), .Z(n13197) );
  XOR U11928 ( .A(n13199), .B(n13200), .Z(n11901) );
  NOR U11929 ( .A(n13201), .B(n13199), .Z(n13200) );
  XOR U11930 ( .A(n13202), .B(n13203), .Z(n11904) );
  NOR U11931 ( .A(n13204), .B(n13202), .Z(n13203) );
  XOR U11932 ( .A(n13205), .B(n13206), .Z(n11907) );
  NOR U11933 ( .A(n13207), .B(n13205), .Z(n13206) );
  XOR U11934 ( .A(n13208), .B(n13209), .Z(n11910) );
  NOR U11935 ( .A(n13210), .B(n13208), .Z(n13209) );
  XOR U11936 ( .A(n13211), .B(n13212), .Z(n11913) );
  NOR U11937 ( .A(n13213), .B(n13211), .Z(n13212) );
  XOR U11938 ( .A(n13214), .B(n13215), .Z(n11916) );
  NOR U11939 ( .A(n13216), .B(n13214), .Z(n13215) );
  XOR U11940 ( .A(n13217), .B(n13218), .Z(n11919) );
  NOR U11941 ( .A(n13219), .B(n13217), .Z(n13218) );
  XOR U11942 ( .A(n13220), .B(n13221), .Z(n11922) );
  NOR U11943 ( .A(n13222), .B(n13220), .Z(n13221) );
  XOR U11944 ( .A(n13223), .B(n13224), .Z(n11925) );
  NOR U11945 ( .A(n13225), .B(n13223), .Z(n13224) );
  XOR U11946 ( .A(n13226), .B(n13227), .Z(n11928) );
  NOR U11947 ( .A(n13228), .B(n13226), .Z(n13227) );
  XOR U11948 ( .A(n13229), .B(n13230), .Z(n11931) );
  NOR U11949 ( .A(n13231), .B(n13229), .Z(n13230) );
  XOR U11950 ( .A(n13232), .B(n13233), .Z(n11934) );
  NOR U11951 ( .A(n13234), .B(n13232), .Z(n13233) );
  XOR U11952 ( .A(n13235), .B(n13236), .Z(n11937) );
  NOR U11953 ( .A(n13237), .B(n13235), .Z(n13236) );
  XOR U11954 ( .A(n13238), .B(n13239), .Z(n11940) );
  NOR U11955 ( .A(n13240), .B(n13238), .Z(n13239) );
  XOR U11956 ( .A(n13241), .B(n13242), .Z(n11943) );
  NOR U11957 ( .A(n13243), .B(n13241), .Z(n13242) );
  XOR U11958 ( .A(n13244), .B(n13245), .Z(n11946) );
  NOR U11959 ( .A(n13246), .B(n13244), .Z(n13245) );
  XOR U11960 ( .A(n13247), .B(n13248), .Z(n11949) );
  NOR U11961 ( .A(n13249), .B(n13247), .Z(n13248) );
  XOR U11962 ( .A(n13250), .B(n13251), .Z(n11952) );
  NOR U11963 ( .A(n13252), .B(n13250), .Z(n13251) );
  XOR U11964 ( .A(n13253), .B(n13254), .Z(n11955) );
  NOR U11965 ( .A(n13255), .B(n13253), .Z(n13254) );
  XOR U11966 ( .A(n13256), .B(n13257), .Z(n11958) );
  NOR U11967 ( .A(n13258), .B(n13256), .Z(n13257) );
  XOR U11968 ( .A(n13259), .B(n13260), .Z(n11961) );
  NOR U11969 ( .A(n13261), .B(n13259), .Z(n13260) );
  XOR U11970 ( .A(n13262), .B(n13263), .Z(n11964) );
  NOR U11971 ( .A(n13264), .B(n13262), .Z(n13263) );
  XOR U11972 ( .A(n13265), .B(n13266), .Z(n11967) );
  NOR U11973 ( .A(n13267), .B(n13265), .Z(n13266) );
  XOR U11974 ( .A(n13268), .B(n13269), .Z(n11970) );
  NOR U11975 ( .A(n13270), .B(n13268), .Z(n13269) );
  XOR U11976 ( .A(n13271), .B(n13272), .Z(n11973) );
  NOR U11977 ( .A(n13273), .B(n13271), .Z(n13272) );
  XOR U11978 ( .A(n13274), .B(n13275), .Z(n11976) );
  NOR U11979 ( .A(n13276), .B(n13274), .Z(n13275) );
  XOR U11980 ( .A(n13277), .B(n13278), .Z(n11979) );
  NOR U11981 ( .A(n13279), .B(n13277), .Z(n13278) );
  XOR U11982 ( .A(n13280), .B(n13281), .Z(n11982) );
  NOR U11983 ( .A(n13282), .B(n13280), .Z(n13281) );
  XOR U11984 ( .A(n13283), .B(n13284), .Z(n11985) );
  NOR U11985 ( .A(n13285), .B(n13283), .Z(n13284) );
  XOR U11986 ( .A(n13286), .B(n13287), .Z(n11988) );
  NOR U11987 ( .A(n13288), .B(n13286), .Z(n13287) );
  XOR U11988 ( .A(n13289), .B(n13290), .Z(n11991) );
  NOR U11989 ( .A(n13291), .B(n13289), .Z(n13290) );
  XOR U11990 ( .A(n13292), .B(n13293), .Z(n11994) );
  NOR U11991 ( .A(n13294), .B(n13292), .Z(n13293) );
  XOR U11992 ( .A(n13295), .B(n13296), .Z(n11997) );
  NOR U11993 ( .A(n13297), .B(n13295), .Z(n13296) );
  XOR U11994 ( .A(n13298), .B(n13299), .Z(n12000) );
  NOR U11995 ( .A(n13300), .B(n13298), .Z(n13299) );
  XOR U11996 ( .A(n13301), .B(n13302), .Z(n12003) );
  NOR U11997 ( .A(n13303), .B(n13301), .Z(n13302) );
  XOR U11998 ( .A(n13304), .B(n13305), .Z(n12006) );
  NOR U11999 ( .A(n13306), .B(n13304), .Z(n13305) );
  XOR U12000 ( .A(n13307), .B(n13308), .Z(n12009) );
  NOR U12001 ( .A(n13309), .B(n13307), .Z(n13308) );
  XOR U12002 ( .A(n13310), .B(n13311), .Z(n12012) );
  NOR U12003 ( .A(n13312), .B(n13310), .Z(n13311) );
  XOR U12004 ( .A(n13313), .B(n13314), .Z(n12015) );
  NOR U12005 ( .A(n13315), .B(n13313), .Z(n13314) );
  XOR U12006 ( .A(n13316), .B(n13317), .Z(n12018) );
  NOR U12007 ( .A(n13318), .B(n13316), .Z(n13317) );
  XOR U12008 ( .A(n13319), .B(n13320), .Z(n12021) );
  NOR U12009 ( .A(n13321), .B(n13319), .Z(n13320) );
  XOR U12010 ( .A(n13322), .B(n13323), .Z(n12024) );
  NOR U12011 ( .A(n13324), .B(n13322), .Z(n13323) );
  XOR U12012 ( .A(n13325), .B(n13326), .Z(n12027) );
  NOR U12013 ( .A(n13327), .B(n13325), .Z(n13326) );
  XOR U12014 ( .A(n13328), .B(n13329), .Z(n12030) );
  NOR U12015 ( .A(n13330), .B(n13328), .Z(n13329) );
  XOR U12016 ( .A(n13331), .B(n13332), .Z(n12033) );
  NOR U12017 ( .A(n13333), .B(n13331), .Z(n13332) );
  XOR U12018 ( .A(n13334), .B(n13335), .Z(n12036) );
  NOR U12019 ( .A(n13336), .B(n13334), .Z(n13335) );
  XOR U12020 ( .A(n13337), .B(n13338), .Z(n12039) );
  NOR U12021 ( .A(n13339), .B(n13337), .Z(n13338) );
  XOR U12022 ( .A(n13340), .B(n13341), .Z(n12042) );
  NOR U12023 ( .A(n13342), .B(n13340), .Z(n13341) );
  XOR U12024 ( .A(n13343), .B(n13344), .Z(n12045) );
  NOR U12025 ( .A(n13345), .B(n13343), .Z(n13344) );
  XOR U12026 ( .A(n13346), .B(n13347), .Z(n12048) );
  NOR U12027 ( .A(n13348), .B(n13346), .Z(n13347) );
  XOR U12028 ( .A(n13349), .B(n13350), .Z(n12051) );
  NOR U12029 ( .A(n13351), .B(n13349), .Z(n13350) );
  XOR U12030 ( .A(n13352), .B(n13353), .Z(n12054) );
  NOR U12031 ( .A(n13354), .B(n13352), .Z(n13353) );
  XOR U12032 ( .A(n13355), .B(n13356), .Z(n12057) );
  NOR U12033 ( .A(n13357), .B(n13355), .Z(n13356) );
  XOR U12034 ( .A(n13358), .B(n13359), .Z(n12060) );
  NOR U12035 ( .A(n13360), .B(n13358), .Z(n13359) );
  XOR U12036 ( .A(n13361), .B(n13362), .Z(n12063) );
  NOR U12037 ( .A(n13363), .B(n13361), .Z(n13362) );
  XOR U12038 ( .A(n13364), .B(n13365), .Z(n12066) );
  NOR U12039 ( .A(n13366), .B(n13364), .Z(n13365) );
  XOR U12040 ( .A(n13367), .B(n13368), .Z(n12069) );
  NOR U12041 ( .A(n13369), .B(n13367), .Z(n13368) );
  XOR U12042 ( .A(n13370), .B(n13371), .Z(n12072) );
  NOR U12043 ( .A(n13372), .B(n13370), .Z(n13371) );
  XOR U12044 ( .A(n13373), .B(n13374), .Z(n12075) );
  NOR U12045 ( .A(n13375), .B(n13373), .Z(n13374) );
  XOR U12046 ( .A(n13376), .B(n13377), .Z(n12078) );
  NOR U12047 ( .A(n13378), .B(n13376), .Z(n13377) );
  XOR U12048 ( .A(n13379), .B(n13380), .Z(n12081) );
  NOR U12049 ( .A(n13381), .B(n13379), .Z(n13380) );
  XOR U12050 ( .A(n13382), .B(n13383), .Z(n12084) );
  NOR U12051 ( .A(n13384), .B(n13382), .Z(n13383) );
  XOR U12052 ( .A(n13385), .B(n13386), .Z(n12087) );
  NOR U12053 ( .A(n13387), .B(n13385), .Z(n13386) );
  XOR U12054 ( .A(n13388), .B(n13389), .Z(n12090) );
  NOR U12055 ( .A(n13390), .B(n13388), .Z(n13389) );
  XOR U12056 ( .A(n13391), .B(n13392), .Z(n12093) );
  NOR U12057 ( .A(n13393), .B(n13391), .Z(n13392) );
  XOR U12058 ( .A(n13394), .B(n13395), .Z(n12096) );
  NOR U12059 ( .A(n13396), .B(n13394), .Z(n13395) );
  XOR U12060 ( .A(n13397), .B(n13398), .Z(n12099) );
  NOR U12061 ( .A(n13399), .B(n13397), .Z(n13398) );
  XOR U12062 ( .A(n13400), .B(n13401), .Z(n12102) );
  NOR U12063 ( .A(n13402), .B(n13400), .Z(n13401) );
  XOR U12064 ( .A(n13403), .B(n13404), .Z(n12105) );
  NOR U12065 ( .A(n13405), .B(n13403), .Z(n13404) );
  XOR U12066 ( .A(n13406), .B(n13407), .Z(n12108) );
  NOR U12067 ( .A(n13408), .B(n13406), .Z(n13407) );
  XOR U12068 ( .A(n13409), .B(n13410), .Z(n12111) );
  NOR U12069 ( .A(n13411), .B(n13409), .Z(n13410) );
  XOR U12070 ( .A(n13412), .B(n13413), .Z(n12114) );
  NOR U12071 ( .A(n13414), .B(n13412), .Z(n13413) );
  XOR U12072 ( .A(n13415), .B(n13416), .Z(n12117) );
  NOR U12073 ( .A(n13417), .B(n13415), .Z(n13416) );
  XOR U12074 ( .A(n13418), .B(n13419), .Z(n12120) );
  NOR U12075 ( .A(n13420), .B(n13418), .Z(n13419) );
  XOR U12076 ( .A(n13421), .B(n13422), .Z(n12123) );
  NOR U12077 ( .A(n13423), .B(n13421), .Z(n13422) );
  XOR U12078 ( .A(n13424), .B(n13425), .Z(n12126) );
  NOR U12079 ( .A(n13426), .B(n13424), .Z(n13425) );
  XOR U12080 ( .A(n13427), .B(n13428), .Z(n12129) );
  NOR U12081 ( .A(n13429), .B(n13427), .Z(n13428) );
  XOR U12082 ( .A(n13430), .B(n13431), .Z(n12132) );
  NOR U12083 ( .A(n13432), .B(n13430), .Z(n13431) );
  XOR U12084 ( .A(n13433), .B(n13434), .Z(n12135) );
  NOR U12085 ( .A(n13435), .B(n13433), .Z(n13434) );
  XOR U12086 ( .A(n13436), .B(n13437), .Z(n12138) );
  NOR U12087 ( .A(n13438), .B(n13436), .Z(n13437) );
  XOR U12088 ( .A(n13439), .B(n13440), .Z(n12141) );
  NOR U12089 ( .A(n13441), .B(n13439), .Z(n13440) );
  XOR U12090 ( .A(n13442), .B(n13443), .Z(n12144) );
  NOR U12091 ( .A(n13444), .B(n13442), .Z(n13443) );
  XOR U12092 ( .A(n13445), .B(n13446), .Z(n12147) );
  NOR U12093 ( .A(n13447), .B(n13445), .Z(n13446) );
  XOR U12094 ( .A(n13448), .B(n13449), .Z(n12150) );
  NOR U12095 ( .A(n13450), .B(n13448), .Z(n13449) );
  XOR U12096 ( .A(n13451), .B(n13452), .Z(n12153) );
  NOR U12097 ( .A(n13453), .B(n13451), .Z(n13452) );
  XOR U12098 ( .A(n13454), .B(n13455), .Z(n12156) );
  NOR U12099 ( .A(n13456), .B(n13454), .Z(n13455) );
  XOR U12100 ( .A(n13457), .B(n13458), .Z(n12159) );
  NOR U12101 ( .A(n13459), .B(n13457), .Z(n13458) );
  XOR U12102 ( .A(n13460), .B(n13461), .Z(n12162) );
  NOR U12103 ( .A(n13462), .B(n13460), .Z(n13461) );
  XOR U12104 ( .A(n13463), .B(n13464), .Z(n12165) );
  NOR U12105 ( .A(n13465), .B(n13463), .Z(n13464) );
  XOR U12106 ( .A(n13466), .B(n13467), .Z(n12168) );
  NOR U12107 ( .A(n13468), .B(n13466), .Z(n13467) );
  XOR U12108 ( .A(n13469), .B(n13470), .Z(n12171) );
  NOR U12109 ( .A(n13471), .B(n13469), .Z(n13470) );
  XOR U12110 ( .A(n13472), .B(n13473), .Z(n12174) );
  NOR U12111 ( .A(n13474), .B(n13472), .Z(n13473) );
  XOR U12112 ( .A(n13475), .B(n13476), .Z(n12177) );
  NOR U12113 ( .A(n13477), .B(n13475), .Z(n13476) );
  XOR U12114 ( .A(n13478), .B(n13479), .Z(n12180) );
  NOR U12115 ( .A(n13480), .B(n13478), .Z(n13479) );
  XOR U12116 ( .A(n13481), .B(n13482), .Z(n12183) );
  NOR U12117 ( .A(n13483), .B(n13481), .Z(n13482) );
  XOR U12118 ( .A(n13484), .B(n13485), .Z(n12186) );
  NOR U12119 ( .A(n13486), .B(n13484), .Z(n13485) );
  XOR U12120 ( .A(n13487), .B(n13488), .Z(n12189) );
  NOR U12121 ( .A(n13489), .B(n13487), .Z(n13488) );
  XOR U12122 ( .A(n13490), .B(n13491), .Z(n12192) );
  NOR U12123 ( .A(n13492), .B(n13490), .Z(n13491) );
  XOR U12124 ( .A(n13493), .B(n13494), .Z(n12195) );
  NOR U12125 ( .A(n13495), .B(n13493), .Z(n13494) );
  XOR U12126 ( .A(n13496), .B(n13497), .Z(n12198) );
  NOR U12127 ( .A(n13498), .B(n13496), .Z(n13497) );
  XOR U12128 ( .A(n13499), .B(n13500), .Z(n12201) );
  NOR U12129 ( .A(n13501), .B(n13499), .Z(n13500) );
  XOR U12130 ( .A(n13502), .B(n13503), .Z(n12204) );
  NOR U12131 ( .A(n13504), .B(n13502), .Z(n13503) );
  XOR U12132 ( .A(n13505), .B(n13506), .Z(n12207) );
  NOR U12133 ( .A(n13507), .B(n13505), .Z(n13506) );
  XOR U12134 ( .A(n13508), .B(n13509), .Z(n12210) );
  NOR U12135 ( .A(n13510), .B(n13508), .Z(n13509) );
  XOR U12136 ( .A(n13511), .B(n13512), .Z(n12213) );
  NOR U12137 ( .A(n13513), .B(n13511), .Z(n13512) );
  XOR U12138 ( .A(n13514), .B(n13515), .Z(n12216) );
  NOR U12139 ( .A(n13516), .B(n13514), .Z(n13515) );
  XOR U12140 ( .A(n13517), .B(n13518), .Z(n12219) );
  NOR U12141 ( .A(n13519), .B(n13517), .Z(n13518) );
  XOR U12142 ( .A(n13520), .B(n13521), .Z(n12222) );
  NOR U12143 ( .A(n13522), .B(n13520), .Z(n13521) );
  XOR U12144 ( .A(n13523), .B(n13524), .Z(n12225) );
  NOR U12145 ( .A(n13525), .B(n13523), .Z(n13524) );
  XOR U12146 ( .A(n13526), .B(n13527), .Z(n12228) );
  NOR U12147 ( .A(n13528), .B(n13526), .Z(n13527) );
  XOR U12148 ( .A(n13529), .B(n13530), .Z(n12231) );
  NOR U12149 ( .A(n13531), .B(n13529), .Z(n13530) );
  XOR U12150 ( .A(n13532), .B(n13533), .Z(n12234) );
  NOR U12151 ( .A(n13534), .B(n13532), .Z(n13533) );
  XOR U12152 ( .A(n13535), .B(n13536), .Z(n12237) );
  NOR U12153 ( .A(n13537), .B(n13535), .Z(n13536) );
  XOR U12154 ( .A(n13538), .B(n13539), .Z(n12240) );
  NOR U12155 ( .A(n13540), .B(n13538), .Z(n13539) );
  XOR U12156 ( .A(n13541), .B(n13542), .Z(n12243) );
  NOR U12157 ( .A(n13543), .B(n13541), .Z(n13542) );
  XOR U12158 ( .A(n13544), .B(n13545), .Z(n12246) );
  NOR U12159 ( .A(n13546), .B(n13544), .Z(n13545) );
  XOR U12160 ( .A(n13547), .B(n13548), .Z(n12249) );
  NOR U12161 ( .A(n13549), .B(n13547), .Z(n13548) );
  XOR U12162 ( .A(n13550), .B(n13551), .Z(n12252) );
  NOR U12163 ( .A(n75), .B(n13552), .Z(n13551) );
  IV U12164 ( .A(n13550), .Z(n13552) );
  XOR U12165 ( .A(n13553), .B(n13554), .Z(n12255) );
  AND U12166 ( .A(n13555), .B(n13556), .Z(n13554) );
  XOR U12167 ( .A(n13553), .B(n78), .Z(n13556) );
  XOR U12168 ( .A(n12903), .B(n12902), .Z(n78) );
  XNOR U12169 ( .A(n12900), .B(n12899), .Z(n12902) );
  XNOR U12170 ( .A(n12897), .B(n12896), .Z(n12899) );
  XNOR U12171 ( .A(n12894), .B(n12893), .Z(n12896) );
  XNOR U12172 ( .A(n12891), .B(n12890), .Z(n12893) );
  XNOR U12173 ( .A(n12888), .B(n12887), .Z(n12890) );
  XNOR U12174 ( .A(n12885), .B(n12884), .Z(n12887) );
  XNOR U12175 ( .A(n12882), .B(n12881), .Z(n12884) );
  XNOR U12176 ( .A(n12879), .B(n12878), .Z(n12881) );
  XNOR U12177 ( .A(n12876), .B(n12875), .Z(n12878) );
  XNOR U12178 ( .A(n12873), .B(n12872), .Z(n12875) );
  XNOR U12179 ( .A(n12870), .B(n12869), .Z(n12872) );
  XNOR U12180 ( .A(n12867), .B(n12866), .Z(n12869) );
  XNOR U12181 ( .A(n12864), .B(n12863), .Z(n12866) );
  XNOR U12182 ( .A(n12861), .B(n12860), .Z(n12863) );
  XNOR U12183 ( .A(n12858), .B(n12857), .Z(n12860) );
  XNOR U12184 ( .A(n12855), .B(n12854), .Z(n12857) );
  XNOR U12185 ( .A(n12852), .B(n12851), .Z(n12854) );
  XNOR U12186 ( .A(n12849), .B(n12848), .Z(n12851) );
  XNOR U12187 ( .A(n12846), .B(n12845), .Z(n12848) );
  XNOR U12188 ( .A(n12843), .B(n12842), .Z(n12845) );
  XNOR U12189 ( .A(n12840), .B(n12839), .Z(n12842) );
  XNOR U12190 ( .A(n12837), .B(n12836), .Z(n12839) );
  XNOR U12191 ( .A(n12834), .B(n12833), .Z(n12836) );
  XNOR U12192 ( .A(n12831), .B(n12830), .Z(n12833) );
  XNOR U12193 ( .A(n12828), .B(n12827), .Z(n12830) );
  XNOR U12194 ( .A(n12825), .B(n12824), .Z(n12827) );
  XNOR U12195 ( .A(n12822), .B(n12821), .Z(n12824) );
  XNOR U12196 ( .A(n12819), .B(n12818), .Z(n12821) );
  XNOR U12197 ( .A(n12816), .B(n12815), .Z(n12818) );
  XNOR U12198 ( .A(n12813), .B(n12812), .Z(n12815) );
  XNOR U12199 ( .A(n12810), .B(n12809), .Z(n12812) );
  XNOR U12200 ( .A(n12807), .B(n12806), .Z(n12809) );
  XNOR U12201 ( .A(n12804), .B(n12803), .Z(n12806) );
  XNOR U12202 ( .A(n12801), .B(n12800), .Z(n12803) );
  XNOR U12203 ( .A(n12798), .B(n12797), .Z(n12800) );
  XNOR U12204 ( .A(n12795), .B(n12794), .Z(n12797) );
  XNOR U12205 ( .A(n12792), .B(n12791), .Z(n12794) );
  XNOR U12206 ( .A(n12789), .B(n12788), .Z(n12791) );
  XNOR U12207 ( .A(n12786), .B(n12785), .Z(n12788) );
  XNOR U12208 ( .A(n12783), .B(n12782), .Z(n12785) );
  XNOR U12209 ( .A(n12780), .B(n12779), .Z(n12782) );
  XNOR U12210 ( .A(n12777), .B(n12776), .Z(n12779) );
  XNOR U12211 ( .A(n12774), .B(n12773), .Z(n12776) );
  XNOR U12212 ( .A(n12771), .B(n12770), .Z(n12773) );
  XNOR U12213 ( .A(n12768), .B(n12767), .Z(n12770) );
  XNOR U12214 ( .A(n12765), .B(n12764), .Z(n12767) );
  XNOR U12215 ( .A(n12762), .B(n12761), .Z(n12764) );
  XNOR U12216 ( .A(n12759), .B(n12758), .Z(n12761) );
  XNOR U12217 ( .A(n12756), .B(n12755), .Z(n12758) );
  XNOR U12218 ( .A(n12753), .B(n12752), .Z(n12755) );
  XNOR U12219 ( .A(n12750), .B(n12749), .Z(n12752) );
  XNOR U12220 ( .A(n12747), .B(n12746), .Z(n12749) );
  XNOR U12221 ( .A(n12744), .B(n12743), .Z(n12746) );
  XNOR U12222 ( .A(n12741), .B(n12740), .Z(n12743) );
  XNOR U12223 ( .A(n12738), .B(n12737), .Z(n12740) );
  XNOR U12224 ( .A(n12735), .B(n12734), .Z(n12737) );
  XNOR U12225 ( .A(n12732), .B(n12731), .Z(n12734) );
  XNOR U12226 ( .A(n12729), .B(n12728), .Z(n12731) );
  XNOR U12227 ( .A(n12726), .B(n12725), .Z(n12728) );
  XNOR U12228 ( .A(n12723), .B(n12722), .Z(n12725) );
  XNOR U12229 ( .A(n12720), .B(n12719), .Z(n12722) );
  XNOR U12230 ( .A(n12717), .B(n12716), .Z(n12719) );
  XNOR U12231 ( .A(n12714), .B(n12713), .Z(n12716) );
  XNOR U12232 ( .A(n12711), .B(n12710), .Z(n12713) );
  XNOR U12233 ( .A(n12708), .B(n12707), .Z(n12710) );
  XNOR U12234 ( .A(n12705), .B(n12704), .Z(n12707) );
  XNOR U12235 ( .A(n12702), .B(n12701), .Z(n12704) );
  XNOR U12236 ( .A(n12699), .B(n12698), .Z(n12701) );
  XNOR U12237 ( .A(n12696), .B(n12695), .Z(n12698) );
  XNOR U12238 ( .A(n12693), .B(n12692), .Z(n12695) );
  XNOR U12239 ( .A(n12690), .B(n12689), .Z(n12692) );
  XNOR U12240 ( .A(n12687), .B(n12686), .Z(n12689) );
  XNOR U12241 ( .A(n12684), .B(n12683), .Z(n12686) );
  XNOR U12242 ( .A(n12681), .B(n12680), .Z(n12683) );
  XNOR U12243 ( .A(n12678), .B(n12677), .Z(n12680) );
  XNOR U12244 ( .A(n12675), .B(n12674), .Z(n12677) );
  XNOR U12245 ( .A(n12672), .B(n12671), .Z(n12674) );
  XNOR U12246 ( .A(n12669), .B(n12668), .Z(n12671) );
  XNOR U12247 ( .A(n12666), .B(n12665), .Z(n12668) );
  XNOR U12248 ( .A(n12663), .B(n12662), .Z(n12665) );
  XNOR U12249 ( .A(n12660), .B(n12659), .Z(n12662) );
  XNOR U12250 ( .A(n12657), .B(n12656), .Z(n12659) );
  XNOR U12251 ( .A(n12654), .B(n12653), .Z(n12656) );
  XNOR U12252 ( .A(n12651), .B(n12650), .Z(n12653) );
  XNOR U12253 ( .A(n12648), .B(n12647), .Z(n12650) );
  XNOR U12254 ( .A(n12645), .B(n12644), .Z(n12647) );
  XNOR U12255 ( .A(n12642), .B(n12641), .Z(n12644) );
  XNOR U12256 ( .A(n12639), .B(n12638), .Z(n12641) );
  XNOR U12257 ( .A(n12636), .B(n12635), .Z(n12638) );
  XNOR U12258 ( .A(n12633), .B(n12632), .Z(n12635) );
  XNOR U12259 ( .A(n12630), .B(n12629), .Z(n12632) );
  XNOR U12260 ( .A(n12627), .B(n12626), .Z(n12629) );
  XNOR U12261 ( .A(n12624), .B(n12623), .Z(n12626) );
  XNOR U12262 ( .A(n12621), .B(n12620), .Z(n12623) );
  XNOR U12263 ( .A(n12618), .B(n12617), .Z(n12620) );
  XNOR U12264 ( .A(n12615), .B(n12614), .Z(n12617) );
  XNOR U12265 ( .A(n12612), .B(n12611), .Z(n12614) );
  XNOR U12266 ( .A(n12609), .B(n12608), .Z(n12611) );
  XNOR U12267 ( .A(n12606), .B(n12605), .Z(n12608) );
  XNOR U12268 ( .A(n12603), .B(n12602), .Z(n12605) );
  XNOR U12269 ( .A(n12600), .B(n12599), .Z(n12602) );
  XNOR U12270 ( .A(n12597), .B(n12596), .Z(n12599) );
  XNOR U12271 ( .A(n12594), .B(n12593), .Z(n12596) );
  XNOR U12272 ( .A(n12591), .B(n12590), .Z(n12593) );
  XNOR U12273 ( .A(n12588), .B(n12587), .Z(n12590) );
  XNOR U12274 ( .A(n12585), .B(n12584), .Z(n12587) );
  XNOR U12275 ( .A(n12582), .B(n12581), .Z(n12584) );
  XNOR U12276 ( .A(n12579), .B(n12578), .Z(n12581) );
  XNOR U12277 ( .A(n12576), .B(n12575), .Z(n12578) );
  XNOR U12278 ( .A(n12573), .B(n12572), .Z(n12575) );
  XNOR U12279 ( .A(n12570), .B(n12569), .Z(n12572) );
  XNOR U12280 ( .A(n12567), .B(n12566), .Z(n12569) );
  XNOR U12281 ( .A(n12564), .B(n12563), .Z(n12566) );
  XNOR U12282 ( .A(n12561), .B(n12560), .Z(n12563) );
  XNOR U12283 ( .A(n12558), .B(n12557), .Z(n12560) );
  XNOR U12284 ( .A(n12555), .B(n12554), .Z(n12557) );
  XNOR U12285 ( .A(n12552), .B(n12551), .Z(n12554) );
  XNOR U12286 ( .A(n12549), .B(n12548), .Z(n12551) );
  XNOR U12287 ( .A(n12546), .B(n12545), .Z(n12548) );
  XNOR U12288 ( .A(n12543), .B(n12542), .Z(n12545) );
  XNOR U12289 ( .A(n12540), .B(n12539), .Z(n12542) );
  XNOR U12290 ( .A(n12537), .B(n12536), .Z(n12539) );
  XNOR U12291 ( .A(n12534), .B(n12533), .Z(n12536) );
  XNOR U12292 ( .A(n12531), .B(n12530), .Z(n12533) );
  XNOR U12293 ( .A(n12528), .B(n12527), .Z(n12530) );
  XNOR U12294 ( .A(n12525), .B(n12524), .Z(n12527) );
  XNOR U12295 ( .A(n12522), .B(n12521), .Z(n12524) );
  XNOR U12296 ( .A(n12519), .B(n12518), .Z(n12521) );
  XNOR U12297 ( .A(n12516), .B(n12515), .Z(n12518) );
  XNOR U12298 ( .A(n12513), .B(n12512), .Z(n12515) );
  XNOR U12299 ( .A(n12510), .B(n12509), .Z(n12512) );
  XNOR U12300 ( .A(n12507), .B(n12506), .Z(n12509) );
  XNOR U12301 ( .A(n12504), .B(n12503), .Z(n12506) );
  XNOR U12302 ( .A(n12501), .B(n12500), .Z(n12503) );
  XNOR U12303 ( .A(n12498), .B(n12497), .Z(n12500) );
  XOR U12304 ( .A(n13557), .B(n12494), .Z(n12497) );
  XOR U12305 ( .A(n12492), .B(n12491), .Z(n12494) );
  XOR U12306 ( .A(n12489), .B(n12488), .Z(n12491) );
  XOR U12307 ( .A(n12485), .B(n12486), .Z(n12488) );
  AND U12308 ( .A(n13558), .B(n13559), .Z(n12486) );
  XOR U12309 ( .A(n12482), .B(n12483), .Z(n12485) );
  AND U12310 ( .A(n13560), .B(n13561), .Z(n12483) );
  XOR U12311 ( .A(n12479), .B(n12480), .Z(n12482) );
  AND U12312 ( .A(n13562), .B(n13563), .Z(n12480) );
  XOR U12313 ( .A(n12476), .B(n12477), .Z(n12479) );
  AND U12314 ( .A(n13564), .B(n13565), .Z(n12477) );
  XNOR U12315 ( .A(n12259), .B(n12474), .Z(n12476) );
  AND U12316 ( .A(n13566), .B(n13567), .Z(n12474) );
  XOR U12317 ( .A(n12261), .B(n12260), .Z(n12259) );
  AND U12318 ( .A(n13568), .B(n13569), .Z(n12260) );
  XOR U12319 ( .A(n12263), .B(n12262), .Z(n12261) );
  AND U12320 ( .A(n13570), .B(n13571), .Z(n12262) );
  XOR U12321 ( .A(n12265), .B(n12264), .Z(n12263) );
  AND U12322 ( .A(n13572), .B(n13573), .Z(n12264) );
  XOR U12323 ( .A(n12267), .B(n12266), .Z(n12265) );
  AND U12324 ( .A(n13574), .B(n13575), .Z(n12266) );
  XOR U12325 ( .A(n12269), .B(n12268), .Z(n12267) );
  AND U12326 ( .A(n13576), .B(n13577), .Z(n12268) );
  XOR U12327 ( .A(n12271), .B(n12270), .Z(n12269) );
  AND U12328 ( .A(n13578), .B(n13579), .Z(n12270) );
  XOR U12329 ( .A(n12273), .B(n12272), .Z(n12271) );
  AND U12330 ( .A(n13580), .B(n13581), .Z(n12272) );
  XOR U12331 ( .A(n12275), .B(n12274), .Z(n12273) );
  AND U12332 ( .A(n13582), .B(n13583), .Z(n12274) );
  XOR U12333 ( .A(n12277), .B(n12276), .Z(n12275) );
  AND U12334 ( .A(n13584), .B(n13585), .Z(n12276) );
  XOR U12335 ( .A(n12279), .B(n12278), .Z(n12277) );
  AND U12336 ( .A(n13586), .B(n13587), .Z(n12278) );
  XOR U12337 ( .A(n12281), .B(n12280), .Z(n12279) );
  AND U12338 ( .A(n13588), .B(n13589), .Z(n12280) );
  XOR U12339 ( .A(n12283), .B(n12282), .Z(n12281) );
  AND U12340 ( .A(n13590), .B(n13591), .Z(n12282) );
  XOR U12341 ( .A(n12285), .B(n12284), .Z(n12283) );
  AND U12342 ( .A(n13592), .B(n13593), .Z(n12284) );
  XOR U12343 ( .A(n12287), .B(n12286), .Z(n12285) );
  AND U12344 ( .A(n13594), .B(n13595), .Z(n12286) );
  XOR U12345 ( .A(n12289), .B(n12288), .Z(n12287) );
  AND U12346 ( .A(n13596), .B(n13597), .Z(n12288) );
  XOR U12347 ( .A(n12291), .B(n12290), .Z(n12289) );
  AND U12348 ( .A(n13598), .B(n13599), .Z(n12290) );
  XOR U12349 ( .A(n12293), .B(n12292), .Z(n12291) );
  AND U12350 ( .A(n13600), .B(n13601), .Z(n12292) );
  XOR U12351 ( .A(n12295), .B(n12294), .Z(n12293) );
  AND U12352 ( .A(n13602), .B(n13603), .Z(n12294) );
  XOR U12353 ( .A(n12297), .B(n12296), .Z(n12295) );
  AND U12354 ( .A(n13604), .B(n13605), .Z(n12296) );
  XOR U12355 ( .A(n12299), .B(n12298), .Z(n12297) );
  AND U12356 ( .A(n13606), .B(n13607), .Z(n12298) );
  XOR U12357 ( .A(n12301), .B(n12300), .Z(n12299) );
  AND U12358 ( .A(n13608), .B(n13609), .Z(n12300) );
  XOR U12359 ( .A(n12303), .B(n12302), .Z(n12301) );
  AND U12360 ( .A(n13610), .B(n13611), .Z(n12302) );
  XOR U12361 ( .A(n12305), .B(n12304), .Z(n12303) );
  AND U12362 ( .A(n13612), .B(n13613), .Z(n12304) );
  XOR U12363 ( .A(n12307), .B(n12306), .Z(n12305) );
  AND U12364 ( .A(n13614), .B(n13615), .Z(n12306) );
  XOR U12365 ( .A(n12309), .B(n12308), .Z(n12307) );
  AND U12366 ( .A(n13616), .B(n13617), .Z(n12308) );
  XOR U12367 ( .A(n12311), .B(n12310), .Z(n12309) );
  AND U12368 ( .A(n13618), .B(n13619), .Z(n12310) );
  XOR U12369 ( .A(n12313), .B(n12312), .Z(n12311) );
  AND U12370 ( .A(n13620), .B(n13621), .Z(n12312) );
  XOR U12371 ( .A(n12315), .B(n12314), .Z(n12313) );
  AND U12372 ( .A(n13622), .B(n13623), .Z(n12314) );
  XOR U12373 ( .A(n12317), .B(n12316), .Z(n12315) );
  AND U12374 ( .A(n13624), .B(n13625), .Z(n12316) );
  XOR U12375 ( .A(n12319), .B(n12318), .Z(n12317) );
  AND U12376 ( .A(n13626), .B(n13627), .Z(n12318) );
  XOR U12377 ( .A(n12321), .B(n12320), .Z(n12319) );
  AND U12378 ( .A(n13628), .B(n13629), .Z(n12320) );
  XOR U12379 ( .A(n12323), .B(n12322), .Z(n12321) );
  AND U12380 ( .A(n13630), .B(n13631), .Z(n12322) );
  XOR U12381 ( .A(n12325), .B(n12324), .Z(n12323) );
  AND U12382 ( .A(n13632), .B(n13633), .Z(n12324) );
  XOR U12383 ( .A(n12327), .B(n12326), .Z(n12325) );
  AND U12384 ( .A(n13634), .B(n13635), .Z(n12326) );
  XOR U12385 ( .A(n12329), .B(n12328), .Z(n12327) );
  AND U12386 ( .A(n13636), .B(n13637), .Z(n12328) );
  XOR U12387 ( .A(n12331), .B(n12330), .Z(n12329) );
  AND U12388 ( .A(n13638), .B(n13639), .Z(n12330) );
  XOR U12389 ( .A(n12333), .B(n12332), .Z(n12331) );
  AND U12390 ( .A(n13640), .B(n13641), .Z(n12332) );
  XOR U12391 ( .A(n12335), .B(n12334), .Z(n12333) );
  AND U12392 ( .A(n13642), .B(n13643), .Z(n12334) );
  XOR U12393 ( .A(n12337), .B(n12336), .Z(n12335) );
  AND U12394 ( .A(n13644), .B(n13645), .Z(n12336) );
  XOR U12395 ( .A(n12470), .B(n12338), .Z(n12337) );
  AND U12396 ( .A(n13646), .B(n13647), .Z(n12338) );
  XOR U12397 ( .A(n12472), .B(n12471), .Z(n12470) );
  AND U12398 ( .A(n13648), .B(n13649), .Z(n12471) );
  XOR U12399 ( .A(n12453), .B(n12473), .Z(n12472) );
  AND U12400 ( .A(n13650), .B(n13651), .Z(n12473) );
  XOR U12401 ( .A(n12455), .B(n12454), .Z(n12453) );
  AND U12402 ( .A(n13652), .B(n13653), .Z(n12454) );
  XOR U12403 ( .A(n12457), .B(n12456), .Z(n12455) );
  AND U12404 ( .A(n13654), .B(n13655), .Z(n12456) );
  XOR U12405 ( .A(n12461), .B(n12458), .Z(n12457) );
  AND U12406 ( .A(n13656), .B(n13657), .Z(n12458) );
  XOR U12407 ( .A(n12463), .B(n12462), .Z(n12461) );
  AND U12408 ( .A(n13658), .B(n13659), .Z(n12462) );
  XOR U12409 ( .A(n12466), .B(n12464), .Z(n12463) );
  AND U12410 ( .A(n13660), .B(n13661), .Z(n12464) );
  XOR U12411 ( .A(n12468), .B(n12467), .Z(n12466) );
  AND U12412 ( .A(n13662), .B(n13663), .Z(n12467) );
  XOR U12413 ( .A(n12353), .B(n12469), .Z(n12468) );
  AND U12414 ( .A(n13664), .B(n13665), .Z(n12469) );
  XNOR U12415 ( .A(n12360), .B(n12354), .Z(n12353) );
  AND U12416 ( .A(n13666), .B(n13667), .Z(n12354) );
  XOR U12417 ( .A(n12359), .B(n12351), .Z(n12360) );
  AND U12418 ( .A(n13668), .B(n13669), .Z(n12351) );
  XOR U12419 ( .A(n12452), .B(n12350), .Z(n12359) );
  AND U12420 ( .A(n13670), .B(n13671), .Z(n12350) );
  XNOR U12421 ( .A(n12371), .B(n12349), .Z(n12452) );
  AND U12422 ( .A(n13672), .B(n13673), .Z(n12349) );
  XNOR U12423 ( .A(n12378), .B(n12372), .Z(n12371) );
  AND U12424 ( .A(n13674), .B(n13675), .Z(n12372) );
  XOR U12425 ( .A(n12377), .B(n12369), .Z(n12378) );
  AND U12426 ( .A(n13676), .B(n13677), .Z(n12369) );
  XOR U12427 ( .A(n12451), .B(n12368), .Z(n12377) );
  AND U12428 ( .A(n13678), .B(n13679), .Z(n12368) );
  XNOR U12429 ( .A(n12389), .B(n12367), .Z(n12451) );
  AND U12430 ( .A(n13680), .B(n13681), .Z(n12367) );
  XNOR U12431 ( .A(n12396), .B(n12390), .Z(n12389) );
  AND U12432 ( .A(n13682), .B(n13683), .Z(n12390) );
  XOR U12433 ( .A(n12395), .B(n12387), .Z(n12396) );
  AND U12434 ( .A(n13684), .B(n13685), .Z(n12387) );
  XOR U12435 ( .A(n12450), .B(n12386), .Z(n12395) );
  AND U12436 ( .A(n13686), .B(n13687), .Z(n12386) );
  XNOR U12437 ( .A(n12407), .B(n12385), .Z(n12450) );
  AND U12438 ( .A(n13688), .B(n13689), .Z(n12385) );
  XNOR U12439 ( .A(n12414), .B(n12408), .Z(n12407) );
  AND U12440 ( .A(n13690), .B(n13691), .Z(n12408) );
  XOR U12441 ( .A(n12413), .B(n12405), .Z(n12414) );
  AND U12442 ( .A(n13692), .B(n13693), .Z(n12405) );
  XOR U12443 ( .A(n12449), .B(n12404), .Z(n12413) );
  AND U12444 ( .A(n13694), .B(n13695), .Z(n12404) );
  XNOR U12445 ( .A(n13696), .B(n13697), .Z(n12449) );
  XOR U12446 ( .A(n12447), .B(n12448), .Z(n13697) );
  AND U12447 ( .A(n13698), .B(n13699), .Z(n12448) );
  AND U12448 ( .A(n13700), .B(n13701), .Z(n12447) );
  XOR U12449 ( .A(n13702), .B(n12403), .Z(n13696) );
  AND U12450 ( .A(n13703), .B(n13704), .Z(n12403) );
  XOR U12451 ( .A(n13705), .B(n13706), .Z(n13702) );
  XOR U12452 ( .A(n13707), .B(n13708), .Z(n13706) );
  XOR U12453 ( .A(n12440), .B(n12441), .Z(n13708) );
  AND U12454 ( .A(n13709), .B(n13710), .Z(n12441) );
  AND U12455 ( .A(n13711), .B(n13712), .Z(n12440) );
  XOR U12456 ( .A(n12434), .B(n12439), .Z(n13707) );
  AND U12457 ( .A(n13713), .B(n13714), .Z(n12439) );
  AND U12458 ( .A(n13715), .B(n13716), .Z(n12434) );
  XOR U12459 ( .A(n13717), .B(n13718), .Z(n13705) );
  XOR U12460 ( .A(n12442), .B(n12445), .Z(n13718) );
  AND U12461 ( .A(n13719), .B(n13720), .Z(n12445) );
  AND U12462 ( .A(n13721), .B(n13722), .Z(n12442) );
  XOR U12463 ( .A(n13723), .B(n12446), .Z(n13717) );
  AND U12464 ( .A(n13724), .B(n13725), .Z(n12446) );
  XOR U12465 ( .A(n13726), .B(n13727), .Z(n13723) );
  XOR U12466 ( .A(n13728), .B(n13729), .Z(n13727) );
  XOR U12467 ( .A(n12427), .B(n12428), .Z(n13729) );
  AND U12468 ( .A(n13730), .B(n13731), .Z(n12428) );
  AND U12469 ( .A(n13732), .B(n13733), .Z(n12427) );
  XNOR U12470 ( .A(n12425), .B(n12424), .Z(n13728) );
  IV U12471 ( .A(n13734), .Z(n12424) );
  AND U12472 ( .A(n13735), .B(n13736), .Z(n13734) );
  AND U12473 ( .A(n13737), .B(n13738), .Z(n12425) );
  XOR U12474 ( .A(n13739), .B(n13740), .Z(n13726) );
  XOR U12475 ( .A(n12431), .B(n12432), .Z(n13740) );
  AND U12476 ( .A(n13741), .B(n13742), .Z(n12432) );
  AND U12477 ( .A(n13743), .B(n13744), .Z(n12431) );
  XOR U12478 ( .A(n12426), .B(n12433), .Z(n13739) );
  AND U12479 ( .A(n13745), .B(n13746), .Z(n12433) );
  XNOR U12480 ( .A(n13747), .B(n13748), .Z(n12426) );
  AND U12481 ( .A(n13749), .B(n13750), .Z(n13748) );
  NOR U12482 ( .A(n13751), .B(n13752), .Z(n13750) );
  NOR U12483 ( .A(n13753), .B(n13754), .Z(n13749) );
  AND U12484 ( .A(n13755), .B(n13756), .Z(n13754) );
  AND U12485 ( .A(n13757), .B(n13758), .Z(n13747) );
  NOR U12486 ( .A(n13759), .B(n13760), .Z(n13758) );
  AND U12487 ( .A(n13752), .B(n13761), .Z(n13760) );
  AND U12488 ( .A(n13753), .B(n13762), .Z(n13759) );
  NOR U12489 ( .A(n13763), .B(n13764), .Z(n13757) );
  XOR U12490 ( .A(n13765), .B(n13766), .Z(n13764) );
  AND U12491 ( .A(n13767), .B(n13768), .Z(n13766) );
  NOR U12492 ( .A(n13769), .B(n13770), .Z(n13768) );
  NOR U12493 ( .A(n13771), .B(n13772), .Z(n13767) );
  AND U12494 ( .A(n13773), .B(n13774), .Z(n13772) );
  AND U12495 ( .A(n13775), .B(n13776), .Z(n13765) );
  NOR U12496 ( .A(n13777), .B(n13778), .Z(n13776) );
  AND U12497 ( .A(n13770), .B(n13779), .Z(n13778) );
  AND U12498 ( .A(n13771), .B(n13780), .Z(n13777) );
  NOR U12499 ( .A(n13781), .B(n13782), .Z(n13775) );
  AND U12500 ( .A(n13783), .B(n13784), .Z(n13782) );
  AND U12501 ( .A(n13785), .B(n13786), .Z(n13784) );
  AND U12502 ( .A(n13787), .B(n13788), .Z(n13786) );
  NOR U12503 ( .A(n13789), .B(n13790), .Z(n13787) );
  NOR U12504 ( .A(n13791), .B(n13792), .Z(n13785) );
  AND U12505 ( .A(n13793), .B(n13794), .Z(n13783) );
  NOR U12506 ( .A(n13795), .B(n13796), .Z(n13794) );
  NOR U12507 ( .A(n13797), .B(n13798), .Z(n13793) );
  AND U12508 ( .A(n13769), .B(n13799), .Z(n13781) );
  AND U12509 ( .A(n13751), .B(n13800), .Z(n13763) );
  XOR U12510 ( .A(n13801), .B(n13802), .Z(n12489) );
  AND U12511 ( .A(n13801), .B(n13803), .Z(n13802) );
  XNOR U12512 ( .A(n13804), .B(n13805), .Z(n12492) );
  AND U12513 ( .A(n13804), .B(n13806), .Z(n13805) );
  IV U12514 ( .A(n12495), .Z(n13557) );
  XNOR U12515 ( .A(n13807), .B(n13808), .Z(n12495) );
  AND U12516 ( .A(n13807), .B(n13809), .Z(n13808) );
  XNOR U12517 ( .A(n13810), .B(n13811), .Z(n12498) );
  AND U12518 ( .A(n13810), .B(n13812), .Z(n13811) );
  XNOR U12519 ( .A(n13813), .B(n13814), .Z(n12501) );
  AND U12520 ( .A(n13815), .B(n13813), .Z(n13814) );
  XOR U12521 ( .A(n13816), .B(n13817), .Z(n12504) );
  NOR U12522 ( .A(n13818), .B(n13816), .Z(n13817) );
  XOR U12523 ( .A(n13819), .B(n13820), .Z(n12507) );
  NOR U12524 ( .A(n13821), .B(n13819), .Z(n13820) );
  XOR U12525 ( .A(n13822), .B(n13823), .Z(n12510) );
  NOR U12526 ( .A(n13824), .B(n13822), .Z(n13823) );
  XOR U12527 ( .A(n13825), .B(n13826), .Z(n12513) );
  NOR U12528 ( .A(n13827), .B(n13825), .Z(n13826) );
  XOR U12529 ( .A(n13828), .B(n13829), .Z(n12516) );
  NOR U12530 ( .A(n13830), .B(n13828), .Z(n13829) );
  XOR U12531 ( .A(n13831), .B(n13832), .Z(n12519) );
  NOR U12532 ( .A(n13833), .B(n13831), .Z(n13832) );
  XOR U12533 ( .A(n13834), .B(n13835), .Z(n12522) );
  NOR U12534 ( .A(n13836), .B(n13834), .Z(n13835) );
  XOR U12535 ( .A(n13837), .B(n13838), .Z(n12525) );
  NOR U12536 ( .A(n13839), .B(n13837), .Z(n13838) );
  XOR U12537 ( .A(n13840), .B(n13841), .Z(n12528) );
  NOR U12538 ( .A(n13842), .B(n13840), .Z(n13841) );
  XOR U12539 ( .A(n13843), .B(n13844), .Z(n12531) );
  NOR U12540 ( .A(n13845), .B(n13843), .Z(n13844) );
  XOR U12541 ( .A(n13846), .B(n13847), .Z(n12534) );
  NOR U12542 ( .A(n13848), .B(n13846), .Z(n13847) );
  XOR U12543 ( .A(n13849), .B(n13850), .Z(n12537) );
  NOR U12544 ( .A(n13851), .B(n13849), .Z(n13850) );
  XOR U12545 ( .A(n13852), .B(n13853), .Z(n12540) );
  NOR U12546 ( .A(n13854), .B(n13852), .Z(n13853) );
  XOR U12547 ( .A(n13855), .B(n13856), .Z(n12543) );
  NOR U12548 ( .A(n13857), .B(n13855), .Z(n13856) );
  XOR U12549 ( .A(n13858), .B(n13859), .Z(n12546) );
  NOR U12550 ( .A(n13860), .B(n13858), .Z(n13859) );
  XOR U12551 ( .A(n13861), .B(n13862), .Z(n12549) );
  NOR U12552 ( .A(n13863), .B(n13861), .Z(n13862) );
  XOR U12553 ( .A(n13864), .B(n13865), .Z(n12552) );
  NOR U12554 ( .A(n13866), .B(n13864), .Z(n13865) );
  XOR U12555 ( .A(n13867), .B(n13868), .Z(n12555) );
  NOR U12556 ( .A(n13869), .B(n13867), .Z(n13868) );
  XOR U12557 ( .A(n13870), .B(n13871), .Z(n12558) );
  NOR U12558 ( .A(n13872), .B(n13870), .Z(n13871) );
  XOR U12559 ( .A(n13873), .B(n13874), .Z(n12561) );
  NOR U12560 ( .A(n13875), .B(n13873), .Z(n13874) );
  XOR U12561 ( .A(n13876), .B(n13877), .Z(n12564) );
  NOR U12562 ( .A(n13878), .B(n13876), .Z(n13877) );
  XOR U12563 ( .A(n13879), .B(n13880), .Z(n12567) );
  NOR U12564 ( .A(n13881), .B(n13879), .Z(n13880) );
  XOR U12565 ( .A(n13882), .B(n13883), .Z(n12570) );
  NOR U12566 ( .A(n13884), .B(n13882), .Z(n13883) );
  XOR U12567 ( .A(n13885), .B(n13886), .Z(n12573) );
  NOR U12568 ( .A(n13887), .B(n13885), .Z(n13886) );
  XOR U12569 ( .A(n13888), .B(n13889), .Z(n12576) );
  NOR U12570 ( .A(n13890), .B(n13888), .Z(n13889) );
  XOR U12571 ( .A(n13891), .B(n13892), .Z(n12579) );
  NOR U12572 ( .A(n13893), .B(n13891), .Z(n13892) );
  XOR U12573 ( .A(n13894), .B(n13895), .Z(n12582) );
  NOR U12574 ( .A(n13896), .B(n13894), .Z(n13895) );
  XOR U12575 ( .A(n13897), .B(n13898), .Z(n12585) );
  NOR U12576 ( .A(n13899), .B(n13897), .Z(n13898) );
  XOR U12577 ( .A(n13900), .B(n13901), .Z(n12588) );
  NOR U12578 ( .A(n13902), .B(n13900), .Z(n13901) );
  XOR U12579 ( .A(n13903), .B(n13904), .Z(n12591) );
  NOR U12580 ( .A(n13905), .B(n13903), .Z(n13904) );
  XOR U12581 ( .A(n13906), .B(n13907), .Z(n12594) );
  NOR U12582 ( .A(n13908), .B(n13906), .Z(n13907) );
  XOR U12583 ( .A(n13909), .B(n13910), .Z(n12597) );
  NOR U12584 ( .A(n13911), .B(n13909), .Z(n13910) );
  XOR U12585 ( .A(n13912), .B(n13913), .Z(n12600) );
  NOR U12586 ( .A(n13914), .B(n13912), .Z(n13913) );
  XOR U12587 ( .A(n13915), .B(n13916), .Z(n12603) );
  NOR U12588 ( .A(n13917), .B(n13915), .Z(n13916) );
  XOR U12589 ( .A(n13918), .B(n13919), .Z(n12606) );
  NOR U12590 ( .A(n13920), .B(n13918), .Z(n13919) );
  XOR U12591 ( .A(n13921), .B(n13922), .Z(n12609) );
  NOR U12592 ( .A(n13923), .B(n13921), .Z(n13922) );
  XOR U12593 ( .A(n13924), .B(n13925), .Z(n12612) );
  NOR U12594 ( .A(n13926), .B(n13924), .Z(n13925) );
  XOR U12595 ( .A(n13927), .B(n13928), .Z(n12615) );
  NOR U12596 ( .A(n13929), .B(n13927), .Z(n13928) );
  XOR U12597 ( .A(n13930), .B(n13931), .Z(n12618) );
  NOR U12598 ( .A(n13932), .B(n13930), .Z(n13931) );
  XOR U12599 ( .A(n13933), .B(n13934), .Z(n12621) );
  NOR U12600 ( .A(n13935), .B(n13933), .Z(n13934) );
  XOR U12601 ( .A(n13936), .B(n13937), .Z(n12624) );
  NOR U12602 ( .A(n13938), .B(n13936), .Z(n13937) );
  XOR U12603 ( .A(n13939), .B(n13940), .Z(n12627) );
  NOR U12604 ( .A(n13941), .B(n13939), .Z(n13940) );
  XOR U12605 ( .A(n13942), .B(n13943), .Z(n12630) );
  NOR U12606 ( .A(n13944), .B(n13942), .Z(n13943) );
  XOR U12607 ( .A(n13945), .B(n13946), .Z(n12633) );
  NOR U12608 ( .A(n13947), .B(n13945), .Z(n13946) );
  XOR U12609 ( .A(n13948), .B(n13949), .Z(n12636) );
  NOR U12610 ( .A(n13950), .B(n13948), .Z(n13949) );
  XOR U12611 ( .A(n13951), .B(n13952), .Z(n12639) );
  NOR U12612 ( .A(n13953), .B(n13951), .Z(n13952) );
  XOR U12613 ( .A(n13954), .B(n13955), .Z(n12642) );
  NOR U12614 ( .A(n13956), .B(n13954), .Z(n13955) );
  XOR U12615 ( .A(n13957), .B(n13958), .Z(n12645) );
  NOR U12616 ( .A(n13959), .B(n13957), .Z(n13958) );
  XOR U12617 ( .A(n13960), .B(n13961), .Z(n12648) );
  NOR U12618 ( .A(n13962), .B(n13960), .Z(n13961) );
  XOR U12619 ( .A(n13963), .B(n13964), .Z(n12651) );
  NOR U12620 ( .A(n13965), .B(n13963), .Z(n13964) );
  XOR U12621 ( .A(n13966), .B(n13967), .Z(n12654) );
  NOR U12622 ( .A(n13968), .B(n13966), .Z(n13967) );
  XOR U12623 ( .A(n13969), .B(n13970), .Z(n12657) );
  NOR U12624 ( .A(n13971), .B(n13969), .Z(n13970) );
  XOR U12625 ( .A(n13972), .B(n13973), .Z(n12660) );
  NOR U12626 ( .A(n13974), .B(n13972), .Z(n13973) );
  XOR U12627 ( .A(n13975), .B(n13976), .Z(n12663) );
  NOR U12628 ( .A(n13977), .B(n13975), .Z(n13976) );
  XOR U12629 ( .A(n13978), .B(n13979), .Z(n12666) );
  NOR U12630 ( .A(n13980), .B(n13978), .Z(n13979) );
  XOR U12631 ( .A(n13981), .B(n13982), .Z(n12669) );
  NOR U12632 ( .A(n13983), .B(n13981), .Z(n13982) );
  XOR U12633 ( .A(n13984), .B(n13985), .Z(n12672) );
  NOR U12634 ( .A(n13986), .B(n13984), .Z(n13985) );
  XOR U12635 ( .A(n13987), .B(n13988), .Z(n12675) );
  NOR U12636 ( .A(n13989), .B(n13987), .Z(n13988) );
  XOR U12637 ( .A(n13990), .B(n13991), .Z(n12678) );
  NOR U12638 ( .A(n13992), .B(n13990), .Z(n13991) );
  XOR U12639 ( .A(n13993), .B(n13994), .Z(n12681) );
  NOR U12640 ( .A(n13995), .B(n13993), .Z(n13994) );
  XOR U12641 ( .A(n13996), .B(n13997), .Z(n12684) );
  NOR U12642 ( .A(n13998), .B(n13996), .Z(n13997) );
  XOR U12643 ( .A(n13999), .B(n14000), .Z(n12687) );
  NOR U12644 ( .A(n14001), .B(n13999), .Z(n14000) );
  XOR U12645 ( .A(n14002), .B(n14003), .Z(n12690) );
  NOR U12646 ( .A(n14004), .B(n14002), .Z(n14003) );
  XOR U12647 ( .A(n14005), .B(n14006), .Z(n12693) );
  NOR U12648 ( .A(n14007), .B(n14005), .Z(n14006) );
  XOR U12649 ( .A(n14008), .B(n14009), .Z(n12696) );
  NOR U12650 ( .A(n14010), .B(n14008), .Z(n14009) );
  XOR U12651 ( .A(n14011), .B(n14012), .Z(n12699) );
  NOR U12652 ( .A(n14013), .B(n14011), .Z(n14012) );
  XOR U12653 ( .A(n14014), .B(n14015), .Z(n12702) );
  NOR U12654 ( .A(n14016), .B(n14014), .Z(n14015) );
  XOR U12655 ( .A(n14017), .B(n14018), .Z(n12705) );
  NOR U12656 ( .A(n14019), .B(n14017), .Z(n14018) );
  XOR U12657 ( .A(n14020), .B(n14021), .Z(n12708) );
  NOR U12658 ( .A(n14022), .B(n14020), .Z(n14021) );
  XOR U12659 ( .A(n14023), .B(n14024), .Z(n12711) );
  NOR U12660 ( .A(n14025), .B(n14023), .Z(n14024) );
  XOR U12661 ( .A(n14026), .B(n14027), .Z(n12714) );
  NOR U12662 ( .A(n14028), .B(n14026), .Z(n14027) );
  XOR U12663 ( .A(n14029), .B(n14030), .Z(n12717) );
  NOR U12664 ( .A(n14031), .B(n14029), .Z(n14030) );
  XOR U12665 ( .A(n14032), .B(n14033), .Z(n12720) );
  NOR U12666 ( .A(n14034), .B(n14032), .Z(n14033) );
  XOR U12667 ( .A(n14035), .B(n14036), .Z(n12723) );
  NOR U12668 ( .A(n14037), .B(n14035), .Z(n14036) );
  XOR U12669 ( .A(n14038), .B(n14039), .Z(n12726) );
  NOR U12670 ( .A(n14040), .B(n14038), .Z(n14039) );
  XOR U12671 ( .A(n14041), .B(n14042), .Z(n12729) );
  NOR U12672 ( .A(n14043), .B(n14041), .Z(n14042) );
  XOR U12673 ( .A(n14044), .B(n14045), .Z(n12732) );
  NOR U12674 ( .A(n14046), .B(n14044), .Z(n14045) );
  XOR U12675 ( .A(n14047), .B(n14048), .Z(n12735) );
  NOR U12676 ( .A(n14049), .B(n14047), .Z(n14048) );
  XOR U12677 ( .A(n14050), .B(n14051), .Z(n12738) );
  NOR U12678 ( .A(n14052), .B(n14050), .Z(n14051) );
  XOR U12679 ( .A(n14053), .B(n14054), .Z(n12741) );
  NOR U12680 ( .A(n14055), .B(n14053), .Z(n14054) );
  XOR U12681 ( .A(n14056), .B(n14057), .Z(n12744) );
  NOR U12682 ( .A(n14058), .B(n14056), .Z(n14057) );
  XOR U12683 ( .A(n14059), .B(n14060), .Z(n12747) );
  NOR U12684 ( .A(n14061), .B(n14059), .Z(n14060) );
  XOR U12685 ( .A(n14062), .B(n14063), .Z(n12750) );
  NOR U12686 ( .A(n14064), .B(n14062), .Z(n14063) );
  XOR U12687 ( .A(n14065), .B(n14066), .Z(n12753) );
  NOR U12688 ( .A(n14067), .B(n14065), .Z(n14066) );
  XOR U12689 ( .A(n14068), .B(n14069), .Z(n12756) );
  NOR U12690 ( .A(n14070), .B(n14068), .Z(n14069) );
  XOR U12691 ( .A(n14071), .B(n14072), .Z(n12759) );
  NOR U12692 ( .A(n14073), .B(n14071), .Z(n14072) );
  XOR U12693 ( .A(n14074), .B(n14075), .Z(n12762) );
  NOR U12694 ( .A(n14076), .B(n14074), .Z(n14075) );
  XOR U12695 ( .A(n14077), .B(n14078), .Z(n12765) );
  NOR U12696 ( .A(n14079), .B(n14077), .Z(n14078) );
  XOR U12697 ( .A(n14080), .B(n14081), .Z(n12768) );
  NOR U12698 ( .A(n14082), .B(n14080), .Z(n14081) );
  XOR U12699 ( .A(n14083), .B(n14084), .Z(n12771) );
  NOR U12700 ( .A(n14085), .B(n14083), .Z(n14084) );
  XOR U12701 ( .A(n14086), .B(n14087), .Z(n12774) );
  NOR U12702 ( .A(n14088), .B(n14086), .Z(n14087) );
  XOR U12703 ( .A(n14089), .B(n14090), .Z(n12777) );
  NOR U12704 ( .A(n14091), .B(n14089), .Z(n14090) );
  XOR U12705 ( .A(n14092), .B(n14093), .Z(n12780) );
  NOR U12706 ( .A(n14094), .B(n14092), .Z(n14093) );
  XOR U12707 ( .A(n14095), .B(n14096), .Z(n12783) );
  NOR U12708 ( .A(n14097), .B(n14095), .Z(n14096) );
  XOR U12709 ( .A(n14098), .B(n14099), .Z(n12786) );
  NOR U12710 ( .A(n14100), .B(n14098), .Z(n14099) );
  XOR U12711 ( .A(n14101), .B(n14102), .Z(n12789) );
  NOR U12712 ( .A(n14103), .B(n14101), .Z(n14102) );
  XOR U12713 ( .A(n14104), .B(n14105), .Z(n12792) );
  NOR U12714 ( .A(n14106), .B(n14104), .Z(n14105) );
  XOR U12715 ( .A(n14107), .B(n14108), .Z(n12795) );
  NOR U12716 ( .A(n14109), .B(n14107), .Z(n14108) );
  XOR U12717 ( .A(n14110), .B(n14111), .Z(n12798) );
  NOR U12718 ( .A(n14112), .B(n14110), .Z(n14111) );
  XOR U12719 ( .A(n14113), .B(n14114), .Z(n12801) );
  NOR U12720 ( .A(n14115), .B(n14113), .Z(n14114) );
  XOR U12721 ( .A(n14116), .B(n14117), .Z(n12804) );
  NOR U12722 ( .A(n14118), .B(n14116), .Z(n14117) );
  XOR U12723 ( .A(n14119), .B(n14120), .Z(n12807) );
  NOR U12724 ( .A(n14121), .B(n14119), .Z(n14120) );
  XOR U12725 ( .A(n14122), .B(n14123), .Z(n12810) );
  NOR U12726 ( .A(n14124), .B(n14122), .Z(n14123) );
  XOR U12727 ( .A(n14125), .B(n14126), .Z(n12813) );
  NOR U12728 ( .A(n14127), .B(n14125), .Z(n14126) );
  XOR U12729 ( .A(n14128), .B(n14129), .Z(n12816) );
  NOR U12730 ( .A(n14130), .B(n14128), .Z(n14129) );
  XOR U12731 ( .A(n14131), .B(n14132), .Z(n12819) );
  NOR U12732 ( .A(n14133), .B(n14131), .Z(n14132) );
  XOR U12733 ( .A(n14134), .B(n14135), .Z(n12822) );
  NOR U12734 ( .A(n14136), .B(n14134), .Z(n14135) );
  XOR U12735 ( .A(n14137), .B(n14138), .Z(n12825) );
  NOR U12736 ( .A(n14139), .B(n14137), .Z(n14138) );
  XOR U12737 ( .A(n14140), .B(n14141), .Z(n12828) );
  NOR U12738 ( .A(n14142), .B(n14140), .Z(n14141) );
  XOR U12739 ( .A(n14143), .B(n14144), .Z(n12831) );
  NOR U12740 ( .A(n14145), .B(n14143), .Z(n14144) );
  XOR U12741 ( .A(n14146), .B(n14147), .Z(n12834) );
  NOR U12742 ( .A(n14148), .B(n14146), .Z(n14147) );
  XOR U12743 ( .A(n14149), .B(n14150), .Z(n12837) );
  NOR U12744 ( .A(n14151), .B(n14149), .Z(n14150) );
  XOR U12745 ( .A(n14152), .B(n14153), .Z(n12840) );
  NOR U12746 ( .A(n14154), .B(n14152), .Z(n14153) );
  XOR U12747 ( .A(n14155), .B(n14156), .Z(n12843) );
  NOR U12748 ( .A(n14157), .B(n14155), .Z(n14156) );
  XOR U12749 ( .A(n14158), .B(n14159), .Z(n12846) );
  NOR U12750 ( .A(n14160), .B(n14158), .Z(n14159) );
  XOR U12751 ( .A(n14161), .B(n14162), .Z(n12849) );
  NOR U12752 ( .A(n14163), .B(n14161), .Z(n14162) );
  XOR U12753 ( .A(n14164), .B(n14165), .Z(n12852) );
  NOR U12754 ( .A(n14166), .B(n14164), .Z(n14165) );
  XOR U12755 ( .A(n14167), .B(n14168), .Z(n12855) );
  NOR U12756 ( .A(n14169), .B(n14167), .Z(n14168) );
  XOR U12757 ( .A(n14170), .B(n14171), .Z(n12858) );
  NOR U12758 ( .A(n14172), .B(n14170), .Z(n14171) );
  XOR U12759 ( .A(n14173), .B(n14174), .Z(n12861) );
  NOR U12760 ( .A(n14175), .B(n14173), .Z(n14174) );
  XOR U12761 ( .A(n14176), .B(n14177), .Z(n12864) );
  NOR U12762 ( .A(n14178), .B(n14176), .Z(n14177) );
  XOR U12763 ( .A(n14179), .B(n14180), .Z(n12867) );
  NOR U12764 ( .A(n14181), .B(n14179), .Z(n14180) );
  XOR U12765 ( .A(n14182), .B(n14183), .Z(n12870) );
  NOR U12766 ( .A(n14184), .B(n14182), .Z(n14183) );
  XOR U12767 ( .A(n14185), .B(n14186), .Z(n12873) );
  NOR U12768 ( .A(n14187), .B(n14185), .Z(n14186) );
  XOR U12769 ( .A(n14188), .B(n14189), .Z(n12876) );
  NOR U12770 ( .A(n14190), .B(n14188), .Z(n14189) );
  XOR U12771 ( .A(n14191), .B(n14192), .Z(n12879) );
  NOR U12772 ( .A(n14193), .B(n14191), .Z(n14192) );
  XOR U12773 ( .A(n14194), .B(n14195), .Z(n12882) );
  NOR U12774 ( .A(n14196), .B(n14194), .Z(n14195) );
  XOR U12775 ( .A(n14197), .B(n14198), .Z(n12885) );
  NOR U12776 ( .A(n14199), .B(n14197), .Z(n14198) );
  XOR U12777 ( .A(n14200), .B(n14201), .Z(n12888) );
  NOR U12778 ( .A(n14202), .B(n14200), .Z(n14201) );
  XOR U12779 ( .A(n14203), .B(n14204), .Z(n12891) );
  NOR U12780 ( .A(n14205), .B(n14203), .Z(n14204) );
  XOR U12781 ( .A(n14206), .B(n14207), .Z(n12894) );
  NOR U12782 ( .A(n14208), .B(n14206), .Z(n14207) );
  XOR U12783 ( .A(n14209), .B(n14210), .Z(n12897) );
  NOR U12784 ( .A(n14211), .B(n14209), .Z(n14210) );
  XOR U12785 ( .A(n14212), .B(n14213), .Z(n12900) );
  AND U12786 ( .A(n14214), .B(n14212), .Z(n14213) );
  XOR U12787 ( .A(n14215), .B(n14216), .Z(n12903) );
  AND U12788 ( .A(n93), .B(n14215), .Z(n14216) );
  XOR U12789 ( .A(n75), .B(n13553), .Z(n13555) );
  XOR U12790 ( .A(n13550), .B(n13549), .Z(n75) );
  XNOR U12791 ( .A(n13547), .B(n13546), .Z(n13549) );
  XNOR U12792 ( .A(n13544), .B(n13543), .Z(n13546) );
  XNOR U12793 ( .A(n13541), .B(n13540), .Z(n13543) );
  XNOR U12794 ( .A(n13538), .B(n13537), .Z(n13540) );
  XNOR U12795 ( .A(n13535), .B(n13534), .Z(n13537) );
  XNOR U12796 ( .A(n13532), .B(n13531), .Z(n13534) );
  XNOR U12797 ( .A(n13529), .B(n13528), .Z(n13531) );
  XNOR U12798 ( .A(n13526), .B(n13525), .Z(n13528) );
  XNOR U12799 ( .A(n13523), .B(n13522), .Z(n13525) );
  XNOR U12800 ( .A(n13520), .B(n13519), .Z(n13522) );
  XNOR U12801 ( .A(n13517), .B(n13516), .Z(n13519) );
  XNOR U12802 ( .A(n13514), .B(n13513), .Z(n13516) );
  XNOR U12803 ( .A(n13511), .B(n13510), .Z(n13513) );
  XNOR U12804 ( .A(n13508), .B(n13507), .Z(n13510) );
  XNOR U12805 ( .A(n13505), .B(n13504), .Z(n13507) );
  XNOR U12806 ( .A(n13502), .B(n13501), .Z(n13504) );
  XNOR U12807 ( .A(n13499), .B(n13498), .Z(n13501) );
  XNOR U12808 ( .A(n13496), .B(n13495), .Z(n13498) );
  XNOR U12809 ( .A(n13493), .B(n13492), .Z(n13495) );
  XNOR U12810 ( .A(n13490), .B(n13489), .Z(n13492) );
  XNOR U12811 ( .A(n13487), .B(n13486), .Z(n13489) );
  XNOR U12812 ( .A(n13484), .B(n13483), .Z(n13486) );
  XNOR U12813 ( .A(n13481), .B(n13480), .Z(n13483) );
  XNOR U12814 ( .A(n13478), .B(n13477), .Z(n13480) );
  XNOR U12815 ( .A(n13475), .B(n13474), .Z(n13477) );
  XNOR U12816 ( .A(n13472), .B(n13471), .Z(n13474) );
  XNOR U12817 ( .A(n13469), .B(n13468), .Z(n13471) );
  XNOR U12818 ( .A(n13466), .B(n13465), .Z(n13468) );
  XNOR U12819 ( .A(n13463), .B(n13462), .Z(n13465) );
  XNOR U12820 ( .A(n13460), .B(n13459), .Z(n13462) );
  XNOR U12821 ( .A(n13457), .B(n13456), .Z(n13459) );
  XNOR U12822 ( .A(n13454), .B(n13453), .Z(n13456) );
  XNOR U12823 ( .A(n13451), .B(n13450), .Z(n13453) );
  XNOR U12824 ( .A(n13448), .B(n13447), .Z(n13450) );
  XNOR U12825 ( .A(n13445), .B(n13444), .Z(n13447) );
  XNOR U12826 ( .A(n13442), .B(n13441), .Z(n13444) );
  XNOR U12827 ( .A(n13439), .B(n13438), .Z(n13441) );
  XNOR U12828 ( .A(n13436), .B(n13435), .Z(n13438) );
  XNOR U12829 ( .A(n13433), .B(n13432), .Z(n13435) );
  XNOR U12830 ( .A(n13430), .B(n13429), .Z(n13432) );
  XNOR U12831 ( .A(n13427), .B(n13426), .Z(n13429) );
  XNOR U12832 ( .A(n13424), .B(n13423), .Z(n13426) );
  XNOR U12833 ( .A(n13421), .B(n13420), .Z(n13423) );
  XNOR U12834 ( .A(n13418), .B(n13417), .Z(n13420) );
  XNOR U12835 ( .A(n13415), .B(n13414), .Z(n13417) );
  XNOR U12836 ( .A(n13412), .B(n13411), .Z(n13414) );
  XNOR U12837 ( .A(n13409), .B(n13408), .Z(n13411) );
  XNOR U12838 ( .A(n13406), .B(n13405), .Z(n13408) );
  XNOR U12839 ( .A(n13403), .B(n13402), .Z(n13405) );
  XNOR U12840 ( .A(n13400), .B(n13399), .Z(n13402) );
  XNOR U12841 ( .A(n13397), .B(n13396), .Z(n13399) );
  XNOR U12842 ( .A(n13394), .B(n13393), .Z(n13396) );
  XNOR U12843 ( .A(n13391), .B(n13390), .Z(n13393) );
  XNOR U12844 ( .A(n13388), .B(n13387), .Z(n13390) );
  XNOR U12845 ( .A(n13385), .B(n13384), .Z(n13387) );
  XNOR U12846 ( .A(n13382), .B(n13381), .Z(n13384) );
  XNOR U12847 ( .A(n13379), .B(n13378), .Z(n13381) );
  XNOR U12848 ( .A(n13376), .B(n13375), .Z(n13378) );
  XNOR U12849 ( .A(n13373), .B(n13372), .Z(n13375) );
  XNOR U12850 ( .A(n13370), .B(n13369), .Z(n13372) );
  XNOR U12851 ( .A(n13367), .B(n13366), .Z(n13369) );
  XNOR U12852 ( .A(n13364), .B(n13363), .Z(n13366) );
  XNOR U12853 ( .A(n13361), .B(n13360), .Z(n13363) );
  XNOR U12854 ( .A(n13358), .B(n13357), .Z(n13360) );
  XNOR U12855 ( .A(n13355), .B(n13354), .Z(n13357) );
  XNOR U12856 ( .A(n13352), .B(n13351), .Z(n13354) );
  XNOR U12857 ( .A(n13349), .B(n13348), .Z(n13351) );
  XNOR U12858 ( .A(n13346), .B(n13345), .Z(n13348) );
  XNOR U12859 ( .A(n13343), .B(n13342), .Z(n13345) );
  XNOR U12860 ( .A(n13340), .B(n13339), .Z(n13342) );
  XNOR U12861 ( .A(n13337), .B(n13336), .Z(n13339) );
  XNOR U12862 ( .A(n13334), .B(n13333), .Z(n13336) );
  XNOR U12863 ( .A(n13331), .B(n13330), .Z(n13333) );
  XNOR U12864 ( .A(n13328), .B(n13327), .Z(n13330) );
  XNOR U12865 ( .A(n13325), .B(n13324), .Z(n13327) );
  XNOR U12866 ( .A(n13322), .B(n13321), .Z(n13324) );
  XNOR U12867 ( .A(n13319), .B(n13318), .Z(n13321) );
  XNOR U12868 ( .A(n13316), .B(n13315), .Z(n13318) );
  XNOR U12869 ( .A(n13313), .B(n13312), .Z(n13315) );
  XNOR U12870 ( .A(n13310), .B(n13309), .Z(n13312) );
  XNOR U12871 ( .A(n13307), .B(n13306), .Z(n13309) );
  XNOR U12872 ( .A(n13304), .B(n13303), .Z(n13306) );
  XNOR U12873 ( .A(n13301), .B(n13300), .Z(n13303) );
  XNOR U12874 ( .A(n13298), .B(n13297), .Z(n13300) );
  XNOR U12875 ( .A(n13295), .B(n13294), .Z(n13297) );
  XNOR U12876 ( .A(n13292), .B(n13291), .Z(n13294) );
  XNOR U12877 ( .A(n13289), .B(n13288), .Z(n13291) );
  XNOR U12878 ( .A(n13286), .B(n13285), .Z(n13288) );
  XNOR U12879 ( .A(n13283), .B(n13282), .Z(n13285) );
  XNOR U12880 ( .A(n13280), .B(n13279), .Z(n13282) );
  XNOR U12881 ( .A(n13277), .B(n13276), .Z(n13279) );
  XNOR U12882 ( .A(n13274), .B(n13273), .Z(n13276) );
  XNOR U12883 ( .A(n13271), .B(n13270), .Z(n13273) );
  XNOR U12884 ( .A(n13268), .B(n13267), .Z(n13270) );
  XNOR U12885 ( .A(n13265), .B(n13264), .Z(n13267) );
  XNOR U12886 ( .A(n13262), .B(n13261), .Z(n13264) );
  XNOR U12887 ( .A(n13259), .B(n13258), .Z(n13261) );
  XNOR U12888 ( .A(n13256), .B(n13255), .Z(n13258) );
  XNOR U12889 ( .A(n13253), .B(n13252), .Z(n13255) );
  XNOR U12890 ( .A(n13250), .B(n13249), .Z(n13252) );
  XNOR U12891 ( .A(n13247), .B(n13246), .Z(n13249) );
  XNOR U12892 ( .A(n13244), .B(n13243), .Z(n13246) );
  XNOR U12893 ( .A(n13241), .B(n13240), .Z(n13243) );
  XNOR U12894 ( .A(n13238), .B(n13237), .Z(n13240) );
  XNOR U12895 ( .A(n13235), .B(n13234), .Z(n13237) );
  XNOR U12896 ( .A(n13232), .B(n13231), .Z(n13234) );
  XNOR U12897 ( .A(n13229), .B(n13228), .Z(n13231) );
  XNOR U12898 ( .A(n13226), .B(n13225), .Z(n13228) );
  XNOR U12899 ( .A(n13223), .B(n13222), .Z(n13225) );
  XNOR U12900 ( .A(n13220), .B(n13219), .Z(n13222) );
  XNOR U12901 ( .A(n13217), .B(n13216), .Z(n13219) );
  XNOR U12902 ( .A(n13214), .B(n13213), .Z(n13216) );
  XNOR U12903 ( .A(n13211), .B(n13210), .Z(n13213) );
  XNOR U12904 ( .A(n13208), .B(n13207), .Z(n13210) );
  XNOR U12905 ( .A(n13205), .B(n13204), .Z(n13207) );
  XNOR U12906 ( .A(n13202), .B(n13201), .Z(n13204) );
  XNOR U12907 ( .A(n13199), .B(n13198), .Z(n13201) );
  XNOR U12908 ( .A(n13196), .B(n13195), .Z(n13198) );
  XNOR U12909 ( .A(n13193), .B(n13192), .Z(n13195) );
  XNOR U12910 ( .A(n13190), .B(n13189), .Z(n13192) );
  XNOR U12911 ( .A(n13187), .B(n13186), .Z(n13189) );
  XNOR U12912 ( .A(n13184), .B(n13183), .Z(n13186) );
  XNOR U12913 ( .A(n13181), .B(n13180), .Z(n13183) );
  XNOR U12914 ( .A(n13178), .B(n13177), .Z(n13180) );
  XNOR U12915 ( .A(n13175), .B(n13174), .Z(n13177) );
  XNOR U12916 ( .A(n13172), .B(n13171), .Z(n13174) );
  XNOR U12917 ( .A(n13169), .B(n13168), .Z(n13171) );
  XNOR U12918 ( .A(n13166), .B(n13165), .Z(n13168) );
  XNOR U12919 ( .A(n13163), .B(n13162), .Z(n13165) );
  XNOR U12920 ( .A(n13160), .B(n13159), .Z(n13162) );
  XNOR U12921 ( .A(n13157), .B(n13156), .Z(n13159) );
  XNOR U12922 ( .A(n13154), .B(n13153), .Z(n13156) );
  XNOR U12923 ( .A(n13151), .B(n13150), .Z(n13153) );
  XNOR U12924 ( .A(n13148), .B(n13147), .Z(n13150) );
  XNOR U12925 ( .A(n13145), .B(n13144), .Z(n13147) );
  XOR U12926 ( .A(n14217), .B(n13141), .Z(n13144) );
  XOR U12927 ( .A(n13139), .B(n13138), .Z(n13141) );
  XOR U12928 ( .A(n13136), .B(n13135), .Z(n13138) );
  XOR U12929 ( .A(n13132), .B(n13133), .Z(n13135) );
  AND U12930 ( .A(n14218), .B(n14219), .Z(n13133) );
  XOR U12931 ( .A(n13129), .B(n13130), .Z(n13132) );
  AND U12932 ( .A(n14220), .B(n14221), .Z(n13130) );
  XOR U12933 ( .A(n13126), .B(n13127), .Z(n13129) );
  AND U12934 ( .A(n14222), .B(n14223), .Z(n13127) );
  XOR U12935 ( .A(n13123), .B(n13124), .Z(n13126) );
  AND U12936 ( .A(n14224), .B(n14225), .Z(n13124) );
  XNOR U12937 ( .A(n12906), .B(n13121), .Z(n13123) );
  AND U12938 ( .A(n14226), .B(n14227), .Z(n13121) );
  XOR U12939 ( .A(n12908), .B(n12907), .Z(n12906) );
  AND U12940 ( .A(n14228), .B(n14229), .Z(n12907) );
  XOR U12941 ( .A(n12910), .B(n12909), .Z(n12908) );
  AND U12942 ( .A(n14230), .B(n14231), .Z(n12909) );
  XOR U12943 ( .A(n12912), .B(n12911), .Z(n12910) );
  AND U12944 ( .A(n14232), .B(n14233), .Z(n12911) );
  XOR U12945 ( .A(n12914), .B(n12913), .Z(n12912) );
  AND U12946 ( .A(n14234), .B(n14235), .Z(n12913) );
  XOR U12947 ( .A(n12916), .B(n12915), .Z(n12914) );
  AND U12948 ( .A(n14236), .B(n14237), .Z(n12915) );
  XOR U12949 ( .A(n12918), .B(n12917), .Z(n12916) );
  AND U12950 ( .A(n14238), .B(n14239), .Z(n12917) );
  XOR U12951 ( .A(n12920), .B(n12919), .Z(n12918) );
  AND U12952 ( .A(n14240), .B(n14241), .Z(n12919) );
  XOR U12953 ( .A(n12922), .B(n12921), .Z(n12920) );
  AND U12954 ( .A(n14242), .B(n14243), .Z(n12921) );
  XOR U12955 ( .A(n12924), .B(n12923), .Z(n12922) );
  AND U12956 ( .A(n14244), .B(n14245), .Z(n12923) );
  XOR U12957 ( .A(n12926), .B(n12925), .Z(n12924) );
  AND U12958 ( .A(n14246), .B(n14247), .Z(n12925) );
  XOR U12959 ( .A(n12928), .B(n12927), .Z(n12926) );
  AND U12960 ( .A(n14248), .B(n14249), .Z(n12927) );
  XOR U12961 ( .A(n12930), .B(n12929), .Z(n12928) );
  AND U12962 ( .A(n14250), .B(n14251), .Z(n12929) );
  XOR U12963 ( .A(n12932), .B(n12931), .Z(n12930) );
  AND U12964 ( .A(n14252), .B(n14253), .Z(n12931) );
  XOR U12965 ( .A(n12934), .B(n12933), .Z(n12932) );
  AND U12966 ( .A(n14254), .B(n14255), .Z(n12933) );
  XOR U12967 ( .A(n12936), .B(n12935), .Z(n12934) );
  AND U12968 ( .A(n14256), .B(n14257), .Z(n12935) );
  XOR U12969 ( .A(n12938), .B(n12937), .Z(n12936) );
  AND U12970 ( .A(n14258), .B(n14259), .Z(n12937) );
  XOR U12971 ( .A(n12940), .B(n12939), .Z(n12938) );
  AND U12972 ( .A(n14260), .B(n14261), .Z(n12939) );
  XOR U12973 ( .A(n12942), .B(n12941), .Z(n12940) );
  AND U12974 ( .A(n14262), .B(n14263), .Z(n12941) );
  XOR U12975 ( .A(n12944), .B(n12943), .Z(n12942) );
  AND U12976 ( .A(n14264), .B(n14265), .Z(n12943) );
  XOR U12977 ( .A(n12946), .B(n12945), .Z(n12944) );
  AND U12978 ( .A(n14266), .B(n14267), .Z(n12945) );
  XOR U12979 ( .A(n12948), .B(n12947), .Z(n12946) );
  AND U12980 ( .A(n14268), .B(n14269), .Z(n12947) );
  XOR U12981 ( .A(n12950), .B(n12949), .Z(n12948) );
  AND U12982 ( .A(n14270), .B(n14271), .Z(n12949) );
  XOR U12983 ( .A(n12952), .B(n12951), .Z(n12950) );
  AND U12984 ( .A(n14272), .B(n14273), .Z(n12951) );
  XOR U12985 ( .A(n12954), .B(n12953), .Z(n12952) );
  AND U12986 ( .A(n14274), .B(n14275), .Z(n12953) );
  XOR U12987 ( .A(n12956), .B(n12955), .Z(n12954) );
  AND U12988 ( .A(n14276), .B(n14277), .Z(n12955) );
  XOR U12989 ( .A(n12958), .B(n12957), .Z(n12956) );
  AND U12990 ( .A(n14278), .B(n14279), .Z(n12957) );
  XOR U12991 ( .A(n12960), .B(n12959), .Z(n12958) );
  AND U12992 ( .A(n14280), .B(n14281), .Z(n12959) );
  XOR U12993 ( .A(n12962), .B(n12961), .Z(n12960) );
  AND U12994 ( .A(n14282), .B(n14283), .Z(n12961) );
  XOR U12995 ( .A(n12964), .B(n12963), .Z(n12962) );
  AND U12996 ( .A(n14284), .B(n14285), .Z(n12963) );
  XOR U12997 ( .A(n12966), .B(n12965), .Z(n12964) );
  AND U12998 ( .A(n14286), .B(n14287), .Z(n12965) );
  XOR U12999 ( .A(n12968), .B(n12967), .Z(n12966) );
  AND U13000 ( .A(n14288), .B(n14289), .Z(n12967) );
  XOR U13001 ( .A(n12970), .B(n12969), .Z(n12968) );
  AND U13002 ( .A(n14290), .B(n14291), .Z(n12969) );
  XOR U13003 ( .A(n12972), .B(n12971), .Z(n12970) );
  AND U13004 ( .A(n14292), .B(n14293), .Z(n12971) );
  XOR U13005 ( .A(n12974), .B(n12973), .Z(n12972) );
  AND U13006 ( .A(n14294), .B(n14295), .Z(n12973) );
  XOR U13007 ( .A(n12976), .B(n12975), .Z(n12974) );
  AND U13008 ( .A(n14296), .B(n14297), .Z(n12975) );
  XOR U13009 ( .A(n12978), .B(n12977), .Z(n12976) );
  AND U13010 ( .A(n14298), .B(n14299), .Z(n12977) );
  XOR U13011 ( .A(n12980), .B(n12979), .Z(n12978) );
  AND U13012 ( .A(n14300), .B(n14301), .Z(n12979) );
  XOR U13013 ( .A(n12982), .B(n12981), .Z(n12980) );
  AND U13014 ( .A(n14302), .B(n14303), .Z(n12981) );
  XOR U13015 ( .A(n12984), .B(n12983), .Z(n12982) );
  AND U13016 ( .A(n14304), .B(n14305), .Z(n12983) );
  XOR U13017 ( .A(n13117), .B(n12985), .Z(n12984) );
  AND U13018 ( .A(n14306), .B(n14307), .Z(n12985) );
  XOR U13019 ( .A(n13119), .B(n13118), .Z(n13117) );
  AND U13020 ( .A(n14308), .B(n14309), .Z(n13118) );
  XOR U13021 ( .A(n13101), .B(n13120), .Z(n13119) );
  AND U13022 ( .A(n14310), .B(n14311), .Z(n13120) );
  XOR U13023 ( .A(n13103), .B(n13102), .Z(n13101) );
  AND U13024 ( .A(n14312), .B(n14313), .Z(n13102) );
  XOR U13025 ( .A(n13105), .B(n13104), .Z(n13103) );
  AND U13026 ( .A(n14314), .B(n14315), .Z(n13104) );
  XOR U13027 ( .A(n13109), .B(n13106), .Z(n13105) );
  AND U13028 ( .A(n14316), .B(n14317), .Z(n13106) );
  XOR U13029 ( .A(n13111), .B(n13110), .Z(n13109) );
  AND U13030 ( .A(n14318), .B(n14319), .Z(n13110) );
  XOR U13031 ( .A(n13113), .B(n13112), .Z(n13111) );
  AND U13032 ( .A(n14320), .B(n14321), .Z(n13112) );
  XOR U13033 ( .A(n13115), .B(n13114), .Z(n13113) );
  AND U13034 ( .A(n14322), .B(n14323), .Z(n13114) );
  XOR U13035 ( .A(n13099), .B(n13116), .Z(n13115) );
  AND U13036 ( .A(n14324), .B(n14325), .Z(n13116) );
  XNOR U13037 ( .A(n13008), .B(n13100), .Z(n13099) );
  AND U13038 ( .A(n14326), .B(n14327), .Z(n13100) );
  XOR U13039 ( .A(n13007), .B(n12999), .Z(n13008) );
  AND U13040 ( .A(n14328), .B(n14329), .Z(n12999) );
  XNOR U13041 ( .A(n13002), .B(n12998), .Z(n13007) );
  AND U13042 ( .A(n14330), .B(n14331), .Z(n12998) );
  XOR U13043 ( .A(n13028), .B(n13003), .Z(n13002) );
  AND U13044 ( .A(n14332), .B(n14333), .Z(n13003) );
  XNOR U13045 ( .A(n13019), .B(n13029), .Z(n13028) );
  AND U13046 ( .A(n14334), .B(n14335), .Z(n13029) );
  XOR U13047 ( .A(n13017), .B(n13018), .Z(n13019) );
  AND U13048 ( .A(n14336), .B(n14337), .Z(n13018) );
  XNOR U13049 ( .A(n13011), .B(n13016), .Z(n13017) );
  AND U13050 ( .A(n14338), .B(n14339), .Z(n13016) );
  XOR U13051 ( .A(n13030), .B(n13012), .Z(n13011) );
  AND U13052 ( .A(n14340), .B(n14341), .Z(n13012) );
  XNOR U13053 ( .A(n13096), .B(n13031), .Z(n13030) );
  AND U13054 ( .A(n14342), .B(n14343), .Z(n13031) );
  XOR U13055 ( .A(n13095), .B(n13087), .Z(n13096) );
  AND U13056 ( .A(n14344), .B(n14345), .Z(n13087) );
  XNOR U13057 ( .A(n13090), .B(n13086), .Z(n13095) );
  AND U13058 ( .A(n14346), .B(n14347), .Z(n13086) );
  XOR U13059 ( .A(n13034), .B(n13091), .Z(n13090) );
  AND U13060 ( .A(n14348), .B(n14349), .Z(n13091) );
  XNOR U13061 ( .A(n13083), .B(n13035), .Z(n13034) );
  AND U13062 ( .A(n14350), .B(n14351), .Z(n13035) );
  XOR U13063 ( .A(n13082), .B(n13074), .Z(n13083) );
  AND U13064 ( .A(n14352), .B(n14353), .Z(n13074) );
  XNOR U13065 ( .A(n13077), .B(n13073), .Z(n13082) );
  AND U13066 ( .A(n14354), .B(n14355), .Z(n13073) );
  XOR U13067 ( .A(n14356), .B(n14357), .Z(n13077) );
  XOR U13068 ( .A(n13067), .B(n13068), .Z(n14357) );
  AND U13069 ( .A(n14358), .B(n14359), .Z(n13068) );
  AND U13070 ( .A(n14360), .B(n14361), .Z(n13067) );
  XOR U13071 ( .A(n14362), .B(n13078), .Z(n14356) );
  AND U13072 ( .A(n14363), .B(n14364), .Z(n13078) );
  XOR U13073 ( .A(n14365), .B(n14366), .Z(n14362) );
  XOR U13074 ( .A(n14367), .B(n14368), .Z(n14366) );
  XOR U13075 ( .A(n13060), .B(n13061), .Z(n14368) );
  AND U13076 ( .A(n14369), .B(n14370), .Z(n13061) );
  AND U13077 ( .A(n14371), .B(n14372), .Z(n13060) );
  XOR U13078 ( .A(n13054), .B(n13059), .Z(n14367) );
  AND U13079 ( .A(n14373), .B(n14374), .Z(n13059) );
  AND U13080 ( .A(n14375), .B(n14376), .Z(n13054) );
  XOR U13081 ( .A(n14377), .B(n14378), .Z(n14365) );
  XOR U13082 ( .A(n13062), .B(n13065), .Z(n14378) );
  AND U13083 ( .A(n14379), .B(n14380), .Z(n13065) );
  AND U13084 ( .A(n14381), .B(n14382), .Z(n13062) );
  XOR U13085 ( .A(n14383), .B(n13066), .Z(n14377) );
  AND U13086 ( .A(n14384), .B(n14385), .Z(n13066) );
  XOR U13087 ( .A(n14386), .B(n14387), .Z(n14383) );
  XOR U13088 ( .A(n14388), .B(n14389), .Z(n14387) );
  XOR U13089 ( .A(n13047), .B(n13048), .Z(n14389) );
  AND U13090 ( .A(n14390), .B(n14391), .Z(n13048) );
  AND U13091 ( .A(n14392), .B(n14393), .Z(n13047) );
  XOR U13092 ( .A(n13045), .B(n13043), .Z(n14388) );
  AND U13093 ( .A(n14394), .B(n14395), .Z(n13043) );
  AND U13094 ( .A(n14396), .B(n14397), .Z(n13045) );
  XOR U13095 ( .A(n14398), .B(n14399), .Z(n14386) );
  XOR U13096 ( .A(n13051), .B(n13052), .Z(n14399) );
  AND U13097 ( .A(n14400), .B(n14401), .Z(n13052) );
  AND U13098 ( .A(n14402), .B(n14403), .Z(n13051) );
  XOR U13099 ( .A(n13046), .B(n13053), .Z(n14398) );
  AND U13100 ( .A(n14404), .B(n14405), .Z(n13053) );
  XOR U13101 ( .A(n14406), .B(n14407), .Z(n13046) );
  XOR U13102 ( .A(n14408), .B(n14409), .Z(n14407) );
  XOR U13103 ( .A(n14410), .B(n14411), .Z(n14409) );
  NOR U13104 ( .A(n14412), .B(n14413), .Z(n14411) );
  NOR U13105 ( .A(n14414), .B(n14415), .Z(n14410) );
  AND U13106 ( .A(n14416), .B(n14417), .Z(n14415) );
  IV U13107 ( .A(n14418), .Z(n14414) );
  NOR U13108 ( .A(n14419), .B(n14420), .Z(n14418) );
  AND U13109 ( .A(n14412), .B(n14421), .Z(n14420) );
  AND U13110 ( .A(n14413), .B(n14422), .Z(n14419) );
  XOR U13111 ( .A(n14423), .B(n14424), .Z(n14408) );
  NOR U13112 ( .A(n14425), .B(n14426), .Z(n14424) );
  NOR U13113 ( .A(n14427), .B(n14428), .Z(n14423) );
  AND U13114 ( .A(n14429), .B(n14430), .Z(n14428) );
  IV U13115 ( .A(n14431), .Z(n14427) );
  NOR U13116 ( .A(n14432), .B(n14433), .Z(n14431) );
  AND U13117 ( .A(n14425), .B(n14434), .Z(n14433) );
  AND U13118 ( .A(n14426), .B(n14435), .Z(n14432) );
  XOR U13119 ( .A(n14436), .B(n14437), .Z(n14406) );
  AND U13120 ( .A(n14438), .B(n14439), .Z(n14437) );
  XNOR U13121 ( .A(n14440), .B(n14441), .Z(n14436) );
  AND U13122 ( .A(n14442), .B(n14443), .Z(n14441) );
  AND U13123 ( .A(n14444), .B(n14445), .Z(n14440) );
  AND U13124 ( .A(n14446), .B(n14447), .Z(n14445) );
  NOR U13125 ( .A(n14448), .B(n14449), .Z(n14447) );
  IV U13126 ( .A(n14450), .Z(n14448) );
  NOR U13127 ( .A(n14451), .B(n14452), .Z(n14450) );
  NOR U13128 ( .A(n14453), .B(n14454), .Z(n14446) );
  AND U13129 ( .A(n14455), .B(n14456), .Z(n14444) );
  NOR U13130 ( .A(n14457), .B(n14458), .Z(n14456) );
  NOR U13131 ( .A(n14459), .B(n14460), .Z(n14455) );
  XOR U13132 ( .A(n14461), .B(n14462), .Z(n13136) );
  AND U13133 ( .A(n14461), .B(n14463), .Z(n14462) );
  XNOR U13134 ( .A(n14464), .B(n14465), .Z(n13139) );
  AND U13135 ( .A(n14464), .B(n14466), .Z(n14465) );
  IV U13136 ( .A(n13142), .Z(n14217) );
  XNOR U13137 ( .A(n14467), .B(n14468), .Z(n13142) );
  AND U13138 ( .A(n14467), .B(n14469), .Z(n14468) );
  XNOR U13139 ( .A(n14470), .B(n14471), .Z(n13145) );
  AND U13140 ( .A(n14470), .B(n14472), .Z(n14471) );
  XNOR U13141 ( .A(n14473), .B(n14474), .Z(n13148) );
  AND U13142 ( .A(n14475), .B(n14473), .Z(n14474) );
  XOR U13143 ( .A(n14476), .B(n14477), .Z(n13151) );
  NOR U13144 ( .A(n14478), .B(n14476), .Z(n14477) );
  XOR U13145 ( .A(n14479), .B(n14480), .Z(n13154) );
  NOR U13146 ( .A(n14481), .B(n14479), .Z(n14480) );
  XOR U13147 ( .A(n14482), .B(n14483), .Z(n13157) );
  NOR U13148 ( .A(n14484), .B(n14482), .Z(n14483) );
  XOR U13149 ( .A(n14485), .B(n14486), .Z(n13160) );
  NOR U13150 ( .A(n14487), .B(n14485), .Z(n14486) );
  XOR U13151 ( .A(n14488), .B(n14489), .Z(n13163) );
  NOR U13152 ( .A(n14490), .B(n14488), .Z(n14489) );
  XOR U13153 ( .A(n14491), .B(n14492), .Z(n13166) );
  NOR U13154 ( .A(n14493), .B(n14491), .Z(n14492) );
  XOR U13155 ( .A(n14494), .B(n14495), .Z(n13169) );
  NOR U13156 ( .A(n14496), .B(n14494), .Z(n14495) );
  XOR U13157 ( .A(n14497), .B(n14498), .Z(n13172) );
  NOR U13158 ( .A(n14499), .B(n14497), .Z(n14498) );
  XOR U13159 ( .A(n14500), .B(n14501), .Z(n13175) );
  NOR U13160 ( .A(n14502), .B(n14500), .Z(n14501) );
  XOR U13161 ( .A(n14503), .B(n14504), .Z(n13178) );
  NOR U13162 ( .A(n14505), .B(n14503), .Z(n14504) );
  XOR U13163 ( .A(n14506), .B(n14507), .Z(n13181) );
  NOR U13164 ( .A(n14508), .B(n14506), .Z(n14507) );
  XOR U13165 ( .A(n14509), .B(n14510), .Z(n13184) );
  NOR U13166 ( .A(n14511), .B(n14509), .Z(n14510) );
  XOR U13167 ( .A(n14512), .B(n14513), .Z(n13187) );
  NOR U13168 ( .A(n14514), .B(n14512), .Z(n14513) );
  XOR U13169 ( .A(n14515), .B(n14516), .Z(n13190) );
  NOR U13170 ( .A(n14517), .B(n14515), .Z(n14516) );
  XOR U13171 ( .A(n14518), .B(n14519), .Z(n13193) );
  NOR U13172 ( .A(n14520), .B(n14518), .Z(n14519) );
  XOR U13173 ( .A(n14521), .B(n14522), .Z(n13196) );
  NOR U13174 ( .A(n14523), .B(n14521), .Z(n14522) );
  XOR U13175 ( .A(n14524), .B(n14525), .Z(n13199) );
  NOR U13176 ( .A(n14526), .B(n14524), .Z(n14525) );
  XOR U13177 ( .A(n14527), .B(n14528), .Z(n13202) );
  NOR U13178 ( .A(n14529), .B(n14527), .Z(n14528) );
  XOR U13179 ( .A(n14530), .B(n14531), .Z(n13205) );
  NOR U13180 ( .A(n14532), .B(n14530), .Z(n14531) );
  XOR U13181 ( .A(n14533), .B(n14534), .Z(n13208) );
  NOR U13182 ( .A(n14535), .B(n14533), .Z(n14534) );
  XOR U13183 ( .A(n14536), .B(n14537), .Z(n13211) );
  NOR U13184 ( .A(n14538), .B(n14536), .Z(n14537) );
  XOR U13185 ( .A(n14539), .B(n14540), .Z(n13214) );
  NOR U13186 ( .A(n14541), .B(n14539), .Z(n14540) );
  XOR U13187 ( .A(n14542), .B(n14543), .Z(n13217) );
  NOR U13188 ( .A(n14544), .B(n14542), .Z(n14543) );
  XOR U13189 ( .A(n14545), .B(n14546), .Z(n13220) );
  NOR U13190 ( .A(n14547), .B(n14545), .Z(n14546) );
  XOR U13191 ( .A(n14548), .B(n14549), .Z(n13223) );
  NOR U13192 ( .A(n14550), .B(n14548), .Z(n14549) );
  XOR U13193 ( .A(n14551), .B(n14552), .Z(n13226) );
  NOR U13194 ( .A(n14553), .B(n14551), .Z(n14552) );
  XOR U13195 ( .A(n14554), .B(n14555), .Z(n13229) );
  NOR U13196 ( .A(n14556), .B(n14554), .Z(n14555) );
  XOR U13197 ( .A(n14557), .B(n14558), .Z(n13232) );
  NOR U13198 ( .A(n14559), .B(n14557), .Z(n14558) );
  XOR U13199 ( .A(n14560), .B(n14561), .Z(n13235) );
  NOR U13200 ( .A(n14562), .B(n14560), .Z(n14561) );
  XOR U13201 ( .A(n14563), .B(n14564), .Z(n13238) );
  NOR U13202 ( .A(n14565), .B(n14563), .Z(n14564) );
  XOR U13203 ( .A(n14566), .B(n14567), .Z(n13241) );
  NOR U13204 ( .A(n14568), .B(n14566), .Z(n14567) );
  XOR U13205 ( .A(n14569), .B(n14570), .Z(n13244) );
  NOR U13206 ( .A(n14571), .B(n14569), .Z(n14570) );
  XOR U13207 ( .A(n14572), .B(n14573), .Z(n13247) );
  NOR U13208 ( .A(n14574), .B(n14572), .Z(n14573) );
  XOR U13209 ( .A(n14575), .B(n14576), .Z(n13250) );
  NOR U13210 ( .A(n14577), .B(n14575), .Z(n14576) );
  XOR U13211 ( .A(n14578), .B(n14579), .Z(n13253) );
  NOR U13212 ( .A(n14580), .B(n14578), .Z(n14579) );
  XOR U13213 ( .A(n14581), .B(n14582), .Z(n13256) );
  NOR U13214 ( .A(n14583), .B(n14581), .Z(n14582) );
  XOR U13215 ( .A(n14584), .B(n14585), .Z(n13259) );
  NOR U13216 ( .A(n14586), .B(n14584), .Z(n14585) );
  XOR U13217 ( .A(n14587), .B(n14588), .Z(n13262) );
  NOR U13218 ( .A(n14589), .B(n14587), .Z(n14588) );
  XOR U13219 ( .A(n14590), .B(n14591), .Z(n13265) );
  NOR U13220 ( .A(n14592), .B(n14590), .Z(n14591) );
  XOR U13221 ( .A(n14593), .B(n14594), .Z(n13268) );
  NOR U13222 ( .A(n14595), .B(n14593), .Z(n14594) );
  XOR U13223 ( .A(n14596), .B(n14597), .Z(n13271) );
  NOR U13224 ( .A(n14598), .B(n14596), .Z(n14597) );
  XOR U13225 ( .A(n14599), .B(n14600), .Z(n13274) );
  NOR U13226 ( .A(n14601), .B(n14599), .Z(n14600) );
  XOR U13227 ( .A(n14602), .B(n14603), .Z(n13277) );
  NOR U13228 ( .A(n14604), .B(n14602), .Z(n14603) );
  XOR U13229 ( .A(n14605), .B(n14606), .Z(n13280) );
  NOR U13230 ( .A(n14607), .B(n14605), .Z(n14606) );
  XOR U13231 ( .A(n14608), .B(n14609), .Z(n13283) );
  NOR U13232 ( .A(n14610), .B(n14608), .Z(n14609) );
  XOR U13233 ( .A(n14611), .B(n14612), .Z(n13286) );
  NOR U13234 ( .A(n14613), .B(n14611), .Z(n14612) );
  XOR U13235 ( .A(n14614), .B(n14615), .Z(n13289) );
  NOR U13236 ( .A(n14616), .B(n14614), .Z(n14615) );
  XOR U13237 ( .A(n14617), .B(n14618), .Z(n13292) );
  NOR U13238 ( .A(n14619), .B(n14617), .Z(n14618) );
  XOR U13239 ( .A(n14620), .B(n14621), .Z(n13295) );
  NOR U13240 ( .A(n14622), .B(n14620), .Z(n14621) );
  XOR U13241 ( .A(n14623), .B(n14624), .Z(n13298) );
  NOR U13242 ( .A(n14625), .B(n14623), .Z(n14624) );
  XOR U13243 ( .A(n14626), .B(n14627), .Z(n13301) );
  NOR U13244 ( .A(n14628), .B(n14626), .Z(n14627) );
  XOR U13245 ( .A(n14629), .B(n14630), .Z(n13304) );
  NOR U13246 ( .A(n14631), .B(n14629), .Z(n14630) );
  XOR U13247 ( .A(n14632), .B(n14633), .Z(n13307) );
  NOR U13248 ( .A(n14634), .B(n14632), .Z(n14633) );
  XOR U13249 ( .A(n14635), .B(n14636), .Z(n13310) );
  NOR U13250 ( .A(n14637), .B(n14635), .Z(n14636) );
  XOR U13251 ( .A(n14638), .B(n14639), .Z(n13313) );
  NOR U13252 ( .A(n14640), .B(n14638), .Z(n14639) );
  XOR U13253 ( .A(n14641), .B(n14642), .Z(n13316) );
  NOR U13254 ( .A(n14643), .B(n14641), .Z(n14642) );
  XOR U13255 ( .A(n14644), .B(n14645), .Z(n13319) );
  NOR U13256 ( .A(n14646), .B(n14644), .Z(n14645) );
  XOR U13257 ( .A(n14647), .B(n14648), .Z(n13322) );
  NOR U13258 ( .A(n14649), .B(n14647), .Z(n14648) );
  XOR U13259 ( .A(n14650), .B(n14651), .Z(n13325) );
  NOR U13260 ( .A(n14652), .B(n14650), .Z(n14651) );
  XOR U13261 ( .A(n14653), .B(n14654), .Z(n13328) );
  NOR U13262 ( .A(n14655), .B(n14653), .Z(n14654) );
  XOR U13263 ( .A(n14656), .B(n14657), .Z(n13331) );
  NOR U13264 ( .A(n14658), .B(n14656), .Z(n14657) );
  XOR U13265 ( .A(n14659), .B(n14660), .Z(n13334) );
  NOR U13266 ( .A(n14661), .B(n14659), .Z(n14660) );
  XOR U13267 ( .A(n14662), .B(n14663), .Z(n13337) );
  NOR U13268 ( .A(n14664), .B(n14662), .Z(n14663) );
  XOR U13269 ( .A(n14665), .B(n14666), .Z(n13340) );
  NOR U13270 ( .A(n14667), .B(n14665), .Z(n14666) );
  XOR U13271 ( .A(n14668), .B(n14669), .Z(n13343) );
  NOR U13272 ( .A(n14670), .B(n14668), .Z(n14669) );
  XOR U13273 ( .A(n14671), .B(n14672), .Z(n13346) );
  NOR U13274 ( .A(n14673), .B(n14671), .Z(n14672) );
  XOR U13275 ( .A(n14674), .B(n14675), .Z(n13349) );
  NOR U13276 ( .A(n14676), .B(n14674), .Z(n14675) );
  XOR U13277 ( .A(n14677), .B(n14678), .Z(n13352) );
  NOR U13278 ( .A(n14679), .B(n14677), .Z(n14678) );
  XOR U13279 ( .A(n14680), .B(n14681), .Z(n13355) );
  NOR U13280 ( .A(n14682), .B(n14680), .Z(n14681) );
  XOR U13281 ( .A(n14683), .B(n14684), .Z(n13358) );
  NOR U13282 ( .A(n14685), .B(n14683), .Z(n14684) );
  XOR U13283 ( .A(n14686), .B(n14687), .Z(n13361) );
  NOR U13284 ( .A(n14688), .B(n14686), .Z(n14687) );
  XOR U13285 ( .A(n14689), .B(n14690), .Z(n13364) );
  NOR U13286 ( .A(n14691), .B(n14689), .Z(n14690) );
  XOR U13287 ( .A(n14692), .B(n14693), .Z(n13367) );
  NOR U13288 ( .A(n14694), .B(n14692), .Z(n14693) );
  XOR U13289 ( .A(n14695), .B(n14696), .Z(n13370) );
  NOR U13290 ( .A(n14697), .B(n14695), .Z(n14696) );
  XOR U13291 ( .A(n14698), .B(n14699), .Z(n13373) );
  NOR U13292 ( .A(n14700), .B(n14698), .Z(n14699) );
  XOR U13293 ( .A(n14701), .B(n14702), .Z(n13376) );
  NOR U13294 ( .A(n14703), .B(n14701), .Z(n14702) );
  XOR U13295 ( .A(n14704), .B(n14705), .Z(n13379) );
  NOR U13296 ( .A(n14706), .B(n14704), .Z(n14705) );
  XOR U13297 ( .A(n14707), .B(n14708), .Z(n13382) );
  NOR U13298 ( .A(n14709), .B(n14707), .Z(n14708) );
  XOR U13299 ( .A(n14710), .B(n14711), .Z(n13385) );
  NOR U13300 ( .A(n14712), .B(n14710), .Z(n14711) );
  XOR U13301 ( .A(n14713), .B(n14714), .Z(n13388) );
  NOR U13302 ( .A(n14715), .B(n14713), .Z(n14714) );
  XOR U13303 ( .A(n14716), .B(n14717), .Z(n13391) );
  NOR U13304 ( .A(n14718), .B(n14716), .Z(n14717) );
  XOR U13305 ( .A(n14719), .B(n14720), .Z(n13394) );
  NOR U13306 ( .A(n14721), .B(n14719), .Z(n14720) );
  XOR U13307 ( .A(n14722), .B(n14723), .Z(n13397) );
  NOR U13308 ( .A(n14724), .B(n14722), .Z(n14723) );
  XOR U13309 ( .A(n14725), .B(n14726), .Z(n13400) );
  NOR U13310 ( .A(n14727), .B(n14725), .Z(n14726) );
  XOR U13311 ( .A(n14728), .B(n14729), .Z(n13403) );
  NOR U13312 ( .A(n14730), .B(n14728), .Z(n14729) );
  XOR U13313 ( .A(n14731), .B(n14732), .Z(n13406) );
  NOR U13314 ( .A(n14733), .B(n14731), .Z(n14732) );
  XOR U13315 ( .A(n14734), .B(n14735), .Z(n13409) );
  NOR U13316 ( .A(n14736), .B(n14734), .Z(n14735) );
  XOR U13317 ( .A(n14737), .B(n14738), .Z(n13412) );
  NOR U13318 ( .A(n14739), .B(n14737), .Z(n14738) );
  XOR U13319 ( .A(n14740), .B(n14741), .Z(n13415) );
  NOR U13320 ( .A(n14742), .B(n14740), .Z(n14741) );
  XOR U13321 ( .A(n14743), .B(n14744), .Z(n13418) );
  NOR U13322 ( .A(n14745), .B(n14743), .Z(n14744) );
  XOR U13323 ( .A(n14746), .B(n14747), .Z(n13421) );
  NOR U13324 ( .A(n14748), .B(n14746), .Z(n14747) );
  XOR U13325 ( .A(n14749), .B(n14750), .Z(n13424) );
  NOR U13326 ( .A(n14751), .B(n14749), .Z(n14750) );
  XOR U13327 ( .A(n14752), .B(n14753), .Z(n13427) );
  NOR U13328 ( .A(n14754), .B(n14752), .Z(n14753) );
  XOR U13329 ( .A(n14755), .B(n14756), .Z(n13430) );
  NOR U13330 ( .A(n14757), .B(n14755), .Z(n14756) );
  XOR U13331 ( .A(n14758), .B(n14759), .Z(n13433) );
  NOR U13332 ( .A(n14760), .B(n14758), .Z(n14759) );
  XOR U13333 ( .A(n14761), .B(n14762), .Z(n13436) );
  NOR U13334 ( .A(n14763), .B(n14761), .Z(n14762) );
  XOR U13335 ( .A(n14764), .B(n14765), .Z(n13439) );
  NOR U13336 ( .A(n14766), .B(n14764), .Z(n14765) );
  XOR U13337 ( .A(n14767), .B(n14768), .Z(n13442) );
  NOR U13338 ( .A(n14769), .B(n14767), .Z(n14768) );
  XOR U13339 ( .A(n14770), .B(n14771), .Z(n13445) );
  NOR U13340 ( .A(n14772), .B(n14770), .Z(n14771) );
  XOR U13341 ( .A(n14773), .B(n14774), .Z(n13448) );
  NOR U13342 ( .A(n14775), .B(n14773), .Z(n14774) );
  XOR U13343 ( .A(n14776), .B(n14777), .Z(n13451) );
  NOR U13344 ( .A(n14778), .B(n14776), .Z(n14777) );
  XOR U13345 ( .A(n14779), .B(n14780), .Z(n13454) );
  NOR U13346 ( .A(n14781), .B(n14779), .Z(n14780) );
  XOR U13347 ( .A(n14782), .B(n14783), .Z(n13457) );
  NOR U13348 ( .A(n14784), .B(n14782), .Z(n14783) );
  XOR U13349 ( .A(n14785), .B(n14786), .Z(n13460) );
  NOR U13350 ( .A(n14787), .B(n14785), .Z(n14786) );
  XOR U13351 ( .A(n14788), .B(n14789), .Z(n13463) );
  NOR U13352 ( .A(n14790), .B(n14788), .Z(n14789) );
  XOR U13353 ( .A(n14791), .B(n14792), .Z(n13466) );
  NOR U13354 ( .A(n14793), .B(n14791), .Z(n14792) );
  XOR U13355 ( .A(n14794), .B(n14795), .Z(n13469) );
  NOR U13356 ( .A(n14796), .B(n14794), .Z(n14795) );
  XOR U13357 ( .A(n14797), .B(n14798), .Z(n13472) );
  NOR U13358 ( .A(n14799), .B(n14797), .Z(n14798) );
  XOR U13359 ( .A(n14800), .B(n14801), .Z(n13475) );
  NOR U13360 ( .A(n14802), .B(n14800), .Z(n14801) );
  XOR U13361 ( .A(n14803), .B(n14804), .Z(n13478) );
  NOR U13362 ( .A(n14805), .B(n14803), .Z(n14804) );
  XOR U13363 ( .A(n14806), .B(n14807), .Z(n13481) );
  NOR U13364 ( .A(n14808), .B(n14806), .Z(n14807) );
  XOR U13365 ( .A(n14809), .B(n14810), .Z(n13484) );
  NOR U13366 ( .A(n14811), .B(n14809), .Z(n14810) );
  XOR U13367 ( .A(n14812), .B(n14813), .Z(n13487) );
  NOR U13368 ( .A(n14814), .B(n14812), .Z(n14813) );
  XOR U13369 ( .A(n14815), .B(n14816), .Z(n13490) );
  NOR U13370 ( .A(n14817), .B(n14815), .Z(n14816) );
  XOR U13371 ( .A(n14818), .B(n14819), .Z(n13493) );
  NOR U13372 ( .A(n14820), .B(n14818), .Z(n14819) );
  XOR U13373 ( .A(n14821), .B(n14822), .Z(n13496) );
  NOR U13374 ( .A(n14823), .B(n14821), .Z(n14822) );
  XOR U13375 ( .A(n14824), .B(n14825), .Z(n13499) );
  NOR U13376 ( .A(n14826), .B(n14824), .Z(n14825) );
  XOR U13377 ( .A(n14827), .B(n14828), .Z(n13502) );
  NOR U13378 ( .A(n14829), .B(n14827), .Z(n14828) );
  XOR U13379 ( .A(n14830), .B(n14831), .Z(n13505) );
  NOR U13380 ( .A(n14832), .B(n14830), .Z(n14831) );
  XOR U13381 ( .A(n14833), .B(n14834), .Z(n13508) );
  NOR U13382 ( .A(n14835), .B(n14833), .Z(n14834) );
  XOR U13383 ( .A(n14836), .B(n14837), .Z(n13511) );
  NOR U13384 ( .A(n14838), .B(n14836), .Z(n14837) );
  XOR U13385 ( .A(n14839), .B(n14840), .Z(n13514) );
  NOR U13386 ( .A(n14841), .B(n14839), .Z(n14840) );
  XOR U13387 ( .A(n14842), .B(n14843), .Z(n13517) );
  NOR U13388 ( .A(n14844), .B(n14842), .Z(n14843) );
  XOR U13389 ( .A(n14845), .B(n14846), .Z(n13520) );
  NOR U13390 ( .A(n14847), .B(n14845), .Z(n14846) );
  XOR U13391 ( .A(n14848), .B(n14849), .Z(n13523) );
  NOR U13392 ( .A(n14850), .B(n14848), .Z(n14849) );
  XOR U13393 ( .A(n14851), .B(n14852), .Z(n13526) );
  NOR U13394 ( .A(n14853), .B(n14851), .Z(n14852) );
  XOR U13395 ( .A(n14854), .B(n14855), .Z(n13529) );
  NOR U13396 ( .A(n14856), .B(n14854), .Z(n14855) );
  XOR U13397 ( .A(n14857), .B(n14858), .Z(n13532) );
  NOR U13398 ( .A(n14859), .B(n14857), .Z(n14858) );
  XOR U13399 ( .A(n14860), .B(n14861), .Z(n13535) );
  NOR U13400 ( .A(n14862), .B(n14860), .Z(n14861) );
  XOR U13401 ( .A(n14863), .B(n14864), .Z(n13538) );
  NOR U13402 ( .A(n14865), .B(n14863), .Z(n14864) );
  XOR U13403 ( .A(n14866), .B(n14867), .Z(n13541) );
  NOR U13404 ( .A(n14868), .B(n14866), .Z(n14867) );
  XOR U13405 ( .A(n14869), .B(n14870), .Z(n13544) );
  NOR U13406 ( .A(n14871), .B(n14869), .Z(n14870) );
  XOR U13407 ( .A(n14872), .B(n14873), .Z(n13547) );
  NOR U13408 ( .A(n14874), .B(n14872), .Z(n14873) );
  XOR U13409 ( .A(n14875), .B(n14876), .Z(n13550) );
  NOR U13410 ( .A(n90), .B(n14877), .Z(n14876) );
  IV U13411 ( .A(n14875), .Z(n14877) );
  XOR U13412 ( .A(n14878), .B(n14879), .Z(n13553) );
  AND U13413 ( .A(n14880), .B(n14881), .Z(n14879) );
  XOR U13414 ( .A(n14878), .B(n93), .Z(n14881) );
  XOR U13415 ( .A(n14215), .B(n14214), .Z(n93) );
  XNOR U13416 ( .A(n14212), .B(n14211), .Z(n14214) );
  XNOR U13417 ( .A(n14209), .B(n14208), .Z(n14211) );
  XNOR U13418 ( .A(n14206), .B(n14205), .Z(n14208) );
  XNOR U13419 ( .A(n14203), .B(n14202), .Z(n14205) );
  XNOR U13420 ( .A(n14200), .B(n14199), .Z(n14202) );
  XNOR U13421 ( .A(n14197), .B(n14196), .Z(n14199) );
  XNOR U13422 ( .A(n14194), .B(n14193), .Z(n14196) );
  XNOR U13423 ( .A(n14191), .B(n14190), .Z(n14193) );
  XNOR U13424 ( .A(n14188), .B(n14187), .Z(n14190) );
  XNOR U13425 ( .A(n14185), .B(n14184), .Z(n14187) );
  XNOR U13426 ( .A(n14182), .B(n14181), .Z(n14184) );
  XNOR U13427 ( .A(n14179), .B(n14178), .Z(n14181) );
  XNOR U13428 ( .A(n14176), .B(n14175), .Z(n14178) );
  XNOR U13429 ( .A(n14173), .B(n14172), .Z(n14175) );
  XNOR U13430 ( .A(n14170), .B(n14169), .Z(n14172) );
  XNOR U13431 ( .A(n14167), .B(n14166), .Z(n14169) );
  XNOR U13432 ( .A(n14164), .B(n14163), .Z(n14166) );
  XNOR U13433 ( .A(n14161), .B(n14160), .Z(n14163) );
  XNOR U13434 ( .A(n14158), .B(n14157), .Z(n14160) );
  XNOR U13435 ( .A(n14155), .B(n14154), .Z(n14157) );
  XNOR U13436 ( .A(n14152), .B(n14151), .Z(n14154) );
  XNOR U13437 ( .A(n14149), .B(n14148), .Z(n14151) );
  XNOR U13438 ( .A(n14146), .B(n14145), .Z(n14148) );
  XNOR U13439 ( .A(n14143), .B(n14142), .Z(n14145) );
  XNOR U13440 ( .A(n14140), .B(n14139), .Z(n14142) );
  XNOR U13441 ( .A(n14137), .B(n14136), .Z(n14139) );
  XNOR U13442 ( .A(n14134), .B(n14133), .Z(n14136) );
  XNOR U13443 ( .A(n14131), .B(n14130), .Z(n14133) );
  XNOR U13444 ( .A(n14128), .B(n14127), .Z(n14130) );
  XNOR U13445 ( .A(n14125), .B(n14124), .Z(n14127) );
  XNOR U13446 ( .A(n14122), .B(n14121), .Z(n14124) );
  XNOR U13447 ( .A(n14119), .B(n14118), .Z(n14121) );
  XNOR U13448 ( .A(n14116), .B(n14115), .Z(n14118) );
  XNOR U13449 ( .A(n14113), .B(n14112), .Z(n14115) );
  XNOR U13450 ( .A(n14110), .B(n14109), .Z(n14112) );
  XNOR U13451 ( .A(n14107), .B(n14106), .Z(n14109) );
  XNOR U13452 ( .A(n14104), .B(n14103), .Z(n14106) );
  XNOR U13453 ( .A(n14101), .B(n14100), .Z(n14103) );
  XNOR U13454 ( .A(n14098), .B(n14097), .Z(n14100) );
  XNOR U13455 ( .A(n14095), .B(n14094), .Z(n14097) );
  XNOR U13456 ( .A(n14092), .B(n14091), .Z(n14094) );
  XNOR U13457 ( .A(n14089), .B(n14088), .Z(n14091) );
  XNOR U13458 ( .A(n14086), .B(n14085), .Z(n14088) );
  XNOR U13459 ( .A(n14083), .B(n14082), .Z(n14085) );
  XNOR U13460 ( .A(n14080), .B(n14079), .Z(n14082) );
  XNOR U13461 ( .A(n14077), .B(n14076), .Z(n14079) );
  XNOR U13462 ( .A(n14074), .B(n14073), .Z(n14076) );
  XNOR U13463 ( .A(n14071), .B(n14070), .Z(n14073) );
  XNOR U13464 ( .A(n14068), .B(n14067), .Z(n14070) );
  XNOR U13465 ( .A(n14065), .B(n14064), .Z(n14067) );
  XNOR U13466 ( .A(n14062), .B(n14061), .Z(n14064) );
  XNOR U13467 ( .A(n14059), .B(n14058), .Z(n14061) );
  XNOR U13468 ( .A(n14056), .B(n14055), .Z(n14058) );
  XNOR U13469 ( .A(n14053), .B(n14052), .Z(n14055) );
  XNOR U13470 ( .A(n14050), .B(n14049), .Z(n14052) );
  XNOR U13471 ( .A(n14047), .B(n14046), .Z(n14049) );
  XNOR U13472 ( .A(n14044), .B(n14043), .Z(n14046) );
  XNOR U13473 ( .A(n14041), .B(n14040), .Z(n14043) );
  XNOR U13474 ( .A(n14038), .B(n14037), .Z(n14040) );
  XNOR U13475 ( .A(n14035), .B(n14034), .Z(n14037) );
  XNOR U13476 ( .A(n14032), .B(n14031), .Z(n14034) );
  XNOR U13477 ( .A(n14029), .B(n14028), .Z(n14031) );
  XNOR U13478 ( .A(n14026), .B(n14025), .Z(n14028) );
  XNOR U13479 ( .A(n14023), .B(n14022), .Z(n14025) );
  XNOR U13480 ( .A(n14020), .B(n14019), .Z(n14022) );
  XNOR U13481 ( .A(n14017), .B(n14016), .Z(n14019) );
  XNOR U13482 ( .A(n14014), .B(n14013), .Z(n14016) );
  XNOR U13483 ( .A(n14011), .B(n14010), .Z(n14013) );
  XNOR U13484 ( .A(n14008), .B(n14007), .Z(n14010) );
  XNOR U13485 ( .A(n14005), .B(n14004), .Z(n14007) );
  XNOR U13486 ( .A(n14002), .B(n14001), .Z(n14004) );
  XNOR U13487 ( .A(n13999), .B(n13998), .Z(n14001) );
  XNOR U13488 ( .A(n13996), .B(n13995), .Z(n13998) );
  XNOR U13489 ( .A(n13993), .B(n13992), .Z(n13995) );
  XNOR U13490 ( .A(n13990), .B(n13989), .Z(n13992) );
  XNOR U13491 ( .A(n13987), .B(n13986), .Z(n13989) );
  XNOR U13492 ( .A(n13984), .B(n13983), .Z(n13986) );
  XNOR U13493 ( .A(n13981), .B(n13980), .Z(n13983) );
  XNOR U13494 ( .A(n13978), .B(n13977), .Z(n13980) );
  XNOR U13495 ( .A(n13975), .B(n13974), .Z(n13977) );
  XNOR U13496 ( .A(n13972), .B(n13971), .Z(n13974) );
  XNOR U13497 ( .A(n13969), .B(n13968), .Z(n13971) );
  XNOR U13498 ( .A(n13966), .B(n13965), .Z(n13968) );
  XNOR U13499 ( .A(n13963), .B(n13962), .Z(n13965) );
  XNOR U13500 ( .A(n13960), .B(n13959), .Z(n13962) );
  XNOR U13501 ( .A(n13957), .B(n13956), .Z(n13959) );
  XNOR U13502 ( .A(n13954), .B(n13953), .Z(n13956) );
  XNOR U13503 ( .A(n13951), .B(n13950), .Z(n13953) );
  XNOR U13504 ( .A(n13948), .B(n13947), .Z(n13950) );
  XNOR U13505 ( .A(n13945), .B(n13944), .Z(n13947) );
  XNOR U13506 ( .A(n13942), .B(n13941), .Z(n13944) );
  XNOR U13507 ( .A(n13939), .B(n13938), .Z(n13941) );
  XNOR U13508 ( .A(n13936), .B(n13935), .Z(n13938) );
  XNOR U13509 ( .A(n13933), .B(n13932), .Z(n13935) );
  XNOR U13510 ( .A(n13930), .B(n13929), .Z(n13932) );
  XNOR U13511 ( .A(n13927), .B(n13926), .Z(n13929) );
  XNOR U13512 ( .A(n13924), .B(n13923), .Z(n13926) );
  XNOR U13513 ( .A(n13921), .B(n13920), .Z(n13923) );
  XNOR U13514 ( .A(n13918), .B(n13917), .Z(n13920) );
  XNOR U13515 ( .A(n13915), .B(n13914), .Z(n13917) );
  XNOR U13516 ( .A(n13912), .B(n13911), .Z(n13914) );
  XNOR U13517 ( .A(n13909), .B(n13908), .Z(n13911) );
  XNOR U13518 ( .A(n13906), .B(n13905), .Z(n13908) );
  XNOR U13519 ( .A(n13903), .B(n13902), .Z(n13905) );
  XNOR U13520 ( .A(n13900), .B(n13899), .Z(n13902) );
  XNOR U13521 ( .A(n13897), .B(n13896), .Z(n13899) );
  XNOR U13522 ( .A(n13894), .B(n13893), .Z(n13896) );
  XNOR U13523 ( .A(n13891), .B(n13890), .Z(n13893) );
  XNOR U13524 ( .A(n13888), .B(n13887), .Z(n13890) );
  XNOR U13525 ( .A(n13885), .B(n13884), .Z(n13887) );
  XNOR U13526 ( .A(n13882), .B(n13881), .Z(n13884) );
  XNOR U13527 ( .A(n13879), .B(n13878), .Z(n13881) );
  XNOR U13528 ( .A(n13876), .B(n13875), .Z(n13878) );
  XNOR U13529 ( .A(n13873), .B(n13872), .Z(n13875) );
  XNOR U13530 ( .A(n13870), .B(n13869), .Z(n13872) );
  XNOR U13531 ( .A(n13867), .B(n13866), .Z(n13869) );
  XNOR U13532 ( .A(n13864), .B(n13863), .Z(n13866) );
  XNOR U13533 ( .A(n13861), .B(n13860), .Z(n13863) );
  XNOR U13534 ( .A(n13858), .B(n13857), .Z(n13860) );
  XNOR U13535 ( .A(n13855), .B(n13854), .Z(n13857) );
  XNOR U13536 ( .A(n13852), .B(n13851), .Z(n13854) );
  XNOR U13537 ( .A(n13849), .B(n13848), .Z(n13851) );
  XNOR U13538 ( .A(n13846), .B(n13845), .Z(n13848) );
  XNOR U13539 ( .A(n13843), .B(n13842), .Z(n13845) );
  XNOR U13540 ( .A(n13840), .B(n13839), .Z(n13842) );
  XNOR U13541 ( .A(n13837), .B(n13836), .Z(n13839) );
  XNOR U13542 ( .A(n13834), .B(n13833), .Z(n13836) );
  XNOR U13543 ( .A(n13831), .B(n13830), .Z(n13833) );
  XNOR U13544 ( .A(n13828), .B(n13827), .Z(n13830) );
  XNOR U13545 ( .A(n13825), .B(n13824), .Z(n13827) );
  XNOR U13546 ( .A(n13822), .B(n13821), .Z(n13824) );
  XNOR U13547 ( .A(n13819), .B(n13818), .Z(n13821) );
  XOR U13548 ( .A(n13816), .B(n13815), .Z(n13818) );
  XOR U13549 ( .A(n13813), .B(n13812), .Z(n13815) );
  XOR U13550 ( .A(n13809), .B(n13810), .Z(n13812) );
  AND U13551 ( .A(n14882), .B(n14883), .Z(n13810) );
  XOR U13552 ( .A(n13806), .B(n13807), .Z(n13809) );
  AND U13553 ( .A(n14884), .B(n14885), .Z(n13807) );
  XOR U13554 ( .A(n13803), .B(n13804), .Z(n13806) );
  AND U13555 ( .A(n14886), .B(n14887), .Z(n13804) );
  XNOR U13556 ( .A(n13558), .B(n13801), .Z(n13803) );
  AND U13557 ( .A(n14888), .B(n14889), .Z(n13801) );
  XOR U13558 ( .A(n13560), .B(n13559), .Z(n13558) );
  AND U13559 ( .A(n14890), .B(n14891), .Z(n13559) );
  XOR U13560 ( .A(n13562), .B(n13561), .Z(n13560) );
  AND U13561 ( .A(n14892), .B(n14893), .Z(n13561) );
  XOR U13562 ( .A(n13564), .B(n13563), .Z(n13562) );
  AND U13563 ( .A(n14894), .B(n14895), .Z(n13563) );
  XOR U13564 ( .A(n13566), .B(n13565), .Z(n13564) );
  AND U13565 ( .A(n14896), .B(n14897), .Z(n13565) );
  XOR U13566 ( .A(n13568), .B(n13567), .Z(n13566) );
  AND U13567 ( .A(n14898), .B(n14899), .Z(n13567) );
  XOR U13568 ( .A(n13570), .B(n13569), .Z(n13568) );
  AND U13569 ( .A(n14900), .B(n14901), .Z(n13569) );
  XOR U13570 ( .A(n13572), .B(n13571), .Z(n13570) );
  AND U13571 ( .A(n14902), .B(n14903), .Z(n13571) );
  XOR U13572 ( .A(n13574), .B(n13573), .Z(n13572) );
  AND U13573 ( .A(n14904), .B(n14905), .Z(n13573) );
  XOR U13574 ( .A(n13576), .B(n13575), .Z(n13574) );
  AND U13575 ( .A(n14906), .B(n14907), .Z(n13575) );
  XOR U13576 ( .A(n13578), .B(n13577), .Z(n13576) );
  AND U13577 ( .A(n14908), .B(n14909), .Z(n13577) );
  XOR U13578 ( .A(n13580), .B(n13579), .Z(n13578) );
  AND U13579 ( .A(n14910), .B(n14911), .Z(n13579) );
  XOR U13580 ( .A(n13582), .B(n13581), .Z(n13580) );
  AND U13581 ( .A(n14912), .B(n14913), .Z(n13581) );
  XOR U13582 ( .A(n13584), .B(n13583), .Z(n13582) );
  AND U13583 ( .A(n14914), .B(n14915), .Z(n13583) );
  XOR U13584 ( .A(n13586), .B(n13585), .Z(n13584) );
  AND U13585 ( .A(n14916), .B(n14917), .Z(n13585) );
  XOR U13586 ( .A(n13588), .B(n13587), .Z(n13586) );
  AND U13587 ( .A(n14918), .B(n14919), .Z(n13587) );
  XOR U13588 ( .A(n13590), .B(n13589), .Z(n13588) );
  AND U13589 ( .A(n14920), .B(n14921), .Z(n13589) );
  XOR U13590 ( .A(n13592), .B(n13591), .Z(n13590) );
  AND U13591 ( .A(n14922), .B(n14923), .Z(n13591) );
  XOR U13592 ( .A(n13594), .B(n13593), .Z(n13592) );
  AND U13593 ( .A(n14924), .B(n14925), .Z(n13593) );
  XOR U13594 ( .A(n13596), .B(n13595), .Z(n13594) );
  AND U13595 ( .A(n14926), .B(n14927), .Z(n13595) );
  XOR U13596 ( .A(n13598), .B(n13597), .Z(n13596) );
  AND U13597 ( .A(n14928), .B(n14929), .Z(n13597) );
  XOR U13598 ( .A(n13600), .B(n13599), .Z(n13598) );
  AND U13599 ( .A(n14930), .B(n14931), .Z(n13599) );
  XOR U13600 ( .A(n13602), .B(n13601), .Z(n13600) );
  AND U13601 ( .A(n14932), .B(n14933), .Z(n13601) );
  XOR U13602 ( .A(n13604), .B(n13603), .Z(n13602) );
  AND U13603 ( .A(n14934), .B(n14935), .Z(n13603) );
  XOR U13604 ( .A(n13606), .B(n13605), .Z(n13604) );
  AND U13605 ( .A(n14936), .B(n14937), .Z(n13605) );
  XOR U13606 ( .A(n13608), .B(n13607), .Z(n13606) );
  AND U13607 ( .A(n14938), .B(n14939), .Z(n13607) );
  XOR U13608 ( .A(n13610), .B(n13609), .Z(n13608) );
  AND U13609 ( .A(n14940), .B(n14941), .Z(n13609) );
  XOR U13610 ( .A(n13612), .B(n13611), .Z(n13610) );
  AND U13611 ( .A(n14942), .B(n14943), .Z(n13611) );
  XOR U13612 ( .A(n13614), .B(n13613), .Z(n13612) );
  AND U13613 ( .A(n14944), .B(n14945), .Z(n13613) );
  XOR U13614 ( .A(n13616), .B(n13615), .Z(n13614) );
  AND U13615 ( .A(n14946), .B(n14947), .Z(n13615) );
  XOR U13616 ( .A(n13618), .B(n13617), .Z(n13616) );
  AND U13617 ( .A(n14948), .B(n14949), .Z(n13617) );
  XOR U13618 ( .A(n13620), .B(n13619), .Z(n13618) );
  AND U13619 ( .A(n14950), .B(n14951), .Z(n13619) );
  XOR U13620 ( .A(n13622), .B(n13621), .Z(n13620) );
  AND U13621 ( .A(n14952), .B(n14953), .Z(n13621) );
  XOR U13622 ( .A(n13624), .B(n13623), .Z(n13622) );
  AND U13623 ( .A(n14954), .B(n14955), .Z(n13623) );
  XOR U13624 ( .A(n13626), .B(n13625), .Z(n13624) );
  AND U13625 ( .A(n14956), .B(n14957), .Z(n13625) );
  XOR U13626 ( .A(n13628), .B(n13627), .Z(n13626) );
  AND U13627 ( .A(n14958), .B(n14959), .Z(n13627) );
  XOR U13628 ( .A(n13630), .B(n13629), .Z(n13628) );
  AND U13629 ( .A(n14960), .B(n14961), .Z(n13629) );
  XOR U13630 ( .A(n13632), .B(n13631), .Z(n13630) );
  AND U13631 ( .A(n14962), .B(n14963), .Z(n13631) );
  XOR U13632 ( .A(n13634), .B(n13633), .Z(n13632) );
  AND U13633 ( .A(n14964), .B(n14965), .Z(n13633) );
  XOR U13634 ( .A(n13636), .B(n13635), .Z(n13634) );
  AND U13635 ( .A(n14966), .B(n14967), .Z(n13635) );
  XOR U13636 ( .A(n13638), .B(n13637), .Z(n13636) );
  AND U13637 ( .A(n14968), .B(n14969), .Z(n13637) );
  XOR U13638 ( .A(n13640), .B(n13639), .Z(n13638) );
  AND U13639 ( .A(n14970), .B(n14971), .Z(n13639) );
  XOR U13640 ( .A(n13642), .B(n13641), .Z(n13640) );
  AND U13641 ( .A(n14972), .B(n14973), .Z(n13641) );
  XOR U13642 ( .A(n13644), .B(n13643), .Z(n13642) );
  AND U13643 ( .A(n14974), .B(n14975), .Z(n13643) );
  XOR U13644 ( .A(n13646), .B(n13645), .Z(n13644) );
  AND U13645 ( .A(n14976), .B(n14977), .Z(n13645) );
  XOR U13646 ( .A(n13648), .B(n13647), .Z(n13646) );
  AND U13647 ( .A(n14978), .B(n14979), .Z(n13647) );
  XOR U13648 ( .A(n13650), .B(n13649), .Z(n13648) );
  AND U13649 ( .A(n14980), .B(n14981), .Z(n13649) );
  XOR U13650 ( .A(n13652), .B(n13651), .Z(n13650) );
  AND U13651 ( .A(n14982), .B(n14983), .Z(n13651) );
  XOR U13652 ( .A(n13654), .B(n13653), .Z(n13652) );
  AND U13653 ( .A(n14984), .B(n14985), .Z(n13653) );
  XOR U13654 ( .A(n13656), .B(n13655), .Z(n13654) );
  AND U13655 ( .A(n14986), .B(n14987), .Z(n13655) );
  XOR U13656 ( .A(n13658), .B(n13657), .Z(n13656) );
  AND U13657 ( .A(n14988), .B(n14989), .Z(n13657) );
  XOR U13658 ( .A(n13660), .B(n13659), .Z(n13658) );
  AND U13659 ( .A(n14990), .B(n14991), .Z(n13659) );
  XOR U13660 ( .A(n13662), .B(n13661), .Z(n13660) );
  AND U13661 ( .A(n14992), .B(n14993), .Z(n13661) );
  XOR U13662 ( .A(n13664), .B(n13663), .Z(n13662) );
  AND U13663 ( .A(n14994), .B(n14995), .Z(n13663) );
  XOR U13664 ( .A(n13666), .B(n13665), .Z(n13664) );
  AND U13665 ( .A(n14996), .B(n14997), .Z(n13665) );
  XOR U13666 ( .A(n13668), .B(n13667), .Z(n13666) );
  AND U13667 ( .A(n14998), .B(n14999), .Z(n13667) );
  XOR U13668 ( .A(n13670), .B(n13669), .Z(n13668) );
  AND U13669 ( .A(n15000), .B(n15001), .Z(n13669) );
  XOR U13670 ( .A(n13672), .B(n13671), .Z(n13670) );
  AND U13671 ( .A(n15002), .B(n15003), .Z(n13671) );
  XOR U13672 ( .A(n13674), .B(n13673), .Z(n13672) );
  AND U13673 ( .A(n15004), .B(n15005), .Z(n13673) );
  XOR U13674 ( .A(n13676), .B(n13675), .Z(n13674) );
  AND U13675 ( .A(n15006), .B(n15007), .Z(n13675) );
  XOR U13676 ( .A(n13678), .B(n13677), .Z(n13676) );
  AND U13677 ( .A(n15008), .B(n15009), .Z(n13677) );
  XOR U13678 ( .A(n13680), .B(n13679), .Z(n13678) );
  AND U13679 ( .A(n15010), .B(n15011), .Z(n13679) );
  XOR U13680 ( .A(n13682), .B(n13681), .Z(n13680) );
  AND U13681 ( .A(n15012), .B(n15013), .Z(n13681) );
  XOR U13682 ( .A(n13684), .B(n13683), .Z(n13682) );
  AND U13683 ( .A(n15014), .B(n15015), .Z(n13683) );
  XOR U13684 ( .A(n13686), .B(n13685), .Z(n13684) );
  AND U13685 ( .A(n15016), .B(n15017), .Z(n13685) );
  XOR U13686 ( .A(n13688), .B(n13687), .Z(n13686) );
  AND U13687 ( .A(n15018), .B(n15019), .Z(n13687) );
  XOR U13688 ( .A(n13690), .B(n13689), .Z(n13688) );
  AND U13689 ( .A(n15020), .B(n15021), .Z(n13689) );
  XOR U13690 ( .A(n13692), .B(n13691), .Z(n13690) );
  AND U13691 ( .A(n15022), .B(n15023), .Z(n13691) );
  XOR U13692 ( .A(n13694), .B(n13693), .Z(n13692) );
  AND U13693 ( .A(n15024), .B(n15025), .Z(n13693) );
  XOR U13694 ( .A(n13703), .B(n13695), .Z(n13694) );
  AND U13695 ( .A(n15026), .B(n15027), .Z(n13695) );
  XOR U13696 ( .A(n13698), .B(n13704), .Z(n13703) );
  AND U13697 ( .A(n15028), .B(n15029), .Z(n13704) );
  XOR U13698 ( .A(n13700), .B(n13699), .Z(n13698) );
  AND U13699 ( .A(n15030), .B(n15031), .Z(n13699) );
  XOR U13700 ( .A(n13724), .B(n13701), .Z(n13700) );
  AND U13701 ( .A(n15032), .B(n15033), .Z(n13701) );
  XOR U13702 ( .A(n13719), .B(n13725), .Z(n13724) );
  AND U13703 ( .A(n15034), .B(n15035), .Z(n13725) );
  XOR U13704 ( .A(n13721), .B(n13720), .Z(n13719) );
  AND U13705 ( .A(n15036), .B(n15037), .Z(n13720) );
  XOR U13706 ( .A(n13709), .B(n13722), .Z(n13721) );
  AND U13707 ( .A(n15038), .B(n15039), .Z(n13722) );
  XOR U13708 ( .A(n13711), .B(n13710), .Z(n13709) );
  AND U13709 ( .A(n15040), .B(n15041), .Z(n13710) );
  XOR U13710 ( .A(n13713), .B(n13712), .Z(n13711) );
  AND U13711 ( .A(n15042), .B(n15043), .Z(n13712) );
  XOR U13712 ( .A(n13715), .B(n13714), .Z(n13713) );
  AND U13713 ( .A(n15044), .B(n15045), .Z(n13714) );
  XOR U13714 ( .A(n13745), .B(n13716), .Z(n13715) );
  AND U13715 ( .A(n15046), .B(n15047), .Z(n13716) );
  XOR U13716 ( .A(n13741), .B(n13746), .Z(n13745) );
  AND U13717 ( .A(n15048), .B(n15049), .Z(n13746) );
  XOR U13718 ( .A(n13743), .B(n13742), .Z(n13741) );
  AND U13719 ( .A(n15050), .B(n15051), .Z(n13742) );
  XOR U13720 ( .A(n13730), .B(n13744), .Z(n13743) );
  AND U13721 ( .A(n15052), .B(n15053), .Z(n13744) );
  XOR U13722 ( .A(n13732), .B(n13731), .Z(n13730) );
  AND U13723 ( .A(n15054), .B(n15055), .Z(n13731) );
  XOR U13724 ( .A(n13735), .B(n13733), .Z(n13732) );
  AND U13725 ( .A(n15056), .B(n15057), .Z(n13733) );
  XOR U13726 ( .A(n13737), .B(n13736), .Z(n13735) );
  AND U13727 ( .A(n15058), .B(n15059), .Z(n13736) );
  XOR U13728 ( .A(n13755), .B(n13738), .Z(n13737) );
  AND U13729 ( .A(n15060), .B(n15061), .Z(n13738) );
  XNOR U13730 ( .A(n13762), .B(n13756), .Z(n13755) );
  AND U13731 ( .A(n15062), .B(n15063), .Z(n13756) );
  XOR U13732 ( .A(n13761), .B(n13753), .Z(n13762) );
  AND U13733 ( .A(n15064), .B(n15065), .Z(n13753) );
  XOR U13734 ( .A(n13800), .B(n13752), .Z(n13761) );
  AND U13735 ( .A(n15066), .B(n15067), .Z(n13752) );
  XNOR U13736 ( .A(n13773), .B(n13751), .Z(n13800) );
  AND U13737 ( .A(n15068), .B(n15069), .Z(n13751) );
  XNOR U13738 ( .A(n13780), .B(n13774), .Z(n13773) );
  AND U13739 ( .A(n15070), .B(n15071), .Z(n13774) );
  XOR U13740 ( .A(n13779), .B(n13771), .Z(n13780) );
  AND U13741 ( .A(n15072), .B(n15073), .Z(n13771) );
  XOR U13742 ( .A(n13799), .B(n13770), .Z(n13779) );
  AND U13743 ( .A(n15074), .B(n15075), .Z(n13770) );
  XNOR U13744 ( .A(n15076), .B(n15077), .Z(n13799) );
  XOR U13745 ( .A(n15078), .B(n15079), .Z(n15077) );
  XOR U13746 ( .A(n15080), .B(n15081), .Z(n15079) );
  XNOR U13747 ( .A(n13797), .B(n13790), .Z(n15081) );
  XNOR U13748 ( .A(n15082), .B(n15083), .Z(n13790) );
  AND U13749 ( .A(n15084), .B(n15085), .Z(n15083) );
  NOR U13750 ( .A(n15086), .B(n15087), .Z(n15085) );
  NOR U13751 ( .A(n15088), .B(n15089), .Z(n15084) );
  AND U13752 ( .A(n15090), .B(n15091), .Z(n15089) );
  AND U13753 ( .A(n15092), .B(n15093), .Z(n15082) );
  NOR U13754 ( .A(n15094), .B(n15095), .Z(n15093) );
  AND U13755 ( .A(n15087), .B(n15096), .Z(n15095) );
  AND U13756 ( .A(n15088), .B(n15097), .Z(n15094) );
  NOR U13757 ( .A(n15098), .B(n15099), .Z(n15092) );
  AND U13758 ( .A(n15100), .B(n15101), .Z(n15099) );
  NOR U13759 ( .A(n15102), .B(n15103), .Z(n15101) );
  IV U13760 ( .A(n15104), .Z(n15102) );
  NOR U13761 ( .A(n15105), .B(n15106), .Z(n15104) );
  NOR U13762 ( .A(n15107), .B(n15108), .Z(n15100) );
  AND U13763 ( .A(n15086), .B(n15109), .Z(n15098) );
  AND U13764 ( .A(n15110), .B(n15111), .Z(n13797) );
  XOR U13765 ( .A(n13795), .B(n13796), .Z(n15080) );
  AND U13766 ( .A(n15112), .B(n15113), .Z(n13796) );
  AND U13767 ( .A(n15114), .B(n15115), .Z(n13795) );
  XOR U13768 ( .A(n15116), .B(n15117), .Z(n15078) );
  XOR U13769 ( .A(n13791), .B(n13792), .Z(n15117) );
  AND U13770 ( .A(n15118), .B(n15119), .Z(n13792) );
  AND U13771 ( .A(n15120), .B(n15121), .Z(n13791) );
  XNOR U13772 ( .A(n13789), .B(n13788), .Z(n15116) );
  IV U13773 ( .A(n15122), .Z(n13788) );
  AND U13774 ( .A(n15123), .B(n15124), .Z(n15122) );
  AND U13775 ( .A(n15125), .B(n15126), .Z(n13789) );
  XNOR U13776 ( .A(n13798), .B(n13769), .Z(n15076) );
  AND U13777 ( .A(n15127), .B(n15128), .Z(n13769) );
  AND U13778 ( .A(n15129), .B(n15130), .Z(n13798) );
  XOR U13779 ( .A(n15131), .B(n15132), .Z(n13813) );
  AND U13780 ( .A(n15131), .B(n15133), .Z(n15132) );
  XNOR U13781 ( .A(n15134), .B(n15135), .Z(n13816) );
  AND U13782 ( .A(n15134), .B(n15136), .Z(n15135) );
  XNOR U13783 ( .A(n15137), .B(n15138), .Z(n13819) );
  AND U13784 ( .A(n15137), .B(n15139), .Z(n15138) );
  XNOR U13785 ( .A(n15140), .B(n15141), .Z(n13822) );
  AND U13786 ( .A(n15140), .B(n15142), .Z(n15141) );
  XNOR U13787 ( .A(n15143), .B(n15144), .Z(n13825) );
  AND U13788 ( .A(n15145), .B(n15143), .Z(n15144) );
  XOR U13789 ( .A(n15146), .B(n15147), .Z(n13828) );
  NOR U13790 ( .A(n15148), .B(n15146), .Z(n15147) );
  XOR U13791 ( .A(n15149), .B(n15150), .Z(n13831) );
  NOR U13792 ( .A(n15151), .B(n15149), .Z(n15150) );
  XOR U13793 ( .A(n15152), .B(n15153), .Z(n13834) );
  NOR U13794 ( .A(n15154), .B(n15152), .Z(n15153) );
  XOR U13795 ( .A(n15155), .B(n15156), .Z(n13837) );
  NOR U13796 ( .A(n15157), .B(n15155), .Z(n15156) );
  XOR U13797 ( .A(n15158), .B(n15159), .Z(n13840) );
  NOR U13798 ( .A(n15160), .B(n15158), .Z(n15159) );
  XOR U13799 ( .A(n15161), .B(n15162), .Z(n13843) );
  NOR U13800 ( .A(n15163), .B(n15161), .Z(n15162) );
  XOR U13801 ( .A(n15164), .B(n15165), .Z(n13846) );
  NOR U13802 ( .A(n15166), .B(n15164), .Z(n15165) );
  XOR U13803 ( .A(n15167), .B(n15168), .Z(n13849) );
  NOR U13804 ( .A(n15169), .B(n15167), .Z(n15168) );
  XOR U13805 ( .A(n15170), .B(n15171), .Z(n13852) );
  NOR U13806 ( .A(n15172), .B(n15170), .Z(n15171) );
  XOR U13807 ( .A(n15173), .B(n15174), .Z(n13855) );
  NOR U13808 ( .A(n15175), .B(n15173), .Z(n15174) );
  XOR U13809 ( .A(n15176), .B(n15177), .Z(n13858) );
  NOR U13810 ( .A(n15178), .B(n15176), .Z(n15177) );
  XOR U13811 ( .A(n15179), .B(n15180), .Z(n13861) );
  NOR U13812 ( .A(n15181), .B(n15179), .Z(n15180) );
  XOR U13813 ( .A(n15182), .B(n15183), .Z(n13864) );
  NOR U13814 ( .A(n15184), .B(n15182), .Z(n15183) );
  XOR U13815 ( .A(n15185), .B(n15186), .Z(n13867) );
  NOR U13816 ( .A(n15187), .B(n15185), .Z(n15186) );
  XOR U13817 ( .A(n15188), .B(n15189), .Z(n13870) );
  NOR U13818 ( .A(n15190), .B(n15188), .Z(n15189) );
  XOR U13819 ( .A(n15191), .B(n15192), .Z(n13873) );
  NOR U13820 ( .A(n15193), .B(n15191), .Z(n15192) );
  XOR U13821 ( .A(n15194), .B(n15195), .Z(n13876) );
  NOR U13822 ( .A(n15196), .B(n15194), .Z(n15195) );
  XOR U13823 ( .A(n15197), .B(n15198), .Z(n13879) );
  NOR U13824 ( .A(n15199), .B(n15197), .Z(n15198) );
  XOR U13825 ( .A(n15200), .B(n15201), .Z(n13882) );
  NOR U13826 ( .A(n15202), .B(n15200), .Z(n15201) );
  XOR U13827 ( .A(n15203), .B(n15204), .Z(n13885) );
  NOR U13828 ( .A(n15205), .B(n15203), .Z(n15204) );
  XOR U13829 ( .A(n15206), .B(n15207), .Z(n13888) );
  NOR U13830 ( .A(n15208), .B(n15206), .Z(n15207) );
  XOR U13831 ( .A(n15209), .B(n15210), .Z(n13891) );
  NOR U13832 ( .A(n15211), .B(n15209), .Z(n15210) );
  XOR U13833 ( .A(n15212), .B(n15213), .Z(n13894) );
  NOR U13834 ( .A(n15214), .B(n15212), .Z(n15213) );
  XOR U13835 ( .A(n15215), .B(n15216), .Z(n13897) );
  NOR U13836 ( .A(n15217), .B(n15215), .Z(n15216) );
  XOR U13837 ( .A(n15218), .B(n15219), .Z(n13900) );
  NOR U13838 ( .A(n15220), .B(n15218), .Z(n15219) );
  XOR U13839 ( .A(n15221), .B(n15222), .Z(n13903) );
  NOR U13840 ( .A(n15223), .B(n15221), .Z(n15222) );
  XOR U13841 ( .A(n15224), .B(n15225), .Z(n13906) );
  NOR U13842 ( .A(n15226), .B(n15224), .Z(n15225) );
  XOR U13843 ( .A(n15227), .B(n15228), .Z(n13909) );
  NOR U13844 ( .A(n15229), .B(n15227), .Z(n15228) );
  XOR U13845 ( .A(n15230), .B(n15231), .Z(n13912) );
  NOR U13846 ( .A(n15232), .B(n15230), .Z(n15231) );
  XOR U13847 ( .A(n15233), .B(n15234), .Z(n13915) );
  NOR U13848 ( .A(n15235), .B(n15233), .Z(n15234) );
  XOR U13849 ( .A(n15236), .B(n15237), .Z(n13918) );
  NOR U13850 ( .A(n15238), .B(n15236), .Z(n15237) );
  XOR U13851 ( .A(n15239), .B(n15240), .Z(n13921) );
  NOR U13852 ( .A(n15241), .B(n15239), .Z(n15240) );
  XOR U13853 ( .A(n15242), .B(n15243), .Z(n13924) );
  NOR U13854 ( .A(n15244), .B(n15242), .Z(n15243) );
  XOR U13855 ( .A(n15245), .B(n15246), .Z(n13927) );
  NOR U13856 ( .A(n15247), .B(n15245), .Z(n15246) );
  XOR U13857 ( .A(n15248), .B(n15249), .Z(n13930) );
  NOR U13858 ( .A(n15250), .B(n15248), .Z(n15249) );
  XOR U13859 ( .A(n15251), .B(n15252), .Z(n13933) );
  NOR U13860 ( .A(n15253), .B(n15251), .Z(n15252) );
  XOR U13861 ( .A(n15254), .B(n15255), .Z(n13936) );
  NOR U13862 ( .A(n15256), .B(n15254), .Z(n15255) );
  XOR U13863 ( .A(n15257), .B(n15258), .Z(n13939) );
  NOR U13864 ( .A(n15259), .B(n15257), .Z(n15258) );
  XOR U13865 ( .A(n15260), .B(n15261), .Z(n13942) );
  NOR U13866 ( .A(n15262), .B(n15260), .Z(n15261) );
  XOR U13867 ( .A(n15263), .B(n15264), .Z(n13945) );
  NOR U13868 ( .A(n15265), .B(n15263), .Z(n15264) );
  XOR U13869 ( .A(n15266), .B(n15267), .Z(n13948) );
  NOR U13870 ( .A(n15268), .B(n15266), .Z(n15267) );
  XOR U13871 ( .A(n15269), .B(n15270), .Z(n13951) );
  NOR U13872 ( .A(n15271), .B(n15269), .Z(n15270) );
  XOR U13873 ( .A(n15272), .B(n15273), .Z(n13954) );
  NOR U13874 ( .A(n15274), .B(n15272), .Z(n15273) );
  XOR U13875 ( .A(n15275), .B(n15276), .Z(n13957) );
  NOR U13876 ( .A(n15277), .B(n15275), .Z(n15276) );
  XOR U13877 ( .A(n15278), .B(n15279), .Z(n13960) );
  NOR U13878 ( .A(n15280), .B(n15278), .Z(n15279) );
  XOR U13879 ( .A(n15281), .B(n15282), .Z(n13963) );
  NOR U13880 ( .A(n15283), .B(n15281), .Z(n15282) );
  XOR U13881 ( .A(n15284), .B(n15285), .Z(n13966) );
  NOR U13882 ( .A(n15286), .B(n15284), .Z(n15285) );
  XOR U13883 ( .A(n15287), .B(n15288), .Z(n13969) );
  NOR U13884 ( .A(n15289), .B(n15287), .Z(n15288) );
  XOR U13885 ( .A(n15290), .B(n15291), .Z(n13972) );
  NOR U13886 ( .A(n15292), .B(n15290), .Z(n15291) );
  XOR U13887 ( .A(n15293), .B(n15294), .Z(n13975) );
  NOR U13888 ( .A(n15295), .B(n15293), .Z(n15294) );
  XOR U13889 ( .A(n15296), .B(n15297), .Z(n13978) );
  NOR U13890 ( .A(n15298), .B(n15296), .Z(n15297) );
  XOR U13891 ( .A(n15299), .B(n15300), .Z(n13981) );
  NOR U13892 ( .A(n15301), .B(n15299), .Z(n15300) );
  XOR U13893 ( .A(n15302), .B(n15303), .Z(n13984) );
  NOR U13894 ( .A(n15304), .B(n15302), .Z(n15303) );
  XOR U13895 ( .A(n15305), .B(n15306), .Z(n13987) );
  NOR U13896 ( .A(n15307), .B(n15305), .Z(n15306) );
  XOR U13897 ( .A(n15308), .B(n15309), .Z(n13990) );
  NOR U13898 ( .A(n15310), .B(n15308), .Z(n15309) );
  XOR U13899 ( .A(n15311), .B(n15312), .Z(n13993) );
  NOR U13900 ( .A(n15313), .B(n15311), .Z(n15312) );
  XOR U13901 ( .A(n15314), .B(n15315), .Z(n13996) );
  NOR U13902 ( .A(n15316), .B(n15314), .Z(n15315) );
  XOR U13903 ( .A(n15317), .B(n15318), .Z(n13999) );
  NOR U13904 ( .A(n15319), .B(n15317), .Z(n15318) );
  XOR U13905 ( .A(n15320), .B(n15321), .Z(n14002) );
  NOR U13906 ( .A(n15322), .B(n15320), .Z(n15321) );
  XOR U13907 ( .A(n15323), .B(n15324), .Z(n14005) );
  NOR U13908 ( .A(n15325), .B(n15323), .Z(n15324) );
  XOR U13909 ( .A(n15326), .B(n15327), .Z(n14008) );
  NOR U13910 ( .A(n15328), .B(n15326), .Z(n15327) );
  XOR U13911 ( .A(n15329), .B(n15330), .Z(n14011) );
  NOR U13912 ( .A(n15331), .B(n15329), .Z(n15330) );
  XOR U13913 ( .A(n15332), .B(n15333), .Z(n14014) );
  NOR U13914 ( .A(n15334), .B(n15332), .Z(n15333) );
  XOR U13915 ( .A(n15335), .B(n15336), .Z(n14017) );
  NOR U13916 ( .A(n15337), .B(n15335), .Z(n15336) );
  XOR U13917 ( .A(n15338), .B(n15339), .Z(n14020) );
  NOR U13918 ( .A(n15340), .B(n15338), .Z(n15339) );
  XOR U13919 ( .A(n15341), .B(n15342), .Z(n14023) );
  NOR U13920 ( .A(n15343), .B(n15341), .Z(n15342) );
  XOR U13921 ( .A(n15344), .B(n15345), .Z(n14026) );
  NOR U13922 ( .A(n15346), .B(n15344), .Z(n15345) );
  XOR U13923 ( .A(n15347), .B(n15348), .Z(n14029) );
  NOR U13924 ( .A(n15349), .B(n15347), .Z(n15348) );
  XOR U13925 ( .A(n15350), .B(n15351), .Z(n14032) );
  NOR U13926 ( .A(n15352), .B(n15350), .Z(n15351) );
  XOR U13927 ( .A(n15353), .B(n15354), .Z(n14035) );
  NOR U13928 ( .A(n15355), .B(n15353), .Z(n15354) );
  XOR U13929 ( .A(n15356), .B(n15357), .Z(n14038) );
  NOR U13930 ( .A(n15358), .B(n15356), .Z(n15357) );
  XOR U13931 ( .A(n15359), .B(n15360), .Z(n14041) );
  NOR U13932 ( .A(n15361), .B(n15359), .Z(n15360) );
  XOR U13933 ( .A(n15362), .B(n15363), .Z(n14044) );
  NOR U13934 ( .A(n15364), .B(n15362), .Z(n15363) );
  XOR U13935 ( .A(n15365), .B(n15366), .Z(n14047) );
  NOR U13936 ( .A(n15367), .B(n15365), .Z(n15366) );
  XOR U13937 ( .A(n15368), .B(n15369), .Z(n14050) );
  NOR U13938 ( .A(n15370), .B(n15368), .Z(n15369) );
  XOR U13939 ( .A(n15371), .B(n15372), .Z(n14053) );
  NOR U13940 ( .A(n15373), .B(n15371), .Z(n15372) );
  XOR U13941 ( .A(n15374), .B(n15375), .Z(n14056) );
  NOR U13942 ( .A(n15376), .B(n15374), .Z(n15375) );
  XOR U13943 ( .A(n15377), .B(n15378), .Z(n14059) );
  NOR U13944 ( .A(n15379), .B(n15377), .Z(n15378) );
  XOR U13945 ( .A(n15380), .B(n15381), .Z(n14062) );
  NOR U13946 ( .A(n15382), .B(n15380), .Z(n15381) );
  XOR U13947 ( .A(n15383), .B(n15384), .Z(n14065) );
  NOR U13948 ( .A(n15385), .B(n15383), .Z(n15384) );
  XOR U13949 ( .A(n15386), .B(n15387), .Z(n14068) );
  NOR U13950 ( .A(n15388), .B(n15386), .Z(n15387) );
  XOR U13951 ( .A(n15389), .B(n15390), .Z(n14071) );
  NOR U13952 ( .A(n15391), .B(n15389), .Z(n15390) );
  XOR U13953 ( .A(n15392), .B(n15393), .Z(n14074) );
  NOR U13954 ( .A(n15394), .B(n15392), .Z(n15393) );
  XOR U13955 ( .A(n15395), .B(n15396), .Z(n14077) );
  NOR U13956 ( .A(n15397), .B(n15395), .Z(n15396) );
  XOR U13957 ( .A(n15398), .B(n15399), .Z(n14080) );
  NOR U13958 ( .A(n15400), .B(n15398), .Z(n15399) );
  XOR U13959 ( .A(n15401), .B(n15402), .Z(n14083) );
  NOR U13960 ( .A(n15403), .B(n15401), .Z(n15402) );
  XOR U13961 ( .A(n15404), .B(n15405), .Z(n14086) );
  NOR U13962 ( .A(n15406), .B(n15404), .Z(n15405) );
  XOR U13963 ( .A(n15407), .B(n15408), .Z(n14089) );
  NOR U13964 ( .A(n15409), .B(n15407), .Z(n15408) );
  XOR U13965 ( .A(n15410), .B(n15411), .Z(n14092) );
  NOR U13966 ( .A(n15412), .B(n15410), .Z(n15411) );
  XOR U13967 ( .A(n15413), .B(n15414), .Z(n14095) );
  NOR U13968 ( .A(n15415), .B(n15413), .Z(n15414) );
  XOR U13969 ( .A(n15416), .B(n15417), .Z(n14098) );
  NOR U13970 ( .A(n15418), .B(n15416), .Z(n15417) );
  XOR U13971 ( .A(n15419), .B(n15420), .Z(n14101) );
  NOR U13972 ( .A(n15421), .B(n15419), .Z(n15420) );
  XOR U13973 ( .A(n15422), .B(n15423), .Z(n14104) );
  NOR U13974 ( .A(n15424), .B(n15422), .Z(n15423) );
  XOR U13975 ( .A(n15425), .B(n15426), .Z(n14107) );
  NOR U13976 ( .A(n15427), .B(n15425), .Z(n15426) );
  XOR U13977 ( .A(n15428), .B(n15429), .Z(n14110) );
  NOR U13978 ( .A(n15430), .B(n15428), .Z(n15429) );
  XOR U13979 ( .A(n15431), .B(n15432), .Z(n14113) );
  NOR U13980 ( .A(n15433), .B(n15431), .Z(n15432) );
  XOR U13981 ( .A(n15434), .B(n15435), .Z(n14116) );
  NOR U13982 ( .A(n15436), .B(n15434), .Z(n15435) );
  XOR U13983 ( .A(n15437), .B(n15438), .Z(n14119) );
  NOR U13984 ( .A(n15439), .B(n15437), .Z(n15438) );
  XOR U13985 ( .A(n15440), .B(n15441), .Z(n14122) );
  NOR U13986 ( .A(n15442), .B(n15440), .Z(n15441) );
  XOR U13987 ( .A(n15443), .B(n15444), .Z(n14125) );
  NOR U13988 ( .A(n15445), .B(n15443), .Z(n15444) );
  XOR U13989 ( .A(n15446), .B(n15447), .Z(n14128) );
  NOR U13990 ( .A(n15448), .B(n15446), .Z(n15447) );
  XOR U13991 ( .A(n15449), .B(n15450), .Z(n14131) );
  NOR U13992 ( .A(n15451), .B(n15449), .Z(n15450) );
  XOR U13993 ( .A(n15452), .B(n15453), .Z(n14134) );
  NOR U13994 ( .A(n15454), .B(n15452), .Z(n15453) );
  XOR U13995 ( .A(n15455), .B(n15456), .Z(n14137) );
  NOR U13996 ( .A(n15457), .B(n15455), .Z(n15456) );
  XOR U13997 ( .A(n15458), .B(n15459), .Z(n14140) );
  NOR U13998 ( .A(n15460), .B(n15458), .Z(n15459) );
  XOR U13999 ( .A(n15461), .B(n15462), .Z(n14143) );
  NOR U14000 ( .A(n15463), .B(n15461), .Z(n15462) );
  XOR U14001 ( .A(n15464), .B(n15465), .Z(n14146) );
  NOR U14002 ( .A(n15466), .B(n15464), .Z(n15465) );
  XOR U14003 ( .A(n15467), .B(n15468), .Z(n14149) );
  NOR U14004 ( .A(n15469), .B(n15467), .Z(n15468) );
  XOR U14005 ( .A(n15470), .B(n15471), .Z(n14152) );
  NOR U14006 ( .A(n15472), .B(n15470), .Z(n15471) );
  XOR U14007 ( .A(n15473), .B(n15474), .Z(n14155) );
  NOR U14008 ( .A(n15475), .B(n15473), .Z(n15474) );
  XOR U14009 ( .A(n15476), .B(n15477), .Z(n14158) );
  NOR U14010 ( .A(n15478), .B(n15476), .Z(n15477) );
  XOR U14011 ( .A(n15479), .B(n15480), .Z(n14161) );
  NOR U14012 ( .A(n15481), .B(n15479), .Z(n15480) );
  XOR U14013 ( .A(n15482), .B(n15483), .Z(n14164) );
  NOR U14014 ( .A(n15484), .B(n15482), .Z(n15483) );
  XOR U14015 ( .A(n15485), .B(n15486), .Z(n14167) );
  NOR U14016 ( .A(n15487), .B(n15485), .Z(n15486) );
  XOR U14017 ( .A(n15488), .B(n15489), .Z(n14170) );
  NOR U14018 ( .A(n15490), .B(n15488), .Z(n15489) );
  XOR U14019 ( .A(n15491), .B(n15492), .Z(n14173) );
  NOR U14020 ( .A(n15493), .B(n15491), .Z(n15492) );
  XOR U14021 ( .A(n15494), .B(n15495), .Z(n14176) );
  NOR U14022 ( .A(n15496), .B(n15494), .Z(n15495) );
  XOR U14023 ( .A(n15497), .B(n15498), .Z(n14179) );
  NOR U14024 ( .A(n15499), .B(n15497), .Z(n15498) );
  XOR U14025 ( .A(n15500), .B(n15501), .Z(n14182) );
  NOR U14026 ( .A(n15502), .B(n15500), .Z(n15501) );
  XOR U14027 ( .A(n15503), .B(n15504), .Z(n14185) );
  NOR U14028 ( .A(n15505), .B(n15503), .Z(n15504) );
  XOR U14029 ( .A(n15506), .B(n15507), .Z(n14188) );
  NOR U14030 ( .A(n15508), .B(n15506), .Z(n15507) );
  XOR U14031 ( .A(n15509), .B(n15510), .Z(n14191) );
  NOR U14032 ( .A(n15511), .B(n15509), .Z(n15510) );
  XOR U14033 ( .A(n15512), .B(n15513), .Z(n14194) );
  NOR U14034 ( .A(n15514), .B(n15512), .Z(n15513) );
  XOR U14035 ( .A(n15515), .B(n15516), .Z(n14197) );
  NOR U14036 ( .A(n15517), .B(n15515), .Z(n15516) );
  XOR U14037 ( .A(n15518), .B(n15519), .Z(n14200) );
  NOR U14038 ( .A(n15520), .B(n15518), .Z(n15519) );
  XOR U14039 ( .A(n15521), .B(n15522), .Z(n14203) );
  NOR U14040 ( .A(n15523), .B(n15521), .Z(n15522) );
  XOR U14041 ( .A(n15524), .B(n15525), .Z(n14206) );
  NOR U14042 ( .A(n15526), .B(n15524), .Z(n15525) );
  XOR U14043 ( .A(n15527), .B(n15528), .Z(n14209) );
  NOR U14044 ( .A(n15529), .B(n15527), .Z(n15528) );
  XNOR U14045 ( .A(n15530), .B(n15531), .Z(n14212) );
  NOR U14046 ( .A(n15532), .B(n15530), .Z(n15531) );
  XOR U14047 ( .A(n15533), .B(n15534), .Z(n14215) );
  AND U14048 ( .A(n108), .B(n15533), .Z(n15534) );
  XOR U14049 ( .A(n90), .B(n14878), .Z(n14880) );
  XOR U14050 ( .A(n14875), .B(n14874), .Z(n90) );
  XNOR U14051 ( .A(n14872), .B(n14871), .Z(n14874) );
  XNOR U14052 ( .A(n14869), .B(n14868), .Z(n14871) );
  XNOR U14053 ( .A(n14866), .B(n14865), .Z(n14868) );
  XNOR U14054 ( .A(n14863), .B(n14862), .Z(n14865) );
  XNOR U14055 ( .A(n14860), .B(n14859), .Z(n14862) );
  XNOR U14056 ( .A(n14857), .B(n14856), .Z(n14859) );
  XNOR U14057 ( .A(n14854), .B(n14853), .Z(n14856) );
  XNOR U14058 ( .A(n14851), .B(n14850), .Z(n14853) );
  XNOR U14059 ( .A(n14848), .B(n14847), .Z(n14850) );
  XNOR U14060 ( .A(n14845), .B(n14844), .Z(n14847) );
  XNOR U14061 ( .A(n14842), .B(n14841), .Z(n14844) );
  XNOR U14062 ( .A(n14839), .B(n14838), .Z(n14841) );
  XNOR U14063 ( .A(n14836), .B(n14835), .Z(n14838) );
  XNOR U14064 ( .A(n14833), .B(n14832), .Z(n14835) );
  XNOR U14065 ( .A(n14830), .B(n14829), .Z(n14832) );
  XNOR U14066 ( .A(n14827), .B(n14826), .Z(n14829) );
  XNOR U14067 ( .A(n14824), .B(n14823), .Z(n14826) );
  XNOR U14068 ( .A(n14821), .B(n14820), .Z(n14823) );
  XNOR U14069 ( .A(n14818), .B(n14817), .Z(n14820) );
  XNOR U14070 ( .A(n14815), .B(n14814), .Z(n14817) );
  XNOR U14071 ( .A(n14812), .B(n14811), .Z(n14814) );
  XNOR U14072 ( .A(n14809), .B(n14808), .Z(n14811) );
  XNOR U14073 ( .A(n14806), .B(n14805), .Z(n14808) );
  XNOR U14074 ( .A(n14803), .B(n14802), .Z(n14805) );
  XNOR U14075 ( .A(n14800), .B(n14799), .Z(n14802) );
  XNOR U14076 ( .A(n14797), .B(n14796), .Z(n14799) );
  XNOR U14077 ( .A(n14794), .B(n14793), .Z(n14796) );
  XNOR U14078 ( .A(n14791), .B(n14790), .Z(n14793) );
  XNOR U14079 ( .A(n14788), .B(n14787), .Z(n14790) );
  XNOR U14080 ( .A(n14785), .B(n14784), .Z(n14787) );
  XNOR U14081 ( .A(n14782), .B(n14781), .Z(n14784) );
  XNOR U14082 ( .A(n14779), .B(n14778), .Z(n14781) );
  XNOR U14083 ( .A(n14776), .B(n14775), .Z(n14778) );
  XNOR U14084 ( .A(n14773), .B(n14772), .Z(n14775) );
  XNOR U14085 ( .A(n14770), .B(n14769), .Z(n14772) );
  XNOR U14086 ( .A(n14767), .B(n14766), .Z(n14769) );
  XNOR U14087 ( .A(n14764), .B(n14763), .Z(n14766) );
  XNOR U14088 ( .A(n14761), .B(n14760), .Z(n14763) );
  XNOR U14089 ( .A(n14758), .B(n14757), .Z(n14760) );
  XNOR U14090 ( .A(n14755), .B(n14754), .Z(n14757) );
  XNOR U14091 ( .A(n14752), .B(n14751), .Z(n14754) );
  XNOR U14092 ( .A(n14749), .B(n14748), .Z(n14751) );
  XNOR U14093 ( .A(n14746), .B(n14745), .Z(n14748) );
  XNOR U14094 ( .A(n14743), .B(n14742), .Z(n14745) );
  XNOR U14095 ( .A(n14740), .B(n14739), .Z(n14742) );
  XNOR U14096 ( .A(n14737), .B(n14736), .Z(n14739) );
  XNOR U14097 ( .A(n14734), .B(n14733), .Z(n14736) );
  XNOR U14098 ( .A(n14731), .B(n14730), .Z(n14733) );
  XNOR U14099 ( .A(n14728), .B(n14727), .Z(n14730) );
  XNOR U14100 ( .A(n14725), .B(n14724), .Z(n14727) );
  XNOR U14101 ( .A(n14722), .B(n14721), .Z(n14724) );
  XNOR U14102 ( .A(n14719), .B(n14718), .Z(n14721) );
  XNOR U14103 ( .A(n14716), .B(n14715), .Z(n14718) );
  XNOR U14104 ( .A(n14713), .B(n14712), .Z(n14715) );
  XNOR U14105 ( .A(n14710), .B(n14709), .Z(n14712) );
  XNOR U14106 ( .A(n14707), .B(n14706), .Z(n14709) );
  XNOR U14107 ( .A(n14704), .B(n14703), .Z(n14706) );
  XNOR U14108 ( .A(n14701), .B(n14700), .Z(n14703) );
  XNOR U14109 ( .A(n14698), .B(n14697), .Z(n14700) );
  XNOR U14110 ( .A(n14695), .B(n14694), .Z(n14697) );
  XNOR U14111 ( .A(n14692), .B(n14691), .Z(n14694) );
  XNOR U14112 ( .A(n14689), .B(n14688), .Z(n14691) );
  XNOR U14113 ( .A(n14686), .B(n14685), .Z(n14688) );
  XNOR U14114 ( .A(n14683), .B(n14682), .Z(n14685) );
  XNOR U14115 ( .A(n14680), .B(n14679), .Z(n14682) );
  XNOR U14116 ( .A(n14677), .B(n14676), .Z(n14679) );
  XNOR U14117 ( .A(n14674), .B(n14673), .Z(n14676) );
  XNOR U14118 ( .A(n14671), .B(n14670), .Z(n14673) );
  XNOR U14119 ( .A(n14668), .B(n14667), .Z(n14670) );
  XNOR U14120 ( .A(n14665), .B(n14664), .Z(n14667) );
  XNOR U14121 ( .A(n14662), .B(n14661), .Z(n14664) );
  XNOR U14122 ( .A(n14659), .B(n14658), .Z(n14661) );
  XNOR U14123 ( .A(n14656), .B(n14655), .Z(n14658) );
  XNOR U14124 ( .A(n14653), .B(n14652), .Z(n14655) );
  XNOR U14125 ( .A(n14650), .B(n14649), .Z(n14652) );
  XNOR U14126 ( .A(n14647), .B(n14646), .Z(n14649) );
  XNOR U14127 ( .A(n14644), .B(n14643), .Z(n14646) );
  XNOR U14128 ( .A(n14641), .B(n14640), .Z(n14643) );
  XNOR U14129 ( .A(n14638), .B(n14637), .Z(n14640) );
  XNOR U14130 ( .A(n14635), .B(n14634), .Z(n14637) );
  XNOR U14131 ( .A(n14632), .B(n14631), .Z(n14634) );
  XNOR U14132 ( .A(n14629), .B(n14628), .Z(n14631) );
  XNOR U14133 ( .A(n14626), .B(n14625), .Z(n14628) );
  XNOR U14134 ( .A(n14623), .B(n14622), .Z(n14625) );
  XNOR U14135 ( .A(n14620), .B(n14619), .Z(n14622) );
  XNOR U14136 ( .A(n14617), .B(n14616), .Z(n14619) );
  XNOR U14137 ( .A(n14614), .B(n14613), .Z(n14616) );
  XNOR U14138 ( .A(n14611), .B(n14610), .Z(n14613) );
  XNOR U14139 ( .A(n14608), .B(n14607), .Z(n14610) );
  XNOR U14140 ( .A(n14605), .B(n14604), .Z(n14607) );
  XNOR U14141 ( .A(n14602), .B(n14601), .Z(n14604) );
  XNOR U14142 ( .A(n14599), .B(n14598), .Z(n14601) );
  XNOR U14143 ( .A(n14596), .B(n14595), .Z(n14598) );
  XNOR U14144 ( .A(n14593), .B(n14592), .Z(n14595) );
  XNOR U14145 ( .A(n14590), .B(n14589), .Z(n14592) );
  XNOR U14146 ( .A(n14587), .B(n14586), .Z(n14589) );
  XNOR U14147 ( .A(n14584), .B(n14583), .Z(n14586) );
  XNOR U14148 ( .A(n14581), .B(n14580), .Z(n14583) );
  XNOR U14149 ( .A(n14578), .B(n14577), .Z(n14580) );
  XNOR U14150 ( .A(n14575), .B(n14574), .Z(n14577) );
  XNOR U14151 ( .A(n14572), .B(n14571), .Z(n14574) );
  XNOR U14152 ( .A(n14569), .B(n14568), .Z(n14571) );
  XNOR U14153 ( .A(n14566), .B(n14565), .Z(n14568) );
  XNOR U14154 ( .A(n14563), .B(n14562), .Z(n14565) );
  XNOR U14155 ( .A(n14560), .B(n14559), .Z(n14562) );
  XNOR U14156 ( .A(n14557), .B(n14556), .Z(n14559) );
  XNOR U14157 ( .A(n14554), .B(n14553), .Z(n14556) );
  XNOR U14158 ( .A(n14551), .B(n14550), .Z(n14553) );
  XNOR U14159 ( .A(n14548), .B(n14547), .Z(n14550) );
  XNOR U14160 ( .A(n14545), .B(n14544), .Z(n14547) );
  XNOR U14161 ( .A(n14542), .B(n14541), .Z(n14544) );
  XNOR U14162 ( .A(n14539), .B(n14538), .Z(n14541) );
  XNOR U14163 ( .A(n14536), .B(n14535), .Z(n14538) );
  XNOR U14164 ( .A(n14533), .B(n14532), .Z(n14535) );
  XNOR U14165 ( .A(n14530), .B(n14529), .Z(n14532) );
  XNOR U14166 ( .A(n14527), .B(n14526), .Z(n14529) );
  XNOR U14167 ( .A(n14524), .B(n14523), .Z(n14526) );
  XNOR U14168 ( .A(n14521), .B(n14520), .Z(n14523) );
  XNOR U14169 ( .A(n14518), .B(n14517), .Z(n14520) );
  XNOR U14170 ( .A(n14515), .B(n14514), .Z(n14517) );
  XNOR U14171 ( .A(n14512), .B(n14511), .Z(n14514) );
  XNOR U14172 ( .A(n14509), .B(n14508), .Z(n14511) );
  XNOR U14173 ( .A(n14506), .B(n14505), .Z(n14508) );
  XNOR U14174 ( .A(n14503), .B(n14502), .Z(n14505) );
  XNOR U14175 ( .A(n14500), .B(n14499), .Z(n14502) );
  XNOR U14176 ( .A(n14497), .B(n14496), .Z(n14499) );
  XNOR U14177 ( .A(n14494), .B(n14493), .Z(n14496) );
  XNOR U14178 ( .A(n14491), .B(n14490), .Z(n14493) );
  XNOR U14179 ( .A(n14488), .B(n14487), .Z(n14490) );
  XNOR U14180 ( .A(n14485), .B(n14484), .Z(n14487) );
  XNOR U14181 ( .A(n14482), .B(n14481), .Z(n14484) );
  XNOR U14182 ( .A(n14479), .B(n14478), .Z(n14481) );
  XOR U14183 ( .A(n14476), .B(n14475), .Z(n14478) );
  XOR U14184 ( .A(n14473), .B(n14472), .Z(n14475) );
  XOR U14185 ( .A(n14469), .B(n14470), .Z(n14472) );
  AND U14186 ( .A(n15535), .B(n15536), .Z(n14470) );
  XOR U14187 ( .A(n14466), .B(n14467), .Z(n14469) );
  AND U14188 ( .A(n15537), .B(n15538), .Z(n14467) );
  XOR U14189 ( .A(n14463), .B(n14464), .Z(n14466) );
  AND U14190 ( .A(n15539), .B(n15540), .Z(n14464) );
  XNOR U14191 ( .A(n14218), .B(n14461), .Z(n14463) );
  AND U14192 ( .A(n15541), .B(n15542), .Z(n14461) );
  XOR U14193 ( .A(n14220), .B(n14219), .Z(n14218) );
  AND U14194 ( .A(n15543), .B(n15544), .Z(n14219) );
  XOR U14195 ( .A(n14222), .B(n14221), .Z(n14220) );
  AND U14196 ( .A(n15545), .B(n15546), .Z(n14221) );
  XOR U14197 ( .A(n14224), .B(n14223), .Z(n14222) );
  AND U14198 ( .A(n15547), .B(n15548), .Z(n14223) );
  XOR U14199 ( .A(n14226), .B(n14225), .Z(n14224) );
  AND U14200 ( .A(n15549), .B(n15550), .Z(n14225) );
  XOR U14201 ( .A(n14228), .B(n14227), .Z(n14226) );
  AND U14202 ( .A(n15551), .B(n15552), .Z(n14227) );
  XOR U14203 ( .A(n14230), .B(n14229), .Z(n14228) );
  AND U14204 ( .A(n15553), .B(n15554), .Z(n14229) );
  XOR U14205 ( .A(n14232), .B(n14231), .Z(n14230) );
  AND U14206 ( .A(n15555), .B(n15556), .Z(n14231) );
  XOR U14207 ( .A(n14234), .B(n14233), .Z(n14232) );
  AND U14208 ( .A(n15557), .B(n15558), .Z(n14233) );
  XOR U14209 ( .A(n14236), .B(n14235), .Z(n14234) );
  AND U14210 ( .A(n15559), .B(n15560), .Z(n14235) );
  XOR U14211 ( .A(n14238), .B(n14237), .Z(n14236) );
  AND U14212 ( .A(n15561), .B(n15562), .Z(n14237) );
  XOR U14213 ( .A(n14240), .B(n14239), .Z(n14238) );
  AND U14214 ( .A(n15563), .B(n15564), .Z(n14239) );
  XOR U14215 ( .A(n14242), .B(n14241), .Z(n14240) );
  AND U14216 ( .A(n15565), .B(n15566), .Z(n14241) );
  XOR U14217 ( .A(n14244), .B(n14243), .Z(n14242) );
  AND U14218 ( .A(n15567), .B(n15568), .Z(n14243) );
  XOR U14219 ( .A(n14246), .B(n14245), .Z(n14244) );
  AND U14220 ( .A(n15569), .B(n15570), .Z(n14245) );
  XOR U14221 ( .A(n14248), .B(n14247), .Z(n14246) );
  AND U14222 ( .A(n15571), .B(n15572), .Z(n14247) );
  XOR U14223 ( .A(n14250), .B(n14249), .Z(n14248) );
  AND U14224 ( .A(n15573), .B(n15574), .Z(n14249) );
  XOR U14225 ( .A(n14252), .B(n14251), .Z(n14250) );
  AND U14226 ( .A(n15575), .B(n15576), .Z(n14251) );
  XOR U14227 ( .A(n14254), .B(n14253), .Z(n14252) );
  AND U14228 ( .A(n15577), .B(n15578), .Z(n14253) );
  XOR U14229 ( .A(n14256), .B(n14255), .Z(n14254) );
  AND U14230 ( .A(n15579), .B(n15580), .Z(n14255) );
  XOR U14231 ( .A(n14258), .B(n14257), .Z(n14256) );
  AND U14232 ( .A(n15581), .B(n15582), .Z(n14257) );
  XOR U14233 ( .A(n14260), .B(n14259), .Z(n14258) );
  AND U14234 ( .A(n15583), .B(n15584), .Z(n14259) );
  XOR U14235 ( .A(n14262), .B(n14261), .Z(n14260) );
  AND U14236 ( .A(n15585), .B(n15586), .Z(n14261) );
  XOR U14237 ( .A(n14264), .B(n14263), .Z(n14262) );
  AND U14238 ( .A(n15587), .B(n15588), .Z(n14263) );
  XOR U14239 ( .A(n14266), .B(n14265), .Z(n14264) );
  AND U14240 ( .A(n15589), .B(n15590), .Z(n14265) );
  XOR U14241 ( .A(n14268), .B(n14267), .Z(n14266) );
  AND U14242 ( .A(n15591), .B(n15592), .Z(n14267) );
  XOR U14243 ( .A(n14270), .B(n14269), .Z(n14268) );
  AND U14244 ( .A(n15593), .B(n15594), .Z(n14269) );
  XOR U14245 ( .A(n14272), .B(n14271), .Z(n14270) );
  AND U14246 ( .A(n15595), .B(n15596), .Z(n14271) );
  XOR U14247 ( .A(n14274), .B(n14273), .Z(n14272) );
  AND U14248 ( .A(n15597), .B(n15598), .Z(n14273) );
  XOR U14249 ( .A(n14276), .B(n14275), .Z(n14274) );
  AND U14250 ( .A(n15599), .B(n15600), .Z(n14275) );
  XOR U14251 ( .A(n14278), .B(n14277), .Z(n14276) );
  AND U14252 ( .A(n15601), .B(n15602), .Z(n14277) );
  XOR U14253 ( .A(n14280), .B(n14279), .Z(n14278) );
  AND U14254 ( .A(n15603), .B(n15604), .Z(n14279) );
  XOR U14255 ( .A(n14282), .B(n14281), .Z(n14280) );
  AND U14256 ( .A(n15605), .B(n15606), .Z(n14281) );
  XOR U14257 ( .A(n14284), .B(n14283), .Z(n14282) );
  AND U14258 ( .A(n15607), .B(n15608), .Z(n14283) );
  XOR U14259 ( .A(n14286), .B(n14285), .Z(n14284) );
  AND U14260 ( .A(n15609), .B(n15610), .Z(n14285) );
  XOR U14261 ( .A(n14288), .B(n14287), .Z(n14286) );
  AND U14262 ( .A(n15611), .B(n15612), .Z(n14287) );
  XOR U14263 ( .A(n14290), .B(n14289), .Z(n14288) );
  AND U14264 ( .A(n15613), .B(n15614), .Z(n14289) );
  XOR U14265 ( .A(n14292), .B(n14291), .Z(n14290) );
  AND U14266 ( .A(n15615), .B(n15616), .Z(n14291) );
  XOR U14267 ( .A(n14294), .B(n14293), .Z(n14292) );
  AND U14268 ( .A(n15617), .B(n15618), .Z(n14293) );
  XOR U14269 ( .A(n14296), .B(n14295), .Z(n14294) );
  AND U14270 ( .A(n15619), .B(n15620), .Z(n14295) );
  XOR U14271 ( .A(n14298), .B(n14297), .Z(n14296) );
  AND U14272 ( .A(n15621), .B(n15622), .Z(n14297) );
  XOR U14273 ( .A(n14300), .B(n14299), .Z(n14298) );
  AND U14274 ( .A(n15623), .B(n15624), .Z(n14299) );
  XOR U14275 ( .A(n14302), .B(n14301), .Z(n14300) );
  AND U14276 ( .A(n15625), .B(n15626), .Z(n14301) );
  XOR U14277 ( .A(n14304), .B(n14303), .Z(n14302) );
  AND U14278 ( .A(n15627), .B(n15628), .Z(n14303) );
  XOR U14279 ( .A(n14306), .B(n14305), .Z(n14304) );
  AND U14280 ( .A(n15629), .B(n15630), .Z(n14305) );
  XOR U14281 ( .A(n14308), .B(n14307), .Z(n14306) );
  AND U14282 ( .A(n15631), .B(n15632), .Z(n14307) );
  XOR U14283 ( .A(n14310), .B(n14309), .Z(n14308) );
  AND U14284 ( .A(n15633), .B(n15634), .Z(n14309) );
  XOR U14285 ( .A(n14312), .B(n14311), .Z(n14310) );
  AND U14286 ( .A(n15635), .B(n15636), .Z(n14311) );
  XOR U14287 ( .A(n14314), .B(n14313), .Z(n14312) );
  AND U14288 ( .A(n15637), .B(n15638), .Z(n14313) );
  XOR U14289 ( .A(n14316), .B(n14315), .Z(n14314) );
  AND U14290 ( .A(n15639), .B(n15640), .Z(n14315) );
  XOR U14291 ( .A(n14318), .B(n14317), .Z(n14316) );
  AND U14292 ( .A(n15641), .B(n15642), .Z(n14317) );
  XOR U14293 ( .A(n14320), .B(n14319), .Z(n14318) );
  AND U14294 ( .A(n15643), .B(n15644), .Z(n14319) );
  XOR U14295 ( .A(n14322), .B(n14321), .Z(n14320) );
  AND U14296 ( .A(n15645), .B(n15646), .Z(n14321) );
  XOR U14297 ( .A(n14324), .B(n14323), .Z(n14322) );
  AND U14298 ( .A(n15647), .B(n15648), .Z(n14323) );
  XOR U14299 ( .A(n14326), .B(n14325), .Z(n14324) );
  AND U14300 ( .A(n15649), .B(n15650), .Z(n14325) );
  XOR U14301 ( .A(n14328), .B(n14327), .Z(n14326) );
  AND U14302 ( .A(n15651), .B(n15652), .Z(n14327) );
  XOR U14303 ( .A(n14330), .B(n14329), .Z(n14328) );
  AND U14304 ( .A(n15653), .B(n15654), .Z(n14329) );
  XOR U14305 ( .A(n14332), .B(n14331), .Z(n14330) );
  AND U14306 ( .A(n15655), .B(n15656), .Z(n14331) );
  XOR U14307 ( .A(n14334), .B(n14333), .Z(n14332) );
  AND U14308 ( .A(n15657), .B(n15658), .Z(n14333) );
  XOR U14309 ( .A(n14336), .B(n14335), .Z(n14334) );
  AND U14310 ( .A(n15659), .B(n15660), .Z(n14335) );
  XOR U14311 ( .A(n14338), .B(n14337), .Z(n14336) );
  AND U14312 ( .A(n15661), .B(n15662), .Z(n14337) );
  XOR U14313 ( .A(n14340), .B(n14339), .Z(n14338) );
  AND U14314 ( .A(n15663), .B(n15664), .Z(n14339) );
  XOR U14315 ( .A(n14342), .B(n14341), .Z(n14340) );
  AND U14316 ( .A(n15665), .B(n15666), .Z(n14341) );
  XOR U14317 ( .A(n14344), .B(n14343), .Z(n14342) );
  AND U14318 ( .A(n15667), .B(n15668), .Z(n14343) );
  XOR U14319 ( .A(n14346), .B(n14345), .Z(n14344) );
  AND U14320 ( .A(n15669), .B(n15670), .Z(n14345) );
  XOR U14321 ( .A(n14348), .B(n14347), .Z(n14346) );
  AND U14322 ( .A(n15671), .B(n15672), .Z(n14347) );
  XOR U14323 ( .A(n14350), .B(n14349), .Z(n14348) );
  AND U14324 ( .A(n15673), .B(n15674), .Z(n14349) );
  XOR U14325 ( .A(n14352), .B(n14351), .Z(n14350) );
  AND U14326 ( .A(n15675), .B(n15676), .Z(n14351) );
  XOR U14327 ( .A(n14354), .B(n14353), .Z(n14352) );
  AND U14328 ( .A(n15677), .B(n15678), .Z(n14353) );
  XOR U14329 ( .A(n14363), .B(n14355), .Z(n14354) );
  AND U14330 ( .A(n15679), .B(n15680), .Z(n14355) );
  XOR U14331 ( .A(n14358), .B(n14364), .Z(n14363) );
  AND U14332 ( .A(n15681), .B(n15682), .Z(n14364) );
  XOR U14333 ( .A(n14360), .B(n14359), .Z(n14358) );
  AND U14334 ( .A(n15683), .B(n15684), .Z(n14359) );
  XOR U14335 ( .A(n14384), .B(n14361), .Z(n14360) );
  AND U14336 ( .A(n15685), .B(n15686), .Z(n14361) );
  XOR U14337 ( .A(n14379), .B(n14385), .Z(n14384) );
  AND U14338 ( .A(n15687), .B(n15688), .Z(n14385) );
  XOR U14339 ( .A(n14381), .B(n14380), .Z(n14379) );
  AND U14340 ( .A(n15689), .B(n15690), .Z(n14380) );
  XOR U14341 ( .A(n14369), .B(n14382), .Z(n14381) );
  AND U14342 ( .A(n15691), .B(n15692), .Z(n14382) );
  XOR U14343 ( .A(n14371), .B(n14370), .Z(n14369) );
  AND U14344 ( .A(n15693), .B(n15694), .Z(n14370) );
  XOR U14345 ( .A(n14373), .B(n14372), .Z(n14371) );
  AND U14346 ( .A(n15695), .B(n15696), .Z(n14372) );
  XOR U14347 ( .A(n14375), .B(n14374), .Z(n14373) );
  AND U14348 ( .A(n15697), .B(n15698), .Z(n14374) );
  XOR U14349 ( .A(n14404), .B(n14376), .Z(n14375) );
  AND U14350 ( .A(n15699), .B(n15700), .Z(n14376) );
  XOR U14351 ( .A(n14400), .B(n14405), .Z(n14404) );
  AND U14352 ( .A(n15701), .B(n15702), .Z(n14405) );
  XOR U14353 ( .A(n14402), .B(n14401), .Z(n14400) );
  AND U14354 ( .A(n15703), .B(n15704), .Z(n14401) );
  XOR U14355 ( .A(n14390), .B(n14403), .Z(n14402) );
  AND U14356 ( .A(n15705), .B(n15706), .Z(n14403) );
  XOR U14357 ( .A(n14392), .B(n14391), .Z(n14390) );
  AND U14358 ( .A(n15707), .B(n15708), .Z(n14391) );
  XOR U14359 ( .A(n14394), .B(n14393), .Z(n14392) );
  AND U14360 ( .A(n15709), .B(n15710), .Z(n14393) );
  XOR U14361 ( .A(n14396), .B(n14395), .Z(n14394) );
  AND U14362 ( .A(n15711), .B(n15712), .Z(n14395) );
  XOR U14363 ( .A(n14438), .B(n14397), .Z(n14396) );
  AND U14364 ( .A(n15713), .B(n15714), .Z(n14397) );
  XNOR U14365 ( .A(n14435), .B(n14439), .Z(n14438) );
  AND U14366 ( .A(n15715), .B(n15716), .Z(n14439) );
  XOR U14367 ( .A(n14434), .B(n14426), .Z(n14435) );
  AND U14368 ( .A(n15717), .B(n15718), .Z(n14426) );
  XNOR U14369 ( .A(n14429), .B(n14425), .Z(n14434) );
  AND U14370 ( .A(n15719), .B(n15720), .Z(n14425) );
  XOR U14371 ( .A(n14442), .B(n14430), .Z(n14429) );
  AND U14372 ( .A(n15721), .B(n15722), .Z(n14430) );
  XNOR U14373 ( .A(n14422), .B(n14443), .Z(n14442) );
  AND U14374 ( .A(n15723), .B(n15724), .Z(n14443) );
  XOR U14375 ( .A(n14421), .B(n14413), .Z(n14422) );
  AND U14376 ( .A(n15725), .B(n15726), .Z(n14413) );
  XNOR U14377 ( .A(n14416), .B(n14412), .Z(n14421) );
  AND U14378 ( .A(n15727), .B(n15728), .Z(n14412) );
  XOR U14379 ( .A(n15729), .B(n15730), .Z(n14416) );
  XOR U14380 ( .A(n15731), .B(n15732), .Z(n15730) );
  XOR U14381 ( .A(n15733), .B(n15734), .Z(n15732) );
  XNOR U14382 ( .A(n14459), .B(n14452), .Z(n15734) );
  XOR U14383 ( .A(n15735), .B(n15736), .Z(n14452) );
  XOR U14384 ( .A(n15737), .B(n15738), .Z(n15736) );
  NOR U14385 ( .A(n15739), .B(n15740), .Z(n15738) );
  NOR U14386 ( .A(n15741), .B(n15742), .Z(n15737) );
  AND U14387 ( .A(n15743), .B(n15744), .Z(n15742) );
  IV U14388 ( .A(n15745), .Z(n15741) );
  NOR U14389 ( .A(n15746), .B(n15747), .Z(n15745) );
  AND U14390 ( .A(n15739), .B(n15748), .Z(n15747) );
  AND U14391 ( .A(n15740), .B(n15749), .Z(n15746) );
  XNOR U14392 ( .A(n15750), .B(n15751), .Z(n15735) );
  AND U14393 ( .A(n15752), .B(n15753), .Z(n15751) );
  AND U14394 ( .A(n15754), .B(n15755), .Z(n15750) );
  NOR U14395 ( .A(n15756), .B(n15757), .Z(n15755) );
  IV U14396 ( .A(n15758), .Z(n15756) );
  NOR U14397 ( .A(n15759), .B(n15760), .Z(n15758) );
  NOR U14398 ( .A(n15761), .B(n15762), .Z(n15754) );
  AND U14399 ( .A(n15763), .B(n15764), .Z(n14459) );
  XOR U14400 ( .A(n14457), .B(n14458), .Z(n15733) );
  AND U14401 ( .A(n15765), .B(n15766), .Z(n14458) );
  AND U14402 ( .A(n15767), .B(n15768), .Z(n14457) );
  XOR U14403 ( .A(n15769), .B(n15770), .Z(n15731) );
  XOR U14404 ( .A(n14453), .B(n14454), .Z(n15770) );
  AND U14405 ( .A(n15771), .B(n15772), .Z(n14454) );
  AND U14406 ( .A(n15773), .B(n15774), .Z(n14453) );
  XOR U14407 ( .A(n14451), .B(n14449), .Z(n15769) );
  AND U14408 ( .A(n15775), .B(n15776), .Z(n14449) );
  AND U14409 ( .A(n15777), .B(n15778), .Z(n14451) );
  XNOR U14410 ( .A(n14460), .B(n14417), .Z(n15729) );
  AND U14411 ( .A(n15779), .B(n15780), .Z(n14417) );
  AND U14412 ( .A(n15781), .B(n15782), .Z(n14460) );
  XOR U14413 ( .A(n15783), .B(n15784), .Z(n14473) );
  AND U14414 ( .A(n15783), .B(n15785), .Z(n15784) );
  XNOR U14415 ( .A(n15786), .B(n15787), .Z(n14476) );
  AND U14416 ( .A(n15786), .B(n15788), .Z(n15787) );
  XNOR U14417 ( .A(n15789), .B(n15790), .Z(n14479) );
  AND U14418 ( .A(n15789), .B(n15791), .Z(n15790) );
  XNOR U14419 ( .A(n15792), .B(n15793), .Z(n14482) );
  AND U14420 ( .A(n15792), .B(n15794), .Z(n15793) );
  XNOR U14421 ( .A(n15795), .B(n15796), .Z(n14485) );
  AND U14422 ( .A(n15797), .B(n15795), .Z(n15796) );
  XOR U14423 ( .A(n15798), .B(n15799), .Z(n14488) );
  NOR U14424 ( .A(n15800), .B(n15798), .Z(n15799) );
  XOR U14425 ( .A(n15801), .B(n15802), .Z(n14491) );
  NOR U14426 ( .A(n15803), .B(n15801), .Z(n15802) );
  XOR U14427 ( .A(n15804), .B(n15805), .Z(n14494) );
  NOR U14428 ( .A(n15806), .B(n15804), .Z(n15805) );
  XOR U14429 ( .A(n15807), .B(n15808), .Z(n14497) );
  NOR U14430 ( .A(n15809), .B(n15807), .Z(n15808) );
  XOR U14431 ( .A(n15810), .B(n15811), .Z(n14500) );
  NOR U14432 ( .A(n15812), .B(n15810), .Z(n15811) );
  XOR U14433 ( .A(n15813), .B(n15814), .Z(n14503) );
  NOR U14434 ( .A(n15815), .B(n15813), .Z(n15814) );
  XOR U14435 ( .A(n15816), .B(n15817), .Z(n14506) );
  NOR U14436 ( .A(n15818), .B(n15816), .Z(n15817) );
  XOR U14437 ( .A(n15819), .B(n15820), .Z(n14509) );
  NOR U14438 ( .A(n15821), .B(n15819), .Z(n15820) );
  XOR U14439 ( .A(n15822), .B(n15823), .Z(n14512) );
  NOR U14440 ( .A(n15824), .B(n15822), .Z(n15823) );
  XOR U14441 ( .A(n15825), .B(n15826), .Z(n14515) );
  NOR U14442 ( .A(n15827), .B(n15825), .Z(n15826) );
  XOR U14443 ( .A(n15828), .B(n15829), .Z(n14518) );
  NOR U14444 ( .A(n15830), .B(n15828), .Z(n15829) );
  XOR U14445 ( .A(n15831), .B(n15832), .Z(n14521) );
  NOR U14446 ( .A(n15833), .B(n15831), .Z(n15832) );
  XOR U14447 ( .A(n15834), .B(n15835), .Z(n14524) );
  NOR U14448 ( .A(n15836), .B(n15834), .Z(n15835) );
  XOR U14449 ( .A(n15837), .B(n15838), .Z(n14527) );
  NOR U14450 ( .A(n15839), .B(n15837), .Z(n15838) );
  XOR U14451 ( .A(n15840), .B(n15841), .Z(n14530) );
  NOR U14452 ( .A(n15842), .B(n15840), .Z(n15841) );
  XOR U14453 ( .A(n15843), .B(n15844), .Z(n14533) );
  NOR U14454 ( .A(n15845), .B(n15843), .Z(n15844) );
  XOR U14455 ( .A(n15846), .B(n15847), .Z(n14536) );
  NOR U14456 ( .A(n15848), .B(n15846), .Z(n15847) );
  XOR U14457 ( .A(n15849), .B(n15850), .Z(n14539) );
  NOR U14458 ( .A(n15851), .B(n15849), .Z(n15850) );
  XOR U14459 ( .A(n15852), .B(n15853), .Z(n14542) );
  NOR U14460 ( .A(n15854), .B(n15852), .Z(n15853) );
  XOR U14461 ( .A(n15855), .B(n15856), .Z(n14545) );
  NOR U14462 ( .A(n15857), .B(n15855), .Z(n15856) );
  XOR U14463 ( .A(n15858), .B(n15859), .Z(n14548) );
  NOR U14464 ( .A(n15860), .B(n15858), .Z(n15859) );
  XOR U14465 ( .A(n15861), .B(n15862), .Z(n14551) );
  NOR U14466 ( .A(n15863), .B(n15861), .Z(n15862) );
  XOR U14467 ( .A(n15864), .B(n15865), .Z(n14554) );
  NOR U14468 ( .A(n15866), .B(n15864), .Z(n15865) );
  XOR U14469 ( .A(n15867), .B(n15868), .Z(n14557) );
  NOR U14470 ( .A(n15869), .B(n15867), .Z(n15868) );
  XOR U14471 ( .A(n15870), .B(n15871), .Z(n14560) );
  NOR U14472 ( .A(n15872), .B(n15870), .Z(n15871) );
  XOR U14473 ( .A(n15873), .B(n15874), .Z(n14563) );
  NOR U14474 ( .A(n15875), .B(n15873), .Z(n15874) );
  XOR U14475 ( .A(n15876), .B(n15877), .Z(n14566) );
  NOR U14476 ( .A(n15878), .B(n15876), .Z(n15877) );
  XOR U14477 ( .A(n15879), .B(n15880), .Z(n14569) );
  NOR U14478 ( .A(n15881), .B(n15879), .Z(n15880) );
  XOR U14479 ( .A(n15882), .B(n15883), .Z(n14572) );
  NOR U14480 ( .A(n15884), .B(n15882), .Z(n15883) );
  XOR U14481 ( .A(n15885), .B(n15886), .Z(n14575) );
  NOR U14482 ( .A(n15887), .B(n15885), .Z(n15886) );
  XOR U14483 ( .A(n15888), .B(n15889), .Z(n14578) );
  NOR U14484 ( .A(n15890), .B(n15888), .Z(n15889) );
  XOR U14485 ( .A(n15891), .B(n15892), .Z(n14581) );
  NOR U14486 ( .A(n15893), .B(n15891), .Z(n15892) );
  XOR U14487 ( .A(n15894), .B(n15895), .Z(n14584) );
  NOR U14488 ( .A(n15896), .B(n15894), .Z(n15895) );
  XOR U14489 ( .A(n15897), .B(n15898), .Z(n14587) );
  NOR U14490 ( .A(n15899), .B(n15897), .Z(n15898) );
  XOR U14491 ( .A(n15900), .B(n15901), .Z(n14590) );
  NOR U14492 ( .A(n15902), .B(n15900), .Z(n15901) );
  XOR U14493 ( .A(n15903), .B(n15904), .Z(n14593) );
  NOR U14494 ( .A(n15905), .B(n15903), .Z(n15904) );
  XOR U14495 ( .A(n15906), .B(n15907), .Z(n14596) );
  NOR U14496 ( .A(n15908), .B(n15906), .Z(n15907) );
  XOR U14497 ( .A(n15909), .B(n15910), .Z(n14599) );
  NOR U14498 ( .A(n15911), .B(n15909), .Z(n15910) );
  XOR U14499 ( .A(n15912), .B(n15913), .Z(n14602) );
  NOR U14500 ( .A(n15914), .B(n15912), .Z(n15913) );
  XOR U14501 ( .A(n15915), .B(n15916), .Z(n14605) );
  NOR U14502 ( .A(n15917), .B(n15915), .Z(n15916) );
  XOR U14503 ( .A(n15918), .B(n15919), .Z(n14608) );
  NOR U14504 ( .A(n15920), .B(n15918), .Z(n15919) );
  XOR U14505 ( .A(n15921), .B(n15922), .Z(n14611) );
  NOR U14506 ( .A(n15923), .B(n15921), .Z(n15922) );
  XOR U14507 ( .A(n15924), .B(n15925), .Z(n14614) );
  NOR U14508 ( .A(n15926), .B(n15924), .Z(n15925) );
  XOR U14509 ( .A(n15927), .B(n15928), .Z(n14617) );
  NOR U14510 ( .A(n15929), .B(n15927), .Z(n15928) );
  XOR U14511 ( .A(n15930), .B(n15931), .Z(n14620) );
  NOR U14512 ( .A(n15932), .B(n15930), .Z(n15931) );
  XOR U14513 ( .A(n15933), .B(n15934), .Z(n14623) );
  NOR U14514 ( .A(n15935), .B(n15933), .Z(n15934) );
  XOR U14515 ( .A(n15936), .B(n15937), .Z(n14626) );
  NOR U14516 ( .A(n15938), .B(n15936), .Z(n15937) );
  XOR U14517 ( .A(n15939), .B(n15940), .Z(n14629) );
  NOR U14518 ( .A(n15941), .B(n15939), .Z(n15940) );
  XOR U14519 ( .A(n15942), .B(n15943), .Z(n14632) );
  NOR U14520 ( .A(n15944), .B(n15942), .Z(n15943) );
  XOR U14521 ( .A(n15945), .B(n15946), .Z(n14635) );
  NOR U14522 ( .A(n15947), .B(n15945), .Z(n15946) );
  XOR U14523 ( .A(n15948), .B(n15949), .Z(n14638) );
  NOR U14524 ( .A(n15950), .B(n15948), .Z(n15949) );
  XOR U14525 ( .A(n15951), .B(n15952), .Z(n14641) );
  NOR U14526 ( .A(n15953), .B(n15951), .Z(n15952) );
  XOR U14527 ( .A(n15954), .B(n15955), .Z(n14644) );
  NOR U14528 ( .A(n15956), .B(n15954), .Z(n15955) );
  XOR U14529 ( .A(n15957), .B(n15958), .Z(n14647) );
  NOR U14530 ( .A(n15959), .B(n15957), .Z(n15958) );
  XOR U14531 ( .A(n15960), .B(n15961), .Z(n14650) );
  NOR U14532 ( .A(n15962), .B(n15960), .Z(n15961) );
  XOR U14533 ( .A(n15963), .B(n15964), .Z(n14653) );
  NOR U14534 ( .A(n15965), .B(n15963), .Z(n15964) );
  XOR U14535 ( .A(n15966), .B(n15967), .Z(n14656) );
  NOR U14536 ( .A(n15968), .B(n15966), .Z(n15967) );
  XOR U14537 ( .A(n15969), .B(n15970), .Z(n14659) );
  NOR U14538 ( .A(n15971), .B(n15969), .Z(n15970) );
  XOR U14539 ( .A(n15972), .B(n15973), .Z(n14662) );
  NOR U14540 ( .A(n15974), .B(n15972), .Z(n15973) );
  XOR U14541 ( .A(n15975), .B(n15976), .Z(n14665) );
  NOR U14542 ( .A(n15977), .B(n15975), .Z(n15976) );
  XOR U14543 ( .A(n15978), .B(n15979), .Z(n14668) );
  NOR U14544 ( .A(n15980), .B(n15978), .Z(n15979) );
  XOR U14545 ( .A(n15981), .B(n15982), .Z(n14671) );
  NOR U14546 ( .A(n15983), .B(n15981), .Z(n15982) );
  XOR U14547 ( .A(n15984), .B(n15985), .Z(n14674) );
  NOR U14548 ( .A(n15986), .B(n15984), .Z(n15985) );
  XOR U14549 ( .A(n15987), .B(n15988), .Z(n14677) );
  NOR U14550 ( .A(n15989), .B(n15987), .Z(n15988) );
  XOR U14551 ( .A(n15990), .B(n15991), .Z(n14680) );
  NOR U14552 ( .A(n15992), .B(n15990), .Z(n15991) );
  XOR U14553 ( .A(n15993), .B(n15994), .Z(n14683) );
  NOR U14554 ( .A(n15995), .B(n15993), .Z(n15994) );
  XOR U14555 ( .A(n15996), .B(n15997), .Z(n14686) );
  NOR U14556 ( .A(n15998), .B(n15996), .Z(n15997) );
  XOR U14557 ( .A(n15999), .B(n16000), .Z(n14689) );
  NOR U14558 ( .A(n16001), .B(n15999), .Z(n16000) );
  XOR U14559 ( .A(n16002), .B(n16003), .Z(n14692) );
  NOR U14560 ( .A(n16004), .B(n16002), .Z(n16003) );
  XOR U14561 ( .A(n16005), .B(n16006), .Z(n14695) );
  NOR U14562 ( .A(n16007), .B(n16005), .Z(n16006) );
  XOR U14563 ( .A(n16008), .B(n16009), .Z(n14698) );
  NOR U14564 ( .A(n16010), .B(n16008), .Z(n16009) );
  XOR U14565 ( .A(n16011), .B(n16012), .Z(n14701) );
  NOR U14566 ( .A(n16013), .B(n16011), .Z(n16012) );
  XOR U14567 ( .A(n16014), .B(n16015), .Z(n14704) );
  NOR U14568 ( .A(n16016), .B(n16014), .Z(n16015) );
  XOR U14569 ( .A(n16017), .B(n16018), .Z(n14707) );
  NOR U14570 ( .A(n16019), .B(n16017), .Z(n16018) );
  XOR U14571 ( .A(n16020), .B(n16021), .Z(n14710) );
  NOR U14572 ( .A(n16022), .B(n16020), .Z(n16021) );
  XOR U14573 ( .A(n16023), .B(n16024), .Z(n14713) );
  NOR U14574 ( .A(n16025), .B(n16023), .Z(n16024) );
  XOR U14575 ( .A(n16026), .B(n16027), .Z(n14716) );
  NOR U14576 ( .A(n16028), .B(n16026), .Z(n16027) );
  XOR U14577 ( .A(n16029), .B(n16030), .Z(n14719) );
  NOR U14578 ( .A(n16031), .B(n16029), .Z(n16030) );
  XOR U14579 ( .A(n16032), .B(n16033), .Z(n14722) );
  NOR U14580 ( .A(n16034), .B(n16032), .Z(n16033) );
  XOR U14581 ( .A(n16035), .B(n16036), .Z(n14725) );
  NOR U14582 ( .A(n16037), .B(n16035), .Z(n16036) );
  XOR U14583 ( .A(n16038), .B(n16039), .Z(n14728) );
  NOR U14584 ( .A(n16040), .B(n16038), .Z(n16039) );
  XOR U14585 ( .A(n16041), .B(n16042), .Z(n14731) );
  NOR U14586 ( .A(n16043), .B(n16041), .Z(n16042) );
  XOR U14587 ( .A(n16044), .B(n16045), .Z(n14734) );
  NOR U14588 ( .A(n16046), .B(n16044), .Z(n16045) );
  XOR U14589 ( .A(n16047), .B(n16048), .Z(n14737) );
  NOR U14590 ( .A(n16049), .B(n16047), .Z(n16048) );
  XOR U14591 ( .A(n16050), .B(n16051), .Z(n14740) );
  NOR U14592 ( .A(n16052), .B(n16050), .Z(n16051) );
  XOR U14593 ( .A(n16053), .B(n16054), .Z(n14743) );
  NOR U14594 ( .A(n16055), .B(n16053), .Z(n16054) );
  XOR U14595 ( .A(n16056), .B(n16057), .Z(n14746) );
  NOR U14596 ( .A(n16058), .B(n16056), .Z(n16057) );
  XOR U14597 ( .A(n16059), .B(n16060), .Z(n14749) );
  NOR U14598 ( .A(n16061), .B(n16059), .Z(n16060) );
  XOR U14599 ( .A(n16062), .B(n16063), .Z(n14752) );
  NOR U14600 ( .A(n16064), .B(n16062), .Z(n16063) );
  XOR U14601 ( .A(n16065), .B(n16066), .Z(n14755) );
  NOR U14602 ( .A(n16067), .B(n16065), .Z(n16066) );
  XOR U14603 ( .A(n16068), .B(n16069), .Z(n14758) );
  NOR U14604 ( .A(n16070), .B(n16068), .Z(n16069) );
  XOR U14605 ( .A(n16071), .B(n16072), .Z(n14761) );
  NOR U14606 ( .A(n16073), .B(n16071), .Z(n16072) );
  XOR U14607 ( .A(n16074), .B(n16075), .Z(n14764) );
  NOR U14608 ( .A(n16076), .B(n16074), .Z(n16075) );
  XOR U14609 ( .A(n16077), .B(n16078), .Z(n14767) );
  NOR U14610 ( .A(n16079), .B(n16077), .Z(n16078) );
  XOR U14611 ( .A(n16080), .B(n16081), .Z(n14770) );
  NOR U14612 ( .A(n16082), .B(n16080), .Z(n16081) );
  XOR U14613 ( .A(n16083), .B(n16084), .Z(n14773) );
  NOR U14614 ( .A(n16085), .B(n16083), .Z(n16084) );
  XOR U14615 ( .A(n16086), .B(n16087), .Z(n14776) );
  NOR U14616 ( .A(n16088), .B(n16086), .Z(n16087) );
  XOR U14617 ( .A(n16089), .B(n16090), .Z(n14779) );
  NOR U14618 ( .A(n16091), .B(n16089), .Z(n16090) );
  XOR U14619 ( .A(n16092), .B(n16093), .Z(n14782) );
  NOR U14620 ( .A(n16094), .B(n16092), .Z(n16093) );
  XOR U14621 ( .A(n16095), .B(n16096), .Z(n14785) );
  NOR U14622 ( .A(n16097), .B(n16095), .Z(n16096) );
  XOR U14623 ( .A(n16098), .B(n16099), .Z(n14788) );
  NOR U14624 ( .A(n16100), .B(n16098), .Z(n16099) );
  XOR U14625 ( .A(n16101), .B(n16102), .Z(n14791) );
  NOR U14626 ( .A(n16103), .B(n16101), .Z(n16102) );
  XOR U14627 ( .A(n16104), .B(n16105), .Z(n14794) );
  NOR U14628 ( .A(n16106), .B(n16104), .Z(n16105) );
  XOR U14629 ( .A(n16107), .B(n16108), .Z(n14797) );
  NOR U14630 ( .A(n16109), .B(n16107), .Z(n16108) );
  XOR U14631 ( .A(n16110), .B(n16111), .Z(n14800) );
  NOR U14632 ( .A(n16112), .B(n16110), .Z(n16111) );
  XOR U14633 ( .A(n16113), .B(n16114), .Z(n14803) );
  NOR U14634 ( .A(n16115), .B(n16113), .Z(n16114) );
  XOR U14635 ( .A(n16116), .B(n16117), .Z(n14806) );
  NOR U14636 ( .A(n16118), .B(n16116), .Z(n16117) );
  XOR U14637 ( .A(n16119), .B(n16120), .Z(n14809) );
  NOR U14638 ( .A(n16121), .B(n16119), .Z(n16120) );
  XOR U14639 ( .A(n16122), .B(n16123), .Z(n14812) );
  NOR U14640 ( .A(n16124), .B(n16122), .Z(n16123) );
  XOR U14641 ( .A(n16125), .B(n16126), .Z(n14815) );
  NOR U14642 ( .A(n16127), .B(n16125), .Z(n16126) );
  XOR U14643 ( .A(n16128), .B(n16129), .Z(n14818) );
  NOR U14644 ( .A(n16130), .B(n16128), .Z(n16129) );
  XOR U14645 ( .A(n16131), .B(n16132), .Z(n14821) );
  NOR U14646 ( .A(n16133), .B(n16131), .Z(n16132) );
  XOR U14647 ( .A(n16134), .B(n16135), .Z(n14824) );
  NOR U14648 ( .A(n16136), .B(n16134), .Z(n16135) );
  XOR U14649 ( .A(n16137), .B(n16138), .Z(n14827) );
  NOR U14650 ( .A(n16139), .B(n16137), .Z(n16138) );
  XOR U14651 ( .A(n16140), .B(n16141), .Z(n14830) );
  NOR U14652 ( .A(n16142), .B(n16140), .Z(n16141) );
  XOR U14653 ( .A(n16143), .B(n16144), .Z(n14833) );
  NOR U14654 ( .A(n16145), .B(n16143), .Z(n16144) );
  XOR U14655 ( .A(n16146), .B(n16147), .Z(n14836) );
  NOR U14656 ( .A(n16148), .B(n16146), .Z(n16147) );
  XOR U14657 ( .A(n16149), .B(n16150), .Z(n14839) );
  NOR U14658 ( .A(n16151), .B(n16149), .Z(n16150) );
  XOR U14659 ( .A(n16152), .B(n16153), .Z(n14842) );
  NOR U14660 ( .A(n16154), .B(n16152), .Z(n16153) );
  XOR U14661 ( .A(n16155), .B(n16156), .Z(n14845) );
  NOR U14662 ( .A(n16157), .B(n16155), .Z(n16156) );
  XOR U14663 ( .A(n16158), .B(n16159), .Z(n14848) );
  NOR U14664 ( .A(n16160), .B(n16158), .Z(n16159) );
  XOR U14665 ( .A(n16161), .B(n16162), .Z(n14851) );
  NOR U14666 ( .A(n16163), .B(n16161), .Z(n16162) );
  XOR U14667 ( .A(n16164), .B(n16165), .Z(n14854) );
  NOR U14668 ( .A(n16166), .B(n16164), .Z(n16165) );
  XOR U14669 ( .A(n16167), .B(n16168), .Z(n14857) );
  NOR U14670 ( .A(n16169), .B(n16167), .Z(n16168) );
  XOR U14671 ( .A(n16170), .B(n16171), .Z(n14860) );
  NOR U14672 ( .A(n16172), .B(n16170), .Z(n16171) );
  XOR U14673 ( .A(n16173), .B(n16174), .Z(n14863) );
  NOR U14674 ( .A(n16175), .B(n16173), .Z(n16174) );
  XOR U14675 ( .A(n16176), .B(n16177), .Z(n14866) );
  NOR U14676 ( .A(n16178), .B(n16176), .Z(n16177) );
  XOR U14677 ( .A(n16179), .B(n16180), .Z(n14869) );
  NOR U14678 ( .A(n16181), .B(n16179), .Z(n16180) );
  XOR U14679 ( .A(n16182), .B(n16183), .Z(n14872) );
  NOR U14680 ( .A(n16184), .B(n16182), .Z(n16183) );
  XOR U14681 ( .A(n16185), .B(n16186), .Z(n14875) );
  NOR U14682 ( .A(n105), .B(n16187), .Z(n16186) );
  XOR U14683 ( .A(n16188), .B(n16189), .Z(n14878) );
  AND U14684 ( .A(n16190), .B(n16191), .Z(n16189) );
  XOR U14685 ( .A(n16188), .B(n108), .Z(n16191) );
  XNOR U14686 ( .A(n15533), .B(n15532), .Z(n108) );
  XNOR U14687 ( .A(n15530), .B(n15529), .Z(n15532) );
  XNOR U14688 ( .A(n15527), .B(n15526), .Z(n15529) );
  XNOR U14689 ( .A(n15524), .B(n15523), .Z(n15526) );
  XNOR U14690 ( .A(n15521), .B(n15520), .Z(n15523) );
  XNOR U14691 ( .A(n15518), .B(n15517), .Z(n15520) );
  XNOR U14692 ( .A(n15515), .B(n15514), .Z(n15517) );
  XNOR U14693 ( .A(n15512), .B(n15511), .Z(n15514) );
  XNOR U14694 ( .A(n15509), .B(n15508), .Z(n15511) );
  XNOR U14695 ( .A(n15506), .B(n15505), .Z(n15508) );
  XNOR U14696 ( .A(n15503), .B(n15502), .Z(n15505) );
  XNOR U14697 ( .A(n15500), .B(n15499), .Z(n15502) );
  XNOR U14698 ( .A(n15497), .B(n15496), .Z(n15499) );
  XNOR U14699 ( .A(n15494), .B(n15493), .Z(n15496) );
  XNOR U14700 ( .A(n15491), .B(n15490), .Z(n15493) );
  XNOR U14701 ( .A(n15488), .B(n15487), .Z(n15490) );
  XNOR U14702 ( .A(n15485), .B(n15484), .Z(n15487) );
  XNOR U14703 ( .A(n15482), .B(n15481), .Z(n15484) );
  XNOR U14704 ( .A(n15479), .B(n15478), .Z(n15481) );
  XNOR U14705 ( .A(n15476), .B(n15475), .Z(n15478) );
  XNOR U14706 ( .A(n15473), .B(n15472), .Z(n15475) );
  XNOR U14707 ( .A(n15470), .B(n15469), .Z(n15472) );
  XNOR U14708 ( .A(n15467), .B(n15466), .Z(n15469) );
  XNOR U14709 ( .A(n15464), .B(n15463), .Z(n15466) );
  XNOR U14710 ( .A(n15461), .B(n15460), .Z(n15463) );
  XNOR U14711 ( .A(n15458), .B(n15457), .Z(n15460) );
  XNOR U14712 ( .A(n15455), .B(n15454), .Z(n15457) );
  XNOR U14713 ( .A(n15452), .B(n15451), .Z(n15454) );
  XNOR U14714 ( .A(n15449), .B(n15448), .Z(n15451) );
  XNOR U14715 ( .A(n15446), .B(n15445), .Z(n15448) );
  XNOR U14716 ( .A(n15443), .B(n15442), .Z(n15445) );
  XNOR U14717 ( .A(n15440), .B(n15439), .Z(n15442) );
  XNOR U14718 ( .A(n15437), .B(n15436), .Z(n15439) );
  XNOR U14719 ( .A(n15434), .B(n15433), .Z(n15436) );
  XNOR U14720 ( .A(n15431), .B(n15430), .Z(n15433) );
  XNOR U14721 ( .A(n15428), .B(n15427), .Z(n15430) );
  XNOR U14722 ( .A(n15425), .B(n15424), .Z(n15427) );
  XNOR U14723 ( .A(n15422), .B(n15421), .Z(n15424) );
  XNOR U14724 ( .A(n15419), .B(n15418), .Z(n15421) );
  XNOR U14725 ( .A(n15416), .B(n15415), .Z(n15418) );
  XNOR U14726 ( .A(n15413), .B(n15412), .Z(n15415) );
  XNOR U14727 ( .A(n15410), .B(n15409), .Z(n15412) );
  XNOR U14728 ( .A(n15407), .B(n15406), .Z(n15409) );
  XNOR U14729 ( .A(n15404), .B(n15403), .Z(n15406) );
  XNOR U14730 ( .A(n15401), .B(n15400), .Z(n15403) );
  XNOR U14731 ( .A(n15398), .B(n15397), .Z(n15400) );
  XNOR U14732 ( .A(n15395), .B(n15394), .Z(n15397) );
  XNOR U14733 ( .A(n15392), .B(n15391), .Z(n15394) );
  XNOR U14734 ( .A(n15389), .B(n15388), .Z(n15391) );
  XNOR U14735 ( .A(n15386), .B(n15385), .Z(n15388) );
  XNOR U14736 ( .A(n15383), .B(n15382), .Z(n15385) );
  XNOR U14737 ( .A(n15380), .B(n15379), .Z(n15382) );
  XNOR U14738 ( .A(n15377), .B(n15376), .Z(n15379) );
  XNOR U14739 ( .A(n15374), .B(n15373), .Z(n15376) );
  XNOR U14740 ( .A(n15371), .B(n15370), .Z(n15373) );
  XNOR U14741 ( .A(n15368), .B(n15367), .Z(n15370) );
  XNOR U14742 ( .A(n15365), .B(n15364), .Z(n15367) );
  XNOR U14743 ( .A(n15362), .B(n15361), .Z(n15364) );
  XNOR U14744 ( .A(n15359), .B(n15358), .Z(n15361) );
  XNOR U14745 ( .A(n15356), .B(n15355), .Z(n15358) );
  XNOR U14746 ( .A(n15353), .B(n15352), .Z(n15355) );
  XNOR U14747 ( .A(n15350), .B(n15349), .Z(n15352) );
  XNOR U14748 ( .A(n15347), .B(n15346), .Z(n15349) );
  XNOR U14749 ( .A(n15344), .B(n15343), .Z(n15346) );
  XNOR U14750 ( .A(n15341), .B(n15340), .Z(n15343) );
  XNOR U14751 ( .A(n15338), .B(n15337), .Z(n15340) );
  XNOR U14752 ( .A(n15335), .B(n15334), .Z(n15337) );
  XNOR U14753 ( .A(n15332), .B(n15331), .Z(n15334) );
  XNOR U14754 ( .A(n15329), .B(n15328), .Z(n15331) );
  XNOR U14755 ( .A(n15326), .B(n15325), .Z(n15328) );
  XNOR U14756 ( .A(n15323), .B(n15322), .Z(n15325) );
  XNOR U14757 ( .A(n15320), .B(n15319), .Z(n15322) );
  XNOR U14758 ( .A(n15317), .B(n15316), .Z(n15319) );
  XNOR U14759 ( .A(n15314), .B(n15313), .Z(n15316) );
  XNOR U14760 ( .A(n15311), .B(n15310), .Z(n15313) );
  XNOR U14761 ( .A(n15308), .B(n15307), .Z(n15310) );
  XNOR U14762 ( .A(n15305), .B(n15304), .Z(n15307) );
  XNOR U14763 ( .A(n15302), .B(n15301), .Z(n15304) );
  XNOR U14764 ( .A(n15299), .B(n15298), .Z(n15301) );
  XNOR U14765 ( .A(n15296), .B(n15295), .Z(n15298) );
  XNOR U14766 ( .A(n15293), .B(n15292), .Z(n15295) );
  XNOR U14767 ( .A(n15290), .B(n15289), .Z(n15292) );
  XNOR U14768 ( .A(n15287), .B(n15286), .Z(n15289) );
  XNOR U14769 ( .A(n15284), .B(n15283), .Z(n15286) );
  XNOR U14770 ( .A(n15281), .B(n15280), .Z(n15283) );
  XNOR U14771 ( .A(n15278), .B(n15277), .Z(n15280) );
  XNOR U14772 ( .A(n15275), .B(n15274), .Z(n15277) );
  XNOR U14773 ( .A(n15272), .B(n15271), .Z(n15274) );
  XNOR U14774 ( .A(n15269), .B(n15268), .Z(n15271) );
  XNOR U14775 ( .A(n15266), .B(n15265), .Z(n15268) );
  XNOR U14776 ( .A(n15263), .B(n15262), .Z(n15265) );
  XNOR U14777 ( .A(n15260), .B(n15259), .Z(n15262) );
  XNOR U14778 ( .A(n15257), .B(n15256), .Z(n15259) );
  XNOR U14779 ( .A(n15254), .B(n15253), .Z(n15256) );
  XNOR U14780 ( .A(n15251), .B(n15250), .Z(n15253) );
  XNOR U14781 ( .A(n15248), .B(n15247), .Z(n15250) );
  XNOR U14782 ( .A(n15245), .B(n15244), .Z(n15247) );
  XNOR U14783 ( .A(n15242), .B(n15241), .Z(n15244) );
  XNOR U14784 ( .A(n15239), .B(n15238), .Z(n15241) );
  XNOR U14785 ( .A(n15236), .B(n15235), .Z(n15238) );
  XNOR U14786 ( .A(n15233), .B(n15232), .Z(n15235) );
  XNOR U14787 ( .A(n15230), .B(n15229), .Z(n15232) );
  XNOR U14788 ( .A(n15227), .B(n15226), .Z(n15229) );
  XNOR U14789 ( .A(n15224), .B(n15223), .Z(n15226) );
  XNOR U14790 ( .A(n15221), .B(n15220), .Z(n15223) );
  XNOR U14791 ( .A(n15218), .B(n15217), .Z(n15220) );
  XNOR U14792 ( .A(n15215), .B(n15214), .Z(n15217) );
  XNOR U14793 ( .A(n15212), .B(n15211), .Z(n15214) );
  XNOR U14794 ( .A(n15209), .B(n15208), .Z(n15211) );
  XNOR U14795 ( .A(n15206), .B(n15205), .Z(n15208) );
  XNOR U14796 ( .A(n15203), .B(n15202), .Z(n15205) );
  XNOR U14797 ( .A(n15200), .B(n15199), .Z(n15202) );
  XNOR U14798 ( .A(n15197), .B(n15196), .Z(n15199) );
  XNOR U14799 ( .A(n15194), .B(n15193), .Z(n15196) );
  XNOR U14800 ( .A(n15191), .B(n15190), .Z(n15193) );
  XNOR U14801 ( .A(n15188), .B(n15187), .Z(n15190) );
  XNOR U14802 ( .A(n15185), .B(n15184), .Z(n15187) );
  XNOR U14803 ( .A(n15182), .B(n15181), .Z(n15184) );
  XNOR U14804 ( .A(n15179), .B(n15178), .Z(n15181) );
  XNOR U14805 ( .A(n15176), .B(n15175), .Z(n15178) );
  XNOR U14806 ( .A(n15173), .B(n15172), .Z(n15175) );
  XNOR U14807 ( .A(n15170), .B(n15169), .Z(n15172) );
  XNOR U14808 ( .A(n15167), .B(n15166), .Z(n15169) );
  XNOR U14809 ( .A(n15164), .B(n15163), .Z(n15166) );
  XNOR U14810 ( .A(n15161), .B(n15160), .Z(n15163) );
  XNOR U14811 ( .A(n15158), .B(n15157), .Z(n15160) );
  XNOR U14812 ( .A(n15155), .B(n15154), .Z(n15157) );
  XNOR U14813 ( .A(n15152), .B(n15151), .Z(n15154) );
  XNOR U14814 ( .A(n15149), .B(n15148), .Z(n15151) );
  XOR U14815 ( .A(n15146), .B(n15145), .Z(n15148) );
  XOR U14816 ( .A(n15143), .B(n15142), .Z(n15145) );
  XOR U14817 ( .A(n15139), .B(n15140), .Z(n15142) );
  AND U14818 ( .A(n16192), .B(n16193), .Z(n15140) );
  XOR U14819 ( .A(n15136), .B(n15137), .Z(n15139) );
  AND U14820 ( .A(n16194), .B(n16195), .Z(n15137) );
  XOR U14821 ( .A(n15133), .B(n15134), .Z(n15136) );
  AND U14822 ( .A(n16196), .B(n16197), .Z(n15134) );
  XNOR U14823 ( .A(n14882), .B(n15131), .Z(n15133) );
  AND U14824 ( .A(n16198), .B(n16199), .Z(n15131) );
  XOR U14825 ( .A(n14884), .B(n14883), .Z(n14882) );
  AND U14826 ( .A(n16200), .B(n16201), .Z(n14883) );
  XOR U14827 ( .A(n14886), .B(n14885), .Z(n14884) );
  AND U14828 ( .A(n16202), .B(n16203), .Z(n14885) );
  XOR U14829 ( .A(n14888), .B(n14887), .Z(n14886) );
  AND U14830 ( .A(n16204), .B(n16205), .Z(n14887) );
  XOR U14831 ( .A(n14890), .B(n14889), .Z(n14888) );
  AND U14832 ( .A(n16206), .B(n16207), .Z(n14889) );
  XOR U14833 ( .A(n14892), .B(n14891), .Z(n14890) );
  AND U14834 ( .A(n16208), .B(n16209), .Z(n14891) );
  XOR U14835 ( .A(n14894), .B(n14893), .Z(n14892) );
  AND U14836 ( .A(n16210), .B(n16211), .Z(n14893) );
  XOR U14837 ( .A(n14896), .B(n14895), .Z(n14894) );
  AND U14838 ( .A(n16212), .B(n16213), .Z(n14895) );
  XOR U14839 ( .A(n14898), .B(n14897), .Z(n14896) );
  AND U14840 ( .A(n16214), .B(n16215), .Z(n14897) );
  XOR U14841 ( .A(n14900), .B(n14899), .Z(n14898) );
  AND U14842 ( .A(n16216), .B(n16217), .Z(n14899) );
  XOR U14843 ( .A(n14902), .B(n14901), .Z(n14900) );
  AND U14844 ( .A(n16218), .B(n16219), .Z(n14901) );
  XOR U14845 ( .A(n14904), .B(n14903), .Z(n14902) );
  AND U14846 ( .A(n16220), .B(n16221), .Z(n14903) );
  XOR U14847 ( .A(n14906), .B(n14905), .Z(n14904) );
  AND U14848 ( .A(n16222), .B(n16223), .Z(n14905) );
  XOR U14849 ( .A(n14908), .B(n14907), .Z(n14906) );
  AND U14850 ( .A(n16224), .B(n16225), .Z(n14907) );
  XOR U14851 ( .A(n14910), .B(n14909), .Z(n14908) );
  AND U14852 ( .A(n16226), .B(n16227), .Z(n14909) );
  XOR U14853 ( .A(n14912), .B(n14911), .Z(n14910) );
  AND U14854 ( .A(n16228), .B(n16229), .Z(n14911) );
  XOR U14855 ( .A(n14914), .B(n14913), .Z(n14912) );
  AND U14856 ( .A(n16230), .B(n16231), .Z(n14913) );
  XOR U14857 ( .A(n14916), .B(n14915), .Z(n14914) );
  AND U14858 ( .A(n16232), .B(n16233), .Z(n14915) );
  XOR U14859 ( .A(n14918), .B(n14917), .Z(n14916) );
  AND U14860 ( .A(n16234), .B(n16235), .Z(n14917) );
  XOR U14861 ( .A(n14920), .B(n14919), .Z(n14918) );
  AND U14862 ( .A(n16236), .B(n16237), .Z(n14919) );
  XOR U14863 ( .A(n14922), .B(n14921), .Z(n14920) );
  AND U14864 ( .A(n16238), .B(n16239), .Z(n14921) );
  XOR U14865 ( .A(n14924), .B(n14923), .Z(n14922) );
  AND U14866 ( .A(n16240), .B(n16241), .Z(n14923) );
  XOR U14867 ( .A(n14926), .B(n14925), .Z(n14924) );
  AND U14868 ( .A(n16242), .B(n16243), .Z(n14925) );
  XOR U14869 ( .A(n14928), .B(n14927), .Z(n14926) );
  AND U14870 ( .A(n16244), .B(n16245), .Z(n14927) );
  XOR U14871 ( .A(n14930), .B(n14929), .Z(n14928) );
  AND U14872 ( .A(n16246), .B(n16247), .Z(n14929) );
  XOR U14873 ( .A(n14932), .B(n14931), .Z(n14930) );
  AND U14874 ( .A(n16248), .B(n16249), .Z(n14931) );
  XOR U14875 ( .A(n14934), .B(n14933), .Z(n14932) );
  AND U14876 ( .A(n16250), .B(n16251), .Z(n14933) );
  XOR U14877 ( .A(n14936), .B(n14935), .Z(n14934) );
  AND U14878 ( .A(n16252), .B(n16253), .Z(n14935) );
  XOR U14879 ( .A(n14938), .B(n14937), .Z(n14936) );
  AND U14880 ( .A(n16254), .B(n16255), .Z(n14937) );
  XOR U14881 ( .A(n14940), .B(n14939), .Z(n14938) );
  AND U14882 ( .A(n16256), .B(n16257), .Z(n14939) );
  XOR U14883 ( .A(n14942), .B(n14941), .Z(n14940) );
  AND U14884 ( .A(n16258), .B(n16259), .Z(n14941) );
  XOR U14885 ( .A(n14944), .B(n14943), .Z(n14942) );
  AND U14886 ( .A(n16260), .B(n16261), .Z(n14943) );
  XOR U14887 ( .A(n14946), .B(n14945), .Z(n14944) );
  AND U14888 ( .A(n16262), .B(n16263), .Z(n14945) );
  XOR U14889 ( .A(n14948), .B(n14947), .Z(n14946) );
  AND U14890 ( .A(n16264), .B(n16265), .Z(n14947) );
  XOR U14891 ( .A(n14950), .B(n14949), .Z(n14948) );
  AND U14892 ( .A(n16266), .B(n16267), .Z(n14949) );
  XOR U14893 ( .A(n14952), .B(n14951), .Z(n14950) );
  AND U14894 ( .A(n16268), .B(n16269), .Z(n14951) );
  XOR U14895 ( .A(n14954), .B(n14953), .Z(n14952) );
  AND U14896 ( .A(n16270), .B(n16271), .Z(n14953) );
  XOR U14897 ( .A(n14956), .B(n14955), .Z(n14954) );
  AND U14898 ( .A(n16272), .B(n16273), .Z(n14955) );
  XOR U14899 ( .A(n14958), .B(n14957), .Z(n14956) );
  AND U14900 ( .A(n16274), .B(n16275), .Z(n14957) );
  XOR U14901 ( .A(n14960), .B(n14959), .Z(n14958) );
  AND U14902 ( .A(n16276), .B(n16277), .Z(n14959) );
  XOR U14903 ( .A(n14962), .B(n14961), .Z(n14960) );
  AND U14904 ( .A(n16278), .B(n16279), .Z(n14961) );
  XOR U14905 ( .A(n14964), .B(n14963), .Z(n14962) );
  AND U14906 ( .A(n16280), .B(n16281), .Z(n14963) );
  XOR U14907 ( .A(n14966), .B(n14965), .Z(n14964) );
  AND U14908 ( .A(n16282), .B(n16283), .Z(n14965) );
  XOR U14909 ( .A(n14968), .B(n14967), .Z(n14966) );
  AND U14910 ( .A(n16284), .B(n16285), .Z(n14967) );
  XOR U14911 ( .A(n14970), .B(n14969), .Z(n14968) );
  AND U14912 ( .A(n16286), .B(n16287), .Z(n14969) );
  XOR U14913 ( .A(n14972), .B(n14971), .Z(n14970) );
  AND U14914 ( .A(n16288), .B(n16289), .Z(n14971) );
  XOR U14915 ( .A(n14974), .B(n14973), .Z(n14972) );
  AND U14916 ( .A(n16290), .B(n16291), .Z(n14973) );
  XOR U14917 ( .A(n14976), .B(n14975), .Z(n14974) );
  AND U14918 ( .A(n16292), .B(n16293), .Z(n14975) );
  XOR U14919 ( .A(n14978), .B(n14977), .Z(n14976) );
  AND U14920 ( .A(n16294), .B(n16295), .Z(n14977) );
  XOR U14921 ( .A(n14980), .B(n14979), .Z(n14978) );
  AND U14922 ( .A(n16296), .B(n16297), .Z(n14979) );
  XOR U14923 ( .A(n14982), .B(n14981), .Z(n14980) );
  AND U14924 ( .A(n16298), .B(n16299), .Z(n14981) );
  XOR U14925 ( .A(n14984), .B(n14983), .Z(n14982) );
  AND U14926 ( .A(n16300), .B(n16301), .Z(n14983) );
  XOR U14927 ( .A(n14986), .B(n14985), .Z(n14984) );
  AND U14928 ( .A(n16302), .B(n16303), .Z(n14985) );
  XOR U14929 ( .A(n14988), .B(n14987), .Z(n14986) );
  AND U14930 ( .A(n16304), .B(n16305), .Z(n14987) );
  XOR U14931 ( .A(n14990), .B(n14989), .Z(n14988) );
  AND U14932 ( .A(n16306), .B(n16307), .Z(n14989) );
  XOR U14933 ( .A(n14992), .B(n14991), .Z(n14990) );
  AND U14934 ( .A(n16308), .B(n16309), .Z(n14991) );
  XOR U14935 ( .A(n14994), .B(n14993), .Z(n14992) );
  AND U14936 ( .A(n16310), .B(n16311), .Z(n14993) );
  XOR U14937 ( .A(n14996), .B(n14995), .Z(n14994) );
  AND U14938 ( .A(n16312), .B(n16313), .Z(n14995) );
  XOR U14939 ( .A(n14998), .B(n14997), .Z(n14996) );
  AND U14940 ( .A(n16314), .B(n16315), .Z(n14997) );
  XOR U14941 ( .A(n15000), .B(n14999), .Z(n14998) );
  AND U14942 ( .A(n16316), .B(n16317), .Z(n14999) );
  XOR U14943 ( .A(n15002), .B(n15001), .Z(n15000) );
  AND U14944 ( .A(n16318), .B(n16319), .Z(n15001) );
  XOR U14945 ( .A(n15004), .B(n15003), .Z(n15002) );
  AND U14946 ( .A(n16320), .B(n16321), .Z(n15003) );
  XOR U14947 ( .A(n15006), .B(n15005), .Z(n15004) );
  AND U14948 ( .A(n16322), .B(n16323), .Z(n15005) );
  XOR U14949 ( .A(n15008), .B(n15007), .Z(n15006) );
  AND U14950 ( .A(n16324), .B(n16325), .Z(n15007) );
  XOR U14951 ( .A(n15010), .B(n15009), .Z(n15008) );
  AND U14952 ( .A(n16326), .B(n16327), .Z(n15009) );
  XOR U14953 ( .A(n15012), .B(n15011), .Z(n15010) );
  AND U14954 ( .A(n16328), .B(n16329), .Z(n15011) );
  XOR U14955 ( .A(n15014), .B(n15013), .Z(n15012) );
  AND U14956 ( .A(n16330), .B(n16331), .Z(n15013) );
  XOR U14957 ( .A(n15016), .B(n15015), .Z(n15014) );
  AND U14958 ( .A(n16332), .B(n16333), .Z(n15015) );
  XOR U14959 ( .A(n15018), .B(n15017), .Z(n15016) );
  AND U14960 ( .A(n16334), .B(n16335), .Z(n15017) );
  XOR U14961 ( .A(n15020), .B(n15019), .Z(n15018) );
  AND U14962 ( .A(n16336), .B(n16337), .Z(n15019) );
  XOR U14963 ( .A(n15022), .B(n15021), .Z(n15020) );
  AND U14964 ( .A(n16338), .B(n16339), .Z(n15021) );
  XOR U14965 ( .A(n15024), .B(n15023), .Z(n15022) );
  AND U14966 ( .A(n16340), .B(n16341), .Z(n15023) );
  XOR U14967 ( .A(n15026), .B(n15025), .Z(n15024) );
  AND U14968 ( .A(n16342), .B(n16343), .Z(n15025) );
  XOR U14969 ( .A(n15028), .B(n15027), .Z(n15026) );
  AND U14970 ( .A(n16344), .B(n16345), .Z(n15027) );
  XOR U14971 ( .A(n15030), .B(n15029), .Z(n15028) );
  AND U14972 ( .A(n16346), .B(n16347), .Z(n15029) );
  XOR U14973 ( .A(n15032), .B(n15031), .Z(n15030) );
  AND U14974 ( .A(n16348), .B(n16349), .Z(n15031) );
  XOR U14975 ( .A(n15034), .B(n15033), .Z(n15032) );
  AND U14976 ( .A(n16350), .B(n16351), .Z(n15033) );
  XOR U14977 ( .A(n15036), .B(n15035), .Z(n15034) );
  AND U14978 ( .A(n16352), .B(n16353), .Z(n15035) );
  XOR U14979 ( .A(n15038), .B(n15037), .Z(n15036) );
  AND U14980 ( .A(n16354), .B(n16355), .Z(n15037) );
  XOR U14981 ( .A(n15040), .B(n15039), .Z(n15038) );
  AND U14982 ( .A(n16356), .B(n16357), .Z(n15039) );
  XOR U14983 ( .A(n15042), .B(n15041), .Z(n15040) );
  AND U14984 ( .A(n16358), .B(n16359), .Z(n15041) );
  XOR U14985 ( .A(n15044), .B(n15043), .Z(n15042) );
  AND U14986 ( .A(n16360), .B(n16361), .Z(n15043) );
  XOR U14987 ( .A(n15046), .B(n15045), .Z(n15044) );
  AND U14988 ( .A(n16362), .B(n16363), .Z(n15045) );
  XOR U14989 ( .A(n15048), .B(n15047), .Z(n15046) );
  AND U14990 ( .A(n16364), .B(n16365), .Z(n15047) );
  XOR U14991 ( .A(n15050), .B(n15049), .Z(n15048) );
  AND U14992 ( .A(n16366), .B(n16367), .Z(n15049) );
  XOR U14993 ( .A(n15052), .B(n15051), .Z(n15050) );
  AND U14994 ( .A(n16368), .B(n16369), .Z(n15051) );
  XOR U14995 ( .A(n15054), .B(n15053), .Z(n15052) );
  AND U14996 ( .A(n16370), .B(n16371), .Z(n15053) );
  XOR U14997 ( .A(n15056), .B(n15055), .Z(n15054) );
  AND U14998 ( .A(n16372), .B(n16373), .Z(n15055) );
  XOR U14999 ( .A(n15058), .B(n15057), .Z(n15056) );
  AND U15000 ( .A(n16374), .B(n16375), .Z(n15057) );
  XOR U15001 ( .A(n15060), .B(n15059), .Z(n15058) );
  AND U15002 ( .A(n16376), .B(n16377), .Z(n15059) );
  XOR U15003 ( .A(n15062), .B(n15061), .Z(n15060) );
  AND U15004 ( .A(n16378), .B(n16379), .Z(n15061) );
  XOR U15005 ( .A(n15064), .B(n15063), .Z(n15062) );
  AND U15006 ( .A(n16380), .B(n16381), .Z(n15063) );
  XOR U15007 ( .A(n15066), .B(n15065), .Z(n15064) );
  AND U15008 ( .A(n16382), .B(n16383), .Z(n15065) );
  XOR U15009 ( .A(n15068), .B(n15067), .Z(n15066) );
  AND U15010 ( .A(n16384), .B(n16385), .Z(n15067) );
  XOR U15011 ( .A(n15070), .B(n15069), .Z(n15068) );
  AND U15012 ( .A(n16386), .B(n16387), .Z(n15069) );
  XOR U15013 ( .A(n15072), .B(n15071), .Z(n15070) );
  AND U15014 ( .A(n16388), .B(n16389), .Z(n15071) );
  XOR U15015 ( .A(n15074), .B(n15073), .Z(n15072) );
  AND U15016 ( .A(n16390), .B(n16391), .Z(n15073) );
  XOR U15017 ( .A(n15127), .B(n15075), .Z(n15074) );
  AND U15018 ( .A(n16392), .B(n16393), .Z(n15075) );
  XOR U15019 ( .A(n15129), .B(n15128), .Z(n15127) );
  AND U15020 ( .A(n16394), .B(n16395), .Z(n15128) );
  XOR U15021 ( .A(n15110), .B(n15130), .Z(n15129) );
  AND U15022 ( .A(n16396), .B(n16397), .Z(n15130) );
  XOR U15023 ( .A(n15112), .B(n15111), .Z(n15110) );
  AND U15024 ( .A(n16398), .B(n16399), .Z(n15111) );
  XOR U15025 ( .A(n15114), .B(n15113), .Z(n15112) );
  AND U15026 ( .A(n16400), .B(n16401), .Z(n15113) );
  XOR U15027 ( .A(n15118), .B(n15115), .Z(n15114) );
  AND U15028 ( .A(n16402), .B(n16403), .Z(n15115) );
  XOR U15029 ( .A(n15120), .B(n15119), .Z(n15118) );
  AND U15030 ( .A(n16404), .B(n16405), .Z(n15119) );
  XOR U15031 ( .A(n15123), .B(n15121), .Z(n15120) );
  AND U15032 ( .A(n16406), .B(n16407), .Z(n15121) );
  XOR U15033 ( .A(n15125), .B(n15124), .Z(n15123) );
  AND U15034 ( .A(n16408), .B(n16409), .Z(n15124) );
  XOR U15035 ( .A(n15090), .B(n15126), .Z(n15125) );
  AND U15036 ( .A(n16410), .B(n16411), .Z(n15126) );
  XNOR U15037 ( .A(n15097), .B(n15091), .Z(n15090) );
  AND U15038 ( .A(n16412), .B(n16413), .Z(n15091) );
  XOR U15039 ( .A(n15096), .B(n15088), .Z(n15097) );
  AND U15040 ( .A(n16414), .B(n16415), .Z(n15088) );
  XOR U15041 ( .A(n15109), .B(n15087), .Z(n15096) );
  AND U15042 ( .A(n16416), .B(n16417), .Z(n15087) );
  XNOR U15043 ( .A(n16418), .B(n16419), .Z(n15109) );
  XOR U15044 ( .A(n15107), .B(n16420), .Z(n16419) );
  XOR U15045 ( .A(n15105), .B(n15103), .Z(n16420) );
  AND U15046 ( .A(n16421), .B(n16422), .Z(n15103) );
  AND U15047 ( .A(n16423), .B(n16424), .Z(n15105) );
  AND U15048 ( .A(n16425), .B(n16426), .Z(n15107) );
  XNOR U15049 ( .A(n16427), .B(n15106), .Z(n16418) );
  XOR U15050 ( .A(n16428), .B(n16429), .Z(n15106) );
  XOR U15051 ( .A(n16430), .B(n16431), .Z(n16429) );
  AND U15052 ( .A(n16432), .B(n16433), .Z(n16431) );
  XNOR U15053 ( .A(n16434), .B(n16435), .Z(n16428) );
  NOR U15054 ( .A(n16436), .B(n16437), .Z(n16435) );
  AND U15055 ( .A(n16438), .B(n16439), .Z(n16437) );
  IV U15056 ( .A(n16440), .Z(n16436) );
  NOR U15057 ( .A(n16430), .B(n16441), .Z(n16440) );
  AND U15058 ( .A(n16442), .B(n16443), .Z(n16441) );
  NOR U15059 ( .A(n16432), .B(n16442), .Z(n16434) );
  XNOR U15060 ( .A(n15108), .B(n15086), .Z(n16427) );
  AND U15061 ( .A(n16444), .B(n16445), .Z(n15086) );
  AND U15062 ( .A(n16446), .B(n16447), .Z(n15108) );
  XOR U15063 ( .A(n16448), .B(n16449), .Z(n15143) );
  NOR U15064 ( .A(n16450), .B(n16451), .Z(n16449) );
  IV U15065 ( .A(n16448), .Z(n16450) );
  XOR U15066 ( .A(n16452), .B(n16453), .Z(n15146) );
  NOR U15067 ( .A(n16452), .B(n16454), .Z(n16453) );
  XNOR U15068 ( .A(n16455), .B(n16456), .Z(n15149) );
  AND U15069 ( .A(n16455), .B(n16457), .Z(n16456) );
  XNOR U15070 ( .A(n16458), .B(n16459), .Z(n15152) );
  AND U15071 ( .A(n16458), .B(n16460), .Z(n16459) );
  XNOR U15072 ( .A(n16461), .B(n16462), .Z(n15155) );
  AND U15073 ( .A(n16461), .B(n16463), .Z(n16462) );
  XNOR U15074 ( .A(n16464), .B(n16465), .Z(n15158) );
  AND U15075 ( .A(n16464), .B(n16466), .Z(n16465) );
  XNOR U15076 ( .A(n16467), .B(n16468), .Z(n15161) );
  AND U15077 ( .A(n16467), .B(n16469), .Z(n16468) );
  XNOR U15078 ( .A(n16470), .B(n16471), .Z(n15164) );
  AND U15079 ( .A(n16470), .B(n16472), .Z(n16471) );
  XNOR U15080 ( .A(n16473), .B(n16474), .Z(n15167) );
  AND U15081 ( .A(n16473), .B(n16475), .Z(n16474) );
  XNOR U15082 ( .A(n16476), .B(n16477), .Z(n15170) );
  AND U15083 ( .A(n16476), .B(n16478), .Z(n16477) );
  XNOR U15084 ( .A(n16479), .B(n16480), .Z(n15173) );
  AND U15085 ( .A(n16479), .B(n16481), .Z(n16480) );
  XNOR U15086 ( .A(n16482), .B(n16483), .Z(n15176) );
  AND U15087 ( .A(n16482), .B(n16484), .Z(n16483) );
  XNOR U15088 ( .A(n16485), .B(n16486), .Z(n15179) );
  AND U15089 ( .A(n16485), .B(n16487), .Z(n16486) );
  XNOR U15090 ( .A(n16488), .B(n16489), .Z(n15182) );
  AND U15091 ( .A(n16488), .B(n16490), .Z(n16489) );
  XNOR U15092 ( .A(n16491), .B(n16492), .Z(n15185) );
  AND U15093 ( .A(n16491), .B(n16493), .Z(n16492) );
  XNOR U15094 ( .A(n16494), .B(n16495), .Z(n15188) );
  AND U15095 ( .A(n16494), .B(n16496), .Z(n16495) );
  XNOR U15096 ( .A(n16497), .B(n16498), .Z(n15191) );
  AND U15097 ( .A(n16497), .B(n16499), .Z(n16498) );
  XNOR U15098 ( .A(n16500), .B(n16501), .Z(n15194) );
  AND U15099 ( .A(n16500), .B(n16502), .Z(n16501) );
  XNOR U15100 ( .A(n16503), .B(n16504), .Z(n15197) );
  AND U15101 ( .A(n16503), .B(n16505), .Z(n16504) );
  XNOR U15102 ( .A(n16506), .B(n16507), .Z(n15200) );
  AND U15103 ( .A(n16506), .B(n16508), .Z(n16507) );
  XNOR U15104 ( .A(n16509), .B(n16510), .Z(n15203) );
  AND U15105 ( .A(n16509), .B(n16511), .Z(n16510) );
  XNOR U15106 ( .A(n16512), .B(n16513), .Z(n15206) );
  AND U15107 ( .A(n16512), .B(n16514), .Z(n16513) );
  XNOR U15108 ( .A(n16515), .B(n16516), .Z(n15209) );
  AND U15109 ( .A(n16515), .B(n16517), .Z(n16516) );
  XNOR U15110 ( .A(n16518), .B(n16519), .Z(n15212) );
  AND U15111 ( .A(n16518), .B(n16520), .Z(n16519) );
  XNOR U15112 ( .A(n16521), .B(n16522), .Z(n15215) );
  AND U15113 ( .A(n16521), .B(n16523), .Z(n16522) );
  XNOR U15114 ( .A(n16524), .B(n16525), .Z(n15218) );
  AND U15115 ( .A(n16524), .B(n16526), .Z(n16525) );
  XNOR U15116 ( .A(n16527), .B(n16528), .Z(n15221) );
  AND U15117 ( .A(n16527), .B(n16529), .Z(n16528) );
  XNOR U15118 ( .A(n16530), .B(n16531), .Z(n15224) );
  AND U15119 ( .A(n16530), .B(n16532), .Z(n16531) );
  XNOR U15120 ( .A(n16533), .B(n16534), .Z(n15227) );
  AND U15121 ( .A(n16533), .B(n16535), .Z(n16534) );
  XNOR U15122 ( .A(n16536), .B(n16537), .Z(n15230) );
  AND U15123 ( .A(n16536), .B(n16538), .Z(n16537) );
  XNOR U15124 ( .A(n16539), .B(n16540), .Z(n15233) );
  AND U15125 ( .A(n16539), .B(n16541), .Z(n16540) );
  XNOR U15126 ( .A(n16542), .B(n16543), .Z(n15236) );
  AND U15127 ( .A(n16542), .B(n16544), .Z(n16543) );
  XNOR U15128 ( .A(n16545), .B(n16546), .Z(n15239) );
  AND U15129 ( .A(n16545), .B(n16547), .Z(n16546) );
  XNOR U15130 ( .A(n16548), .B(n16549), .Z(n15242) );
  AND U15131 ( .A(n16548), .B(n16550), .Z(n16549) );
  XNOR U15132 ( .A(n16551), .B(n16552), .Z(n15245) );
  AND U15133 ( .A(n16551), .B(n16553), .Z(n16552) );
  XNOR U15134 ( .A(n16554), .B(n16555), .Z(n15248) );
  AND U15135 ( .A(n16554), .B(n16556), .Z(n16555) );
  XNOR U15136 ( .A(n16557), .B(n16558), .Z(n15251) );
  AND U15137 ( .A(n16557), .B(n16559), .Z(n16558) );
  XNOR U15138 ( .A(n16560), .B(n16561), .Z(n15254) );
  AND U15139 ( .A(n16560), .B(n16562), .Z(n16561) );
  XNOR U15140 ( .A(n16563), .B(n16564), .Z(n15257) );
  AND U15141 ( .A(n16563), .B(n16565), .Z(n16564) );
  XNOR U15142 ( .A(n16566), .B(n16567), .Z(n15260) );
  AND U15143 ( .A(n16566), .B(n16568), .Z(n16567) );
  XNOR U15144 ( .A(n16569), .B(n16570), .Z(n15263) );
  AND U15145 ( .A(n16569), .B(n16571), .Z(n16570) );
  XNOR U15146 ( .A(n16572), .B(n16573), .Z(n15266) );
  AND U15147 ( .A(n16572), .B(n16574), .Z(n16573) );
  XNOR U15148 ( .A(n16575), .B(n16576), .Z(n15269) );
  AND U15149 ( .A(n16575), .B(n16577), .Z(n16576) );
  XNOR U15150 ( .A(n16578), .B(n16579), .Z(n15272) );
  AND U15151 ( .A(n16578), .B(n16580), .Z(n16579) );
  XNOR U15152 ( .A(n16581), .B(n16582), .Z(n15275) );
  AND U15153 ( .A(n16581), .B(n16583), .Z(n16582) );
  XNOR U15154 ( .A(n16584), .B(n16585), .Z(n15278) );
  AND U15155 ( .A(n16584), .B(n16586), .Z(n16585) );
  XNOR U15156 ( .A(n16587), .B(n16588), .Z(n15281) );
  AND U15157 ( .A(n16587), .B(n16589), .Z(n16588) );
  XNOR U15158 ( .A(n16590), .B(n16591), .Z(n15284) );
  AND U15159 ( .A(n16590), .B(n16592), .Z(n16591) );
  XNOR U15160 ( .A(n16593), .B(n16594), .Z(n15287) );
  AND U15161 ( .A(n16593), .B(n16595), .Z(n16594) );
  XNOR U15162 ( .A(n16596), .B(n16597), .Z(n15290) );
  AND U15163 ( .A(n16596), .B(n16598), .Z(n16597) );
  XNOR U15164 ( .A(n16599), .B(n16600), .Z(n15293) );
  AND U15165 ( .A(n16599), .B(n16601), .Z(n16600) );
  XNOR U15166 ( .A(n16602), .B(n16603), .Z(n15296) );
  AND U15167 ( .A(n16602), .B(n16604), .Z(n16603) );
  XNOR U15168 ( .A(n16605), .B(n16606), .Z(n15299) );
  AND U15169 ( .A(n16605), .B(n16607), .Z(n16606) );
  XNOR U15170 ( .A(n16608), .B(n16609), .Z(n15302) );
  AND U15171 ( .A(n16608), .B(n16610), .Z(n16609) );
  XNOR U15172 ( .A(n16611), .B(n16612), .Z(n15305) );
  AND U15173 ( .A(n16611), .B(n16613), .Z(n16612) );
  XNOR U15174 ( .A(n16614), .B(n16615), .Z(n15308) );
  AND U15175 ( .A(n16614), .B(n16616), .Z(n16615) );
  XNOR U15176 ( .A(n16617), .B(n16618), .Z(n15311) );
  AND U15177 ( .A(n16617), .B(n16619), .Z(n16618) );
  XNOR U15178 ( .A(n16620), .B(n16621), .Z(n15314) );
  AND U15179 ( .A(n16620), .B(n16622), .Z(n16621) );
  XNOR U15180 ( .A(n16623), .B(n16624), .Z(n15317) );
  AND U15181 ( .A(n16623), .B(n16625), .Z(n16624) );
  XNOR U15182 ( .A(n16626), .B(n16627), .Z(n15320) );
  AND U15183 ( .A(n16626), .B(n16628), .Z(n16627) );
  XNOR U15184 ( .A(n16629), .B(n16630), .Z(n15323) );
  AND U15185 ( .A(n16629), .B(n16631), .Z(n16630) );
  XNOR U15186 ( .A(n16632), .B(n16633), .Z(n15326) );
  AND U15187 ( .A(n16632), .B(n16634), .Z(n16633) );
  XNOR U15188 ( .A(n16635), .B(n16636), .Z(n15329) );
  AND U15189 ( .A(n16635), .B(n16637), .Z(n16636) );
  XNOR U15190 ( .A(n16638), .B(n16639), .Z(n15332) );
  AND U15191 ( .A(n16638), .B(n16640), .Z(n16639) );
  XNOR U15192 ( .A(n16641), .B(n16642), .Z(n15335) );
  AND U15193 ( .A(n16641), .B(n16643), .Z(n16642) );
  XNOR U15194 ( .A(n16644), .B(n16645), .Z(n15338) );
  AND U15195 ( .A(n16644), .B(n16646), .Z(n16645) );
  XNOR U15196 ( .A(n16647), .B(n16648), .Z(n15341) );
  AND U15197 ( .A(n16647), .B(n16649), .Z(n16648) );
  XNOR U15198 ( .A(n16650), .B(n16651), .Z(n15344) );
  AND U15199 ( .A(n16650), .B(n16652), .Z(n16651) );
  XNOR U15200 ( .A(n16653), .B(n16654), .Z(n15347) );
  AND U15201 ( .A(n16653), .B(n16655), .Z(n16654) );
  XNOR U15202 ( .A(n16656), .B(n16657), .Z(n15350) );
  AND U15203 ( .A(n16656), .B(n16658), .Z(n16657) );
  XNOR U15204 ( .A(n16659), .B(n16660), .Z(n15353) );
  AND U15205 ( .A(n16659), .B(n16661), .Z(n16660) );
  XNOR U15206 ( .A(n16662), .B(n16663), .Z(n15356) );
  AND U15207 ( .A(n16662), .B(n16664), .Z(n16663) );
  XNOR U15208 ( .A(n16665), .B(n16666), .Z(n15359) );
  AND U15209 ( .A(n16665), .B(n16667), .Z(n16666) );
  XNOR U15210 ( .A(n16668), .B(n16669), .Z(n15362) );
  AND U15211 ( .A(n16668), .B(n16670), .Z(n16669) );
  XNOR U15212 ( .A(n16671), .B(n16672), .Z(n15365) );
  AND U15213 ( .A(n16671), .B(n16673), .Z(n16672) );
  XNOR U15214 ( .A(n16674), .B(n16675), .Z(n15368) );
  AND U15215 ( .A(n16674), .B(n16676), .Z(n16675) );
  XNOR U15216 ( .A(n16677), .B(n16678), .Z(n15371) );
  AND U15217 ( .A(n16677), .B(n16679), .Z(n16678) );
  XNOR U15218 ( .A(n16680), .B(n16681), .Z(n15374) );
  AND U15219 ( .A(n16680), .B(n16682), .Z(n16681) );
  XNOR U15220 ( .A(n16683), .B(n16684), .Z(n15377) );
  AND U15221 ( .A(n16683), .B(n16685), .Z(n16684) );
  XNOR U15222 ( .A(n16686), .B(n16687), .Z(n15380) );
  AND U15223 ( .A(n16686), .B(n16688), .Z(n16687) );
  XNOR U15224 ( .A(n16689), .B(n16690), .Z(n15383) );
  AND U15225 ( .A(n16689), .B(n16691), .Z(n16690) );
  XNOR U15226 ( .A(n16692), .B(n16693), .Z(n15386) );
  AND U15227 ( .A(n16692), .B(n16694), .Z(n16693) );
  XNOR U15228 ( .A(n16695), .B(n16696), .Z(n15389) );
  AND U15229 ( .A(n16695), .B(n16697), .Z(n16696) );
  XNOR U15230 ( .A(n16698), .B(n16699), .Z(n15392) );
  AND U15231 ( .A(n16698), .B(n16700), .Z(n16699) );
  XNOR U15232 ( .A(n16701), .B(n16702), .Z(n15395) );
  AND U15233 ( .A(n16701), .B(n16703), .Z(n16702) );
  XNOR U15234 ( .A(n16704), .B(n16705), .Z(n15398) );
  AND U15235 ( .A(n16704), .B(n16706), .Z(n16705) );
  XNOR U15236 ( .A(n16707), .B(n16708), .Z(n15401) );
  AND U15237 ( .A(n16707), .B(n16709), .Z(n16708) );
  XNOR U15238 ( .A(n16710), .B(n16711), .Z(n15404) );
  AND U15239 ( .A(n16710), .B(n16712), .Z(n16711) );
  XNOR U15240 ( .A(n16713), .B(n16714), .Z(n15407) );
  AND U15241 ( .A(n16713), .B(n16715), .Z(n16714) );
  XNOR U15242 ( .A(n16716), .B(n16717), .Z(n15410) );
  AND U15243 ( .A(n16716), .B(n16718), .Z(n16717) );
  XNOR U15244 ( .A(n16719), .B(n16720), .Z(n15413) );
  AND U15245 ( .A(n16719), .B(n16721), .Z(n16720) );
  XNOR U15246 ( .A(n16722), .B(n16723), .Z(n15416) );
  AND U15247 ( .A(n16722), .B(n16724), .Z(n16723) );
  XNOR U15248 ( .A(n16725), .B(n16726), .Z(n15419) );
  AND U15249 ( .A(n16725), .B(n16727), .Z(n16726) );
  XNOR U15250 ( .A(n16728), .B(n16729), .Z(n15422) );
  AND U15251 ( .A(n16728), .B(n16730), .Z(n16729) );
  XNOR U15252 ( .A(n16731), .B(n16732), .Z(n15425) );
  AND U15253 ( .A(n16731), .B(n16733), .Z(n16732) );
  XNOR U15254 ( .A(n16734), .B(n16735), .Z(n15428) );
  AND U15255 ( .A(n16734), .B(n16736), .Z(n16735) );
  XNOR U15256 ( .A(n16737), .B(n16738), .Z(n15431) );
  AND U15257 ( .A(n16737), .B(n16739), .Z(n16738) );
  XNOR U15258 ( .A(n16740), .B(n16741), .Z(n15434) );
  AND U15259 ( .A(n16740), .B(n16742), .Z(n16741) );
  XNOR U15260 ( .A(n16743), .B(n16744), .Z(n15437) );
  AND U15261 ( .A(n16743), .B(n16745), .Z(n16744) );
  XNOR U15262 ( .A(n16746), .B(n16747), .Z(n15440) );
  AND U15263 ( .A(n16746), .B(n16748), .Z(n16747) );
  XNOR U15264 ( .A(n16749), .B(n16750), .Z(n15443) );
  AND U15265 ( .A(n16749), .B(n16751), .Z(n16750) );
  XNOR U15266 ( .A(n16752), .B(n16753), .Z(n15446) );
  AND U15267 ( .A(n16752), .B(n16754), .Z(n16753) );
  XNOR U15268 ( .A(n16755), .B(n16756), .Z(n15449) );
  AND U15269 ( .A(n16755), .B(n16757), .Z(n16756) );
  XNOR U15270 ( .A(n16758), .B(n16759), .Z(n15452) );
  AND U15271 ( .A(n16758), .B(n16760), .Z(n16759) );
  XNOR U15272 ( .A(n16761), .B(n16762), .Z(n15455) );
  AND U15273 ( .A(n16761), .B(n16763), .Z(n16762) );
  XNOR U15274 ( .A(n16764), .B(n16765), .Z(n15458) );
  AND U15275 ( .A(n16764), .B(n16766), .Z(n16765) );
  XNOR U15276 ( .A(n16767), .B(n16768), .Z(n15461) );
  AND U15277 ( .A(n16767), .B(n16769), .Z(n16768) );
  XNOR U15278 ( .A(n16770), .B(n16771), .Z(n15464) );
  AND U15279 ( .A(n16770), .B(n16772), .Z(n16771) );
  XNOR U15280 ( .A(n16773), .B(n16774), .Z(n15467) );
  AND U15281 ( .A(n16773), .B(n16775), .Z(n16774) );
  XNOR U15282 ( .A(n16776), .B(n16777), .Z(n15470) );
  AND U15283 ( .A(n16776), .B(n16778), .Z(n16777) );
  XNOR U15284 ( .A(n16779), .B(n16780), .Z(n15473) );
  AND U15285 ( .A(n16779), .B(n16781), .Z(n16780) );
  XNOR U15286 ( .A(n16782), .B(n16783), .Z(n15476) );
  AND U15287 ( .A(n16782), .B(n16784), .Z(n16783) );
  XNOR U15288 ( .A(n16785), .B(n16786), .Z(n15479) );
  AND U15289 ( .A(n16785), .B(n16787), .Z(n16786) );
  XNOR U15290 ( .A(n16788), .B(n16789), .Z(n15482) );
  AND U15291 ( .A(n16788), .B(n16790), .Z(n16789) );
  XNOR U15292 ( .A(n16791), .B(n16792), .Z(n15485) );
  AND U15293 ( .A(n16791), .B(n16793), .Z(n16792) );
  XNOR U15294 ( .A(n16794), .B(n16795), .Z(n15488) );
  AND U15295 ( .A(n16794), .B(n16796), .Z(n16795) );
  XNOR U15296 ( .A(n16797), .B(n16798), .Z(n15491) );
  AND U15297 ( .A(n16797), .B(n16799), .Z(n16798) );
  XNOR U15298 ( .A(n16800), .B(n16801), .Z(n15494) );
  AND U15299 ( .A(n16800), .B(n16802), .Z(n16801) );
  XNOR U15300 ( .A(n16803), .B(n16804), .Z(n15497) );
  AND U15301 ( .A(n16803), .B(n16805), .Z(n16804) );
  XNOR U15302 ( .A(n16806), .B(n16807), .Z(n15500) );
  AND U15303 ( .A(n16806), .B(n16808), .Z(n16807) );
  XNOR U15304 ( .A(n16809), .B(n16810), .Z(n15503) );
  AND U15305 ( .A(n16809), .B(n16811), .Z(n16810) );
  XNOR U15306 ( .A(n16812), .B(n16813), .Z(n15506) );
  AND U15307 ( .A(n16812), .B(n16814), .Z(n16813) );
  XNOR U15308 ( .A(n16815), .B(n16816), .Z(n15509) );
  AND U15309 ( .A(n16815), .B(n16817), .Z(n16816) );
  XNOR U15310 ( .A(n16818), .B(n16819), .Z(n15512) );
  AND U15311 ( .A(n16818), .B(n16820), .Z(n16819) );
  XNOR U15312 ( .A(n16821), .B(n16822), .Z(n15515) );
  AND U15313 ( .A(n16821), .B(n16823), .Z(n16822) );
  XNOR U15314 ( .A(n16824), .B(n16825), .Z(n15518) );
  AND U15315 ( .A(n16824), .B(n16826), .Z(n16825) );
  XNOR U15316 ( .A(n16827), .B(n16828), .Z(n15521) );
  AND U15317 ( .A(n16827), .B(n16829), .Z(n16828) );
  XNOR U15318 ( .A(n16830), .B(n16831), .Z(n15524) );
  AND U15319 ( .A(n16830), .B(n16832), .Z(n16831) );
  XNOR U15320 ( .A(n16833), .B(n16834), .Z(n15527) );
  AND U15321 ( .A(n16833), .B(n16835), .Z(n16834) );
  XNOR U15322 ( .A(n16836), .B(n16837), .Z(n15530) );
  AND U15323 ( .A(n16836), .B(n16838), .Z(n16837) );
  XOR U15324 ( .A(n16839), .B(n16840), .Z(n15533) );
  AND U15325 ( .A(n16839), .B(n123), .Z(n16840) );
  XOR U15326 ( .A(n105), .B(n16188), .Z(n16190) );
  XOR U15327 ( .A(n16185), .B(n16184), .Z(n105) );
  XNOR U15328 ( .A(n16182), .B(n16181), .Z(n16184) );
  XNOR U15329 ( .A(n16179), .B(n16178), .Z(n16181) );
  XNOR U15330 ( .A(n16176), .B(n16175), .Z(n16178) );
  XNOR U15331 ( .A(n16173), .B(n16172), .Z(n16175) );
  XNOR U15332 ( .A(n16170), .B(n16169), .Z(n16172) );
  XNOR U15333 ( .A(n16167), .B(n16166), .Z(n16169) );
  XNOR U15334 ( .A(n16164), .B(n16163), .Z(n16166) );
  XNOR U15335 ( .A(n16161), .B(n16160), .Z(n16163) );
  XNOR U15336 ( .A(n16158), .B(n16157), .Z(n16160) );
  XNOR U15337 ( .A(n16155), .B(n16154), .Z(n16157) );
  XNOR U15338 ( .A(n16152), .B(n16151), .Z(n16154) );
  XNOR U15339 ( .A(n16149), .B(n16148), .Z(n16151) );
  XNOR U15340 ( .A(n16146), .B(n16145), .Z(n16148) );
  XNOR U15341 ( .A(n16143), .B(n16142), .Z(n16145) );
  XNOR U15342 ( .A(n16140), .B(n16139), .Z(n16142) );
  XNOR U15343 ( .A(n16137), .B(n16136), .Z(n16139) );
  XNOR U15344 ( .A(n16134), .B(n16133), .Z(n16136) );
  XNOR U15345 ( .A(n16131), .B(n16130), .Z(n16133) );
  XNOR U15346 ( .A(n16128), .B(n16127), .Z(n16130) );
  XNOR U15347 ( .A(n16125), .B(n16124), .Z(n16127) );
  XNOR U15348 ( .A(n16122), .B(n16121), .Z(n16124) );
  XNOR U15349 ( .A(n16119), .B(n16118), .Z(n16121) );
  XNOR U15350 ( .A(n16116), .B(n16115), .Z(n16118) );
  XNOR U15351 ( .A(n16113), .B(n16112), .Z(n16115) );
  XNOR U15352 ( .A(n16110), .B(n16109), .Z(n16112) );
  XNOR U15353 ( .A(n16107), .B(n16106), .Z(n16109) );
  XNOR U15354 ( .A(n16104), .B(n16103), .Z(n16106) );
  XNOR U15355 ( .A(n16101), .B(n16100), .Z(n16103) );
  XNOR U15356 ( .A(n16098), .B(n16097), .Z(n16100) );
  XNOR U15357 ( .A(n16095), .B(n16094), .Z(n16097) );
  XNOR U15358 ( .A(n16092), .B(n16091), .Z(n16094) );
  XNOR U15359 ( .A(n16089), .B(n16088), .Z(n16091) );
  XNOR U15360 ( .A(n16086), .B(n16085), .Z(n16088) );
  XNOR U15361 ( .A(n16083), .B(n16082), .Z(n16085) );
  XNOR U15362 ( .A(n16080), .B(n16079), .Z(n16082) );
  XNOR U15363 ( .A(n16077), .B(n16076), .Z(n16079) );
  XNOR U15364 ( .A(n16074), .B(n16073), .Z(n16076) );
  XNOR U15365 ( .A(n16071), .B(n16070), .Z(n16073) );
  XNOR U15366 ( .A(n16068), .B(n16067), .Z(n16070) );
  XNOR U15367 ( .A(n16065), .B(n16064), .Z(n16067) );
  XNOR U15368 ( .A(n16062), .B(n16061), .Z(n16064) );
  XNOR U15369 ( .A(n16059), .B(n16058), .Z(n16061) );
  XNOR U15370 ( .A(n16056), .B(n16055), .Z(n16058) );
  XNOR U15371 ( .A(n16053), .B(n16052), .Z(n16055) );
  XNOR U15372 ( .A(n16050), .B(n16049), .Z(n16052) );
  XNOR U15373 ( .A(n16047), .B(n16046), .Z(n16049) );
  XNOR U15374 ( .A(n16044), .B(n16043), .Z(n16046) );
  XNOR U15375 ( .A(n16041), .B(n16040), .Z(n16043) );
  XNOR U15376 ( .A(n16038), .B(n16037), .Z(n16040) );
  XNOR U15377 ( .A(n16035), .B(n16034), .Z(n16037) );
  XNOR U15378 ( .A(n16032), .B(n16031), .Z(n16034) );
  XNOR U15379 ( .A(n16029), .B(n16028), .Z(n16031) );
  XNOR U15380 ( .A(n16026), .B(n16025), .Z(n16028) );
  XNOR U15381 ( .A(n16023), .B(n16022), .Z(n16025) );
  XNOR U15382 ( .A(n16020), .B(n16019), .Z(n16022) );
  XNOR U15383 ( .A(n16017), .B(n16016), .Z(n16019) );
  XNOR U15384 ( .A(n16014), .B(n16013), .Z(n16016) );
  XNOR U15385 ( .A(n16011), .B(n16010), .Z(n16013) );
  XNOR U15386 ( .A(n16008), .B(n16007), .Z(n16010) );
  XNOR U15387 ( .A(n16005), .B(n16004), .Z(n16007) );
  XNOR U15388 ( .A(n16002), .B(n16001), .Z(n16004) );
  XNOR U15389 ( .A(n15999), .B(n15998), .Z(n16001) );
  XNOR U15390 ( .A(n15996), .B(n15995), .Z(n15998) );
  XNOR U15391 ( .A(n15993), .B(n15992), .Z(n15995) );
  XNOR U15392 ( .A(n15990), .B(n15989), .Z(n15992) );
  XNOR U15393 ( .A(n15987), .B(n15986), .Z(n15989) );
  XNOR U15394 ( .A(n15984), .B(n15983), .Z(n15986) );
  XNOR U15395 ( .A(n15981), .B(n15980), .Z(n15983) );
  XNOR U15396 ( .A(n15978), .B(n15977), .Z(n15980) );
  XNOR U15397 ( .A(n15975), .B(n15974), .Z(n15977) );
  XNOR U15398 ( .A(n15972), .B(n15971), .Z(n15974) );
  XNOR U15399 ( .A(n15969), .B(n15968), .Z(n15971) );
  XNOR U15400 ( .A(n15966), .B(n15965), .Z(n15968) );
  XNOR U15401 ( .A(n15963), .B(n15962), .Z(n15965) );
  XNOR U15402 ( .A(n15960), .B(n15959), .Z(n15962) );
  XNOR U15403 ( .A(n15957), .B(n15956), .Z(n15959) );
  XNOR U15404 ( .A(n15954), .B(n15953), .Z(n15956) );
  XNOR U15405 ( .A(n15951), .B(n15950), .Z(n15953) );
  XNOR U15406 ( .A(n15948), .B(n15947), .Z(n15950) );
  XNOR U15407 ( .A(n15945), .B(n15944), .Z(n15947) );
  XNOR U15408 ( .A(n15942), .B(n15941), .Z(n15944) );
  XNOR U15409 ( .A(n15939), .B(n15938), .Z(n15941) );
  XNOR U15410 ( .A(n15936), .B(n15935), .Z(n15938) );
  XNOR U15411 ( .A(n15933), .B(n15932), .Z(n15935) );
  XNOR U15412 ( .A(n15930), .B(n15929), .Z(n15932) );
  XNOR U15413 ( .A(n15927), .B(n15926), .Z(n15929) );
  XNOR U15414 ( .A(n15924), .B(n15923), .Z(n15926) );
  XNOR U15415 ( .A(n15921), .B(n15920), .Z(n15923) );
  XNOR U15416 ( .A(n15918), .B(n15917), .Z(n15920) );
  XNOR U15417 ( .A(n15915), .B(n15914), .Z(n15917) );
  XNOR U15418 ( .A(n15912), .B(n15911), .Z(n15914) );
  XNOR U15419 ( .A(n15909), .B(n15908), .Z(n15911) );
  XNOR U15420 ( .A(n15906), .B(n15905), .Z(n15908) );
  XNOR U15421 ( .A(n15903), .B(n15902), .Z(n15905) );
  XNOR U15422 ( .A(n15900), .B(n15899), .Z(n15902) );
  XNOR U15423 ( .A(n15897), .B(n15896), .Z(n15899) );
  XNOR U15424 ( .A(n15894), .B(n15893), .Z(n15896) );
  XNOR U15425 ( .A(n15891), .B(n15890), .Z(n15893) );
  XNOR U15426 ( .A(n15888), .B(n15887), .Z(n15890) );
  XNOR U15427 ( .A(n15885), .B(n15884), .Z(n15887) );
  XNOR U15428 ( .A(n15882), .B(n15881), .Z(n15884) );
  XNOR U15429 ( .A(n15879), .B(n15878), .Z(n15881) );
  XNOR U15430 ( .A(n15876), .B(n15875), .Z(n15878) );
  XNOR U15431 ( .A(n15873), .B(n15872), .Z(n15875) );
  XNOR U15432 ( .A(n15870), .B(n15869), .Z(n15872) );
  XNOR U15433 ( .A(n15867), .B(n15866), .Z(n15869) );
  XNOR U15434 ( .A(n15864), .B(n15863), .Z(n15866) );
  XNOR U15435 ( .A(n15861), .B(n15860), .Z(n15863) );
  XNOR U15436 ( .A(n15858), .B(n15857), .Z(n15860) );
  XNOR U15437 ( .A(n15855), .B(n15854), .Z(n15857) );
  XNOR U15438 ( .A(n15852), .B(n15851), .Z(n15854) );
  XNOR U15439 ( .A(n15849), .B(n15848), .Z(n15851) );
  XNOR U15440 ( .A(n15846), .B(n15845), .Z(n15848) );
  XNOR U15441 ( .A(n15843), .B(n15842), .Z(n15845) );
  XNOR U15442 ( .A(n15840), .B(n15839), .Z(n15842) );
  XNOR U15443 ( .A(n15837), .B(n15836), .Z(n15839) );
  XNOR U15444 ( .A(n15834), .B(n15833), .Z(n15836) );
  XNOR U15445 ( .A(n15831), .B(n15830), .Z(n15833) );
  XNOR U15446 ( .A(n15828), .B(n15827), .Z(n15830) );
  XNOR U15447 ( .A(n15825), .B(n15824), .Z(n15827) );
  XNOR U15448 ( .A(n15822), .B(n15821), .Z(n15824) );
  XNOR U15449 ( .A(n15819), .B(n15818), .Z(n15821) );
  XNOR U15450 ( .A(n15816), .B(n15815), .Z(n15818) );
  XNOR U15451 ( .A(n15813), .B(n15812), .Z(n15815) );
  XNOR U15452 ( .A(n15810), .B(n15809), .Z(n15812) );
  XNOR U15453 ( .A(n15807), .B(n15806), .Z(n15809) );
  XNOR U15454 ( .A(n15804), .B(n15803), .Z(n15806) );
  XNOR U15455 ( .A(n15801), .B(n15800), .Z(n15803) );
  XOR U15456 ( .A(n15798), .B(n15797), .Z(n15800) );
  XOR U15457 ( .A(n15795), .B(n15794), .Z(n15797) );
  XOR U15458 ( .A(n15791), .B(n15792), .Z(n15794) );
  AND U15459 ( .A(n16841), .B(n16842), .Z(n15792) );
  XOR U15460 ( .A(n15788), .B(n15789), .Z(n15791) );
  AND U15461 ( .A(n16843), .B(n16844), .Z(n15789) );
  XOR U15462 ( .A(n15785), .B(n15786), .Z(n15788) );
  AND U15463 ( .A(n16845), .B(n16846), .Z(n15786) );
  XNOR U15464 ( .A(n15535), .B(n15783), .Z(n15785) );
  AND U15465 ( .A(n16847), .B(n16848), .Z(n15783) );
  XOR U15466 ( .A(n15537), .B(n15536), .Z(n15535) );
  AND U15467 ( .A(n16849), .B(n16850), .Z(n15536) );
  XOR U15468 ( .A(n15539), .B(n15538), .Z(n15537) );
  AND U15469 ( .A(n16851), .B(n16852), .Z(n15538) );
  XOR U15470 ( .A(n15541), .B(n15540), .Z(n15539) );
  AND U15471 ( .A(n16853), .B(n16854), .Z(n15540) );
  XOR U15472 ( .A(n15543), .B(n15542), .Z(n15541) );
  AND U15473 ( .A(n16855), .B(n16856), .Z(n15542) );
  XOR U15474 ( .A(n15545), .B(n15544), .Z(n15543) );
  AND U15475 ( .A(n16857), .B(n16858), .Z(n15544) );
  XOR U15476 ( .A(n15547), .B(n15546), .Z(n15545) );
  AND U15477 ( .A(n16859), .B(n16860), .Z(n15546) );
  XOR U15478 ( .A(n15549), .B(n15548), .Z(n15547) );
  AND U15479 ( .A(n16861), .B(n16862), .Z(n15548) );
  XOR U15480 ( .A(n15551), .B(n15550), .Z(n15549) );
  AND U15481 ( .A(n16863), .B(n16864), .Z(n15550) );
  XOR U15482 ( .A(n15553), .B(n15552), .Z(n15551) );
  AND U15483 ( .A(n16865), .B(n16866), .Z(n15552) );
  XOR U15484 ( .A(n15555), .B(n15554), .Z(n15553) );
  AND U15485 ( .A(n16867), .B(n16868), .Z(n15554) );
  XOR U15486 ( .A(n15557), .B(n15556), .Z(n15555) );
  AND U15487 ( .A(n16869), .B(n16870), .Z(n15556) );
  XOR U15488 ( .A(n15559), .B(n15558), .Z(n15557) );
  AND U15489 ( .A(n16871), .B(n16872), .Z(n15558) );
  XOR U15490 ( .A(n15561), .B(n15560), .Z(n15559) );
  AND U15491 ( .A(n16873), .B(n16874), .Z(n15560) );
  XOR U15492 ( .A(n15563), .B(n15562), .Z(n15561) );
  AND U15493 ( .A(n16875), .B(n16876), .Z(n15562) );
  XOR U15494 ( .A(n15565), .B(n15564), .Z(n15563) );
  AND U15495 ( .A(n16877), .B(n16878), .Z(n15564) );
  XOR U15496 ( .A(n15567), .B(n15566), .Z(n15565) );
  AND U15497 ( .A(n16879), .B(n16880), .Z(n15566) );
  XOR U15498 ( .A(n15569), .B(n15568), .Z(n15567) );
  AND U15499 ( .A(n16881), .B(n16882), .Z(n15568) );
  XOR U15500 ( .A(n15571), .B(n15570), .Z(n15569) );
  AND U15501 ( .A(n16883), .B(n16884), .Z(n15570) );
  XOR U15502 ( .A(n15573), .B(n15572), .Z(n15571) );
  AND U15503 ( .A(n16885), .B(n16886), .Z(n15572) );
  XOR U15504 ( .A(n15575), .B(n15574), .Z(n15573) );
  AND U15505 ( .A(n16887), .B(n16888), .Z(n15574) );
  XOR U15506 ( .A(n15577), .B(n15576), .Z(n15575) );
  AND U15507 ( .A(n16889), .B(n16890), .Z(n15576) );
  XOR U15508 ( .A(n15579), .B(n15578), .Z(n15577) );
  AND U15509 ( .A(n16891), .B(n16892), .Z(n15578) );
  XOR U15510 ( .A(n15581), .B(n15580), .Z(n15579) );
  AND U15511 ( .A(n16893), .B(n16894), .Z(n15580) );
  XOR U15512 ( .A(n15583), .B(n15582), .Z(n15581) );
  AND U15513 ( .A(n16895), .B(n16896), .Z(n15582) );
  XOR U15514 ( .A(n15585), .B(n15584), .Z(n15583) );
  AND U15515 ( .A(n16897), .B(n16898), .Z(n15584) );
  XOR U15516 ( .A(n15587), .B(n15586), .Z(n15585) );
  AND U15517 ( .A(n16899), .B(n16900), .Z(n15586) );
  XOR U15518 ( .A(n15589), .B(n15588), .Z(n15587) );
  AND U15519 ( .A(n16901), .B(n16902), .Z(n15588) );
  XOR U15520 ( .A(n15591), .B(n15590), .Z(n15589) );
  AND U15521 ( .A(n16903), .B(n16904), .Z(n15590) );
  XOR U15522 ( .A(n15593), .B(n15592), .Z(n15591) );
  AND U15523 ( .A(n16905), .B(n16906), .Z(n15592) );
  XOR U15524 ( .A(n15595), .B(n15594), .Z(n15593) );
  AND U15525 ( .A(n16907), .B(n16908), .Z(n15594) );
  XOR U15526 ( .A(n15597), .B(n15596), .Z(n15595) );
  AND U15527 ( .A(n16909), .B(n16910), .Z(n15596) );
  XOR U15528 ( .A(n15599), .B(n15598), .Z(n15597) );
  AND U15529 ( .A(n16911), .B(n16912), .Z(n15598) );
  XOR U15530 ( .A(n15601), .B(n15600), .Z(n15599) );
  AND U15531 ( .A(n16913), .B(n16914), .Z(n15600) );
  XOR U15532 ( .A(n15603), .B(n15602), .Z(n15601) );
  AND U15533 ( .A(n16915), .B(n16916), .Z(n15602) );
  XOR U15534 ( .A(n15605), .B(n15604), .Z(n15603) );
  AND U15535 ( .A(n16917), .B(n16918), .Z(n15604) );
  XOR U15536 ( .A(n15607), .B(n15606), .Z(n15605) );
  AND U15537 ( .A(n16919), .B(n16920), .Z(n15606) );
  XOR U15538 ( .A(n15609), .B(n15608), .Z(n15607) );
  AND U15539 ( .A(n16921), .B(n16922), .Z(n15608) );
  XOR U15540 ( .A(n15611), .B(n15610), .Z(n15609) );
  AND U15541 ( .A(n16923), .B(n16924), .Z(n15610) );
  XOR U15542 ( .A(n15613), .B(n15612), .Z(n15611) );
  AND U15543 ( .A(n16925), .B(n16926), .Z(n15612) );
  XOR U15544 ( .A(n15615), .B(n15614), .Z(n15613) );
  AND U15545 ( .A(n16927), .B(n16928), .Z(n15614) );
  XOR U15546 ( .A(n15617), .B(n15616), .Z(n15615) );
  AND U15547 ( .A(n16929), .B(n16930), .Z(n15616) );
  XOR U15548 ( .A(n15619), .B(n15618), .Z(n15617) );
  AND U15549 ( .A(n16931), .B(n16932), .Z(n15618) );
  XOR U15550 ( .A(n15621), .B(n15620), .Z(n15619) );
  AND U15551 ( .A(n16933), .B(n16934), .Z(n15620) );
  XOR U15552 ( .A(n15623), .B(n15622), .Z(n15621) );
  AND U15553 ( .A(n16935), .B(n16936), .Z(n15622) );
  XOR U15554 ( .A(n15625), .B(n15624), .Z(n15623) );
  AND U15555 ( .A(n16937), .B(n16938), .Z(n15624) );
  XOR U15556 ( .A(n15627), .B(n15626), .Z(n15625) );
  AND U15557 ( .A(n16939), .B(n16940), .Z(n15626) );
  XOR U15558 ( .A(n15629), .B(n15628), .Z(n15627) );
  AND U15559 ( .A(n16941), .B(n16942), .Z(n15628) );
  XOR U15560 ( .A(n15631), .B(n15630), .Z(n15629) );
  AND U15561 ( .A(n16943), .B(n16944), .Z(n15630) );
  XOR U15562 ( .A(n15633), .B(n15632), .Z(n15631) );
  AND U15563 ( .A(n16945), .B(n16946), .Z(n15632) );
  XOR U15564 ( .A(n15635), .B(n15634), .Z(n15633) );
  AND U15565 ( .A(n16947), .B(n16948), .Z(n15634) );
  XOR U15566 ( .A(n15637), .B(n15636), .Z(n15635) );
  AND U15567 ( .A(n16949), .B(n16950), .Z(n15636) );
  XOR U15568 ( .A(n15639), .B(n15638), .Z(n15637) );
  AND U15569 ( .A(n16951), .B(n16952), .Z(n15638) );
  XOR U15570 ( .A(n15641), .B(n15640), .Z(n15639) );
  AND U15571 ( .A(n16953), .B(n16954), .Z(n15640) );
  XOR U15572 ( .A(n15643), .B(n15642), .Z(n15641) );
  AND U15573 ( .A(n16955), .B(n16956), .Z(n15642) );
  XOR U15574 ( .A(n15645), .B(n15644), .Z(n15643) );
  AND U15575 ( .A(n16957), .B(n16958), .Z(n15644) );
  XOR U15576 ( .A(n15647), .B(n15646), .Z(n15645) );
  AND U15577 ( .A(n16959), .B(n16960), .Z(n15646) );
  XOR U15578 ( .A(n15649), .B(n15648), .Z(n15647) );
  AND U15579 ( .A(n16961), .B(n16962), .Z(n15648) );
  XOR U15580 ( .A(n15651), .B(n15650), .Z(n15649) );
  AND U15581 ( .A(n16963), .B(n16964), .Z(n15650) );
  XOR U15582 ( .A(n15653), .B(n15652), .Z(n15651) );
  AND U15583 ( .A(n16965), .B(n16966), .Z(n15652) );
  XOR U15584 ( .A(n15655), .B(n15654), .Z(n15653) );
  AND U15585 ( .A(n16967), .B(n16968), .Z(n15654) );
  XOR U15586 ( .A(n15657), .B(n15656), .Z(n15655) );
  AND U15587 ( .A(n16969), .B(n16970), .Z(n15656) );
  XOR U15588 ( .A(n15659), .B(n15658), .Z(n15657) );
  AND U15589 ( .A(n16971), .B(n16972), .Z(n15658) );
  XOR U15590 ( .A(n15661), .B(n15660), .Z(n15659) );
  AND U15591 ( .A(n16973), .B(n16974), .Z(n15660) );
  XOR U15592 ( .A(n15663), .B(n15662), .Z(n15661) );
  AND U15593 ( .A(n16975), .B(n16976), .Z(n15662) );
  XOR U15594 ( .A(n15665), .B(n15664), .Z(n15663) );
  AND U15595 ( .A(n16977), .B(n16978), .Z(n15664) );
  XOR U15596 ( .A(n15667), .B(n15666), .Z(n15665) );
  AND U15597 ( .A(n16979), .B(n16980), .Z(n15666) );
  XOR U15598 ( .A(n15669), .B(n15668), .Z(n15667) );
  AND U15599 ( .A(n16981), .B(n16982), .Z(n15668) );
  XOR U15600 ( .A(n15671), .B(n15670), .Z(n15669) );
  AND U15601 ( .A(n16983), .B(n16984), .Z(n15670) );
  XOR U15602 ( .A(n15673), .B(n15672), .Z(n15671) );
  AND U15603 ( .A(n16985), .B(n16986), .Z(n15672) );
  XOR U15604 ( .A(n15675), .B(n15674), .Z(n15673) );
  AND U15605 ( .A(n16987), .B(n16988), .Z(n15674) );
  XOR U15606 ( .A(n15677), .B(n15676), .Z(n15675) );
  AND U15607 ( .A(n16989), .B(n16990), .Z(n15676) );
  XOR U15608 ( .A(n15679), .B(n15678), .Z(n15677) );
  AND U15609 ( .A(n16991), .B(n16992), .Z(n15678) );
  XOR U15610 ( .A(n15681), .B(n15680), .Z(n15679) );
  AND U15611 ( .A(n16993), .B(n16994), .Z(n15680) );
  XOR U15612 ( .A(n15683), .B(n15682), .Z(n15681) );
  AND U15613 ( .A(n16995), .B(n16996), .Z(n15682) );
  XOR U15614 ( .A(n15685), .B(n15684), .Z(n15683) );
  AND U15615 ( .A(n16997), .B(n16998), .Z(n15684) );
  XOR U15616 ( .A(n15687), .B(n15686), .Z(n15685) );
  AND U15617 ( .A(n16999), .B(n17000), .Z(n15686) );
  XOR U15618 ( .A(n15689), .B(n15688), .Z(n15687) );
  AND U15619 ( .A(n17001), .B(n17002), .Z(n15688) );
  XOR U15620 ( .A(n15691), .B(n15690), .Z(n15689) );
  AND U15621 ( .A(n17003), .B(n17004), .Z(n15690) );
  XOR U15622 ( .A(n15693), .B(n15692), .Z(n15691) );
  AND U15623 ( .A(n17005), .B(n17006), .Z(n15692) );
  XOR U15624 ( .A(n15695), .B(n15694), .Z(n15693) );
  AND U15625 ( .A(n17007), .B(n17008), .Z(n15694) );
  XOR U15626 ( .A(n15697), .B(n15696), .Z(n15695) );
  AND U15627 ( .A(n17009), .B(n17010), .Z(n15696) );
  XOR U15628 ( .A(n15699), .B(n15698), .Z(n15697) );
  AND U15629 ( .A(n17011), .B(n17012), .Z(n15698) );
  XOR U15630 ( .A(n15701), .B(n15700), .Z(n15699) );
  AND U15631 ( .A(n17013), .B(n17014), .Z(n15700) );
  XOR U15632 ( .A(n15703), .B(n15702), .Z(n15701) );
  AND U15633 ( .A(n17015), .B(n17016), .Z(n15702) );
  XOR U15634 ( .A(n15705), .B(n15704), .Z(n15703) );
  AND U15635 ( .A(n17017), .B(n17018), .Z(n15704) );
  XOR U15636 ( .A(n15707), .B(n15706), .Z(n15705) );
  AND U15637 ( .A(n17019), .B(n17020), .Z(n15706) );
  XOR U15638 ( .A(n15709), .B(n15708), .Z(n15707) );
  AND U15639 ( .A(n17021), .B(n17022), .Z(n15708) );
  XOR U15640 ( .A(n15711), .B(n15710), .Z(n15709) );
  AND U15641 ( .A(n17023), .B(n17024), .Z(n15710) );
  XOR U15642 ( .A(n15713), .B(n15712), .Z(n15711) );
  AND U15643 ( .A(n17025), .B(n17026), .Z(n15712) );
  XOR U15644 ( .A(n15715), .B(n15714), .Z(n15713) );
  AND U15645 ( .A(n17027), .B(n17028), .Z(n15714) );
  XOR U15646 ( .A(n15717), .B(n15716), .Z(n15715) );
  AND U15647 ( .A(n17029), .B(n17030), .Z(n15716) );
  XOR U15648 ( .A(n15719), .B(n15718), .Z(n15717) );
  AND U15649 ( .A(n17031), .B(n17032), .Z(n15718) );
  XOR U15650 ( .A(n15721), .B(n15720), .Z(n15719) );
  AND U15651 ( .A(n17033), .B(n17034), .Z(n15720) );
  XOR U15652 ( .A(n15723), .B(n15722), .Z(n15721) );
  AND U15653 ( .A(n17035), .B(n17036), .Z(n15722) );
  XOR U15654 ( .A(n15725), .B(n15724), .Z(n15723) );
  AND U15655 ( .A(n17037), .B(n17038), .Z(n15724) );
  XOR U15656 ( .A(n15727), .B(n15726), .Z(n15725) );
  AND U15657 ( .A(n17039), .B(n17040), .Z(n15726) );
  XOR U15658 ( .A(n15779), .B(n15728), .Z(n15727) );
  AND U15659 ( .A(n17041), .B(n17042), .Z(n15728) );
  XOR U15660 ( .A(n15781), .B(n15780), .Z(n15779) );
  AND U15661 ( .A(n17043), .B(n17044), .Z(n15780) );
  XOR U15662 ( .A(n15763), .B(n15782), .Z(n15781) );
  AND U15663 ( .A(n17045), .B(n17046), .Z(n15782) );
  XOR U15664 ( .A(n15765), .B(n15764), .Z(n15763) );
  AND U15665 ( .A(n17047), .B(n17048), .Z(n15764) );
  XOR U15666 ( .A(n15767), .B(n15766), .Z(n15765) );
  AND U15667 ( .A(n17049), .B(n17050), .Z(n15766) );
  XOR U15668 ( .A(n15771), .B(n15768), .Z(n15767) );
  AND U15669 ( .A(n17051), .B(n17052), .Z(n15768) );
  XOR U15670 ( .A(n15773), .B(n15772), .Z(n15771) );
  AND U15671 ( .A(n17053), .B(n17054), .Z(n15772) );
  XOR U15672 ( .A(n15775), .B(n15774), .Z(n15773) );
  AND U15673 ( .A(n17055), .B(n17056), .Z(n15774) );
  XOR U15674 ( .A(n15777), .B(n15776), .Z(n15775) );
  AND U15675 ( .A(n17057), .B(n17058), .Z(n15776) );
  XOR U15676 ( .A(n15752), .B(n15778), .Z(n15777) );
  AND U15677 ( .A(n17059), .B(n17060), .Z(n15778) );
  XNOR U15678 ( .A(n15749), .B(n15753), .Z(n15752) );
  AND U15679 ( .A(n17061), .B(n17062), .Z(n15753) );
  XOR U15680 ( .A(n15748), .B(n15740), .Z(n15749) );
  AND U15681 ( .A(n17063), .B(n17064), .Z(n15740) );
  XNOR U15682 ( .A(n15743), .B(n15739), .Z(n15748) );
  AND U15683 ( .A(n17065), .B(n17066), .Z(n15739) );
  XOR U15684 ( .A(n17067), .B(n17068), .Z(n15743) );
  XOR U15685 ( .A(n15761), .B(n17069), .Z(n17068) );
  XOR U15686 ( .A(n15759), .B(n15757), .Z(n17069) );
  AND U15687 ( .A(n17070), .B(n17071), .Z(n15757) );
  AND U15688 ( .A(n17072), .B(n17073), .Z(n15759) );
  AND U15689 ( .A(n17074), .B(n17075), .Z(n15761) );
  XNOR U15690 ( .A(n17076), .B(n15760), .Z(n17067) );
  XOR U15691 ( .A(n17077), .B(n17078), .Z(n15760) );
  XOR U15692 ( .A(n17079), .B(n17080), .Z(n17078) );
  AND U15693 ( .A(n17081), .B(n17082), .Z(n17080) );
  XNOR U15694 ( .A(n17083), .B(n17084), .Z(n17077) );
  NOR U15695 ( .A(n17085), .B(n17086), .Z(n17084) );
  AND U15696 ( .A(n17087), .B(n17088), .Z(n17086) );
  IV U15697 ( .A(n17089), .Z(n17085) );
  NOR U15698 ( .A(n17079), .B(n17090), .Z(n17089) );
  AND U15699 ( .A(n17091), .B(n17092), .Z(n17090) );
  NOR U15700 ( .A(n17081), .B(n17091), .Z(n17083) );
  XNOR U15701 ( .A(n15762), .B(n15744), .Z(n17076) );
  AND U15702 ( .A(n17093), .B(n17094), .Z(n15744) );
  AND U15703 ( .A(n17095), .B(n17096), .Z(n15762) );
  XOR U15704 ( .A(n17097), .B(n17098), .Z(n15795) );
  NOR U15705 ( .A(n17099), .B(n17100), .Z(n17098) );
  IV U15706 ( .A(n17097), .Z(n17099) );
  XOR U15707 ( .A(n17101), .B(n17102), .Z(n15798) );
  NOR U15708 ( .A(n17101), .B(n17103), .Z(n17102) );
  XNOR U15709 ( .A(n17104), .B(n17105), .Z(n15801) );
  AND U15710 ( .A(n17104), .B(n17106), .Z(n17105) );
  XNOR U15711 ( .A(n17107), .B(n17108), .Z(n15804) );
  AND U15712 ( .A(n17107), .B(n17109), .Z(n17108) );
  XNOR U15713 ( .A(n17110), .B(n17111), .Z(n15807) );
  AND U15714 ( .A(n17110), .B(n17112), .Z(n17111) );
  XNOR U15715 ( .A(n17113), .B(n17114), .Z(n15810) );
  AND U15716 ( .A(n17113), .B(n17115), .Z(n17114) );
  XNOR U15717 ( .A(n17116), .B(n17117), .Z(n15813) );
  AND U15718 ( .A(n17116), .B(n17118), .Z(n17117) );
  XNOR U15719 ( .A(n17119), .B(n17120), .Z(n15816) );
  AND U15720 ( .A(n17119), .B(n17121), .Z(n17120) );
  XNOR U15721 ( .A(n17122), .B(n17123), .Z(n15819) );
  AND U15722 ( .A(n17122), .B(n17124), .Z(n17123) );
  XNOR U15723 ( .A(n17125), .B(n17126), .Z(n15822) );
  AND U15724 ( .A(n17125), .B(n17127), .Z(n17126) );
  XNOR U15725 ( .A(n17128), .B(n17129), .Z(n15825) );
  AND U15726 ( .A(n17128), .B(n17130), .Z(n17129) );
  XNOR U15727 ( .A(n17131), .B(n17132), .Z(n15828) );
  AND U15728 ( .A(n17131), .B(n17133), .Z(n17132) );
  XNOR U15729 ( .A(n17134), .B(n17135), .Z(n15831) );
  AND U15730 ( .A(n17134), .B(n17136), .Z(n17135) );
  XNOR U15731 ( .A(n17137), .B(n17138), .Z(n15834) );
  AND U15732 ( .A(n17137), .B(n17139), .Z(n17138) );
  XNOR U15733 ( .A(n17140), .B(n17141), .Z(n15837) );
  AND U15734 ( .A(n17140), .B(n17142), .Z(n17141) );
  XNOR U15735 ( .A(n17143), .B(n17144), .Z(n15840) );
  AND U15736 ( .A(n17143), .B(n17145), .Z(n17144) );
  XNOR U15737 ( .A(n17146), .B(n17147), .Z(n15843) );
  AND U15738 ( .A(n17146), .B(n17148), .Z(n17147) );
  XNOR U15739 ( .A(n17149), .B(n17150), .Z(n15846) );
  AND U15740 ( .A(n17149), .B(n17151), .Z(n17150) );
  XNOR U15741 ( .A(n17152), .B(n17153), .Z(n15849) );
  AND U15742 ( .A(n17152), .B(n17154), .Z(n17153) );
  XNOR U15743 ( .A(n17155), .B(n17156), .Z(n15852) );
  AND U15744 ( .A(n17155), .B(n17157), .Z(n17156) );
  XNOR U15745 ( .A(n17158), .B(n17159), .Z(n15855) );
  AND U15746 ( .A(n17158), .B(n17160), .Z(n17159) );
  XNOR U15747 ( .A(n17161), .B(n17162), .Z(n15858) );
  AND U15748 ( .A(n17161), .B(n17163), .Z(n17162) );
  XNOR U15749 ( .A(n17164), .B(n17165), .Z(n15861) );
  AND U15750 ( .A(n17164), .B(n17166), .Z(n17165) );
  XNOR U15751 ( .A(n17167), .B(n17168), .Z(n15864) );
  AND U15752 ( .A(n17167), .B(n17169), .Z(n17168) );
  XNOR U15753 ( .A(n17170), .B(n17171), .Z(n15867) );
  AND U15754 ( .A(n17170), .B(n17172), .Z(n17171) );
  XNOR U15755 ( .A(n17173), .B(n17174), .Z(n15870) );
  AND U15756 ( .A(n17173), .B(n17175), .Z(n17174) );
  XNOR U15757 ( .A(n17176), .B(n17177), .Z(n15873) );
  AND U15758 ( .A(n17176), .B(n17178), .Z(n17177) );
  XNOR U15759 ( .A(n17179), .B(n17180), .Z(n15876) );
  AND U15760 ( .A(n17179), .B(n17181), .Z(n17180) );
  XNOR U15761 ( .A(n17182), .B(n17183), .Z(n15879) );
  AND U15762 ( .A(n17182), .B(n17184), .Z(n17183) );
  XNOR U15763 ( .A(n17185), .B(n17186), .Z(n15882) );
  AND U15764 ( .A(n17185), .B(n17187), .Z(n17186) );
  XNOR U15765 ( .A(n17188), .B(n17189), .Z(n15885) );
  AND U15766 ( .A(n17188), .B(n17190), .Z(n17189) );
  XNOR U15767 ( .A(n17191), .B(n17192), .Z(n15888) );
  AND U15768 ( .A(n17191), .B(n17193), .Z(n17192) );
  XNOR U15769 ( .A(n17194), .B(n17195), .Z(n15891) );
  AND U15770 ( .A(n17194), .B(n17196), .Z(n17195) );
  XNOR U15771 ( .A(n17197), .B(n17198), .Z(n15894) );
  AND U15772 ( .A(n17197), .B(n17199), .Z(n17198) );
  XNOR U15773 ( .A(n17200), .B(n17201), .Z(n15897) );
  AND U15774 ( .A(n17200), .B(n17202), .Z(n17201) );
  XNOR U15775 ( .A(n17203), .B(n17204), .Z(n15900) );
  AND U15776 ( .A(n17203), .B(n17205), .Z(n17204) );
  XNOR U15777 ( .A(n17206), .B(n17207), .Z(n15903) );
  AND U15778 ( .A(n17206), .B(n17208), .Z(n17207) );
  XNOR U15779 ( .A(n17209), .B(n17210), .Z(n15906) );
  AND U15780 ( .A(n17209), .B(n17211), .Z(n17210) );
  XNOR U15781 ( .A(n17212), .B(n17213), .Z(n15909) );
  AND U15782 ( .A(n17212), .B(n17214), .Z(n17213) );
  XNOR U15783 ( .A(n17215), .B(n17216), .Z(n15912) );
  AND U15784 ( .A(n17215), .B(n17217), .Z(n17216) );
  XNOR U15785 ( .A(n17218), .B(n17219), .Z(n15915) );
  AND U15786 ( .A(n17218), .B(n17220), .Z(n17219) );
  XNOR U15787 ( .A(n17221), .B(n17222), .Z(n15918) );
  AND U15788 ( .A(n17221), .B(n17223), .Z(n17222) );
  XNOR U15789 ( .A(n17224), .B(n17225), .Z(n15921) );
  AND U15790 ( .A(n17224), .B(n17226), .Z(n17225) );
  XNOR U15791 ( .A(n17227), .B(n17228), .Z(n15924) );
  AND U15792 ( .A(n17227), .B(n17229), .Z(n17228) );
  XNOR U15793 ( .A(n17230), .B(n17231), .Z(n15927) );
  AND U15794 ( .A(n17230), .B(n17232), .Z(n17231) );
  XNOR U15795 ( .A(n17233), .B(n17234), .Z(n15930) );
  AND U15796 ( .A(n17233), .B(n17235), .Z(n17234) );
  XNOR U15797 ( .A(n17236), .B(n17237), .Z(n15933) );
  AND U15798 ( .A(n17236), .B(n17238), .Z(n17237) );
  XNOR U15799 ( .A(n17239), .B(n17240), .Z(n15936) );
  AND U15800 ( .A(n17239), .B(n17241), .Z(n17240) );
  XNOR U15801 ( .A(n17242), .B(n17243), .Z(n15939) );
  AND U15802 ( .A(n17242), .B(n17244), .Z(n17243) );
  XNOR U15803 ( .A(n17245), .B(n17246), .Z(n15942) );
  AND U15804 ( .A(n17245), .B(n17247), .Z(n17246) );
  XNOR U15805 ( .A(n17248), .B(n17249), .Z(n15945) );
  AND U15806 ( .A(n17248), .B(n17250), .Z(n17249) );
  XNOR U15807 ( .A(n17251), .B(n17252), .Z(n15948) );
  AND U15808 ( .A(n17251), .B(n17253), .Z(n17252) );
  XNOR U15809 ( .A(n17254), .B(n17255), .Z(n15951) );
  AND U15810 ( .A(n17254), .B(n17256), .Z(n17255) );
  XNOR U15811 ( .A(n17257), .B(n17258), .Z(n15954) );
  AND U15812 ( .A(n17257), .B(n17259), .Z(n17258) );
  XNOR U15813 ( .A(n17260), .B(n17261), .Z(n15957) );
  AND U15814 ( .A(n17260), .B(n17262), .Z(n17261) );
  XNOR U15815 ( .A(n17263), .B(n17264), .Z(n15960) );
  AND U15816 ( .A(n17263), .B(n17265), .Z(n17264) );
  XNOR U15817 ( .A(n17266), .B(n17267), .Z(n15963) );
  AND U15818 ( .A(n17266), .B(n17268), .Z(n17267) );
  XNOR U15819 ( .A(n17269), .B(n17270), .Z(n15966) );
  AND U15820 ( .A(n17269), .B(n17271), .Z(n17270) );
  XNOR U15821 ( .A(n17272), .B(n17273), .Z(n15969) );
  AND U15822 ( .A(n17272), .B(n17274), .Z(n17273) );
  XNOR U15823 ( .A(n17275), .B(n17276), .Z(n15972) );
  AND U15824 ( .A(n17275), .B(n17277), .Z(n17276) );
  XNOR U15825 ( .A(n17278), .B(n17279), .Z(n15975) );
  AND U15826 ( .A(n17278), .B(n17280), .Z(n17279) );
  XNOR U15827 ( .A(n17281), .B(n17282), .Z(n15978) );
  AND U15828 ( .A(n17281), .B(n17283), .Z(n17282) );
  XNOR U15829 ( .A(n17284), .B(n17285), .Z(n15981) );
  AND U15830 ( .A(n17284), .B(n17286), .Z(n17285) );
  XNOR U15831 ( .A(n17287), .B(n17288), .Z(n15984) );
  AND U15832 ( .A(n17287), .B(n17289), .Z(n17288) );
  XNOR U15833 ( .A(n17290), .B(n17291), .Z(n15987) );
  AND U15834 ( .A(n17290), .B(n17292), .Z(n17291) );
  XNOR U15835 ( .A(n17293), .B(n17294), .Z(n15990) );
  AND U15836 ( .A(n17293), .B(n17295), .Z(n17294) );
  XNOR U15837 ( .A(n17296), .B(n17297), .Z(n15993) );
  AND U15838 ( .A(n17296), .B(n17298), .Z(n17297) );
  XNOR U15839 ( .A(n17299), .B(n17300), .Z(n15996) );
  AND U15840 ( .A(n17299), .B(n17301), .Z(n17300) );
  XNOR U15841 ( .A(n17302), .B(n17303), .Z(n15999) );
  AND U15842 ( .A(n17302), .B(n17304), .Z(n17303) );
  XNOR U15843 ( .A(n17305), .B(n17306), .Z(n16002) );
  AND U15844 ( .A(n17305), .B(n17307), .Z(n17306) );
  XNOR U15845 ( .A(n17308), .B(n17309), .Z(n16005) );
  AND U15846 ( .A(n17308), .B(n17310), .Z(n17309) );
  XNOR U15847 ( .A(n17311), .B(n17312), .Z(n16008) );
  AND U15848 ( .A(n17311), .B(n17313), .Z(n17312) );
  XNOR U15849 ( .A(n17314), .B(n17315), .Z(n16011) );
  AND U15850 ( .A(n17314), .B(n17316), .Z(n17315) );
  XNOR U15851 ( .A(n17317), .B(n17318), .Z(n16014) );
  AND U15852 ( .A(n17317), .B(n17319), .Z(n17318) );
  XNOR U15853 ( .A(n17320), .B(n17321), .Z(n16017) );
  AND U15854 ( .A(n17320), .B(n17322), .Z(n17321) );
  XNOR U15855 ( .A(n17323), .B(n17324), .Z(n16020) );
  AND U15856 ( .A(n17323), .B(n17325), .Z(n17324) );
  XNOR U15857 ( .A(n17326), .B(n17327), .Z(n16023) );
  AND U15858 ( .A(n17326), .B(n17328), .Z(n17327) );
  XNOR U15859 ( .A(n17329), .B(n17330), .Z(n16026) );
  AND U15860 ( .A(n17329), .B(n17331), .Z(n17330) );
  XNOR U15861 ( .A(n17332), .B(n17333), .Z(n16029) );
  AND U15862 ( .A(n17332), .B(n17334), .Z(n17333) );
  XNOR U15863 ( .A(n17335), .B(n17336), .Z(n16032) );
  AND U15864 ( .A(n17335), .B(n17337), .Z(n17336) );
  XNOR U15865 ( .A(n17338), .B(n17339), .Z(n16035) );
  AND U15866 ( .A(n17338), .B(n17340), .Z(n17339) );
  XNOR U15867 ( .A(n17341), .B(n17342), .Z(n16038) );
  AND U15868 ( .A(n17341), .B(n17343), .Z(n17342) );
  XNOR U15869 ( .A(n17344), .B(n17345), .Z(n16041) );
  AND U15870 ( .A(n17344), .B(n17346), .Z(n17345) );
  XNOR U15871 ( .A(n17347), .B(n17348), .Z(n16044) );
  AND U15872 ( .A(n17347), .B(n17349), .Z(n17348) );
  XNOR U15873 ( .A(n17350), .B(n17351), .Z(n16047) );
  AND U15874 ( .A(n17350), .B(n17352), .Z(n17351) );
  XNOR U15875 ( .A(n17353), .B(n17354), .Z(n16050) );
  AND U15876 ( .A(n17353), .B(n17355), .Z(n17354) );
  XNOR U15877 ( .A(n17356), .B(n17357), .Z(n16053) );
  AND U15878 ( .A(n17356), .B(n17358), .Z(n17357) );
  XNOR U15879 ( .A(n17359), .B(n17360), .Z(n16056) );
  AND U15880 ( .A(n17359), .B(n17361), .Z(n17360) );
  XNOR U15881 ( .A(n17362), .B(n17363), .Z(n16059) );
  AND U15882 ( .A(n17362), .B(n17364), .Z(n17363) );
  XNOR U15883 ( .A(n17365), .B(n17366), .Z(n16062) );
  AND U15884 ( .A(n17365), .B(n17367), .Z(n17366) );
  XNOR U15885 ( .A(n17368), .B(n17369), .Z(n16065) );
  AND U15886 ( .A(n17368), .B(n17370), .Z(n17369) );
  XNOR U15887 ( .A(n17371), .B(n17372), .Z(n16068) );
  AND U15888 ( .A(n17371), .B(n17373), .Z(n17372) );
  XNOR U15889 ( .A(n17374), .B(n17375), .Z(n16071) );
  AND U15890 ( .A(n17374), .B(n17376), .Z(n17375) );
  XNOR U15891 ( .A(n17377), .B(n17378), .Z(n16074) );
  AND U15892 ( .A(n17377), .B(n17379), .Z(n17378) );
  XNOR U15893 ( .A(n17380), .B(n17381), .Z(n16077) );
  AND U15894 ( .A(n17380), .B(n17382), .Z(n17381) );
  XNOR U15895 ( .A(n17383), .B(n17384), .Z(n16080) );
  AND U15896 ( .A(n17383), .B(n17385), .Z(n17384) );
  XNOR U15897 ( .A(n17386), .B(n17387), .Z(n16083) );
  AND U15898 ( .A(n17386), .B(n17388), .Z(n17387) );
  XNOR U15899 ( .A(n17389), .B(n17390), .Z(n16086) );
  AND U15900 ( .A(n17389), .B(n17391), .Z(n17390) );
  XNOR U15901 ( .A(n17392), .B(n17393), .Z(n16089) );
  AND U15902 ( .A(n17392), .B(n17394), .Z(n17393) );
  XNOR U15903 ( .A(n17395), .B(n17396), .Z(n16092) );
  AND U15904 ( .A(n17395), .B(n17397), .Z(n17396) );
  XNOR U15905 ( .A(n17398), .B(n17399), .Z(n16095) );
  AND U15906 ( .A(n17398), .B(n17400), .Z(n17399) );
  XNOR U15907 ( .A(n17401), .B(n17402), .Z(n16098) );
  AND U15908 ( .A(n17401), .B(n17403), .Z(n17402) );
  XNOR U15909 ( .A(n17404), .B(n17405), .Z(n16101) );
  AND U15910 ( .A(n17404), .B(n17406), .Z(n17405) );
  XNOR U15911 ( .A(n17407), .B(n17408), .Z(n16104) );
  AND U15912 ( .A(n17407), .B(n17409), .Z(n17408) );
  XNOR U15913 ( .A(n17410), .B(n17411), .Z(n16107) );
  AND U15914 ( .A(n17410), .B(n17412), .Z(n17411) );
  XNOR U15915 ( .A(n17413), .B(n17414), .Z(n16110) );
  AND U15916 ( .A(n17413), .B(n17415), .Z(n17414) );
  XNOR U15917 ( .A(n17416), .B(n17417), .Z(n16113) );
  AND U15918 ( .A(n17416), .B(n17418), .Z(n17417) );
  XNOR U15919 ( .A(n17419), .B(n17420), .Z(n16116) );
  AND U15920 ( .A(n17419), .B(n17421), .Z(n17420) );
  XNOR U15921 ( .A(n17422), .B(n17423), .Z(n16119) );
  AND U15922 ( .A(n17422), .B(n17424), .Z(n17423) );
  XNOR U15923 ( .A(n17425), .B(n17426), .Z(n16122) );
  AND U15924 ( .A(n17425), .B(n17427), .Z(n17426) );
  XNOR U15925 ( .A(n17428), .B(n17429), .Z(n16125) );
  AND U15926 ( .A(n17428), .B(n17430), .Z(n17429) );
  XNOR U15927 ( .A(n17431), .B(n17432), .Z(n16128) );
  AND U15928 ( .A(n17431), .B(n17433), .Z(n17432) );
  XNOR U15929 ( .A(n17434), .B(n17435), .Z(n16131) );
  AND U15930 ( .A(n17434), .B(n17436), .Z(n17435) );
  XNOR U15931 ( .A(n17437), .B(n17438), .Z(n16134) );
  AND U15932 ( .A(n17437), .B(n17439), .Z(n17438) );
  XNOR U15933 ( .A(n17440), .B(n17441), .Z(n16137) );
  AND U15934 ( .A(n17440), .B(n17442), .Z(n17441) );
  XNOR U15935 ( .A(n17443), .B(n17444), .Z(n16140) );
  AND U15936 ( .A(n17443), .B(n17445), .Z(n17444) );
  XNOR U15937 ( .A(n17446), .B(n17447), .Z(n16143) );
  AND U15938 ( .A(n17446), .B(n17448), .Z(n17447) );
  XNOR U15939 ( .A(n17449), .B(n17450), .Z(n16146) );
  AND U15940 ( .A(n17449), .B(n17451), .Z(n17450) );
  XNOR U15941 ( .A(n17452), .B(n17453), .Z(n16149) );
  AND U15942 ( .A(n17452), .B(n17454), .Z(n17453) );
  XNOR U15943 ( .A(n17455), .B(n17456), .Z(n16152) );
  AND U15944 ( .A(n17455), .B(n17457), .Z(n17456) );
  XNOR U15945 ( .A(n17458), .B(n17459), .Z(n16155) );
  AND U15946 ( .A(n17458), .B(n17460), .Z(n17459) );
  XNOR U15947 ( .A(n17461), .B(n17462), .Z(n16158) );
  AND U15948 ( .A(n17461), .B(n17463), .Z(n17462) );
  XNOR U15949 ( .A(n17464), .B(n17465), .Z(n16161) );
  AND U15950 ( .A(n17464), .B(n17466), .Z(n17465) );
  XNOR U15951 ( .A(n17467), .B(n17468), .Z(n16164) );
  AND U15952 ( .A(n17467), .B(n17469), .Z(n17468) );
  XNOR U15953 ( .A(n17470), .B(n17471), .Z(n16167) );
  AND U15954 ( .A(n17470), .B(n17472), .Z(n17471) );
  XNOR U15955 ( .A(n17473), .B(n17474), .Z(n16170) );
  AND U15956 ( .A(n17473), .B(n17475), .Z(n17474) );
  XNOR U15957 ( .A(n17476), .B(n17477), .Z(n16173) );
  AND U15958 ( .A(n17476), .B(n17478), .Z(n17477) );
  XNOR U15959 ( .A(n17479), .B(n17480), .Z(n16176) );
  AND U15960 ( .A(n17479), .B(n17481), .Z(n17480) );
  XNOR U15961 ( .A(n17482), .B(n17483), .Z(n16179) );
  AND U15962 ( .A(n17482), .B(n17484), .Z(n17483) );
  XNOR U15963 ( .A(n17485), .B(n17486), .Z(n16182) );
  AND U15964 ( .A(n17485), .B(n17487), .Z(n17486) );
  IV U15965 ( .A(n16187), .Z(n16185) );
  XNOR U15966 ( .A(n17488), .B(n17489), .Z(n16187) );
  AND U15967 ( .A(n17488), .B(n119), .Z(n17489) );
  XOR U15968 ( .A(n17490), .B(n17491), .Z(n16188) );
  AND U15969 ( .A(n17492), .B(n17493), .Z(n17491) );
  XOR U15970 ( .A(n123), .B(n17490), .Z(n17493) );
  XOR U15971 ( .A(n16838), .B(n16839), .Z(n123) );
  AND U15972 ( .A(n17494), .B(n17495), .Z(n16839) );
  XOR U15973 ( .A(n16835), .B(n16836), .Z(n16838) );
  AND U15974 ( .A(n17496), .B(n17497), .Z(n16836) );
  XOR U15975 ( .A(n16832), .B(n16833), .Z(n16835) );
  AND U15976 ( .A(n17498), .B(n17499), .Z(n16833) );
  XOR U15977 ( .A(n16829), .B(n16830), .Z(n16832) );
  AND U15978 ( .A(n17500), .B(n17501), .Z(n16830) );
  XOR U15979 ( .A(n16826), .B(n16827), .Z(n16829) );
  AND U15980 ( .A(n17502), .B(n17503), .Z(n16827) );
  XOR U15981 ( .A(n16823), .B(n16824), .Z(n16826) );
  AND U15982 ( .A(n17504), .B(n17505), .Z(n16824) );
  XOR U15983 ( .A(n16820), .B(n16821), .Z(n16823) );
  AND U15984 ( .A(n17506), .B(n17507), .Z(n16821) );
  XOR U15985 ( .A(n16817), .B(n16818), .Z(n16820) );
  AND U15986 ( .A(n17508), .B(n17509), .Z(n16818) );
  XOR U15987 ( .A(n16814), .B(n16815), .Z(n16817) );
  AND U15988 ( .A(n17510), .B(n17511), .Z(n16815) );
  XOR U15989 ( .A(n16811), .B(n16812), .Z(n16814) );
  AND U15990 ( .A(n17512), .B(n17513), .Z(n16812) );
  XOR U15991 ( .A(n16808), .B(n16809), .Z(n16811) );
  AND U15992 ( .A(n17514), .B(n17515), .Z(n16809) );
  XOR U15993 ( .A(n16805), .B(n16806), .Z(n16808) );
  AND U15994 ( .A(n17516), .B(n17517), .Z(n16806) );
  XOR U15995 ( .A(n16802), .B(n16803), .Z(n16805) );
  AND U15996 ( .A(n17518), .B(n17519), .Z(n16803) );
  XOR U15997 ( .A(n16799), .B(n16800), .Z(n16802) );
  AND U15998 ( .A(n17520), .B(n17521), .Z(n16800) );
  XOR U15999 ( .A(n16796), .B(n16797), .Z(n16799) );
  AND U16000 ( .A(n17522), .B(n17523), .Z(n16797) );
  XOR U16001 ( .A(n16793), .B(n16794), .Z(n16796) );
  AND U16002 ( .A(n17524), .B(n17525), .Z(n16794) );
  XOR U16003 ( .A(n16790), .B(n16791), .Z(n16793) );
  AND U16004 ( .A(n17526), .B(n17527), .Z(n16791) );
  XOR U16005 ( .A(n16787), .B(n16788), .Z(n16790) );
  AND U16006 ( .A(n17528), .B(n17529), .Z(n16788) );
  XOR U16007 ( .A(n16784), .B(n16785), .Z(n16787) );
  AND U16008 ( .A(n17530), .B(n17531), .Z(n16785) );
  XOR U16009 ( .A(n16781), .B(n16782), .Z(n16784) );
  AND U16010 ( .A(n17532), .B(n17533), .Z(n16782) );
  XOR U16011 ( .A(n16778), .B(n16779), .Z(n16781) );
  AND U16012 ( .A(n17534), .B(n17535), .Z(n16779) );
  XOR U16013 ( .A(n16775), .B(n16776), .Z(n16778) );
  AND U16014 ( .A(n17536), .B(n17537), .Z(n16776) );
  XOR U16015 ( .A(n16772), .B(n16773), .Z(n16775) );
  AND U16016 ( .A(n17538), .B(n17539), .Z(n16773) );
  XOR U16017 ( .A(n16769), .B(n16770), .Z(n16772) );
  AND U16018 ( .A(n17540), .B(n17541), .Z(n16770) );
  XOR U16019 ( .A(n16766), .B(n16767), .Z(n16769) );
  AND U16020 ( .A(n17542), .B(n17543), .Z(n16767) );
  XOR U16021 ( .A(n16763), .B(n16764), .Z(n16766) );
  AND U16022 ( .A(n17544), .B(n17545), .Z(n16764) );
  XOR U16023 ( .A(n16760), .B(n16761), .Z(n16763) );
  AND U16024 ( .A(n17546), .B(n17547), .Z(n16761) );
  XOR U16025 ( .A(n16757), .B(n16758), .Z(n16760) );
  AND U16026 ( .A(n17548), .B(n17549), .Z(n16758) );
  XOR U16027 ( .A(n16754), .B(n16755), .Z(n16757) );
  AND U16028 ( .A(n17550), .B(n17551), .Z(n16755) );
  XOR U16029 ( .A(n16751), .B(n16752), .Z(n16754) );
  AND U16030 ( .A(n17552), .B(n17553), .Z(n16752) );
  XOR U16031 ( .A(n16748), .B(n16749), .Z(n16751) );
  AND U16032 ( .A(n17554), .B(n17555), .Z(n16749) );
  XOR U16033 ( .A(n16745), .B(n16746), .Z(n16748) );
  AND U16034 ( .A(n17556), .B(n17557), .Z(n16746) );
  XOR U16035 ( .A(n16742), .B(n16743), .Z(n16745) );
  AND U16036 ( .A(n17558), .B(n17559), .Z(n16743) );
  XOR U16037 ( .A(n16739), .B(n16740), .Z(n16742) );
  AND U16038 ( .A(n17560), .B(n17561), .Z(n16740) );
  XOR U16039 ( .A(n16736), .B(n16737), .Z(n16739) );
  AND U16040 ( .A(n17562), .B(n17563), .Z(n16737) );
  XOR U16041 ( .A(n16733), .B(n16734), .Z(n16736) );
  AND U16042 ( .A(n17564), .B(n17565), .Z(n16734) );
  XOR U16043 ( .A(n16730), .B(n16731), .Z(n16733) );
  AND U16044 ( .A(n17566), .B(n17567), .Z(n16731) );
  XOR U16045 ( .A(n16727), .B(n16728), .Z(n16730) );
  AND U16046 ( .A(n17568), .B(n17569), .Z(n16728) );
  XOR U16047 ( .A(n16724), .B(n16725), .Z(n16727) );
  AND U16048 ( .A(n17570), .B(n17571), .Z(n16725) );
  XOR U16049 ( .A(n16721), .B(n16722), .Z(n16724) );
  AND U16050 ( .A(n17572), .B(n17573), .Z(n16722) );
  XOR U16051 ( .A(n16718), .B(n16719), .Z(n16721) );
  AND U16052 ( .A(n17574), .B(n17575), .Z(n16719) );
  XOR U16053 ( .A(n16715), .B(n16716), .Z(n16718) );
  AND U16054 ( .A(n17576), .B(n17577), .Z(n16716) );
  XOR U16055 ( .A(n16712), .B(n16713), .Z(n16715) );
  AND U16056 ( .A(n17578), .B(n17579), .Z(n16713) );
  XOR U16057 ( .A(n16709), .B(n16710), .Z(n16712) );
  AND U16058 ( .A(n17580), .B(n17581), .Z(n16710) );
  XOR U16059 ( .A(n16706), .B(n16707), .Z(n16709) );
  AND U16060 ( .A(n17582), .B(n17583), .Z(n16707) );
  XOR U16061 ( .A(n16703), .B(n16704), .Z(n16706) );
  AND U16062 ( .A(n17584), .B(n17585), .Z(n16704) );
  XOR U16063 ( .A(n16700), .B(n16701), .Z(n16703) );
  AND U16064 ( .A(n17586), .B(n17587), .Z(n16701) );
  XOR U16065 ( .A(n16697), .B(n16698), .Z(n16700) );
  AND U16066 ( .A(n17588), .B(n17589), .Z(n16698) );
  XOR U16067 ( .A(n16694), .B(n16695), .Z(n16697) );
  AND U16068 ( .A(n17590), .B(n17591), .Z(n16695) );
  XOR U16069 ( .A(n16691), .B(n16692), .Z(n16694) );
  AND U16070 ( .A(n17592), .B(n17593), .Z(n16692) );
  XOR U16071 ( .A(n16688), .B(n16689), .Z(n16691) );
  AND U16072 ( .A(n17594), .B(n17595), .Z(n16689) );
  XOR U16073 ( .A(n16685), .B(n16686), .Z(n16688) );
  AND U16074 ( .A(n17596), .B(n17597), .Z(n16686) );
  XOR U16075 ( .A(n16682), .B(n16683), .Z(n16685) );
  AND U16076 ( .A(n17598), .B(n17599), .Z(n16683) );
  XOR U16077 ( .A(n16679), .B(n16680), .Z(n16682) );
  AND U16078 ( .A(n17600), .B(n17601), .Z(n16680) );
  XOR U16079 ( .A(n16676), .B(n16677), .Z(n16679) );
  AND U16080 ( .A(n17602), .B(n17603), .Z(n16677) );
  XOR U16081 ( .A(n16673), .B(n16674), .Z(n16676) );
  AND U16082 ( .A(n17604), .B(n17605), .Z(n16674) );
  XOR U16083 ( .A(n16670), .B(n16671), .Z(n16673) );
  AND U16084 ( .A(n17606), .B(n17607), .Z(n16671) );
  XOR U16085 ( .A(n16667), .B(n16668), .Z(n16670) );
  AND U16086 ( .A(n17608), .B(n17609), .Z(n16668) );
  XOR U16087 ( .A(n16664), .B(n16665), .Z(n16667) );
  AND U16088 ( .A(n17610), .B(n17611), .Z(n16665) );
  XOR U16089 ( .A(n16661), .B(n16662), .Z(n16664) );
  AND U16090 ( .A(n17612), .B(n17613), .Z(n16662) );
  XOR U16091 ( .A(n16658), .B(n16659), .Z(n16661) );
  AND U16092 ( .A(n17614), .B(n17615), .Z(n16659) );
  XOR U16093 ( .A(n16655), .B(n16656), .Z(n16658) );
  AND U16094 ( .A(n17616), .B(n17617), .Z(n16656) );
  XOR U16095 ( .A(n16652), .B(n16653), .Z(n16655) );
  AND U16096 ( .A(n17618), .B(n17619), .Z(n16653) );
  XOR U16097 ( .A(n16649), .B(n16650), .Z(n16652) );
  AND U16098 ( .A(n17620), .B(n17621), .Z(n16650) );
  XOR U16099 ( .A(n16646), .B(n16647), .Z(n16649) );
  AND U16100 ( .A(n17622), .B(n17623), .Z(n16647) );
  XOR U16101 ( .A(n16643), .B(n16644), .Z(n16646) );
  AND U16102 ( .A(n17624), .B(n17625), .Z(n16644) );
  XOR U16103 ( .A(n16640), .B(n16641), .Z(n16643) );
  AND U16104 ( .A(n17626), .B(n17627), .Z(n16641) );
  XOR U16105 ( .A(n16637), .B(n16638), .Z(n16640) );
  AND U16106 ( .A(n17628), .B(n17629), .Z(n16638) );
  XOR U16107 ( .A(n16634), .B(n16635), .Z(n16637) );
  AND U16108 ( .A(n17630), .B(n17631), .Z(n16635) );
  XOR U16109 ( .A(n16631), .B(n16632), .Z(n16634) );
  AND U16110 ( .A(n17632), .B(n17633), .Z(n16632) );
  XOR U16111 ( .A(n16628), .B(n16629), .Z(n16631) );
  AND U16112 ( .A(n17634), .B(n17635), .Z(n16629) );
  XOR U16113 ( .A(n16625), .B(n16626), .Z(n16628) );
  AND U16114 ( .A(n17636), .B(n17637), .Z(n16626) );
  XOR U16115 ( .A(n16622), .B(n16623), .Z(n16625) );
  AND U16116 ( .A(n17638), .B(n17639), .Z(n16623) );
  XOR U16117 ( .A(n16619), .B(n16620), .Z(n16622) );
  AND U16118 ( .A(n17640), .B(n17641), .Z(n16620) );
  XOR U16119 ( .A(n16616), .B(n16617), .Z(n16619) );
  AND U16120 ( .A(n17642), .B(n17643), .Z(n16617) );
  XOR U16121 ( .A(n16613), .B(n16614), .Z(n16616) );
  AND U16122 ( .A(n17644), .B(n17645), .Z(n16614) );
  XOR U16123 ( .A(n16610), .B(n16611), .Z(n16613) );
  AND U16124 ( .A(n17646), .B(n17647), .Z(n16611) );
  XOR U16125 ( .A(n16607), .B(n16608), .Z(n16610) );
  AND U16126 ( .A(n17648), .B(n17649), .Z(n16608) );
  XOR U16127 ( .A(n16604), .B(n16605), .Z(n16607) );
  AND U16128 ( .A(n17650), .B(n17651), .Z(n16605) );
  XOR U16129 ( .A(n16601), .B(n16602), .Z(n16604) );
  AND U16130 ( .A(n17652), .B(n17653), .Z(n16602) );
  XOR U16131 ( .A(n16598), .B(n16599), .Z(n16601) );
  AND U16132 ( .A(n17654), .B(n17655), .Z(n16599) );
  XOR U16133 ( .A(n16595), .B(n16596), .Z(n16598) );
  AND U16134 ( .A(n17656), .B(n17657), .Z(n16596) );
  XOR U16135 ( .A(n16592), .B(n16593), .Z(n16595) );
  AND U16136 ( .A(n17658), .B(n17659), .Z(n16593) );
  XOR U16137 ( .A(n16589), .B(n16590), .Z(n16592) );
  AND U16138 ( .A(n17660), .B(n17661), .Z(n16590) );
  XOR U16139 ( .A(n16586), .B(n16587), .Z(n16589) );
  AND U16140 ( .A(n17662), .B(n17663), .Z(n16587) );
  XOR U16141 ( .A(n16583), .B(n16584), .Z(n16586) );
  AND U16142 ( .A(n17664), .B(n17665), .Z(n16584) );
  XOR U16143 ( .A(n16580), .B(n16581), .Z(n16583) );
  AND U16144 ( .A(n17666), .B(n17667), .Z(n16581) );
  XOR U16145 ( .A(n16577), .B(n16578), .Z(n16580) );
  AND U16146 ( .A(n17668), .B(n17669), .Z(n16578) );
  XOR U16147 ( .A(n16574), .B(n16575), .Z(n16577) );
  AND U16148 ( .A(n17670), .B(n17671), .Z(n16575) );
  XOR U16149 ( .A(n16571), .B(n16572), .Z(n16574) );
  AND U16150 ( .A(n17672), .B(n17673), .Z(n16572) );
  XOR U16151 ( .A(n16568), .B(n16569), .Z(n16571) );
  AND U16152 ( .A(n17674), .B(n17675), .Z(n16569) );
  XOR U16153 ( .A(n16565), .B(n16566), .Z(n16568) );
  AND U16154 ( .A(n17676), .B(n17677), .Z(n16566) );
  XOR U16155 ( .A(n16562), .B(n16563), .Z(n16565) );
  AND U16156 ( .A(n17678), .B(n17679), .Z(n16563) );
  XOR U16157 ( .A(n16559), .B(n16560), .Z(n16562) );
  AND U16158 ( .A(n17680), .B(n17681), .Z(n16560) );
  XOR U16159 ( .A(n16556), .B(n16557), .Z(n16559) );
  AND U16160 ( .A(n17682), .B(n17683), .Z(n16557) );
  XOR U16161 ( .A(n16553), .B(n16554), .Z(n16556) );
  AND U16162 ( .A(n17684), .B(n17685), .Z(n16554) );
  XOR U16163 ( .A(n16550), .B(n16551), .Z(n16553) );
  AND U16164 ( .A(n17686), .B(n17687), .Z(n16551) );
  XOR U16165 ( .A(n16547), .B(n16548), .Z(n16550) );
  AND U16166 ( .A(n17688), .B(n17689), .Z(n16548) );
  XOR U16167 ( .A(n16544), .B(n16545), .Z(n16547) );
  AND U16168 ( .A(n17690), .B(n17691), .Z(n16545) );
  XOR U16169 ( .A(n16541), .B(n16542), .Z(n16544) );
  AND U16170 ( .A(n17692), .B(n17693), .Z(n16542) );
  XOR U16171 ( .A(n16538), .B(n16539), .Z(n16541) );
  AND U16172 ( .A(n17694), .B(n17695), .Z(n16539) );
  XOR U16173 ( .A(n16535), .B(n16536), .Z(n16538) );
  AND U16174 ( .A(n17696), .B(n17697), .Z(n16536) );
  XOR U16175 ( .A(n16532), .B(n16533), .Z(n16535) );
  AND U16176 ( .A(n17698), .B(n17699), .Z(n16533) );
  XOR U16177 ( .A(n16529), .B(n16530), .Z(n16532) );
  AND U16178 ( .A(n17700), .B(n17701), .Z(n16530) );
  XOR U16179 ( .A(n16526), .B(n16527), .Z(n16529) );
  AND U16180 ( .A(n17702), .B(n17703), .Z(n16527) );
  XOR U16181 ( .A(n16523), .B(n16524), .Z(n16526) );
  AND U16182 ( .A(n17704), .B(n17705), .Z(n16524) );
  XOR U16183 ( .A(n16520), .B(n16521), .Z(n16523) );
  AND U16184 ( .A(n17706), .B(n17707), .Z(n16521) );
  XOR U16185 ( .A(n16517), .B(n16518), .Z(n16520) );
  AND U16186 ( .A(n17708), .B(n17709), .Z(n16518) );
  XOR U16187 ( .A(n16514), .B(n16515), .Z(n16517) );
  AND U16188 ( .A(n17710), .B(n17711), .Z(n16515) );
  XOR U16189 ( .A(n16511), .B(n16512), .Z(n16514) );
  AND U16190 ( .A(n17712), .B(n17713), .Z(n16512) );
  XOR U16191 ( .A(n16508), .B(n16509), .Z(n16511) );
  AND U16192 ( .A(n17714), .B(n17715), .Z(n16509) );
  XOR U16193 ( .A(n16505), .B(n16506), .Z(n16508) );
  AND U16194 ( .A(n17716), .B(n17717), .Z(n16506) );
  XOR U16195 ( .A(n16502), .B(n16503), .Z(n16505) );
  AND U16196 ( .A(n17718), .B(n17719), .Z(n16503) );
  XOR U16197 ( .A(n16499), .B(n16500), .Z(n16502) );
  AND U16198 ( .A(n17720), .B(n17721), .Z(n16500) );
  XOR U16199 ( .A(n16496), .B(n16497), .Z(n16499) );
  AND U16200 ( .A(n17722), .B(n17723), .Z(n16497) );
  XOR U16201 ( .A(n16493), .B(n16494), .Z(n16496) );
  AND U16202 ( .A(n17724), .B(n17725), .Z(n16494) );
  XOR U16203 ( .A(n16490), .B(n16491), .Z(n16493) );
  AND U16204 ( .A(n17726), .B(n17727), .Z(n16491) );
  XOR U16205 ( .A(n16487), .B(n16488), .Z(n16490) );
  AND U16206 ( .A(n17728), .B(n17729), .Z(n16488) );
  XOR U16207 ( .A(n16484), .B(n16485), .Z(n16487) );
  AND U16208 ( .A(n17730), .B(n17731), .Z(n16485) );
  XOR U16209 ( .A(n16481), .B(n16482), .Z(n16484) );
  AND U16210 ( .A(n17732), .B(n17733), .Z(n16482) );
  XOR U16211 ( .A(n16478), .B(n16479), .Z(n16481) );
  AND U16212 ( .A(n17734), .B(n17735), .Z(n16479) );
  XOR U16213 ( .A(n16475), .B(n16476), .Z(n16478) );
  AND U16214 ( .A(n17736), .B(n17737), .Z(n16476) );
  XOR U16215 ( .A(n16472), .B(n16473), .Z(n16475) );
  AND U16216 ( .A(n17738), .B(n17739), .Z(n16473) );
  XOR U16217 ( .A(n16469), .B(n16470), .Z(n16472) );
  AND U16218 ( .A(n17740), .B(n17741), .Z(n16470) );
  XOR U16219 ( .A(n16466), .B(n16467), .Z(n16469) );
  AND U16220 ( .A(n17742), .B(n17743), .Z(n16467) );
  XOR U16221 ( .A(n16463), .B(n16464), .Z(n16466) );
  AND U16222 ( .A(n17744), .B(n17745), .Z(n16464) );
  XOR U16223 ( .A(n16460), .B(n16461), .Z(n16463) );
  AND U16224 ( .A(n17746), .B(n17747), .Z(n16461) );
  XOR U16225 ( .A(n16457), .B(n16458), .Z(n16460) );
  AND U16226 ( .A(n17748), .B(n17749), .Z(n16458) );
  XNOR U16227 ( .A(n16454), .B(n16455), .Z(n16457) );
  AND U16228 ( .A(n17750), .B(n17751), .Z(n16455) );
  XOR U16229 ( .A(n17752), .B(n16452), .Z(n16454) );
  IV U16230 ( .A(n17753), .Z(n16452) );
  AND U16231 ( .A(n17754), .B(n17755), .Z(n17753) );
  IV U16232 ( .A(n16451), .Z(n17752) );
  XOR U16233 ( .A(n16192), .B(n16448), .Z(n16451) );
  AND U16234 ( .A(n17756), .B(n17757), .Z(n16448) );
  XOR U16235 ( .A(n16194), .B(n16193), .Z(n16192) );
  AND U16236 ( .A(n17758), .B(n17759), .Z(n16193) );
  XOR U16237 ( .A(n16196), .B(n16195), .Z(n16194) );
  AND U16238 ( .A(n17760), .B(n17761), .Z(n16195) );
  XOR U16239 ( .A(n16198), .B(n16197), .Z(n16196) );
  AND U16240 ( .A(n17762), .B(n17763), .Z(n16197) );
  XOR U16241 ( .A(n16200), .B(n16199), .Z(n16198) );
  AND U16242 ( .A(n17764), .B(n17765), .Z(n16199) );
  XOR U16243 ( .A(n16202), .B(n16201), .Z(n16200) );
  AND U16244 ( .A(n17766), .B(n17767), .Z(n16201) );
  XOR U16245 ( .A(n16204), .B(n16203), .Z(n16202) );
  AND U16246 ( .A(n17768), .B(n17769), .Z(n16203) );
  XOR U16247 ( .A(n16206), .B(n16205), .Z(n16204) );
  AND U16248 ( .A(n17770), .B(n17771), .Z(n16205) );
  XOR U16249 ( .A(n16208), .B(n16207), .Z(n16206) );
  AND U16250 ( .A(n17772), .B(n17773), .Z(n16207) );
  XOR U16251 ( .A(n16210), .B(n16209), .Z(n16208) );
  AND U16252 ( .A(n17774), .B(n17775), .Z(n16209) );
  XOR U16253 ( .A(n16212), .B(n16211), .Z(n16210) );
  AND U16254 ( .A(n17776), .B(n17777), .Z(n16211) );
  XOR U16255 ( .A(n16214), .B(n16213), .Z(n16212) );
  AND U16256 ( .A(n17778), .B(n17779), .Z(n16213) );
  XOR U16257 ( .A(n16216), .B(n16215), .Z(n16214) );
  AND U16258 ( .A(n17780), .B(n17781), .Z(n16215) );
  XOR U16259 ( .A(n16218), .B(n16217), .Z(n16216) );
  AND U16260 ( .A(n17782), .B(n17783), .Z(n16217) );
  XOR U16261 ( .A(n16220), .B(n16219), .Z(n16218) );
  AND U16262 ( .A(n17784), .B(n17785), .Z(n16219) );
  XOR U16263 ( .A(n16222), .B(n16221), .Z(n16220) );
  AND U16264 ( .A(n17786), .B(n17787), .Z(n16221) );
  XOR U16265 ( .A(n16224), .B(n16223), .Z(n16222) );
  AND U16266 ( .A(n17788), .B(n17789), .Z(n16223) );
  XOR U16267 ( .A(n16226), .B(n16225), .Z(n16224) );
  AND U16268 ( .A(n17790), .B(n17791), .Z(n16225) );
  XOR U16269 ( .A(n16228), .B(n16227), .Z(n16226) );
  AND U16270 ( .A(n17792), .B(n17793), .Z(n16227) );
  XOR U16271 ( .A(n16230), .B(n16229), .Z(n16228) );
  AND U16272 ( .A(n17794), .B(n17795), .Z(n16229) );
  XOR U16273 ( .A(n16232), .B(n16231), .Z(n16230) );
  AND U16274 ( .A(n17796), .B(n17797), .Z(n16231) );
  XOR U16275 ( .A(n16234), .B(n16233), .Z(n16232) );
  AND U16276 ( .A(n17798), .B(n17799), .Z(n16233) );
  XOR U16277 ( .A(n16236), .B(n16235), .Z(n16234) );
  AND U16278 ( .A(n17800), .B(n17801), .Z(n16235) );
  XOR U16279 ( .A(n16238), .B(n16237), .Z(n16236) );
  AND U16280 ( .A(n17802), .B(n17803), .Z(n16237) );
  XOR U16281 ( .A(n16240), .B(n16239), .Z(n16238) );
  AND U16282 ( .A(n17804), .B(n17805), .Z(n16239) );
  XOR U16283 ( .A(n16242), .B(n16241), .Z(n16240) );
  AND U16284 ( .A(n17806), .B(n17807), .Z(n16241) );
  XOR U16285 ( .A(n16244), .B(n16243), .Z(n16242) );
  AND U16286 ( .A(n17808), .B(n17809), .Z(n16243) );
  XOR U16287 ( .A(n16246), .B(n16245), .Z(n16244) );
  AND U16288 ( .A(n17810), .B(n17811), .Z(n16245) );
  XOR U16289 ( .A(n16248), .B(n16247), .Z(n16246) );
  AND U16290 ( .A(n17812), .B(n17813), .Z(n16247) );
  XOR U16291 ( .A(n16250), .B(n16249), .Z(n16248) );
  AND U16292 ( .A(n17814), .B(n17815), .Z(n16249) );
  XOR U16293 ( .A(n16252), .B(n16251), .Z(n16250) );
  AND U16294 ( .A(n17816), .B(n17817), .Z(n16251) );
  XOR U16295 ( .A(n16254), .B(n16253), .Z(n16252) );
  AND U16296 ( .A(n17818), .B(n17819), .Z(n16253) );
  XOR U16297 ( .A(n16256), .B(n16255), .Z(n16254) );
  AND U16298 ( .A(n17820), .B(n17821), .Z(n16255) );
  XOR U16299 ( .A(n16258), .B(n16257), .Z(n16256) );
  AND U16300 ( .A(n17822), .B(n17823), .Z(n16257) );
  XOR U16301 ( .A(n16260), .B(n16259), .Z(n16258) );
  AND U16302 ( .A(n17824), .B(n17825), .Z(n16259) );
  XOR U16303 ( .A(n16262), .B(n16261), .Z(n16260) );
  AND U16304 ( .A(n17826), .B(n17827), .Z(n16261) );
  XOR U16305 ( .A(n16264), .B(n16263), .Z(n16262) );
  AND U16306 ( .A(n17828), .B(n17829), .Z(n16263) );
  XOR U16307 ( .A(n16266), .B(n16265), .Z(n16264) );
  AND U16308 ( .A(n17830), .B(n17831), .Z(n16265) );
  XOR U16309 ( .A(n16268), .B(n16267), .Z(n16266) );
  AND U16310 ( .A(n17832), .B(n17833), .Z(n16267) );
  XOR U16311 ( .A(n16270), .B(n16269), .Z(n16268) );
  AND U16312 ( .A(n17834), .B(n17835), .Z(n16269) );
  XOR U16313 ( .A(n16272), .B(n16271), .Z(n16270) );
  AND U16314 ( .A(n17836), .B(n17837), .Z(n16271) );
  XOR U16315 ( .A(n16274), .B(n16273), .Z(n16272) );
  AND U16316 ( .A(n17838), .B(n17839), .Z(n16273) );
  XOR U16317 ( .A(n16276), .B(n16275), .Z(n16274) );
  AND U16318 ( .A(n17840), .B(n17841), .Z(n16275) );
  XOR U16319 ( .A(n16278), .B(n16277), .Z(n16276) );
  AND U16320 ( .A(n17842), .B(n17843), .Z(n16277) );
  XOR U16321 ( .A(n16280), .B(n16279), .Z(n16278) );
  AND U16322 ( .A(n17844), .B(n17845), .Z(n16279) );
  XOR U16323 ( .A(n16282), .B(n16281), .Z(n16280) );
  AND U16324 ( .A(n17846), .B(n17847), .Z(n16281) );
  XOR U16325 ( .A(n16284), .B(n16283), .Z(n16282) );
  AND U16326 ( .A(n17848), .B(n17849), .Z(n16283) );
  XOR U16327 ( .A(n16286), .B(n16285), .Z(n16284) );
  AND U16328 ( .A(n17850), .B(n17851), .Z(n16285) );
  XOR U16329 ( .A(n16288), .B(n16287), .Z(n16286) );
  AND U16330 ( .A(n17852), .B(n17853), .Z(n16287) );
  XOR U16331 ( .A(n16290), .B(n16289), .Z(n16288) );
  AND U16332 ( .A(n17854), .B(n17855), .Z(n16289) );
  XOR U16333 ( .A(n16292), .B(n16291), .Z(n16290) );
  AND U16334 ( .A(n17856), .B(n17857), .Z(n16291) );
  XOR U16335 ( .A(n16294), .B(n16293), .Z(n16292) );
  AND U16336 ( .A(n17858), .B(n17859), .Z(n16293) );
  XOR U16337 ( .A(n16296), .B(n16295), .Z(n16294) );
  AND U16338 ( .A(n17860), .B(n17861), .Z(n16295) );
  XOR U16339 ( .A(n16298), .B(n16297), .Z(n16296) );
  AND U16340 ( .A(n17862), .B(n17863), .Z(n16297) );
  XOR U16341 ( .A(n16300), .B(n16299), .Z(n16298) );
  AND U16342 ( .A(n17864), .B(n17865), .Z(n16299) );
  XOR U16343 ( .A(n16302), .B(n16301), .Z(n16300) );
  AND U16344 ( .A(n17866), .B(n17867), .Z(n16301) );
  XOR U16345 ( .A(n16304), .B(n16303), .Z(n16302) );
  AND U16346 ( .A(n17868), .B(n17869), .Z(n16303) );
  XOR U16347 ( .A(n16306), .B(n16305), .Z(n16304) );
  AND U16348 ( .A(n17870), .B(n17871), .Z(n16305) );
  XOR U16349 ( .A(n16308), .B(n16307), .Z(n16306) );
  AND U16350 ( .A(n17872), .B(n17873), .Z(n16307) );
  XOR U16351 ( .A(n16310), .B(n16309), .Z(n16308) );
  AND U16352 ( .A(n17874), .B(n17875), .Z(n16309) );
  XOR U16353 ( .A(n16312), .B(n16311), .Z(n16310) );
  AND U16354 ( .A(n17876), .B(n17877), .Z(n16311) );
  XOR U16355 ( .A(n16314), .B(n16313), .Z(n16312) );
  AND U16356 ( .A(n17878), .B(n17879), .Z(n16313) );
  XOR U16357 ( .A(n16316), .B(n16315), .Z(n16314) );
  AND U16358 ( .A(n17880), .B(n17881), .Z(n16315) );
  XOR U16359 ( .A(n16318), .B(n16317), .Z(n16316) );
  AND U16360 ( .A(n17882), .B(n17883), .Z(n16317) );
  XOR U16361 ( .A(n16320), .B(n16319), .Z(n16318) );
  AND U16362 ( .A(n17884), .B(n17885), .Z(n16319) );
  XOR U16363 ( .A(n16322), .B(n16321), .Z(n16320) );
  AND U16364 ( .A(n17886), .B(n17887), .Z(n16321) );
  XOR U16365 ( .A(n16324), .B(n16323), .Z(n16322) );
  AND U16366 ( .A(n17888), .B(n17889), .Z(n16323) );
  XOR U16367 ( .A(n16326), .B(n16325), .Z(n16324) );
  AND U16368 ( .A(n17890), .B(n17891), .Z(n16325) );
  XOR U16369 ( .A(n16328), .B(n16327), .Z(n16326) );
  AND U16370 ( .A(n17892), .B(n17893), .Z(n16327) );
  XOR U16371 ( .A(n16330), .B(n16329), .Z(n16328) );
  AND U16372 ( .A(n17894), .B(n17895), .Z(n16329) );
  XOR U16373 ( .A(n16332), .B(n16331), .Z(n16330) );
  AND U16374 ( .A(n17896), .B(n17897), .Z(n16331) );
  XOR U16375 ( .A(n16334), .B(n16333), .Z(n16332) );
  AND U16376 ( .A(n17898), .B(n17899), .Z(n16333) );
  XOR U16377 ( .A(n16336), .B(n16335), .Z(n16334) );
  AND U16378 ( .A(n17900), .B(n17901), .Z(n16335) );
  XOR U16379 ( .A(n16338), .B(n16337), .Z(n16336) );
  AND U16380 ( .A(n17902), .B(n17903), .Z(n16337) );
  XOR U16381 ( .A(n16340), .B(n16339), .Z(n16338) );
  AND U16382 ( .A(n17904), .B(n17905), .Z(n16339) );
  XOR U16383 ( .A(n16342), .B(n16341), .Z(n16340) );
  AND U16384 ( .A(n17906), .B(n17907), .Z(n16341) );
  XOR U16385 ( .A(n16344), .B(n16343), .Z(n16342) );
  AND U16386 ( .A(n17908), .B(n17909), .Z(n16343) );
  XOR U16387 ( .A(n16346), .B(n16345), .Z(n16344) );
  AND U16388 ( .A(n17910), .B(n17911), .Z(n16345) );
  XOR U16389 ( .A(n16348), .B(n16347), .Z(n16346) );
  AND U16390 ( .A(n17912), .B(n17913), .Z(n16347) );
  XOR U16391 ( .A(n16350), .B(n16349), .Z(n16348) );
  AND U16392 ( .A(n17914), .B(n17915), .Z(n16349) );
  XOR U16393 ( .A(n16352), .B(n16351), .Z(n16350) );
  AND U16394 ( .A(n17916), .B(n17917), .Z(n16351) );
  XOR U16395 ( .A(n16354), .B(n16353), .Z(n16352) );
  AND U16396 ( .A(n17918), .B(n17919), .Z(n16353) );
  XOR U16397 ( .A(n16356), .B(n16355), .Z(n16354) );
  AND U16398 ( .A(n17920), .B(n17921), .Z(n16355) );
  XOR U16399 ( .A(n16358), .B(n16357), .Z(n16356) );
  AND U16400 ( .A(n17922), .B(n17923), .Z(n16357) );
  XOR U16401 ( .A(n16360), .B(n16359), .Z(n16358) );
  AND U16402 ( .A(n17924), .B(n17925), .Z(n16359) );
  XOR U16403 ( .A(n16362), .B(n16361), .Z(n16360) );
  AND U16404 ( .A(n17926), .B(n17927), .Z(n16361) );
  XOR U16405 ( .A(n16364), .B(n16363), .Z(n16362) );
  AND U16406 ( .A(n17928), .B(n17929), .Z(n16363) );
  XOR U16407 ( .A(n16366), .B(n16365), .Z(n16364) );
  AND U16408 ( .A(n17930), .B(n17931), .Z(n16365) );
  XOR U16409 ( .A(n16368), .B(n16367), .Z(n16366) );
  AND U16410 ( .A(n17932), .B(n17933), .Z(n16367) );
  XOR U16411 ( .A(n16370), .B(n16369), .Z(n16368) );
  AND U16412 ( .A(n17934), .B(n17935), .Z(n16369) );
  XOR U16413 ( .A(n16372), .B(n16371), .Z(n16370) );
  AND U16414 ( .A(n17936), .B(n17937), .Z(n16371) );
  XOR U16415 ( .A(n16374), .B(n16373), .Z(n16372) );
  AND U16416 ( .A(n17938), .B(n17939), .Z(n16373) );
  XOR U16417 ( .A(n16376), .B(n16375), .Z(n16374) );
  AND U16418 ( .A(n17940), .B(n17941), .Z(n16375) );
  XOR U16419 ( .A(n16378), .B(n16377), .Z(n16376) );
  AND U16420 ( .A(n17942), .B(n17943), .Z(n16377) );
  XOR U16421 ( .A(n16380), .B(n16379), .Z(n16378) );
  AND U16422 ( .A(n17944), .B(n17945), .Z(n16379) );
  XOR U16423 ( .A(n16382), .B(n16381), .Z(n16380) );
  AND U16424 ( .A(n17946), .B(n17947), .Z(n16381) );
  XOR U16425 ( .A(n16384), .B(n16383), .Z(n16382) );
  AND U16426 ( .A(n17948), .B(n17949), .Z(n16383) );
  XOR U16427 ( .A(n16386), .B(n16385), .Z(n16384) );
  AND U16428 ( .A(n17950), .B(n17951), .Z(n16385) );
  XOR U16429 ( .A(n16388), .B(n16387), .Z(n16386) );
  AND U16430 ( .A(n17952), .B(n17953), .Z(n16387) );
  XOR U16431 ( .A(n16390), .B(n16389), .Z(n16388) );
  AND U16432 ( .A(n17954), .B(n17955), .Z(n16389) );
  XOR U16433 ( .A(n16392), .B(n16391), .Z(n16390) );
  AND U16434 ( .A(n17956), .B(n17957), .Z(n16391) );
  XOR U16435 ( .A(n16394), .B(n16393), .Z(n16392) );
  AND U16436 ( .A(n17958), .B(n17959), .Z(n16393) );
  XOR U16437 ( .A(n16396), .B(n16395), .Z(n16394) );
  AND U16438 ( .A(n17960), .B(n17961), .Z(n16395) );
  XOR U16439 ( .A(n16398), .B(n16397), .Z(n16396) );
  AND U16440 ( .A(n17962), .B(n17963), .Z(n16397) );
  XOR U16441 ( .A(n16400), .B(n16399), .Z(n16398) );
  AND U16442 ( .A(n17964), .B(n17965), .Z(n16399) );
  XOR U16443 ( .A(n16402), .B(n16401), .Z(n16400) );
  AND U16444 ( .A(n17966), .B(n17967), .Z(n16401) );
  XOR U16445 ( .A(n16404), .B(n16403), .Z(n16402) );
  AND U16446 ( .A(n17968), .B(n17969), .Z(n16403) );
  XOR U16447 ( .A(n16406), .B(n16405), .Z(n16404) );
  AND U16448 ( .A(n17970), .B(n17971), .Z(n16405) );
  XOR U16449 ( .A(n16408), .B(n16407), .Z(n16406) );
  AND U16450 ( .A(n17972), .B(n17973), .Z(n16407) );
  XOR U16451 ( .A(n16410), .B(n16409), .Z(n16408) );
  AND U16452 ( .A(n17974), .B(n17975), .Z(n16409) );
  XOR U16453 ( .A(n16412), .B(n16411), .Z(n16410) );
  AND U16454 ( .A(n17976), .B(n17977), .Z(n16411) );
  XOR U16455 ( .A(n16414), .B(n16413), .Z(n16412) );
  AND U16456 ( .A(n17978), .B(n17979), .Z(n16413) );
  XOR U16457 ( .A(n16416), .B(n16415), .Z(n16414) );
  AND U16458 ( .A(n17980), .B(n17981), .Z(n16415) );
  XOR U16459 ( .A(n16444), .B(n16417), .Z(n16416) );
  AND U16460 ( .A(n17982), .B(n17983), .Z(n16417) );
  XOR U16461 ( .A(n16446), .B(n16445), .Z(n16444) );
  AND U16462 ( .A(n17984), .B(n17985), .Z(n16445) );
  XOR U16463 ( .A(n16425), .B(n16447), .Z(n16446) );
  AND U16464 ( .A(n17986), .B(n17987), .Z(n16447) );
  XOR U16465 ( .A(n16421), .B(n16426), .Z(n16425) );
  AND U16466 ( .A(n17988), .B(n17989), .Z(n16426) );
  XOR U16467 ( .A(n16423), .B(n16422), .Z(n16421) );
  AND U16468 ( .A(n17990), .B(n17991), .Z(n16422) );
  XNOR U16469 ( .A(n16433), .B(n16424), .Z(n16423) );
  AND U16470 ( .A(n17992), .B(n17993), .Z(n16424) );
  XOR U16471 ( .A(n16443), .B(n16432), .Z(n16433) );
  AND U16472 ( .A(n17994), .B(n17995), .Z(n16432) );
  XNOR U16473 ( .A(n17996), .B(n16438), .Z(n16443) );
  XOR U16474 ( .A(n16439), .B(n17997), .Z(n16438) );
  AND U16475 ( .A(n17998), .B(n17999), .Z(n17997) );
  XOR U16476 ( .A(n18000), .B(n18001), .Z(n16439) );
  NOR U16477 ( .A(n18002), .B(n18003), .Z(n18001) );
  AND U16478 ( .A(n18004), .B(n18005), .Z(n18003) );
  AND U16479 ( .A(n18006), .B(n18007), .Z(n18002) );
  XNOR U16480 ( .A(n18004), .B(n18005), .Z(n18000) );
  XNOR U16481 ( .A(n16430), .B(n16442), .Z(n17996) );
  AND U16482 ( .A(n18008), .B(n18009), .Z(n16442) );
  AND U16483 ( .A(n18010), .B(n18011), .Z(n16430) );
  XNOR U16484 ( .A(n17490), .B(n119), .Z(n17492) );
  XOR U16485 ( .A(n17487), .B(n17488), .Z(n119) );
  AND U16486 ( .A(n18012), .B(n18013), .Z(n17488) );
  XOR U16487 ( .A(n17484), .B(n17485), .Z(n17487) );
  AND U16488 ( .A(n18014), .B(n18015), .Z(n17485) );
  XOR U16489 ( .A(n17481), .B(n17482), .Z(n17484) );
  AND U16490 ( .A(n18016), .B(n18017), .Z(n17482) );
  XOR U16491 ( .A(n17478), .B(n17479), .Z(n17481) );
  AND U16492 ( .A(n18018), .B(n18019), .Z(n17479) );
  XOR U16493 ( .A(n17475), .B(n17476), .Z(n17478) );
  AND U16494 ( .A(n18020), .B(n18021), .Z(n17476) );
  XOR U16495 ( .A(n17472), .B(n17473), .Z(n17475) );
  AND U16496 ( .A(n18022), .B(n18023), .Z(n17473) );
  XOR U16497 ( .A(n17469), .B(n17470), .Z(n17472) );
  AND U16498 ( .A(n18024), .B(n18025), .Z(n17470) );
  XOR U16499 ( .A(n17466), .B(n17467), .Z(n17469) );
  AND U16500 ( .A(n18026), .B(n18027), .Z(n17467) );
  XOR U16501 ( .A(n17463), .B(n17464), .Z(n17466) );
  AND U16502 ( .A(n18028), .B(n18029), .Z(n17464) );
  XOR U16503 ( .A(n17460), .B(n17461), .Z(n17463) );
  AND U16504 ( .A(n18030), .B(n18031), .Z(n17461) );
  XOR U16505 ( .A(n17457), .B(n17458), .Z(n17460) );
  AND U16506 ( .A(n18032), .B(n18033), .Z(n17458) );
  XOR U16507 ( .A(n17454), .B(n17455), .Z(n17457) );
  AND U16508 ( .A(n18034), .B(n18035), .Z(n17455) );
  XOR U16509 ( .A(n17451), .B(n17452), .Z(n17454) );
  AND U16510 ( .A(n18036), .B(n18037), .Z(n17452) );
  XOR U16511 ( .A(n17448), .B(n17449), .Z(n17451) );
  AND U16512 ( .A(n18038), .B(n18039), .Z(n17449) );
  XOR U16513 ( .A(n17445), .B(n17446), .Z(n17448) );
  AND U16514 ( .A(n18040), .B(n18041), .Z(n17446) );
  XOR U16515 ( .A(n17442), .B(n17443), .Z(n17445) );
  AND U16516 ( .A(n18042), .B(n18043), .Z(n17443) );
  XOR U16517 ( .A(n17439), .B(n17440), .Z(n17442) );
  AND U16518 ( .A(n18044), .B(n18045), .Z(n17440) );
  XOR U16519 ( .A(n17436), .B(n17437), .Z(n17439) );
  AND U16520 ( .A(n18046), .B(n18047), .Z(n17437) );
  XOR U16521 ( .A(n17433), .B(n17434), .Z(n17436) );
  AND U16522 ( .A(n18048), .B(n18049), .Z(n17434) );
  XOR U16523 ( .A(n17430), .B(n17431), .Z(n17433) );
  AND U16524 ( .A(n18050), .B(n18051), .Z(n17431) );
  XOR U16525 ( .A(n17427), .B(n17428), .Z(n17430) );
  AND U16526 ( .A(n18052), .B(n18053), .Z(n17428) );
  XOR U16527 ( .A(n17424), .B(n17425), .Z(n17427) );
  AND U16528 ( .A(n18054), .B(n18055), .Z(n17425) );
  XOR U16529 ( .A(n17421), .B(n17422), .Z(n17424) );
  AND U16530 ( .A(n18056), .B(n18057), .Z(n17422) );
  XOR U16531 ( .A(n17418), .B(n17419), .Z(n17421) );
  AND U16532 ( .A(n18058), .B(n18059), .Z(n17419) );
  XOR U16533 ( .A(n17415), .B(n17416), .Z(n17418) );
  AND U16534 ( .A(n18060), .B(n18061), .Z(n17416) );
  XOR U16535 ( .A(n17412), .B(n17413), .Z(n17415) );
  AND U16536 ( .A(n18062), .B(n18063), .Z(n17413) );
  XOR U16537 ( .A(n17409), .B(n17410), .Z(n17412) );
  AND U16538 ( .A(n18064), .B(n18065), .Z(n17410) );
  XOR U16539 ( .A(n17406), .B(n17407), .Z(n17409) );
  AND U16540 ( .A(n18066), .B(n18067), .Z(n17407) );
  XOR U16541 ( .A(n17403), .B(n17404), .Z(n17406) );
  AND U16542 ( .A(n18068), .B(n18069), .Z(n17404) );
  XOR U16543 ( .A(n17400), .B(n17401), .Z(n17403) );
  AND U16544 ( .A(n18070), .B(n18071), .Z(n17401) );
  XOR U16545 ( .A(n17397), .B(n17398), .Z(n17400) );
  AND U16546 ( .A(n18072), .B(n18073), .Z(n17398) );
  XOR U16547 ( .A(n17394), .B(n17395), .Z(n17397) );
  AND U16548 ( .A(n18074), .B(n18075), .Z(n17395) );
  XOR U16549 ( .A(n17391), .B(n17392), .Z(n17394) );
  AND U16550 ( .A(n18076), .B(n18077), .Z(n17392) );
  XOR U16551 ( .A(n17388), .B(n17389), .Z(n17391) );
  AND U16552 ( .A(n18078), .B(n18079), .Z(n17389) );
  XOR U16553 ( .A(n17385), .B(n17386), .Z(n17388) );
  AND U16554 ( .A(n18080), .B(n18081), .Z(n17386) );
  XOR U16555 ( .A(n17382), .B(n17383), .Z(n17385) );
  AND U16556 ( .A(n18082), .B(n18083), .Z(n17383) );
  XOR U16557 ( .A(n17379), .B(n17380), .Z(n17382) );
  AND U16558 ( .A(n18084), .B(n18085), .Z(n17380) );
  XOR U16559 ( .A(n17376), .B(n17377), .Z(n17379) );
  AND U16560 ( .A(n18086), .B(n18087), .Z(n17377) );
  XOR U16561 ( .A(n17373), .B(n17374), .Z(n17376) );
  AND U16562 ( .A(n18088), .B(n18089), .Z(n17374) );
  XOR U16563 ( .A(n17370), .B(n17371), .Z(n17373) );
  AND U16564 ( .A(n18090), .B(n18091), .Z(n17371) );
  XOR U16565 ( .A(n17367), .B(n17368), .Z(n17370) );
  AND U16566 ( .A(n18092), .B(n18093), .Z(n17368) );
  XOR U16567 ( .A(n17364), .B(n17365), .Z(n17367) );
  AND U16568 ( .A(n18094), .B(n18095), .Z(n17365) );
  XOR U16569 ( .A(n17361), .B(n17362), .Z(n17364) );
  AND U16570 ( .A(n18096), .B(n18097), .Z(n17362) );
  XOR U16571 ( .A(n17358), .B(n17359), .Z(n17361) );
  AND U16572 ( .A(n18098), .B(n18099), .Z(n17359) );
  XOR U16573 ( .A(n17355), .B(n17356), .Z(n17358) );
  AND U16574 ( .A(n18100), .B(n18101), .Z(n17356) );
  XOR U16575 ( .A(n17352), .B(n17353), .Z(n17355) );
  AND U16576 ( .A(n18102), .B(n18103), .Z(n17353) );
  XOR U16577 ( .A(n17349), .B(n17350), .Z(n17352) );
  AND U16578 ( .A(n18104), .B(n18105), .Z(n17350) );
  XOR U16579 ( .A(n17346), .B(n17347), .Z(n17349) );
  AND U16580 ( .A(n18106), .B(n18107), .Z(n17347) );
  XOR U16581 ( .A(n17343), .B(n17344), .Z(n17346) );
  AND U16582 ( .A(n18108), .B(n18109), .Z(n17344) );
  XOR U16583 ( .A(n17340), .B(n17341), .Z(n17343) );
  AND U16584 ( .A(n18110), .B(n18111), .Z(n17341) );
  XOR U16585 ( .A(n17337), .B(n17338), .Z(n17340) );
  AND U16586 ( .A(n18112), .B(n18113), .Z(n17338) );
  XOR U16587 ( .A(n17334), .B(n17335), .Z(n17337) );
  AND U16588 ( .A(n18114), .B(n18115), .Z(n17335) );
  XOR U16589 ( .A(n17331), .B(n17332), .Z(n17334) );
  AND U16590 ( .A(n18116), .B(n18117), .Z(n17332) );
  XOR U16591 ( .A(n17328), .B(n17329), .Z(n17331) );
  AND U16592 ( .A(n18118), .B(n18119), .Z(n17329) );
  XOR U16593 ( .A(n17325), .B(n17326), .Z(n17328) );
  AND U16594 ( .A(n18120), .B(n18121), .Z(n17326) );
  XOR U16595 ( .A(n17322), .B(n17323), .Z(n17325) );
  AND U16596 ( .A(n18122), .B(n18123), .Z(n17323) );
  XOR U16597 ( .A(n17319), .B(n17320), .Z(n17322) );
  AND U16598 ( .A(n18124), .B(n18125), .Z(n17320) );
  XOR U16599 ( .A(n17316), .B(n17317), .Z(n17319) );
  AND U16600 ( .A(n18126), .B(n18127), .Z(n17317) );
  XOR U16601 ( .A(n17313), .B(n17314), .Z(n17316) );
  AND U16602 ( .A(n18128), .B(n18129), .Z(n17314) );
  XOR U16603 ( .A(n17310), .B(n17311), .Z(n17313) );
  AND U16604 ( .A(n18130), .B(n18131), .Z(n17311) );
  XOR U16605 ( .A(n17307), .B(n17308), .Z(n17310) );
  AND U16606 ( .A(n18132), .B(n18133), .Z(n17308) );
  XOR U16607 ( .A(n17304), .B(n17305), .Z(n17307) );
  AND U16608 ( .A(n18134), .B(n18135), .Z(n17305) );
  XOR U16609 ( .A(n17301), .B(n17302), .Z(n17304) );
  AND U16610 ( .A(n18136), .B(n18137), .Z(n17302) );
  XOR U16611 ( .A(n17298), .B(n17299), .Z(n17301) );
  AND U16612 ( .A(n18138), .B(n18139), .Z(n17299) );
  XOR U16613 ( .A(n17295), .B(n17296), .Z(n17298) );
  AND U16614 ( .A(n18140), .B(n18141), .Z(n17296) );
  XOR U16615 ( .A(n17292), .B(n17293), .Z(n17295) );
  AND U16616 ( .A(n18142), .B(n18143), .Z(n17293) );
  XOR U16617 ( .A(n17289), .B(n17290), .Z(n17292) );
  AND U16618 ( .A(n18144), .B(n18145), .Z(n17290) );
  XOR U16619 ( .A(n17286), .B(n17287), .Z(n17289) );
  AND U16620 ( .A(n18146), .B(n18147), .Z(n17287) );
  XOR U16621 ( .A(n17283), .B(n17284), .Z(n17286) );
  AND U16622 ( .A(n18148), .B(n18149), .Z(n17284) );
  XOR U16623 ( .A(n17280), .B(n17281), .Z(n17283) );
  AND U16624 ( .A(n18150), .B(n18151), .Z(n17281) );
  XOR U16625 ( .A(n17277), .B(n17278), .Z(n17280) );
  AND U16626 ( .A(n18152), .B(n18153), .Z(n17278) );
  XOR U16627 ( .A(n17274), .B(n17275), .Z(n17277) );
  AND U16628 ( .A(n18154), .B(n18155), .Z(n17275) );
  XOR U16629 ( .A(n17271), .B(n17272), .Z(n17274) );
  AND U16630 ( .A(n18156), .B(n18157), .Z(n17272) );
  XOR U16631 ( .A(n17268), .B(n17269), .Z(n17271) );
  AND U16632 ( .A(n18158), .B(n18159), .Z(n17269) );
  XOR U16633 ( .A(n17265), .B(n17266), .Z(n17268) );
  AND U16634 ( .A(n18160), .B(n18161), .Z(n17266) );
  XOR U16635 ( .A(n17262), .B(n17263), .Z(n17265) );
  AND U16636 ( .A(n18162), .B(n18163), .Z(n17263) );
  XOR U16637 ( .A(n17259), .B(n17260), .Z(n17262) );
  AND U16638 ( .A(n18164), .B(n18165), .Z(n17260) );
  XOR U16639 ( .A(n17256), .B(n17257), .Z(n17259) );
  AND U16640 ( .A(n18166), .B(n18167), .Z(n17257) );
  XOR U16641 ( .A(n17253), .B(n17254), .Z(n17256) );
  AND U16642 ( .A(n18168), .B(n18169), .Z(n17254) );
  XOR U16643 ( .A(n17250), .B(n17251), .Z(n17253) );
  AND U16644 ( .A(n18170), .B(n18171), .Z(n17251) );
  XOR U16645 ( .A(n17247), .B(n17248), .Z(n17250) );
  AND U16646 ( .A(n18172), .B(n18173), .Z(n17248) );
  XOR U16647 ( .A(n17244), .B(n17245), .Z(n17247) );
  AND U16648 ( .A(n18174), .B(n18175), .Z(n17245) );
  XOR U16649 ( .A(n17241), .B(n17242), .Z(n17244) );
  AND U16650 ( .A(n18176), .B(n18177), .Z(n17242) );
  XOR U16651 ( .A(n17238), .B(n17239), .Z(n17241) );
  AND U16652 ( .A(n18178), .B(n18179), .Z(n17239) );
  XOR U16653 ( .A(n17235), .B(n17236), .Z(n17238) );
  AND U16654 ( .A(n18180), .B(n18181), .Z(n17236) );
  XOR U16655 ( .A(n17232), .B(n17233), .Z(n17235) );
  AND U16656 ( .A(n18182), .B(n18183), .Z(n17233) );
  XOR U16657 ( .A(n17229), .B(n17230), .Z(n17232) );
  AND U16658 ( .A(n18184), .B(n18185), .Z(n17230) );
  XOR U16659 ( .A(n17226), .B(n17227), .Z(n17229) );
  AND U16660 ( .A(n18186), .B(n18187), .Z(n17227) );
  XOR U16661 ( .A(n17223), .B(n17224), .Z(n17226) );
  AND U16662 ( .A(n18188), .B(n18189), .Z(n17224) );
  XOR U16663 ( .A(n17220), .B(n17221), .Z(n17223) );
  AND U16664 ( .A(n18190), .B(n18191), .Z(n17221) );
  XOR U16665 ( .A(n17217), .B(n17218), .Z(n17220) );
  AND U16666 ( .A(n18192), .B(n18193), .Z(n17218) );
  XOR U16667 ( .A(n17214), .B(n17215), .Z(n17217) );
  AND U16668 ( .A(n18194), .B(n18195), .Z(n17215) );
  XOR U16669 ( .A(n17211), .B(n17212), .Z(n17214) );
  AND U16670 ( .A(n18196), .B(n18197), .Z(n17212) );
  XOR U16671 ( .A(n17208), .B(n17209), .Z(n17211) );
  AND U16672 ( .A(n18198), .B(n18199), .Z(n17209) );
  XOR U16673 ( .A(n17205), .B(n17206), .Z(n17208) );
  AND U16674 ( .A(n18200), .B(n18201), .Z(n17206) );
  XOR U16675 ( .A(n17202), .B(n17203), .Z(n17205) );
  AND U16676 ( .A(n18202), .B(n18203), .Z(n17203) );
  XOR U16677 ( .A(n17199), .B(n17200), .Z(n17202) );
  AND U16678 ( .A(n18204), .B(n18205), .Z(n17200) );
  XOR U16679 ( .A(n17196), .B(n17197), .Z(n17199) );
  AND U16680 ( .A(n18206), .B(n18207), .Z(n17197) );
  XOR U16681 ( .A(n17193), .B(n17194), .Z(n17196) );
  AND U16682 ( .A(n18208), .B(n18209), .Z(n17194) );
  XOR U16683 ( .A(n17190), .B(n17191), .Z(n17193) );
  AND U16684 ( .A(n18210), .B(n18211), .Z(n17191) );
  XOR U16685 ( .A(n17187), .B(n17188), .Z(n17190) );
  AND U16686 ( .A(n18212), .B(n18213), .Z(n17188) );
  XOR U16687 ( .A(n17184), .B(n17185), .Z(n17187) );
  AND U16688 ( .A(n18214), .B(n18215), .Z(n17185) );
  XOR U16689 ( .A(n17181), .B(n17182), .Z(n17184) );
  AND U16690 ( .A(n18216), .B(n18217), .Z(n17182) );
  XOR U16691 ( .A(n17178), .B(n17179), .Z(n17181) );
  AND U16692 ( .A(n18218), .B(n18219), .Z(n17179) );
  XOR U16693 ( .A(n17175), .B(n17176), .Z(n17178) );
  AND U16694 ( .A(n18220), .B(n18221), .Z(n17176) );
  XOR U16695 ( .A(n17172), .B(n17173), .Z(n17175) );
  AND U16696 ( .A(n18222), .B(n18223), .Z(n17173) );
  XOR U16697 ( .A(n17169), .B(n17170), .Z(n17172) );
  AND U16698 ( .A(n18224), .B(n18225), .Z(n17170) );
  XOR U16699 ( .A(n17166), .B(n17167), .Z(n17169) );
  AND U16700 ( .A(n18226), .B(n18227), .Z(n17167) );
  XOR U16701 ( .A(n17163), .B(n17164), .Z(n17166) );
  AND U16702 ( .A(n18228), .B(n18229), .Z(n17164) );
  XOR U16703 ( .A(n17160), .B(n17161), .Z(n17163) );
  AND U16704 ( .A(n18230), .B(n18231), .Z(n17161) );
  XOR U16705 ( .A(n17157), .B(n17158), .Z(n17160) );
  AND U16706 ( .A(n18232), .B(n18233), .Z(n17158) );
  XOR U16707 ( .A(n17154), .B(n17155), .Z(n17157) );
  AND U16708 ( .A(n18234), .B(n18235), .Z(n17155) );
  XOR U16709 ( .A(n17151), .B(n17152), .Z(n17154) );
  AND U16710 ( .A(n18236), .B(n18237), .Z(n17152) );
  XOR U16711 ( .A(n17148), .B(n17149), .Z(n17151) );
  AND U16712 ( .A(n18238), .B(n18239), .Z(n17149) );
  XOR U16713 ( .A(n17145), .B(n17146), .Z(n17148) );
  AND U16714 ( .A(n18240), .B(n18241), .Z(n17146) );
  XOR U16715 ( .A(n17142), .B(n17143), .Z(n17145) );
  AND U16716 ( .A(n18242), .B(n18243), .Z(n17143) );
  XOR U16717 ( .A(n17139), .B(n17140), .Z(n17142) );
  AND U16718 ( .A(n18244), .B(n18245), .Z(n17140) );
  XOR U16719 ( .A(n17136), .B(n17137), .Z(n17139) );
  AND U16720 ( .A(n18246), .B(n18247), .Z(n17137) );
  XOR U16721 ( .A(n17133), .B(n17134), .Z(n17136) );
  AND U16722 ( .A(n18248), .B(n18249), .Z(n17134) );
  XOR U16723 ( .A(n17130), .B(n17131), .Z(n17133) );
  AND U16724 ( .A(n18250), .B(n18251), .Z(n17131) );
  XOR U16725 ( .A(n17127), .B(n17128), .Z(n17130) );
  AND U16726 ( .A(n18252), .B(n18253), .Z(n17128) );
  XOR U16727 ( .A(n17124), .B(n17125), .Z(n17127) );
  AND U16728 ( .A(n18254), .B(n18255), .Z(n17125) );
  XOR U16729 ( .A(n17121), .B(n17122), .Z(n17124) );
  AND U16730 ( .A(n18256), .B(n18257), .Z(n17122) );
  XOR U16731 ( .A(n17118), .B(n17119), .Z(n17121) );
  AND U16732 ( .A(n18258), .B(n18259), .Z(n17119) );
  XOR U16733 ( .A(n17115), .B(n17116), .Z(n17118) );
  AND U16734 ( .A(n18260), .B(n18261), .Z(n17116) );
  XOR U16735 ( .A(n17112), .B(n17113), .Z(n17115) );
  AND U16736 ( .A(n18262), .B(n18263), .Z(n17113) );
  XOR U16737 ( .A(n17109), .B(n17110), .Z(n17112) );
  AND U16738 ( .A(n18264), .B(n18265), .Z(n17110) );
  XOR U16739 ( .A(n17106), .B(n17107), .Z(n17109) );
  AND U16740 ( .A(n18266), .B(n18267), .Z(n17107) );
  XNOR U16741 ( .A(n17103), .B(n17104), .Z(n17106) );
  AND U16742 ( .A(n18268), .B(n18269), .Z(n17104) );
  XOR U16743 ( .A(n18270), .B(n17101), .Z(n17103) );
  IV U16744 ( .A(n18271), .Z(n17101) );
  AND U16745 ( .A(n18272), .B(n18273), .Z(n18271) );
  IV U16746 ( .A(n17100), .Z(n18270) );
  XOR U16747 ( .A(n16841), .B(n17097), .Z(n17100) );
  AND U16748 ( .A(n18274), .B(n18275), .Z(n17097) );
  XOR U16749 ( .A(n16843), .B(n16842), .Z(n16841) );
  AND U16750 ( .A(n18276), .B(n18277), .Z(n16842) );
  XOR U16751 ( .A(n16845), .B(n16844), .Z(n16843) );
  AND U16752 ( .A(n18278), .B(n18279), .Z(n16844) );
  XOR U16753 ( .A(n16847), .B(n16846), .Z(n16845) );
  AND U16754 ( .A(n18280), .B(n18281), .Z(n16846) );
  XOR U16755 ( .A(n16849), .B(n16848), .Z(n16847) );
  AND U16756 ( .A(n18282), .B(n18283), .Z(n16848) );
  XOR U16757 ( .A(n16851), .B(n16850), .Z(n16849) );
  AND U16758 ( .A(n18284), .B(n18285), .Z(n16850) );
  XOR U16759 ( .A(n16853), .B(n16852), .Z(n16851) );
  AND U16760 ( .A(n18286), .B(n18287), .Z(n16852) );
  XOR U16761 ( .A(n16855), .B(n16854), .Z(n16853) );
  AND U16762 ( .A(n18288), .B(n18289), .Z(n16854) );
  XOR U16763 ( .A(n16857), .B(n16856), .Z(n16855) );
  AND U16764 ( .A(n18290), .B(n18291), .Z(n16856) );
  XOR U16765 ( .A(n16859), .B(n16858), .Z(n16857) );
  AND U16766 ( .A(n18292), .B(n18293), .Z(n16858) );
  XOR U16767 ( .A(n16861), .B(n16860), .Z(n16859) );
  AND U16768 ( .A(n18294), .B(n18295), .Z(n16860) );
  XOR U16769 ( .A(n16863), .B(n16862), .Z(n16861) );
  AND U16770 ( .A(n18296), .B(n18297), .Z(n16862) );
  XOR U16771 ( .A(n16865), .B(n16864), .Z(n16863) );
  AND U16772 ( .A(n18298), .B(n18299), .Z(n16864) );
  XOR U16773 ( .A(n16867), .B(n16866), .Z(n16865) );
  AND U16774 ( .A(n18300), .B(n18301), .Z(n16866) );
  XOR U16775 ( .A(n16869), .B(n16868), .Z(n16867) );
  AND U16776 ( .A(n18302), .B(n18303), .Z(n16868) );
  XOR U16777 ( .A(n16871), .B(n16870), .Z(n16869) );
  AND U16778 ( .A(n18304), .B(n18305), .Z(n16870) );
  XOR U16779 ( .A(n16873), .B(n16872), .Z(n16871) );
  AND U16780 ( .A(n18306), .B(n18307), .Z(n16872) );
  XOR U16781 ( .A(n16875), .B(n16874), .Z(n16873) );
  AND U16782 ( .A(n18308), .B(n18309), .Z(n16874) );
  XOR U16783 ( .A(n16877), .B(n16876), .Z(n16875) );
  AND U16784 ( .A(n18310), .B(n18311), .Z(n16876) );
  XOR U16785 ( .A(n16879), .B(n16878), .Z(n16877) );
  AND U16786 ( .A(n18312), .B(n18313), .Z(n16878) );
  XOR U16787 ( .A(n16881), .B(n16880), .Z(n16879) );
  AND U16788 ( .A(n18314), .B(n18315), .Z(n16880) );
  XOR U16789 ( .A(n16883), .B(n16882), .Z(n16881) );
  AND U16790 ( .A(n18316), .B(n18317), .Z(n16882) );
  XOR U16791 ( .A(n16885), .B(n16884), .Z(n16883) );
  AND U16792 ( .A(n18318), .B(n18319), .Z(n16884) );
  XOR U16793 ( .A(n16887), .B(n16886), .Z(n16885) );
  AND U16794 ( .A(n18320), .B(n18321), .Z(n16886) );
  XOR U16795 ( .A(n16889), .B(n16888), .Z(n16887) );
  AND U16796 ( .A(n18322), .B(n18323), .Z(n16888) );
  XOR U16797 ( .A(n16891), .B(n16890), .Z(n16889) );
  AND U16798 ( .A(n18324), .B(n18325), .Z(n16890) );
  XOR U16799 ( .A(n16893), .B(n16892), .Z(n16891) );
  AND U16800 ( .A(n18326), .B(n18327), .Z(n16892) );
  XOR U16801 ( .A(n16895), .B(n16894), .Z(n16893) );
  AND U16802 ( .A(n18328), .B(n18329), .Z(n16894) );
  XOR U16803 ( .A(n16897), .B(n16896), .Z(n16895) );
  AND U16804 ( .A(n18330), .B(n18331), .Z(n16896) );
  XOR U16805 ( .A(n16899), .B(n16898), .Z(n16897) );
  AND U16806 ( .A(n18332), .B(n18333), .Z(n16898) );
  XOR U16807 ( .A(n16901), .B(n16900), .Z(n16899) );
  AND U16808 ( .A(n18334), .B(n18335), .Z(n16900) );
  XOR U16809 ( .A(n16903), .B(n16902), .Z(n16901) );
  AND U16810 ( .A(n18336), .B(n18337), .Z(n16902) );
  XOR U16811 ( .A(n16905), .B(n16904), .Z(n16903) );
  AND U16812 ( .A(n18338), .B(n18339), .Z(n16904) );
  XOR U16813 ( .A(n16907), .B(n16906), .Z(n16905) );
  AND U16814 ( .A(n18340), .B(n18341), .Z(n16906) );
  XOR U16815 ( .A(n16909), .B(n16908), .Z(n16907) );
  AND U16816 ( .A(n18342), .B(n18343), .Z(n16908) );
  XOR U16817 ( .A(n16911), .B(n16910), .Z(n16909) );
  AND U16818 ( .A(n18344), .B(n18345), .Z(n16910) );
  XOR U16819 ( .A(n16913), .B(n16912), .Z(n16911) );
  AND U16820 ( .A(n18346), .B(n18347), .Z(n16912) );
  XOR U16821 ( .A(n16915), .B(n16914), .Z(n16913) );
  AND U16822 ( .A(n18348), .B(n18349), .Z(n16914) );
  XOR U16823 ( .A(n16917), .B(n16916), .Z(n16915) );
  AND U16824 ( .A(n18350), .B(n18351), .Z(n16916) );
  XOR U16825 ( .A(n16919), .B(n16918), .Z(n16917) );
  AND U16826 ( .A(n18352), .B(n18353), .Z(n16918) );
  XOR U16827 ( .A(n16921), .B(n16920), .Z(n16919) );
  AND U16828 ( .A(n18354), .B(n18355), .Z(n16920) );
  XOR U16829 ( .A(n16923), .B(n16922), .Z(n16921) );
  AND U16830 ( .A(n18356), .B(n18357), .Z(n16922) );
  XOR U16831 ( .A(n16925), .B(n16924), .Z(n16923) );
  AND U16832 ( .A(n18358), .B(n18359), .Z(n16924) );
  XOR U16833 ( .A(n16927), .B(n16926), .Z(n16925) );
  AND U16834 ( .A(n18360), .B(n18361), .Z(n16926) );
  XOR U16835 ( .A(n16929), .B(n16928), .Z(n16927) );
  AND U16836 ( .A(n18362), .B(n18363), .Z(n16928) );
  XOR U16837 ( .A(n16931), .B(n16930), .Z(n16929) );
  AND U16838 ( .A(n18364), .B(n18365), .Z(n16930) );
  XOR U16839 ( .A(n16933), .B(n16932), .Z(n16931) );
  AND U16840 ( .A(n18366), .B(n18367), .Z(n16932) );
  XOR U16841 ( .A(n16935), .B(n16934), .Z(n16933) );
  AND U16842 ( .A(n18368), .B(n18369), .Z(n16934) );
  XOR U16843 ( .A(n16937), .B(n16936), .Z(n16935) );
  AND U16844 ( .A(n18370), .B(n18371), .Z(n16936) );
  XOR U16845 ( .A(n16939), .B(n16938), .Z(n16937) );
  AND U16846 ( .A(n18372), .B(n18373), .Z(n16938) );
  XOR U16847 ( .A(n16941), .B(n16940), .Z(n16939) );
  AND U16848 ( .A(n18374), .B(n18375), .Z(n16940) );
  XOR U16849 ( .A(n16943), .B(n16942), .Z(n16941) );
  AND U16850 ( .A(n18376), .B(n18377), .Z(n16942) );
  XOR U16851 ( .A(n16945), .B(n16944), .Z(n16943) );
  AND U16852 ( .A(n18378), .B(n18379), .Z(n16944) );
  XOR U16853 ( .A(n16947), .B(n16946), .Z(n16945) );
  AND U16854 ( .A(n18380), .B(n18381), .Z(n16946) );
  XOR U16855 ( .A(n16949), .B(n16948), .Z(n16947) );
  AND U16856 ( .A(n18382), .B(n18383), .Z(n16948) );
  XOR U16857 ( .A(n16951), .B(n16950), .Z(n16949) );
  AND U16858 ( .A(n18384), .B(n18385), .Z(n16950) );
  XOR U16859 ( .A(n16953), .B(n16952), .Z(n16951) );
  AND U16860 ( .A(n18386), .B(n18387), .Z(n16952) );
  XOR U16861 ( .A(n16955), .B(n16954), .Z(n16953) );
  AND U16862 ( .A(n18388), .B(n18389), .Z(n16954) );
  XOR U16863 ( .A(n16957), .B(n16956), .Z(n16955) );
  AND U16864 ( .A(n18390), .B(n18391), .Z(n16956) );
  XOR U16865 ( .A(n16959), .B(n16958), .Z(n16957) );
  AND U16866 ( .A(n18392), .B(n18393), .Z(n16958) );
  XOR U16867 ( .A(n16961), .B(n16960), .Z(n16959) );
  AND U16868 ( .A(n18394), .B(n18395), .Z(n16960) );
  XOR U16869 ( .A(n16963), .B(n16962), .Z(n16961) );
  AND U16870 ( .A(n18396), .B(n18397), .Z(n16962) );
  XOR U16871 ( .A(n16965), .B(n16964), .Z(n16963) );
  AND U16872 ( .A(n18398), .B(n18399), .Z(n16964) );
  XOR U16873 ( .A(n16967), .B(n16966), .Z(n16965) );
  AND U16874 ( .A(n18400), .B(n18401), .Z(n16966) );
  XOR U16875 ( .A(n16969), .B(n16968), .Z(n16967) );
  AND U16876 ( .A(n18402), .B(n18403), .Z(n16968) );
  XOR U16877 ( .A(n16971), .B(n16970), .Z(n16969) );
  AND U16878 ( .A(n18404), .B(n18405), .Z(n16970) );
  XOR U16879 ( .A(n16973), .B(n16972), .Z(n16971) );
  AND U16880 ( .A(n18406), .B(n18407), .Z(n16972) );
  XOR U16881 ( .A(n16975), .B(n16974), .Z(n16973) );
  AND U16882 ( .A(n18408), .B(n18409), .Z(n16974) );
  XOR U16883 ( .A(n16977), .B(n16976), .Z(n16975) );
  AND U16884 ( .A(n18410), .B(n18411), .Z(n16976) );
  XOR U16885 ( .A(n16979), .B(n16978), .Z(n16977) );
  AND U16886 ( .A(n18412), .B(n18413), .Z(n16978) );
  XOR U16887 ( .A(n16981), .B(n16980), .Z(n16979) );
  AND U16888 ( .A(n18414), .B(n18415), .Z(n16980) );
  XOR U16889 ( .A(n16983), .B(n16982), .Z(n16981) );
  AND U16890 ( .A(n18416), .B(n18417), .Z(n16982) );
  XOR U16891 ( .A(n16985), .B(n16984), .Z(n16983) );
  AND U16892 ( .A(n18418), .B(n18419), .Z(n16984) );
  XOR U16893 ( .A(n16987), .B(n16986), .Z(n16985) );
  AND U16894 ( .A(n18420), .B(n18421), .Z(n16986) );
  XOR U16895 ( .A(n16989), .B(n16988), .Z(n16987) );
  AND U16896 ( .A(n18422), .B(n18423), .Z(n16988) );
  XOR U16897 ( .A(n16991), .B(n16990), .Z(n16989) );
  AND U16898 ( .A(n18424), .B(n18425), .Z(n16990) );
  XOR U16899 ( .A(n16993), .B(n16992), .Z(n16991) );
  AND U16900 ( .A(n18426), .B(n18427), .Z(n16992) );
  XOR U16901 ( .A(n16995), .B(n16994), .Z(n16993) );
  AND U16902 ( .A(n18428), .B(n18429), .Z(n16994) );
  XOR U16903 ( .A(n16997), .B(n16996), .Z(n16995) );
  AND U16904 ( .A(n18430), .B(n18431), .Z(n16996) );
  XOR U16905 ( .A(n16999), .B(n16998), .Z(n16997) );
  AND U16906 ( .A(n18432), .B(n18433), .Z(n16998) );
  XOR U16907 ( .A(n17001), .B(n17000), .Z(n16999) );
  AND U16908 ( .A(n18434), .B(n18435), .Z(n17000) );
  XOR U16909 ( .A(n17003), .B(n17002), .Z(n17001) );
  AND U16910 ( .A(n18436), .B(n18437), .Z(n17002) );
  XOR U16911 ( .A(n17005), .B(n17004), .Z(n17003) );
  AND U16912 ( .A(n18438), .B(n18439), .Z(n17004) );
  XOR U16913 ( .A(n17007), .B(n17006), .Z(n17005) );
  AND U16914 ( .A(n18440), .B(n18441), .Z(n17006) );
  XOR U16915 ( .A(n17009), .B(n17008), .Z(n17007) );
  AND U16916 ( .A(n18442), .B(n18443), .Z(n17008) );
  XOR U16917 ( .A(n17011), .B(n17010), .Z(n17009) );
  AND U16918 ( .A(n18444), .B(n18445), .Z(n17010) );
  XOR U16919 ( .A(n17013), .B(n17012), .Z(n17011) );
  AND U16920 ( .A(n18446), .B(n18447), .Z(n17012) );
  XOR U16921 ( .A(n17015), .B(n17014), .Z(n17013) );
  AND U16922 ( .A(n18448), .B(n18449), .Z(n17014) );
  XOR U16923 ( .A(n17017), .B(n17016), .Z(n17015) );
  AND U16924 ( .A(n18450), .B(n18451), .Z(n17016) );
  XOR U16925 ( .A(n17019), .B(n17018), .Z(n17017) );
  AND U16926 ( .A(n18452), .B(n18453), .Z(n17018) );
  XOR U16927 ( .A(n17021), .B(n17020), .Z(n17019) );
  AND U16928 ( .A(n18454), .B(n18455), .Z(n17020) );
  XOR U16929 ( .A(n17023), .B(n17022), .Z(n17021) );
  AND U16930 ( .A(n18456), .B(n18457), .Z(n17022) );
  XOR U16931 ( .A(n17025), .B(n17024), .Z(n17023) );
  AND U16932 ( .A(n18458), .B(n18459), .Z(n17024) );
  XOR U16933 ( .A(n17027), .B(n17026), .Z(n17025) );
  AND U16934 ( .A(n18460), .B(n18461), .Z(n17026) );
  XOR U16935 ( .A(n17029), .B(n17028), .Z(n17027) );
  AND U16936 ( .A(n18462), .B(n18463), .Z(n17028) );
  XOR U16937 ( .A(n17031), .B(n17030), .Z(n17029) );
  AND U16938 ( .A(n18464), .B(n18465), .Z(n17030) );
  XOR U16939 ( .A(n17033), .B(n17032), .Z(n17031) );
  AND U16940 ( .A(n18466), .B(n18467), .Z(n17032) );
  XOR U16941 ( .A(n17035), .B(n17034), .Z(n17033) );
  AND U16942 ( .A(n18468), .B(n18469), .Z(n17034) );
  XOR U16943 ( .A(n17037), .B(n17036), .Z(n17035) );
  AND U16944 ( .A(n18470), .B(n18471), .Z(n17036) );
  XOR U16945 ( .A(n17039), .B(n17038), .Z(n17037) );
  AND U16946 ( .A(n18472), .B(n18473), .Z(n17038) );
  XOR U16947 ( .A(n17041), .B(n17040), .Z(n17039) );
  AND U16948 ( .A(n18474), .B(n18475), .Z(n17040) );
  XOR U16949 ( .A(n17043), .B(n17042), .Z(n17041) );
  AND U16950 ( .A(n18476), .B(n18477), .Z(n17042) );
  XOR U16951 ( .A(n17045), .B(n17044), .Z(n17043) );
  AND U16952 ( .A(n18478), .B(n18479), .Z(n17044) );
  XOR U16953 ( .A(n17047), .B(n17046), .Z(n17045) );
  AND U16954 ( .A(n18480), .B(n18481), .Z(n17046) );
  XOR U16955 ( .A(n17049), .B(n17048), .Z(n17047) );
  AND U16956 ( .A(n18482), .B(n18483), .Z(n17048) );
  XOR U16957 ( .A(n17051), .B(n17050), .Z(n17049) );
  AND U16958 ( .A(n18484), .B(n18485), .Z(n17050) );
  XOR U16959 ( .A(n17053), .B(n17052), .Z(n17051) );
  AND U16960 ( .A(n18486), .B(n18487), .Z(n17052) );
  XOR U16961 ( .A(n17055), .B(n17054), .Z(n17053) );
  AND U16962 ( .A(n18488), .B(n18489), .Z(n17054) );
  XOR U16963 ( .A(n17057), .B(n17056), .Z(n17055) );
  AND U16964 ( .A(n18490), .B(n18491), .Z(n17056) );
  XOR U16965 ( .A(n17059), .B(n17058), .Z(n17057) );
  AND U16966 ( .A(n18492), .B(n18493), .Z(n17058) );
  XOR U16967 ( .A(n17061), .B(n17060), .Z(n17059) );
  AND U16968 ( .A(n18494), .B(n18495), .Z(n17060) );
  XOR U16969 ( .A(n17063), .B(n17062), .Z(n17061) );
  AND U16970 ( .A(n18496), .B(n18497), .Z(n17062) );
  XOR U16971 ( .A(n17065), .B(n17064), .Z(n17063) );
  AND U16972 ( .A(n18498), .B(n18499), .Z(n17064) );
  XOR U16973 ( .A(n17093), .B(n17066), .Z(n17065) );
  AND U16974 ( .A(n18500), .B(n18501), .Z(n17066) );
  XOR U16975 ( .A(n17095), .B(n17094), .Z(n17093) );
  AND U16976 ( .A(n18502), .B(n18503), .Z(n17094) );
  XOR U16977 ( .A(n17074), .B(n17096), .Z(n17095) );
  AND U16978 ( .A(n18504), .B(n18505), .Z(n17096) );
  XOR U16979 ( .A(n17070), .B(n17075), .Z(n17074) );
  AND U16980 ( .A(n18506), .B(n18507), .Z(n17075) );
  XOR U16981 ( .A(n17072), .B(n17071), .Z(n17070) );
  AND U16982 ( .A(n18508), .B(n18509), .Z(n17071) );
  XNOR U16983 ( .A(n17082), .B(n17073), .Z(n17072) );
  AND U16984 ( .A(n18510), .B(n18511), .Z(n17073) );
  XOR U16985 ( .A(n17092), .B(n17081), .Z(n17082) );
  AND U16986 ( .A(n18512), .B(n18513), .Z(n17081) );
  XNOR U16987 ( .A(n18514), .B(n17087), .Z(n17092) );
  XOR U16988 ( .A(n17088), .B(n18515), .Z(n17087) );
  AND U16989 ( .A(n18516), .B(n18517), .Z(n18515) );
  XOR U16990 ( .A(n18518), .B(n18519), .Z(n17088) );
  NOR U16991 ( .A(n18520), .B(n18521), .Z(n18519) );
  AND U16992 ( .A(n18522), .B(n18523), .Z(n18521) );
  AND U16993 ( .A(n18524), .B(n18525), .Z(n18520) );
  XNOR U16994 ( .A(n18522), .B(n18523), .Z(n18518) );
  XNOR U16995 ( .A(n17079), .B(n17091), .Z(n18514) );
  AND U16996 ( .A(n18526), .B(n18527), .Z(n17091) );
  AND U16997 ( .A(n18528), .B(n18529), .Z(n17079) );
  NOR U16998 ( .A(n9586), .B(n9589), .Z(n17490) );
  XNOR U16999 ( .A(n17495), .B(n17494), .Z(n9589) );
  NOR U17000 ( .A(n9075), .B(p_input[511]), .Z(n17494) );
  XOR U17001 ( .A(n17497), .B(n17496), .Z(n17495) );
  NOR U17002 ( .A(n9077), .B(p_input[509]), .Z(n17496) );
  XOR U17003 ( .A(n17499), .B(n17498), .Z(n17497) );
  NOR U17004 ( .A(n9079), .B(p_input[507]), .Z(n17498) );
  XOR U17005 ( .A(n17501), .B(n17500), .Z(n17499) );
  NOR U17006 ( .A(n9081), .B(p_input[505]), .Z(n17500) );
  XOR U17007 ( .A(n17503), .B(n17502), .Z(n17501) );
  NOR U17008 ( .A(n9083), .B(p_input[503]), .Z(n17502) );
  XOR U17009 ( .A(n17505), .B(n17504), .Z(n17503) );
  NOR U17010 ( .A(n9085), .B(p_input[501]), .Z(n17504) );
  XOR U17011 ( .A(n17507), .B(n17506), .Z(n17505) );
  NOR U17012 ( .A(n9087), .B(p_input[499]), .Z(n17506) );
  XOR U17013 ( .A(n17509), .B(n17508), .Z(n17507) );
  NOR U17014 ( .A(n9089), .B(p_input[497]), .Z(n17508) );
  XOR U17015 ( .A(n17511), .B(n17510), .Z(n17509) );
  NOR U17016 ( .A(n9091), .B(p_input[495]), .Z(n17510) );
  XOR U17017 ( .A(n17513), .B(n17512), .Z(n17511) );
  NOR U17018 ( .A(n9093), .B(p_input[493]), .Z(n17512) );
  XOR U17019 ( .A(n17515), .B(n17514), .Z(n17513) );
  NOR U17020 ( .A(n9095), .B(p_input[491]), .Z(n17514) );
  XOR U17021 ( .A(n17517), .B(n17516), .Z(n17515) );
  NOR U17022 ( .A(n9097), .B(p_input[489]), .Z(n17516) );
  XOR U17023 ( .A(n17519), .B(n17518), .Z(n17517) );
  NOR U17024 ( .A(n9099), .B(p_input[487]), .Z(n17518) );
  XOR U17025 ( .A(n17521), .B(n17520), .Z(n17519) );
  NOR U17026 ( .A(n9101), .B(p_input[485]), .Z(n17520) );
  XOR U17027 ( .A(n17523), .B(n17522), .Z(n17521) );
  NOR U17028 ( .A(n9103), .B(p_input[483]), .Z(n17522) );
  XOR U17029 ( .A(n17525), .B(n17524), .Z(n17523) );
  NOR U17030 ( .A(n9105), .B(p_input[481]), .Z(n17524) );
  XOR U17031 ( .A(n17527), .B(n17526), .Z(n17525) );
  NOR U17032 ( .A(n9107), .B(p_input[479]), .Z(n17526) );
  XOR U17033 ( .A(n17529), .B(n17528), .Z(n17527) );
  NOR U17034 ( .A(n9109), .B(p_input[477]), .Z(n17528) );
  XOR U17035 ( .A(n17531), .B(n17530), .Z(n17529) );
  NOR U17036 ( .A(n9111), .B(p_input[475]), .Z(n17530) );
  XOR U17037 ( .A(n17533), .B(n17532), .Z(n17531) );
  NOR U17038 ( .A(n9113), .B(p_input[473]), .Z(n17532) );
  XOR U17039 ( .A(n17535), .B(n17534), .Z(n17533) );
  NOR U17040 ( .A(n9115), .B(p_input[471]), .Z(n17534) );
  XOR U17041 ( .A(n17537), .B(n17536), .Z(n17535) );
  NOR U17042 ( .A(n9117), .B(p_input[469]), .Z(n17536) );
  XOR U17043 ( .A(n17539), .B(n17538), .Z(n17537) );
  NOR U17044 ( .A(n9119), .B(p_input[467]), .Z(n17538) );
  XOR U17045 ( .A(n17541), .B(n17540), .Z(n17539) );
  NOR U17046 ( .A(n9121), .B(p_input[465]), .Z(n17540) );
  XOR U17047 ( .A(n17543), .B(n17542), .Z(n17541) );
  NOR U17048 ( .A(n9123), .B(p_input[463]), .Z(n17542) );
  XOR U17049 ( .A(n17545), .B(n17544), .Z(n17543) );
  NOR U17050 ( .A(n9125), .B(p_input[461]), .Z(n17544) );
  XOR U17051 ( .A(n17547), .B(n17546), .Z(n17545) );
  NOR U17052 ( .A(n9127), .B(p_input[459]), .Z(n17546) );
  XOR U17053 ( .A(n17549), .B(n17548), .Z(n17547) );
  NOR U17054 ( .A(n9129), .B(p_input[457]), .Z(n17548) );
  XOR U17055 ( .A(n17551), .B(n17550), .Z(n17549) );
  NOR U17056 ( .A(n9131), .B(p_input[455]), .Z(n17550) );
  XOR U17057 ( .A(n17553), .B(n17552), .Z(n17551) );
  NOR U17058 ( .A(n9133), .B(p_input[453]), .Z(n17552) );
  XOR U17059 ( .A(n17555), .B(n17554), .Z(n17553) );
  NOR U17060 ( .A(n9135), .B(p_input[451]), .Z(n17554) );
  XOR U17061 ( .A(n17557), .B(n17556), .Z(n17555) );
  NOR U17062 ( .A(n9137), .B(p_input[449]), .Z(n17556) );
  XOR U17063 ( .A(n17559), .B(n17558), .Z(n17557) );
  NOR U17064 ( .A(n9139), .B(p_input[447]), .Z(n17558) );
  XOR U17065 ( .A(n17561), .B(n17560), .Z(n17559) );
  NOR U17066 ( .A(n9141), .B(p_input[445]), .Z(n17560) );
  XOR U17067 ( .A(n17563), .B(n17562), .Z(n17561) );
  NOR U17068 ( .A(n9143), .B(p_input[443]), .Z(n17562) );
  XOR U17069 ( .A(n17565), .B(n17564), .Z(n17563) );
  NOR U17070 ( .A(n9145), .B(p_input[441]), .Z(n17564) );
  XOR U17071 ( .A(n17567), .B(n17566), .Z(n17565) );
  NOR U17072 ( .A(n9147), .B(p_input[439]), .Z(n17566) );
  XOR U17073 ( .A(n17569), .B(n17568), .Z(n17567) );
  NOR U17074 ( .A(n9149), .B(p_input[437]), .Z(n17568) );
  XOR U17075 ( .A(n17571), .B(n17570), .Z(n17569) );
  NOR U17076 ( .A(n9151), .B(p_input[435]), .Z(n17570) );
  XOR U17077 ( .A(n17573), .B(n17572), .Z(n17571) );
  NOR U17078 ( .A(n9153), .B(p_input[433]), .Z(n17572) );
  XOR U17079 ( .A(n17575), .B(n17574), .Z(n17573) );
  NOR U17080 ( .A(n9155), .B(p_input[431]), .Z(n17574) );
  XOR U17081 ( .A(n17577), .B(n17576), .Z(n17575) );
  NOR U17082 ( .A(n9157), .B(p_input[429]), .Z(n17576) );
  XOR U17083 ( .A(n17579), .B(n17578), .Z(n17577) );
  NOR U17084 ( .A(n9159), .B(p_input[427]), .Z(n17578) );
  XOR U17085 ( .A(n17581), .B(n17580), .Z(n17579) );
  NOR U17086 ( .A(n9161), .B(p_input[425]), .Z(n17580) );
  XOR U17087 ( .A(n17583), .B(n17582), .Z(n17581) );
  NOR U17088 ( .A(n9163), .B(p_input[423]), .Z(n17582) );
  XOR U17089 ( .A(n17585), .B(n17584), .Z(n17583) );
  NOR U17090 ( .A(n9165), .B(p_input[421]), .Z(n17584) );
  XOR U17091 ( .A(n17587), .B(n17586), .Z(n17585) );
  NOR U17092 ( .A(n9167), .B(p_input[419]), .Z(n17586) );
  XOR U17093 ( .A(n17589), .B(n17588), .Z(n17587) );
  NOR U17094 ( .A(n9169), .B(p_input[417]), .Z(n17588) );
  XOR U17095 ( .A(n17591), .B(n17590), .Z(n17589) );
  NOR U17096 ( .A(n9171), .B(p_input[415]), .Z(n17590) );
  XOR U17097 ( .A(n17593), .B(n17592), .Z(n17591) );
  NOR U17098 ( .A(n9173), .B(p_input[413]), .Z(n17592) );
  XOR U17099 ( .A(n17595), .B(n17594), .Z(n17593) );
  NOR U17100 ( .A(n9175), .B(p_input[411]), .Z(n17594) );
  XOR U17101 ( .A(n17597), .B(n17596), .Z(n17595) );
  NOR U17102 ( .A(n9177), .B(p_input[409]), .Z(n17596) );
  XOR U17103 ( .A(n17599), .B(n17598), .Z(n17597) );
  NOR U17104 ( .A(n9179), .B(p_input[407]), .Z(n17598) );
  XOR U17105 ( .A(n17601), .B(n17600), .Z(n17599) );
  NOR U17106 ( .A(n9181), .B(p_input[405]), .Z(n17600) );
  XOR U17107 ( .A(n17603), .B(n17602), .Z(n17601) );
  NOR U17108 ( .A(n9183), .B(p_input[403]), .Z(n17602) );
  XOR U17109 ( .A(n17605), .B(n17604), .Z(n17603) );
  NOR U17110 ( .A(n9185), .B(p_input[401]), .Z(n17604) );
  XOR U17111 ( .A(n17607), .B(n17606), .Z(n17605) );
  NOR U17112 ( .A(n9187), .B(p_input[399]), .Z(n17606) );
  XOR U17113 ( .A(n17609), .B(n17608), .Z(n17607) );
  NOR U17114 ( .A(n9189), .B(p_input[397]), .Z(n17608) );
  XOR U17115 ( .A(n17611), .B(n17610), .Z(n17609) );
  NOR U17116 ( .A(n9191), .B(p_input[395]), .Z(n17610) );
  XOR U17117 ( .A(n17613), .B(n17612), .Z(n17611) );
  NOR U17118 ( .A(n9193), .B(p_input[393]), .Z(n17612) );
  XOR U17119 ( .A(n17615), .B(n17614), .Z(n17613) );
  NOR U17120 ( .A(n9195), .B(p_input[391]), .Z(n17614) );
  XOR U17121 ( .A(n17617), .B(n17616), .Z(n17615) );
  NOR U17122 ( .A(n9197), .B(p_input[389]), .Z(n17616) );
  XOR U17123 ( .A(n17619), .B(n17618), .Z(n17617) );
  NOR U17124 ( .A(n9199), .B(p_input[387]), .Z(n17618) );
  XOR U17125 ( .A(n17621), .B(n17620), .Z(n17619) );
  NOR U17126 ( .A(n9201), .B(p_input[385]), .Z(n17620) );
  XOR U17127 ( .A(n17623), .B(n17622), .Z(n17621) );
  NOR U17128 ( .A(n9203), .B(p_input[383]), .Z(n17622) );
  XOR U17129 ( .A(n17625), .B(n17624), .Z(n17623) );
  NOR U17130 ( .A(n9205), .B(p_input[381]), .Z(n17624) );
  XOR U17131 ( .A(n17627), .B(n17626), .Z(n17625) );
  NOR U17132 ( .A(n9207), .B(p_input[379]), .Z(n17626) );
  XOR U17133 ( .A(n17629), .B(n17628), .Z(n17627) );
  NOR U17134 ( .A(n9209), .B(p_input[377]), .Z(n17628) );
  XOR U17135 ( .A(n17631), .B(n17630), .Z(n17629) );
  NOR U17136 ( .A(n9211), .B(p_input[375]), .Z(n17630) );
  XOR U17137 ( .A(n17633), .B(n17632), .Z(n17631) );
  NOR U17138 ( .A(n9213), .B(p_input[373]), .Z(n17632) );
  XOR U17139 ( .A(n17635), .B(n17634), .Z(n17633) );
  NOR U17140 ( .A(n9215), .B(p_input[371]), .Z(n17634) );
  XOR U17141 ( .A(n17637), .B(n17636), .Z(n17635) );
  NOR U17142 ( .A(n9217), .B(p_input[369]), .Z(n17636) );
  XOR U17143 ( .A(n17639), .B(n17638), .Z(n17637) );
  NOR U17144 ( .A(n9219), .B(p_input[367]), .Z(n17638) );
  XOR U17145 ( .A(n17641), .B(n17640), .Z(n17639) );
  NOR U17146 ( .A(n9221), .B(p_input[365]), .Z(n17640) );
  XOR U17147 ( .A(n17643), .B(n17642), .Z(n17641) );
  NOR U17148 ( .A(n9223), .B(p_input[363]), .Z(n17642) );
  XOR U17149 ( .A(n17645), .B(n17644), .Z(n17643) );
  NOR U17150 ( .A(n9225), .B(p_input[361]), .Z(n17644) );
  XOR U17151 ( .A(n17647), .B(n17646), .Z(n17645) );
  NOR U17152 ( .A(n9227), .B(p_input[359]), .Z(n17646) );
  XOR U17153 ( .A(n17649), .B(n17648), .Z(n17647) );
  NOR U17154 ( .A(n9229), .B(p_input[357]), .Z(n17648) );
  XOR U17155 ( .A(n17651), .B(n17650), .Z(n17649) );
  NOR U17156 ( .A(n9231), .B(p_input[355]), .Z(n17650) );
  XOR U17157 ( .A(n17653), .B(n17652), .Z(n17651) );
  NOR U17158 ( .A(n9233), .B(p_input[353]), .Z(n17652) );
  XOR U17159 ( .A(n17655), .B(n17654), .Z(n17653) );
  NOR U17160 ( .A(n9235), .B(p_input[351]), .Z(n17654) );
  XOR U17161 ( .A(n17657), .B(n17656), .Z(n17655) );
  NOR U17162 ( .A(n9237), .B(p_input[349]), .Z(n17656) );
  XOR U17163 ( .A(n17659), .B(n17658), .Z(n17657) );
  NOR U17164 ( .A(n9239), .B(p_input[347]), .Z(n17658) );
  XOR U17165 ( .A(n17661), .B(n17660), .Z(n17659) );
  NOR U17166 ( .A(n9241), .B(p_input[345]), .Z(n17660) );
  XOR U17167 ( .A(n17663), .B(n17662), .Z(n17661) );
  NOR U17168 ( .A(n9243), .B(p_input[343]), .Z(n17662) );
  XOR U17169 ( .A(n17665), .B(n17664), .Z(n17663) );
  NOR U17170 ( .A(n9245), .B(p_input[341]), .Z(n17664) );
  XOR U17171 ( .A(n17667), .B(n17666), .Z(n17665) );
  NOR U17172 ( .A(n9247), .B(p_input[339]), .Z(n17666) );
  XOR U17173 ( .A(n17669), .B(n17668), .Z(n17667) );
  NOR U17174 ( .A(n9249), .B(p_input[337]), .Z(n17668) );
  XOR U17175 ( .A(n17671), .B(n17670), .Z(n17669) );
  NOR U17176 ( .A(n9251), .B(p_input[335]), .Z(n17670) );
  XOR U17177 ( .A(n17673), .B(n17672), .Z(n17671) );
  NOR U17178 ( .A(n9253), .B(p_input[333]), .Z(n17672) );
  XOR U17179 ( .A(n17675), .B(n17674), .Z(n17673) );
  NOR U17180 ( .A(n9255), .B(p_input[331]), .Z(n17674) );
  XOR U17181 ( .A(n17677), .B(n17676), .Z(n17675) );
  NOR U17182 ( .A(n9257), .B(p_input[329]), .Z(n17676) );
  XOR U17183 ( .A(n17679), .B(n17678), .Z(n17677) );
  NOR U17184 ( .A(n9259), .B(p_input[327]), .Z(n17678) );
  XOR U17185 ( .A(n17681), .B(n17680), .Z(n17679) );
  NOR U17186 ( .A(n9261), .B(p_input[325]), .Z(n17680) );
  XOR U17187 ( .A(n17683), .B(n17682), .Z(n17681) );
  NOR U17188 ( .A(n9263), .B(p_input[323]), .Z(n17682) );
  XOR U17189 ( .A(n17685), .B(n17684), .Z(n17683) );
  NOR U17190 ( .A(n9265), .B(p_input[321]), .Z(n17684) );
  XOR U17191 ( .A(n17687), .B(n17686), .Z(n17685) );
  NOR U17192 ( .A(n9267), .B(p_input[319]), .Z(n17686) );
  XOR U17193 ( .A(n17689), .B(n17688), .Z(n17687) );
  NOR U17194 ( .A(n9269), .B(p_input[317]), .Z(n17688) );
  XOR U17195 ( .A(n17691), .B(n17690), .Z(n17689) );
  NOR U17196 ( .A(n9271), .B(p_input[315]), .Z(n17690) );
  XOR U17197 ( .A(n17693), .B(n17692), .Z(n17691) );
  NOR U17198 ( .A(n9273), .B(p_input[313]), .Z(n17692) );
  XOR U17199 ( .A(n17695), .B(n17694), .Z(n17693) );
  NOR U17200 ( .A(n9275), .B(p_input[311]), .Z(n17694) );
  XOR U17201 ( .A(n17697), .B(n17696), .Z(n17695) );
  NOR U17202 ( .A(n9277), .B(p_input[309]), .Z(n17696) );
  XOR U17203 ( .A(n17699), .B(n17698), .Z(n17697) );
  NOR U17204 ( .A(n9279), .B(p_input[307]), .Z(n17698) );
  XOR U17205 ( .A(n17701), .B(n17700), .Z(n17699) );
  NOR U17206 ( .A(n9281), .B(p_input[305]), .Z(n17700) );
  XOR U17207 ( .A(n17703), .B(n17702), .Z(n17701) );
  NOR U17208 ( .A(n9283), .B(p_input[303]), .Z(n17702) );
  XOR U17209 ( .A(n17705), .B(n17704), .Z(n17703) );
  NOR U17210 ( .A(n9285), .B(p_input[301]), .Z(n17704) );
  XOR U17211 ( .A(n17707), .B(n17706), .Z(n17705) );
  NOR U17212 ( .A(n9287), .B(p_input[299]), .Z(n17706) );
  XOR U17213 ( .A(n17709), .B(n17708), .Z(n17707) );
  NOR U17214 ( .A(n9289), .B(p_input[297]), .Z(n17708) );
  XOR U17215 ( .A(n17711), .B(n17710), .Z(n17709) );
  NOR U17216 ( .A(n9291), .B(p_input[295]), .Z(n17710) );
  XOR U17217 ( .A(n17713), .B(n17712), .Z(n17711) );
  NOR U17218 ( .A(n9293), .B(p_input[293]), .Z(n17712) );
  XOR U17219 ( .A(n17715), .B(n17714), .Z(n17713) );
  NOR U17220 ( .A(n9295), .B(p_input[291]), .Z(n17714) );
  XOR U17221 ( .A(n17717), .B(n17716), .Z(n17715) );
  NOR U17222 ( .A(n9297), .B(p_input[289]), .Z(n17716) );
  XOR U17223 ( .A(n17719), .B(n17718), .Z(n17717) );
  NOR U17224 ( .A(n9299), .B(p_input[287]), .Z(n17718) );
  XOR U17225 ( .A(n17721), .B(n17720), .Z(n17719) );
  NOR U17226 ( .A(n9301), .B(p_input[285]), .Z(n17720) );
  XOR U17227 ( .A(n17723), .B(n17722), .Z(n17721) );
  NOR U17228 ( .A(n9303), .B(p_input[283]), .Z(n17722) );
  XOR U17229 ( .A(n17725), .B(n17724), .Z(n17723) );
  NOR U17230 ( .A(n9305), .B(p_input[281]), .Z(n17724) );
  XOR U17231 ( .A(n17727), .B(n17726), .Z(n17725) );
  NOR U17232 ( .A(n9307), .B(p_input[279]), .Z(n17726) );
  XOR U17233 ( .A(n17729), .B(n17728), .Z(n17727) );
  NOR U17234 ( .A(n9309), .B(p_input[277]), .Z(n17728) );
  XOR U17235 ( .A(n17731), .B(n17730), .Z(n17729) );
  NOR U17236 ( .A(n9311), .B(p_input[275]), .Z(n17730) );
  XOR U17237 ( .A(n17733), .B(n17732), .Z(n17731) );
  NOR U17238 ( .A(n9313), .B(p_input[273]), .Z(n17732) );
  XOR U17239 ( .A(n17735), .B(n17734), .Z(n17733) );
  NOR U17240 ( .A(n9315), .B(p_input[271]), .Z(n17734) );
  XOR U17241 ( .A(n17737), .B(n17736), .Z(n17735) );
  NOR U17242 ( .A(n9317), .B(p_input[269]), .Z(n17736) );
  XOR U17243 ( .A(n17739), .B(n17738), .Z(n17737) );
  NOR U17244 ( .A(n9319), .B(p_input[267]), .Z(n17738) );
  XOR U17245 ( .A(n17741), .B(n17740), .Z(n17739) );
  NOR U17246 ( .A(n9321), .B(p_input[265]), .Z(n17740) );
  XOR U17247 ( .A(n17743), .B(n17742), .Z(n17741) );
  NOR U17248 ( .A(n9323), .B(p_input[263]), .Z(n17742) );
  XOR U17249 ( .A(n17745), .B(n17744), .Z(n17743) );
  NOR U17250 ( .A(n9325), .B(p_input[261]), .Z(n17744) );
  XOR U17251 ( .A(n17747), .B(n17746), .Z(n17745) );
  NOR U17252 ( .A(n9327), .B(p_input[259]), .Z(n17746) );
  XOR U17253 ( .A(n17749), .B(n17748), .Z(n17747) );
  NOR U17254 ( .A(n9329), .B(p_input[257]), .Z(n17748) );
  XOR U17255 ( .A(n17751), .B(n17750), .Z(n17749) );
  NOR U17256 ( .A(n9331), .B(p_input[255]), .Z(n17750) );
  XOR U17257 ( .A(n17755), .B(n17754), .Z(n17751) );
  NOR U17258 ( .A(n9333), .B(p_input[253]), .Z(n17754) );
  XOR U17259 ( .A(n17757), .B(n17756), .Z(n17755) );
  NOR U17260 ( .A(n9335), .B(p_input[251]), .Z(n17756) );
  XOR U17261 ( .A(n17759), .B(n17758), .Z(n17757) );
  NOR U17262 ( .A(n9337), .B(p_input[249]), .Z(n17758) );
  XOR U17263 ( .A(n17761), .B(n17760), .Z(n17759) );
  NOR U17264 ( .A(n9339), .B(p_input[247]), .Z(n17760) );
  XOR U17265 ( .A(n17763), .B(n17762), .Z(n17761) );
  NOR U17266 ( .A(n9341), .B(p_input[245]), .Z(n17762) );
  XOR U17267 ( .A(n17765), .B(n17764), .Z(n17763) );
  NOR U17268 ( .A(n9343), .B(p_input[243]), .Z(n17764) );
  XOR U17269 ( .A(n17767), .B(n17766), .Z(n17765) );
  NOR U17270 ( .A(n9345), .B(p_input[241]), .Z(n17766) );
  XOR U17271 ( .A(n17769), .B(n17768), .Z(n17767) );
  NOR U17272 ( .A(n9347), .B(p_input[239]), .Z(n17768) );
  XOR U17273 ( .A(n17771), .B(n17770), .Z(n17769) );
  NOR U17274 ( .A(n9349), .B(p_input[237]), .Z(n17770) );
  XOR U17275 ( .A(n17773), .B(n17772), .Z(n17771) );
  NOR U17276 ( .A(n9351), .B(p_input[235]), .Z(n17772) );
  XOR U17277 ( .A(n17775), .B(n17774), .Z(n17773) );
  NOR U17278 ( .A(n9353), .B(p_input[233]), .Z(n17774) );
  XOR U17279 ( .A(n17777), .B(n17776), .Z(n17775) );
  NOR U17280 ( .A(n9355), .B(p_input[231]), .Z(n17776) );
  XOR U17281 ( .A(n17779), .B(n17778), .Z(n17777) );
  NOR U17282 ( .A(n9357), .B(p_input[229]), .Z(n17778) );
  XOR U17283 ( .A(n17781), .B(n17780), .Z(n17779) );
  NOR U17284 ( .A(n9359), .B(p_input[227]), .Z(n17780) );
  XOR U17285 ( .A(n17783), .B(n17782), .Z(n17781) );
  NOR U17286 ( .A(n9361), .B(p_input[225]), .Z(n17782) );
  XOR U17287 ( .A(n17785), .B(n17784), .Z(n17783) );
  NOR U17288 ( .A(n9363), .B(p_input[223]), .Z(n17784) );
  XOR U17289 ( .A(n17787), .B(n17786), .Z(n17785) );
  NOR U17290 ( .A(n9365), .B(p_input[221]), .Z(n17786) );
  XOR U17291 ( .A(n17789), .B(n17788), .Z(n17787) );
  NOR U17292 ( .A(n9367), .B(p_input[219]), .Z(n17788) );
  XOR U17293 ( .A(n17791), .B(n17790), .Z(n17789) );
  NOR U17294 ( .A(n9369), .B(p_input[217]), .Z(n17790) );
  XOR U17295 ( .A(n17793), .B(n17792), .Z(n17791) );
  NOR U17296 ( .A(n9371), .B(p_input[215]), .Z(n17792) );
  XOR U17297 ( .A(n17795), .B(n17794), .Z(n17793) );
  NOR U17298 ( .A(n9373), .B(p_input[213]), .Z(n17794) );
  XOR U17299 ( .A(n17797), .B(n17796), .Z(n17795) );
  NOR U17300 ( .A(n9375), .B(p_input[211]), .Z(n17796) );
  XOR U17301 ( .A(n17799), .B(n17798), .Z(n17797) );
  NOR U17302 ( .A(n9377), .B(p_input[209]), .Z(n17798) );
  XOR U17303 ( .A(n17801), .B(n17800), .Z(n17799) );
  NOR U17304 ( .A(n9379), .B(p_input[207]), .Z(n17800) );
  XOR U17305 ( .A(n17803), .B(n17802), .Z(n17801) );
  NOR U17306 ( .A(n9381), .B(p_input[205]), .Z(n17802) );
  XOR U17307 ( .A(n17805), .B(n17804), .Z(n17803) );
  NOR U17308 ( .A(n9383), .B(p_input[203]), .Z(n17804) );
  XOR U17309 ( .A(n17807), .B(n17806), .Z(n17805) );
  NOR U17310 ( .A(n9385), .B(p_input[201]), .Z(n17806) );
  XOR U17311 ( .A(n17809), .B(n17808), .Z(n17807) );
  NOR U17312 ( .A(n9387), .B(p_input[199]), .Z(n17808) );
  XOR U17313 ( .A(n17811), .B(n17810), .Z(n17809) );
  NOR U17314 ( .A(n9389), .B(p_input[197]), .Z(n17810) );
  XOR U17315 ( .A(n17813), .B(n17812), .Z(n17811) );
  NOR U17316 ( .A(n9391), .B(p_input[195]), .Z(n17812) );
  XOR U17317 ( .A(n17815), .B(n17814), .Z(n17813) );
  NOR U17318 ( .A(n9393), .B(p_input[193]), .Z(n17814) );
  XOR U17319 ( .A(n17817), .B(n17816), .Z(n17815) );
  NOR U17320 ( .A(n9395), .B(p_input[191]), .Z(n17816) );
  XOR U17321 ( .A(n17819), .B(n17818), .Z(n17817) );
  NOR U17322 ( .A(n9397), .B(p_input[189]), .Z(n17818) );
  XOR U17323 ( .A(n17821), .B(n17820), .Z(n17819) );
  NOR U17324 ( .A(n9399), .B(p_input[187]), .Z(n17820) );
  XOR U17325 ( .A(n17823), .B(n17822), .Z(n17821) );
  NOR U17326 ( .A(n9401), .B(p_input[185]), .Z(n17822) );
  XOR U17327 ( .A(n17825), .B(n17824), .Z(n17823) );
  NOR U17328 ( .A(n9403), .B(p_input[183]), .Z(n17824) );
  XOR U17329 ( .A(n17827), .B(n17826), .Z(n17825) );
  NOR U17330 ( .A(n9405), .B(p_input[181]), .Z(n17826) );
  XOR U17331 ( .A(n17829), .B(n17828), .Z(n17827) );
  NOR U17332 ( .A(n9407), .B(p_input[179]), .Z(n17828) );
  XOR U17333 ( .A(n17831), .B(n17830), .Z(n17829) );
  NOR U17334 ( .A(n9409), .B(p_input[177]), .Z(n17830) );
  XOR U17335 ( .A(n17833), .B(n17832), .Z(n17831) );
  NOR U17336 ( .A(n9411), .B(p_input[175]), .Z(n17832) );
  XOR U17337 ( .A(n17835), .B(n17834), .Z(n17833) );
  NOR U17338 ( .A(n9413), .B(p_input[173]), .Z(n17834) );
  XOR U17339 ( .A(n17837), .B(n17836), .Z(n17835) );
  NOR U17340 ( .A(n9415), .B(p_input[171]), .Z(n17836) );
  XOR U17341 ( .A(n17839), .B(n17838), .Z(n17837) );
  NOR U17342 ( .A(n9417), .B(p_input[169]), .Z(n17838) );
  XOR U17343 ( .A(n17841), .B(n17840), .Z(n17839) );
  NOR U17344 ( .A(n9419), .B(p_input[167]), .Z(n17840) );
  XOR U17345 ( .A(n17843), .B(n17842), .Z(n17841) );
  NOR U17346 ( .A(n9421), .B(p_input[165]), .Z(n17842) );
  XOR U17347 ( .A(n17845), .B(n17844), .Z(n17843) );
  NOR U17348 ( .A(n9423), .B(p_input[163]), .Z(n17844) );
  XOR U17349 ( .A(n17847), .B(n17846), .Z(n17845) );
  NOR U17350 ( .A(n9425), .B(p_input[161]), .Z(n17846) );
  XOR U17351 ( .A(n17849), .B(n17848), .Z(n17847) );
  NOR U17352 ( .A(n9427), .B(p_input[159]), .Z(n17848) );
  XOR U17353 ( .A(n17851), .B(n17850), .Z(n17849) );
  NOR U17354 ( .A(n9429), .B(p_input[157]), .Z(n17850) );
  XOR U17355 ( .A(n17853), .B(n17852), .Z(n17851) );
  NOR U17356 ( .A(n9431), .B(p_input[155]), .Z(n17852) );
  XOR U17357 ( .A(n17855), .B(n17854), .Z(n17853) );
  NOR U17358 ( .A(n9433), .B(p_input[153]), .Z(n17854) );
  XOR U17359 ( .A(n17857), .B(n17856), .Z(n17855) );
  NOR U17360 ( .A(n9435), .B(p_input[151]), .Z(n17856) );
  XOR U17361 ( .A(n17859), .B(n17858), .Z(n17857) );
  NOR U17362 ( .A(n9437), .B(p_input[149]), .Z(n17858) );
  XOR U17363 ( .A(n17861), .B(n17860), .Z(n17859) );
  NOR U17364 ( .A(n9439), .B(p_input[147]), .Z(n17860) );
  XOR U17365 ( .A(n17863), .B(n17862), .Z(n17861) );
  NOR U17366 ( .A(n9441), .B(p_input[145]), .Z(n17862) );
  XOR U17367 ( .A(n17865), .B(n17864), .Z(n17863) );
  NOR U17368 ( .A(n9443), .B(p_input[143]), .Z(n17864) );
  XOR U17369 ( .A(n17867), .B(n17866), .Z(n17865) );
  NOR U17370 ( .A(n9445), .B(p_input[141]), .Z(n17866) );
  XOR U17371 ( .A(n17869), .B(n17868), .Z(n17867) );
  NOR U17372 ( .A(n9447), .B(p_input[139]), .Z(n17868) );
  XOR U17373 ( .A(n17871), .B(n17870), .Z(n17869) );
  NOR U17374 ( .A(n9449), .B(p_input[137]), .Z(n17870) );
  XOR U17375 ( .A(n17873), .B(n17872), .Z(n17871) );
  NOR U17376 ( .A(n9451), .B(p_input[135]), .Z(n17872) );
  XOR U17377 ( .A(n17875), .B(n17874), .Z(n17873) );
  NOR U17378 ( .A(n9453), .B(p_input[133]), .Z(n17874) );
  XOR U17379 ( .A(n17877), .B(n17876), .Z(n17875) );
  NOR U17380 ( .A(n9455), .B(p_input[131]), .Z(n17876) );
  XOR U17381 ( .A(n17879), .B(n17878), .Z(n17877) );
  NOR U17382 ( .A(n9457), .B(p_input[129]), .Z(n17878) );
  XOR U17383 ( .A(n17881), .B(n17880), .Z(n17879) );
  NOR U17384 ( .A(n9459), .B(p_input[127]), .Z(n17880) );
  XOR U17385 ( .A(n17883), .B(n17882), .Z(n17881) );
  NOR U17386 ( .A(n9461), .B(p_input[125]), .Z(n17882) );
  XOR U17387 ( .A(n17885), .B(n17884), .Z(n17883) );
  NOR U17388 ( .A(n9463), .B(p_input[123]), .Z(n17884) );
  XOR U17389 ( .A(n17887), .B(n17886), .Z(n17885) );
  NOR U17390 ( .A(n9465), .B(p_input[121]), .Z(n17886) );
  XOR U17391 ( .A(n17889), .B(n17888), .Z(n17887) );
  NOR U17392 ( .A(n9467), .B(p_input[119]), .Z(n17888) );
  XOR U17393 ( .A(n17891), .B(n17890), .Z(n17889) );
  NOR U17394 ( .A(n9469), .B(p_input[117]), .Z(n17890) );
  XOR U17395 ( .A(n17893), .B(n17892), .Z(n17891) );
  NOR U17396 ( .A(n9471), .B(p_input[115]), .Z(n17892) );
  XOR U17397 ( .A(n17895), .B(n17894), .Z(n17893) );
  NOR U17398 ( .A(n9473), .B(p_input[113]), .Z(n17894) );
  XOR U17399 ( .A(n17897), .B(n17896), .Z(n17895) );
  NOR U17400 ( .A(n9475), .B(p_input[111]), .Z(n17896) );
  XOR U17401 ( .A(n17899), .B(n17898), .Z(n17897) );
  NOR U17402 ( .A(n9477), .B(p_input[109]), .Z(n17898) );
  XOR U17403 ( .A(n17901), .B(n17900), .Z(n17899) );
  NOR U17404 ( .A(n9479), .B(p_input[107]), .Z(n17900) );
  XOR U17405 ( .A(n17903), .B(n17902), .Z(n17901) );
  NOR U17406 ( .A(n9481), .B(p_input[105]), .Z(n17902) );
  XOR U17407 ( .A(n17905), .B(n17904), .Z(n17903) );
  NOR U17408 ( .A(n9483), .B(p_input[103]), .Z(n17904) );
  XOR U17409 ( .A(n17907), .B(n17906), .Z(n17905) );
  NOR U17410 ( .A(n9485), .B(p_input[101]), .Z(n17906) );
  XOR U17411 ( .A(n17909), .B(n17908), .Z(n17907) );
  NOR U17412 ( .A(n9487), .B(p_input[99]), .Z(n17908) );
  XOR U17413 ( .A(n17911), .B(n17910), .Z(n17909) );
  NOR U17414 ( .A(n9489), .B(p_input[97]), .Z(n17910) );
  XOR U17415 ( .A(n17913), .B(n17912), .Z(n17911) );
  NOR U17416 ( .A(n9491), .B(p_input[95]), .Z(n17912) );
  XOR U17417 ( .A(n17915), .B(n17914), .Z(n17913) );
  NOR U17418 ( .A(n9493), .B(p_input[93]), .Z(n17914) );
  XOR U17419 ( .A(n17917), .B(n17916), .Z(n17915) );
  NOR U17420 ( .A(n9495), .B(p_input[91]), .Z(n17916) );
  XOR U17421 ( .A(n17919), .B(n17918), .Z(n17917) );
  NOR U17422 ( .A(n9497), .B(p_input[89]), .Z(n17918) );
  XOR U17423 ( .A(n17921), .B(n17920), .Z(n17919) );
  NOR U17424 ( .A(n9499), .B(p_input[87]), .Z(n17920) );
  XOR U17425 ( .A(n17923), .B(n17922), .Z(n17921) );
  NOR U17426 ( .A(n9501), .B(p_input[85]), .Z(n17922) );
  XOR U17427 ( .A(n17925), .B(n17924), .Z(n17923) );
  NOR U17428 ( .A(n9503), .B(p_input[83]), .Z(n17924) );
  XOR U17429 ( .A(n17927), .B(n17926), .Z(n17925) );
  NOR U17430 ( .A(n9505), .B(p_input[81]), .Z(n17926) );
  XOR U17431 ( .A(n17929), .B(n17928), .Z(n17927) );
  NOR U17432 ( .A(n9507), .B(p_input[79]), .Z(n17928) );
  XOR U17433 ( .A(n17931), .B(n17930), .Z(n17929) );
  NOR U17434 ( .A(n9509), .B(p_input[77]), .Z(n17930) );
  XOR U17435 ( .A(n17933), .B(n17932), .Z(n17931) );
  NOR U17436 ( .A(n9511), .B(p_input[75]), .Z(n17932) );
  XOR U17437 ( .A(n17935), .B(n17934), .Z(n17933) );
  NOR U17438 ( .A(n9513), .B(p_input[73]), .Z(n17934) );
  XOR U17439 ( .A(n17937), .B(n17936), .Z(n17935) );
  NOR U17440 ( .A(n9515), .B(p_input[71]), .Z(n17936) );
  XOR U17441 ( .A(n17939), .B(n17938), .Z(n17937) );
  NOR U17442 ( .A(n9517), .B(p_input[69]), .Z(n17938) );
  XOR U17443 ( .A(n17941), .B(n17940), .Z(n17939) );
  NOR U17444 ( .A(n9519), .B(p_input[67]), .Z(n17940) );
  XOR U17445 ( .A(n17943), .B(n17942), .Z(n17941) );
  NOR U17446 ( .A(n9521), .B(p_input[65]), .Z(n17942) );
  XOR U17447 ( .A(n17945), .B(n17944), .Z(n17943) );
  NOR U17448 ( .A(n9523), .B(p_input[63]), .Z(n17944) );
  XOR U17449 ( .A(n17947), .B(n17946), .Z(n17945) );
  NOR U17450 ( .A(n9525), .B(p_input[61]), .Z(n17946) );
  XOR U17451 ( .A(n17949), .B(n17948), .Z(n17947) );
  NOR U17452 ( .A(n9527), .B(p_input[59]), .Z(n17948) );
  XOR U17453 ( .A(n17951), .B(n17950), .Z(n17949) );
  NOR U17454 ( .A(n9529), .B(p_input[57]), .Z(n17950) );
  XOR U17455 ( .A(n17953), .B(n17952), .Z(n17951) );
  NOR U17456 ( .A(n9531), .B(p_input[55]), .Z(n17952) );
  XOR U17457 ( .A(n17955), .B(n17954), .Z(n17953) );
  NOR U17458 ( .A(n9533), .B(p_input[53]), .Z(n17954) );
  XOR U17459 ( .A(n17957), .B(n17956), .Z(n17955) );
  NOR U17460 ( .A(n9535), .B(p_input[51]), .Z(n17956) );
  XOR U17461 ( .A(n17959), .B(n17958), .Z(n17957) );
  NOR U17462 ( .A(n9537), .B(p_input[49]), .Z(n17958) );
  XOR U17463 ( .A(n17961), .B(n17960), .Z(n17959) );
  NOR U17464 ( .A(n9539), .B(p_input[47]), .Z(n17960) );
  XOR U17465 ( .A(n17963), .B(n17962), .Z(n17961) );
  NOR U17466 ( .A(n9541), .B(p_input[45]), .Z(n17962) );
  XOR U17467 ( .A(n17965), .B(n17964), .Z(n17963) );
  NOR U17468 ( .A(n9543), .B(p_input[43]), .Z(n17964) );
  XOR U17469 ( .A(n17967), .B(n17966), .Z(n17965) );
  NOR U17470 ( .A(n9545), .B(p_input[41]), .Z(n17966) );
  XOR U17471 ( .A(n17969), .B(n17968), .Z(n17967) );
  NOR U17472 ( .A(n9547), .B(p_input[39]), .Z(n17968) );
  XOR U17473 ( .A(n17971), .B(n17970), .Z(n17969) );
  NOR U17474 ( .A(n9549), .B(p_input[37]), .Z(n17970) );
  XOR U17475 ( .A(n17973), .B(n17972), .Z(n17971) );
  NOR U17476 ( .A(n9551), .B(p_input[35]), .Z(n17972) );
  XOR U17477 ( .A(n17975), .B(n17974), .Z(n17973) );
  NOR U17478 ( .A(n9553), .B(p_input[33]), .Z(n17974) );
  XOR U17479 ( .A(n17977), .B(n17976), .Z(n17975) );
  NOR U17480 ( .A(n9555), .B(p_input[31]), .Z(n17976) );
  XOR U17481 ( .A(n17979), .B(n17978), .Z(n17977) );
  NOR U17482 ( .A(n9557), .B(p_input[29]), .Z(n17978) );
  XOR U17483 ( .A(n17981), .B(n17980), .Z(n17979) );
  NOR U17484 ( .A(n9559), .B(p_input[27]), .Z(n17980) );
  XOR U17485 ( .A(n17983), .B(n17982), .Z(n17981) );
  NOR U17486 ( .A(n9561), .B(p_input[25]), .Z(n17982) );
  XOR U17487 ( .A(n17985), .B(n17984), .Z(n17983) );
  NOR U17488 ( .A(n9563), .B(p_input[23]), .Z(n17984) );
  XOR U17489 ( .A(n17987), .B(n17986), .Z(n17985) );
  NOR U17490 ( .A(n9565), .B(p_input[21]), .Z(n17986) );
  XOR U17491 ( .A(n17989), .B(n17988), .Z(n17987) );
  NOR U17492 ( .A(n9567), .B(p_input[19]), .Z(n17988) );
  XOR U17493 ( .A(n17991), .B(n17990), .Z(n17989) );
  NOR U17494 ( .A(n9569), .B(p_input[17]), .Z(n17990) );
  XOR U17495 ( .A(n17993), .B(n17992), .Z(n17991) );
  NOR U17496 ( .A(n9571), .B(p_input[15]), .Z(n17992) );
  XOR U17497 ( .A(n17995), .B(n17994), .Z(n17993) );
  NOR U17498 ( .A(n9573), .B(p_input[13]), .Z(n17994) );
  XOR U17499 ( .A(n18009), .B(n18008), .Z(n17995) );
  NOR U17500 ( .A(n9575), .B(p_input[11]), .Z(n18008) );
  XOR U17501 ( .A(n18011), .B(n18010), .Z(n18009) );
  NOR U17502 ( .A(n9577), .B(p_input[9]), .Z(n18010) );
  XOR U17503 ( .A(n17999), .B(n17998), .Z(n18011) );
  NOR U17504 ( .A(n9579), .B(p_input[7]), .Z(n17998) );
  XOR U17505 ( .A(n18006), .B(n18007), .Z(n17999) );
  XOR U17506 ( .A(n18004), .B(n18005), .Z(n18007) );
  NOR U17507 ( .A(n9581), .B(p_input[3]), .Z(n18005) );
  NOR U17508 ( .A(n9583), .B(p_input[1]), .Z(n18004) );
  NOR U17509 ( .A(n9585), .B(p_input[5]), .Z(n18006) );
  XOR U17510 ( .A(n18013), .B(n18012), .Z(n9586) );
  AND U17511 ( .A(n9074), .B(n9075), .Z(n18012) );
  IV U17512 ( .A(p_input[510]), .Z(n9075) );
  IV U17513 ( .A(p_input[511]), .Z(n9074) );
  XOR U17514 ( .A(n18015), .B(n18014), .Z(n18013) );
  AND U17515 ( .A(n9076), .B(n9077), .Z(n18014) );
  IV U17516 ( .A(p_input[508]), .Z(n9077) );
  IV U17517 ( .A(p_input[509]), .Z(n9076) );
  XOR U17518 ( .A(n18017), .B(n18016), .Z(n18015) );
  AND U17519 ( .A(n9078), .B(n9079), .Z(n18016) );
  IV U17520 ( .A(p_input[506]), .Z(n9079) );
  IV U17521 ( .A(p_input[507]), .Z(n9078) );
  XOR U17522 ( .A(n18019), .B(n18018), .Z(n18017) );
  AND U17523 ( .A(n9080), .B(n9081), .Z(n18018) );
  IV U17524 ( .A(p_input[504]), .Z(n9081) );
  IV U17525 ( .A(p_input[505]), .Z(n9080) );
  XOR U17526 ( .A(n18021), .B(n18020), .Z(n18019) );
  AND U17527 ( .A(n9082), .B(n9083), .Z(n18020) );
  IV U17528 ( .A(p_input[502]), .Z(n9083) );
  IV U17529 ( .A(p_input[503]), .Z(n9082) );
  XOR U17530 ( .A(n18023), .B(n18022), .Z(n18021) );
  AND U17531 ( .A(n9084), .B(n9085), .Z(n18022) );
  IV U17532 ( .A(p_input[500]), .Z(n9085) );
  IV U17533 ( .A(p_input[501]), .Z(n9084) );
  XOR U17534 ( .A(n18025), .B(n18024), .Z(n18023) );
  AND U17535 ( .A(n9086), .B(n9087), .Z(n18024) );
  IV U17536 ( .A(p_input[498]), .Z(n9087) );
  IV U17537 ( .A(p_input[499]), .Z(n9086) );
  XOR U17538 ( .A(n18027), .B(n18026), .Z(n18025) );
  AND U17539 ( .A(n9088), .B(n9089), .Z(n18026) );
  IV U17540 ( .A(p_input[496]), .Z(n9089) );
  IV U17541 ( .A(p_input[497]), .Z(n9088) );
  XOR U17542 ( .A(n18029), .B(n18028), .Z(n18027) );
  AND U17543 ( .A(n9090), .B(n9091), .Z(n18028) );
  IV U17544 ( .A(p_input[494]), .Z(n9091) );
  IV U17545 ( .A(p_input[495]), .Z(n9090) );
  XOR U17546 ( .A(n18031), .B(n18030), .Z(n18029) );
  AND U17547 ( .A(n9092), .B(n9093), .Z(n18030) );
  IV U17548 ( .A(p_input[492]), .Z(n9093) );
  IV U17549 ( .A(p_input[493]), .Z(n9092) );
  XOR U17550 ( .A(n18033), .B(n18032), .Z(n18031) );
  AND U17551 ( .A(n9094), .B(n9095), .Z(n18032) );
  IV U17552 ( .A(p_input[490]), .Z(n9095) );
  IV U17553 ( .A(p_input[491]), .Z(n9094) );
  XOR U17554 ( .A(n18035), .B(n18034), .Z(n18033) );
  AND U17555 ( .A(n9096), .B(n9097), .Z(n18034) );
  IV U17556 ( .A(p_input[488]), .Z(n9097) );
  IV U17557 ( .A(p_input[489]), .Z(n9096) );
  XOR U17558 ( .A(n18037), .B(n18036), .Z(n18035) );
  AND U17559 ( .A(n9098), .B(n9099), .Z(n18036) );
  IV U17560 ( .A(p_input[486]), .Z(n9099) );
  IV U17561 ( .A(p_input[487]), .Z(n9098) );
  XOR U17562 ( .A(n18039), .B(n18038), .Z(n18037) );
  AND U17563 ( .A(n9100), .B(n9101), .Z(n18038) );
  IV U17564 ( .A(p_input[484]), .Z(n9101) );
  IV U17565 ( .A(p_input[485]), .Z(n9100) );
  XOR U17566 ( .A(n18041), .B(n18040), .Z(n18039) );
  AND U17567 ( .A(n9102), .B(n9103), .Z(n18040) );
  IV U17568 ( .A(p_input[482]), .Z(n9103) );
  IV U17569 ( .A(p_input[483]), .Z(n9102) );
  XOR U17570 ( .A(n18043), .B(n18042), .Z(n18041) );
  AND U17571 ( .A(n9104), .B(n9105), .Z(n18042) );
  IV U17572 ( .A(p_input[480]), .Z(n9105) );
  IV U17573 ( .A(p_input[481]), .Z(n9104) );
  XOR U17574 ( .A(n18045), .B(n18044), .Z(n18043) );
  AND U17575 ( .A(n9106), .B(n9107), .Z(n18044) );
  IV U17576 ( .A(p_input[478]), .Z(n9107) );
  IV U17577 ( .A(p_input[479]), .Z(n9106) );
  XOR U17578 ( .A(n18047), .B(n18046), .Z(n18045) );
  AND U17579 ( .A(n9108), .B(n9109), .Z(n18046) );
  IV U17580 ( .A(p_input[476]), .Z(n9109) );
  IV U17581 ( .A(p_input[477]), .Z(n9108) );
  XOR U17582 ( .A(n18049), .B(n18048), .Z(n18047) );
  AND U17583 ( .A(n9110), .B(n9111), .Z(n18048) );
  IV U17584 ( .A(p_input[474]), .Z(n9111) );
  IV U17585 ( .A(p_input[475]), .Z(n9110) );
  XOR U17586 ( .A(n18051), .B(n18050), .Z(n18049) );
  AND U17587 ( .A(n9112), .B(n9113), .Z(n18050) );
  IV U17588 ( .A(p_input[472]), .Z(n9113) );
  IV U17589 ( .A(p_input[473]), .Z(n9112) );
  XOR U17590 ( .A(n18053), .B(n18052), .Z(n18051) );
  AND U17591 ( .A(n9114), .B(n9115), .Z(n18052) );
  IV U17592 ( .A(p_input[470]), .Z(n9115) );
  IV U17593 ( .A(p_input[471]), .Z(n9114) );
  XOR U17594 ( .A(n18055), .B(n18054), .Z(n18053) );
  AND U17595 ( .A(n9116), .B(n9117), .Z(n18054) );
  IV U17596 ( .A(p_input[468]), .Z(n9117) );
  IV U17597 ( .A(p_input[469]), .Z(n9116) );
  XOR U17598 ( .A(n18057), .B(n18056), .Z(n18055) );
  AND U17599 ( .A(n9118), .B(n9119), .Z(n18056) );
  IV U17600 ( .A(p_input[466]), .Z(n9119) );
  IV U17601 ( .A(p_input[467]), .Z(n9118) );
  XOR U17602 ( .A(n18059), .B(n18058), .Z(n18057) );
  AND U17603 ( .A(n9120), .B(n9121), .Z(n18058) );
  IV U17604 ( .A(p_input[464]), .Z(n9121) );
  IV U17605 ( .A(p_input[465]), .Z(n9120) );
  XOR U17606 ( .A(n18061), .B(n18060), .Z(n18059) );
  AND U17607 ( .A(n9122), .B(n9123), .Z(n18060) );
  IV U17608 ( .A(p_input[462]), .Z(n9123) );
  IV U17609 ( .A(p_input[463]), .Z(n9122) );
  XOR U17610 ( .A(n18063), .B(n18062), .Z(n18061) );
  AND U17611 ( .A(n9124), .B(n9125), .Z(n18062) );
  IV U17612 ( .A(p_input[460]), .Z(n9125) );
  IV U17613 ( .A(p_input[461]), .Z(n9124) );
  XOR U17614 ( .A(n18065), .B(n18064), .Z(n18063) );
  AND U17615 ( .A(n9126), .B(n9127), .Z(n18064) );
  IV U17616 ( .A(p_input[458]), .Z(n9127) );
  IV U17617 ( .A(p_input[459]), .Z(n9126) );
  XOR U17618 ( .A(n18067), .B(n18066), .Z(n18065) );
  AND U17619 ( .A(n9128), .B(n9129), .Z(n18066) );
  IV U17620 ( .A(p_input[456]), .Z(n9129) );
  IV U17621 ( .A(p_input[457]), .Z(n9128) );
  XOR U17622 ( .A(n18069), .B(n18068), .Z(n18067) );
  AND U17623 ( .A(n9130), .B(n9131), .Z(n18068) );
  IV U17624 ( .A(p_input[454]), .Z(n9131) );
  IV U17625 ( .A(p_input[455]), .Z(n9130) );
  XOR U17626 ( .A(n18071), .B(n18070), .Z(n18069) );
  AND U17627 ( .A(n9132), .B(n9133), .Z(n18070) );
  IV U17628 ( .A(p_input[452]), .Z(n9133) );
  IV U17629 ( .A(p_input[453]), .Z(n9132) );
  XOR U17630 ( .A(n18073), .B(n18072), .Z(n18071) );
  AND U17631 ( .A(n9134), .B(n9135), .Z(n18072) );
  IV U17632 ( .A(p_input[450]), .Z(n9135) );
  IV U17633 ( .A(p_input[451]), .Z(n9134) );
  XOR U17634 ( .A(n18075), .B(n18074), .Z(n18073) );
  AND U17635 ( .A(n9136), .B(n9137), .Z(n18074) );
  IV U17636 ( .A(p_input[448]), .Z(n9137) );
  IV U17637 ( .A(p_input[449]), .Z(n9136) );
  XOR U17638 ( .A(n18077), .B(n18076), .Z(n18075) );
  AND U17639 ( .A(n9138), .B(n9139), .Z(n18076) );
  IV U17640 ( .A(p_input[446]), .Z(n9139) );
  IV U17641 ( .A(p_input[447]), .Z(n9138) );
  XOR U17642 ( .A(n18079), .B(n18078), .Z(n18077) );
  AND U17643 ( .A(n9140), .B(n9141), .Z(n18078) );
  IV U17644 ( .A(p_input[444]), .Z(n9141) );
  IV U17645 ( .A(p_input[445]), .Z(n9140) );
  XOR U17646 ( .A(n18081), .B(n18080), .Z(n18079) );
  AND U17647 ( .A(n9142), .B(n9143), .Z(n18080) );
  IV U17648 ( .A(p_input[442]), .Z(n9143) );
  IV U17649 ( .A(p_input[443]), .Z(n9142) );
  XOR U17650 ( .A(n18083), .B(n18082), .Z(n18081) );
  AND U17651 ( .A(n9144), .B(n9145), .Z(n18082) );
  IV U17652 ( .A(p_input[440]), .Z(n9145) );
  IV U17653 ( .A(p_input[441]), .Z(n9144) );
  XOR U17654 ( .A(n18085), .B(n18084), .Z(n18083) );
  AND U17655 ( .A(n9146), .B(n9147), .Z(n18084) );
  IV U17656 ( .A(p_input[438]), .Z(n9147) );
  IV U17657 ( .A(p_input[439]), .Z(n9146) );
  XOR U17658 ( .A(n18087), .B(n18086), .Z(n18085) );
  AND U17659 ( .A(n9148), .B(n9149), .Z(n18086) );
  IV U17660 ( .A(p_input[436]), .Z(n9149) );
  IV U17661 ( .A(p_input[437]), .Z(n9148) );
  XOR U17662 ( .A(n18089), .B(n18088), .Z(n18087) );
  AND U17663 ( .A(n9150), .B(n9151), .Z(n18088) );
  IV U17664 ( .A(p_input[434]), .Z(n9151) );
  IV U17665 ( .A(p_input[435]), .Z(n9150) );
  XOR U17666 ( .A(n18091), .B(n18090), .Z(n18089) );
  AND U17667 ( .A(n9152), .B(n9153), .Z(n18090) );
  IV U17668 ( .A(p_input[432]), .Z(n9153) );
  IV U17669 ( .A(p_input[433]), .Z(n9152) );
  XOR U17670 ( .A(n18093), .B(n18092), .Z(n18091) );
  AND U17671 ( .A(n9154), .B(n9155), .Z(n18092) );
  IV U17672 ( .A(p_input[430]), .Z(n9155) );
  IV U17673 ( .A(p_input[431]), .Z(n9154) );
  XOR U17674 ( .A(n18095), .B(n18094), .Z(n18093) );
  AND U17675 ( .A(n9156), .B(n9157), .Z(n18094) );
  IV U17676 ( .A(p_input[428]), .Z(n9157) );
  IV U17677 ( .A(p_input[429]), .Z(n9156) );
  XOR U17678 ( .A(n18097), .B(n18096), .Z(n18095) );
  AND U17679 ( .A(n9158), .B(n9159), .Z(n18096) );
  IV U17680 ( .A(p_input[426]), .Z(n9159) );
  IV U17681 ( .A(p_input[427]), .Z(n9158) );
  XOR U17682 ( .A(n18099), .B(n18098), .Z(n18097) );
  AND U17683 ( .A(n9160), .B(n9161), .Z(n18098) );
  IV U17684 ( .A(p_input[424]), .Z(n9161) );
  IV U17685 ( .A(p_input[425]), .Z(n9160) );
  XOR U17686 ( .A(n18101), .B(n18100), .Z(n18099) );
  AND U17687 ( .A(n9162), .B(n9163), .Z(n18100) );
  IV U17688 ( .A(p_input[422]), .Z(n9163) );
  IV U17689 ( .A(p_input[423]), .Z(n9162) );
  XOR U17690 ( .A(n18103), .B(n18102), .Z(n18101) );
  AND U17691 ( .A(n9164), .B(n9165), .Z(n18102) );
  IV U17692 ( .A(p_input[420]), .Z(n9165) );
  IV U17693 ( .A(p_input[421]), .Z(n9164) );
  XOR U17694 ( .A(n18105), .B(n18104), .Z(n18103) );
  AND U17695 ( .A(n9166), .B(n9167), .Z(n18104) );
  IV U17696 ( .A(p_input[418]), .Z(n9167) );
  IV U17697 ( .A(p_input[419]), .Z(n9166) );
  XOR U17698 ( .A(n18107), .B(n18106), .Z(n18105) );
  AND U17699 ( .A(n9168), .B(n9169), .Z(n18106) );
  IV U17700 ( .A(p_input[416]), .Z(n9169) );
  IV U17701 ( .A(p_input[417]), .Z(n9168) );
  XOR U17702 ( .A(n18109), .B(n18108), .Z(n18107) );
  AND U17703 ( .A(n9170), .B(n9171), .Z(n18108) );
  IV U17704 ( .A(p_input[414]), .Z(n9171) );
  IV U17705 ( .A(p_input[415]), .Z(n9170) );
  XOR U17706 ( .A(n18111), .B(n18110), .Z(n18109) );
  AND U17707 ( .A(n9172), .B(n9173), .Z(n18110) );
  IV U17708 ( .A(p_input[412]), .Z(n9173) );
  IV U17709 ( .A(p_input[413]), .Z(n9172) );
  XOR U17710 ( .A(n18113), .B(n18112), .Z(n18111) );
  AND U17711 ( .A(n9174), .B(n9175), .Z(n18112) );
  IV U17712 ( .A(p_input[410]), .Z(n9175) );
  IV U17713 ( .A(p_input[411]), .Z(n9174) );
  XOR U17714 ( .A(n18115), .B(n18114), .Z(n18113) );
  AND U17715 ( .A(n9176), .B(n9177), .Z(n18114) );
  IV U17716 ( .A(p_input[408]), .Z(n9177) );
  IV U17717 ( .A(p_input[409]), .Z(n9176) );
  XOR U17718 ( .A(n18117), .B(n18116), .Z(n18115) );
  AND U17719 ( .A(n9178), .B(n9179), .Z(n18116) );
  IV U17720 ( .A(p_input[406]), .Z(n9179) );
  IV U17721 ( .A(p_input[407]), .Z(n9178) );
  XOR U17722 ( .A(n18119), .B(n18118), .Z(n18117) );
  AND U17723 ( .A(n9180), .B(n9181), .Z(n18118) );
  IV U17724 ( .A(p_input[404]), .Z(n9181) );
  IV U17725 ( .A(p_input[405]), .Z(n9180) );
  XOR U17726 ( .A(n18121), .B(n18120), .Z(n18119) );
  AND U17727 ( .A(n9182), .B(n9183), .Z(n18120) );
  IV U17728 ( .A(p_input[402]), .Z(n9183) );
  IV U17729 ( .A(p_input[403]), .Z(n9182) );
  XOR U17730 ( .A(n18123), .B(n18122), .Z(n18121) );
  AND U17731 ( .A(n9184), .B(n9185), .Z(n18122) );
  IV U17732 ( .A(p_input[400]), .Z(n9185) );
  IV U17733 ( .A(p_input[401]), .Z(n9184) );
  XOR U17734 ( .A(n18125), .B(n18124), .Z(n18123) );
  AND U17735 ( .A(n9186), .B(n9187), .Z(n18124) );
  IV U17736 ( .A(p_input[398]), .Z(n9187) );
  IV U17737 ( .A(p_input[399]), .Z(n9186) );
  XOR U17738 ( .A(n18127), .B(n18126), .Z(n18125) );
  AND U17739 ( .A(n9188), .B(n9189), .Z(n18126) );
  IV U17740 ( .A(p_input[396]), .Z(n9189) );
  IV U17741 ( .A(p_input[397]), .Z(n9188) );
  XOR U17742 ( .A(n18129), .B(n18128), .Z(n18127) );
  AND U17743 ( .A(n9190), .B(n9191), .Z(n18128) );
  IV U17744 ( .A(p_input[394]), .Z(n9191) );
  IV U17745 ( .A(p_input[395]), .Z(n9190) );
  XOR U17746 ( .A(n18131), .B(n18130), .Z(n18129) );
  AND U17747 ( .A(n9192), .B(n9193), .Z(n18130) );
  IV U17748 ( .A(p_input[392]), .Z(n9193) );
  IV U17749 ( .A(p_input[393]), .Z(n9192) );
  XOR U17750 ( .A(n18133), .B(n18132), .Z(n18131) );
  AND U17751 ( .A(n9194), .B(n9195), .Z(n18132) );
  IV U17752 ( .A(p_input[390]), .Z(n9195) );
  IV U17753 ( .A(p_input[391]), .Z(n9194) );
  XOR U17754 ( .A(n18135), .B(n18134), .Z(n18133) );
  AND U17755 ( .A(n9196), .B(n9197), .Z(n18134) );
  IV U17756 ( .A(p_input[388]), .Z(n9197) );
  IV U17757 ( .A(p_input[389]), .Z(n9196) );
  XOR U17758 ( .A(n18137), .B(n18136), .Z(n18135) );
  AND U17759 ( .A(n9198), .B(n9199), .Z(n18136) );
  IV U17760 ( .A(p_input[386]), .Z(n9199) );
  IV U17761 ( .A(p_input[387]), .Z(n9198) );
  XOR U17762 ( .A(n18139), .B(n18138), .Z(n18137) );
  AND U17763 ( .A(n9200), .B(n9201), .Z(n18138) );
  IV U17764 ( .A(p_input[384]), .Z(n9201) );
  IV U17765 ( .A(p_input[385]), .Z(n9200) );
  XOR U17766 ( .A(n18141), .B(n18140), .Z(n18139) );
  AND U17767 ( .A(n9202), .B(n9203), .Z(n18140) );
  IV U17768 ( .A(p_input[382]), .Z(n9203) );
  IV U17769 ( .A(p_input[383]), .Z(n9202) );
  XOR U17770 ( .A(n18143), .B(n18142), .Z(n18141) );
  AND U17771 ( .A(n9204), .B(n9205), .Z(n18142) );
  IV U17772 ( .A(p_input[380]), .Z(n9205) );
  IV U17773 ( .A(p_input[381]), .Z(n9204) );
  XOR U17774 ( .A(n18145), .B(n18144), .Z(n18143) );
  AND U17775 ( .A(n9206), .B(n9207), .Z(n18144) );
  IV U17776 ( .A(p_input[378]), .Z(n9207) );
  IV U17777 ( .A(p_input[379]), .Z(n9206) );
  XOR U17778 ( .A(n18147), .B(n18146), .Z(n18145) );
  AND U17779 ( .A(n9208), .B(n9209), .Z(n18146) );
  IV U17780 ( .A(p_input[376]), .Z(n9209) );
  IV U17781 ( .A(p_input[377]), .Z(n9208) );
  XOR U17782 ( .A(n18149), .B(n18148), .Z(n18147) );
  AND U17783 ( .A(n9210), .B(n9211), .Z(n18148) );
  IV U17784 ( .A(p_input[374]), .Z(n9211) );
  IV U17785 ( .A(p_input[375]), .Z(n9210) );
  XOR U17786 ( .A(n18151), .B(n18150), .Z(n18149) );
  AND U17787 ( .A(n9212), .B(n9213), .Z(n18150) );
  IV U17788 ( .A(p_input[372]), .Z(n9213) );
  IV U17789 ( .A(p_input[373]), .Z(n9212) );
  XOR U17790 ( .A(n18153), .B(n18152), .Z(n18151) );
  AND U17791 ( .A(n9214), .B(n9215), .Z(n18152) );
  IV U17792 ( .A(p_input[370]), .Z(n9215) );
  IV U17793 ( .A(p_input[371]), .Z(n9214) );
  XOR U17794 ( .A(n18155), .B(n18154), .Z(n18153) );
  AND U17795 ( .A(n9216), .B(n9217), .Z(n18154) );
  IV U17796 ( .A(p_input[368]), .Z(n9217) );
  IV U17797 ( .A(p_input[369]), .Z(n9216) );
  XOR U17798 ( .A(n18157), .B(n18156), .Z(n18155) );
  AND U17799 ( .A(n9218), .B(n9219), .Z(n18156) );
  IV U17800 ( .A(p_input[366]), .Z(n9219) );
  IV U17801 ( .A(p_input[367]), .Z(n9218) );
  XOR U17802 ( .A(n18159), .B(n18158), .Z(n18157) );
  AND U17803 ( .A(n9220), .B(n9221), .Z(n18158) );
  IV U17804 ( .A(p_input[364]), .Z(n9221) );
  IV U17805 ( .A(p_input[365]), .Z(n9220) );
  XOR U17806 ( .A(n18161), .B(n18160), .Z(n18159) );
  AND U17807 ( .A(n9222), .B(n9223), .Z(n18160) );
  IV U17808 ( .A(p_input[362]), .Z(n9223) );
  IV U17809 ( .A(p_input[363]), .Z(n9222) );
  XOR U17810 ( .A(n18163), .B(n18162), .Z(n18161) );
  AND U17811 ( .A(n9224), .B(n9225), .Z(n18162) );
  IV U17812 ( .A(p_input[360]), .Z(n9225) );
  IV U17813 ( .A(p_input[361]), .Z(n9224) );
  XOR U17814 ( .A(n18165), .B(n18164), .Z(n18163) );
  AND U17815 ( .A(n9226), .B(n9227), .Z(n18164) );
  IV U17816 ( .A(p_input[358]), .Z(n9227) );
  IV U17817 ( .A(p_input[359]), .Z(n9226) );
  XOR U17818 ( .A(n18167), .B(n18166), .Z(n18165) );
  AND U17819 ( .A(n9228), .B(n9229), .Z(n18166) );
  IV U17820 ( .A(p_input[356]), .Z(n9229) );
  IV U17821 ( .A(p_input[357]), .Z(n9228) );
  XOR U17822 ( .A(n18169), .B(n18168), .Z(n18167) );
  AND U17823 ( .A(n9230), .B(n9231), .Z(n18168) );
  IV U17824 ( .A(p_input[354]), .Z(n9231) );
  IV U17825 ( .A(p_input[355]), .Z(n9230) );
  XOR U17826 ( .A(n18171), .B(n18170), .Z(n18169) );
  AND U17827 ( .A(n9232), .B(n9233), .Z(n18170) );
  IV U17828 ( .A(p_input[352]), .Z(n9233) );
  IV U17829 ( .A(p_input[353]), .Z(n9232) );
  XOR U17830 ( .A(n18173), .B(n18172), .Z(n18171) );
  AND U17831 ( .A(n9234), .B(n9235), .Z(n18172) );
  IV U17832 ( .A(p_input[350]), .Z(n9235) );
  IV U17833 ( .A(p_input[351]), .Z(n9234) );
  XOR U17834 ( .A(n18175), .B(n18174), .Z(n18173) );
  AND U17835 ( .A(n9236), .B(n9237), .Z(n18174) );
  IV U17836 ( .A(p_input[348]), .Z(n9237) );
  IV U17837 ( .A(p_input[349]), .Z(n9236) );
  XOR U17838 ( .A(n18177), .B(n18176), .Z(n18175) );
  AND U17839 ( .A(n9238), .B(n9239), .Z(n18176) );
  IV U17840 ( .A(p_input[346]), .Z(n9239) );
  IV U17841 ( .A(p_input[347]), .Z(n9238) );
  XOR U17842 ( .A(n18179), .B(n18178), .Z(n18177) );
  AND U17843 ( .A(n9240), .B(n9241), .Z(n18178) );
  IV U17844 ( .A(p_input[344]), .Z(n9241) );
  IV U17845 ( .A(p_input[345]), .Z(n9240) );
  XOR U17846 ( .A(n18181), .B(n18180), .Z(n18179) );
  AND U17847 ( .A(n9242), .B(n9243), .Z(n18180) );
  IV U17848 ( .A(p_input[342]), .Z(n9243) );
  IV U17849 ( .A(p_input[343]), .Z(n9242) );
  XOR U17850 ( .A(n18183), .B(n18182), .Z(n18181) );
  AND U17851 ( .A(n9244), .B(n9245), .Z(n18182) );
  IV U17852 ( .A(p_input[340]), .Z(n9245) );
  IV U17853 ( .A(p_input[341]), .Z(n9244) );
  XOR U17854 ( .A(n18185), .B(n18184), .Z(n18183) );
  AND U17855 ( .A(n9246), .B(n9247), .Z(n18184) );
  IV U17856 ( .A(p_input[338]), .Z(n9247) );
  IV U17857 ( .A(p_input[339]), .Z(n9246) );
  XOR U17858 ( .A(n18187), .B(n18186), .Z(n18185) );
  AND U17859 ( .A(n9248), .B(n9249), .Z(n18186) );
  IV U17860 ( .A(p_input[336]), .Z(n9249) );
  IV U17861 ( .A(p_input[337]), .Z(n9248) );
  XOR U17862 ( .A(n18189), .B(n18188), .Z(n18187) );
  AND U17863 ( .A(n9250), .B(n9251), .Z(n18188) );
  IV U17864 ( .A(p_input[334]), .Z(n9251) );
  IV U17865 ( .A(p_input[335]), .Z(n9250) );
  XOR U17866 ( .A(n18191), .B(n18190), .Z(n18189) );
  AND U17867 ( .A(n9252), .B(n9253), .Z(n18190) );
  IV U17868 ( .A(p_input[332]), .Z(n9253) );
  IV U17869 ( .A(p_input[333]), .Z(n9252) );
  XOR U17870 ( .A(n18193), .B(n18192), .Z(n18191) );
  AND U17871 ( .A(n9254), .B(n9255), .Z(n18192) );
  IV U17872 ( .A(p_input[330]), .Z(n9255) );
  IV U17873 ( .A(p_input[331]), .Z(n9254) );
  XOR U17874 ( .A(n18195), .B(n18194), .Z(n18193) );
  AND U17875 ( .A(n9256), .B(n9257), .Z(n18194) );
  IV U17876 ( .A(p_input[328]), .Z(n9257) );
  IV U17877 ( .A(p_input[329]), .Z(n9256) );
  XOR U17878 ( .A(n18197), .B(n18196), .Z(n18195) );
  AND U17879 ( .A(n9258), .B(n9259), .Z(n18196) );
  IV U17880 ( .A(p_input[326]), .Z(n9259) );
  IV U17881 ( .A(p_input[327]), .Z(n9258) );
  XOR U17882 ( .A(n18199), .B(n18198), .Z(n18197) );
  AND U17883 ( .A(n9260), .B(n9261), .Z(n18198) );
  IV U17884 ( .A(p_input[324]), .Z(n9261) );
  IV U17885 ( .A(p_input[325]), .Z(n9260) );
  XOR U17886 ( .A(n18201), .B(n18200), .Z(n18199) );
  AND U17887 ( .A(n9262), .B(n9263), .Z(n18200) );
  IV U17888 ( .A(p_input[322]), .Z(n9263) );
  IV U17889 ( .A(p_input[323]), .Z(n9262) );
  XOR U17890 ( .A(n18203), .B(n18202), .Z(n18201) );
  AND U17891 ( .A(n9264), .B(n9265), .Z(n18202) );
  IV U17892 ( .A(p_input[320]), .Z(n9265) );
  IV U17893 ( .A(p_input[321]), .Z(n9264) );
  XOR U17894 ( .A(n18205), .B(n18204), .Z(n18203) );
  AND U17895 ( .A(n9266), .B(n9267), .Z(n18204) );
  IV U17896 ( .A(p_input[318]), .Z(n9267) );
  IV U17897 ( .A(p_input[319]), .Z(n9266) );
  XOR U17898 ( .A(n18207), .B(n18206), .Z(n18205) );
  AND U17899 ( .A(n9268), .B(n9269), .Z(n18206) );
  IV U17900 ( .A(p_input[316]), .Z(n9269) );
  IV U17901 ( .A(p_input[317]), .Z(n9268) );
  XOR U17902 ( .A(n18209), .B(n18208), .Z(n18207) );
  AND U17903 ( .A(n9270), .B(n9271), .Z(n18208) );
  IV U17904 ( .A(p_input[314]), .Z(n9271) );
  IV U17905 ( .A(p_input[315]), .Z(n9270) );
  XOR U17906 ( .A(n18211), .B(n18210), .Z(n18209) );
  AND U17907 ( .A(n9272), .B(n9273), .Z(n18210) );
  IV U17908 ( .A(p_input[312]), .Z(n9273) );
  IV U17909 ( .A(p_input[313]), .Z(n9272) );
  XOR U17910 ( .A(n18213), .B(n18212), .Z(n18211) );
  AND U17911 ( .A(n9274), .B(n9275), .Z(n18212) );
  IV U17912 ( .A(p_input[310]), .Z(n9275) );
  IV U17913 ( .A(p_input[311]), .Z(n9274) );
  XOR U17914 ( .A(n18215), .B(n18214), .Z(n18213) );
  AND U17915 ( .A(n9276), .B(n9277), .Z(n18214) );
  IV U17916 ( .A(p_input[308]), .Z(n9277) );
  IV U17917 ( .A(p_input[309]), .Z(n9276) );
  XOR U17918 ( .A(n18217), .B(n18216), .Z(n18215) );
  AND U17919 ( .A(n9278), .B(n9279), .Z(n18216) );
  IV U17920 ( .A(p_input[306]), .Z(n9279) );
  IV U17921 ( .A(p_input[307]), .Z(n9278) );
  XOR U17922 ( .A(n18219), .B(n18218), .Z(n18217) );
  AND U17923 ( .A(n9280), .B(n9281), .Z(n18218) );
  IV U17924 ( .A(p_input[304]), .Z(n9281) );
  IV U17925 ( .A(p_input[305]), .Z(n9280) );
  XOR U17926 ( .A(n18221), .B(n18220), .Z(n18219) );
  AND U17927 ( .A(n9282), .B(n9283), .Z(n18220) );
  IV U17928 ( .A(p_input[302]), .Z(n9283) );
  IV U17929 ( .A(p_input[303]), .Z(n9282) );
  XOR U17930 ( .A(n18223), .B(n18222), .Z(n18221) );
  AND U17931 ( .A(n9284), .B(n9285), .Z(n18222) );
  IV U17932 ( .A(p_input[300]), .Z(n9285) );
  IV U17933 ( .A(p_input[301]), .Z(n9284) );
  XOR U17934 ( .A(n18225), .B(n18224), .Z(n18223) );
  AND U17935 ( .A(n9286), .B(n9287), .Z(n18224) );
  IV U17936 ( .A(p_input[298]), .Z(n9287) );
  IV U17937 ( .A(p_input[299]), .Z(n9286) );
  XOR U17938 ( .A(n18227), .B(n18226), .Z(n18225) );
  AND U17939 ( .A(n9288), .B(n9289), .Z(n18226) );
  IV U17940 ( .A(p_input[296]), .Z(n9289) );
  IV U17941 ( .A(p_input[297]), .Z(n9288) );
  XOR U17942 ( .A(n18229), .B(n18228), .Z(n18227) );
  AND U17943 ( .A(n9290), .B(n9291), .Z(n18228) );
  IV U17944 ( .A(p_input[294]), .Z(n9291) );
  IV U17945 ( .A(p_input[295]), .Z(n9290) );
  XOR U17946 ( .A(n18231), .B(n18230), .Z(n18229) );
  AND U17947 ( .A(n9292), .B(n9293), .Z(n18230) );
  IV U17948 ( .A(p_input[292]), .Z(n9293) );
  IV U17949 ( .A(p_input[293]), .Z(n9292) );
  XOR U17950 ( .A(n18233), .B(n18232), .Z(n18231) );
  AND U17951 ( .A(n9294), .B(n9295), .Z(n18232) );
  IV U17952 ( .A(p_input[290]), .Z(n9295) );
  IV U17953 ( .A(p_input[291]), .Z(n9294) );
  XOR U17954 ( .A(n18235), .B(n18234), .Z(n18233) );
  AND U17955 ( .A(n9296), .B(n9297), .Z(n18234) );
  IV U17956 ( .A(p_input[288]), .Z(n9297) );
  IV U17957 ( .A(p_input[289]), .Z(n9296) );
  XOR U17958 ( .A(n18237), .B(n18236), .Z(n18235) );
  AND U17959 ( .A(n9298), .B(n9299), .Z(n18236) );
  IV U17960 ( .A(p_input[286]), .Z(n9299) );
  IV U17961 ( .A(p_input[287]), .Z(n9298) );
  XOR U17962 ( .A(n18239), .B(n18238), .Z(n18237) );
  AND U17963 ( .A(n9300), .B(n9301), .Z(n18238) );
  IV U17964 ( .A(p_input[284]), .Z(n9301) );
  IV U17965 ( .A(p_input[285]), .Z(n9300) );
  XOR U17966 ( .A(n18241), .B(n18240), .Z(n18239) );
  AND U17967 ( .A(n9302), .B(n9303), .Z(n18240) );
  IV U17968 ( .A(p_input[282]), .Z(n9303) );
  IV U17969 ( .A(p_input[283]), .Z(n9302) );
  XOR U17970 ( .A(n18243), .B(n18242), .Z(n18241) );
  AND U17971 ( .A(n9304), .B(n9305), .Z(n18242) );
  IV U17972 ( .A(p_input[280]), .Z(n9305) );
  IV U17973 ( .A(p_input[281]), .Z(n9304) );
  XOR U17974 ( .A(n18245), .B(n18244), .Z(n18243) );
  AND U17975 ( .A(n9306), .B(n9307), .Z(n18244) );
  IV U17976 ( .A(p_input[278]), .Z(n9307) );
  IV U17977 ( .A(p_input[279]), .Z(n9306) );
  XOR U17978 ( .A(n18247), .B(n18246), .Z(n18245) );
  AND U17979 ( .A(n9308), .B(n9309), .Z(n18246) );
  IV U17980 ( .A(p_input[276]), .Z(n9309) );
  IV U17981 ( .A(p_input[277]), .Z(n9308) );
  XOR U17982 ( .A(n18249), .B(n18248), .Z(n18247) );
  AND U17983 ( .A(n9310), .B(n9311), .Z(n18248) );
  IV U17984 ( .A(p_input[274]), .Z(n9311) );
  IV U17985 ( .A(p_input[275]), .Z(n9310) );
  XOR U17986 ( .A(n18251), .B(n18250), .Z(n18249) );
  AND U17987 ( .A(n9312), .B(n9313), .Z(n18250) );
  IV U17988 ( .A(p_input[272]), .Z(n9313) );
  IV U17989 ( .A(p_input[273]), .Z(n9312) );
  XOR U17990 ( .A(n18253), .B(n18252), .Z(n18251) );
  AND U17991 ( .A(n9314), .B(n9315), .Z(n18252) );
  IV U17992 ( .A(p_input[270]), .Z(n9315) );
  IV U17993 ( .A(p_input[271]), .Z(n9314) );
  XOR U17994 ( .A(n18255), .B(n18254), .Z(n18253) );
  AND U17995 ( .A(n9316), .B(n9317), .Z(n18254) );
  IV U17996 ( .A(p_input[268]), .Z(n9317) );
  IV U17997 ( .A(p_input[269]), .Z(n9316) );
  XOR U17998 ( .A(n18257), .B(n18256), .Z(n18255) );
  AND U17999 ( .A(n9318), .B(n9319), .Z(n18256) );
  IV U18000 ( .A(p_input[266]), .Z(n9319) );
  IV U18001 ( .A(p_input[267]), .Z(n9318) );
  XOR U18002 ( .A(n18259), .B(n18258), .Z(n18257) );
  AND U18003 ( .A(n9320), .B(n9321), .Z(n18258) );
  IV U18004 ( .A(p_input[264]), .Z(n9321) );
  IV U18005 ( .A(p_input[265]), .Z(n9320) );
  XOR U18006 ( .A(n18261), .B(n18260), .Z(n18259) );
  AND U18007 ( .A(n9322), .B(n9323), .Z(n18260) );
  IV U18008 ( .A(p_input[262]), .Z(n9323) );
  IV U18009 ( .A(p_input[263]), .Z(n9322) );
  XOR U18010 ( .A(n18263), .B(n18262), .Z(n18261) );
  AND U18011 ( .A(n9324), .B(n9325), .Z(n18262) );
  IV U18012 ( .A(p_input[260]), .Z(n9325) );
  IV U18013 ( .A(p_input[261]), .Z(n9324) );
  XOR U18014 ( .A(n18265), .B(n18264), .Z(n18263) );
  AND U18015 ( .A(n9326), .B(n9327), .Z(n18264) );
  IV U18016 ( .A(p_input[258]), .Z(n9327) );
  IV U18017 ( .A(p_input[259]), .Z(n9326) );
  XOR U18018 ( .A(n18267), .B(n18266), .Z(n18265) );
  AND U18019 ( .A(n9328), .B(n9329), .Z(n18266) );
  IV U18020 ( .A(p_input[256]), .Z(n9329) );
  IV U18021 ( .A(p_input[257]), .Z(n9328) );
  XOR U18022 ( .A(n18269), .B(n18268), .Z(n18267) );
  AND U18023 ( .A(n9330), .B(n9331), .Z(n18268) );
  IV U18024 ( .A(p_input[254]), .Z(n9331) );
  IV U18025 ( .A(p_input[255]), .Z(n9330) );
  XOR U18026 ( .A(n18273), .B(n18272), .Z(n18269) );
  AND U18027 ( .A(n9332), .B(n9333), .Z(n18272) );
  IV U18028 ( .A(p_input[252]), .Z(n9333) );
  IV U18029 ( .A(p_input[253]), .Z(n9332) );
  XOR U18030 ( .A(n18275), .B(n18274), .Z(n18273) );
  AND U18031 ( .A(n9334), .B(n9335), .Z(n18274) );
  IV U18032 ( .A(p_input[250]), .Z(n9335) );
  IV U18033 ( .A(p_input[251]), .Z(n9334) );
  XOR U18034 ( .A(n18277), .B(n18276), .Z(n18275) );
  AND U18035 ( .A(n9336), .B(n9337), .Z(n18276) );
  IV U18036 ( .A(p_input[248]), .Z(n9337) );
  IV U18037 ( .A(p_input[249]), .Z(n9336) );
  XOR U18038 ( .A(n18279), .B(n18278), .Z(n18277) );
  AND U18039 ( .A(n9338), .B(n9339), .Z(n18278) );
  IV U18040 ( .A(p_input[246]), .Z(n9339) );
  IV U18041 ( .A(p_input[247]), .Z(n9338) );
  XOR U18042 ( .A(n18281), .B(n18280), .Z(n18279) );
  AND U18043 ( .A(n9340), .B(n9341), .Z(n18280) );
  IV U18044 ( .A(p_input[244]), .Z(n9341) );
  IV U18045 ( .A(p_input[245]), .Z(n9340) );
  XOR U18046 ( .A(n18283), .B(n18282), .Z(n18281) );
  AND U18047 ( .A(n9342), .B(n9343), .Z(n18282) );
  IV U18048 ( .A(p_input[242]), .Z(n9343) );
  IV U18049 ( .A(p_input[243]), .Z(n9342) );
  XOR U18050 ( .A(n18285), .B(n18284), .Z(n18283) );
  AND U18051 ( .A(n9344), .B(n9345), .Z(n18284) );
  IV U18052 ( .A(p_input[240]), .Z(n9345) );
  IV U18053 ( .A(p_input[241]), .Z(n9344) );
  XOR U18054 ( .A(n18287), .B(n18286), .Z(n18285) );
  AND U18055 ( .A(n9346), .B(n9347), .Z(n18286) );
  IV U18056 ( .A(p_input[238]), .Z(n9347) );
  IV U18057 ( .A(p_input[239]), .Z(n9346) );
  XOR U18058 ( .A(n18289), .B(n18288), .Z(n18287) );
  AND U18059 ( .A(n9348), .B(n9349), .Z(n18288) );
  IV U18060 ( .A(p_input[236]), .Z(n9349) );
  IV U18061 ( .A(p_input[237]), .Z(n9348) );
  XOR U18062 ( .A(n18291), .B(n18290), .Z(n18289) );
  AND U18063 ( .A(n9350), .B(n9351), .Z(n18290) );
  IV U18064 ( .A(p_input[234]), .Z(n9351) );
  IV U18065 ( .A(p_input[235]), .Z(n9350) );
  XOR U18066 ( .A(n18293), .B(n18292), .Z(n18291) );
  AND U18067 ( .A(n9352), .B(n9353), .Z(n18292) );
  IV U18068 ( .A(p_input[232]), .Z(n9353) );
  IV U18069 ( .A(p_input[233]), .Z(n9352) );
  XOR U18070 ( .A(n18295), .B(n18294), .Z(n18293) );
  AND U18071 ( .A(n9354), .B(n9355), .Z(n18294) );
  IV U18072 ( .A(p_input[230]), .Z(n9355) );
  IV U18073 ( .A(p_input[231]), .Z(n9354) );
  XOR U18074 ( .A(n18297), .B(n18296), .Z(n18295) );
  AND U18075 ( .A(n9356), .B(n9357), .Z(n18296) );
  IV U18076 ( .A(p_input[228]), .Z(n9357) );
  IV U18077 ( .A(p_input[229]), .Z(n9356) );
  XOR U18078 ( .A(n18299), .B(n18298), .Z(n18297) );
  AND U18079 ( .A(n9358), .B(n9359), .Z(n18298) );
  IV U18080 ( .A(p_input[226]), .Z(n9359) );
  IV U18081 ( .A(p_input[227]), .Z(n9358) );
  XOR U18082 ( .A(n18301), .B(n18300), .Z(n18299) );
  AND U18083 ( .A(n9360), .B(n9361), .Z(n18300) );
  IV U18084 ( .A(p_input[224]), .Z(n9361) );
  IV U18085 ( .A(p_input[225]), .Z(n9360) );
  XOR U18086 ( .A(n18303), .B(n18302), .Z(n18301) );
  AND U18087 ( .A(n9362), .B(n9363), .Z(n18302) );
  IV U18088 ( .A(p_input[222]), .Z(n9363) );
  IV U18089 ( .A(p_input[223]), .Z(n9362) );
  XOR U18090 ( .A(n18305), .B(n18304), .Z(n18303) );
  AND U18091 ( .A(n9364), .B(n9365), .Z(n18304) );
  IV U18092 ( .A(p_input[220]), .Z(n9365) );
  IV U18093 ( .A(p_input[221]), .Z(n9364) );
  XOR U18094 ( .A(n18307), .B(n18306), .Z(n18305) );
  AND U18095 ( .A(n9366), .B(n9367), .Z(n18306) );
  IV U18096 ( .A(p_input[218]), .Z(n9367) );
  IV U18097 ( .A(p_input[219]), .Z(n9366) );
  XOR U18098 ( .A(n18309), .B(n18308), .Z(n18307) );
  AND U18099 ( .A(n9368), .B(n9369), .Z(n18308) );
  IV U18100 ( .A(p_input[216]), .Z(n9369) );
  IV U18101 ( .A(p_input[217]), .Z(n9368) );
  XOR U18102 ( .A(n18311), .B(n18310), .Z(n18309) );
  AND U18103 ( .A(n9370), .B(n9371), .Z(n18310) );
  IV U18104 ( .A(p_input[214]), .Z(n9371) );
  IV U18105 ( .A(p_input[215]), .Z(n9370) );
  XOR U18106 ( .A(n18313), .B(n18312), .Z(n18311) );
  AND U18107 ( .A(n9372), .B(n9373), .Z(n18312) );
  IV U18108 ( .A(p_input[212]), .Z(n9373) );
  IV U18109 ( .A(p_input[213]), .Z(n9372) );
  XOR U18110 ( .A(n18315), .B(n18314), .Z(n18313) );
  AND U18111 ( .A(n9374), .B(n9375), .Z(n18314) );
  IV U18112 ( .A(p_input[210]), .Z(n9375) );
  IV U18113 ( .A(p_input[211]), .Z(n9374) );
  XOR U18114 ( .A(n18317), .B(n18316), .Z(n18315) );
  AND U18115 ( .A(n9376), .B(n9377), .Z(n18316) );
  IV U18116 ( .A(p_input[208]), .Z(n9377) );
  IV U18117 ( .A(p_input[209]), .Z(n9376) );
  XOR U18118 ( .A(n18319), .B(n18318), .Z(n18317) );
  AND U18119 ( .A(n9378), .B(n9379), .Z(n18318) );
  IV U18120 ( .A(p_input[206]), .Z(n9379) );
  IV U18121 ( .A(p_input[207]), .Z(n9378) );
  XOR U18122 ( .A(n18321), .B(n18320), .Z(n18319) );
  AND U18123 ( .A(n9380), .B(n9381), .Z(n18320) );
  IV U18124 ( .A(p_input[204]), .Z(n9381) );
  IV U18125 ( .A(p_input[205]), .Z(n9380) );
  XOR U18126 ( .A(n18323), .B(n18322), .Z(n18321) );
  AND U18127 ( .A(n9382), .B(n9383), .Z(n18322) );
  IV U18128 ( .A(p_input[202]), .Z(n9383) );
  IV U18129 ( .A(p_input[203]), .Z(n9382) );
  XOR U18130 ( .A(n18325), .B(n18324), .Z(n18323) );
  AND U18131 ( .A(n9384), .B(n9385), .Z(n18324) );
  IV U18132 ( .A(p_input[200]), .Z(n9385) );
  IV U18133 ( .A(p_input[201]), .Z(n9384) );
  XOR U18134 ( .A(n18327), .B(n18326), .Z(n18325) );
  AND U18135 ( .A(n9386), .B(n9387), .Z(n18326) );
  IV U18136 ( .A(p_input[198]), .Z(n9387) );
  IV U18137 ( .A(p_input[199]), .Z(n9386) );
  XOR U18138 ( .A(n18329), .B(n18328), .Z(n18327) );
  AND U18139 ( .A(n9388), .B(n9389), .Z(n18328) );
  IV U18140 ( .A(p_input[196]), .Z(n9389) );
  IV U18141 ( .A(p_input[197]), .Z(n9388) );
  XOR U18142 ( .A(n18331), .B(n18330), .Z(n18329) );
  AND U18143 ( .A(n9390), .B(n9391), .Z(n18330) );
  IV U18144 ( .A(p_input[194]), .Z(n9391) );
  IV U18145 ( .A(p_input[195]), .Z(n9390) );
  XOR U18146 ( .A(n18333), .B(n18332), .Z(n18331) );
  AND U18147 ( .A(n9392), .B(n9393), .Z(n18332) );
  IV U18148 ( .A(p_input[192]), .Z(n9393) );
  IV U18149 ( .A(p_input[193]), .Z(n9392) );
  XOR U18150 ( .A(n18335), .B(n18334), .Z(n18333) );
  AND U18151 ( .A(n9394), .B(n9395), .Z(n18334) );
  IV U18152 ( .A(p_input[190]), .Z(n9395) );
  IV U18153 ( .A(p_input[191]), .Z(n9394) );
  XOR U18154 ( .A(n18337), .B(n18336), .Z(n18335) );
  AND U18155 ( .A(n9396), .B(n9397), .Z(n18336) );
  IV U18156 ( .A(p_input[188]), .Z(n9397) );
  IV U18157 ( .A(p_input[189]), .Z(n9396) );
  XOR U18158 ( .A(n18339), .B(n18338), .Z(n18337) );
  AND U18159 ( .A(n9398), .B(n9399), .Z(n18338) );
  IV U18160 ( .A(p_input[186]), .Z(n9399) );
  IV U18161 ( .A(p_input[187]), .Z(n9398) );
  XOR U18162 ( .A(n18341), .B(n18340), .Z(n18339) );
  AND U18163 ( .A(n9400), .B(n9401), .Z(n18340) );
  IV U18164 ( .A(p_input[184]), .Z(n9401) );
  IV U18165 ( .A(p_input[185]), .Z(n9400) );
  XOR U18166 ( .A(n18343), .B(n18342), .Z(n18341) );
  AND U18167 ( .A(n9402), .B(n9403), .Z(n18342) );
  IV U18168 ( .A(p_input[182]), .Z(n9403) );
  IV U18169 ( .A(p_input[183]), .Z(n9402) );
  XOR U18170 ( .A(n18345), .B(n18344), .Z(n18343) );
  AND U18171 ( .A(n9404), .B(n9405), .Z(n18344) );
  IV U18172 ( .A(p_input[180]), .Z(n9405) );
  IV U18173 ( .A(p_input[181]), .Z(n9404) );
  XOR U18174 ( .A(n18347), .B(n18346), .Z(n18345) );
  AND U18175 ( .A(n9406), .B(n9407), .Z(n18346) );
  IV U18176 ( .A(p_input[178]), .Z(n9407) );
  IV U18177 ( .A(p_input[179]), .Z(n9406) );
  XOR U18178 ( .A(n18349), .B(n18348), .Z(n18347) );
  AND U18179 ( .A(n9408), .B(n9409), .Z(n18348) );
  IV U18180 ( .A(p_input[176]), .Z(n9409) );
  IV U18181 ( .A(p_input[177]), .Z(n9408) );
  XOR U18182 ( .A(n18351), .B(n18350), .Z(n18349) );
  AND U18183 ( .A(n9410), .B(n9411), .Z(n18350) );
  IV U18184 ( .A(p_input[174]), .Z(n9411) );
  IV U18185 ( .A(p_input[175]), .Z(n9410) );
  XOR U18186 ( .A(n18353), .B(n18352), .Z(n18351) );
  AND U18187 ( .A(n9412), .B(n9413), .Z(n18352) );
  IV U18188 ( .A(p_input[172]), .Z(n9413) );
  IV U18189 ( .A(p_input[173]), .Z(n9412) );
  XOR U18190 ( .A(n18355), .B(n18354), .Z(n18353) );
  AND U18191 ( .A(n9414), .B(n9415), .Z(n18354) );
  IV U18192 ( .A(p_input[170]), .Z(n9415) );
  IV U18193 ( .A(p_input[171]), .Z(n9414) );
  XOR U18194 ( .A(n18357), .B(n18356), .Z(n18355) );
  AND U18195 ( .A(n9416), .B(n9417), .Z(n18356) );
  IV U18196 ( .A(p_input[168]), .Z(n9417) );
  IV U18197 ( .A(p_input[169]), .Z(n9416) );
  XOR U18198 ( .A(n18359), .B(n18358), .Z(n18357) );
  AND U18199 ( .A(n9418), .B(n9419), .Z(n18358) );
  IV U18200 ( .A(p_input[166]), .Z(n9419) );
  IV U18201 ( .A(p_input[167]), .Z(n9418) );
  XOR U18202 ( .A(n18361), .B(n18360), .Z(n18359) );
  AND U18203 ( .A(n9420), .B(n9421), .Z(n18360) );
  IV U18204 ( .A(p_input[164]), .Z(n9421) );
  IV U18205 ( .A(p_input[165]), .Z(n9420) );
  XOR U18206 ( .A(n18363), .B(n18362), .Z(n18361) );
  AND U18207 ( .A(n9422), .B(n9423), .Z(n18362) );
  IV U18208 ( .A(p_input[162]), .Z(n9423) );
  IV U18209 ( .A(p_input[163]), .Z(n9422) );
  XOR U18210 ( .A(n18365), .B(n18364), .Z(n18363) );
  AND U18211 ( .A(n9424), .B(n9425), .Z(n18364) );
  IV U18212 ( .A(p_input[160]), .Z(n9425) );
  IV U18213 ( .A(p_input[161]), .Z(n9424) );
  XOR U18214 ( .A(n18367), .B(n18366), .Z(n18365) );
  AND U18215 ( .A(n9426), .B(n9427), .Z(n18366) );
  IV U18216 ( .A(p_input[158]), .Z(n9427) );
  IV U18217 ( .A(p_input[159]), .Z(n9426) );
  XOR U18218 ( .A(n18369), .B(n18368), .Z(n18367) );
  AND U18219 ( .A(n9428), .B(n9429), .Z(n18368) );
  IV U18220 ( .A(p_input[156]), .Z(n9429) );
  IV U18221 ( .A(p_input[157]), .Z(n9428) );
  XOR U18222 ( .A(n18371), .B(n18370), .Z(n18369) );
  AND U18223 ( .A(n9430), .B(n9431), .Z(n18370) );
  IV U18224 ( .A(p_input[154]), .Z(n9431) );
  IV U18225 ( .A(p_input[155]), .Z(n9430) );
  XOR U18226 ( .A(n18373), .B(n18372), .Z(n18371) );
  AND U18227 ( .A(n9432), .B(n9433), .Z(n18372) );
  IV U18228 ( .A(p_input[152]), .Z(n9433) );
  IV U18229 ( .A(p_input[153]), .Z(n9432) );
  XOR U18230 ( .A(n18375), .B(n18374), .Z(n18373) );
  AND U18231 ( .A(n9434), .B(n9435), .Z(n18374) );
  IV U18232 ( .A(p_input[150]), .Z(n9435) );
  IV U18233 ( .A(p_input[151]), .Z(n9434) );
  XOR U18234 ( .A(n18377), .B(n18376), .Z(n18375) );
  AND U18235 ( .A(n9436), .B(n9437), .Z(n18376) );
  IV U18236 ( .A(p_input[148]), .Z(n9437) );
  IV U18237 ( .A(p_input[149]), .Z(n9436) );
  XOR U18238 ( .A(n18379), .B(n18378), .Z(n18377) );
  AND U18239 ( .A(n9438), .B(n9439), .Z(n18378) );
  IV U18240 ( .A(p_input[146]), .Z(n9439) );
  IV U18241 ( .A(p_input[147]), .Z(n9438) );
  XOR U18242 ( .A(n18381), .B(n18380), .Z(n18379) );
  AND U18243 ( .A(n9440), .B(n9441), .Z(n18380) );
  IV U18244 ( .A(p_input[144]), .Z(n9441) );
  IV U18245 ( .A(p_input[145]), .Z(n9440) );
  XOR U18246 ( .A(n18383), .B(n18382), .Z(n18381) );
  AND U18247 ( .A(n9442), .B(n9443), .Z(n18382) );
  IV U18248 ( .A(p_input[142]), .Z(n9443) );
  IV U18249 ( .A(p_input[143]), .Z(n9442) );
  XOR U18250 ( .A(n18385), .B(n18384), .Z(n18383) );
  AND U18251 ( .A(n9444), .B(n9445), .Z(n18384) );
  IV U18252 ( .A(p_input[140]), .Z(n9445) );
  IV U18253 ( .A(p_input[141]), .Z(n9444) );
  XOR U18254 ( .A(n18387), .B(n18386), .Z(n18385) );
  AND U18255 ( .A(n9446), .B(n9447), .Z(n18386) );
  IV U18256 ( .A(p_input[138]), .Z(n9447) );
  IV U18257 ( .A(p_input[139]), .Z(n9446) );
  XOR U18258 ( .A(n18389), .B(n18388), .Z(n18387) );
  AND U18259 ( .A(n9448), .B(n9449), .Z(n18388) );
  IV U18260 ( .A(p_input[136]), .Z(n9449) );
  IV U18261 ( .A(p_input[137]), .Z(n9448) );
  XOR U18262 ( .A(n18391), .B(n18390), .Z(n18389) );
  AND U18263 ( .A(n9450), .B(n9451), .Z(n18390) );
  IV U18264 ( .A(p_input[134]), .Z(n9451) );
  IV U18265 ( .A(p_input[135]), .Z(n9450) );
  XOR U18266 ( .A(n18393), .B(n18392), .Z(n18391) );
  AND U18267 ( .A(n9452), .B(n9453), .Z(n18392) );
  IV U18268 ( .A(p_input[132]), .Z(n9453) );
  IV U18269 ( .A(p_input[133]), .Z(n9452) );
  XOR U18270 ( .A(n18395), .B(n18394), .Z(n18393) );
  AND U18271 ( .A(n9454), .B(n9455), .Z(n18394) );
  IV U18272 ( .A(p_input[130]), .Z(n9455) );
  IV U18273 ( .A(p_input[131]), .Z(n9454) );
  XOR U18274 ( .A(n18397), .B(n18396), .Z(n18395) );
  AND U18275 ( .A(n9456), .B(n9457), .Z(n18396) );
  IV U18276 ( .A(p_input[128]), .Z(n9457) );
  IV U18277 ( .A(p_input[129]), .Z(n9456) );
  XOR U18278 ( .A(n18399), .B(n18398), .Z(n18397) );
  AND U18279 ( .A(n9458), .B(n9459), .Z(n18398) );
  IV U18280 ( .A(p_input[126]), .Z(n9459) );
  IV U18281 ( .A(p_input[127]), .Z(n9458) );
  XOR U18282 ( .A(n18401), .B(n18400), .Z(n18399) );
  AND U18283 ( .A(n9460), .B(n9461), .Z(n18400) );
  IV U18284 ( .A(p_input[124]), .Z(n9461) );
  IV U18285 ( .A(p_input[125]), .Z(n9460) );
  XOR U18286 ( .A(n18403), .B(n18402), .Z(n18401) );
  AND U18287 ( .A(n9462), .B(n9463), .Z(n18402) );
  IV U18288 ( .A(p_input[122]), .Z(n9463) );
  IV U18289 ( .A(p_input[123]), .Z(n9462) );
  XOR U18290 ( .A(n18405), .B(n18404), .Z(n18403) );
  AND U18291 ( .A(n9464), .B(n9465), .Z(n18404) );
  IV U18292 ( .A(p_input[120]), .Z(n9465) );
  IV U18293 ( .A(p_input[121]), .Z(n9464) );
  XOR U18294 ( .A(n18407), .B(n18406), .Z(n18405) );
  AND U18295 ( .A(n9466), .B(n9467), .Z(n18406) );
  IV U18296 ( .A(p_input[118]), .Z(n9467) );
  IV U18297 ( .A(p_input[119]), .Z(n9466) );
  XOR U18298 ( .A(n18409), .B(n18408), .Z(n18407) );
  AND U18299 ( .A(n9468), .B(n9469), .Z(n18408) );
  IV U18300 ( .A(p_input[116]), .Z(n9469) );
  IV U18301 ( .A(p_input[117]), .Z(n9468) );
  XOR U18302 ( .A(n18411), .B(n18410), .Z(n18409) );
  AND U18303 ( .A(n9470), .B(n9471), .Z(n18410) );
  IV U18304 ( .A(p_input[114]), .Z(n9471) );
  IV U18305 ( .A(p_input[115]), .Z(n9470) );
  XOR U18306 ( .A(n18413), .B(n18412), .Z(n18411) );
  AND U18307 ( .A(n9472), .B(n9473), .Z(n18412) );
  IV U18308 ( .A(p_input[112]), .Z(n9473) );
  IV U18309 ( .A(p_input[113]), .Z(n9472) );
  XOR U18310 ( .A(n18415), .B(n18414), .Z(n18413) );
  AND U18311 ( .A(n9474), .B(n9475), .Z(n18414) );
  IV U18312 ( .A(p_input[110]), .Z(n9475) );
  IV U18313 ( .A(p_input[111]), .Z(n9474) );
  XOR U18314 ( .A(n18417), .B(n18416), .Z(n18415) );
  AND U18315 ( .A(n9476), .B(n9477), .Z(n18416) );
  IV U18316 ( .A(p_input[108]), .Z(n9477) );
  IV U18317 ( .A(p_input[109]), .Z(n9476) );
  XOR U18318 ( .A(n18419), .B(n18418), .Z(n18417) );
  AND U18319 ( .A(n9478), .B(n9479), .Z(n18418) );
  IV U18320 ( .A(p_input[106]), .Z(n9479) );
  IV U18321 ( .A(p_input[107]), .Z(n9478) );
  XOR U18322 ( .A(n18421), .B(n18420), .Z(n18419) );
  AND U18323 ( .A(n9480), .B(n9481), .Z(n18420) );
  IV U18324 ( .A(p_input[104]), .Z(n9481) );
  IV U18325 ( .A(p_input[105]), .Z(n9480) );
  XOR U18326 ( .A(n18423), .B(n18422), .Z(n18421) );
  AND U18327 ( .A(n9482), .B(n9483), .Z(n18422) );
  IV U18328 ( .A(p_input[102]), .Z(n9483) );
  IV U18329 ( .A(p_input[103]), .Z(n9482) );
  XOR U18330 ( .A(n18425), .B(n18424), .Z(n18423) );
  AND U18331 ( .A(n9484), .B(n9485), .Z(n18424) );
  IV U18332 ( .A(p_input[100]), .Z(n9485) );
  IV U18333 ( .A(p_input[101]), .Z(n9484) );
  XOR U18334 ( .A(n18427), .B(n18426), .Z(n18425) );
  AND U18335 ( .A(n9486), .B(n9487), .Z(n18426) );
  IV U18336 ( .A(p_input[98]), .Z(n9487) );
  IV U18337 ( .A(p_input[99]), .Z(n9486) );
  XOR U18338 ( .A(n18429), .B(n18428), .Z(n18427) );
  AND U18339 ( .A(n9488), .B(n9489), .Z(n18428) );
  IV U18340 ( .A(p_input[96]), .Z(n9489) );
  IV U18341 ( .A(p_input[97]), .Z(n9488) );
  XOR U18342 ( .A(n18431), .B(n18430), .Z(n18429) );
  AND U18343 ( .A(n9490), .B(n9491), .Z(n18430) );
  IV U18344 ( .A(p_input[94]), .Z(n9491) );
  IV U18345 ( .A(p_input[95]), .Z(n9490) );
  XOR U18346 ( .A(n18433), .B(n18432), .Z(n18431) );
  AND U18347 ( .A(n9492), .B(n9493), .Z(n18432) );
  IV U18348 ( .A(p_input[92]), .Z(n9493) );
  IV U18349 ( .A(p_input[93]), .Z(n9492) );
  XOR U18350 ( .A(n18435), .B(n18434), .Z(n18433) );
  AND U18351 ( .A(n9494), .B(n9495), .Z(n18434) );
  IV U18352 ( .A(p_input[90]), .Z(n9495) );
  IV U18353 ( .A(p_input[91]), .Z(n9494) );
  XOR U18354 ( .A(n18437), .B(n18436), .Z(n18435) );
  AND U18355 ( .A(n9496), .B(n9497), .Z(n18436) );
  IV U18356 ( .A(p_input[88]), .Z(n9497) );
  IV U18357 ( .A(p_input[89]), .Z(n9496) );
  XOR U18358 ( .A(n18439), .B(n18438), .Z(n18437) );
  AND U18359 ( .A(n9498), .B(n9499), .Z(n18438) );
  IV U18360 ( .A(p_input[86]), .Z(n9499) );
  IV U18361 ( .A(p_input[87]), .Z(n9498) );
  XOR U18362 ( .A(n18441), .B(n18440), .Z(n18439) );
  AND U18363 ( .A(n9500), .B(n9501), .Z(n18440) );
  IV U18364 ( .A(p_input[84]), .Z(n9501) );
  IV U18365 ( .A(p_input[85]), .Z(n9500) );
  XOR U18366 ( .A(n18443), .B(n18442), .Z(n18441) );
  AND U18367 ( .A(n9502), .B(n9503), .Z(n18442) );
  IV U18368 ( .A(p_input[82]), .Z(n9503) );
  IV U18369 ( .A(p_input[83]), .Z(n9502) );
  XOR U18370 ( .A(n18445), .B(n18444), .Z(n18443) );
  AND U18371 ( .A(n9504), .B(n9505), .Z(n18444) );
  IV U18372 ( .A(p_input[80]), .Z(n9505) );
  IV U18373 ( .A(p_input[81]), .Z(n9504) );
  XOR U18374 ( .A(n18447), .B(n18446), .Z(n18445) );
  AND U18375 ( .A(n9506), .B(n9507), .Z(n18446) );
  IV U18376 ( .A(p_input[78]), .Z(n9507) );
  IV U18377 ( .A(p_input[79]), .Z(n9506) );
  XOR U18378 ( .A(n18449), .B(n18448), .Z(n18447) );
  AND U18379 ( .A(n9508), .B(n9509), .Z(n18448) );
  IV U18380 ( .A(p_input[76]), .Z(n9509) );
  IV U18381 ( .A(p_input[77]), .Z(n9508) );
  XOR U18382 ( .A(n18451), .B(n18450), .Z(n18449) );
  AND U18383 ( .A(n9510), .B(n9511), .Z(n18450) );
  IV U18384 ( .A(p_input[74]), .Z(n9511) );
  IV U18385 ( .A(p_input[75]), .Z(n9510) );
  XOR U18386 ( .A(n18453), .B(n18452), .Z(n18451) );
  AND U18387 ( .A(n9512), .B(n9513), .Z(n18452) );
  IV U18388 ( .A(p_input[72]), .Z(n9513) );
  IV U18389 ( .A(p_input[73]), .Z(n9512) );
  XOR U18390 ( .A(n18455), .B(n18454), .Z(n18453) );
  AND U18391 ( .A(n9514), .B(n9515), .Z(n18454) );
  IV U18392 ( .A(p_input[70]), .Z(n9515) );
  IV U18393 ( .A(p_input[71]), .Z(n9514) );
  XOR U18394 ( .A(n18457), .B(n18456), .Z(n18455) );
  AND U18395 ( .A(n9516), .B(n9517), .Z(n18456) );
  IV U18396 ( .A(p_input[68]), .Z(n9517) );
  IV U18397 ( .A(p_input[69]), .Z(n9516) );
  XOR U18398 ( .A(n18459), .B(n18458), .Z(n18457) );
  AND U18399 ( .A(n9518), .B(n9519), .Z(n18458) );
  IV U18400 ( .A(p_input[66]), .Z(n9519) );
  IV U18401 ( .A(p_input[67]), .Z(n9518) );
  XOR U18402 ( .A(n18461), .B(n18460), .Z(n18459) );
  AND U18403 ( .A(n9520), .B(n9521), .Z(n18460) );
  IV U18404 ( .A(p_input[64]), .Z(n9521) );
  IV U18405 ( .A(p_input[65]), .Z(n9520) );
  XOR U18406 ( .A(n18463), .B(n18462), .Z(n18461) );
  AND U18407 ( .A(n9522), .B(n9523), .Z(n18462) );
  IV U18408 ( .A(p_input[62]), .Z(n9523) );
  IV U18409 ( .A(p_input[63]), .Z(n9522) );
  XOR U18410 ( .A(n18465), .B(n18464), .Z(n18463) );
  AND U18411 ( .A(n9524), .B(n9525), .Z(n18464) );
  IV U18412 ( .A(p_input[60]), .Z(n9525) );
  IV U18413 ( .A(p_input[61]), .Z(n9524) );
  XOR U18414 ( .A(n18467), .B(n18466), .Z(n18465) );
  AND U18415 ( .A(n9526), .B(n9527), .Z(n18466) );
  IV U18416 ( .A(p_input[58]), .Z(n9527) );
  IV U18417 ( .A(p_input[59]), .Z(n9526) );
  XOR U18418 ( .A(n18469), .B(n18468), .Z(n18467) );
  AND U18419 ( .A(n9528), .B(n9529), .Z(n18468) );
  IV U18420 ( .A(p_input[56]), .Z(n9529) );
  IV U18421 ( .A(p_input[57]), .Z(n9528) );
  XOR U18422 ( .A(n18471), .B(n18470), .Z(n18469) );
  AND U18423 ( .A(n9530), .B(n9531), .Z(n18470) );
  IV U18424 ( .A(p_input[54]), .Z(n9531) );
  IV U18425 ( .A(p_input[55]), .Z(n9530) );
  XOR U18426 ( .A(n18473), .B(n18472), .Z(n18471) );
  AND U18427 ( .A(n9532), .B(n9533), .Z(n18472) );
  IV U18428 ( .A(p_input[52]), .Z(n9533) );
  IV U18429 ( .A(p_input[53]), .Z(n9532) );
  XOR U18430 ( .A(n18475), .B(n18474), .Z(n18473) );
  AND U18431 ( .A(n9534), .B(n9535), .Z(n18474) );
  IV U18432 ( .A(p_input[50]), .Z(n9535) );
  IV U18433 ( .A(p_input[51]), .Z(n9534) );
  XOR U18434 ( .A(n18477), .B(n18476), .Z(n18475) );
  AND U18435 ( .A(n9536), .B(n9537), .Z(n18476) );
  IV U18436 ( .A(p_input[48]), .Z(n9537) );
  IV U18437 ( .A(p_input[49]), .Z(n9536) );
  XOR U18438 ( .A(n18479), .B(n18478), .Z(n18477) );
  AND U18439 ( .A(n9538), .B(n9539), .Z(n18478) );
  IV U18440 ( .A(p_input[46]), .Z(n9539) );
  IV U18441 ( .A(p_input[47]), .Z(n9538) );
  XOR U18442 ( .A(n18481), .B(n18480), .Z(n18479) );
  AND U18443 ( .A(n9540), .B(n9541), .Z(n18480) );
  IV U18444 ( .A(p_input[44]), .Z(n9541) );
  IV U18445 ( .A(p_input[45]), .Z(n9540) );
  XOR U18446 ( .A(n18483), .B(n18482), .Z(n18481) );
  AND U18447 ( .A(n9542), .B(n9543), .Z(n18482) );
  IV U18448 ( .A(p_input[42]), .Z(n9543) );
  IV U18449 ( .A(p_input[43]), .Z(n9542) );
  XOR U18450 ( .A(n18485), .B(n18484), .Z(n18483) );
  AND U18451 ( .A(n9544), .B(n9545), .Z(n18484) );
  IV U18452 ( .A(p_input[40]), .Z(n9545) );
  IV U18453 ( .A(p_input[41]), .Z(n9544) );
  XOR U18454 ( .A(n18487), .B(n18486), .Z(n18485) );
  AND U18455 ( .A(n9546), .B(n9547), .Z(n18486) );
  IV U18456 ( .A(p_input[38]), .Z(n9547) );
  IV U18457 ( .A(p_input[39]), .Z(n9546) );
  XOR U18458 ( .A(n18489), .B(n18488), .Z(n18487) );
  AND U18459 ( .A(n9548), .B(n9549), .Z(n18488) );
  IV U18460 ( .A(p_input[36]), .Z(n9549) );
  IV U18461 ( .A(p_input[37]), .Z(n9548) );
  XOR U18462 ( .A(n18491), .B(n18490), .Z(n18489) );
  AND U18463 ( .A(n9550), .B(n9551), .Z(n18490) );
  IV U18464 ( .A(p_input[34]), .Z(n9551) );
  IV U18465 ( .A(p_input[35]), .Z(n9550) );
  XOR U18466 ( .A(n18493), .B(n18492), .Z(n18491) );
  AND U18467 ( .A(n9552), .B(n9553), .Z(n18492) );
  IV U18468 ( .A(p_input[32]), .Z(n9553) );
  IV U18469 ( .A(p_input[33]), .Z(n9552) );
  XOR U18470 ( .A(n18495), .B(n18494), .Z(n18493) );
  AND U18471 ( .A(n9554), .B(n9555), .Z(n18494) );
  IV U18472 ( .A(p_input[30]), .Z(n9555) );
  IV U18473 ( .A(p_input[31]), .Z(n9554) );
  XOR U18474 ( .A(n18497), .B(n18496), .Z(n18495) );
  AND U18475 ( .A(n9556), .B(n9557), .Z(n18496) );
  IV U18476 ( .A(p_input[28]), .Z(n9557) );
  IV U18477 ( .A(p_input[29]), .Z(n9556) );
  XOR U18478 ( .A(n18499), .B(n18498), .Z(n18497) );
  AND U18479 ( .A(n9558), .B(n9559), .Z(n18498) );
  IV U18480 ( .A(p_input[26]), .Z(n9559) );
  IV U18481 ( .A(p_input[27]), .Z(n9558) );
  XOR U18482 ( .A(n18501), .B(n18500), .Z(n18499) );
  AND U18483 ( .A(n9560), .B(n9561), .Z(n18500) );
  IV U18484 ( .A(p_input[24]), .Z(n9561) );
  IV U18485 ( .A(p_input[25]), .Z(n9560) );
  XOR U18486 ( .A(n18503), .B(n18502), .Z(n18501) );
  AND U18487 ( .A(n9562), .B(n9563), .Z(n18502) );
  IV U18488 ( .A(p_input[22]), .Z(n9563) );
  IV U18489 ( .A(p_input[23]), .Z(n9562) );
  XOR U18490 ( .A(n18505), .B(n18504), .Z(n18503) );
  AND U18491 ( .A(n9564), .B(n9565), .Z(n18504) );
  IV U18492 ( .A(p_input[20]), .Z(n9565) );
  IV U18493 ( .A(p_input[21]), .Z(n9564) );
  XOR U18494 ( .A(n18507), .B(n18506), .Z(n18505) );
  AND U18495 ( .A(n9566), .B(n9567), .Z(n18506) );
  IV U18496 ( .A(p_input[18]), .Z(n9567) );
  IV U18497 ( .A(p_input[19]), .Z(n9566) );
  XOR U18498 ( .A(n18509), .B(n18508), .Z(n18507) );
  AND U18499 ( .A(n9568), .B(n9569), .Z(n18508) );
  IV U18500 ( .A(p_input[16]), .Z(n9569) );
  IV U18501 ( .A(p_input[17]), .Z(n9568) );
  XOR U18502 ( .A(n18511), .B(n18510), .Z(n18509) );
  AND U18503 ( .A(n9570), .B(n9571), .Z(n18510) );
  IV U18504 ( .A(p_input[14]), .Z(n9571) );
  IV U18505 ( .A(p_input[15]), .Z(n9570) );
  XOR U18506 ( .A(n18513), .B(n18512), .Z(n18511) );
  AND U18507 ( .A(n9572), .B(n9573), .Z(n18512) );
  IV U18508 ( .A(p_input[12]), .Z(n9573) );
  IV U18509 ( .A(p_input[13]), .Z(n9572) );
  XOR U18510 ( .A(n18527), .B(n18526), .Z(n18513) );
  AND U18511 ( .A(n9574), .B(n9575), .Z(n18526) );
  IV U18512 ( .A(p_input[10]), .Z(n9575) );
  IV U18513 ( .A(p_input[11]), .Z(n9574) );
  XOR U18514 ( .A(n18529), .B(n18528), .Z(n18527) );
  AND U18515 ( .A(n9576), .B(n9577), .Z(n18528) );
  IV U18516 ( .A(p_input[8]), .Z(n9577) );
  IV U18517 ( .A(p_input[9]), .Z(n9576) );
  XOR U18518 ( .A(n18517), .B(n18516), .Z(n18529) );
  AND U18519 ( .A(n9578), .B(n9579), .Z(n18516) );
  IV U18520 ( .A(p_input[6]), .Z(n9579) );
  IV U18521 ( .A(p_input[7]), .Z(n9578) );
  XOR U18522 ( .A(n18524), .B(n18525), .Z(n18517) );
  XOR U18523 ( .A(n18522), .B(n18523), .Z(n18525) );
  AND U18524 ( .A(n9580), .B(n9581), .Z(n18523) );
  IV U18525 ( .A(p_input[2]), .Z(n9581) );
  IV U18526 ( .A(p_input[3]), .Z(n9580) );
  AND U18527 ( .A(n9582), .B(n9583), .Z(n18522) );
  IV U18528 ( .A(p_input[0]), .Z(n9583) );
  IV U18529 ( .A(p_input[1]), .Z(n9582) );
  AND U18530 ( .A(n9584), .B(n9585), .Z(n18524) );
  IV U18531 ( .A(p_input[4]), .Z(n9585) );
  IV U18532 ( .A(p_input[5]), .Z(n9584) );
endmodule

