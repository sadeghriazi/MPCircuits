
module knn_comb_BMR_W32_K3_N4 ( p_input, o );
  input [159:0] p_input;
  output [95:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/min_val_out[0][16] , \knn_comb_/min_val_out[0][17] ,
         \knn_comb_/min_val_out[0][18] , \knn_comb_/min_val_out[0][19] ,
         \knn_comb_/min_val_out[0][20] , \knn_comb_/min_val_out[0][21] ,
         \knn_comb_/min_val_out[0][22] , \knn_comb_/min_val_out[0][23] ,
         \knn_comb_/min_val_out[0][24] , \knn_comb_/min_val_out[0][25] ,
         \knn_comb_/min_val_out[0][26] , \knn_comb_/min_val_out[0][27] ,
         \knn_comb_/min_val_out[0][28] , \knn_comb_/min_val_out[0][29] ,
         \knn_comb_/min_val_out[0][30] , \knn_comb_/min_val_out[0][31] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][31] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775;
  assign \knn_comb_/min_val_out[0][0]  = p_input[96];
  assign \knn_comb_/min_val_out[0][1]  = p_input[97];
  assign \knn_comb_/min_val_out[0][2]  = p_input[98];
  assign \knn_comb_/min_val_out[0][3]  = p_input[99];
  assign \knn_comb_/min_val_out[0][4]  = p_input[100];
  assign \knn_comb_/min_val_out[0][5]  = p_input[101];
  assign \knn_comb_/min_val_out[0][6]  = p_input[102];
  assign \knn_comb_/min_val_out[0][7]  = p_input[103];
  assign \knn_comb_/min_val_out[0][8]  = p_input[104];
  assign \knn_comb_/min_val_out[0][9]  = p_input[105];
  assign \knn_comb_/min_val_out[0][10]  = p_input[106];
  assign \knn_comb_/min_val_out[0][11]  = p_input[107];
  assign \knn_comb_/min_val_out[0][12]  = p_input[108];
  assign \knn_comb_/min_val_out[0][13]  = p_input[109];
  assign \knn_comb_/min_val_out[0][14]  = p_input[110];
  assign \knn_comb_/min_val_out[0][15]  = p_input[111];
  assign \knn_comb_/min_val_out[0][16]  = p_input[112];
  assign \knn_comb_/min_val_out[0][17]  = p_input[113];
  assign \knn_comb_/min_val_out[0][18]  = p_input[114];
  assign \knn_comb_/min_val_out[0][19]  = p_input[115];
  assign \knn_comb_/min_val_out[0][20]  = p_input[116];
  assign \knn_comb_/min_val_out[0][21]  = p_input[117];
  assign \knn_comb_/min_val_out[0][22]  = p_input[118];
  assign \knn_comb_/min_val_out[0][23]  = p_input[119];
  assign \knn_comb_/min_val_out[0][24]  = p_input[120];
  assign \knn_comb_/min_val_out[0][25]  = p_input[121];
  assign \knn_comb_/min_val_out[0][26]  = p_input[122];
  assign \knn_comb_/min_val_out[0][27]  = p_input[123];
  assign \knn_comb_/min_val_out[0][28]  = p_input[124];
  assign \knn_comb_/min_val_out[0][29]  = p_input[125];
  assign \knn_comb_/min_val_out[0][30]  = p_input[126];
  assign \knn_comb_/min_val_out[0][31]  = p_input[127];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][0]  = p_input[32];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][1]  = p_input[33];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][2]  = p_input[34];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][3]  = p_input[35];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][4]  = p_input[36];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][5]  = p_input[37];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][6]  = p_input[38];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][7]  = p_input[39];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][8]  = p_input[40];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][9]  = p_input[41];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][10]  = p_input[42];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][11]  = p_input[43];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][12]  = p_input[44];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][13]  = p_input[45];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][14]  = p_input[46];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][15]  = p_input[47];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][16]  = p_input[48];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][17]  = p_input[49];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][18]  = p_input[50];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][19]  = p_input[51];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][20]  = p_input[52];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][21]  = p_input[53];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][22]  = p_input[54];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][23]  = p_input[55];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][24]  = p_input[56];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][25]  = p_input[57];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][26]  = p_input[58];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][27]  = p_input[59];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][28]  = p_input[60];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][29]  = p_input[61];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][30]  = p_input[62];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][31]  = p_input[63];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[64];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[65];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[66];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[67];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[68];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[69];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[70];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[71];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[72];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[73];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[74];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[75];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[76];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[77];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[78];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[79];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][16]  = p_input[80];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][17]  = p_input[81];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][18]  = p_input[82];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][19]  = p_input[83];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][20]  = p_input[84];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][21]  = p_input[85];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][22]  = p_input[86];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][23]  = p_input[87];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][24]  = p_input[88];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][25]  = p_input[89];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][26]  = p_input[90];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][27]  = p_input[91];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][28]  = p_input[92];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][29]  = p_input[93];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][30]  = p_input[94];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][31]  = p_input[95];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[95]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[94]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[93]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[92]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[91]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[90]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[8]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[89]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[88]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[87]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[86]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[85]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[84]) );
  XOR U15 ( .A(n29), .B(n30), .Z(o[83]) );
  XOR U16 ( .A(n31), .B(n32), .Z(o[82]) );
  XOR U17 ( .A(n33), .B(n34), .Z(o[81]) );
  XOR U18 ( .A(n35), .B(n36), .Z(o[80]) );
  XOR U19 ( .A(n37), .B(n38), .Z(o[7]) );
  XOR U20 ( .A(n39), .B(n40), .Z(o[79]) );
  XOR U21 ( .A(n41), .B(n42), .Z(o[78]) );
  XOR U22 ( .A(n43), .B(n44), .Z(o[77]) );
  XOR U23 ( .A(n45), .B(n46), .Z(o[76]) );
  XOR U24 ( .A(n47), .B(n48), .Z(o[75]) );
  XOR U25 ( .A(n49), .B(n50), .Z(o[74]) );
  XOR U26 ( .A(n51), .B(n52), .Z(o[73]) );
  XOR U27 ( .A(n53), .B(n54), .Z(o[72]) );
  XOR U28 ( .A(n55), .B(n56), .Z(o[71]) );
  XOR U29 ( .A(n57), .B(n58), .Z(o[70]) );
  XOR U30 ( .A(n59), .B(n60), .Z(o[6]) );
  XOR U31 ( .A(n61), .B(n62), .Z(o[69]) );
  XOR U32 ( .A(n63), .B(n64), .Z(o[68]) );
  XOR U33 ( .A(n65), .B(n66), .Z(o[67]) );
  XOR U34 ( .A(n67), .B(n68), .Z(o[66]) );
  XOR U35 ( .A(n69), .B(n70), .Z(o[65]) );
  XOR U36 ( .A(n71), .B(n72), .Z(o[64]) );
  XOR U37 ( .A(n73), .B(n74), .Z(o[63]) );
  XOR U38 ( .A(n75), .B(n76), .Z(o[62]) );
  XOR U39 ( .A(n77), .B(n78), .Z(o[61]) );
  XOR U40 ( .A(n79), .B(n80), .Z(o[60]) );
  XOR U41 ( .A(n81), .B(n82), .Z(o[5]) );
  XOR U42 ( .A(n83), .B(n84), .Z(o[59]) );
  XOR U43 ( .A(n85), .B(n86), .Z(o[58]) );
  XOR U44 ( .A(n87), .B(n88), .Z(o[57]) );
  XOR U45 ( .A(n89), .B(n90), .Z(o[56]) );
  XOR U46 ( .A(n91), .B(n92), .Z(o[55]) );
  XOR U47 ( .A(n93), .B(n94), .Z(o[54]) );
  XOR U48 ( .A(n95), .B(n96), .Z(o[53]) );
  XOR U49 ( .A(n97), .B(n98), .Z(o[52]) );
  XOR U50 ( .A(n99), .B(n100), .Z(o[51]) );
  XOR U51 ( .A(n101), .B(n102), .Z(o[50]) );
  XOR U52 ( .A(n103), .B(n104), .Z(o[4]) );
  XOR U53 ( .A(n105), .B(n106), .Z(o[49]) );
  XOR U54 ( .A(n107), .B(n108), .Z(o[48]) );
  XOR U55 ( .A(n109), .B(n110), .Z(o[47]) );
  XOR U56 ( .A(n111), .B(n112), .Z(o[46]) );
  XOR U57 ( .A(n113), .B(n114), .Z(o[45]) );
  XOR U58 ( .A(n115), .B(n116), .Z(o[44]) );
  XOR U59 ( .A(n117), .B(n118), .Z(o[43]) );
  XOR U60 ( .A(n119), .B(n120), .Z(o[42]) );
  XOR U61 ( .A(n1), .B(n121), .Z(o[41]) );
  AND U62 ( .A(n122), .B(n123), .Z(n1) );
  XOR U63 ( .A(n2), .B(n121), .Z(n123) );
  XOR U64 ( .A(n124), .B(n51), .Z(n121) );
  AND U65 ( .A(n125), .B(n126), .Z(n51) );
  XNOR U66 ( .A(n127), .B(n52), .Z(n126) );
  XOR U67 ( .A(n128), .B(n129), .Z(n52) );
  AND U68 ( .A(n130), .B(n131), .Z(n129) );
  XOR U69 ( .A(p_input[9]), .B(n128), .Z(n131) );
  XOR U70 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n132), .Z(
        n128) );
  AND U71 ( .A(n133), .B(n134), .Z(n132) );
  IV U72 ( .A(n124), .Z(n127) );
  XOR U73 ( .A(n135), .B(n136), .Z(n124) );
  AND U74 ( .A(n137), .B(n138), .Z(n136) );
  XOR U75 ( .A(n139), .B(n140), .Z(n2) );
  AND U76 ( .A(n141), .B(n138), .Z(n140) );
  XNOR U77 ( .A(n142), .B(n135), .Z(n138) );
  XNOR U78 ( .A(n143), .B(n144), .Z(n135) );
  AND U79 ( .A(n145), .B(n134), .Z(n144) );
  XNOR U80 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n143), .Z(
        n134) );
  XNOR U81 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .B(n146), .Z(
        n143) );
  AND U82 ( .A(n147), .B(n148), .Z(n146) );
  IV U83 ( .A(n142), .Z(n139) );
  XNOR U84 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n149), .Z(n142) );
  AND U85 ( .A(n150), .B(n148), .Z(n149) );
  XOR U86 ( .A(\knn_comb_/min_val_out[0][9] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n148) );
  XOR U87 ( .A(n15), .B(n151), .Z(o[40]) );
  AND U88 ( .A(n122), .B(n152), .Z(n15) );
  XOR U89 ( .A(n16), .B(n151), .Z(n152) );
  XOR U90 ( .A(n153), .B(n53), .Z(n151) );
  AND U91 ( .A(n125), .B(n154), .Z(n53) );
  XNOR U92 ( .A(n155), .B(n54), .Z(n154) );
  XOR U93 ( .A(n156), .B(n157), .Z(n54) );
  AND U94 ( .A(n130), .B(n158), .Z(n157) );
  XOR U95 ( .A(p_input[8]), .B(n156), .Z(n158) );
  XOR U96 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n159), .Z(
        n156) );
  AND U97 ( .A(n133), .B(n160), .Z(n159) );
  IV U98 ( .A(n153), .Z(n155) );
  XOR U99 ( .A(n161), .B(n162), .Z(n153) );
  AND U100 ( .A(n137), .B(n163), .Z(n162) );
  XOR U101 ( .A(n164), .B(n165), .Z(n16) );
  AND U102 ( .A(n141), .B(n163), .Z(n165) );
  XNOR U103 ( .A(n166), .B(n161), .Z(n163) );
  XNOR U104 ( .A(n167), .B(n168), .Z(n161) );
  AND U105 ( .A(n145), .B(n160), .Z(n168) );
  XNOR U106 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n167), .Z(
        n160) );
  XNOR U107 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n169), .Z(
        n167) );
  AND U108 ( .A(n147), .B(n170), .Z(n169) );
  IV U109 ( .A(n166), .Z(n164) );
  XNOR U110 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n171), .Z(n166) );
  AND U111 ( .A(n150), .B(n170), .Z(n171) );
  XOR U112 ( .A(\knn_comb_/min_val_out[0][8] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n170) );
  XOR U113 ( .A(n172), .B(n173), .Z(o[3]) );
  XOR U114 ( .A(n37), .B(n174), .Z(o[39]) );
  AND U115 ( .A(n122), .B(n175), .Z(n37) );
  XOR U116 ( .A(n38), .B(n174), .Z(n175) );
  XOR U117 ( .A(n176), .B(n55), .Z(n174) );
  AND U118 ( .A(n125), .B(n177), .Z(n55) );
  XNOR U119 ( .A(n178), .B(n56), .Z(n177) );
  XOR U120 ( .A(n179), .B(n180), .Z(n56) );
  AND U121 ( .A(n130), .B(n181), .Z(n180) );
  XOR U122 ( .A(p_input[7]), .B(n179), .Z(n181) );
  XOR U123 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n182), .Z(
        n179) );
  AND U124 ( .A(n133), .B(n183), .Z(n182) );
  IV U125 ( .A(n176), .Z(n178) );
  XOR U126 ( .A(n184), .B(n185), .Z(n176) );
  AND U127 ( .A(n137), .B(n186), .Z(n185) );
  XOR U128 ( .A(n187), .B(n188), .Z(n38) );
  AND U129 ( .A(n141), .B(n186), .Z(n188) );
  XNOR U130 ( .A(n189), .B(n184), .Z(n186) );
  XNOR U131 ( .A(n190), .B(n191), .Z(n184) );
  AND U132 ( .A(n145), .B(n183), .Z(n191) );
  XNOR U133 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n190), .Z(
        n183) );
  XNOR U134 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(n192), .Z(
        n190) );
  AND U135 ( .A(n147), .B(n193), .Z(n192) );
  IV U136 ( .A(n189), .Z(n187) );
  XNOR U137 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n194), .Z(n189) );
  AND U138 ( .A(n150), .B(n193), .Z(n194) );
  XOR U139 ( .A(\knn_comb_/min_val_out[0][7] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n193) );
  XOR U140 ( .A(n59), .B(n195), .Z(o[38]) );
  AND U141 ( .A(n122), .B(n196), .Z(n59) );
  XOR U142 ( .A(n60), .B(n195), .Z(n196) );
  XOR U143 ( .A(n197), .B(n57), .Z(n195) );
  AND U144 ( .A(n125), .B(n198), .Z(n57) );
  XOR U145 ( .A(n58), .B(n197), .Z(n198) );
  XOR U146 ( .A(n199), .B(n200), .Z(n58) );
  AND U147 ( .A(n130), .B(n201), .Z(n200) );
  XOR U148 ( .A(p_input[6]), .B(n199), .Z(n201) );
  XOR U149 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n202), .Z(
        n199) );
  AND U150 ( .A(n133), .B(n203), .Z(n202) );
  XOR U151 ( .A(n204), .B(n205), .Z(n197) );
  AND U152 ( .A(n137), .B(n206), .Z(n205) );
  XOR U153 ( .A(n207), .B(n208), .Z(n60) );
  AND U154 ( .A(n141), .B(n206), .Z(n208) );
  XNOR U155 ( .A(n209), .B(n207), .Z(n206) );
  IV U156 ( .A(n204), .Z(n209) );
  XOR U157 ( .A(n210), .B(n211), .Z(n204) );
  AND U158 ( .A(n145), .B(n203), .Z(n211) );
  XOR U159 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n210), .Z(
        n203) );
  XOR U160 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(n212), .Z(
        n210) );
  AND U161 ( .A(n147), .B(n213), .Z(n212) );
  XOR U162 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n214), .Z(n207) );
  AND U163 ( .A(n150), .B(n213), .Z(n214) );
  XOR U164 ( .A(\knn_comb_/min_val_out[0][6] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n213) );
  XOR U165 ( .A(n81), .B(n215), .Z(o[37]) );
  AND U166 ( .A(n122), .B(n216), .Z(n81) );
  XOR U167 ( .A(n82), .B(n215), .Z(n216) );
  XOR U168 ( .A(n217), .B(n61), .Z(n215) );
  AND U169 ( .A(n125), .B(n218), .Z(n61) );
  XOR U170 ( .A(n62), .B(n217), .Z(n218) );
  XOR U171 ( .A(n219), .B(n220), .Z(n62) );
  AND U172 ( .A(n130), .B(n221), .Z(n220) );
  XOR U173 ( .A(p_input[5]), .B(n219), .Z(n221) );
  XOR U174 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n222), .Z(
        n219) );
  AND U175 ( .A(n133), .B(n223), .Z(n222) );
  XOR U176 ( .A(n224), .B(n225), .Z(n217) );
  AND U177 ( .A(n137), .B(n226), .Z(n225) );
  XOR U178 ( .A(n227), .B(n228), .Z(n82) );
  AND U179 ( .A(n141), .B(n226), .Z(n228) );
  XNOR U180 ( .A(n229), .B(n227), .Z(n226) );
  IV U181 ( .A(n224), .Z(n229) );
  XOR U182 ( .A(n230), .B(n231), .Z(n224) );
  AND U183 ( .A(n145), .B(n223), .Z(n231) );
  XOR U184 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n230), .Z(
        n223) );
  XOR U185 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n232), .Z(
        n230) );
  AND U186 ( .A(n147), .B(n233), .Z(n232) );
  XOR U187 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n234), .Z(n227) );
  AND U188 ( .A(n150), .B(n233), .Z(n234) );
  XOR U189 ( .A(n235), .B(n236), .Z(n233) );
  IV U190 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n236) );
  IV U191 ( .A(\knn_comb_/min_val_out[0][5] ), .Z(n235) );
  XOR U192 ( .A(n103), .B(n237), .Z(o[36]) );
  AND U193 ( .A(n122), .B(n238), .Z(n103) );
  XOR U194 ( .A(n104), .B(n237), .Z(n238) );
  XOR U195 ( .A(n239), .B(n63), .Z(n237) );
  AND U196 ( .A(n125), .B(n240), .Z(n63) );
  XOR U197 ( .A(n64), .B(n239), .Z(n240) );
  XOR U198 ( .A(n241), .B(n242), .Z(n64) );
  AND U199 ( .A(n130), .B(n243), .Z(n242) );
  XOR U200 ( .A(p_input[4]), .B(n241), .Z(n243) );
  XOR U201 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n244), .Z(
        n241) );
  AND U202 ( .A(n133), .B(n245), .Z(n244) );
  XOR U203 ( .A(n246), .B(n247), .Z(n239) );
  AND U204 ( .A(n137), .B(n248), .Z(n247) );
  XOR U205 ( .A(n249), .B(n250), .Z(n104) );
  AND U206 ( .A(n141), .B(n248), .Z(n250) );
  XNOR U207 ( .A(n251), .B(n249), .Z(n248) );
  IV U208 ( .A(n246), .Z(n251) );
  XOR U209 ( .A(n252), .B(n253), .Z(n246) );
  AND U210 ( .A(n145), .B(n245), .Z(n253) );
  XOR U211 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n252), .Z(
        n245) );
  XOR U212 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n254), .Z(
        n252) );
  AND U213 ( .A(n147), .B(n255), .Z(n254) );
  XOR U214 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n256), .Z(n249) );
  AND U215 ( .A(n150), .B(n255), .Z(n256) );
  XOR U216 ( .A(\knn_comb_/min_val_out[0][4] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n255) );
  XOR U217 ( .A(n172), .B(n257), .Z(o[35]) );
  AND U218 ( .A(n122), .B(n258), .Z(n172) );
  XOR U219 ( .A(n173), .B(n257), .Z(n258) );
  XOR U220 ( .A(n259), .B(n65), .Z(n257) );
  AND U221 ( .A(n125), .B(n260), .Z(n65) );
  XOR U222 ( .A(n66), .B(n259), .Z(n260) );
  XOR U223 ( .A(n261), .B(n262), .Z(n66) );
  AND U224 ( .A(n130), .B(n263), .Z(n262) );
  XOR U225 ( .A(p_input[3]), .B(n261), .Z(n263) );
  XOR U226 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n264), .Z(
        n261) );
  AND U227 ( .A(n133), .B(n265), .Z(n264) );
  XOR U228 ( .A(n266), .B(n267), .Z(n259) );
  AND U229 ( .A(n137), .B(n268), .Z(n267) );
  XOR U230 ( .A(n269), .B(n270), .Z(n173) );
  AND U231 ( .A(n141), .B(n268), .Z(n270) );
  XNOR U232 ( .A(n271), .B(n269), .Z(n268) );
  IV U233 ( .A(n266), .Z(n271) );
  XOR U234 ( .A(n272), .B(n273), .Z(n266) );
  AND U235 ( .A(n145), .B(n265), .Z(n273) );
  XOR U236 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n272), .Z(
        n265) );
  XOR U237 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(n274), .Z(
        n272) );
  AND U238 ( .A(n147), .B(n275), .Z(n274) );
  XOR U239 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n276), .Z(n269) );
  AND U240 ( .A(n150), .B(n275), .Z(n276) );
  XOR U241 ( .A(\knn_comb_/min_val_out[0][3] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n275) );
  XOR U242 ( .A(n277), .B(n278), .Z(o[34]) );
  XOR U243 ( .A(n279), .B(n280), .Z(o[33]) );
  XOR U244 ( .A(n281), .B(n282), .Z(o[32]) );
  XOR U245 ( .A(n73), .B(n283), .Z(o[31]) );
  AND U246 ( .A(n122), .B(n284), .Z(n73) );
  XOR U247 ( .A(n74), .B(n283), .Z(n284) );
  XOR U248 ( .A(n285), .B(n286), .Z(n283) );
  AND U249 ( .A(n141), .B(n287), .Z(n286) );
  XOR U250 ( .A(n288), .B(n3), .Z(n74) );
  AND U251 ( .A(n125), .B(n289), .Z(n3) );
  XOR U252 ( .A(n4), .B(n288), .Z(n289) );
  XOR U253 ( .A(n290), .B(n291), .Z(n4) );
  AND U254 ( .A(n130), .B(n292), .Z(n291) );
  XOR U255 ( .A(p_input[31]), .B(n290), .Z(n292) );
  XOR U256 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ), .B(n293), .Z(
        n290) );
  AND U257 ( .A(n133), .B(n294), .Z(n293) );
  XOR U258 ( .A(n295), .B(n296), .Z(n288) );
  AND U259 ( .A(n137), .B(n287), .Z(n296) );
  XNOR U260 ( .A(n297), .B(n285), .Z(n287) );
  XOR U261 ( .A(\knn_comb_/min_val_out[0][31] ), .B(n298), .Z(n285) );
  AND U262 ( .A(n150), .B(n299), .Z(n298) );
  IV U263 ( .A(n295), .Z(n297) );
  XOR U264 ( .A(n300), .B(n301), .Z(n295) );
  AND U265 ( .A(n145), .B(n294), .Z(n301) );
  XOR U266 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ), .B(n300), .Z(
        n294) );
  XOR U267 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .B(n302), .Z(
        n300) );
  AND U268 ( .A(n147), .B(n299), .Z(n302) );
  XOR U269 ( .A(n303), .B(n304), .Z(n299) );
  IV U270 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .Z(n304) );
  IV U271 ( .A(\knn_comb_/min_val_out[0][31] ), .Z(n303) );
  XOR U272 ( .A(n75), .B(n305), .Z(o[30]) );
  AND U273 ( .A(n122), .B(n306), .Z(n75) );
  XOR U274 ( .A(n76), .B(n305), .Z(n306) );
  XOR U275 ( .A(n307), .B(n308), .Z(n305) );
  AND U276 ( .A(n141), .B(n309), .Z(n308) );
  XOR U277 ( .A(n310), .B(n5), .Z(n76) );
  AND U278 ( .A(n125), .B(n311), .Z(n5) );
  XOR U279 ( .A(n6), .B(n310), .Z(n311) );
  XOR U280 ( .A(n312), .B(n313), .Z(n6) );
  AND U281 ( .A(n130), .B(n314), .Z(n313) );
  XOR U282 ( .A(p_input[30]), .B(n312), .Z(n314) );
  XOR U283 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ), .B(n315), .Z(
        n312) );
  AND U284 ( .A(n133), .B(n316), .Z(n315) );
  XOR U285 ( .A(n317), .B(n318), .Z(n310) );
  AND U286 ( .A(n137), .B(n309), .Z(n318) );
  XNOR U287 ( .A(n319), .B(n307), .Z(n309) );
  XOR U288 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n320), .Z(n307) );
  AND U289 ( .A(n150), .B(n321), .Z(n320) );
  IV U290 ( .A(n317), .Z(n319) );
  XOR U291 ( .A(n322), .B(n323), .Z(n317) );
  AND U292 ( .A(n145), .B(n316), .Z(n323) );
  XOR U293 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ), .B(n322), .Z(
        n316) );
  XOR U294 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .B(n324), .Z(
        n322) );
  AND U295 ( .A(n147), .B(n321), .Z(n324) );
  XOR U296 ( .A(n325), .B(n326), .Z(n321) );
  IV U297 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .Z(n326) );
  IV U298 ( .A(\knn_comb_/min_val_out[0][30] ), .Z(n325) );
  XOR U299 ( .A(n277), .B(n327), .Z(o[2]) );
  AND U300 ( .A(n122), .B(n328), .Z(n277) );
  XOR U301 ( .A(n278), .B(n327), .Z(n328) );
  XOR U302 ( .A(n329), .B(n330), .Z(n327) );
  AND U303 ( .A(n141), .B(n331), .Z(n330) );
  XOR U304 ( .A(n332), .B(n67), .Z(n278) );
  AND U305 ( .A(n125), .B(n333), .Z(n67) );
  XOR U306 ( .A(n68), .B(n332), .Z(n333) );
  XOR U307 ( .A(n334), .B(n335), .Z(n68) );
  AND U308 ( .A(n130), .B(n336), .Z(n335) );
  XOR U309 ( .A(p_input[2]), .B(n334), .Z(n336) );
  XOR U310 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n337), .Z(
        n334) );
  AND U311 ( .A(n133), .B(n338), .Z(n337) );
  XOR U312 ( .A(n339), .B(n340), .Z(n332) );
  AND U313 ( .A(n137), .B(n331), .Z(n340) );
  XNOR U314 ( .A(n341), .B(n329), .Z(n331) );
  XOR U315 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n342), .Z(n329) );
  AND U316 ( .A(n150), .B(n343), .Z(n342) );
  IV U317 ( .A(n339), .Z(n341) );
  XOR U318 ( .A(n344), .B(n345), .Z(n339) );
  AND U319 ( .A(n145), .B(n338), .Z(n345) );
  XOR U320 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n344), .Z(
        n338) );
  XOR U321 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(n346), .Z(
        n344) );
  AND U322 ( .A(n147), .B(n343), .Z(n346) );
  XOR U323 ( .A(\knn_comb_/min_val_out[0][2] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n343) );
  XOR U324 ( .A(n77), .B(n347), .Z(o[29]) );
  AND U325 ( .A(n122), .B(n348), .Z(n77) );
  XOR U326 ( .A(n78), .B(n347), .Z(n348) );
  XOR U327 ( .A(n349), .B(n350), .Z(n347) );
  AND U328 ( .A(n141), .B(n351), .Z(n350) );
  XOR U329 ( .A(n352), .B(n7), .Z(n78) );
  AND U330 ( .A(n125), .B(n353), .Z(n7) );
  XOR U331 ( .A(n8), .B(n352), .Z(n353) );
  XOR U332 ( .A(n354), .B(n355), .Z(n8) );
  AND U333 ( .A(n130), .B(n356), .Z(n355) );
  XOR U334 ( .A(p_input[29]), .B(n354), .Z(n356) );
  XOR U335 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ), .B(n357), .Z(
        n354) );
  AND U336 ( .A(n133), .B(n358), .Z(n357) );
  XOR U337 ( .A(n359), .B(n360), .Z(n352) );
  AND U338 ( .A(n137), .B(n351), .Z(n360) );
  XNOR U339 ( .A(n361), .B(n349), .Z(n351) );
  XOR U340 ( .A(\knn_comb_/min_val_out[0][29] ), .B(n362), .Z(n349) );
  AND U341 ( .A(n150), .B(n363), .Z(n362) );
  IV U342 ( .A(n359), .Z(n361) );
  XOR U343 ( .A(n364), .B(n365), .Z(n359) );
  AND U344 ( .A(n145), .B(n358), .Z(n365) );
  XOR U345 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ), .B(n364), .Z(
        n358) );
  XOR U346 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .B(n366), .Z(
        n364) );
  AND U347 ( .A(n147), .B(n363), .Z(n366) );
  XOR U348 ( .A(\knn_comb_/min_val_out[0][29] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .Z(n363) );
  XOR U349 ( .A(n79), .B(n367), .Z(o[28]) );
  AND U350 ( .A(n122), .B(n368), .Z(n79) );
  XOR U351 ( .A(n80), .B(n367), .Z(n368) );
  XOR U352 ( .A(n369), .B(n370), .Z(n367) );
  AND U353 ( .A(n141), .B(n371), .Z(n370) );
  XOR U354 ( .A(n372), .B(n9), .Z(n80) );
  AND U355 ( .A(n125), .B(n373), .Z(n9) );
  XOR U356 ( .A(n10), .B(n372), .Z(n373) );
  XOR U357 ( .A(n374), .B(n375), .Z(n10) );
  AND U358 ( .A(n130), .B(n376), .Z(n375) );
  XOR U359 ( .A(p_input[28]), .B(n374), .Z(n376) );
  XOR U360 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ), .B(n377), .Z(
        n374) );
  AND U361 ( .A(n133), .B(n378), .Z(n377) );
  XOR U362 ( .A(n379), .B(n380), .Z(n372) );
  AND U363 ( .A(n137), .B(n371), .Z(n380) );
  XNOR U364 ( .A(n381), .B(n369), .Z(n371) );
  XOR U365 ( .A(\knn_comb_/min_val_out[0][28] ), .B(n382), .Z(n369) );
  AND U366 ( .A(n150), .B(n383), .Z(n382) );
  IV U367 ( .A(n379), .Z(n381) );
  XOR U368 ( .A(n384), .B(n385), .Z(n379) );
  AND U369 ( .A(n145), .B(n378), .Z(n385) );
  XOR U370 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ), .B(n384), .Z(
        n378) );
  XOR U371 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .B(n386), .Z(
        n384) );
  AND U372 ( .A(n147), .B(n383), .Z(n386) );
  XOR U373 ( .A(\knn_comb_/min_val_out[0][28] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .Z(n383) );
  XOR U374 ( .A(n83), .B(n387), .Z(o[27]) );
  AND U375 ( .A(n122), .B(n388), .Z(n83) );
  XOR U376 ( .A(n84), .B(n387), .Z(n388) );
  XOR U377 ( .A(n389), .B(n390), .Z(n387) );
  AND U378 ( .A(n141), .B(n391), .Z(n390) );
  XOR U379 ( .A(n392), .B(n11), .Z(n84) );
  AND U380 ( .A(n125), .B(n393), .Z(n11) );
  XOR U381 ( .A(n12), .B(n392), .Z(n393) );
  XOR U382 ( .A(n394), .B(n395), .Z(n12) );
  AND U383 ( .A(n130), .B(n396), .Z(n395) );
  XOR U384 ( .A(p_input[27]), .B(n394), .Z(n396) );
  XOR U385 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ), .B(n397), .Z(
        n394) );
  AND U386 ( .A(n133), .B(n398), .Z(n397) );
  XOR U387 ( .A(n399), .B(n400), .Z(n392) );
  AND U388 ( .A(n137), .B(n391), .Z(n400) );
  XNOR U389 ( .A(n401), .B(n389), .Z(n391) );
  XOR U390 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n402), .Z(n389) );
  AND U391 ( .A(n150), .B(n403), .Z(n402) );
  IV U392 ( .A(n399), .Z(n401) );
  XOR U393 ( .A(n404), .B(n405), .Z(n399) );
  AND U394 ( .A(n145), .B(n398), .Z(n405) );
  XOR U395 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ), .B(n404), .Z(
        n398) );
  XOR U396 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .B(n406), .Z(
        n404) );
  AND U397 ( .A(n147), .B(n403), .Z(n406) );
  XOR U398 ( .A(n407), .B(n408), .Z(n403) );
  IV U399 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .Z(n408) );
  IV U400 ( .A(\knn_comb_/min_val_out[0][27] ), .Z(n407) );
  XOR U401 ( .A(n85), .B(n409), .Z(o[26]) );
  AND U402 ( .A(n122), .B(n410), .Z(n85) );
  XOR U403 ( .A(n86), .B(n409), .Z(n410) );
  XOR U404 ( .A(n411), .B(n412), .Z(n409) );
  AND U405 ( .A(n141), .B(n413), .Z(n412) );
  XOR U406 ( .A(n414), .B(n13), .Z(n86) );
  AND U407 ( .A(n125), .B(n415), .Z(n13) );
  XOR U408 ( .A(n14), .B(n414), .Z(n415) );
  XOR U409 ( .A(n416), .B(n417), .Z(n14) );
  AND U410 ( .A(n130), .B(n418), .Z(n417) );
  XOR U411 ( .A(p_input[26]), .B(n416), .Z(n418) );
  XOR U412 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ), .B(n419), .Z(
        n416) );
  AND U413 ( .A(n133), .B(n420), .Z(n419) );
  XOR U414 ( .A(n421), .B(n422), .Z(n414) );
  AND U415 ( .A(n137), .B(n413), .Z(n422) );
  XNOR U416 ( .A(n423), .B(n411), .Z(n413) );
  XOR U417 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n424), .Z(n411) );
  AND U418 ( .A(n150), .B(n425), .Z(n424) );
  IV U419 ( .A(n421), .Z(n423) );
  XOR U420 ( .A(n426), .B(n427), .Z(n421) );
  AND U421 ( .A(n145), .B(n420), .Z(n427) );
  XOR U422 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ), .B(n426), .Z(
        n420) );
  XOR U423 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .B(n428), .Z(
        n426) );
  AND U424 ( .A(n147), .B(n425), .Z(n428) );
  XOR U425 ( .A(\knn_comb_/min_val_out[0][26] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .Z(n425) );
  XOR U426 ( .A(n87), .B(n429), .Z(o[25]) );
  AND U427 ( .A(n122), .B(n430), .Z(n87) );
  XOR U428 ( .A(n88), .B(n429), .Z(n430) );
  XOR U429 ( .A(n431), .B(n432), .Z(n429) );
  AND U430 ( .A(n141), .B(n433), .Z(n432) );
  XOR U431 ( .A(n434), .B(n17), .Z(n88) );
  AND U432 ( .A(n125), .B(n435), .Z(n17) );
  XOR U433 ( .A(n18), .B(n434), .Z(n435) );
  XOR U434 ( .A(n436), .B(n437), .Z(n18) );
  AND U435 ( .A(n130), .B(n438), .Z(n437) );
  XOR U436 ( .A(p_input[25]), .B(n436), .Z(n438) );
  XOR U437 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ), .B(n439), .Z(
        n436) );
  AND U438 ( .A(n133), .B(n440), .Z(n439) );
  XOR U439 ( .A(n441), .B(n442), .Z(n434) );
  AND U440 ( .A(n137), .B(n433), .Z(n442) );
  XNOR U441 ( .A(n443), .B(n431), .Z(n433) );
  XOR U442 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n444), .Z(n431) );
  AND U443 ( .A(n150), .B(n445), .Z(n444) );
  IV U444 ( .A(n441), .Z(n443) );
  XOR U445 ( .A(n446), .B(n447), .Z(n441) );
  AND U446 ( .A(n145), .B(n440), .Z(n447) );
  XOR U447 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ), .B(n446), .Z(
        n440) );
  XOR U448 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .B(n448), .Z(
        n446) );
  AND U449 ( .A(n147), .B(n445), .Z(n448) );
  XOR U450 ( .A(\knn_comb_/min_val_out[0][25] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .Z(n445) );
  XOR U451 ( .A(n89), .B(n449), .Z(o[24]) );
  AND U452 ( .A(n122), .B(n450), .Z(n89) );
  XOR U453 ( .A(n90), .B(n449), .Z(n450) );
  XOR U454 ( .A(n451), .B(n452), .Z(n449) );
  AND U455 ( .A(n141), .B(n453), .Z(n452) );
  XOR U456 ( .A(n454), .B(n19), .Z(n90) );
  AND U457 ( .A(n125), .B(n455), .Z(n19) );
  XOR U458 ( .A(n20), .B(n454), .Z(n455) );
  XOR U459 ( .A(n456), .B(n457), .Z(n20) );
  AND U460 ( .A(n130), .B(n458), .Z(n457) );
  XOR U461 ( .A(p_input[24]), .B(n456), .Z(n458) );
  XOR U462 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ), .B(n459), .Z(
        n456) );
  AND U463 ( .A(n133), .B(n460), .Z(n459) );
  XOR U464 ( .A(n461), .B(n462), .Z(n454) );
  AND U465 ( .A(n137), .B(n453), .Z(n462) );
  XNOR U466 ( .A(n463), .B(n451), .Z(n453) );
  XOR U467 ( .A(\knn_comb_/min_val_out[0][24] ), .B(n464), .Z(n451) );
  AND U468 ( .A(n150), .B(n465), .Z(n464) );
  IV U469 ( .A(n461), .Z(n463) );
  XOR U470 ( .A(n466), .B(n467), .Z(n461) );
  AND U471 ( .A(n145), .B(n460), .Z(n467) );
  XOR U472 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ), .B(n466), .Z(
        n460) );
  XOR U473 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .B(n468), .Z(
        n466) );
  AND U474 ( .A(n147), .B(n465), .Z(n468) );
  XOR U475 ( .A(\knn_comb_/min_val_out[0][24] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .Z(n465) );
  XOR U476 ( .A(n91), .B(n469), .Z(o[23]) );
  AND U477 ( .A(n122), .B(n470), .Z(n91) );
  XOR U478 ( .A(n92), .B(n469), .Z(n470) );
  XOR U479 ( .A(n471), .B(n472), .Z(n469) );
  AND U480 ( .A(n141), .B(n473), .Z(n472) );
  XOR U481 ( .A(n474), .B(n21), .Z(n92) );
  AND U482 ( .A(n125), .B(n475), .Z(n21) );
  XOR U483 ( .A(n22), .B(n474), .Z(n475) );
  XOR U484 ( .A(n476), .B(n477), .Z(n22) );
  AND U485 ( .A(n130), .B(n478), .Z(n477) );
  XOR U486 ( .A(p_input[23]), .B(n476), .Z(n478) );
  XOR U487 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ), .B(n479), .Z(
        n476) );
  AND U488 ( .A(n133), .B(n480), .Z(n479) );
  XOR U489 ( .A(n481), .B(n482), .Z(n474) );
  AND U490 ( .A(n137), .B(n473), .Z(n482) );
  XNOR U491 ( .A(n483), .B(n471), .Z(n473) );
  XOR U492 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n484), .Z(n471) );
  AND U493 ( .A(n150), .B(n485), .Z(n484) );
  IV U494 ( .A(n481), .Z(n483) );
  XOR U495 ( .A(n486), .B(n487), .Z(n481) );
  AND U496 ( .A(n145), .B(n480), .Z(n487) );
  XOR U497 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ), .B(n486), .Z(
        n480) );
  XOR U498 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .B(n488), .Z(
        n486) );
  AND U499 ( .A(n147), .B(n485), .Z(n488) );
  XOR U500 ( .A(n489), .B(n490), .Z(n485) );
  IV U501 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .Z(n490) );
  IV U502 ( .A(\knn_comb_/min_val_out[0][23] ), .Z(n489) );
  XOR U503 ( .A(n93), .B(n491), .Z(o[22]) );
  AND U504 ( .A(n122), .B(n492), .Z(n93) );
  XOR U505 ( .A(n94), .B(n491), .Z(n492) );
  XOR U506 ( .A(n493), .B(n494), .Z(n491) );
  AND U507 ( .A(n141), .B(n495), .Z(n494) );
  XOR U508 ( .A(n496), .B(n23), .Z(n94) );
  AND U509 ( .A(n125), .B(n497), .Z(n23) );
  XOR U510 ( .A(n24), .B(n496), .Z(n497) );
  XOR U511 ( .A(n498), .B(n499), .Z(n24) );
  AND U512 ( .A(n130), .B(n500), .Z(n499) );
  XOR U513 ( .A(p_input[22]), .B(n498), .Z(n500) );
  XOR U514 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ), .B(n501), .Z(
        n498) );
  AND U515 ( .A(n133), .B(n502), .Z(n501) );
  XOR U516 ( .A(n503), .B(n504), .Z(n496) );
  AND U517 ( .A(n137), .B(n495), .Z(n504) );
  XNOR U518 ( .A(n505), .B(n493), .Z(n495) );
  XOR U519 ( .A(\knn_comb_/min_val_out[0][22] ), .B(n506), .Z(n493) );
  AND U520 ( .A(n150), .B(n507), .Z(n506) );
  IV U521 ( .A(n503), .Z(n505) );
  XOR U522 ( .A(n508), .B(n509), .Z(n503) );
  AND U523 ( .A(n145), .B(n502), .Z(n509) );
  XOR U524 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ), .B(n508), .Z(
        n502) );
  XOR U525 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .B(n510), .Z(
        n508) );
  AND U526 ( .A(n147), .B(n507), .Z(n510) );
  XOR U527 ( .A(\knn_comb_/min_val_out[0][22] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .Z(n507) );
  XOR U528 ( .A(n95), .B(n511), .Z(o[21]) );
  AND U529 ( .A(n122), .B(n512), .Z(n95) );
  XOR U530 ( .A(n96), .B(n511), .Z(n512) );
  XOR U531 ( .A(n513), .B(n514), .Z(n511) );
  AND U532 ( .A(n141), .B(n515), .Z(n514) );
  XOR U533 ( .A(n516), .B(n25), .Z(n96) );
  AND U534 ( .A(n125), .B(n517), .Z(n25) );
  XOR U535 ( .A(n26), .B(n516), .Z(n517) );
  XOR U536 ( .A(n518), .B(n519), .Z(n26) );
  AND U537 ( .A(n130), .B(n520), .Z(n519) );
  XOR U538 ( .A(p_input[21]), .B(n518), .Z(n520) );
  XOR U539 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ), .B(n521), .Z(
        n518) );
  AND U540 ( .A(n133), .B(n522), .Z(n521) );
  XOR U541 ( .A(n523), .B(n524), .Z(n516) );
  AND U542 ( .A(n137), .B(n515), .Z(n524) );
  XNOR U543 ( .A(n525), .B(n513), .Z(n515) );
  XOR U544 ( .A(\knn_comb_/min_val_out[0][21] ), .B(n526), .Z(n513) );
  AND U545 ( .A(n150), .B(n527), .Z(n526) );
  IV U546 ( .A(n523), .Z(n525) );
  XOR U547 ( .A(n528), .B(n529), .Z(n523) );
  AND U548 ( .A(n145), .B(n522), .Z(n529) );
  XOR U549 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ), .B(n528), .Z(
        n522) );
  XOR U550 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .B(n530), .Z(
        n528) );
  AND U551 ( .A(n147), .B(n527), .Z(n530) );
  XOR U552 ( .A(\knn_comb_/min_val_out[0][21] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .Z(n527) );
  XOR U553 ( .A(n97), .B(n531), .Z(o[20]) );
  AND U554 ( .A(n122), .B(n532), .Z(n97) );
  XOR U555 ( .A(n98), .B(n531), .Z(n532) );
  XOR U556 ( .A(n533), .B(n534), .Z(n531) );
  AND U557 ( .A(n141), .B(n535), .Z(n534) );
  XOR U558 ( .A(n536), .B(n27), .Z(n98) );
  AND U559 ( .A(n125), .B(n537), .Z(n27) );
  XOR U560 ( .A(n28), .B(n536), .Z(n537) );
  XOR U561 ( .A(n538), .B(n539), .Z(n28) );
  AND U562 ( .A(n130), .B(n540), .Z(n539) );
  XOR U563 ( .A(p_input[20]), .B(n538), .Z(n540) );
  XOR U564 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ), .B(n541), .Z(
        n538) );
  AND U565 ( .A(n133), .B(n542), .Z(n541) );
  XOR U566 ( .A(n543), .B(n544), .Z(n536) );
  AND U567 ( .A(n137), .B(n535), .Z(n544) );
  XNOR U568 ( .A(n545), .B(n533), .Z(n535) );
  XOR U569 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n546), .Z(n533) );
  AND U570 ( .A(n150), .B(n547), .Z(n546) );
  IV U571 ( .A(n543), .Z(n545) );
  XOR U572 ( .A(n548), .B(n549), .Z(n543) );
  AND U573 ( .A(n145), .B(n542), .Z(n549) );
  XOR U574 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ), .B(n548), .Z(
        n542) );
  XOR U575 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .B(n550), .Z(
        n548) );
  AND U576 ( .A(n147), .B(n547), .Z(n550) );
  XOR U577 ( .A(n551), .B(n552), .Z(n547) );
  IV U578 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .Z(n552) );
  IV U579 ( .A(\knn_comb_/min_val_out[0][20] ), .Z(n551) );
  XOR U580 ( .A(n279), .B(n553), .Z(o[1]) );
  AND U581 ( .A(n122), .B(n554), .Z(n279) );
  XOR U582 ( .A(n280), .B(n553), .Z(n554) );
  XOR U583 ( .A(n555), .B(n556), .Z(n553) );
  AND U584 ( .A(n141), .B(n557), .Z(n556) );
  XOR U585 ( .A(n558), .B(n69), .Z(n280) );
  AND U586 ( .A(n125), .B(n559), .Z(n69) );
  XOR U587 ( .A(n70), .B(n558), .Z(n559) );
  XOR U588 ( .A(n560), .B(n561), .Z(n70) );
  AND U589 ( .A(n130), .B(n562), .Z(n561) );
  XOR U590 ( .A(p_input[1]), .B(n560), .Z(n562) );
  XOR U591 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n563), .Z(
        n560) );
  AND U592 ( .A(n133), .B(n564), .Z(n563) );
  XOR U593 ( .A(n565), .B(n566), .Z(n558) );
  AND U594 ( .A(n137), .B(n557), .Z(n566) );
  XNOR U595 ( .A(n567), .B(n555), .Z(n557) );
  XOR U596 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n568), .Z(n555) );
  AND U597 ( .A(n150), .B(n569), .Z(n568) );
  IV U598 ( .A(n565), .Z(n567) );
  XOR U599 ( .A(n570), .B(n571), .Z(n565) );
  AND U600 ( .A(n145), .B(n564), .Z(n571) );
  XOR U601 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n570), .Z(
        n564) );
  XOR U602 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(n572), .Z(
        n570) );
  AND U603 ( .A(n147), .B(n569), .Z(n572) );
  XOR U604 ( .A(\knn_comb_/min_val_out[0][1] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n569) );
  XOR U605 ( .A(n99), .B(n573), .Z(o[19]) );
  AND U606 ( .A(n122), .B(n574), .Z(n99) );
  XOR U607 ( .A(n100), .B(n573), .Z(n574) );
  XOR U608 ( .A(n575), .B(n576), .Z(n573) );
  AND U609 ( .A(n141), .B(n577), .Z(n576) );
  XOR U610 ( .A(n578), .B(n29), .Z(n100) );
  AND U611 ( .A(n125), .B(n579), .Z(n29) );
  XOR U612 ( .A(n30), .B(n578), .Z(n579) );
  XOR U613 ( .A(n580), .B(n581), .Z(n30) );
  AND U614 ( .A(n130), .B(n582), .Z(n581) );
  XOR U615 ( .A(p_input[19]), .B(n580), .Z(n582) );
  XOR U616 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ), .B(n583), .Z(
        n580) );
  AND U617 ( .A(n133), .B(n584), .Z(n583) );
  XOR U618 ( .A(n585), .B(n586), .Z(n578) );
  AND U619 ( .A(n137), .B(n577), .Z(n586) );
  XNOR U620 ( .A(n587), .B(n575), .Z(n577) );
  XOR U621 ( .A(\knn_comb_/min_val_out[0][19] ), .B(n588), .Z(n575) );
  AND U622 ( .A(n150), .B(n589), .Z(n588) );
  IV U623 ( .A(n585), .Z(n587) );
  XOR U624 ( .A(n590), .B(n591), .Z(n585) );
  AND U625 ( .A(n145), .B(n584), .Z(n591) );
  XOR U626 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ), .B(n590), .Z(
        n584) );
  XOR U627 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .B(n592), .Z(
        n590) );
  AND U628 ( .A(n147), .B(n589), .Z(n592) );
  XOR U629 ( .A(\knn_comb_/min_val_out[0][19] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .Z(n589) );
  XOR U630 ( .A(n101), .B(n593), .Z(o[18]) );
  AND U631 ( .A(n122), .B(n594), .Z(n101) );
  XOR U632 ( .A(n102), .B(n593), .Z(n594) );
  XOR U633 ( .A(n595), .B(n596), .Z(n593) );
  AND U634 ( .A(n141), .B(n597), .Z(n596) );
  XOR U635 ( .A(n598), .B(n31), .Z(n102) );
  AND U636 ( .A(n125), .B(n599), .Z(n31) );
  XOR U637 ( .A(n32), .B(n598), .Z(n599) );
  XOR U638 ( .A(n600), .B(n601), .Z(n32) );
  AND U639 ( .A(n130), .B(n602), .Z(n601) );
  XOR U640 ( .A(p_input[18]), .B(n600), .Z(n602) );
  XOR U641 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ), .B(n603), .Z(
        n600) );
  AND U642 ( .A(n133), .B(n604), .Z(n603) );
  XOR U643 ( .A(n605), .B(n606), .Z(n598) );
  AND U644 ( .A(n137), .B(n597), .Z(n606) );
  XNOR U645 ( .A(n607), .B(n595), .Z(n597) );
  XOR U646 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n608), .Z(n595) );
  AND U647 ( .A(n150), .B(n609), .Z(n608) );
  IV U648 ( .A(n605), .Z(n607) );
  XOR U649 ( .A(n610), .B(n611), .Z(n605) );
  AND U650 ( .A(n145), .B(n604), .Z(n611) );
  XOR U651 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ), .B(n610), .Z(
        n604) );
  XOR U652 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .B(n612), .Z(
        n610) );
  AND U653 ( .A(n147), .B(n609), .Z(n612) );
  XOR U654 ( .A(\knn_comb_/min_val_out[0][18] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .Z(n609) );
  XOR U655 ( .A(n105), .B(n613), .Z(o[17]) );
  AND U656 ( .A(n122), .B(n614), .Z(n105) );
  XOR U657 ( .A(n106), .B(n613), .Z(n614) );
  XOR U658 ( .A(n615), .B(n616), .Z(n613) );
  AND U659 ( .A(n141), .B(n617), .Z(n616) );
  XOR U660 ( .A(n618), .B(n33), .Z(n106) );
  AND U661 ( .A(n125), .B(n619), .Z(n33) );
  XOR U662 ( .A(n34), .B(n618), .Z(n619) );
  XOR U663 ( .A(n620), .B(n621), .Z(n34) );
  AND U664 ( .A(n130), .B(n622), .Z(n621) );
  XOR U665 ( .A(p_input[17]), .B(n620), .Z(n622) );
  XOR U666 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ), .B(n623), .Z(
        n620) );
  AND U667 ( .A(n133), .B(n624), .Z(n623) );
  XOR U668 ( .A(n625), .B(n626), .Z(n618) );
  AND U669 ( .A(n137), .B(n617), .Z(n626) );
  XNOR U670 ( .A(n627), .B(n615), .Z(n617) );
  XOR U671 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n628), .Z(n615) );
  AND U672 ( .A(n150), .B(n629), .Z(n628) );
  IV U673 ( .A(n625), .Z(n627) );
  XOR U674 ( .A(n630), .B(n631), .Z(n625) );
  AND U675 ( .A(n145), .B(n624), .Z(n631) );
  XOR U676 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ), .B(n630), .Z(
        n624) );
  XOR U677 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .B(n632), .Z(
        n630) );
  AND U678 ( .A(n147), .B(n629), .Z(n632) );
  XOR U679 ( .A(\knn_comb_/min_val_out[0][17] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .Z(n629) );
  XOR U680 ( .A(n107), .B(n633), .Z(o[16]) );
  AND U681 ( .A(n122), .B(n634), .Z(n107) );
  XOR U682 ( .A(n108), .B(n633), .Z(n634) );
  XOR U683 ( .A(n635), .B(n636), .Z(n633) );
  AND U684 ( .A(n141), .B(n637), .Z(n636) );
  XOR U685 ( .A(n638), .B(n35), .Z(n108) );
  AND U686 ( .A(n125), .B(n639), .Z(n35) );
  XOR U687 ( .A(n36), .B(n638), .Z(n639) );
  XOR U688 ( .A(n640), .B(n641), .Z(n36) );
  AND U689 ( .A(n130), .B(n642), .Z(n641) );
  XOR U690 ( .A(p_input[16]), .B(n640), .Z(n642) );
  XOR U691 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ), .B(n643), .Z(
        n640) );
  AND U692 ( .A(n133), .B(n644), .Z(n643) );
  XOR U693 ( .A(n645), .B(n646), .Z(n638) );
  AND U694 ( .A(n137), .B(n637), .Z(n646) );
  XNOR U695 ( .A(n647), .B(n635), .Z(n637) );
  XOR U696 ( .A(\knn_comb_/min_val_out[0][16] ), .B(n648), .Z(n635) );
  AND U697 ( .A(n150), .B(n649), .Z(n648) );
  IV U698 ( .A(n645), .Z(n647) );
  XOR U699 ( .A(n650), .B(n651), .Z(n645) );
  AND U700 ( .A(n145), .B(n644), .Z(n651) );
  XOR U701 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ), .B(n650), .Z(
        n644) );
  XOR U702 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .B(n652), .Z(
        n650) );
  AND U703 ( .A(n147), .B(n649), .Z(n652) );
  XOR U704 ( .A(n653), .B(n654), .Z(n649) );
  IV U705 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .Z(n654) );
  IV U706 ( .A(\knn_comb_/min_val_out[0][16] ), .Z(n653) );
  XOR U707 ( .A(n109), .B(n655), .Z(o[15]) );
  AND U708 ( .A(n122), .B(n656), .Z(n109) );
  XOR U709 ( .A(n110), .B(n655), .Z(n656) );
  XOR U710 ( .A(n657), .B(n658), .Z(n655) );
  AND U711 ( .A(n141), .B(n659), .Z(n658) );
  XOR U712 ( .A(n660), .B(n39), .Z(n110) );
  AND U713 ( .A(n125), .B(n661), .Z(n39) );
  XOR U714 ( .A(n40), .B(n660), .Z(n661) );
  XOR U715 ( .A(n662), .B(n663), .Z(n40) );
  AND U716 ( .A(n130), .B(n664), .Z(n663) );
  XOR U717 ( .A(p_input[15]), .B(n662), .Z(n664) );
  XOR U718 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n665), .Z(
        n662) );
  AND U719 ( .A(n133), .B(n666), .Z(n665) );
  XOR U720 ( .A(n667), .B(n668), .Z(n660) );
  AND U721 ( .A(n137), .B(n659), .Z(n668) );
  XNOR U722 ( .A(n669), .B(n657), .Z(n659) );
  XOR U723 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n670), .Z(n657) );
  AND U724 ( .A(n150), .B(n671), .Z(n670) );
  IV U725 ( .A(n667), .Z(n669) );
  XOR U726 ( .A(n672), .B(n673), .Z(n667) );
  AND U727 ( .A(n145), .B(n666), .Z(n673) );
  XOR U728 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n672), .Z(
        n666) );
  XOR U729 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n674), .Z(
        n672) );
  AND U730 ( .A(n147), .B(n671), .Z(n674) );
  XOR U731 ( .A(n675), .B(n676), .Z(n671) );
  IV U732 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n676) );
  IV U733 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n675) );
  XOR U734 ( .A(n111), .B(n677), .Z(o[14]) );
  AND U735 ( .A(n122), .B(n678), .Z(n111) );
  XOR U736 ( .A(n112), .B(n677), .Z(n678) );
  XOR U737 ( .A(n679), .B(n680), .Z(n677) );
  AND U738 ( .A(n141), .B(n681), .Z(n680) );
  XOR U739 ( .A(n682), .B(n41), .Z(n112) );
  AND U740 ( .A(n125), .B(n683), .Z(n41) );
  XOR U741 ( .A(n42), .B(n682), .Z(n683) );
  XOR U742 ( .A(n684), .B(n685), .Z(n42) );
  AND U743 ( .A(n130), .B(n686), .Z(n685) );
  XOR U744 ( .A(p_input[14]), .B(n684), .Z(n686) );
  XOR U745 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n687), .Z(
        n684) );
  AND U746 ( .A(n133), .B(n688), .Z(n687) );
  XOR U747 ( .A(n689), .B(n690), .Z(n682) );
  AND U748 ( .A(n137), .B(n681), .Z(n690) );
  XNOR U749 ( .A(n691), .B(n679), .Z(n681) );
  XOR U750 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n692), .Z(n679) );
  AND U751 ( .A(n150), .B(n693), .Z(n692) );
  IV U752 ( .A(n689), .Z(n691) );
  XOR U753 ( .A(n694), .B(n695), .Z(n689) );
  AND U754 ( .A(n145), .B(n688), .Z(n695) );
  XOR U755 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n694), .Z(
        n688) );
  XOR U756 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n696), .Z(
        n694) );
  AND U757 ( .A(n147), .B(n693), .Z(n696) );
  XOR U758 ( .A(\knn_comb_/min_val_out[0][14] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n693) );
  XOR U759 ( .A(n113), .B(n697), .Z(o[13]) );
  AND U760 ( .A(n122), .B(n698), .Z(n113) );
  XOR U761 ( .A(n114), .B(n697), .Z(n698) );
  XOR U762 ( .A(n699), .B(n700), .Z(n697) );
  AND U763 ( .A(n141), .B(n701), .Z(n700) );
  XOR U764 ( .A(n702), .B(n43), .Z(n114) );
  AND U765 ( .A(n125), .B(n703), .Z(n43) );
  XOR U766 ( .A(n44), .B(n702), .Z(n703) );
  XOR U767 ( .A(n704), .B(n705), .Z(n44) );
  AND U768 ( .A(n130), .B(n706), .Z(n705) );
  XOR U769 ( .A(p_input[13]), .B(n704), .Z(n706) );
  XOR U770 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n707), .Z(
        n704) );
  AND U771 ( .A(n133), .B(n708), .Z(n707) );
  XOR U772 ( .A(n709), .B(n710), .Z(n702) );
  AND U773 ( .A(n137), .B(n701), .Z(n710) );
  XNOR U774 ( .A(n711), .B(n699), .Z(n701) );
  XOR U775 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n712), .Z(n699) );
  AND U776 ( .A(n150), .B(n713), .Z(n712) );
  IV U777 ( .A(n709), .Z(n711) );
  XOR U778 ( .A(n714), .B(n715), .Z(n709) );
  AND U779 ( .A(n145), .B(n708), .Z(n715) );
  XOR U780 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n714), .Z(
        n708) );
  XOR U781 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(n716), .Z(
        n714) );
  AND U782 ( .A(n147), .B(n713), .Z(n716) );
  XOR U783 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n713) );
  XOR U784 ( .A(n115), .B(n717), .Z(o[12]) );
  AND U785 ( .A(n122), .B(n718), .Z(n115) );
  XOR U786 ( .A(n116), .B(n717), .Z(n718) );
  XOR U787 ( .A(n719), .B(n720), .Z(n717) );
  AND U788 ( .A(n141), .B(n721), .Z(n720) );
  XOR U789 ( .A(n722), .B(n45), .Z(n116) );
  AND U790 ( .A(n125), .B(n723), .Z(n45) );
  XOR U791 ( .A(n46), .B(n722), .Z(n723) );
  XOR U792 ( .A(n724), .B(n725), .Z(n46) );
  AND U793 ( .A(n130), .B(n726), .Z(n725) );
  XOR U794 ( .A(p_input[12]), .B(n724), .Z(n726) );
  XOR U795 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n727), .Z(
        n724) );
  AND U796 ( .A(n133), .B(n728), .Z(n727) );
  XOR U797 ( .A(n729), .B(n730), .Z(n722) );
  AND U798 ( .A(n137), .B(n721), .Z(n730) );
  XNOR U799 ( .A(n731), .B(n719), .Z(n721) );
  XOR U800 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n732), .Z(n719) );
  AND U801 ( .A(n150), .B(n733), .Z(n732) );
  IV U802 ( .A(n729), .Z(n731) );
  XOR U803 ( .A(n734), .B(n735), .Z(n729) );
  AND U804 ( .A(n145), .B(n728), .Z(n735) );
  XOR U805 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n734), .Z(
        n728) );
  XOR U806 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n736), .Z(
        n734) );
  AND U807 ( .A(n147), .B(n733), .Z(n736) );
  XOR U808 ( .A(n737), .B(n738), .Z(n733) );
  IV U809 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n738) );
  IV U810 ( .A(\knn_comb_/min_val_out[0][12] ), .Z(n737) );
  XOR U811 ( .A(n117), .B(n739), .Z(o[11]) );
  AND U812 ( .A(n122), .B(n740), .Z(n117) );
  XOR U813 ( .A(n118), .B(n739), .Z(n740) );
  XOR U814 ( .A(n741), .B(n742), .Z(n739) );
  AND U815 ( .A(n141), .B(n743), .Z(n742) );
  XOR U816 ( .A(n744), .B(n47), .Z(n118) );
  AND U817 ( .A(n125), .B(n745), .Z(n47) );
  XOR U818 ( .A(n48), .B(n744), .Z(n745) );
  XOR U819 ( .A(n746), .B(n747), .Z(n48) );
  AND U820 ( .A(n130), .B(n748), .Z(n747) );
  XOR U821 ( .A(p_input[11]), .B(n746), .Z(n748) );
  XOR U822 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n749), .Z(
        n746) );
  AND U823 ( .A(n133), .B(n750), .Z(n749) );
  XOR U824 ( .A(n751), .B(n752), .Z(n744) );
  AND U825 ( .A(n137), .B(n743), .Z(n752) );
  XNOR U826 ( .A(n753), .B(n741), .Z(n743) );
  XOR U827 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n754), .Z(n741) );
  AND U828 ( .A(n150), .B(n755), .Z(n754) );
  IV U829 ( .A(n751), .Z(n753) );
  XOR U830 ( .A(n756), .B(n757), .Z(n751) );
  AND U831 ( .A(n145), .B(n750), .Z(n757) );
  XOR U832 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n756), .Z(
        n750) );
  XOR U833 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n758), .Z(
        n756) );
  AND U834 ( .A(n147), .B(n755), .Z(n758) );
  XOR U835 ( .A(\knn_comb_/min_val_out[0][11] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n755) );
  XOR U836 ( .A(n119), .B(n759), .Z(o[10]) );
  AND U837 ( .A(n122), .B(n760), .Z(n119) );
  XOR U838 ( .A(n120), .B(n759), .Z(n760) );
  XOR U839 ( .A(n761), .B(n762), .Z(n759) );
  AND U840 ( .A(n141), .B(n763), .Z(n762) );
  XOR U841 ( .A(n764), .B(n49), .Z(n120) );
  AND U842 ( .A(n125), .B(n765), .Z(n49) );
  XOR U843 ( .A(n50), .B(n764), .Z(n765) );
  XOR U844 ( .A(n766), .B(n767), .Z(n50) );
  AND U845 ( .A(n130), .B(n768), .Z(n767) );
  XOR U846 ( .A(p_input[10]), .B(n766), .Z(n768) );
  XOR U847 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n769), .Z(
        n766) );
  AND U848 ( .A(n133), .B(n770), .Z(n769) );
  XOR U849 ( .A(n771), .B(n772), .Z(n764) );
  AND U850 ( .A(n137), .B(n763), .Z(n772) );
  XNOR U851 ( .A(n773), .B(n761), .Z(n763) );
  XOR U852 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n774), .Z(n761) );
  AND U853 ( .A(n150), .B(n775), .Z(n774) );
  IV U854 ( .A(n771), .Z(n773) );
  XOR U855 ( .A(n776), .B(n777), .Z(n771) );
  AND U856 ( .A(n145), .B(n770), .Z(n777) );
  XOR U857 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n776), .Z(
        n770) );
  XOR U858 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(n778), .Z(
        n776) );
  AND U859 ( .A(n147), .B(n775), .Z(n778) );
  XOR U860 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n775) );
  XOR U861 ( .A(n281), .B(n779), .Z(o[0]) );
  AND U862 ( .A(n122), .B(n780), .Z(n281) );
  XOR U863 ( .A(n282), .B(n779), .Z(n780) );
  XOR U864 ( .A(n781), .B(n782), .Z(n779) );
  AND U865 ( .A(n141), .B(n783), .Z(n782) );
  XOR U866 ( .A(n784), .B(n71), .Z(n282) );
  AND U867 ( .A(n125), .B(n785), .Z(n71) );
  XOR U868 ( .A(n72), .B(n784), .Z(n785) );
  XOR U869 ( .A(n786), .B(n787), .Z(n72) );
  AND U870 ( .A(n130), .B(n788), .Z(n787) );
  XOR U871 ( .A(p_input[0]), .B(n786), .Z(n788) );
  XOR U872 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n789), .Z(
        n786) );
  AND U873 ( .A(n133), .B(n790), .Z(n789) );
  XOR U874 ( .A(n791), .B(n792), .Z(n784) );
  AND U875 ( .A(n137), .B(n783), .Z(n792) );
  XNOR U876 ( .A(n793), .B(n781), .Z(n783) );
  XOR U877 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n794), .Z(n781) );
  AND U878 ( .A(n150), .B(n795), .Z(n794) );
  IV U879 ( .A(n791), .Z(n793) );
  XOR U880 ( .A(n796), .B(n797), .Z(n791) );
  AND U881 ( .A(n145), .B(n790), .Z(n797) );
  XOR U882 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n796), .Z(
        n790) );
  XOR U883 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(n798), .Z(
        n796) );
  AND U884 ( .A(n147), .B(n795), .Z(n798) );
  XOR U885 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n795) );
  XNOR U886 ( .A(n799), .B(n800), .Z(n122) );
  NOR U887 ( .A(n801), .B(n802), .Z(n800) );
  XOR U888 ( .A(n803), .B(n799), .Z(n802) );
  AND U889 ( .A(n804), .B(n805), .Z(n803) );
  NOR U890 ( .A(n799), .B(n806), .Z(n801) );
  NOR U891 ( .A(n807), .B(n808), .Z(n806) );
  IV U892 ( .A(n809), .Z(n807) );
  XOR U893 ( .A(n810), .B(n811), .Z(n799) );
  AND U894 ( .A(n812), .B(n813), .Z(n811) );
  XNOR U895 ( .A(n814), .B(n810), .Z(n813) );
  XNOR U896 ( .A(n815), .B(n816), .Z(n814) );
  AND U897 ( .A(n125), .B(n817), .Z(n816) );
  XNOR U898 ( .A(n815), .B(n818), .Z(n817) );
  XNOR U899 ( .A(n810), .B(n819), .Z(n812) );
  XOR U900 ( .A(n820), .B(n821), .Z(n819) );
  AND U901 ( .A(n141), .B(n822), .Z(n821) );
  XOR U902 ( .A(n823), .B(n824), .Z(n810) );
  AND U903 ( .A(n825), .B(n826), .Z(n824) );
  XOR U904 ( .A(n827), .B(n823), .Z(n826) );
  XNOR U905 ( .A(n828), .B(n829), .Z(n827) );
  AND U906 ( .A(n125), .B(n830), .Z(n829) );
  XNOR U907 ( .A(n831), .B(n828), .Z(n830) );
  XNOR U908 ( .A(n823), .B(n832), .Z(n825) );
  XOR U909 ( .A(n833), .B(n834), .Z(n832) );
  AND U910 ( .A(n141), .B(n835), .Z(n834) );
  XOR U911 ( .A(n836), .B(n837), .Z(n823) );
  AND U912 ( .A(n838), .B(n839), .Z(n837) );
  XOR U913 ( .A(n840), .B(n836), .Z(n839) );
  XNOR U914 ( .A(n841), .B(n842), .Z(n840) );
  AND U915 ( .A(n125), .B(n843), .Z(n842) );
  XNOR U916 ( .A(n844), .B(n841), .Z(n843) );
  XNOR U917 ( .A(n836), .B(n845), .Z(n838) );
  XOR U918 ( .A(n846), .B(n847), .Z(n845) );
  AND U919 ( .A(n141), .B(n848), .Z(n847) );
  XOR U920 ( .A(n849), .B(n850), .Z(n836) );
  AND U921 ( .A(n851), .B(n852), .Z(n850) );
  XOR U922 ( .A(n849), .B(n853), .Z(n852) );
  XOR U923 ( .A(n854), .B(n855), .Z(n853) );
  AND U924 ( .A(n125), .B(n856), .Z(n855) );
  XOR U925 ( .A(n857), .B(n854), .Z(n856) );
  XNOR U926 ( .A(n858), .B(n849), .Z(n851) );
  XNOR U927 ( .A(n859), .B(n860), .Z(n858) );
  AND U928 ( .A(n141), .B(n861), .Z(n860) );
  AND U929 ( .A(n862), .B(n863), .Z(n849) );
  XNOR U930 ( .A(n864), .B(n865), .Z(n863) );
  AND U931 ( .A(n125), .B(n866), .Z(n865) );
  XNOR U932 ( .A(n867), .B(n864), .Z(n866) );
  XNOR U933 ( .A(n868), .B(n869), .Z(n125) );
  NOR U934 ( .A(n870), .B(n871), .Z(n869) );
  XNOR U935 ( .A(n868), .B(n808), .Z(n871) );
  NOR U936 ( .A(n804), .B(n805), .Z(n808) );
  NOR U937 ( .A(n868), .B(n809), .Z(n870) );
  AND U938 ( .A(n872), .B(n873), .Z(n809) );
  IV U939 ( .A(n874), .Z(n872) );
  XOR U940 ( .A(n875), .B(n876), .Z(n868) );
  AND U941 ( .A(n877), .B(n878), .Z(n876) );
  XNOR U942 ( .A(n875), .B(n818), .Z(n878) );
  XOR U943 ( .A(n879), .B(n880), .Z(n818) );
  AND U944 ( .A(n130), .B(n881), .Z(n880) );
  XOR U945 ( .A(n882), .B(n879), .Z(n881) );
  XNOR U946 ( .A(n875), .B(n815), .Z(n877) );
  XNOR U947 ( .A(n883), .B(n884), .Z(n815) );
  AND U948 ( .A(n137), .B(n822), .Z(n884) );
  XOR U949 ( .A(n883), .B(n885), .Z(n822) );
  XOR U950 ( .A(n886), .B(n887), .Z(n875) );
  AND U951 ( .A(n888), .B(n889), .Z(n887) );
  XOR U952 ( .A(n831), .B(n886), .Z(n889) );
  XOR U953 ( .A(n890), .B(n891), .Z(n831) );
  AND U954 ( .A(n130), .B(n892), .Z(n891) );
  XNOR U955 ( .A(n893), .B(n890), .Z(n892) );
  XOR U956 ( .A(n886), .B(n828), .Z(n888) );
  XOR U957 ( .A(n894), .B(n895), .Z(n828) );
  AND U958 ( .A(n137), .B(n835), .Z(n895) );
  XOR U959 ( .A(n894), .B(n896), .Z(n835) );
  XOR U960 ( .A(n897), .B(n898), .Z(n886) );
  AND U961 ( .A(n899), .B(n900), .Z(n898) );
  XOR U962 ( .A(n844), .B(n897), .Z(n900) );
  XOR U963 ( .A(n901), .B(n902), .Z(n844) );
  AND U964 ( .A(n130), .B(n903), .Z(n902) );
  XOR U965 ( .A(n904), .B(n901), .Z(n903) );
  XOR U966 ( .A(n897), .B(n841), .Z(n899) );
  XOR U967 ( .A(n905), .B(n906), .Z(n841) );
  AND U968 ( .A(n137), .B(n848), .Z(n906) );
  XOR U969 ( .A(n905), .B(n907), .Z(n848) );
  XOR U970 ( .A(n908), .B(n909), .Z(n897) );
  AND U971 ( .A(n910), .B(n911), .Z(n909) );
  XOR U972 ( .A(n908), .B(n857), .Z(n911) );
  XOR U973 ( .A(n912), .B(n913), .Z(n857) );
  AND U974 ( .A(n130), .B(n914), .Z(n913) );
  XNOR U975 ( .A(n915), .B(n912), .Z(n914) );
  XNOR U976 ( .A(n854), .B(n908), .Z(n910) );
  XNOR U977 ( .A(n916), .B(n917), .Z(n854) );
  AND U978 ( .A(n137), .B(n861), .Z(n917) );
  XOR U979 ( .A(n916), .B(n859), .Z(n861) );
  AND U980 ( .A(n864), .B(n867), .Z(n908) );
  XOR U981 ( .A(n918), .B(n919), .Z(n867) );
  AND U982 ( .A(n130), .B(n920), .Z(n919) );
  XNOR U983 ( .A(n921), .B(n918), .Z(n920) );
  XNOR U984 ( .A(n922), .B(n923), .Z(n130) );
  NOR U985 ( .A(n924), .B(n925), .Z(n923) );
  XNOR U986 ( .A(n922), .B(n874), .Z(n925) );
  NOR U987 ( .A(n926), .B(n927), .Z(n874) );
  NOR U988 ( .A(n922), .B(n873), .Z(n924) );
  AND U989 ( .A(n882), .B(n928), .Z(n873) );
  XOR U990 ( .A(n929), .B(n930), .Z(n922) );
  AND U991 ( .A(n931), .B(n932), .Z(n930) );
  XNOR U992 ( .A(n929), .B(n882), .Z(n932) );
  XNOR U993 ( .A(n933), .B(n934), .Z(n882) );
  XOR U994 ( .A(n935), .B(n928), .Z(n934) );
  AND U995 ( .A(n893), .B(n936), .Z(n928) );
  AND U996 ( .A(n937), .B(n938), .Z(n935) );
  XOR U997 ( .A(n939), .B(n933), .Z(n937) );
  XOR U998 ( .A(n879), .B(n929), .Z(n931) );
  AND U999 ( .A(n940), .B(n941), .Z(n879) );
  XOR U1000 ( .A(n942), .B(n943), .Z(n929) );
  AND U1001 ( .A(n944), .B(n945), .Z(n943) );
  XNOR U1002 ( .A(n942), .B(n893), .Z(n945) );
  XOR U1003 ( .A(n946), .B(n938), .Z(n893) );
  XNOR U1004 ( .A(n947), .B(n933), .Z(n938) );
  XOR U1005 ( .A(n948), .B(n949), .Z(n933) );
  AND U1006 ( .A(n950), .B(n951), .Z(n949) );
  XOR U1007 ( .A(n952), .B(n948), .Z(n950) );
  XNOR U1008 ( .A(n953), .B(n954), .Z(n947) );
  AND U1009 ( .A(n955), .B(n956), .Z(n954) );
  XOR U1010 ( .A(n953), .B(n957), .Z(n955) );
  XNOR U1011 ( .A(n939), .B(n936), .Z(n946) );
  AND U1012 ( .A(n958), .B(n959), .Z(n936) );
  XOR U1013 ( .A(n960), .B(n961), .Z(n939) );
  AND U1014 ( .A(n962), .B(n963), .Z(n961) );
  XOR U1015 ( .A(n960), .B(n964), .Z(n962) );
  XNOR U1016 ( .A(n890), .B(n942), .Z(n944) );
  XNOR U1017 ( .A(n965), .B(n966), .Z(n890) );
  AND U1018 ( .A(n133), .B(n967), .Z(n966) );
  XOR U1019 ( .A(n968), .B(n969), .Z(n942) );
  AND U1020 ( .A(n970), .B(n971), .Z(n969) );
  XNOR U1021 ( .A(n968), .B(n958), .Z(n971) );
  IV U1022 ( .A(n904), .Z(n958) );
  XNOR U1023 ( .A(n972), .B(n951), .Z(n904) );
  XNOR U1024 ( .A(n973), .B(n957), .Z(n951) );
  XOR U1025 ( .A(n974), .B(n975), .Z(n957) );
  AND U1026 ( .A(n976), .B(n977), .Z(n975) );
  XOR U1027 ( .A(n974), .B(n978), .Z(n976) );
  XNOR U1028 ( .A(n956), .B(n948), .Z(n973) );
  XOR U1029 ( .A(n979), .B(n980), .Z(n948) );
  AND U1030 ( .A(n981), .B(n982), .Z(n980) );
  XNOR U1031 ( .A(n983), .B(n979), .Z(n981) );
  XNOR U1032 ( .A(n984), .B(n953), .Z(n956) );
  XOR U1033 ( .A(n985), .B(n986), .Z(n953) );
  AND U1034 ( .A(n987), .B(n988), .Z(n986) );
  XOR U1035 ( .A(n985), .B(n989), .Z(n987) );
  XNOR U1036 ( .A(n990), .B(n991), .Z(n984) );
  AND U1037 ( .A(n992), .B(n993), .Z(n991) );
  XNOR U1038 ( .A(n990), .B(n994), .Z(n992) );
  XNOR U1039 ( .A(n952), .B(n959), .Z(n972) );
  AND U1040 ( .A(n915), .B(n995), .Z(n959) );
  XOR U1041 ( .A(n964), .B(n963), .Z(n952) );
  XNOR U1042 ( .A(n996), .B(n960), .Z(n963) );
  XOR U1043 ( .A(n997), .B(n998), .Z(n960) );
  AND U1044 ( .A(n999), .B(n1000), .Z(n998) );
  XOR U1045 ( .A(n997), .B(n1001), .Z(n999) );
  XNOR U1046 ( .A(n1002), .B(n1003), .Z(n996) );
  AND U1047 ( .A(n1004), .B(n1005), .Z(n1003) );
  XOR U1048 ( .A(n1002), .B(n1006), .Z(n1004) );
  XOR U1049 ( .A(n1007), .B(n1008), .Z(n964) );
  AND U1050 ( .A(n1009), .B(n1010), .Z(n1008) );
  XOR U1051 ( .A(n1007), .B(n1011), .Z(n1009) );
  XNOR U1052 ( .A(n901), .B(n968), .Z(n970) );
  XNOR U1053 ( .A(n1012), .B(n1013), .Z(n901) );
  AND U1054 ( .A(n133), .B(n1014), .Z(n1013) );
  XNOR U1055 ( .A(n1015), .B(n1016), .Z(n1014) );
  XOR U1056 ( .A(n1017), .B(n1018), .Z(n968) );
  AND U1057 ( .A(n1019), .B(n1020), .Z(n1018) );
  XNOR U1058 ( .A(n1017), .B(n915), .Z(n1020) );
  XOR U1059 ( .A(n1021), .B(n982), .Z(n915) );
  XNOR U1060 ( .A(n1022), .B(n989), .Z(n982) );
  XOR U1061 ( .A(n978), .B(n977), .Z(n989) );
  XNOR U1062 ( .A(n1023), .B(n974), .Z(n977) );
  XOR U1063 ( .A(n1024), .B(n1025), .Z(n974) );
  AND U1064 ( .A(n1026), .B(n1027), .Z(n1025) );
  XOR U1065 ( .A(n1024), .B(n1028), .Z(n1026) );
  XNOR U1066 ( .A(n1029), .B(n1030), .Z(n1023) );
  NOR U1067 ( .A(n1031), .B(n1032), .Z(n1030) );
  XNOR U1068 ( .A(n1029), .B(n1033), .Z(n1031) );
  XOR U1069 ( .A(n1034), .B(n1035), .Z(n978) );
  NOR U1070 ( .A(n1036), .B(n1037), .Z(n1035) );
  XNOR U1071 ( .A(n1034), .B(n1038), .Z(n1036) );
  XNOR U1072 ( .A(n988), .B(n979), .Z(n1022) );
  XOR U1073 ( .A(n1039), .B(n1040), .Z(n979) );
  NOR U1074 ( .A(n1041), .B(n1042), .Z(n1040) );
  XNOR U1075 ( .A(n1039), .B(n1043), .Z(n1041) );
  XOR U1076 ( .A(n1044), .B(n994), .Z(n988) );
  XNOR U1077 ( .A(n1045), .B(n1046), .Z(n994) );
  NOR U1078 ( .A(n1047), .B(n1048), .Z(n1046) );
  XNOR U1079 ( .A(n1045), .B(n1049), .Z(n1047) );
  XNOR U1080 ( .A(n993), .B(n985), .Z(n1044) );
  XOR U1081 ( .A(n1050), .B(n1051), .Z(n985) );
  AND U1082 ( .A(n1052), .B(n1053), .Z(n1051) );
  XOR U1083 ( .A(n1050), .B(n1054), .Z(n1052) );
  XNOR U1084 ( .A(n1055), .B(n990), .Z(n993) );
  XOR U1085 ( .A(n1056), .B(n1057), .Z(n990) );
  AND U1086 ( .A(n1058), .B(n1059), .Z(n1057) );
  XOR U1087 ( .A(n1056), .B(n1060), .Z(n1058) );
  XNOR U1088 ( .A(n1061), .B(n1062), .Z(n1055) );
  NOR U1089 ( .A(n1063), .B(n1064), .Z(n1062) );
  XOR U1090 ( .A(n1061), .B(n1065), .Z(n1063) );
  XOR U1091 ( .A(n983), .B(n995), .Z(n1021) );
  AND U1092 ( .A(n921), .B(n1066), .Z(n995) );
  XNOR U1093 ( .A(n1001), .B(n1000), .Z(n983) );
  XNOR U1094 ( .A(n1067), .B(n1006), .Z(n1000) );
  XOR U1095 ( .A(n1068), .B(n1069), .Z(n1006) );
  NOR U1096 ( .A(n1070), .B(n1071), .Z(n1069) );
  XNOR U1097 ( .A(n1068), .B(n1072), .Z(n1070) );
  XNOR U1098 ( .A(n1005), .B(n997), .Z(n1067) );
  XOR U1099 ( .A(n1073), .B(n1074), .Z(n997) );
  AND U1100 ( .A(n1075), .B(n1076), .Z(n1074) );
  XNOR U1101 ( .A(n1073), .B(n1077), .Z(n1075) );
  XNOR U1102 ( .A(n1078), .B(n1002), .Z(n1005) );
  XOR U1103 ( .A(n1079), .B(n1080), .Z(n1002) );
  AND U1104 ( .A(n1081), .B(n1082), .Z(n1080) );
  XOR U1105 ( .A(n1079), .B(n1083), .Z(n1081) );
  XNOR U1106 ( .A(n1084), .B(n1085), .Z(n1078) );
  NOR U1107 ( .A(n1086), .B(n1087), .Z(n1085) );
  XOR U1108 ( .A(n1084), .B(n1088), .Z(n1086) );
  XOR U1109 ( .A(n1011), .B(n1010), .Z(n1001) );
  XNOR U1110 ( .A(n1089), .B(n1007), .Z(n1010) );
  XOR U1111 ( .A(n1090), .B(n1091), .Z(n1007) );
  AND U1112 ( .A(n1092), .B(n1093), .Z(n1091) );
  XOR U1113 ( .A(n1090), .B(n1094), .Z(n1092) );
  XNOR U1114 ( .A(n1095), .B(n1096), .Z(n1089) );
  NOR U1115 ( .A(n1097), .B(n1098), .Z(n1096) );
  XNOR U1116 ( .A(n1095), .B(n1099), .Z(n1097) );
  XOR U1117 ( .A(n1100), .B(n1101), .Z(n1011) );
  NOR U1118 ( .A(n1102), .B(n1103), .Z(n1101) );
  XNOR U1119 ( .A(n1100), .B(n1104), .Z(n1102) );
  XNOR U1120 ( .A(n912), .B(n1017), .Z(n1019) );
  XNOR U1121 ( .A(n1105), .B(n1106), .Z(n912) );
  AND U1122 ( .A(n133), .B(n1107), .Z(n1106) );
  NOR U1123 ( .A(n918), .B(n921), .Z(n1017) );
  XOR U1124 ( .A(n1108), .B(n1066), .Z(n921) );
  XOR U1125 ( .A(p_input[0]), .B(p_input[128]), .Z(n1066) );
  XOR U1126 ( .A(n1043), .B(n1042), .Z(n1108) );
  XOR U1127 ( .A(n1109), .B(n1054), .Z(n1042) );
  XOR U1128 ( .A(n1028), .B(n1027), .Z(n1054) );
  XNOR U1129 ( .A(n1110), .B(n1033), .Z(n1027) );
  XOR U1130 ( .A(p_input[152]), .B(p_input[24]), .Z(n1033) );
  XOR U1131 ( .A(n1024), .B(n1032), .Z(n1110) );
  XOR U1132 ( .A(n1111), .B(n1029), .Z(n1032) );
  XOR U1133 ( .A(p_input[150]), .B(p_input[22]), .Z(n1029) );
  XNOR U1134 ( .A(p_input[151]), .B(p_input[23]), .Z(n1111) );
  XOR U1135 ( .A(p_input[146]), .B(p_input[18]), .Z(n1024) );
  XNOR U1136 ( .A(n1038), .B(n1037), .Z(n1028) );
  XOR U1137 ( .A(n1112), .B(n1034), .Z(n1037) );
  XOR U1138 ( .A(p_input[147]), .B(p_input[19]), .Z(n1034) );
  XNOR U1139 ( .A(p_input[148]), .B(p_input[20]), .Z(n1112) );
  XOR U1140 ( .A(p_input[149]), .B(p_input[21]), .Z(n1038) );
  XNOR U1141 ( .A(n1053), .B(n1039), .Z(n1109) );
  XOR U1142 ( .A(p_input[129]), .B(p_input[1]), .Z(n1039) );
  XNOR U1143 ( .A(n1113), .B(n1060), .Z(n1053) );
  XNOR U1144 ( .A(n1049), .B(n1048), .Z(n1060) );
  XOR U1145 ( .A(n1114), .B(n1045), .Z(n1048) );
  XOR U1146 ( .A(p_input[154]), .B(p_input[26]), .Z(n1045) );
  XNOR U1147 ( .A(p_input[155]), .B(p_input[27]), .Z(n1114) );
  XOR U1148 ( .A(p_input[156]), .B(p_input[28]), .Z(n1049) );
  XNOR U1149 ( .A(n1059), .B(n1050), .Z(n1113) );
  XOR U1150 ( .A(p_input[145]), .B(p_input[17]), .Z(n1050) );
  XOR U1151 ( .A(n1115), .B(n1065), .Z(n1059) );
  XNOR U1152 ( .A(p_input[159]), .B(p_input[31]), .Z(n1065) );
  XOR U1153 ( .A(n1056), .B(n1064), .Z(n1115) );
  XOR U1154 ( .A(n1116), .B(n1061), .Z(n1064) );
  XOR U1155 ( .A(p_input[157]), .B(p_input[29]), .Z(n1061) );
  XNOR U1156 ( .A(p_input[158]), .B(p_input[30]), .Z(n1116) );
  XOR U1157 ( .A(p_input[153]), .B(p_input[25]), .Z(n1056) );
  XNOR U1158 ( .A(n1077), .B(n1076), .Z(n1043) );
  XNOR U1159 ( .A(n1117), .B(n1083), .Z(n1076) );
  XNOR U1160 ( .A(n1072), .B(n1071), .Z(n1083) );
  XOR U1161 ( .A(n1118), .B(n1068), .Z(n1071) );
  XOR U1162 ( .A(p_input[11]), .B(p_input[139]), .Z(n1068) );
  XNOR U1163 ( .A(p_input[12]), .B(p_input[140]), .Z(n1118) );
  XOR U1164 ( .A(p_input[13]), .B(p_input[141]), .Z(n1072) );
  XNOR U1165 ( .A(n1082), .B(n1073), .Z(n1117) );
  XOR U1166 ( .A(p_input[130]), .B(p_input[2]), .Z(n1073) );
  XOR U1167 ( .A(n1119), .B(n1088), .Z(n1082) );
  XNOR U1168 ( .A(p_input[144]), .B(p_input[16]), .Z(n1088) );
  XOR U1169 ( .A(n1079), .B(n1087), .Z(n1119) );
  XOR U1170 ( .A(n1120), .B(n1084), .Z(n1087) );
  XOR U1171 ( .A(p_input[142]), .B(p_input[14]), .Z(n1084) );
  XNOR U1172 ( .A(p_input[143]), .B(p_input[15]), .Z(n1120) );
  XOR U1173 ( .A(p_input[10]), .B(p_input[138]), .Z(n1079) );
  XNOR U1174 ( .A(n1094), .B(n1093), .Z(n1077) );
  XNOR U1175 ( .A(n1121), .B(n1099), .Z(n1093) );
  XOR U1176 ( .A(p_input[137]), .B(p_input[9]), .Z(n1099) );
  XOR U1177 ( .A(n1090), .B(n1098), .Z(n1121) );
  XOR U1178 ( .A(n1122), .B(n1095), .Z(n1098) );
  XOR U1179 ( .A(p_input[135]), .B(p_input[7]), .Z(n1095) );
  XNOR U1180 ( .A(p_input[136]), .B(p_input[8]), .Z(n1122) );
  XOR U1181 ( .A(p_input[131]), .B(p_input[3]), .Z(n1090) );
  XNOR U1182 ( .A(n1104), .B(n1103), .Z(n1094) );
  XOR U1183 ( .A(n1123), .B(n1100), .Z(n1103) );
  XOR U1184 ( .A(p_input[132]), .B(p_input[4]), .Z(n1100) );
  XNOR U1185 ( .A(p_input[133]), .B(p_input[5]), .Z(n1123) );
  XOR U1186 ( .A(p_input[134]), .B(p_input[6]), .Z(n1104) );
  XOR U1187 ( .A(n1124), .B(n1125), .Z(n918) );
  AND U1188 ( .A(n133), .B(n1126), .Z(n1125) );
  XNOR U1189 ( .A(n1127), .B(n1128), .Z(n133) );
  NOR U1190 ( .A(n1129), .B(n1130), .Z(n1128) );
  XOR U1191 ( .A(n1127), .B(n926), .Z(n1130) );
  XNOR U1192 ( .A(n1131), .B(n1132), .Z(n864) );
  AND U1193 ( .A(n137), .B(n1133), .Z(n1132) );
  XNOR U1194 ( .A(n1134), .B(n1135), .Z(n137) );
  NOR U1195 ( .A(n1136), .B(n1137), .Z(n1135) );
  XOR U1196 ( .A(n805), .B(n1134), .Z(n1137) );
  NOR U1197 ( .A(n1134), .B(n804), .Z(n1136) );
  XOR U1198 ( .A(n1138), .B(n1139), .Z(n1134) );
  AND U1199 ( .A(n1140), .B(n1141), .Z(n1139) );
  XNOR U1200 ( .A(n883), .B(n1138), .Z(n1141) );
  XOR U1201 ( .A(n1138), .B(n885), .Z(n1140) );
  XOR U1202 ( .A(n1142), .B(n1143), .Z(n1138) );
  AND U1203 ( .A(n1144), .B(n1145), .Z(n1143) );
  XNOR U1204 ( .A(n894), .B(n1142), .Z(n1145) );
  XOR U1205 ( .A(n1142), .B(n896), .Z(n1144) );
  IV U1206 ( .A(n833), .Z(n896) );
  XOR U1207 ( .A(n1146), .B(n1147), .Z(n1142) );
  AND U1208 ( .A(n1148), .B(n1149), .Z(n1147) );
  XOR U1209 ( .A(n1146), .B(n907), .Z(n1148) );
  XOR U1210 ( .A(n1150), .B(n1151), .Z(n862) );
  AND U1211 ( .A(n141), .B(n1133), .Z(n1151) );
  XNOR U1212 ( .A(n1131), .B(n1150), .Z(n1133) );
  XNOR U1213 ( .A(n1152), .B(n1153), .Z(n141) );
  NOR U1214 ( .A(n1154), .B(n1155), .Z(n1153) );
  XNOR U1215 ( .A(n805), .B(n1156), .Z(n1155) );
  IV U1216 ( .A(n1152), .Z(n1156) );
  AND U1217 ( .A(n1157), .B(n1158), .Z(n805) );
  NOR U1218 ( .A(n1152), .B(n804), .Z(n1154) );
  AND U1219 ( .A(n926), .B(n927), .Z(n804) );
  IV U1220 ( .A(n1159), .Z(n926) );
  XOR U1221 ( .A(n1160), .B(n1161), .Z(n1152) );
  AND U1222 ( .A(n1162), .B(n1163), .Z(n1161) );
  XNOR U1223 ( .A(n1160), .B(n883), .Z(n1163) );
  XOR U1224 ( .A(n940), .B(n1164), .Z(n883) );
  AND U1225 ( .A(n145), .B(n1165), .Z(n1164) );
  XOR U1226 ( .A(n941), .B(n940), .Z(n1165) );
  XNOR U1227 ( .A(n820), .B(n1160), .Z(n1162) );
  IV U1228 ( .A(n885), .Z(n820) );
  XOR U1229 ( .A(n1166), .B(n1167), .Z(n885) );
  AND U1230 ( .A(n150), .B(n1168), .Z(n1167) );
  XOR U1231 ( .A(n1169), .B(n1170), .Z(n1160) );
  AND U1232 ( .A(n1171), .B(n1172), .Z(n1170) );
  XNOR U1233 ( .A(n1169), .B(n894), .Z(n1172) );
  XOR U1234 ( .A(n1173), .B(n1174), .Z(n894) );
  AND U1235 ( .A(n145), .B(n967), .Z(n1174) );
  XOR U1236 ( .A(n965), .B(n1173), .Z(n967) );
  XNOR U1237 ( .A(n833), .B(n1169), .Z(n1171) );
  XNOR U1238 ( .A(n1175), .B(n1176), .Z(n833) );
  AND U1239 ( .A(n150), .B(n1177), .Z(n1176) );
  XOR U1240 ( .A(n1146), .B(n1178), .Z(n1169) );
  AND U1241 ( .A(n1179), .B(n1149), .Z(n1178) );
  XNOR U1242 ( .A(n905), .B(n1146), .Z(n1149) );
  XOR U1243 ( .A(n1016), .B(n1180), .Z(n905) );
  AND U1244 ( .A(n145), .B(n1181), .Z(n1180) );
  XOR U1245 ( .A(n1012), .B(n1016), .Z(n1181) );
  XNOR U1246 ( .A(n846), .B(n1146), .Z(n1179) );
  IV U1247 ( .A(n907), .Z(n846) );
  XOR U1248 ( .A(n1182), .B(n1183), .Z(n907) );
  AND U1249 ( .A(n150), .B(n1184), .Z(n1183) );
  XOR U1250 ( .A(n1185), .B(n1186), .Z(n1146) );
  AND U1251 ( .A(n1187), .B(n1188), .Z(n1186) );
  XNOR U1252 ( .A(n1185), .B(n916), .Z(n1188) );
  XNOR U1253 ( .A(n1189), .B(n1190), .Z(n916) );
  AND U1254 ( .A(n145), .B(n1107), .Z(n1190) );
  XOR U1255 ( .A(n1105), .B(n1191), .Z(n1107) );
  IV U1256 ( .A(n1189), .Z(n1191) );
  XNOR U1257 ( .A(n1192), .B(n1185), .Z(n1187) );
  IV U1258 ( .A(n859), .Z(n1192) );
  XOR U1259 ( .A(n1193), .B(n1194), .Z(n859) );
  AND U1260 ( .A(n150), .B(n1195), .Z(n1194) );
  AND U1261 ( .A(n1150), .B(n1131), .Z(n1185) );
  XNOR U1262 ( .A(n1196), .B(n1197), .Z(n1131) );
  AND U1263 ( .A(n145), .B(n1126), .Z(n1197) );
  XNOR U1264 ( .A(n1124), .B(n1196), .Z(n1126) );
  XNOR U1265 ( .A(n1127), .B(n1198), .Z(n145) );
  NOR U1266 ( .A(n1129), .B(n1199), .Z(n1198) );
  XNOR U1267 ( .A(n1127), .B(n1159), .Z(n1199) );
  NOR U1268 ( .A(n1157), .B(n1158), .Z(n1159) );
  NOR U1269 ( .A(n1127), .B(n927), .Z(n1129) );
  AND U1270 ( .A(n941), .B(n1200), .Z(n927) );
  XOR U1271 ( .A(n1201), .B(n1202), .Z(n1127) );
  AND U1272 ( .A(n1203), .B(n1204), .Z(n1202) );
  XNOR U1273 ( .A(n941), .B(n1201), .Z(n1204) );
  XNOR U1274 ( .A(n1205), .B(n1206), .Z(n941) );
  XOR U1275 ( .A(n1207), .B(n1200), .Z(n1206) );
  AND U1276 ( .A(n965), .B(n1208), .Z(n1200) );
  AND U1277 ( .A(n1209), .B(n1210), .Z(n1207) );
  XOR U1278 ( .A(n1211), .B(n1205), .Z(n1209) );
  XOR U1279 ( .A(n1201), .B(n940), .Z(n1203) );
  XOR U1280 ( .A(n1212), .B(n1213), .Z(n940) );
  AND U1281 ( .A(n147), .B(n1168), .Z(n1213) );
  XOR U1282 ( .A(n1212), .B(n1166), .Z(n1168) );
  XOR U1283 ( .A(n1214), .B(n1215), .Z(n1201) );
  AND U1284 ( .A(n1216), .B(n1217), .Z(n1215) );
  XNOR U1285 ( .A(n965), .B(n1214), .Z(n1217) );
  XOR U1286 ( .A(n1218), .B(n1210), .Z(n965) );
  XNOR U1287 ( .A(n1219), .B(n1205), .Z(n1210) );
  XOR U1288 ( .A(n1220), .B(n1221), .Z(n1205) );
  AND U1289 ( .A(n1222), .B(n1223), .Z(n1221) );
  XOR U1290 ( .A(n1224), .B(n1220), .Z(n1222) );
  XNOR U1291 ( .A(n1225), .B(n1226), .Z(n1219) );
  AND U1292 ( .A(n1227), .B(n1228), .Z(n1226) );
  XOR U1293 ( .A(n1225), .B(n1229), .Z(n1227) );
  XNOR U1294 ( .A(n1211), .B(n1208), .Z(n1218) );
  AND U1295 ( .A(n1012), .B(n1230), .Z(n1208) );
  XOR U1296 ( .A(n1231), .B(n1232), .Z(n1211) );
  AND U1297 ( .A(n1233), .B(n1234), .Z(n1232) );
  XOR U1298 ( .A(n1231), .B(n1235), .Z(n1233) );
  XOR U1299 ( .A(n1214), .B(n1173), .Z(n1216) );
  XOR U1300 ( .A(n1236), .B(n1237), .Z(n1173) );
  AND U1301 ( .A(n147), .B(n1177), .Z(n1237) );
  XOR U1302 ( .A(n1236), .B(n1175), .Z(n1177) );
  XOR U1303 ( .A(n1238), .B(n1239), .Z(n1214) );
  AND U1304 ( .A(n1240), .B(n1241), .Z(n1239) );
  XNOR U1305 ( .A(n1012), .B(n1238), .Z(n1241) );
  IV U1306 ( .A(n1015), .Z(n1012) );
  XNOR U1307 ( .A(n1242), .B(n1223), .Z(n1015) );
  XNOR U1308 ( .A(n1243), .B(n1229), .Z(n1223) );
  XOR U1309 ( .A(n1244), .B(n1245), .Z(n1229) );
  AND U1310 ( .A(n1246), .B(n1247), .Z(n1245) );
  XOR U1311 ( .A(n1244), .B(n1248), .Z(n1246) );
  XNOR U1312 ( .A(n1228), .B(n1220), .Z(n1243) );
  XOR U1313 ( .A(n1249), .B(n1250), .Z(n1220) );
  AND U1314 ( .A(n1251), .B(n1252), .Z(n1250) );
  XNOR U1315 ( .A(n1253), .B(n1249), .Z(n1251) );
  XNOR U1316 ( .A(n1254), .B(n1225), .Z(n1228) );
  XOR U1317 ( .A(n1255), .B(n1256), .Z(n1225) );
  AND U1318 ( .A(n1257), .B(n1258), .Z(n1256) );
  XOR U1319 ( .A(n1255), .B(n1259), .Z(n1257) );
  XNOR U1320 ( .A(n1260), .B(n1261), .Z(n1254) );
  AND U1321 ( .A(n1262), .B(n1263), .Z(n1261) );
  XNOR U1322 ( .A(n1260), .B(n1264), .Z(n1262) );
  XNOR U1323 ( .A(n1224), .B(n1230), .Z(n1242) );
  AND U1324 ( .A(n1105), .B(n1265), .Z(n1230) );
  XOR U1325 ( .A(n1235), .B(n1234), .Z(n1224) );
  XNOR U1326 ( .A(n1266), .B(n1231), .Z(n1234) );
  XOR U1327 ( .A(n1267), .B(n1268), .Z(n1231) );
  AND U1328 ( .A(n1269), .B(n1270), .Z(n1268) );
  XOR U1329 ( .A(n1267), .B(n1271), .Z(n1269) );
  XNOR U1330 ( .A(n1272), .B(n1273), .Z(n1266) );
  AND U1331 ( .A(n1274), .B(n1275), .Z(n1273) );
  XOR U1332 ( .A(n1272), .B(n1276), .Z(n1274) );
  XOR U1333 ( .A(n1277), .B(n1278), .Z(n1235) );
  AND U1334 ( .A(n1279), .B(n1280), .Z(n1278) );
  XOR U1335 ( .A(n1277), .B(n1281), .Z(n1279) );
  XOR U1336 ( .A(n1238), .B(n1016), .Z(n1240) );
  XOR U1337 ( .A(n1282), .B(n1283), .Z(n1016) );
  AND U1338 ( .A(n147), .B(n1184), .Z(n1283) );
  XOR U1339 ( .A(n1282), .B(n1182), .Z(n1184) );
  XOR U1340 ( .A(n1284), .B(n1285), .Z(n1238) );
  AND U1341 ( .A(n1286), .B(n1287), .Z(n1285) );
  XNOR U1342 ( .A(n1284), .B(n1105), .Z(n1287) );
  XOR U1343 ( .A(n1288), .B(n1252), .Z(n1105) );
  XNOR U1344 ( .A(n1289), .B(n1259), .Z(n1252) );
  XOR U1345 ( .A(n1248), .B(n1247), .Z(n1259) );
  XNOR U1346 ( .A(n1290), .B(n1244), .Z(n1247) );
  XOR U1347 ( .A(n1291), .B(n1292), .Z(n1244) );
  AND U1348 ( .A(n1293), .B(n1294), .Z(n1292) );
  XNOR U1349 ( .A(n1295), .B(n1296), .Z(n1293) );
  XNOR U1350 ( .A(n1297), .B(n1298), .Z(n1290) );
  AND U1351 ( .A(n1299), .B(n1300), .Z(n1298) );
  XNOR U1352 ( .A(n1297), .B(n1301), .Z(n1299) );
  XOR U1353 ( .A(n1302), .B(n1303), .Z(n1248) );
  AND U1354 ( .A(n1304), .B(n1305), .Z(n1303) );
  XOR U1355 ( .A(n1302), .B(n1306), .Z(n1304) );
  XNOR U1356 ( .A(n1258), .B(n1249), .Z(n1289) );
  XOR U1357 ( .A(n1307), .B(n1308), .Z(n1249) );
  NOR U1358 ( .A(n1309), .B(n1310), .Z(n1308) );
  XNOR U1359 ( .A(n1307), .B(n1311), .Z(n1309) );
  XOR U1360 ( .A(n1312), .B(n1264), .Z(n1258) );
  XNOR U1361 ( .A(n1313), .B(n1314), .Z(n1264) );
  AND U1362 ( .A(n1315), .B(n1316), .Z(n1314) );
  XOR U1363 ( .A(n1313), .B(n1317), .Z(n1315) );
  XNOR U1364 ( .A(n1263), .B(n1255), .Z(n1312) );
  XOR U1365 ( .A(n1318), .B(n1319), .Z(n1255) );
  AND U1366 ( .A(n1320), .B(n1321), .Z(n1319) );
  XOR U1367 ( .A(n1318), .B(n1322), .Z(n1320) );
  XNOR U1368 ( .A(n1323), .B(n1260), .Z(n1263) );
  XOR U1369 ( .A(n1324), .B(n1325), .Z(n1260) );
  AND U1370 ( .A(n1326), .B(n1327), .Z(n1325) );
  XNOR U1371 ( .A(n1328), .B(n1329), .Z(n1326) );
  XNOR U1372 ( .A(n1330), .B(n1331), .Z(n1323) );
  AND U1373 ( .A(n1332), .B(n1333), .Z(n1331) );
  XNOR U1374 ( .A(n1330), .B(n1334), .Z(n1332) );
  XOR U1375 ( .A(n1253), .B(n1265), .Z(n1288) );
  NOR U1376 ( .A(n1124), .B(n1335), .Z(n1265) );
  XNOR U1377 ( .A(n1271), .B(n1270), .Z(n1253) );
  XNOR U1378 ( .A(n1336), .B(n1276), .Z(n1270) );
  XOR U1379 ( .A(n1337), .B(n1338), .Z(n1276) );
  NOR U1380 ( .A(n1339), .B(n1340), .Z(n1338) );
  XNOR U1381 ( .A(n1337), .B(n1341), .Z(n1339) );
  XNOR U1382 ( .A(n1275), .B(n1267), .Z(n1336) );
  XOR U1383 ( .A(n1342), .B(n1343), .Z(n1267) );
  AND U1384 ( .A(n1344), .B(n1345), .Z(n1343) );
  XNOR U1385 ( .A(n1342), .B(n1346), .Z(n1344) );
  XNOR U1386 ( .A(n1347), .B(n1272), .Z(n1275) );
  XOR U1387 ( .A(n1348), .B(n1349), .Z(n1272) );
  AND U1388 ( .A(n1350), .B(n1351), .Z(n1349) );
  XOR U1389 ( .A(n1348), .B(n1352), .Z(n1350) );
  XNOR U1390 ( .A(n1353), .B(n1354), .Z(n1347) );
  AND U1391 ( .A(n1355), .B(n1356), .Z(n1354) );
  XNOR U1392 ( .A(n1353), .B(n1357), .Z(n1355) );
  XOR U1393 ( .A(n1281), .B(n1280), .Z(n1271) );
  XNOR U1394 ( .A(n1358), .B(n1277), .Z(n1280) );
  XOR U1395 ( .A(n1359), .B(n1360), .Z(n1277) );
  AND U1396 ( .A(n1361), .B(n1362), .Z(n1360) );
  XNOR U1397 ( .A(n1363), .B(n1364), .Z(n1361) );
  XNOR U1398 ( .A(n1365), .B(n1366), .Z(n1358) );
  AND U1399 ( .A(n1367), .B(n1368), .Z(n1366) );
  XNOR U1400 ( .A(n1365), .B(n1369), .Z(n1367) );
  XOR U1401 ( .A(n1370), .B(n1371), .Z(n1281) );
  AND U1402 ( .A(n1372), .B(n1373), .Z(n1371) );
  XOR U1403 ( .A(n1370), .B(n1374), .Z(n1372) );
  XNOR U1404 ( .A(n1189), .B(n1284), .Z(n1286) );
  XNOR U1405 ( .A(n1375), .B(n1376), .Z(n1189) );
  AND U1406 ( .A(n147), .B(n1195), .Z(n1376) );
  XOR U1407 ( .A(n1375), .B(n1193), .Z(n1195) );
  AND U1408 ( .A(n1196), .B(n1124), .Z(n1284) );
  XOR U1409 ( .A(n1377), .B(n1335), .Z(n1124) );
  XNOR U1410 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(
        p_input[128]), .Z(n1335) );
  XOR U1411 ( .A(n1311), .B(n1310), .Z(n1377) );
  XOR U1412 ( .A(n1378), .B(n1322), .Z(n1310) );
  XOR U1413 ( .A(n1296), .B(n1294), .Z(n1322) );
  XOR U1414 ( .A(n1379), .B(n1301), .Z(n1294) );
  XNOR U1415 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ), .B(
        p_input[152]), .Z(n1301) );
  XNOR U1416 ( .A(n1291), .B(n1300), .Z(n1379) );
  XNOR U1417 ( .A(n1380), .B(n1297), .Z(n1300) );
  XOR U1418 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ), .B(
        p_input[150]), .Z(n1297) );
  XNOR U1419 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ), .B(
        p_input[151]), .Z(n1380) );
  IV U1420 ( .A(n1295), .Z(n1291) );
  XNOR U1421 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ), .B(
        p_input[146]), .Z(n1295) );
  XOR U1422 ( .A(n1306), .B(n1305), .Z(n1296) );
  XNOR U1423 ( .A(n1381), .B(n1302), .Z(n1305) );
  XOR U1424 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ), .B(
        p_input[147]), .Z(n1302) );
  XNOR U1425 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ), .B(
        p_input[148]), .Z(n1381) );
  XOR U1426 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ), .B(
        p_input[149]), .Z(n1306) );
  XNOR U1427 ( .A(n1321), .B(n1307), .Z(n1378) );
  XOR U1428 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(
        p_input[129]), .Z(n1307) );
  XNOR U1429 ( .A(n1382), .B(n1329), .Z(n1321) );
  XOR U1430 ( .A(n1317), .B(n1316), .Z(n1329) );
  XNOR U1431 ( .A(n1383), .B(n1313), .Z(n1316) );
  XOR U1432 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ), .B(
        p_input[154]), .Z(n1313) );
  XNOR U1433 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ), .B(
        p_input[155]), .Z(n1383) );
  XOR U1434 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ), .B(
        p_input[156]), .Z(n1317) );
  XNOR U1435 ( .A(n1327), .B(n1318), .Z(n1382) );
  XOR U1436 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ), .B(
        p_input[145]), .Z(n1318) );
  XOR U1437 ( .A(n1384), .B(n1334), .Z(n1327) );
  XNOR U1438 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ), .B(
        p_input[159]), .Z(n1334) );
  XNOR U1439 ( .A(n1324), .B(n1333), .Z(n1384) );
  XNOR U1440 ( .A(n1385), .B(n1330), .Z(n1333) );
  XOR U1441 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ), .B(
        p_input[157]), .Z(n1330) );
  XNOR U1442 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ), .B(
        p_input[158]), .Z(n1385) );
  IV U1443 ( .A(n1328), .Z(n1324) );
  XNOR U1444 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ), .B(
        p_input[153]), .Z(n1328) );
  XNOR U1445 ( .A(n1346), .B(n1345), .Z(n1311) );
  XNOR U1446 ( .A(n1386), .B(n1352), .Z(n1345) );
  XNOR U1447 ( .A(n1341), .B(n1340), .Z(n1352) );
  XOR U1448 ( .A(n1387), .B(n1337), .Z(n1340) );
  XOR U1449 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(
        p_input[139]), .Z(n1337) );
  XOR U1450 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n1388), 
        .Z(n1387) );
  XOR U1451 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(
        p_input[141]), .Z(n1341) );
  XNOR U1452 ( .A(n1351), .B(n1342), .Z(n1386) );
  XOR U1453 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(
        p_input[130]), .Z(n1342) );
  XOR U1454 ( .A(n1389), .B(n1357), .Z(n1351) );
  XNOR U1455 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ), .B(
        p_input[144]), .Z(n1357) );
  XNOR U1456 ( .A(n1348), .B(n1356), .Z(n1389) );
  XNOR U1457 ( .A(n1390), .B(n1353), .Z(n1356) );
  XOR U1458 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(
        p_input[142]), .Z(n1353) );
  XNOR U1459 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(
        p_input[143]), .Z(n1390) );
  XOR U1460 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(
        p_input[138]), .Z(n1348) );
  XNOR U1461 ( .A(n1364), .B(n1362), .Z(n1346) );
  XOR U1462 ( .A(n1391), .B(n1369), .Z(n1362) );
  XNOR U1463 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(
        p_input[137]), .Z(n1369) );
  XNOR U1464 ( .A(n1359), .B(n1368), .Z(n1391) );
  XNOR U1465 ( .A(n1392), .B(n1365), .Z(n1368) );
  XOR U1466 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(
        p_input[135]), .Z(n1365) );
  XNOR U1467 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(
        p_input[136]), .Z(n1392) );
  IV U1468 ( .A(n1363), .Z(n1359) );
  XNOR U1469 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(
        p_input[131]), .Z(n1363) );
  XOR U1470 ( .A(n1374), .B(n1373), .Z(n1364) );
  XNOR U1471 ( .A(n1393), .B(n1370), .Z(n1373) );
  XOR U1472 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(
        p_input[132]), .Z(n1370) );
  XNOR U1473 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(
        p_input[133]), .Z(n1393) );
  XOR U1474 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(
        p_input[134]), .Z(n1374) );
  XNOR U1475 ( .A(n1394), .B(n1395), .Z(n1196) );
  AND U1476 ( .A(n147), .B(n1396), .Z(n1395) );
  XNOR U1477 ( .A(n1397), .B(n1398), .Z(n147) );
  NOR U1478 ( .A(n1399), .B(n1400), .Z(n1398) );
  XOR U1479 ( .A(n1158), .B(n1397), .Z(n1400) );
  NOR U1480 ( .A(n1397), .B(n1157), .Z(n1399) );
  XOR U1481 ( .A(n1401), .B(n1402), .Z(n1397) );
  AND U1482 ( .A(n1403), .B(n1404), .Z(n1402) );
  XNOR U1483 ( .A(n1212), .B(n1401), .Z(n1404) );
  XOR U1484 ( .A(n1401), .B(n1166), .Z(n1403) );
  XOR U1485 ( .A(n1405), .B(n1406), .Z(n1401) );
  AND U1486 ( .A(n1407), .B(n1408), .Z(n1406) );
  XNOR U1487 ( .A(n1236), .B(n1405), .Z(n1408) );
  XOR U1488 ( .A(n1405), .B(n1175), .Z(n1407) );
  XOR U1489 ( .A(n1409), .B(n1410), .Z(n1405) );
  AND U1490 ( .A(n1411), .B(n1412), .Z(n1410) );
  XOR U1491 ( .A(n1409), .B(n1182), .Z(n1411) );
  XOR U1492 ( .A(n1413), .B(n1414), .Z(n1150) );
  AND U1493 ( .A(n150), .B(n1396), .Z(n1414) );
  XOR U1494 ( .A(n1415), .B(n1413), .Z(n1396) );
  XNOR U1495 ( .A(n1416), .B(n1417), .Z(n150) );
  NOR U1496 ( .A(n1418), .B(n1419), .Z(n1417) );
  XNOR U1497 ( .A(n1158), .B(n1420), .Z(n1419) );
  IV U1498 ( .A(n1416), .Z(n1420) );
  AND U1499 ( .A(n1166), .B(n1421), .Z(n1158) );
  NOR U1500 ( .A(n1416), .B(n1157), .Z(n1418) );
  AND U1501 ( .A(n1212), .B(n1422), .Z(n1157) );
  XOR U1502 ( .A(n1423), .B(n1424), .Z(n1416) );
  AND U1503 ( .A(n1425), .B(n1426), .Z(n1424) );
  XNOR U1504 ( .A(n1423), .B(n1212), .Z(n1426) );
  XNOR U1505 ( .A(n1427), .B(n1428), .Z(n1212) );
  XOR U1506 ( .A(n1429), .B(n1422), .Z(n1428) );
  AND U1507 ( .A(n1236), .B(n1430), .Z(n1422) );
  AND U1508 ( .A(n1431), .B(n1432), .Z(n1429) );
  XOR U1509 ( .A(n1433), .B(n1427), .Z(n1431) );
  XNOR U1510 ( .A(n1434), .B(n1423), .Z(n1425) );
  IV U1511 ( .A(n1166), .Z(n1434) );
  XNOR U1512 ( .A(n1435), .B(n1436), .Z(n1166) );
  XOR U1513 ( .A(n1437), .B(n1421), .Z(n1436) );
  AND U1514 ( .A(n1175), .B(n1438), .Z(n1421) );
  AND U1515 ( .A(n1439), .B(n1440), .Z(n1437) );
  XNOR U1516 ( .A(n1435), .B(n1441), .Z(n1439) );
  XOR U1517 ( .A(n1442), .B(n1443), .Z(n1423) );
  AND U1518 ( .A(n1444), .B(n1445), .Z(n1443) );
  XNOR U1519 ( .A(n1442), .B(n1236), .Z(n1445) );
  XOR U1520 ( .A(n1446), .B(n1432), .Z(n1236) );
  XNOR U1521 ( .A(n1447), .B(n1427), .Z(n1432) );
  XOR U1522 ( .A(n1448), .B(n1449), .Z(n1427) );
  AND U1523 ( .A(n1450), .B(n1451), .Z(n1449) );
  XOR U1524 ( .A(n1452), .B(n1448), .Z(n1450) );
  XNOR U1525 ( .A(n1453), .B(n1454), .Z(n1447) );
  AND U1526 ( .A(n1455), .B(n1456), .Z(n1454) );
  XOR U1527 ( .A(n1453), .B(n1457), .Z(n1455) );
  XNOR U1528 ( .A(n1433), .B(n1430), .Z(n1446) );
  AND U1529 ( .A(n1282), .B(n1458), .Z(n1430) );
  XOR U1530 ( .A(n1459), .B(n1460), .Z(n1433) );
  AND U1531 ( .A(n1461), .B(n1462), .Z(n1460) );
  XOR U1532 ( .A(n1459), .B(n1463), .Z(n1461) );
  XOR U1533 ( .A(n1175), .B(n1442), .Z(n1444) );
  XNOR U1534 ( .A(n1464), .B(n1441), .Z(n1175) );
  XNOR U1535 ( .A(n1465), .B(n1466), .Z(n1441) );
  AND U1536 ( .A(n1467), .B(n1468), .Z(n1466) );
  XOR U1537 ( .A(n1465), .B(n1469), .Z(n1467) );
  XNOR U1538 ( .A(n1440), .B(n1438), .Z(n1464) );
  AND U1539 ( .A(n1182), .B(n1470), .Z(n1438) );
  XNOR U1540 ( .A(n1471), .B(n1435), .Z(n1440) );
  XOR U1541 ( .A(n1472), .B(n1473), .Z(n1435) );
  AND U1542 ( .A(n1474), .B(n1475), .Z(n1473) );
  XOR U1543 ( .A(n1472), .B(n1476), .Z(n1474) );
  XNOR U1544 ( .A(n1477), .B(n1478), .Z(n1471) );
  AND U1545 ( .A(n1479), .B(n1480), .Z(n1478) );
  XNOR U1546 ( .A(n1477), .B(n1481), .Z(n1479) );
  XOR U1547 ( .A(n1409), .B(n1482), .Z(n1442) );
  AND U1548 ( .A(n1483), .B(n1412), .Z(n1482) );
  XNOR U1549 ( .A(n1282), .B(n1409), .Z(n1412) );
  XOR U1550 ( .A(n1484), .B(n1451), .Z(n1282) );
  XNOR U1551 ( .A(n1485), .B(n1457), .Z(n1451) );
  XOR U1552 ( .A(n1486), .B(n1487), .Z(n1457) );
  AND U1553 ( .A(n1488), .B(n1489), .Z(n1487) );
  XOR U1554 ( .A(n1486), .B(n1490), .Z(n1488) );
  XNOR U1555 ( .A(n1456), .B(n1448), .Z(n1485) );
  XOR U1556 ( .A(n1491), .B(n1492), .Z(n1448) );
  AND U1557 ( .A(n1493), .B(n1494), .Z(n1492) );
  XNOR U1558 ( .A(n1495), .B(n1491), .Z(n1493) );
  XNOR U1559 ( .A(n1496), .B(n1453), .Z(n1456) );
  XOR U1560 ( .A(n1497), .B(n1498), .Z(n1453) );
  AND U1561 ( .A(n1499), .B(n1500), .Z(n1498) );
  XOR U1562 ( .A(n1497), .B(n1501), .Z(n1499) );
  XNOR U1563 ( .A(n1502), .B(n1503), .Z(n1496) );
  AND U1564 ( .A(n1504), .B(n1505), .Z(n1503) );
  XNOR U1565 ( .A(n1502), .B(n1506), .Z(n1504) );
  XNOR U1566 ( .A(n1452), .B(n1458), .Z(n1484) );
  AND U1567 ( .A(n1375), .B(n1507), .Z(n1458) );
  XOR U1568 ( .A(n1463), .B(n1462), .Z(n1452) );
  XNOR U1569 ( .A(n1508), .B(n1459), .Z(n1462) );
  XOR U1570 ( .A(n1509), .B(n1510), .Z(n1459) );
  AND U1571 ( .A(n1511), .B(n1512), .Z(n1510) );
  XOR U1572 ( .A(n1509), .B(n1513), .Z(n1511) );
  XNOR U1573 ( .A(n1514), .B(n1515), .Z(n1508) );
  AND U1574 ( .A(n1516), .B(n1517), .Z(n1515) );
  XOR U1575 ( .A(n1514), .B(n1518), .Z(n1516) );
  XOR U1576 ( .A(n1519), .B(n1520), .Z(n1463) );
  AND U1577 ( .A(n1521), .B(n1522), .Z(n1520) );
  XOR U1578 ( .A(n1519), .B(n1523), .Z(n1521) );
  XNOR U1579 ( .A(n1524), .B(n1409), .Z(n1483) );
  IV U1580 ( .A(n1182), .Z(n1524) );
  XOR U1581 ( .A(n1525), .B(n1476), .Z(n1182) );
  XOR U1582 ( .A(n1469), .B(n1468), .Z(n1476) );
  XNOR U1583 ( .A(n1526), .B(n1465), .Z(n1468) );
  XOR U1584 ( .A(n1527), .B(n1528), .Z(n1465) );
  AND U1585 ( .A(n1529), .B(n1530), .Z(n1528) );
  XOR U1586 ( .A(n1527), .B(n1531), .Z(n1529) );
  XNOR U1587 ( .A(n1532), .B(n1533), .Z(n1526) );
  AND U1588 ( .A(n1534), .B(n1535), .Z(n1533) );
  XOR U1589 ( .A(n1532), .B(n1536), .Z(n1534) );
  XOR U1590 ( .A(n1537), .B(n1538), .Z(n1469) );
  AND U1591 ( .A(n1539), .B(n1540), .Z(n1538) );
  XOR U1592 ( .A(n1537), .B(n1541), .Z(n1539) );
  XNOR U1593 ( .A(n1475), .B(n1470), .Z(n1525) );
  AND U1594 ( .A(n1193), .B(n1542), .Z(n1470) );
  XOR U1595 ( .A(n1543), .B(n1481), .Z(n1475) );
  XNOR U1596 ( .A(n1544), .B(n1545), .Z(n1481) );
  AND U1597 ( .A(n1546), .B(n1547), .Z(n1545) );
  XOR U1598 ( .A(n1544), .B(n1548), .Z(n1546) );
  XNOR U1599 ( .A(n1480), .B(n1472), .Z(n1543) );
  XOR U1600 ( .A(n1549), .B(n1550), .Z(n1472) );
  AND U1601 ( .A(n1551), .B(n1552), .Z(n1550) );
  XOR U1602 ( .A(n1549), .B(n1553), .Z(n1551) );
  XNOR U1603 ( .A(n1554), .B(n1477), .Z(n1480) );
  XOR U1604 ( .A(n1555), .B(n1556), .Z(n1477) );
  AND U1605 ( .A(n1557), .B(n1558), .Z(n1556) );
  XOR U1606 ( .A(n1555), .B(n1559), .Z(n1557) );
  XNOR U1607 ( .A(n1560), .B(n1561), .Z(n1554) );
  AND U1608 ( .A(n1562), .B(n1563), .Z(n1561) );
  XNOR U1609 ( .A(n1560), .B(n1564), .Z(n1562) );
  XOR U1610 ( .A(n1565), .B(n1566), .Z(n1409) );
  AND U1611 ( .A(n1567), .B(n1568), .Z(n1566) );
  XNOR U1612 ( .A(n1565), .B(n1375), .Z(n1568) );
  XOR U1613 ( .A(n1569), .B(n1494), .Z(n1375) );
  XNOR U1614 ( .A(n1570), .B(n1501), .Z(n1494) );
  XOR U1615 ( .A(n1490), .B(n1489), .Z(n1501) );
  XNOR U1616 ( .A(n1571), .B(n1486), .Z(n1489) );
  XOR U1617 ( .A(n1572), .B(n1573), .Z(n1486) );
  AND U1618 ( .A(n1574), .B(n1575), .Z(n1573) );
  XOR U1619 ( .A(n1572), .B(n1576), .Z(n1574) );
  XNOR U1620 ( .A(n1577), .B(n1578), .Z(n1571) );
  NOR U1621 ( .A(n1579), .B(n1580), .Z(n1578) );
  XNOR U1622 ( .A(n1577), .B(n1581), .Z(n1579) );
  XOR U1623 ( .A(n1582), .B(n1583), .Z(n1490) );
  NOR U1624 ( .A(n1584), .B(n1585), .Z(n1583) );
  XNOR U1625 ( .A(n1582), .B(n1586), .Z(n1584) );
  XNOR U1626 ( .A(n1500), .B(n1491), .Z(n1570) );
  XOR U1627 ( .A(n1587), .B(n1588), .Z(n1491) );
  NOR U1628 ( .A(n1589), .B(n1590), .Z(n1588) );
  XNOR U1629 ( .A(n1587), .B(n1591), .Z(n1589) );
  XOR U1630 ( .A(n1592), .B(n1506), .Z(n1500) );
  XNOR U1631 ( .A(n1593), .B(n1594), .Z(n1506) );
  NOR U1632 ( .A(n1595), .B(n1596), .Z(n1594) );
  XNOR U1633 ( .A(n1593), .B(n1597), .Z(n1595) );
  XNOR U1634 ( .A(n1505), .B(n1497), .Z(n1592) );
  XOR U1635 ( .A(n1598), .B(n1599), .Z(n1497) );
  AND U1636 ( .A(n1600), .B(n1601), .Z(n1599) );
  XOR U1637 ( .A(n1598), .B(n1602), .Z(n1600) );
  XNOR U1638 ( .A(n1603), .B(n1502), .Z(n1505) );
  XOR U1639 ( .A(n1604), .B(n1605), .Z(n1502) );
  AND U1640 ( .A(n1606), .B(n1607), .Z(n1605) );
  XOR U1641 ( .A(n1604), .B(n1608), .Z(n1606) );
  XNOR U1642 ( .A(n1609), .B(n1610), .Z(n1603) );
  NOR U1643 ( .A(n1611), .B(n1612), .Z(n1610) );
  XOR U1644 ( .A(n1609), .B(n1613), .Z(n1611) );
  XOR U1645 ( .A(n1495), .B(n1507), .Z(n1569) );
  AND U1646 ( .A(n1415), .B(n1614), .Z(n1507) );
  IV U1647 ( .A(n1394), .Z(n1415) );
  XNOR U1648 ( .A(n1513), .B(n1512), .Z(n1495) );
  XNOR U1649 ( .A(n1615), .B(n1518), .Z(n1512) );
  XOR U1650 ( .A(n1616), .B(n1617), .Z(n1518) );
  NOR U1651 ( .A(n1618), .B(n1619), .Z(n1617) );
  XNOR U1652 ( .A(n1616), .B(n1620), .Z(n1618) );
  XNOR U1653 ( .A(n1517), .B(n1509), .Z(n1615) );
  XOR U1654 ( .A(n1621), .B(n1622), .Z(n1509) );
  AND U1655 ( .A(n1623), .B(n1624), .Z(n1622) );
  XNOR U1656 ( .A(n1621), .B(n1625), .Z(n1623) );
  XNOR U1657 ( .A(n1626), .B(n1514), .Z(n1517) );
  XOR U1658 ( .A(n1627), .B(n1628), .Z(n1514) );
  AND U1659 ( .A(n1629), .B(n1630), .Z(n1628) );
  XOR U1660 ( .A(n1627), .B(n1631), .Z(n1629) );
  XNOR U1661 ( .A(n1632), .B(n1633), .Z(n1626) );
  NOR U1662 ( .A(n1634), .B(n1635), .Z(n1633) );
  XOR U1663 ( .A(n1632), .B(n1636), .Z(n1634) );
  XOR U1664 ( .A(n1523), .B(n1522), .Z(n1513) );
  XNOR U1665 ( .A(n1637), .B(n1519), .Z(n1522) );
  XOR U1666 ( .A(n1638), .B(n1639), .Z(n1519) );
  AND U1667 ( .A(n1640), .B(n1641), .Z(n1639) );
  XOR U1668 ( .A(n1638), .B(n1642), .Z(n1640) );
  XNOR U1669 ( .A(n1643), .B(n1644), .Z(n1637) );
  NOR U1670 ( .A(n1645), .B(n1646), .Z(n1644) );
  XNOR U1671 ( .A(n1643), .B(n1647), .Z(n1645) );
  XOR U1672 ( .A(n1648), .B(n1649), .Z(n1523) );
  NOR U1673 ( .A(n1650), .B(n1651), .Z(n1649) );
  XNOR U1674 ( .A(n1648), .B(n1652), .Z(n1650) );
  XNOR U1675 ( .A(n1653), .B(n1565), .Z(n1567) );
  IV U1676 ( .A(n1193), .Z(n1653) );
  XOR U1677 ( .A(n1654), .B(n1553), .Z(n1193) );
  XOR U1678 ( .A(n1531), .B(n1530), .Z(n1553) );
  XNOR U1679 ( .A(n1655), .B(n1536), .Z(n1530) );
  XOR U1680 ( .A(n1656), .B(n1657), .Z(n1536) );
  NOR U1681 ( .A(n1658), .B(n1659), .Z(n1657) );
  XNOR U1682 ( .A(n1656), .B(n1660), .Z(n1658) );
  XNOR U1683 ( .A(n1535), .B(n1527), .Z(n1655) );
  XOR U1684 ( .A(n1661), .B(n1662), .Z(n1527) );
  AND U1685 ( .A(n1663), .B(n1664), .Z(n1662) );
  XNOR U1686 ( .A(n1661), .B(n1665), .Z(n1663) );
  XNOR U1687 ( .A(n1666), .B(n1532), .Z(n1535) );
  XOR U1688 ( .A(n1667), .B(n1668), .Z(n1532) );
  AND U1689 ( .A(n1669), .B(n1670), .Z(n1668) );
  XOR U1690 ( .A(n1667), .B(n1671), .Z(n1669) );
  XNOR U1691 ( .A(n1672), .B(n1673), .Z(n1666) );
  NOR U1692 ( .A(n1674), .B(n1675), .Z(n1673) );
  XOR U1693 ( .A(n1672), .B(n1676), .Z(n1674) );
  XOR U1694 ( .A(n1541), .B(n1540), .Z(n1531) );
  XNOR U1695 ( .A(n1677), .B(n1537), .Z(n1540) );
  XOR U1696 ( .A(n1678), .B(n1679), .Z(n1537) );
  AND U1697 ( .A(n1680), .B(n1681), .Z(n1679) );
  XOR U1698 ( .A(n1678), .B(n1682), .Z(n1680) );
  XNOR U1699 ( .A(n1683), .B(n1684), .Z(n1677) );
  NOR U1700 ( .A(n1685), .B(n1686), .Z(n1684) );
  XNOR U1701 ( .A(n1683), .B(n1687), .Z(n1685) );
  XOR U1702 ( .A(n1688), .B(n1689), .Z(n1541) );
  NOR U1703 ( .A(n1690), .B(n1691), .Z(n1689) );
  XNOR U1704 ( .A(n1688), .B(n1692), .Z(n1690) );
  XNOR U1705 ( .A(n1552), .B(n1542), .Z(n1654) );
  AND U1706 ( .A(n1413), .B(n1693), .Z(n1542) );
  XNOR U1707 ( .A(n1694), .B(n1559), .Z(n1552) );
  XOR U1708 ( .A(n1548), .B(n1547), .Z(n1559) );
  XNOR U1709 ( .A(n1695), .B(n1544), .Z(n1547) );
  XOR U1710 ( .A(n1696), .B(n1697), .Z(n1544) );
  AND U1711 ( .A(n1698), .B(n1699), .Z(n1697) );
  XOR U1712 ( .A(n1696), .B(n1700), .Z(n1698) );
  XNOR U1713 ( .A(n1701), .B(n1702), .Z(n1695) );
  NOR U1714 ( .A(n1703), .B(n1704), .Z(n1702) );
  XNOR U1715 ( .A(n1701), .B(n1705), .Z(n1703) );
  XOR U1716 ( .A(n1706), .B(n1707), .Z(n1548) );
  NOR U1717 ( .A(n1708), .B(n1709), .Z(n1707) );
  XNOR U1718 ( .A(n1706), .B(n1710), .Z(n1708) );
  XNOR U1719 ( .A(n1558), .B(n1549), .Z(n1694) );
  XOR U1720 ( .A(n1711), .B(n1712), .Z(n1549) );
  NOR U1721 ( .A(n1713), .B(n1714), .Z(n1712) );
  XNOR U1722 ( .A(n1711), .B(n1715), .Z(n1713) );
  XOR U1723 ( .A(n1716), .B(n1564), .Z(n1558) );
  XNOR U1724 ( .A(n1717), .B(n1718), .Z(n1564) );
  NOR U1725 ( .A(n1719), .B(n1720), .Z(n1718) );
  XNOR U1726 ( .A(n1717), .B(n1721), .Z(n1719) );
  XNOR U1727 ( .A(n1563), .B(n1555), .Z(n1716) );
  XOR U1728 ( .A(n1722), .B(n1723), .Z(n1555) );
  AND U1729 ( .A(n1724), .B(n1725), .Z(n1723) );
  XOR U1730 ( .A(n1722), .B(n1726), .Z(n1724) );
  XNOR U1731 ( .A(n1727), .B(n1560), .Z(n1563) );
  XOR U1732 ( .A(n1728), .B(n1729), .Z(n1560) );
  AND U1733 ( .A(n1730), .B(n1731), .Z(n1729) );
  XOR U1734 ( .A(n1728), .B(n1732), .Z(n1730) );
  XNOR U1735 ( .A(n1733), .B(n1734), .Z(n1727) );
  NOR U1736 ( .A(n1735), .B(n1736), .Z(n1734) );
  XOR U1737 ( .A(n1733), .B(n1737), .Z(n1735) );
  AND U1738 ( .A(n1413), .B(n1394), .Z(n1565) );
  XNOR U1739 ( .A(n1738), .B(n1614), .Z(n1394) );
  XOR U1740 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(
        p_input[128]), .Z(n1614) );
  XOR U1741 ( .A(n1591), .B(n1590), .Z(n1738) );
  XOR U1742 ( .A(n1739), .B(n1602), .Z(n1590) );
  XOR U1743 ( .A(n1576), .B(n1575), .Z(n1602) );
  XNOR U1744 ( .A(n1740), .B(n1581), .Z(n1575) );
  XOR U1745 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .B(
        p_input[152]), .Z(n1581) );
  XOR U1746 ( .A(n1572), .B(n1580), .Z(n1740) );
  XOR U1747 ( .A(n1741), .B(n1577), .Z(n1580) );
  XOR U1748 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .B(
        p_input[150]), .Z(n1577) );
  XOR U1749 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .B(n1742), 
        .Z(n1741) );
  XOR U1750 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .B(
        p_input[146]), .Z(n1572) );
  XNOR U1751 ( .A(n1586), .B(n1585), .Z(n1576) );
  XOR U1752 ( .A(n1743), .B(n1582), .Z(n1585) );
  XOR U1753 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .B(
        p_input[147]), .Z(n1582) );
  XOR U1754 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .B(n1744), 
        .Z(n1743) );
  XOR U1755 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .B(
        p_input[149]), .Z(n1586) );
  XNOR U1756 ( .A(n1601), .B(n1587), .Z(n1739) );
  XOR U1757 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(
        p_input[129]), .Z(n1587) );
  XNOR U1758 ( .A(n1745), .B(n1608), .Z(n1601) );
  XNOR U1759 ( .A(n1597), .B(n1596), .Z(n1608) );
  XOR U1760 ( .A(n1746), .B(n1593), .Z(n1596) );
  XOR U1761 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .B(
        p_input[154]), .Z(n1593) );
  XOR U1762 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .B(n1747), 
        .Z(n1746) );
  XOR U1763 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .B(
        p_input[156]), .Z(n1597) );
  XNOR U1764 ( .A(n1607), .B(n1598), .Z(n1745) );
  XOR U1765 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .B(
        p_input[145]), .Z(n1598) );
  XOR U1766 ( .A(n1748), .B(n1613), .Z(n1607) );
  XNOR U1767 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .B(
        p_input[159]), .Z(n1613) );
  XOR U1768 ( .A(n1604), .B(n1612), .Z(n1748) );
  XOR U1769 ( .A(n1749), .B(n1609), .Z(n1612) );
  XOR U1770 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .B(
        p_input[157]), .Z(n1609) );
  XOR U1771 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .B(n1750), 
        .Z(n1749) );
  XOR U1772 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .B(
        p_input[153]), .Z(n1604) );
  XNOR U1773 ( .A(n1625), .B(n1624), .Z(n1591) );
  XNOR U1774 ( .A(n1751), .B(n1631), .Z(n1624) );
  XNOR U1775 ( .A(n1620), .B(n1619), .Z(n1631) );
  XOR U1776 ( .A(n1752), .B(n1616), .Z(n1619) );
  XOR U1777 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(
        p_input[139]), .Z(n1616) );
  XOR U1778 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n1388), 
        .Z(n1752) );
  XOR U1779 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(
        p_input[141]), .Z(n1620) );
  XNOR U1780 ( .A(n1630), .B(n1621), .Z(n1751) );
  XOR U1781 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(
        p_input[130]), .Z(n1621) );
  XOR U1782 ( .A(n1753), .B(n1636), .Z(n1630) );
  XNOR U1783 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .B(
        p_input[144]), .Z(n1636) );
  XOR U1784 ( .A(n1627), .B(n1635), .Z(n1753) );
  XOR U1785 ( .A(n1754), .B(n1632), .Z(n1635) );
  XOR U1786 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(
        p_input[142]), .Z(n1632) );
  XOR U1787 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n1755), 
        .Z(n1754) );
  XOR U1788 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(
        p_input[138]), .Z(n1627) );
  XNOR U1789 ( .A(n1642), .B(n1641), .Z(n1625) );
  XNOR U1790 ( .A(n1756), .B(n1647), .Z(n1641) );
  XOR U1791 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .B(
        p_input[137]), .Z(n1647) );
  XOR U1792 ( .A(n1638), .B(n1646), .Z(n1756) );
  XOR U1793 ( .A(n1757), .B(n1643), .Z(n1646) );
  XOR U1794 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(
        p_input[135]), .Z(n1643) );
  XNOR U1795 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(
        p_input[136]), .Z(n1757) );
  XOR U1796 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(
        p_input[131]), .Z(n1638) );
  XNOR U1797 ( .A(n1652), .B(n1651), .Z(n1642) );
  XOR U1798 ( .A(n1758), .B(n1648), .Z(n1651) );
  XOR U1799 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(
        p_input[132]), .Z(n1648) );
  XOR U1800 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n1759), 
        .Z(n1758) );
  XOR U1801 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(
        p_input[134]), .Z(n1652) );
  XOR U1802 ( .A(n1760), .B(n1715), .Z(n1413) );
  XNOR U1803 ( .A(n1665), .B(n1664), .Z(n1715) );
  XNOR U1804 ( .A(n1761), .B(n1671), .Z(n1664) );
  XNOR U1805 ( .A(n1660), .B(n1659), .Z(n1671) );
  XOR U1806 ( .A(n1762), .B(n1656), .Z(n1659) );
  XOR U1807 ( .A(\knn_comb_/min_val_out[0][11] ), .B(p_input[139]), .Z(n1656)
         );
  XOR U1808 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n1388), .Z(n1762) );
  IV U1809 ( .A(p_input[140]), .Z(n1388) );
  XOR U1810 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[141]), .Z(n1660)
         );
  XNOR U1811 ( .A(n1670), .B(n1661), .Z(n1761) );
  XOR U1812 ( .A(\knn_comb_/min_val_out[0][2] ), .B(p_input[130]), .Z(n1661)
         );
  XOR U1813 ( .A(n1763), .B(n1676), .Z(n1670) );
  XNOR U1814 ( .A(\knn_comb_/min_val_out[0][16] ), .B(p_input[144]), .Z(n1676)
         );
  XOR U1815 ( .A(n1667), .B(n1675), .Z(n1763) );
  XOR U1816 ( .A(n1764), .B(n1672), .Z(n1675) );
  XOR U1817 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[142]), .Z(n1672)
         );
  XOR U1818 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n1755), .Z(n1764) );
  IV U1819 ( .A(p_input[143]), .Z(n1755) );
  XOR U1820 ( .A(\knn_comb_/min_val_out[0][10] ), .B(p_input[138]), .Z(n1667)
         );
  XNOR U1821 ( .A(n1682), .B(n1681), .Z(n1665) );
  XNOR U1822 ( .A(n1765), .B(n1687), .Z(n1681) );
  XOR U1823 ( .A(\knn_comb_/min_val_out[0][9] ), .B(p_input[137]), .Z(n1687)
         );
  XOR U1824 ( .A(n1678), .B(n1686), .Z(n1765) );
  XOR U1825 ( .A(n1766), .B(n1683), .Z(n1686) );
  XOR U1826 ( .A(\knn_comb_/min_val_out[0][7] ), .B(p_input[135]), .Z(n1683)
         );
  XNOR U1827 ( .A(\knn_comb_/min_val_out[0][8] ), .B(p_input[136]), .Z(n1766)
         );
  XOR U1828 ( .A(\knn_comb_/min_val_out[0][3] ), .B(p_input[131]), .Z(n1678)
         );
  XNOR U1829 ( .A(n1692), .B(n1691), .Z(n1682) );
  XOR U1830 ( .A(n1767), .B(n1688), .Z(n1691) );
  XOR U1831 ( .A(\knn_comb_/min_val_out[0][4] ), .B(p_input[132]), .Z(n1688)
         );
  XOR U1832 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n1759), .Z(n1767) );
  IV U1833 ( .A(p_input[133]), .Z(n1759) );
  XOR U1834 ( .A(\knn_comb_/min_val_out[0][6] ), .B(p_input[134]), .Z(n1692)
         );
  XOR U1835 ( .A(n1714), .B(n1693), .Z(n1760) );
  XOR U1836 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[128]), .Z(n1693)
         );
  XOR U1837 ( .A(n1768), .B(n1726), .Z(n1714) );
  XOR U1838 ( .A(n1700), .B(n1699), .Z(n1726) );
  XNOR U1839 ( .A(n1769), .B(n1705), .Z(n1699) );
  XOR U1840 ( .A(\knn_comb_/min_val_out[0][24] ), .B(p_input[152]), .Z(n1705)
         );
  XOR U1841 ( .A(n1696), .B(n1704), .Z(n1769) );
  XOR U1842 ( .A(n1770), .B(n1701), .Z(n1704) );
  XOR U1843 ( .A(\knn_comb_/min_val_out[0][22] ), .B(p_input[150]), .Z(n1701)
         );
  XOR U1844 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n1742), .Z(n1770) );
  IV U1845 ( .A(p_input[151]), .Z(n1742) );
  XOR U1846 ( .A(\knn_comb_/min_val_out[0][18] ), .B(p_input[146]), .Z(n1696)
         );
  XNOR U1847 ( .A(n1710), .B(n1709), .Z(n1700) );
  XOR U1848 ( .A(n1771), .B(n1706), .Z(n1709) );
  XOR U1849 ( .A(\knn_comb_/min_val_out[0][19] ), .B(p_input[147]), .Z(n1706)
         );
  XOR U1850 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n1744), .Z(n1771) );
  IV U1851 ( .A(p_input[148]), .Z(n1744) );
  XOR U1852 ( .A(\knn_comb_/min_val_out[0][21] ), .B(p_input[149]), .Z(n1710)
         );
  XNOR U1853 ( .A(n1725), .B(n1711), .Z(n1768) );
  XOR U1854 ( .A(\knn_comb_/min_val_out[0][1] ), .B(p_input[129]), .Z(n1711)
         );
  XNOR U1855 ( .A(n1772), .B(n1732), .Z(n1725) );
  XNOR U1856 ( .A(n1721), .B(n1720), .Z(n1732) );
  XOR U1857 ( .A(n1773), .B(n1717), .Z(n1720) );
  XOR U1858 ( .A(\knn_comb_/min_val_out[0][26] ), .B(p_input[154]), .Z(n1717)
         );
  XOR U1859 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n1747), .Z(n1773) );
  IV U1860 ( .A(p_input[155]), .Z(n1747) );
  XOR U1861 ( .A(\knn_comb_/min_val_out[0][28] ), .B(p_input[156]), .Z(n1721)
         );
  XNOR U1862 ( .A(n1731), .B(n1722), .Z(n1772) );
  XOR U1863 ( .A(\knn_comb_/min_val_out[0][17] ), .B(p_input[145]), .Z(n1722)
         );
  XOR U1864 ( .A(n1774), .B(n1737), .Z(n1731) );
  XNOR U1865 ( .A(\knn_comb_/min_val_out[0][31] ), .B(p_input[159]), .Z(n1737)
         );
  XOR U1866 ( .A(n1728), .B(n1736), .Z(n1774) );
  XOR U1867 ( .A(n1775), .B(n1733), .Z(n1736) );
  XOR U1868 ( .A(\knn_comb_/min_val_out[0][29] ), .B(p_input[157]), .Z(n1733)
         );
  XOR U1869 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n1750), .Z(n1775) );
  IV U1870 ( .A(p_input[158]), .Z(n1750) );
  XOR U1871 ( .A(\knn_comb_/min_val_out[0][25] ), .B(p_input[153]), .Z(n1728)
         );
endmodule

