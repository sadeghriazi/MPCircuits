
module auction_BMR_N2_W32 ( p_input, o );
  input [127:0] p_input;
  output [33:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662;

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(o[1]), .B(n3), .Z(n1) );
  XOR U3 ( .A(n2), .B(n4), .Z(n3) );
  XNOR U4 ( .A(n5), .B(n6), .Z(o[8]) );
  AND U5 ( .A(o[1]), .B(n7), .Z(n5) );
  XOR U6 ( .A(n8), .B(n6), .Z(n7) );
  XNOR U7 ( .A(n9), .B(n10), .Z(o[7]) );
  AND U8 ( .A(o[1]), .B(n11), .Z(n9) );
  XOR U9 ( .A(n12), .B(n10), .Z(n11) );
  XNOR U10 ( .A(n13), .B(n14), .Z(o[6]) );
  AND U11 ( .A(o[1]), .B(n15), .Z(n13) );
  XOR U12 ( .A(n16), .B(n14), .Z(n15) );
  XNOR U13 ( .A(n17), .B(n18), .Z(o[5]) );
  AND U14 ( .A(o[1]), .B(n19), .Z(n17) );
  XOR U15 ( .A(n20), .B(n18), .Z(n19) );
  XNOR U16 ( .A(n21), .B(n22), .Z(o[4]) );
  AND U17 ( .A(o[1]), .B(n23), .Z(n21) );
  XOR U18 ( .A(n24), .B(n22), .Z(n23) );
  XOR U19 ( .A(n25), .B(n26), .Z(o[3]) );
  AND U20 ( .A(o[1]), .B(n27), .Z(n25) );
  XOR U21 ( .A(n28), .B(n29), .Z(n27) );
  XOR U22 ( .A(n30), .B(n31), .Z(o[33]) );
  AND U23 ( .A(n32), .B(o[1]), .Z(n30) );
  AND U24 ( .A(n31), .B(n33), .Z(n32) );
  XNOR U25 ( .A(n34), .B(n35), .Z(o[32]) );
  AND U26 ( .A(o[1]), .B(n36), .Z(n34) );
  XOR U27 ( .A(n37), .B(n35), .Z(n36) );
  XNOR U28 ( .A(n38), .B(n39), .Z(o[31]) );
  AND U29 ( .A(o[1]), .B(n40), .Z(n38) );
  XOR U30 ( .A(n41), .B(n39), .Z(n40) );
  XNOR U31 ( .A(n42), .B(n43), .Z(o[30]) );
  AND U32 ( .A(o[1]), .B(n44), .Z(n42) );
  XOR U33 ( .A(n45), .B(n43), .Z(n44) );
  XNOR U34 ( .A(n46), .B(n47), .Z(o[2]) );
  AND U35 ( .A(o[1]), .B(n48), .Z(n46) );
  XNOR U36 ( .A(n49), .B(n47), .Z(n48) );
  XNOR U37 ( .A(n50), .B(n51), .Z(o[29]) );
  AND U38 ( .A(o[1]), .B(n52), .Z(n50) );
  XOR U39 ( .A(n53), .B(n51), .Z(n52) );
  XNOR U40 ( .A(n54), .B(n55), .Z(o[28]) );
  AND U41 ( .A(o[1]), .B(n56), .Z(n54) );
  XOR U42 ( .A(n57), .B(n55), .Z(n56) );
  XNOR U43 ( .A(n58), .B(n59), .Z(o[27]) );
  AND U44 ( .A(o[1]), .B(n60), .Z(n58) );
  XOR U45 ( .A(n61), .B(n59), .Z(n60) );
  XNOR U46 ( .A(n62), .B(n63), .Z(o[26]) );
  AND U47 ( .A(o[1]), .B(n64), .Z(n62) );
  XOR U48 ( .A(n65), .B(n63), .Z(n64) );
  XNOR U49 ( .A(n66), .B(n67), .Z(o[25]) );
  AND U50 ( .A(o[1]), .B(n68), .Z(n66) );
  XOR U51 ( .A(n69), .B(n67), .Z(n68) );
  XNOR U52 ( .A(n70), .B(n71), .Z(o[24]) );
  AND U53 ( .A(o[1]), .B(n72), .Z(n70) );
  XOR U54 ( .A(n73), .B(n71), .Z(n72) );
  XNOR U55 ( .A(n74), .B(n75), .Z(o[23]) );
  AND U56 ( .A(o[1]), .B(n76), .Z(n74) );
  XOR U57 ( .A(n77), .B(n75), .Z(n76) );
  XNOR U58 ( .A(n78), .B(n79), .Z(o[22]) );
  AND U59 ( .A(o[1]), .B(n80), .Z(n78) );
  XOR U60 ( .A(n81), .B(n79), .Z(n80) );
  XNOR U61 ( .A(n82), .B(n83), .Z(o[21]) );
  AND U62 ( .A(o[1]), .B(n84), .Z(n82) );
  XOR U63 ( .A(n85), .B(n83), .Z(n84) );
  XNOR U64 ( .A(n86), .B(n87), .Z(o[20]) );
  AND U65 ( .A(o[1]), .B(n88), .Z(n86) );
  XOR U66 ( .A(n89), .B(n87), .Z(n88) );
  XNOR U67 ( .A(n90), .B(n91), .Z(o[19]) );
  AND U68 ( .A(o[1]), .B(n92), .Z(n90) );
  XOR U69 ( .A(n93), .B(n91), .Z(n92) );
  XNOR U70 ( .A(n94), .B(n95), .Z(o[18]) );
  AND U71 ( .A(o[1]), .B(n96), .Z(n94) );
  XOR U72 ( .A(n97), .B(n95), .Z(n96) );
  XNOR U73 ( .A(n98), .B(n99), .Z(o[17]) );
  AND U74 ( .A(o[1]), .B(n100), .Z(n98) );
  XOR U75 ( .A(n101), .B(n99), .Z(n100) );
  XNOR U76 ( .A(n102), .B(n103), .Z(o[16]) );
  AND U77 ( .A(o[1]), .B(n104), .Z(n102) );
  XOR U78 ( .A(n105), .B(n103), .Z(n104) );
  XNOR U79 ( .A(n106), .B(n107), .Z(o[15]) );
  AND U80 ( .A(o[1]), .B(n108), .Z(n106) );
  XOR U81 ( .A(n109), .B(n107), .Z(n108) );
  XNOR U82 ( .A(n110), .B(n111), .Z(o[14]) );
  AND U83 ( .A(o[1]), .B(n112), .Z(n110) );
  XOR U84 ( .A(n113), .B(n111), .Z(n112) );
  XNOR U85 ( .A(n114), .B(n115), .Z(o[13]) );
  AND U86 ( .A(o[1]), .B(n116), .Z(n114) );
  XOR U87 ( .A(n117), .B(n115), .Z(n116) );
  XNOR U88 ( .A(n118), .B(n119), .Z(o[12]) );
  AND U89 ( .A(o[1]), .B(n120), .Z(n118) );
  XOR U90 ( .A(n121), .B(n119), .Z(n120) );
  XNOR U91 ( .A(n122), .B(n123), .Z(o[11]) );
  AND U92 ( .A(o[1]), .B(n124), .Z(n122) );
  XOR U93 ( .A(n125), .B(n123), .Z(n124) );
  XNOR U94 ( .A(n126), .B(n127), .Z(o[10]) );
  AND U95 ( .A(o[1]), .B(n128), .Z(n126) );
  XOR U96 ( .A(n129), .B(n127), .Z(n128) );
  XOR U97 ( .A(n130), .B(n131), .Z(o[0]) );
  AND U98 ( .A(o[1]), .B(n132), .Z(n131) );
  XOR U99 ( .A(n130), .B(n133), .Z(n132) );
  XOR U100 ( .A(n134), .B(n135), .Z(o[1]) );
  AND U101 ( .A(n136), .B(n137), .Z(n135) );
  XOR U102 ( .A(n33), .B(n134), .Z(n137) );
  IV U103 ( .A(n138), .Z(n33) );
  AND U104 ( .A(p_input[95]), .B(p_input[127]), .Z(n138) );
  XOR U105 ( .A(n134), .B(n31), .Z(n136) );
  AND U106 ( .A(p_input[31]), .B(p_input[63]), .Z(n31) );
  XOR U107 ( .A(n139), .B(n140), .Z(n134) );
  AND U108 ( .A(n141), .B(n142), .Z(n140) );
  XOR U109 ( .A(n139), .B(n37), .Z(n142) );
  XNOR U110 ( .A(p_input[94]), .B(n143), .Z(n37) );
  AND U111 ( .A(n133), .B(n144), .Z(n143) );
  XOR U112 ( .A(p_input[94]), .B(p_input[126]), .Z(n144) );
  XNOR U113 ( .A(n35), .B(n139), .Z(n141) );
  XOR U114 ( .A(n145), .B(n146), .Z(n35) );
  AND U115 ( .A(n130), .B(n147), .Z(n146) );
  XOR U116 ( .A(p_input[62]), .B(p_input[30]), .Z(n147) );
  XOR U117 ( .A(n148), .B(n149), .Z(n139) );
  AND U118 ( .A(n150), .B(n151), .Z(n149) );
  XOR U119 ( .A(n148), .B(n41), .Z(n151) );
  XNOR U120 ( .A(p_input[93]), .B(n152), .Z(n41) );
  AND U121 ( .A(n133), .B(n153), .Z(n152) );
  XOR U122 ( .A(p_input[93]), .B(p_input[125]), .Z(n153) );
  XNOR U123 ( .A(n39), .B(n148), .Z(n150) );
  XOR U124 ( .A(n154), .B(n155), .Z(n39) );
  AND U125 ( .A(n130), .B(n156), .Z(n155) );
  XOR U126 ( .A(p_input[61]), .B(p_input[29]), .Z(n156) );
  XOR U127 ( .A(n157), .B(n158), .Z(n148) );
  AND U128 ( .A(n159), .B(n160), .Z(n158) );
  XOR U129 ( .A(n157), .B(n45), .Z(n160) );
  XNOR U130 ( .A(p_input[92]), .B(n161), .Z(n45) );
  AND U131 ( .A(n133), .B(n162), .Z(n161) );
  XOR U132 ( .A(p_input[92]), .B(p_input[124]), .Z(n162) );
  XNOR U133 ( .A(n43), .B(n157), .Z(n159) );
  XOR U134 ( .A(n163), .B(n164), .Z(n43) );
  AND U135 ( .A(n130), .B(n165), .Z(n164) );
  XOR U136 ( .A(p_input[60]), .B(p_input[28]), .Z(n165) );
  XOR U137 ( .A(n166), .B(n167), .Z(n157) );
  AND U138 ( .A(n168), .B(n169), .Z(n167) );
  XOR U139 ( .A(n166), .B(n53), .Z(n169) );
  XNOR U140 ( .A(p_input[91]), .B(n170), .Z(n53) );
  AND U141 ( .A(n133), .B(n171), .Z(n170) );
  XOR U142 ( .A(p_input[91]), .B(p_input[123]), .Z(n171) );
  XNOR U143 ( .A(n51), .B(n166), .Z(n168) );
  XOR U144 ( .A(n172), .B(n173), .Z(n51) );
  AND U145 ( .A(n130), .B(n174), .Z(n173) );
  XOR U146 ( .A(p_input[59]), .B(p_input[27]), .Z(n174) );
  XOR U147 ( .A(n175), .B(n176), .Z(n166) );
  AND U148 ( .A(n177), .B(n178), .Z(n176) );
  XOR U149 ( .A(n175), .B(n57), .Z(n178) );
  XNOR U150 ( .A(p_input[90]), .B(n179), .Z(n57) );
  AND U151 ( .A(n133), .B(n180), .Z(n179) );
  XOR U152 ( .A(p_input[90]), .B(p_input[122]), .Z(n180) );
  XNOR U153 ( .A(n55), .B(n175), .Z(n177) );
  XOR U154 ( .A(n181), .B(n182), .Z(n55) );
  AND U155 ( .A(n130), .B(n183), .Z(n182) );
  XOR U156 ( .A(p_input[58]), .B(p_input[26]), .Z(n183) );
  XOR U157 ( .A(n184), .B(n185), .Z(n175) );
  AND U158 ( .A(n186), .B(n187), .Z(n185) );
  XOR U159 ( .A(n184), .B(n61), .Z(n187) );
  XNOR U160 ( .A(p_input[89]), .B(n188), .Z(n61) );
  AND U161 ( .A(n133), .B(n189), .Z(n188) );
  XOR U162 ( .A(p_input[89]), .B(p_input[121]), .Z(n189) );
  XNOR U163 ( .A(n59), .B(n184), .Z(n186) );
  XOR U164 ( .A(n190), .B(n191), .Z(n59) );
  AND U165 ( .A(n130), .B(n192), .Z(n191) );
  XOR U166 ( .A(p_input[57]), .B(p_input[25]), .Z(n192) );
  XOR U167 ( .A(n193), .B(n194), .Z(n184) );
  AND U168 ( .A(n195), .B(n196), .Z(n194) );
  XOR U169 ( .A(n193), .B(n65), .Z(n196) );
  XNOR U170 ( .A(p_input[88]), .B(n197), .Z(n65) );
  AND U171 ( .A(n133), .B(n198), .Z(n197) );
  XOR U172 ( .A(p_input[88]), .B(p_input[120]), .Z(n198) );
  XNOR U173 ( .A(n63), .B(n193), .Z(n195) );
  XOR U174 ( .A(n199), .B(n200), .Z(n63) );
  AND U175 ( .A(n130), .B(n201), .Z(n200) );
  XOR U176 ( .A(p_input[56]), .B(p_input[24]), .Z(n201) );
  XOR U177 ( .A(n202), .B(n203), .Z(n193) );
  AND U178 ( .A(n204), .B(n205), .Z(n203) );
  XOR U179 ( .A(n202), .B(n69), .Z(n205) );
  XNOR U180 ( .A(p_input[87]), .B(n206), .Z(n69) );
  AND U181 ( .A(n133), .B(n207), .Z(n206) );
  XOR U182 ( .A(p_input[87]), .B(p_input[119]), .Z(n207) );
  XNOR U183 ( .A(n67), .B(n202), .Z(n204) );
  XOR U184 ( .A(n208), .B(n209), .Z(n67) );
  AND U185 ( .A(n130), .B(n210), .Z(n209) );
  XOR U186 ( .A(p_input[55]), .B(p_input[23]), .Z(n210) );
  XOR U187 ( .A(n211), .B(n212), .Z(n202) );
  AND U188 ( .A(n213), .B(n214), .Z(n212) );
  XOR U189 ( .A(n211), .B(n73), .Z(n214) );
  XNOR U190 ( .A(p_input[86]), .B(n215), .Z(n73) );
  AND U191 ( .A(n133), .B(n216), .Z(n215) );
  XOR U192 ( .A(p_input[86]), .B(p_input[118]), .Z(n216) );
  XNOR U193 ( .A(n71), .B(n211), .Z(n213) );
  XOR U194 ( .A(n217), .B(n218), .Z(n71) );
  AND U195 ( .A(n130), .B(n219), .Z(n218) );
  XOR U196 ( .A(p_input[54]), .B(p_input[22]), .Z(n219) );
  XOR U197 ( .A(n220), .B(n221), .Z(n211) );
  AND U198 ( .A(n222), .B(n223), .Z(n221) );
  XOR U199 ( .A(n220), .B(n77), .Z(n223) );
  XNOR U200 ( .A(p_input[85]), .B(n224), .Z(n77) );
  AND U201 ( .A(n133), .B(n225), .Z(n224) );
  XOR U202 ( .A(p_input[85]), .B(p_input[117]), .Z(n225) );
  XNOR U203 ( .A(n75), .B(n220), .Z(n222) );
  XOR U204 ( .A(n226), .B(n227), .Z(n75) );
  AND U205 ( .A(n130), .B(n228), .Z(n227) );
  XOR U206 ( .A(p_input[53]), .B(p_input[21]), .Z(n228) );
  XOR U207 ( .A(n229), .B(n230), .Z(n220) );
  AND U208 ( .A(n231), .B(n232), .Z(n230) );
  XOR U209 ( .A(n229), .B(n81), .Z(n232) );
  XNOR U210 ( .A(p_input[84]), .B(n233), .Z(n81) );
  AND U211 ( .A(n133), .B(n234), .Z(n233) );
  XOR U212 ( .A(p_input[84]), .B(p_input[116]), .Z(n234) );
  XNOR U213 ( .A(n79), .B(n229), .Z(n231) );
  XOR U214 ( .A(n235), .B(n236), .Z(n79) );
  AND U215 ( .A(n130), .B(n237), .Z(n236) );
  XOR U216 ( .A(p_input[52]), .B(p_input[20]), .Z(n237) );
  XOR U217 ( .A(n238), .B(n239), .Z(n229) );
  AND U218 ( .A(n240), .B(n241), .Z(n239) );
  XOR U219 ( .A(n238), .B(n85), .Z(n241) );
  XNOR U220 ( .A(p_input[83]), .B(n242), .Z(n85) );
  AND U221 ( .A(n133), .B(n243), .Z(n242) );
  XOR U222 ( .A(p_input[83]), .B(p_input[115]), .Z(n243) );
  XNOR U223 ( .A(n83), .B(n238), .Z(n240) );
  XOR U224 ( .A(n244), .B(n245), .Z(n83) );
  AND U225 ( .A(n130), .B(n246), .Z(n245) );
  XOR U226 ( .A(p_input[51]), .B(p_input[19]), .Z(n246) );
  XOR U227 ( .A(n247), .B(n248), .Z(n238) );
  AND U228 ( .A(n249), .B(n250), .Z(n248) );
  XOR U229 ( .A(n247), .B(n89), .Z(n250) );
  XNOR U230 ( .A(p_input[82]), .B(n251), .Z(n89) );
  AND U231 ( .A(n133), .B(n252), .Z(n251) );
  XOR U232 ( .A(p_input[82]), .B(p_input[114]), .Z(n252) );
  XNOR U233 ( .A(n87), .B(n247), .Z(n249) );
  XOR U234 ( .A(n253), .B(n254), .Z(n87) );
  AND U235 ( .A(n130), .B(n255), .Z(n254) );
  XOR U236 ( .A(p_input[50]), .B(p_input[18]), .Z(n255) );
  XOR U237 ( .A(n256), .B(n257), .Z(n247) );
  AND U238 ( .A(n258), .B(n259), .Z(n257) );
  XOR U239 ( .A(n256), .B(n93), .Z(n259) );
  XNOR U240 ( .A(p_input[81]), .B(n260), .Z(n93) );
  AND U241 ( .A(n133), .B(n261), .Z(n260) );
  XOR U242 ( .A(p_input[81]), .B(p_input[113]), .Z(n261) );
  XNOR U243 ( .A(n91), .B(n256), .Z(n258) );
  XOR U244 ( .A(n262), .B(n263), .Z(n91) );
  AND U245 ( .A(n130), .B(n264), .Z(n263) );
  XOR U246 ( .A(p_input[49]), .B(p_input[17]), .Z(n264) );
  XOR U247 ( .A(n265), .B(n266), .Z(n256) );
  AND U248 ( .A(n267), .B(n268), .Z(n266) );
  XOR U249 ( .A(n265), .B(n97), .Z(n268) );
  XNOR U250 ( .A(p_input[80]), .B(n269), .Z(n97) );
  AND U251 ( .A(n133), .B(n270), .Z(n269) );
  XOR U252 ( .A(p_input[80]), .B(p_input[112]), .Z(n270) );
  XNOR U253 ( .A(n95), .B(n265), .Z(n267) );
  XOR U254 ( .A(n271), .B(n272), .Z(n95) );
  AND U255 ( .A(n130), .B(n273), .Z(n272) );
  XOR U256 ( .A(p_input[48]), .B(p_input[16]), .Z(n273) );
  XOR U257 ( .A(n274), .B(n275), .Z(n265) );
  AND U258 ( .A(n276), .B(n277), .Z(n275) );
  XOR U259 ( .A(n274), .B(n101), .Z(n277) );
  XNOR U260 ( .A(p_input[79]), .B(n278), .Z(n101) );
  AND U261 ( .A(n133), .B(n279), .Z(n278) );
  XOR U262 ( .A(p_input[79]), .B(p_input[111]), .Z(n279) );
  XNOR U263 ( .A(n99), .B(n274), .Z(n276) );
  XOR U264 ( .A(n280), .B(n281), .Z(n99) );
  AND U265 ( .A(n130), .B(n282), .Z(n281) );
  XOR U266 ( .A(p_input[47]), .B(p_input[15]), .Z(n282) );
  XOR U267 ( .A(n283), .B(n284), .Z(n274) );
  AND U268 ( .A(n285), .B(n286), .Z(n284) );
  XOR U269 ( .A(n283), .B(n105), .Z(n286) );
  XNOR U270 ( .A(p_input[78]), .B(n287), .Z(n105) );
  AND U271 ( .A(n133), .B(n288), .Z(n287) );
  XOR U272 ( .A(p_input[78]), .B(p_input[110]), .Z(n288) );
  XNOR U273 ( .A(n103), .B(n283), .Z(n285) );
  XOR U274 ( .A(n289), .B(n290), .Z(n103) );
  AND U275 ( .A(n130), .B(n291), .Z(n290) );
  XOR U276 ( .A(p_input[46]), .B(p_input[14]), .Z(n291) );
  XOR U277 ( .A(n292), .B(n293), .Z(n283) );
  AND U278 ( .A(n294), .B(n295), .Z(n293) );
  XOR U279 ( .A(n292), .B(n109), .Z(n295) );
  XNOR U280 ( .A(p_input[77]), .B(n296), .Z(n109) );
  AND U281 ( .A(n133), .B(n297), .Z(n296) );
  XOR U282 ( .A(p_input[77]), .B(p_input[109]), .Z(n297) );
  XNOR U283 ( .A(n107), .B(n292), .Z(n294) );
  XOR U284 ( .A(n298), .B(n299), .Z(n107) );
  AND U285 ( .A(n130), .B(n300), .Z(n299) );
  XOR U286 ( .A(p_input[45]), .B(p_input[13]), .Z(n300) );
  XOR U287 ( .A(n301), .B(n302), .Z(n292) );
  AND U288 ( .A(n303), .B(n304), .Z(n302) );
  XOR U289 ( .A(n301), .B(n113), .Z(n304) );
  XNOR U290 ( .A(p_input[76]), .B(n305), .Z(n113) );
  AND U291 ( .A(n133), .B(n306), .Z(n305) );
  XOR U292 ( .A(p_input[76]), .B(p_input[108]), .Z(n306) );
  XNOR U293 ( .A(n111), .B(n301), .Z(n303) );
  XOR U294 ( .A(n307), .B(n308), .Z(n111) );
  AND U295 ( .A(n130), .B(n309), .Z(n308) );
  XOR U296 ( .A(p_input[44]), .B(p_input[12]), .Z(n309) );
  XOR U297 ( .A(n310), .B(n311), .Z(n301) );
  AND U298 ( .A(n312), .B(n313), .Z(n311) );
  XOR U299 ( .A(n310), .B(n117), .Z(n313) );
  XNOR U300 ( .A(p_input[75]), .B(n314), .Z(n117) );
  AND U301 ( .A(n133), .B(n315), .Z(n314) );
  XOR U302 ( .A(p_input[75]), .B(p_input[107]), .Z(n315) );
  XNOR U303 ( .A(n115), .B(n310), .Z(n312) );
  XOR U304 ( .A(n316), .B(n317), .Z(n115) );
  AND U305 ( .A(n130), .B(n318), .Z(n317) );
  XOR U306 ( .A(p_input[43]), .B(p_input[11]), .Z(n318) );
  XOR U307 ( .A(n319), .B(n320), .Z(n310) );
  AND U308 ( .A(n321), .B(n322), .Z(n320) );
  XOR U309 ( .A(n319), .B(n121), .Z(n322) );
  XNOR U310 ( .A(p_input[74]), .B(n323), .Z(n121) );
  AND U311 ( .A(n133), .B(n324), .Z(n323) );
  XOR U312 ( .A(p_input[74]), .B(p_input[106]), .Z(n324) );
  XNOR U313 ( .A(n119), .B(n319), .Z(n321) );
  XOR U314 ( .A(n325), .B(n326), .Z(n119) );
  AND U315 ( .A(n130), .B(n327), .Z(n326) );
  XOR U316 ( .A(p_input[42]), .B(p_input[10]), .Z(n327) );
  XOR U317 ( .A(n328), .B(n329), .Z(n319) );
  AND U318 ( .A(n330), .B(n331), .Z(n329) );
  XOR U319 ( .A(n328), .B(n125), .Z(n331) );
  XNOR U320 ( .A(p_input[73]), .B(n332), .Z(n125) );
  AND U321 ( .A(n133), .B(n333), .Z(n332) );
  XOR U322 ( .A(p_input[73]), .B(p_input[105]), .Z(n333) );
  XNOR U323 ( .A(n123), .B(n328), .Z(n330) );
  XOR U324 ( .A(n334), .B(n335), .Z(n123) );
  AND U325 ( .A(n130), .B(n336), .Z(n335) );
  XOR U326 ( .A(p_input[9]), .B(p_input[41]), .Z(n336) );
  XOR U327 ( .A(n337), .B(n338), .Z(n328) );
  AND U328 ( .A(n339), .B(n340), .Z(n338) );
  XOR U329 ( .A(n337), .B(n129), .Z(n340) );
  XNOR U330 ( .A(p_input[72]), .B(n341), .Z(n129) );
  AND U331 ( .A(n133), .B(n342), .Z(n341) );
  XOR U332 ( .A(p_input[72]), .B(p_input[104]), .Z(n342) );
  XNOR U333 ( .A(n127), .B(n337), .Z(n339) );
  XOR U334 ( .A(n343), .B(n344), .Z(n127) );
  AND U335 ( .A(n130), .B(n345), .Z(n344) );
  XOR U336 ( .A(p_input[8]), .B(p_input[40]), .Z(n345) );
  XOR U337 ( .A(n346), .B(n347), .Z(n337) );
  AND U338 ( .A(n348), .B(n349), .Z(n347) );
  XOR U339 ( .A(n4), .B(n346), .Z(n349) );
  XNOR U340 ( .A(p_input[71]), .B(n350), .Z(n4) );
  AND U341 ( .A(n133), .B(n351), .Z(n350) );
  XOR U342 ( .A(p_input[71]), .B(p_input[103]), .Z(n351) );
  XNOR U343 ( .A(n346), .B(n2), .Z(n348) );
  XOR U344 ( .A(n352), .B(n353), .Z(n2) );
  AND U345 ( .A(n130), .B(n354), .Z(n353) );
  XOR U346 ( .A(p_input[7]), .B(p_input[39]), .Z(n354) );
  XOR U347 ( .A(n355), .B(n356), .Z(n346) );
  AND U348 ( .A(n357), .B(n358), .Z(n356) );
  XOR U349 ( .A(n355), .B(n8), .Z(n358) );
  XNOR U350 ( .A(p_input[70]), .B(n359), .Z(n8) );
  AND U351 ( .A(n133), .B(n360), .Z(n359) );
  XOR U352 ( .A(p_input[70]), .B(p_input[102]), .Z(n360) );
  XNOR U353 ( .A(n6), .B(n355), .Z(n357) );
  XOR U354 ( .A(n361), .B(n362), .Z(n6) );
  AND U355 ( .A(n130), .B(n363), .Z(n362) );
  XOR U356 ( .A(p_input[6]), .B(p_input[38]), .Z(n363) );
  XOR U357 ( .A(n364), .B(n365), .Z(n355) );
  AND U358 ( .A(n366), .B(n367), .Z(n365) );
  XOR U359 ( .A(n364), .B(n12), .Z(n367) );
  XNOR U360 ( .A(p_input[69]), .B(n368), .Z(n12) );
  AND U361 ( .A(n133), .B(n369), .Z(n368) );
  XOR U362 ( .A(p_input[69]), .B(p_input[101]), .Z(n369) );
  XNOR U363 ( .A(n10), .B(n364), .Z(n366) );
  XOR U364 ( .A(n370), .B(n371), .Z(n10) );
  AND U365 ( .A(n130), .B(n372), .Z(n371) );
  XOR U366 ( .A(p_input[5]), .B(p_input[37]), .Z(n372) );
  XOR U367 ( .A(n373), .B(n374), .Z(n364) );
  AND U368 ( .A(n375), .B(n376), .Z(n374) );
  XOR U369 ( .A(n373), .B(n16), .Z(n376) );
  XNOR U370 ( .A(p_input[68]), .B(n377), .Z(n16) );
  AND U371 ( .A(n133), .B(n378), .Z(n377) );
  XOR U372 ( .A(p_input[68]), .B(p_input[100]), .Z(n378) );
  XNOR U373 ( .A(n14), .B(n373), .Z(n375) );
  XOR U374 ( .A(n379), .B(n380), .Z(n14) );
  AND U375 ( .A(n130), .B(n381), .Z(n380) );
  XOR U376 ( .A(p_input[4]), .B(p_input[36]), .Z(n381) );
  XOR U377 ( .A(n382), .B(n383), .Z(n373) );
  AND U378 ( .A(n384), .B(n385), .Z(n383) );
  XOR U379 ( .A(n382), .B(n20), .Z(n385) );
  XNOR U380 ( .A(p_input[67]), .B(n386), .Z(n20) );
  AND U381 ( .A(n133), .B(n387), .Z(n386) );
  XOR U382 ( .A(p_input[99]), .B(p_input[67]), .Z(n387) );
  XNOR U383 ( .A(n18), .B(n382), .Z(n384) );
  XOR U384 ( .A(n388), .B(n389), .Z(n18) );
  AND U385 ( .A(n130), .B(n390), .Z(n389) );
  XOR U386 ( .A(p_input[3]), .B(p_input[35]), .Z(n390) );
  XOR U387 ( .A(n391), .B(n392), .Z(n382) );
  AND U388 ( .A(n393), .B(n394), .Z(n392) );
  XOR U389 ( .A(n391), .B(n24), .Z(n394) );
  XNOR U390 ( .A(p_input[66]), .B(n395), .Z(n24) );
  AND U391 ( .A(n133), .B(n396), .Z(n395) );
  XOR U392 ( .A(p_input[98]), .B(p_input[66]), .Z(n396) );
  XNOR U393 ( .A(n22), .B(n391), .Z(n393) );
  XOR U394 ( .A(n397), .B(n398), .Z(n22) );
  AND U395 ( .A(n130), .B(n399), .Z(n398) );
  XOR U396 ( .A(p_input[34]), .B(p_input[2]), .Z(n399) );
  XNOR U397 ( .A(n400), .B(n401), .Z(n391) );
  AND U398 ( .A(n402), .B(n403), .Z(n401) );
  XNOR U399 ( .A(n400), .B(n28), .Z(n403) );
  XNOR U400 ( .A(p_input[65]), .B(n404), .Z(n28) );
  AND U401 ( .A(n133), .B(n405), .Z(n404) );
  XNOR U402 ( .A(p_input[97]), .B(n406), .Z(n405) );
  IV U403 ( .A(p_input[65]), .Z(n406) );
  XOR U404 ( .A(n29), .B(n400), .Z(n402) );
  IV U405 ( .A(n26), .Z(n29) );
  XOR U406 ( .A(p_input[1]), .B(n407), .Z(n26) );
  AND U407 ( .A(n130), .B(n408), .Z(n407) );
  XOR U408 ( .A(p_input[33]), .B(p_input[1]), .Z(n408) );
  AND U409 ( .A(n47), .B(n49), .Z(n400) );
  XOR U410 ( .A(p_input[64]), .B(n409), .Z(n49) );
  AND U411 ( .A(n133), .B(n410), .Z(n409) );
  XOR U412 ( .A(p_input[96]), .B(p_input[64]), .Z(n410) );
  XOR U413 ( .A(n411), .B(n412), .Z(n133) );
  AND U414 ( .A(n413), .B(n414), .Z(n412) );
  XNOR U415 ( .A(p_input[127]), .B(n411), .Z(n414) );
  XOR U416 ( .A(n411), .B(p_input[95]), .Z(n413) );
  XOR U417 ( .A(n415), .B(n416), .Z(n411) );
  AND U418 ( .A(n417), .B(n418), .Z(n416) );
  XNOR U419 ( .A(p_input[126]), .B(n415), .Z(n418) );
  XOR U420 ( .A(n415), .B(p_input[94]), .Z(n417) );
  XOR U421 ( .A(n419), .B(n420), .Z(n415) );
  AND U422 ( .A(n421), .B(n422), .Z(n420) );
  XNOR U423 ( .A(p_input[125]), .B(n419), .Z(n422) );
  XOR U424 ( .A(n419), .B(p_input[93]), .Z(n421) );
  XOR U425 ( .A(n423), .B(n424), .Z(n419) );
  AND U426 ( .A(n425), .B(n426), .Z(n424) );
  XNOR U427 ( .A(p_input[124]), .B(n423), .Z(n426) );
  XOR U428 ( .A(n423), .B(p_input[92]), .Z(n425) );
  XOR U429 ( .A(n427), .B(n428), .Z(n423) );
  AND U430 ( .A(n429), .B(n430), .Z(n428) );
  XNOR U431 ( .A(p_input[123]), .B(n427), .Z(n430) );
  XOR U432 ( .A(n427), .B(p_input[91]), .Z(n429) );
  XOR U433 ( .A(n431), .B(n432), .Z(n427) );
  AND U434 ( .A(n433), .B(n434), .Z(n432) );
  XNOR U435 ( .A(p_input[122]), .B(n431), .Z(n434) );
  XOR U436 ( .A(n431), .B(p_input[90]), .Z(n433) );
  XOR U437 ( .A(n435), .B(n436), .Z(n431) );
  AND U438 ( .A(n437), .B(n438), .Z(n436) );
  XNOR U439 ( .A(p_input[121]), .B(n435), .Z(n438) );
  XOR U440 ( .A(n435), .B(p_input[89]), .Z(n437) );
  XOR U441 ( .A(n439), .B(n440), .Z(n435) );
  AND U442 ( .A(n441), .B(n442), .Z(n440) );
  XNOR U443 ( .A(p_input[120]), .B(n439), .Z(n442) );
  XOR U444 ( .A(n439), .B(p_input[88]), .Z(n441) );
  XOR U445 ( .A(n443), .B(n444), .Z(n439) );
  AND U446 ( .A(n445), .B(n446), .Z(n444) );
  XNOR U447 ( .A(p_input[119]), .B(n443), .Z(n446) );
  XOR U448 ( .A(n443), .B(p_input[87]), .Z(n445) );
  XOR U449 ( .A(n447), .B(n448), .Z(n443) );
  AND U450 ( .A(n449), .B(n450), .Z(n448) );
  XNOR U451 ( .A(p_input[118]), .B(n447), .Z(n450) );
  XOR U452 ( .A(n447), .B(p_input[86]), .Z(n449) );
  XOR U453 ( .A(n451), .B(n452), .Z(n447) );
  AND U454 ( .A(n453), .B(n454), .Z(n452) );
  XNOR U455 ( .A(p_input[117]), .B(n451), .Z(n454) );
  XOR U456 ( .A(n451), .B(p_input[85]), .Z(n453) );
  XOR U457 ( .A(n455), .B(n456), .Z(n451) );
  AND U458 ( .A(n457), .B(n458), .Z(n456) );
  XNOR U459 ( .A(p_input[116]), .B(n455), .Z(n458) );
  XOR U460 ( .A(n455), .B(p_input[84]), .Z(n457) );
  XOR U461 ( .A(n459), .B(n460), .Z(n455) );
  AND U462 ( .A(n461), .B(n462), .Z(n460) );
  XNOR U463 ( .A(p_input[115]), .B(n459), .Z(n462) );
  XOR U464 ( .A(n459), .B(p_input[83]), .Z(n461) );
  XOR U465 ( .A(n463), .B(n464), .Z(n459) );
  AND U466 ( .A(n465), .B(n466), .Z(n464) );
  XNOR U467 ( .A(p_input[114]), .B(n463), .Z(n466) );
  XOR U468 ( .A(n463), .B(p_input[82]), .Z(n465) );
  XOR U469 ( .A(n467), .B(n468), .Z(n463) );
  AND U470 ( .A(n469), .B(n470), .Z(n468) );
  XNOR U471 ( .A(p_input[113]), .B(n467), .Z(n470) );
  XOR U472 ( .A(n467), .B(p_input[81]), .Z(n469) );
  XOR U473 ( .A(n471), .B(n472), .Z(n467) );
  AND U474 ( .A(n473), .B(n474), .Z(n472) );
  XNOR U475 ( .A(p_input[112]), .B(n471), .Z(n474) );
  XOR U476 ( .A(n471), .B(p_input[80]), .Z(n473) );
  XOR U477 ( .A(n475), .B(n476), .Z(n471) );
  AND U478 ( .A(n477), .B(n478), .Z(n476) );
  XNOR U479 ( .A(p_input[111]), .B(n475), .Z(n478) );
  XOR U480 ( .A(n475), .B(p_input[79]), .Z(n477) );
  XOR U481 ( .A(n479), .B(n480), .Z(n475) );
  AND U482 ( .A(n481), .B(n482), .Z(n480) );
  XNOR U483 ( .A(p_input[110]), .B(n479), .Z(n482) );
  XOR U484 ( .A(n479), .B(p_input[78]), .Z(n481) );
  XOR U485 ( .A(n483), .B(n484), .Z(n479) );
  AND U486 ( .A(n485), .B(n486), .Z(n484) );
  XNOR U487 ( .A(p_input[109]), .B(n483), .Z(n486) );
  XOR U488 ( .A(n483), .B(p_input[77]), .Z(n485) );
  XOR U489 ( .A(n487), .B(n488), .Z(n483) );
  AND U490 ( .A(n489), .B(n490), .Z(n488) );
  XNOR U491 ( .A(p_input[108]), .B(n487), .Z(n490) );
  XOR U492 ( .A(n487), .B(p_input[76]), .Z(n489) );
  XOR U493 ( .A(n491), .B(n492), .Z(n487) );
  AND U494 ( .A(n493), .B(n494), .Z(n492) );
  XNOR U495 ( .A(p_input[107]), .B(n491), .Z(n494) );
  XOR U496 ( .A(n491), .B(p_input[75]), .Z(n493) );
  XOR U497 ( .A(n495), .B(n496), .Z(n491) );
  AND U498 ( .A(n497), .B(n498), .Z(n496) );
  XNOR U499 ( .A(p_input[106]), .B(n495), .Z(n498) );
  XOR U500 ( .A(n495), .B(p_input[74]), .Z(n497) );
  XOR U501 ( .A(n499), .B(n500), .Z(n495) );
  AND U502 ( .A(n501), .B(n502), .Z(n500) );
  XNOR U503 ( .A(p_input[105]), .B(n499), .Z(n502) );
  XOR U504 ( .A(n499), .B(p_input[73]), .Z(n501) );
  XOR U505 ( .A(n503), .B(n504), .Z(n499) );
  AND U506 ( .A(n505), .B(n506), .Z(n504) );
  XNOR U507 ( .A(p_input[104]), .B(n503), .Z(n506) );
  XOR U508 ( .A(n503), .B(p_input[72]), .Z(n505) );
  XOR U509 ( .A(n507), .B(n508), .Z(n503) );
  AND U510 ( .A(n509), .B(n510), .Z(n508) );
  XNOR U511 ( .A(p_input[103]), .B(n507), .Z(n510) );
  XOR U512 ( .A(n507), .B(p_input[71]), .Z(n509) );
  XOR U513 ( .A(n511), .B(n512), .Z(n507) );
  AND U514 ( .A(n513), .B(n514), .Z(n512) );
  XNOR U515 ( .A(p_input[102]), .B(n511), .Z(n514) );
  XOR U516 ( .A(n511), .B(p_input[70]), .Z(n513) );
  XOR U517 ( .A(n515), .B(n516), .Z(n511) );
  AND U518 ( .A(n517), .B(n518), .Z(n516) );
  XNOR U519 ( .A(p_input[101]), .B(n515), .Z(n518) );
  XOR U520 ( .A(n515), .B(p_input[69]), .Z(n517) );
  XOR U521 ( .A(n519), .B(n520), .Z(n515) );
  AND U522 ( .A(n521), .B(n522), .Z(n520) );
  XNOR U523 ( .A(p_input[100]), .B(n519), .Z(n522) );
  XOR U524 ( .A(n519), .B(p_input[68]), .Z(n521) );
  XOR U525 ( .A(n523), .B(n524), .Z(n519) );
  AND U526 ( .A(n525), .B(n526), .Z(n524) );
  XNOR U527 ( .A(p_input[99]), .B(n523), .Z(n526) );
  XOR U528 ( .A(n523), .B(p_input[67]), .Z(n525) );
  XOR U529 ( .A(n527), .B(n528), .Z(n523) );
  AND U530 ( .A(n529), .B(n530), .Z(n528) );
  XNOR U531 ( .A(p_input[98]), .B(n527), .Z(n530) );
  XOR U532 ( .A(n527), .B(p_input[66]), .Z(n529) );
  XNOR U533 ( .A(n531), .B(n532), .Z(n527) );
  AND U534 ( .A(n533), .B(n534), .Z(n532) );
  XOR U535 ( .A(p_input[97]), .B(n531), .Z(n534) );
  XNOR U536 ( .A(p_input[65]), .B(n531), .Z(n533) );
  AND U537 ( .A(p_input[96]), .B(n535), .Z(n531) );
  IV U538 ( .A(p_input[64]), .Z(n535) );
  XNOR U539 ( .A(p_input[0]), .B(n536), .Z(n47) );
  AND U540 ( .A(n130), .B(n537), .Z(n536) );
  XOR U541 ( .A(p_input[32]), .B(p_input[0]), .Z(n537) );
  XOR U542 ( .A(n538), .B(n539), .Z(n130) );
  AND U543 ( .A(n540), .B(n541), .Z(n539) );
  XNOR U544 ( .A(p_input[63]), .B(n538), .Z(n541) );
  XOR U545 ( .A(n538), .B(p_input[31]), .Z(n540) );
  XOR U546 ( .A(n542), .B(n543), .Z(n538) );
  AND U547 ( .A(n544), .B(n545), .Z(n543) );
  XNOR U548 ( .A(p_input[62]), .B(n542), .Z(n545) );
  XNOR U549 ( .A(n542), .B(n145), .Z(n544) );
  IV U550 ( .A(p_input[30]), .Z(n145) );
  XOR U551 ( .A(n546), .B(n547), .Z(n542) );
  AND U552 ( .A(n548), .B(n549), .Z(n547) );
  XNOR U553 ( .A(p_input[61]), .B(n546), .Z(n549) );
  XNOR U554 ( .A(n546), .B(n154), .Z(n548) );
  IV U555 ( .A(p_input[29]), .Z(n154) );
  XOR U556 ( .A(n550), .B(n551), .Z(n546) );
  AND U557 ( .A(n552), .B(n553), .Z(n551) );
  XNOR U558 ( .A(p_input[60]), .B(n550), .Z(n553) );
  XNOR U559 ( .A(n550), .B(n163), .Z(n552) );
  IV U560 ( .A(p_input[28]), .Z(n163) );
  XOR U561 ( .A(n554), .B(n555), .Z(n550) );
  AND U562 ( .A(n556), .B(n557), .Z(n555) );
  XNOR U563 ( .A(p_input[59]), .B(n554), .Z(n557) );
  XNOR U564 ( .A(n554), .B(n172), .Z(n556) );
  IV U565 ( .A(p_input[27]), .Z(n172) );
  XOR U566 ( .A(n558), .B(n559), .Z(n554) );
  AND U567 ( .A(n560), .B(n561), .Z(n559) );
  XNOR U568 ( .A(p_input[58]), .B(n558), .Z(n561) );
  XNOR U569 ( .A(n558), .B(n181), .Z(n560) );
  IV U570 ( .A(p_input[26]), .Z(n181) );
  XOR U571 ( .A(n562), .B(n563), .Z(n558) );
  AND U572 ( .A(n564), .B(n565), .Z(n563) );
  XNOR U573 ( .A(p_input[57]), .B(n562), .Z(n565) );
  XNOR U574 ( .A(n562), .B(n190), .Z(n564) );
  IV U575 ( .A(p_input[25]), .Z(n190) );
  XOR U576 ( .A(n566), .B(n567), .Z(n562) );
  AND U577 ( .A(n568), .B(n569), .Z(n567) );
  XNOR U578 ( .A(p_input[56]), .B(n566), .Z(n569) );
  XNOR U579 ( .A(n566), .B(n199), .Z(n568) );
  IV U580 ( .A(p_input[24]), .Z(n199) );
  XOR U581 ( .A(n570), .B(n571), .Z(n566) );
  AND U582 ( .A(n572), .B(n573), .Z(n571) );
  XNOR U583 ( .A(p_input[55]), .B(n570), .Z(n573) );
  XNOR U584 ( .A(n570), .B(n208), .Z(n572) );
  IV U585 ( .A(p_input[23]), .Z(n208) );
  XOR U586 ( .A(n574), .B(n575), .Z(n570) );
  AND U587 ( .A(n576), .B(n577), .Z(n575) );
  XNOR U588 ( .A(p_input[54]), .B(n574), .Z(n577) );
  XNOR U589 ( .A(n574), .B(n217), .Z(n576) );
  IV U590 ( .A(p_input[22]), .Z(n217) );
  XOR U591 ( .A(n578), .B(n579), .Z(n574) );
  AND U592 ( .A(n580), .B(n581), .Z(n579) );
  XNOR U593 ( .A(p_input[53]), .B(n578), .Z(n581) );
  XNOR U594 ( .A(n578), .B(n226), .Z(n580) );
  IV U595 ( .A(p_input[21]), .Z(n226) );
  XOR U596 ( .A(n582), .B(n583), .Z(n578) );
  AND U597 ( .A(n584), .B(n585), .Z(n583) );
  XNOR U598 ( .A(p_input[52]), .B(n582), .Z(n585) );
  XNOR U599 ( .A(n582), .B(n235), .Z(n584) );
  IV U600 ( .A(p_input[20]), .Z(n235) );
  XOR U601 ( .A(n586), .B(n587), .Z(n582) );
  AND U602 ( .A(n588), .B(n589), .Z(n587) );
  XNOR U603 ( .A(p_input[51]), .B(n586), .Z(n589) );
  XNOR U604 ( .A(n586), .B(n244), .Z(n588) );
  IV U605 ( .A(p_input[19]), .Z(n244) );
  XOR U606 ( .A(n590), .B(n591), .Z(n586) );
  AND U607 ( .A(n592), .B(n593), .Z(n591) );
  XNOR U608 ( .A(p_input[50]), .B(n590), .Z(n593) );
  XNOR U609 ( .A(n590), .B(n253), .Z(n592) );
  IV U610 ( .A(p_input[18]), .Z(n253) );
  XOR U611 ( .A(n594), .B(n595), .Z(n590) );
  AND U612 ( .A(n596), .B(n597), .Z(n595) );
  XNOR U613 ( .A(p_input[49]), .B(n594), .Z(n597) );
  XNOR U614 ( .A(n594), .B(n262), .Z(n596) );
  IV U615 ( .A(p_input[17]), .Z(n262) );
  XOR U616 ( .A(n598), .B(n599), .Z(n594) );
  AND U617 ( .A(n600), .B(n601), .Z(n599) );
  XNOR U618 ( .A(p_input[48]), .B(n598), .Z(n601) );
  XNOR U619 ( .A(n598), .B(n271), .Z(n600) );
  IV U620 ( .A(p_input[16]), .Z(n271) );
  XOR U621 ( .A(n602), .B(n603), .Z(n598) );
  AND U622 ( .A(n604), .B(n605), .Z(n603) );
  XNOR U623 ( .A(p_input[47]), .B(n602), .Z(n605) );
  XNOR U624 ( .A(n602), .B(n280), .Z(n604) );
  IV U625 ( .A(p_input[15]), .Z(n280) );
  XOR U626 ( .A(n606), .B(n607), .Z(n602) );
  AND U627 ( .A(n608), .B(n609), .Z(n607) );
  XNOR U628 ( .A(p_input[46]), .B(n606), .Z(n609) );
  XNOR U629 ( .A(n606), .B(n289), .Z(n608) );
  IV U630 ( .A(p_input[14]), .Z(n289) );
  XOR U631 ( .A(n610), .B(n611), .Z(n606) );
  AND U632 ( .A(n612), .B(n613), .Z(n611) );
  XNOR U633 ( .A(p_input[45]), .B(n610), .Z(n613) );
  XNOR U634 ( .A(n610), .B(n298), .Z(n612) );
  IV U635 ( .A(p_input[13]), .Z(n298) );
  XOR U636 ( .A(n614), .B(n615), .Z(n610) );
  AND U637 ( .A(n616), .B(n617), .Z(n615) );
  XNOR U638 ( .A(p_input[44]), .B(n614), .Z(n617) );
  XNOR U639 ( .A(n614), .B(n307), .Z(n616) );
  IV U640 ( .A(p_input[12]), .Z(n307) );
  XOR U641 ( .A(n618), .B(n619), .Z(n614) );
  AND U642 ( .A(n620), .B(n621), .Z(n619) );
  XNOR U643 ( .A(p_input[43]), .B(n618), .Z(n621) );
  XNOR U644 ( .A(n618), .B(n316), .Z(n620) );
  IV U645 ( .A(p_input[11]), .Z(n316) );
  XOR U646 ( .A(n622), .B(n623), .Z(n618) );
  AND U647 ( .A(n624), .B(n625), .Z(n623) );
  XNOR U648 ( .A(p_input[42]), .B(n622), .Z(n625) );
  XNOR U649 ( .A(n622), .B(n325), .Z(n624) );
  IV U650 ( .A(p_input[10]), .Z(n325) );
  XOR U651 ( .A(n626), .B(n627), .Z(n622) );
  AND U652 ( .A(n628), .B(n629), .Z(n627) );
  XNOR U653 ( .A(p_input[41]), .B(n626), .Z(n629) );
  XNOR U654 ( .A(n626), .B(n334), .Z(n628) );
  IV U655 ( .A(p_input[9]), .Z(n334) );
  XOR U656 ( .A(n630), .B(n631), .Z(n626) );
  AND U657 ( .A(n632), .B(n633), .Z(n631) );
  XNOR U658 ( .A(p_input[40]), .B(n630), .Z(n633) );
  XNOR U659 ( .A(n630), .B(n343), .Z(n632) );
  IV U660 ( .A(p_input[8]), .Z(n343) );
  XOR U661 ( .A(n634), .B(n635), .Z(n630) );
  AND U662 ( .A(n636), .B(n637), .Z(n635) );
  XNOR U663 ( .A(p_input[39]), .B(n634), .Z(n637) );
  XNOR U664 ( .A(n634), .B(n352), .Z(n636) );
  IV U665 ( .A(p_input[7]), .Z(n352) );
  XOR U666 ( .A(n638), .B(n639), .Z(n634) );
  AND U667 ( .A(n640), .B(n641), .Z(n639) );
  XNOR U668 ( .A(p_input[38]), .B(n638), .Z(n641) );
  XNOR U669 ( .A(n638), .B(n361), .Z(n640) );
  IV U670 ( .A(p_input[6]), .Z(n361) );
  XOR U671 ( .A(n642), .B(n643), .Z(n638) );
  AND U672 ( .A(n644), .B(n645), .Z(n643) );
  XNOR U673 ( .A(p_input[37]), .B(n642), .Z(n645) );
  XNOR U674 ( .A(n642), .B(n370), .Z(n644) );
  IV U675 ( .A(p_input[5]), .Z(n370) );
  XOR U676 ( .A(n646), .B(n647), .Z(n642) );
  AND U677 ( .A(n648), .B(n649), .Z(n647) );
  XNOR U678 ( .A(p_input[36]), .B(n646), .Z(n649) );
  XNOR U679 ( .A(n646), .B(n379), .Z(n648) );
  IV U680 ( .A(p_input[4]), .Z(n379) );
  XOR U681 ( .A(n650), .B(n651), .Z(n646) );
  AND U682 ( .A(n652), .B(n653), .Z(n651) );
  XNOR U683 ( .A(p_input[35]), .B(n650), .Z(n653) );
  XNOR U684 ( .A(n650), .B(n388), .Z(n652) );
  IV U685 ( .A(p_input[3]), .Z(n388) );
  XOR U686 ( .A(n654), .B(n655), .Z(n650) );
  AND U687 ( .A(n656), .B(n657), .Z(n655) );
  XNOR U688 ( .A(p_input[34]), .B(n654), .Z(n657) );
  XNOR U689 ( .A(n654), .B(n397), .Z(n656) );
  IV U690 ( .A(p_input[2]), .Z(n397) );
  XNOR U691 ( .A(n658), .B(n659), .Z(n654) );
  AND U692 ( .A(n660), .B(n661), .Z(n659) );
  XOR U693 ( .A(p_input[33]), .B(n658), .Z(n661) );
  XNOR U694 ( .A(p_input[1]), .B(n658), .Z(n660) );
  AND U695 ( .A(p_input[32]), .B(n662), .Z(n658) );
  IV U696 ( .A(p_input[0]), .Z(n662) );
endmodule

