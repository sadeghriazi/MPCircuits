
module knn_comb_BMR_W16_K3_N8 ( p_input, o );
  input [143:0] p_input;
  output [47:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760;
  assign \knn_comb_/min_val_out[0][0]  = p_input[112];
  assign \knn_comb_/min_val_out[0][1]  = p_input[113];
  assign \knn_comb_/min_val_out[0][2]  = p_input[114];
  assign \knn_comb_/min_val_out[0][3]  = p_input[115];
  assign \knn_comb_/min_val_out[0][4]  = p_input[116];
  assign \knn_comb_/min_val_out[0][5]  = p_input[117];
  assign \knn_comb_/min_val_out[0][6]  = p_input[118];
  assign \knn_comb_/min_val_out[0][7]  = p_input[119];
  assign \knn_comb_/min_val_out[0][8]  = p_input[120];
  assign \knn_comb_/min_val_out[0][9]  = p_input[121];
  assign \knn_comb_/min_val_out[0][10]  = p_input[122];
  assign \knn_comb_/min_val_out[0][11]  = p_input[123];
  assign \knn_comb_/min_val_out[0][12]  = p_input[124];
  assign \knn_comb_/min_val_out[0][13]  = p_input[125];
  assign \knn_comb_/min_val_out[0][14]  = p_input[126];
  assign \knn_comb_/min_val_out[0][15]  = p_input[127];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][0]  = p_input[80];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][1]  = p_input[81];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][2]  = p_input[82];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][3]  = p_input[83];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][4]  = p_input[84];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][5]  = p_input[85];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][6]  = p_input[86];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][7]  = p_input[87];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][8]  = p_input[88];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][9]  = p_input[89];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][10]  = p_input[90];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][11]  = p_input[91];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][12]  = p_input[92];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][13]  = p_input[93];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][14]  = p_input[94];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][15]  = p_input[95];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[96];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[97];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[98];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[99];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[100];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[101];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[102];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[103];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[104];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[105];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[106];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[107];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[108];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[109];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[110];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[111];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[8]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[7]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[6]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[5]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[4]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[47]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[46]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[45]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[44]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[43]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[42]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[41]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[40]) );
  XOR U15 ( .A(n29), .B(n30), .Z(o[3]) );
  XOR U16 ( .A(n31), .B(n32), .Z(o[39]) );
  XOR U17 ( .A(n33), .B(n34), .Z(o[38]) );
  XOR U18 ( .A(n35), .B(n36), .Z(o[37]) );
  XOR U19 ( .A(n37), .B(n38), .Z(o[36]) );
  XOR U20 ( .A(n39), .B(n40), .Z(o[35]) );
  XOR U21 ( .A(n41), .B(n42), .Z(o[34]) );
  XOR U22 ( .A(n43), .B(n44), .Z(o[33]) );
  XOR U23 ( .A(n45), .B(n46), .Z(o[32]) );
  XOR U24 ( .A(n47), .B(n48), .Z(o[31]) );
  XOR U25 ( .A(n49), .B(n50), .Z(o[30]) );
  XOR U26 ( .A(n51), .B(n52), .Z(o[2]) );
  XOR U27 ( .A(n53), .B(n54), .Z(o[29]) );
  XOR U28 ( .A(n55), .B(n56), .Z(o[28]) );
  XOR U29 ( .A(n57), .B(n58), .Z(o[27]) );
  XOR U30 ( .A(n59), .B(n60), .Z(o[26]) );
  XOR U31 ( .A(n1), .B(n61), .Z(o[25]) );
  AND U32 ( .A(n62), .B(n63), .Z(n1) );
  XOR U33 ( .A(n2), .B(n61), .Z(n63) );
  XOR U34 ( .A(n64), .B(n25), .Z(n61) );
  AND U35 ( .A(n65), .B(n66), .Z(n25) );
  XNOR U36 ( .A(n67), .B(n26), .Z(n66) );
  XOR U37 ( .A(n68), .B(n69), .Z(n26) );
  AND U38 ( .A(n70), .B(n71), .Z(n69) );
  XOR U39 ( .A(p_input[9]), .B(n68), .Z(n71) );
  XOR U40 ( .A(n72), .B(n73), .Z(n68) );
  AND U41 ( .A(n74), .B(n75), .Z(n73) );
  IV U42 ( .A(n64), .Z(n67) );
  XOR U43 ( .A(n76), .B(n77), .Z(n64) );
  AND U44 ( .A(n78), .B(n79), .Z(n77) );
  XOR U45 ( .A(n80), .B(n81), .Z(n2) );
  AND U46 ( .A(n82), .B(n79), .Z(n81) );
  XNOR U47 ( .A(n83), .B(n76), .Z(n79) );
  XOR U48 ( .A(n84), .B(n85), .Z(n76) );
  AND U49 ( .A(n86), .B(n75), .Z(n85) );
  XNOR U50 ( .A(n87), .B(n72), .Z(n75) );
  XOR U51 ( .A(n88), .B(n89), .Z(n72) );
  AND U52 ( .A(n90), .B(n91), .Z(n89) );
  XOR U53 ( .A(p_input[25]), .B(n88), .Z(n91) );
  XOR U54 ( .A(n92), .B(n93), .Z(n88) );
  AND U55 ( .A(n94), .B(n95), .Z(n93) );
  IV U56 ( .A(n84), .Z(n87) );
  XOR U57 ( .A(n96), .B(n97), .Z(n84) );
  AND U58 ( .A(n98), .B(n99), .Z(n97) );
  IV U59 ( .A(n80), .Z(n83) );
  XNOR U60 ( .A(n100), .B(n101), .Z(n80) );
  AND U61 ( .A(n102), .B(n99), .Z(n101) );
  XNOR U62 ( .A(n100), .B(n96), .Z(n99) );
  XOR U63 ( .A(n103), .B(n104), .Z(n96) );
  AND U64 ( .A(n105), .B(n95), .Z(n104) );
  XNOR U65 ( .A(n106), .B(n92), .Z(n95) );
  XOR U66 ( .A(n107), .B(n108), .Z(n92) );
  AND U67 ( .A(n109), .B(n110), .Z(n108) );
  XOR U68 ( .A(p_input[41]), .B(n107), .Z(n110) );
  XOR U69 ( .A(n111), .B(n112), .Z(n107) );
  AND U70 ( .A(n113), .B(n114), .Z(n112) );
  IV U71 ( .A(n103), .Z(n106) );
  XOR U72 ( .A(n115), .B(n116), .Z(n103) );
  AND U73 ( .A(n117), .B(n118), .Z(n116) );
  XOR U74 ( .A(n119), .B(n120), .Z(n100) );
  AND U75 ( .A(n121), .B(n118), .Z(n120) );
  XNOR U76 ( .A(n119), .B(n115), .Z(n118) );
  XOR U77 ( .A(n122), .B(n123), .Z(n115) );
  AND U78 ( .A(n124), .B(n114), .Z(n123) );
  XNOR U79 ( .A(n125), .B(n111), .Z(n114) );
  XOR U80 ( .A(n126), .B(n127), .Z(n111) );
  AND U81 ( .A(n128), .B(n129), .Z(n127) );
  XOR U82 ( .A(p_input[57]), .B(n126), .Z(n129) );
  XOR U83 ( .A(n130), .B(n131), .Z(n126) );
  AND U84 ( .A(n132), .B(n133), .Z(n131) );
  IV U85 ( .A(n122), .Z(n125) );
  XOR U86 ( .A(n134), .B(n135), .Z(n122) );
  AND U87 ( .A(n136), .B(n137), .Z(n135) );
  XOR U88 ( .A(n138), .B(n139), .Z(n119) );
  AND U89 ( .A(n140), .B(n137), .Z(n139) );
  XNOR U90 ( .A(n138), .B(n134), .Z(n137) );
  XOR U91 ( .A(n141), .B(n142), .Z(n134) );
  AND U92 ( .A(n143), .B(n133), .Z(n142) );
  XNOR U93 ( .A(n144), .B(n130), .Z(n133) );
  XOR U94 ( .A(n145), .B(n146), .Z(n130) );
  AND U95 ( .A(n147), .B(n148), .Z(n146) );
  XOR U96 ( .A(p_input[73]), .B(n145), .Z(n148) );
  XOR U97 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n149), .Z(
        n145) );
  AND U98 ( .A(n150), .B(n151), .Z(n149) );
  IV U99 ( .A(n141), .Z(n144) );
  XOR U100 ( .A(n152), .B(n153), .Z(n141) );
  AND U101 ( .A(n154), .B(n155), .Z(n153) );
  XOR U102 ( .A(n156), .B(n157), .Z(n138) );
  AND U103 ( .A(n158), .B(n155), .Z(n157) );
  XNOR U104 ( .A(n156), .B(n152), .Z(n155) );
  XNOR U105 ( .A(n159), .B(n160), .Z(n152) );
  AND U106 ( .A(n161), .B(n151), .Z(n160) );
  XNOR U107 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n159), .Z(
        n151) );
  XNOR U108 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .B(n162), .Z(
        n159) );
  AND U109 ( .A(n163), .B(n164), .Z(n162) );
  XNOR U110 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n165), .Z(n156) );
  AND U111 ( .A(n166), .B(n164), .Z(n165) );
  XOR U112 ( .A(n167), .B(n168), .Z(n164) );
  XOR U113 ( .A(n3), .B(n169), .Z(o[24]) );
  AND U114 ( .A(n62), .B(n170), .Z(n3) );
  XOR U115 ( .A(n4), .B(n169), .Z(n170) );
  XOR U116 ( .A(n171), .B(n27), .Z(n169) );
  AND U117 ( .A(n65), .B(n172), .Z(n27) );
  XNOR U118 ( .A(n173), .B(n28), .Z(n172) );
  XOR U119 ( .A(n174), .B(n175), .Z(n28) );
  AND U120 ( .A(n70), .B(n176), .Z(n175) );
  XOR U121 ( .A(p_input[8]), .B(n174), .Z(n176) );
  XOR U122 ( .A(n177), .B(n178), .Z(n174) );
  AND U123 ( .A(n74), .B(n179), .Z(n178) );
  IV U124 ( .A(n171), .Z(n173) );
  XOR U125 ( .A(n180), .B(n181), .Z(n171) );
  AND U126 ( .A(n78), .B(n182), .Z(n181) );
  XOR U127 ( .A(n183), .B(n184), .Z(n4) );
  AND U128 ( .A(n82), .B(n182), .Z(n184) );
  XNOR U129 ( .A(n185), .B(n180), .Z(n182) );
  XOR U130 ( .A(n186), .B(n187), .Z(n180) );
  AND U131 ( .A(n86), .B(n179), .Z(n187) );
  XNOR U132 ( .A(n188), .B(n177), .Z(n179) );
  XOR U133 ( .A(n189), .B(n190), .Z(n177) );
  AND U134 ( .A(n90), .B(n191), .Z(n190) );
  XOR U135 ( .A(p_input[24]), .B(n189), .Z(n191) );
  XOR U136 ( .A(n192), .B(n193), .Z(n189) );
  AND U137 ( .A(n94), .B(n194), .Z(n193) );
  IV U138 ( .A(n186), .Z(n188) );
  XOR U139 ( .A(n195), .B(n196), .Z(n186) );
  AND U140 ( .A(n98), .B(n197), .Z(n196) );
  IV U141 ( .A(n183), .Z(n185) );
  XNOR U142 ( .A(n198), .B(n199), .Z(n183) );
  AND U143 ( .A(n102), .B(n197), .Z(n199) );
  XNOR U144 ( .A(n198), .B(n195), .Z(n197) );
  XOR U145 ( .A(n200), .B(n201), .Z(n195) );
  AND U146 ( .A(n105), .B(n194), .Z(n201) );
  XNOR U147 ( .A(n202), .B(n192), .Z(n194) );
  XOR U148 ( .A(n203), .B(n204), .Z(n192) );
  AND U149 ( .A(n109), .B(n205), .Z(n204) );
  XOR U150 ( .A(p_input[40]), .B(n203), .Z(n205) );
  XOR U151 ( .A(n206), .B(n207), .Z(n203) );
  AND U152 ( .A(n113), .B(n208), .Z(n207) );
  IV U153 ( .A(n200), .Z(n202) );
  XOR U154 ( .A(n209), .B(n210), .Z(n200) );
  AND U155 ( .A(n117), .B(n211), .Z(n210) );
  XOR U156 ( .A(n212), .B(n213), .Z(n198) );
  AND U157 ( .A(n121), .B(n211), .Z(n213) );
  XNOR U158 ( .A(n212), .B(n209), .Z(n211) );
  XOR U159 ( .A(n214), .B(n215), .Z(n209) );
  AND U160 ( .A(n124), .B(n208), .Z(n215) );
  XNOR U161 ( .A(n216), .B(n206), .Z(n208) );
  XOR U162 ( .A(n217), .B(n218), .Z(n206) );
  AND U163 ( .A(n128), .B(n219), .Z(n218) );
  XOR U164 ( .A(p_input[56]), .B(n217), .Z(n219) );
  XOR U165 ( .A(n220), .B(n221), .Z(n217) );
  AND U166 ( .A(n132), .B(n222), .Z(n221) );
  IV U167 ( .A(n214), .Z(n216) );
  XOR U168 ( .A(n223), .B(n224), .Z(n214) );
  AND U169 ( .A(n136), .B(n225), .Z(n224) );
  XOR U170 ( .A(n226), .B(n227), .Z(n212) );
  AND U171 ( .A(n140), .B(n225), .Z(n227) );
  XNOR U172 ( .A(n226), .B(n223), .Z(n225) );
  XOR U173 ( .A(n228), .B(n229), .Z(n223) );
  AND U174 ( .A(n143), .B(n222), .Z(n229) );
  XNOR U175 ( .A(n230), .B(n220), .Z(n222) );
  XOR U176 ( .A(n231), .B(n232), .Z(n220) );
  AND U177 ( .A(n147), .B(n233), .Z(n232) );
  XOR U178 ( .A(p_input[72]), .B(n231), .Z(n233) );
  XOR U179 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n234), .Z(
        n231) );
  AND U180 ( .A(n150), .B(n235), .Z(n234) );
  IV U181 ( .A(n228), .Z(n230) );
  XOR U182 ( .A(n236), .B(n237), .Z(n228) );
  AND U183 ( .A(n154), .B(n238), .Z(n237) );
  XOR U184 ( .A(n239), .B(n240), .Z(n226) );
  AND U185 ( .A(n158), .B(n238), .Z(n240) );
  XNOR U186 ( .A(n239), .B(n236), .Z(n238) );
  XNOR U187 ( .A(n241), .B(n242), .Z(n236) );
  AND U188 ( .A(n161), .B(n235), .Z(n242) );
  XNOR U189 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n241), .Z(
        n235) );
  XNOR U190 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n243), .Z(
        n241) );
  AND U191 ( .A(n163), .B(n244), .Z(n243) );
  XNOR U192 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n245), .Z(n239) );
  AND U193 ( .A(n166), .B(n244), .Z(n245) );
  XOR U194 ( .A(n246), .B(n247), .Z(n244) );
  XOR U195 ( .A(n5), .B(n248), .Z(o[23]) );
  AND U196 ( .A(n62), .B(n249), .Z(n5) );
  XOR U197 ( .A(n6), .B(n248), .Z(n249) );
  XOR U198 ( .A(n250), .B(n31), .Z(n248) );
  AND U199 ( .A(n65), .B(n251), .Z(n31) );
  XNOR U200 ( .A(n252), .B(n32), .Z(n251) );
  XOR U201 ( .A(n253), .B(n254), .Z(n32) );
  AND U202 ( .A(n70), .B(n255), .Z(n254) );
  XOR U203 ( .A(p_input[7]), .B(n253), .Z(n255) );
  XOR U204 ( .A(n256), .B(n257), .Z(n253) );
  AND U205 ( .A(n74), .B(n258), .Z(n257) );
  IV U206 ( .A(n250), .Z(n252) );
  XOR U207 ( .A(n259), .B(n260), .Z(n250) );
  AND U208 ( .A(n78), .B(n261), .Z(n260) );
  XOR U209 ( .A(n262), .B(n263), .Z(n6) );
  AND U210 ( .A(n82), .B(n261), .Z(n263) );
  XNOR U211 ( .A(n264), .B(n259), .Z(n261) );
  XOR U212 ( .A(n265), .B(n266), .Z(n259) );
  AND U213 ( .A(n86), .B(n258), .Z(n266) );
  XNOR U214 ( .A(n267), .B(n256), .Z(n258) );
  XOR U215 ( .A(n268), .B(n269), .Z(n256) );
  AND U216 ( .A(n90), .B(n270), .Z(n269) );
  XOR U217 ( .A(p_input[23]), .B(n268), .Z(n270) );
  XOR U218 ( .A(n271), .B(n272), .Z(n268) );
  AND U219 ( .A(n94), .B(n273), .Z(n272) );
  IV U220 ( .A(n265), .Z(n267) );
  XOR U221 ( .A(n274), .B(n275), .Z(n265) );
  AND U222 ( .A(n98), .B(n276), .Z(n275) );
  IV U223 ( .A(n262), .Z(n264) );
  XNOR U224 ( .A(n277), .B(n278), .Z(n262) );
  AND U225 ( .A(n102), .B(n276), .Z(n278) );
  XNOR U226 ( .A(n277), .B(n274), .Z(n276) );
  XOR U227 ( .A(n279), .B(n280), .Z(n274) );
  AND U228 ( .A(n105), .B(n273), .Z(n280) );
  XNOR U229 ( .A(n281), .B(n271), .Z(n273) );
  XOR U230 ( .A(n282), .B(n283), .Z(n271) );
  AND U231 ( .A(n109), .B(n284), .Z(n283) );
  XOR U232 ( .A(p_input[39]), .B(n282), .Z(n284) );
  XOR U233 ( .A(n285), .B(n286), .Z(n282) );
  AND U234 ( .A(n113), .B(n287), .Z(n286) );
  IV U235 ( .A(n279), .Z(n281) );
  XOR U236 ( .A(n288), .B(n289), .Z(n279) );
  AND U237 ( .A(n117), .B(n290), .Z(n289) );
  XOR U238 ( .A(n291), .B(n292), .Z(n277) );
  AND U239 ( .A(n121), .B(n290), .Z(n292) );
  XNOR U240 ( .A(n291), .B(n288), .Z(n290) );
  XOR U241 ( .A(n293), .B(n294), .Z(n288) );
  AND U242 ( .A(n124), .B(n287), .Z(n294) );
  XNOR U243 ( .A(n295), .B(n285), .Z(n287) );
  XOR U244 ( .A(n296), .B(n297), .Z(n285) );
  AND U245 ( .A(n128), .B(n298), .Z(n297) );
  XOR U246 ( .A(p_input[55]), .B(n296), .Z(n298) );
  XOR U247 ( .A(n299), .B(n300), .Z(n296) );
  AND U248 ( .A(n132), .B(n301), .Z(n300) );
  IV U249 ( .A(n293), .Z(n295) );
  XOR U250 ( .A(n302), .B(n303), .Z(n293) );
  AND U251 ( .A(n136), .B(n304), .Z(n303) );
  XOR U252 ( .A(n305), .B(n306), .Z(n291) );
  AND U253 ( .A(n140), .B(n304), .Z(n306) );
  XNOR U254 ( .A(n305), .B(n302), .Z(n304) );
  XOR U255 ( .A(n307), .B(n308), .Z(n302) );
  AND U256 ( .A(n143), .B(n301), .Z(n308) );
  XNOR U257 ( .A(n309), .B(n299), .Z(n301) );
  XOR U258 ( .A(n310), .B(n311), .Z(n299) );
  AND U259 ( .A(n147), .B(n312), .Z(n311) );
  XOR U260 ( .A(p_input[71]), .B(n310), .Z(n312) );
  XOR U261 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n313), .Z(
        n310) );
  AND U262 ( .A(n150), .B(n314), .Z(n313) );
  IV U263 ( .A(n307), .Z(n309) );
  XOR U264 ( .A(n315), .B(n316), .Z(n307) );
  AND U265 ( .A(n154), .B(n317), .Z(n316) );
  XOR U266 ( .A(n318), .B(n319), .Z(n305) );
  AND U267 ( .A(n158), .B(n317), .Z(n319) );
  XNOR U268 ( .A(n318), .B(n315), .Z(n317) );
  XNOR U269 ( .A(n320), .B(n321), .Z(n315) );
  AND U270 ( .A(n161), .B(n314), .Z(n321) );
  XNOR U271 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n320), .Z(
        n314) );
  XNOR U272 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(n322), .Z(
        n320) );
  AND U273 ( .A(n163), .B(n323), .Z(n322) );
  XNOR U274 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n324), .Z(n318) );
  AND U275 ( .A(n166), .B(n323), .Z(n324) );
  XOR U276 ( .A(n325), .B(n326), .Z(n323) );
  IV U277 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n326) );
  IV U278 ( .A(\knn_comb_/min_val_out[0][7] ), .Z(n325) );
  XOR U279 ( .A(n7), .B(n327), .Z(o[22]) );
  AND U280 ( .A(n62), .B(n328), .Z(n7) );
  XOR U281 ( .A(n8), .B(n327), .Z(n328) );
  XOR U282 ( .A(n329), .B(n33), .Z(n327) );
  AND U283 ( .A(n65), .B(n330), .Z(n33) );
  XNOR U284 ( .A(n331), .B(n34), .Z(n330) );
  XOR U285 ( .A(n332), .B(n333), .Z(n34) );
  AND U286 ( .A(n70), .B(n334), .Z(n333) );
  XOR U287 ( .A(p_input[6]), .B(n332), .Z(n334) );
  XOR U288 ( .A(n335), .B(n336), .Z(n332) );
  AND U289 ( .A(n74), .B(n337), .Z(n336) );
  IV U290 ( .A(n329), .Z(n331) );
  XOR U291 ( .A(n338), .B(n339), .Z(n329) );
  AND U292 ( .A(n78), .B(n340), .Z(n339) );
  XOR U293 ( .A(n341), .B(n342), .Z(n8) );
  AND U294 ( .A(n82), .B(n340), .Z(n342) );
  XNOR U295 ( .A(n343), .B(n338), .Z(n340) );
  XOR U296 ( .A(n344), .B(n345), .Z(n338) );
  AND U297 ( .A(n86), .B(n337), .Z(n345) );
  XNOR U298 ( .A(n346), .B(n335), .Z(n337) );
  XOR U299 ( .A(n347), .B(n348), .Z(n335) );
  AND U300 ( .A(n90), .B(n349), .Z(n348) );
  XOR U301 ( .A(p_input[22]), .B(n347), .Z(n349) );
  XOR U302 ( .A(n350), .B(n351), .Z(n347) );
  AND U303 ( .A(n94), .B(n352), .Z(n351) );
  IV U304 ( .A(n344), .Z(n346) );
  XOR U305 ( .A(n353), .B(n354), .Z(n344) );
  AND U306 ( .A(n98), .B(n355), .Z(n354) );
  IV U307 ( .A(n341), .Z(n343) );
  XNOR U308 ( .A(n356), .B(n357), .Z(n341) );
  AND U309 ( .A(n102), .B(n355), .Z(n357) );
  XNOR U310 ( .A(n356), .B(n353), .Z(n355) );
  XOR U311 ( .A(n358), .B(n359), .Z(n353) );
  AND U312 ( .A(n105), .B(n352), .Z(n359) );
  XNOR U313 ( .A(n360), .B(n350), .Z(n352) );
  XOR U314 ( .A(n361), .B(n362), .Z(n350) );
  AND U315 ( .A(n109), .B(n363), .Z(n362) );
  XOR U316 ( .A(p_input[38]), .B(n361), .Z(n363) );
  XOR U317 ( .A(n364), .B(n365), .Z(n361) );
  AND U318 ( .A(n113), .B(n366), .Z(n365) );
  IV U319 ( .A(n358), .Z(n360) );
  XOR U320 ( .A(n367), .B(n368), .Z(n358) );
  AND U321 ( .A(n117), .B(n369), .Z(n368) );
  XOR U322 ( .A(n370), .B(n371), .Z(n356) );
  AND U323 ( .A(n121), .B(n369), .Z(n371) );
  XNOR U324 ( .A(n370), .B(n367), .Z(n369) );
  XOR U325 ( .A(n372), .B(n373), .Z(n367) );
  AND U326 ( .A(n124), .B(n366), .Z(n373) );
  XNOR U327 ( .A(n374), .B(n364), .Z(n366) );
  XOR U328 ( .A(n375), .B(n376), .Z(n364) );
  AND U329 ( .A(n128), .B(n377), .Z(n376) );
  XOR U330 ( .A(p_input[54]), .B(n375), .Z(n377) );
  XOR U331 ( .A(n378), .B(n379), .Z(n375) );
  AND U332 ( .A(n132), .B(n380), .Z(n379) );
  IV U333 ( .A(n372), .Z(n374) );
  XOR U334 ( .A(n381), .B(n382), .Z(n372) );
  AND U335 ( .A(n136), .B(n383), .Z(n382) );
  XOR U336 ( .A(n384), .B(n385), .Z(n370) );
  AND U337 ( .A(n140), .B(n383), .Z(n385) );
  XNOR U338 ( .A(n384), .B(n381), .Z(n383) );
  XOR U339 ( .A(n386), .B(n387), .Z(n381) );
  AND U340 ( .A(n143), .B(n380), .Z(n387) );
  XNOR U341 ( .A(n388), .B(n378), .Z(n380) );
  XOR U342 ( .A(n389), .B(n390), .Z(n378) );
  AND U343 ( .A(n147), .B(n391), .Z(n390) );
  XOR U344 ( .A(p_input[70]), .B(n389), .Z(n391) );
  XOR U345 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n392), .Z(
        n389) );
  AND U346 ( .A(n150), .B(n393), .Z(n392) );
  IV U347 ( .A(n386), .Z(n388) );
  XOR U348 ( .A(n394), .B(n395), .Z(n386) );
  AND U349 ( .A(n154), .B(n396), .Z(n395) );
  XOR U350 ( .A(n397), .B(n398), .Z(n384) );
  AND U351 ( .A(n158), .B(n396), .Z(n398) );
  XNOR U352 ( .A(n397), .B(n394), .Z(n396) );
  XNOR U353 ( .A(n399), .B(n400), .Z(n394) );
  AND U354 ( .A(n161), .B(n393), .Z(n400) );
  XNOR U355 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n399), .Z(
        n393) );
  XNOR U356 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(n401), .Z(
        n399) );
  AND U357 ( .A(n163), .B(n402), .Z(n401) );
  XNOR U358 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n403), .Z(n397) );
  AND U359 ( .A(n166), .B(n402), .Z(n403) );
  XOR U360 ( .A(n404), .B(n405), .Z(n402) );
  XOR U361 ( .A(n9), .B(n406), .Z(o[21]) );
  AND U362 ( .A(n62), .B(n407), .Z(n9) );
  XOR U363 ( .A(n10), .B(n406), .Z(n407) );
  XOR U364 ( .A(n408), .B(n35), .Z(n406) );
  AND U365 ( .A(n65), .B(n409), .Z(n35) );
  XNOR U366 ( .A(n410), .B(n36), .Z(n409) );
  XOR U367 ( .A(n411), .B(n412), .Z(n36) );
  AND U368 ( .A(n70), .B(n413), .Z(n412) );
  XOR U369 ( .A(p_input[5]), .B(n411), .Z(n413) );
  XOR U370 ( .A(n414), .B(n415), .Z(n411) );
  AND U371 ( .A(n74), .B(n416), .Z(n415) );
  IV U372 ( .A(n408), .Z(n410) );
  XOR U373 ( .A(n417), .B(n418), .Z(n408) );
  AND U374 ( .A(n78), .B(n419), .Z(n418) );
  XOR U375 ( .A(n420), .B(n421), .Z(n10) );
  AND U376 ( .A(n82), .B(n419), .Z(n421) );
  XNOR U377 ( .A(n422), .B(n417), .Z(n419) );
  XOR U378 ( .A(n423), .B(n424), .Z(n417) );
  AND U379 ( .A(n86), .B(n416), .Z(n424) );
  XNOR U380 ( .A(n425), .B(n414), .Z(n416) );
  XOR U381 ( .A(n426), .B(n427), .Z(n414) );
  AND U382 ( .A(n90), .B(n428), .Z(n427) );
  XOR U383 ( .A(p_input[21]), .B(n426), .Z(n428) );
  XOR U384 ( .A(n429), .B(n430), .Z(n426) );
  AND U385 ( .A(n94), .B(n431), .Z(n430) );
  IV U386 ( .A(n423), .Z(n425) );
  XOR U387 ( .A(n432), .B(n433), .Z(n423) );
  AND U388 ( .A(n98), .B(n434), .Z(n433) );
  IV U389 ( .A(n420), .Z(n422) );
  XNOR U390 ( .A(n435), .B(n436), .Z(n420) );
  AND U391 ( .A(n102), .B(n434), .Z(n436) );
  XNOR U392 ( .A(n435), .B(n432), .Z(n434) );
  XOR U393 ( .A(n437), .B(n438), .Z(n432) );
  AND U394 ( .A(n105), .B(n431), .Z(n438) );
  XNOR U395 ( .A(n439), .B(n429), .Z(n431) );
  XOR U396 ( .A(n440), .B(n441), .Z(n429) );
  AND U397 ( .A(n109), .B(n442), .Z(n441) );
  XOR U398 ( .A(p_input[37]), .B(n440), .Z(n442) );
  XOR U399 ( .A(n443), .B(n444), .Z(n440) );
  AND U400 ( .A(n113), .B(n445), .Z(n444) );
  IV U401 ( .A(n437), .Z(n439) );
  XOR U402 ( .A(n446), .B(n447), .Z(n437) );
  AND U403 ( .A(n117), .B(n448), .Z(n447) );
  XOR U404 ( .A(n449), .B(n450), .Z(n435) );
  AND U405 ( .A(n121), .B(n448), .Z(n450) );
  XNOR U406 ( .A(n449), .B(n446), .Z(n448) );
  XOR U407 ( .A(n451), .B(n452), .Z(n446) );
  AND U408 ( .A(n124), .B(n445), .Z(n452) );
  XNOR U409 ( .A(n453), .B(n443), .Z(n445) );
  XOR U410 ( .A(n454), .B(n455), .Z(n443) );
  AND U411 ( .A(n128), .B(n456), .Z(n455) );
  XOR U412 ( .A(p_input[53]), .B(n454), .Z(n456) );
  XOR U413 ( .A(n457), .B(n458), .Z(n454) );
  AND U414 ( .A(n132), .B(n459), .Z(n458) );
  IV U415 ( .A(n451), .Z(n453) );
  XOR U416 ( .A(n460), .B(n461), .Z(n451) );
  AND U417 ( .A(n136), .B(n462), .Z(n461) );
  XOR U418 ( .A(n463), .B(n464), .Z(n449) );
  AND U419 ( .A(n140), .B(n462), .Z(n464) );
  XNOR U420 ( .A(n463), .B(n460), .Z(n462) );
  XOR U421 ( .A(n465), .B(n466), .Z(n460) );
  AND U422 ( .A(n143), .B(n459), .Z(n466) );
  XNOR U423 ( .A(n467), .B(n457), .Z(n459) );
  XOR U424 ( .A(n468), .B(n469), .Z(n457) );
  AND U425 ( .A(n147), .B(n470), .Z(n469) );
  XOR U426 ( .A(p_input[69]), .B(n468), .Z(n470) );
  XOR U427 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n471), .Z(
        n468) );
  AND U428 ( .A(n150), .B(n472), .Z(n471) );
  IV U429 ( .A(n465), .Z(n467) );
  XOR U430 ( .A(n473), .B(n474), .Z(n465) );
  AND U431 ( .A(n154), .B(n475), .Z(n474) );
  XOR U432 ( .A(n476), .B(n477), .Z(n463) );
  AND U433 ( .A(n158), .B(n475), .Z(n477) );
  XNOR U434 ( .A(n476), .B(n473), .Z(n475) );
  XNOR U435 ( .A(n478), .B(n479), .Z(n473) );
  AND U436 ( .A(n161), .B(n472), .Z(n479) );
  XNOR U437 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n478), .Z(
        n472) );
  XNOR U438 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n480), .Z(
        n478) );
  AND U439 ( .A(n163), .B(n481), .Z(n480) );
  XNOR U440 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n482), .Z(n476) );
  AND U441 ( .A(n166), .B(n481), .Z(n482) );
  XOR U442 ( .A(n483), .B(n484), .Z(n481) );
  XOR U443 ( .A(n11), .B(n485), .Z(o[20]) );
  AND U444 ( .A(n62), .B(n486), .Z(n11) );
  XOR U445 ( .A(n12), .B(n485), .Z(n486) );
  XOR U446 ( .A(n487), .B(n37), .Z(n485) );
  AND U447 ( .A(n65), .B(n488), .Z(n37) );
  XNOR U448 ( .A(n489), .B(n38), .Z(n488) );
  XOR U449 ( .A(n490), .B(n491), .Z(n38) );
  AND U450 ( .A(n70), .B(n492), .Z(n491) );
  XOR U451 ( .A(p_input[4]), .B(n490), .Z(n492) );
  XOR U452 ( .A(n493), .B(n494), .Z(n490) );
  AND U453 ( .A(n74), .B(n495), .Z(n494) );
  IV U454 ( .A(n487), .Z(n489) );
  XOR U455 ( .A(n496), .B(n497), .Z(n487) );
  AND U456 ( .A(n78), .B(n498), .Z(n497) );
  XOR U457 ( .A(n499), .B(n500), .Z(n12) );
  AND U458 ( .A(n82), .B(n498), .Z(n500) );
  XNOR U459 ( .A(n501), .B(n496), .Z(n498) );
  XOR U460 ( .A(n502), .B(n503), .Z(n496) );
  AND U461 ( .A(n86), .B(n495), .Z(n503) );
  XNOR U462 ( .A(n504), .B(n493), .Z(n495) );
  XOR U463 ( .A(n505), .B(n506), .Z(n493) );
  AND U464 ( .A(n90), .B(n507), .Z(n506) );
  XOR U465 ( .A(p_input[20]), .B(n505), .Z(n507) );
  XOR U466 ( .A(n508), .B(n509), .Z(n505) );
  AND U467 ( .A(n94), .B(n510), .Z(n509) );
  IV U468 ( .A(n502), .Z(n504) );
  XOR U469 ( .A(n511), .B(n512), .Z(n502) );
  AND U470 ( .A(n98), .B(n513), .Z(n512) );
  IV U471 ( .A(n499), .Z(n501) );
  XNOR U472 ( .A(n514), .B(n515), .Z(n499) );
  AND U473 ( .A(n102), .B(n513), .Z(n515) );
  XNOR U474 ( .A(n514), .B(n511), .Z(n513) );
  XOR U475 ( .A(n516), .B(n517), .Z(n511) );
  AND U476 ( .A(n105), .B(n510), .Z(n517) );
  XNOR U477 ( .A(n518), .B(n508), .Z(n510) );
  XOR U478 ( .A(n519), .B(n520), .Z(n508) );
  AND U479 ( .A(n109), .B(n521), .Z(n520) );
  XOR U480 ( .A(p_input[36]), .B(n519), .Z(n521) );
  XOR U481 ( .A(n522), .B(n523), .Z(n519) );
  AND U482 ( .A(n113), .B(n524), .Z(n523) );
  IV U483 ( .A(n516), .Z(n518) );
  XOR U484 ( .A(n525), .B(n526), .Z(n516) );
  AND U485 ( .A(n117), .B(n527), .Z(n526) );
  XOR U486 ( .A(n528), .B(n529), .Z(n514) );
  AND U487 ( .A(n121), .B(n527), .Z(n529) );
  XNOR U488 ( .A(n528), .B(n525), .Z(n527) );
  XOR U489 ( .A(n530), .B(n531), .Z(n525) );
  AND U490 ( .A(n124), .B(n524), .Z(n531) );
  XNOR U491 ( .A(n532), .B(n522), .Z(n524) );
  XOR U492 ( .A(n533), .B(n534), .Z(n522) );
  AND U493 ( .A(n128), .B(n535), .Z(n534) );
  XOR U494 ( .A(p_input[52]), .B(n533), .Z(n535) );
  XOR U495 ( .A(n536), .B(n537), .Z(n533) );
  AND U496 ( .A(n132), .B(n538), .Z(n537) );
  IV U497 ( .A(n530), .Z(n532) );
  XOR U498 ( .A(n539), .B(n540), .Z(n530) );
  AND U499 ( .A(n136), .B(n541), .Z(n540) );
  XOR U500 ( .A(n542), .B(n543), .Z(n528) );
  AND U501 ( .A(n140), .B(n541), .Z(n543) );
  XNOR U502 ( .A(n542), .B(n539), .Z(n541) );
  XOR U503 ( .A(n544), .B(n545), .Z(n539) );
  AND U504 ( .A(n143), .B(n538), .Z(n545) );
  XNOR U505 ( .A(n546), .B(n536), .Z(n538) );
  XOR U506 ( .A(n547), .B(n548), .Z(n536) );
  AND U507 ( .A(n147), .B(n549), .Z(n548) );
  XOR U508 ( .A(p_input[68]), .B(n547), .Z(n549) );
  XOR U509 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n550), .Z(
        n547) );
  AND U510 ( .A(n150), .B(n551), .Z(n550) );
  IV U511 ( .A(n544), .Z(n546) );
  XOR U512 ( .A(n552), .B(n553), .Z(n544) );
  AND U513 ( .A(n154), .B(n554), .Z(n553) );
  XOR U514 ( .A(n555), .B(n556), .Z(n542) );
  AND U515 ( .A(n158), .B(n554), .Z(n556) );
  XNOR U516 ( .A(n555), .B(n552), .Z(n554) );
  XNOR U517 ( .A(n557), .B(n558), .Z(n552) );
  AND U518 ( .A(n161), .B(n551), .Z(n558) );
  XNOR U519 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n557), .Z(
        n551) );
  XNOR U520 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n559), .Z(
        n557) );
  AND U521 ( .A(n163), .B(n560), .Z(n559) );
  XNOR U522 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n561), .Z(n555) );
  AND U523 ( .A(n166), .B(n560), .Z(n561) );
  XOR U524 ( .A(n562), .B(n563), .Z(n560) );
  IV U525 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n563) );
  IV U526 ( .A(\knn_comb_/min_val_out[0][4] ), .Z(n562) );
  XOR U527 ( .A(n564), .B(n565), .Z(o[1]) );
  XOR U528 ( .A(n29), .B(n566), .Z(o[19]) );
  AND U529 ( .A(n62), .B(n567), .Z(n29) );
  XOR U530 ( .A(n30), .B(n566), .Z(n567) );
  XOR U531 ( .A(n568), .B(n39), .Z(n566) );
  AND U532 ( .A(n65), .B(n569), .Z(n39) );
  XNOR U533 ( .A(n570), .B(n40), .Z(n569) );
  XOR U534 ( .A(n571), .B(n572), .Z(n40) );
  AND U535 ( .A(n70), .B(n573), .Z(n572) );
  XOR U536 ( .A(p_input[3]), .B(n571), .Z(n573) );
  XOR U537 ( .A(n574), .B(n575), .Z(n571) );
  AND U538 ( .A(n74), .B(n576), .Z(n575) );
  IV U539 ( .A(n568), .Z(n570) );
  XOR U540 ( .A(n577), .B(n578), .Z(n568) );
  AND U541 ( .A(n78), .B(n579), .Z(n578) );
  XOR U542 ( .A(n580), .B(n581), .Z(n30) );
  AND U543 ( .A(n82), .B(n579), .Z(n581) );
  XNOR U544 ( .A(n582), .B(n577), .Z(n579) );
  XOR U545 ( .A(n583), .B(n584), .Z(n577) );
  AND U546 ( .A(n86), .B(n576), .Z(n584) );
  XNOR U547 ( .A(n585), .B(n574), .Z(n576) );
  XOR U548 ( .A(n586), .B(n587), .Z(n574) );
  AND U549 ( .A(n90), .B(n588), .Z(n587) );
  XOR U550 ( .A(p_input[19]), .B(n586), .Z(n588) );
  XOR U551 ( .A(n589), .B(n590), .Z(n586) );
  AND U552 ( .A(n94), .B(n591), .Z(n590) );
  IV U553 ( .A(n583), .Z(n585) );
  XOR U554 ( .A(n592), .B(n593), .Z(n583) );
  AND U555 ( .A(n98), .B(n594), .Z(n593) );
  IV U556 ( .A(n580), .Z(n582) );
  XNOR U557 ( .A(n595), .B(n596), .Z(n580) );
  AND U558 ( .A(n102), .B(n594), .Z(n596) );
  XNOR U559 ( .A(n595), .B(n592), .Z(n594) );
  XOR U560 ( .A(n597), .B(n598), .Z(n592) );
  AND U561 ( .A(n105), .B(n591), .Z(n598) );
  XNOR U562 ( .A(n599), .B(n589), .Z(n591) );
  XOR U563 ( .A(n600), .B(n601), .Z(n589) );
  AND U564 ( .A(n109), .B(n602), .Z(n601) );
  XOR U565 ( .A(p_input[35]), .B(n600), .Z(n602) );
  XOR U566 ( .A(n603), .B(n604), .Z(n600) );
  AND U567 ( .A(n113), .B(n605), .Z(n604) );
  IV U568 ( .A(n597), .Z(n599) );
  XOR U569 ( .A(n606), .B(n607), .Z(n597) );
  AND U570 ( .A(n117), .B(n608), .Z(n607) );
  XOR U571 ( .A(n609), .B(n610), .Z(n595) );
  AND U572 ( .A(n121), .B(n608), .Z(n610) );
  XNOR U573 ( .A(n609), .B(n606), .Z(n608) );
  XOR U574 ( .A(n611), .B(n612), .Z(n606) );
  AND U575 ( .A(n124), .B(n605), .Z(n612) );
  XNOR U576 ( .A(n613), .B(n603), .Z(n605) );
  XOR U577 ( .A(n614), .B(n615), .Z(n603) );
  AND U578 ( .A(n128), .B(n616), .Z(n615) );
  XOR U579 ( .A(p_input[51]), .B(n614), .Z(n616) );
  XOR U580 ( .A(n617), .B(n618), .Z(n614) );
  AND U581 ( .A(n132), .B(n619), .Z(n618) );
  IV U582 ( .A(n611), .Z(n613) );
  XOR U583 ( .A(n620), .B(n621), .Z(n611) );
  AND U584 ( .A(n136), .B(n622), .Z(n621) );
  XOR U585 ( .A(n623), .B(n624), .Z(n609) );
  AND U586 ( .A(n140), .B(n622), .Z(n624) );
  XNOR U587 ( .A(n623), .B(n620), .Z(n622) );
  XOR U588 ( .A(n625), .B(n626), .Z(n620) );
  AND U589 ( .A(n143), .B(n619), .Z(n626) );
  XNOR U590 ( .A(n627), .B(n617), .Z(n619) );
  XOR U591 ( .A(n628), .B(n629), .Z(n617) );
  AND U592 ( .A(n147), .B(n630), .Z(n629) );
  XOR U593 ( .A(p_input[67]), .B(n628), .Z(n630) );
  XOR U594 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n631), .Z(
        n628) );
  AND U595 ( .A(n150), .B(n632), .Z(n631) );
  IV U596 ( .A(n625), .Z(n627) );
  XOR U597 ( .A(n633), .B(n634), .Z(n625) );
  AND U598 ( .A(n154), .B(n635), .Z(n634) );
  XOR U599 ( .A(n636), .B(n637), .Z(n623) );
  AND U600 ( .A(n158), .B(n635), .Z(n637) );
  XNOR U601 ( .A(n636), .B(n633), .Z(n635) );
  XNOR U602 ( .A(n638), .B(n639), .Z(n633) );
  AND U603 ( .A(n161), .B(n632), .Z(n639) );
  XNOR U604 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n638), .Z(
        n632) );
  XNOR U605 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(n640), .Z(
        n638) );
  AND U606 ( .A(n163), .B(n641), .Z(n640) );
  XNOR U607 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n642), .Z(n636) );
  AND U608 ( .A(n166), .B(n641), .Z(n642) );
  XOR U609 ( .A(n643), .B(n644), .Z(n641) );
  XOR U610 ( .A(n51), .B(n645), .Z(o[18]) );
  AND U611 ( .A(n62), .B(n646), .Z(n51) );
  XOR U612 ( .A(n52), .B(n645), .Z(n646) );
  XOR U613 ( .A(n647), .B(n41), .Z(n645) );
  AND U614 ( .A(n65), .B(n648), .Z(n41) );
  XOR U615 ( .A(n42), .B(n647), .Z(n648) );
  XOR U616 ( .A(n649), .B(n650), .Z(n42) );
  AND U617 ( .A(n70), .B(n651), .Z(n650) );
  XOR U618 ( .A(p_input[2]), .B(n649), .Z(n651) );
  XNOR U619 ( .A(n652), .B(n653), .Z(n649) );
  AND U620 ( .A(n74), .B(n654), .Z(n653) );
  XOR U621 ( .A(n655), .B(n656), .Z(n647) );
  AND U622 ( .A(n78), .B(n657), .Z(n656) );
  XOR U623 ( .A(n658), .B(n659), .Z(n52) );
  AND U624 ( .A(n82), .B(n657), .Z(n659) );
  XNOR U625 ( .A(n660), .B(n658), .Z(n657) );
  IV U626 ( .A(n655), .Z(n660) );
  XOR U627 ( .A(n661), .B(n662), .Z(n655) );
  AND U628 ( .A(n86), .B(n654), .Z(n662) );
  XNOR U629 ( .A(n652), .B(n661), .Z(n654) );
  XNOR U630 ( .A(n663), .B(n664), .Z(n652) );
  AND U631 ( .A(n90), .B(n665), .Z(n664) );
  XOR U632 ( .A(p_input[18]), .B(n663), .Z(n665) );
  XNOR U633 ( .A(n666), .B(n667), .Z(n663) );
  AND U634 ( .A(n94), .B(n668), .Z(n667) );
  XOR U635 ( .A(n669), .B(n670), .Z(n661) );
  AND U636 ( .A(n98), .B(n671), .Z(n670) );
  XOR U637 ( .A(n672), .B(n673), .Z(n658) );
  AND U638 ( .A(n102), .B(n671), .Z(n673) );
  XNOR U639 ( .A(n674), .B(n672), .Z(n671) );
  IV U640 ( .A(n669), .Z(n674) );
  XOR U641 ( .A(n675), .B(n676), .Z(n669) );
  AND U642 ( .A(n105), .B(n668), .Z(n676) );
  XNOR U643 ( .A(n666), .B(n675), .Z(n668) );
  XNOR U644 ( .A(n677), .B(n678), .Z(n666) );
  AND U645 ( .A(n109), .B(n679), .Z(n678) );
  XOR U646 ( .A(p_input[34]), .B(n677), .Z(n679) );
  XNOR U647 ( .A(n680), .B(n681), .Z(n677) );
  AND U648 ( .A(n113), .B(n682), .Z(n681) );
  XOR U649 ( .A(n683), .B(n684), .Z(n675) );
  AND U650 ( .A(n117), .B(n685), .Z(n684) );
  XOR U651 ( .A(n686), .B(n687), .Z(n672) );
  AND U652 ( .A(n121), .B(n685), .Z(n687) );
  XNOR U653 ( .A(n688), .B(n686), .Z(n685) );
  IV U654 ( .A(n683), .Z(n688) );
  XOR U655 ( .A(n689), .B(n690), .Z(n683) );
  AND U656 ( .A(n124), .B(n682), .Z(n690) );
  XNOR U657 ( .A(n680), .B(n689), .Z(n682) );
  XNOR U658 ( .A(n691), .B(n692), .Z(n680) );
  AND U659 ( .A(n128), .B(n693), .Z(n692) );
  XOR U660 ( .A(p_input[50]), .B(n691), .Z(n693) );
  XNOR U661 ( .A(n694), .B(n695), .Z(n691) );
  AND U662 ( .A(n132), .B(n696), .Z(n695) );
  XOR U663 ( .A(n697), .B(n698), .Z(n689) );
  AND U664 ( .A(n136), .B(n699), .Z(n698) );
  XOR U665 ( .A(n700), .B(n701), .Z(n686) );
  AND U666 ( .A(n140), .B(n699), .Z(n701) );
  XNOR U667 ( .A(n702), .B(n700), .Z(n699) );
  IV U668 ( .A(n697), .Z(n702) );
  XOR U669 ( .A(n703), .B(n704), .Z(n697) );
  AND U670 ( .A(n143), .B(n696), .Z(n704) );
  XNOR U671 ( .A(n694), .B(n703), .Z(n696) );
  XNOR U672 ( .A(n705), .B(n706), .Z(n694) );
  AND U673 ( .A(n147), .B(n707), .Z(n706) );
  XOR U674 ( .A(p_input[66]), .B(n705), .Z(n707) );
  XOR U675 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n708), .Z(
        n705) );
  AND U676 ( .A(n150), .B(n709), .Z(n708) );
  XOR U677 ( .A(n710), .B(n711), .Z(n703) );
  AND U678 ( .A(n154), .B(n712), .Z(n711) );
  XOR U679 ( .A(n713), .B(n714), .Z(n700) );
  AND U680 ( .A(n158), .B(n712), .Z(n714) );
  XNOR U681 ( .A(n715), .B(n713), .Z(n712) );
  IV U682 ( .A(n710), .Z(n715) );
  XOR U683 ( .A(n716), .B(n717), .Z(n710) );
  AND U684 ( .A(n161), .B(n709), .Z(n717) );
  XOR U685 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n716), .Z(
        n709) );
  XOR U686 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(n718), .Z(
        n716) );
  AND U687 ( .A(n163), .B(n719), .Z(n718) );
  XOR U688 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n720), .Z(n713) );
  AND U689 ( .A(n166), .B(n719), .Z(n720) );
  XOR U690 ( .A(\knn_comb_/min_val_out[0][2] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n719) );
  XOR U691 ( .A(n564), .B(n721), .Z(o[17]) );
  AND U692 ( .A(n62), .B(n722), .Z(n564) );
  XOR U693 ( .A(n565), .B(n721), .Z(n722) );
  XOR U694 ( .A(n723), .B(n43), .Z(n721) );
  AND U695 ( .A(n65), .B(n724), .Z(n43) );
  XOR U696 ( .A(n44), .B(n723), .Z(n724) );
  XOR U697 ( .A(n725), .B(n726), .Z(n44) );
  AND U698 ( .A(n70), .B(n727), .Z(n726) );
  XOR U699 ( .A(p_input[1]), .B(n725), .Z(n727) );
  XNOR U700 ( .A(n728), .B(n729), .Z(n725) );
  AND U701 ( .A(n74), .B(n730), .Z(n729) );
  XOR U702 ( .A(n731), .B(n732), .Z(n723) );
  AND U703 ( .A(n78), .B(n733), .Z(n732) );
  XOR U704 ( .A(n734), .B(n735), .Z(n565) );
  AND U705 ( .A(n82), .B(n733), .Z(n735) );
  XNOR U706 ( .A(n736), .B(n734), .Z(n733) );
  IV U707 ( .A(n731), .Z(n736) );
  XOR U708 ( .A(n737), .B(n738), .Z(n731) );
  AND U709 ( .A(n86), .B(n730), .Z(n738) );
  XNOR U710 ( .A(n728), .B(n737), .Z(n730) );
  XNOR U711 ( .A(n739), .B(n740), .Z(n728) );
  AND U712 ( .A(n90), .B(n741), .Z(n740) );
  XOR U713 ( .A(p_input[17]), .B(n739), .Z(n741) );
  XNOR U714 ( .A(n742), .B(n743), .Z(n739) );
  AND U715 ( .A(n94), .B(n744), .Z(n743) );
  XOR U716 ( .A(n745), .B(n746), .Z(n737) );
  AND U717 ( .A(n98), .B(n747), .Z(n746) );
  XOR U718 ( .A(n748), .B(n749), .Z(n734) );
  AND U719 ( .A(n102), .B(n747), .Z(n749) );
  XNOR U720 ( .A(n750), .B(n748), .Z(n747) );
  IV U721 ( .A(n745), .Z(n750) );
  XOR U722 ( .A(n751), .B(n752), .Z(n745) );
  AND U723 ( .A(n105), .B(n744), .Z(n752) );
  XNOR U724 ( .A(n742), .B(n751), .Z(n744) );
  XNOR U725 ( .A(n753), .B(n754), .Z(n742) );
  AND U726 ( .A(n109), .B(n755), .Z(n754) );
  XOR U727 ( .A(p_input[33]), .B(n753), .Z(n755) );
  XNOR U728 ( .A(n756), .B(n757), .Z(n753) );
  AND U729 ( .A(n113), .B(n758), .Z(n757) );
  XOR U730 ( .A(n759), .B(n760), .Z(n751) );
  AND U731 ( .A(n117), .B(n761), .Z(n760) );
  XOR U732 ( .A(n762), .B(n763), .Z(n748) );
  AND U733 ( .A(n121), .B(n761), .Z(n763) );
  XNOR U734 ( .A(n764), .B(n762), .Z(n761) );
  IV U735 ( .A(n759), .Z(n764) );
  XOR U736 ( .A(n765), .B(n766), .Z(n759) );
  AND U737 ( .A(n124), .B(n758), .Z(n766) );
  XNOR U738 ( .A(n756), .B(n765), .Z(n758) );
  XNOR U739 ( .A(n767), .B(n768), .Z(n756) );
  AND U740 ( .A(n128), .B(n769), .Z(n768) );
  XOR U741 ( .A(p_input[49]), .B(n767), .Z(n769) );
  XNOR U742 ( .A(n770), .B(n771), .Z(n767) );
  AND U743 ( .A(n132), .B(n772), .Z(n771) );
  XOR U744 ( .A(n773), .B(n774), .Z(n765) );
  AND U745 ( .A(n136), .B(n775), .Z(n774) );
  XOR U746 ( .A(n776), .B(n777), .Z(n762) );
  AND U747 ( .A(n140), .B(n775), .Z(n777) );
  XNOR U748 ( .A(n778), .B(n776), .Z(n775) );
  IV U749 ( .A(n773), .Z(n778) );
  XOR U750 ( .A(n779), .B(n780), .Z(n773) );
  AND U751 ( .A(n143), .B(n772), .Z(n780) );
  XNOR U752 ( .A(n770), .B(n779), .Z(n772) );
  XNOR U753 ( .A(n781), .B(n782), .Z(n770) );
  AND U754 ( .A(n147), .B(n783), .Z(n782) );
  XOR U755 ( .A(p_input[65]), .B(n781), .Z(n783) );
  XOR U756 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n784), .Z(
        n781) );
  AND U757 ( .A(n150), .B(n785), .Z(n784) );
  XOR U758 ( .A(n786), .B(n787), .Z(n779) );
  AND U759 ( .A(n154), .B(n788), .Z(n787) );
  XOR U760 ( .A(n789), .B(n790), .Z(n776) );
  AND U761 ( .A(n158), .B(n788), .Z(n790) );
  XNOR U762 ( .A(n791), .B(n789), .Z(n788) );
  IV U763 ( .A(n786), .Z(n791) );
  XOR U764 ( .A(n792), .B(n793), .Z(n786) );
  AND U765 ( .A(n161), .B(n785), .Z(n793) );
  XOR U766 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n792), .Z(
        n785) );
  XOR U767 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(n794), .Z(
        n792) );
  AND U768 ( .A(n163), .B(n795), .Z(n794) );
  XOR U769 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n796), .Z(n789) );
  AND U770 ( .A(n166), .B(n795), .Z(n796) );
  XOR U771 ( .A(\knn_comb_/min_val_out[0][1] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n795) );
  XOR U772 ( .A(n797), .B(n798), .Z(o[16]) );
  XOR U773 ( .A(n47), .B(n799), .Z(o[15]) );
  AND U774 ( .A(n62), .B(n800), .Z(n47) );
  XOR U775 ( .A(n48), .B(n799), .Z(n800) );
  XOR U776 ( .A(n801), .B(n802), .Z(n799) );
  AND U777 ( .A(n82), .B(n803), .Z(n802) );
  XOR U778 ( .A(n804), .B(n13), .Z(n48) );
  AND U779 ( .A(n65), .B(n805), .Z(n13) );
  XOR U780 ( .A(n14), .B(n804), .Z(n805) );
  XOR U781 ( .A(n806), .B(n807), .Z(n14) );
  AND U782 ( .A(n70), .B(n808), .Z(n807) );
  XOR U783 ( .A(p_input[15]), .B(n806), .Z(n808) );
  XNOR U784 ( .A(n809), .B(n810), .Z(n806) );
  AND U785 ( .A(n74), .B(n811), .Z(n810) );
  XOR U786 ( .A(n812), .B(n813), .Z(n804) );
  AND U787 ( .A(n78), .B(n803), .Z(n813) );
  XNOR U788 ( .A(n814), .B(n801), .Z(n803) );
  XOR U789 ( .A(n815), .B(n816), .Z(n801) );
  AND U790 ( .A(n102), .B(n817), .Z(n816) );
  IV U791 ( .A(n812), .Z(n814) );
  XOR U792 ( .A(n818), .B(n819), .Z(n812) );
  AND U793 ( .A(n86), .B(n811), .Z(n819) );
  XNOR U794 ( .A(n809), .B(n818), .Z(n811) );
  XNOR U795 ( .A(n820), .B(n821), .Z(n809) );
  AND U796 ( .A(n90), .B(n822), .Z(n821) );
  XOR U797 ( .A(p_input[31]), .B(n820), .Z(n822) );
  XNOR U798 ( .A(n823), .B(n824), .Z(n820) );
  AND U799 ( .A(n94), .B(n825), .Z(n824) );
  XOR U800 ( .A(n826), .B(n827), .Z(n818) );
  AND U801 ( .A(n98), .B(n817), .Z(n827) );
  XNOR U802 ( .A(n828), .B(n815), .Z(n817) );
  XOR U803 ( .A(n829), .B(n830), .Z(n815) );
  AND U804 ( .A(n121), .B(n831), .Z(n830) );
  IV U805 ( .A(n826), .Z(n828) );
  XOR U806 ( .A(n832), .B(n833), .Z(n826) );
  AND U807 ( .A(n105), .B(n825), .Z(n833) );
  XNOR U808 ( .A(n823), .B(n832), .Z(n825) );
  XNOR U809 ( .A(n834), .B(n835), .Z(n823) );
  AND U810 ( .A(n109), .B(n836), .Z(n835) );
  XOR U811 ( .A(p_input[47]), .B(n834), .Z(n836) );
  XNOR U812 ( .A(n837), .B(n838), .Z(n834) );
  AND U813 ( .A(n113), .B(n839), .Z(n838) );
  XOR U814 ( .A(n840), .B(n841), .Z(n832) );
  AND U815 ( .A(n117), .B(n831), .Z(n841) );
  XNOR U816 ( .A(n842), .B(n829), .Z(n831) );
  XOR U817 ( .A(n843), .B(n844), .Z(n829) );
  AND U818 ( .A(n140), .B(n845), .Z(n844) );
  IV U819 ( .A(n840), .Z(n842) );
  XOR U820 ( .A(n846), .B(n847), .Z(n840) );
  AND U821 ( .A(n124), .B(n839), .Z(n847) );
  XNOR U822 ( .A(n837), .B(n846), .Z(n839) );
  XNOR U823 ( .A(n848), .B(n849), .Z(n837) );
  AND U824 ( .A(n128), .B(n850), .Z(n849) );
  XOR U825 ( .A(p_input[63]), .B(n848), .Z(n850) );
  XNOR U826 ( .A(n851), .B(n852), .Z(n848) );
  AND U827 ( .A(n132), .B(n853), .Z(n852) );
  XOR U828 ( .A(n854), .B(n855), .Z(n846) );
  AND U829 ( .A(n136), .B(n845), .Z(n855) );
  XNOR U830 ( .A(n856), .B(n843), .Z(n845) );
  XOR U831 ( .A(n857), .B(n858), .Z(n843) );
  AND U832 ( .A(n158), .B(n859), .Z(n858) );
  IV U833 ( .A(n854), .Z(n856) );
  XOR U834 ( .A(n860), .B(n861), .Z(n854) );
  AND U835 ( .A(n143), .B(n853), .Z(n861) );
  XNOR U836 ( .A(n851), .B(n860), .Z(n853) );
  XNOR U837 ( .A(n862), .B(n863), .Z(n851) );
  AND U838 ( .A(n147), .B(n864), .Z(n863) );
  XOR U839 ( .A(p_input[79]), .B(n862), .Z(n864) );
  XOR U840 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n865), .Z(
        n862) );
  AND U841 ( .A(n150), .B(n866), .Z(n865) );
  XOR U842 ( .A(n867), .B(n868), .Z(n860) );
  AND U843 ( .A(n154), .B(n859), .Z(n868) );
  XNOR U844 ( .A(n869), .B(n857), .Z(n859) );
  XOR U845 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n870), .Z(n857) );
  AND U846 ( .A(n166), .B(n871), .Z(n870) );
  IV U847 ( .A(n867), .Z(n869) );
  XOR U848 ( .A(n872), .B(n873), .Z(n867) );
  AND U849 ( .A(n161), .B(n866), .Z(n873) );
  XOR U850 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n872), .Z(
        n866) );
  XOR U851 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n874), .Z(
        n872) );
  AND U852 ( .A(n163), .B(n871), .Z(n874) );
  XOR U853 ( .A(n875), .B(n876), .Z(n871) );
  IV U854 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n876) );
  IV U855 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n875) );
  XOR U856 ( .A(n49), .B(n877), .Z(o[14]) );
  AND U857 ( .A(n62), .B(n878), .Z(n49) );
  XOR U858 ( .A(n50), .B(n877), .Z(n878) );
  XOR U859 ( .A(n879), .B(n880), .Z(n877) );
  AND U860 ( .A(n82), .B(n881), .Z(n880) );
  XOR U861 ( .A(n882), .B(n15), .Z(n50) );
  AND U862 ( .A(n65), .B(n883), .Z(n15) );
  XOR U863 ( .A(n16), .B(n882), .Z(n883) );
  XOR U864 ( .A(n884), .B(n885), .Z(n16) );
  AND U865 ( .A(n70), .B(n886), .Z(n885) );
  XOR U866 ( .A(p_input[14]), .B(n884), .Z(n886) );
  XNOR U867 ( .A(n887), .B(n888), .Z(n884) );
  AND U868 ( .A(n74), .B(n889), .Z(n888) );
  XOR U869 ( .A(n890), .B(n891), .Z(n882) );
  AND U870 ( .A(n78), .B(n881), .Z(n891) );
  XNOR U871 ( .A(n892), .B(n879), .Z(n881) );
  XOR U872 ( .A(n893), .B(n894), .Z(n879) );
  AND U873 ( .A(n102), .B(n895), .Z(n894) );
  IV U874 ( .A(n890), .Z(n892) );
  XOR U875 ( .A(n896), .B(n897), .Z(n890) );
  AND U876 ( .A(n86), .B(n889), .Z(n897) );
  XNOR U877 ( .A(n887), .B(n896), .Z(n889) );
  XNOR U878 ( .A(n898), .B(n899), .Z(n887) );
  AND U879 ( .A(n90), .B(n900), .Z(n899) );
  XOR U880 ( .A(p_input[30]), .B(n898), .Z(n900) );
  XNOR U881 ( .A(n901), .B(n902), .Z(n898) );
  AND U882 ( .A(n94), .B(n903), .Z(n902) );
  XOR U883 ( .A(n904), .B(n905), .Z(n896) );
  AND U884 ( .A(n98), .B(n895), .Z(n905) );
  XNOR U885 ( .A(n906), .B(n893), .Z(n895) );
  XOR U886 ( .A(n907), .B(n908), .Z(n893) );
  AND U887 ( .A(n121), .B(n909), .Z(n908) );
  IV U888 ( .A(n904), .Z(n906) );
  XOR U889 ( .A(n910), .B(n911), .Z(n904) );
  AND U890 ( .A(n105), .B(n903), .Z(n911) );
  XNOR U891 ( .A(n901), .B(n910), .Z(n903) );
  XNOR U892 ( .A(n912), .B(n913), .Z(n901) );
  AND U893 ( .A(n109), .B(n914), .Z(n913) );
  XOR U894 ( .A(p_input[46]), .B(n912), .Z(n914) );
  XNOR U895 ( .A(n915), .B(n916), .Z(n912) );
  AND U896 ( .A(n113), .B(n917), .Z(n916) );
  XOR U897 ( .A(n918), .B(n919), .Z(n910) );
  AND U898 ( .A(n117), .B(n909), .Z(n919) );
  XNOR U899 ( .A(n920), .B(n907), .Z(n909) );
  XOR U900 ( .A(n921), .B(n922), .Z(n907) );
  AND U901 ( .A(n140), .B(n923), .Z(n922) );
  IV U902 ( .A(n918), .Z(n920) );
  XOR U903 ( .A(n924), .B(n925), .Z(n918) );
  AND U904 ( .A(n124), .B(n917), .Z(n925) );
  XNOR U905 ( .A(n915), .B(n924), .Z(n917) );
  XNOR U906 ( .A(n926), .B(n927), .Z(n915) );
  AND U907 ( .A(n128), .B(n928), .Z(n927) );
  XOR U908 ( .A(p_input[62]), .B(n926), .Z(n928) );
  XNOR U909 ( .A(n929), .B(n930), .Z(n926) );
  AND U910 ( .A(n132), .B(n931), .Z(n930) );
  XOR U911 ( .A(n932), .B(n933), .Z(n924) );
  AND U912 ( .A(n136), .B(n923), .Z(n933) );
  XNOR U913 ( .A(n934), .B(n921), .Z(n923) );
  XOR U914 ( .A(n935), .B(n936), .Z(n921) );
  AND U915 ( .A(n158), .B(n937), .Z(n936) );
  IV U916 ( .A(n932), .Z(n934) );
  XOR U917 ( .A(n938), .B(n939), .Z(n932) );
  AND U918 ( .A(n143), .B(n931), .Z(n939) );
  XNOR U919 ( .A(n929), .B(n938), .Z(n931) );
  XNOR U920 ( .A(n940), .B(n941), .Z(n929) );
  AND U921 ( .A(n147), .B(n942), .Z(n941) );
  XOR U922 ( .A(p_input[78]), .B(n940), .Z(n942) );
  XOR U923 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n943), .Z(
        n940) );
  AND U924 ( .A(n150), .B(n944), .Z(n943) );
  XOR U925 ( .A(n945), .B(n946), .Z(n938) );
  AND U926 ( .A(n154), .B(n937), .Z(n946) );
  XNOR U927 ( .A(n947), .B(n935), .Z(n937) );
  XOR U928 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n948), .Z(n935) );
  AND U929 ( .A(n166), .B(n949), .Z(n948) );
  IV U930 ( .A(n945), .Z(n947) );
  XOR U931 ( .A(n950), .B(n951), .Z(n945) );
  AND U932 ( .A(n161), .B(n944), .Z(n951) );
  XOR U933 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n950), .Z(
        n944) );
  XOR U934 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n952), .Z(
        n950) );
  AND U935 ( .A(n163), .B(n949), .Z(n952) );
  XOR U936 ( .A(n953), .B(n954), .Z(n949) );
  IV U937 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n954) );
  IV U938 ( .A(\knn_comb_/min_val_out[0][14] ), .Z(n953) );
  XOR U939 ( .A(n53), .B(n955), .Z(o[13]) );
  AND U940 ( .A(n62), .B(n956), .Z(n53) );
  XOR U941 ( .A(n54), .B(n955), .Z(n956) );
  XOR U942 ( .A(n957), .B(n958), .Z(n955) );
  AND U943 ( .A(n82), .B(n959), .Z(n958) );
  XOR U944 ( .A(n960), .B(n17), .Z(n54) );
  AND U945 ( .A(n65), .B(n961), .Z(n17) );
  XOR U946 ( .A(n18), .B(n960), .Z(n961) );
  XOR U947 ( .A(n962), .B(n963), .Z(n18) );
  AND U948 ( .A(n70), .B(n964), .Z(n963) );
  XOR U949 ( .A(p_input[13]), .B(n962), .Z(n964) );
  XNOR U950 ( .A(n965), .B(n966), .Z(n962) );
  AND U951 ( .A(n74), .B(n967), .Z(n966) );
  XOR U952 ( .A(n968), .B(n969), .Z(n960) );
  AND U953 ( .A(n78), .B(n959), .Z(n969) );
  XNOR U954 ( .A(n970), .B(n957), .Z(n959) );
  XOR U955 ( .A(n971), .B(n972), .Z(n957) );
  AND U956 ( .A(n102), .B(n973), .Z(n972) );
  IV U957 ( .A(n968), .Z(n970) );
  XOR U958 ( .A(n974), .B(n975), .Z(n968) );
  AND U959 ( .A(n86), .B(n967), .Z(n975) );
  XNOR U960 ( .A(n965), .B(n974), .Z(n967) );
  XNOR U961 ( .A(n976), .B(n977), .Z(n965) );
  AND U962 ( .A(n90), .B(n978), .Z(n977) );
  XOR U963 ( .A(p_input[29]), .B(n976), .Z(n978) );
  XNOR U964 ( .A(n979), .B(n980), .Z(n976) );
  AND U965 ( .A(n94), .B(n981), .Z(n980) );
  XOR U966 ( .A(n982), .B(n983), .Z(n974) );
  AND U967 ( .A(n98), .B(n973), .Z(n983) );
  XNOR U968 ( .A(n984), .B(n971), .Z(n973) );
  XOR U969 ( .A(n985), .B(n986), .Z(n971) );
  AND U970 ( .A(n121), .B(n987), .Z(n986) );
  IV U971 ( .A(n982), .Z(n984) );
  XOR U972 ( .A(n988), .B(n989), .Z(n982) );
  AND U973 ( .A(n105), .B(n981), .Z(n989) );
  XNOR U974 ( .A(n979), .B(n988), .Z(n981) );
  XNOR U975 ( .A(n990), .B(n991), .Z(n979) );
  AND U976 ( .A(n109), .B(n992), .Z(n991) );
  XOR U977 ( .A(p_input[45]), .B(n990), .Z(n992) );
  XNOR U978 ( .A(n993), .B(n994), .Z(n990) );
  AND U979 ( .A(n113), .B(n995), .Z(n994) );
  XOR U980 ( .A(n996), .B(n997), .Z(n988) );
  AND U981 ( .A(n117), .B(n987), .Z(n997) );
  XNOR U982 ( .A(n998), .B(n985), .Z(n987) );
  XOR U983 ( .A(n999), .B(n1000), .Z(n985) );
  AND U984 ( .A(n140), .B(n1001), .Z(n1000) );
  IV U985 ( .A(n996), .Z(n998) );
  XOR U986 ( .A(n1002), .B(n1003), .Z(n996) );
  AND U987 ( .A(n124), .B(n995), .Z(n1003) );
  XNOR U988 ( .A(n993), .B(n1002), .Z(n995) );
  XNOR U989 ( .A(n1004), .B(n1005), .Z(n993) );
  AND U990 ( .A(n128), .B(n1006), .Z(n1005) );
  XOR U991 ( .A(p_input[61]), .B(n1004), .Z(n1006) );
  XNOR U992 ( .A(n1007), .B(n1008), .Z(n1004) );
  AND U993 ( .A(n132), .B(n1009), .Z(n1008) );
  XOR U994 ( .A(n1010), .B(n1011), .Z(n1002) );
  AND U995 ( .A(n136), .B(n1001), .Z(n1011) );
  XNOR U996 ( .A(n1012), .B(n999), .Z(n1001) );
  XOR U997 ( .A(n1013), .B(n1014), .Z(n999) );
  AND U998 ( .A(n158), .B(n1015), .Z(n1014) );
  IV U999 ( .A(n1010), .Z(n1012) );
  XOR U1000 ( .A(n1016), .B(n1017), .Z(n1010) );
  AND U1001 ( .A(n143), .B(n1009), .Z(n1017) );
  XNOR U1002 ( .A(n1007), .B(n1016), .Z(n1009) );
  XNOR U1003 ( .A(n1018), .B(n1019), .Z(n1007) );
  AND U1004 ( .A(n147), .B(n1020), .Z(n1019) );
  XOR U1005 ( .A(p_input[77]), .B(n1018), .Z(n1020) );
  XOR U1006 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n1021), 
        .Z(n1018) );
  AND U1007 ( .A(n150), .B(n1022), .Z(n1021) );
  XOR U1008 ( .A(n1023), .B(n1024), .Z(n1016) );
  AND U1009 ( .A(n154), .B(n1015), .Z(n1024) );
  XNOR U1010 ( .A(n1025), .B(n1013), .Z(n1015) );
  XOR U1011 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n1026), .Z(n1013) );
  AND U1012 ( .A(n166), .B(n1027), .Z(n1026) );
  IV U1013 ( .A(n1023), .Z(n1025) );
  XOR U1014 ( .A(n1028), .B(n1029), .Z(n1023) );
  AND U1015 ( .A(n161), .B(n1022), .Z(n1029) );
  XOR U1016 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n1028), 
        .Z(n1022) );
  XOR U1017 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(n1030), 
        .Z(n1028) );
  AND U1018 ( .A(n163), .B(n1027), .Z(n1030) );
  XOR U1019 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n1027) );
  XOR U1020 ( .A(n55), .B(n1031), .Z(o[12]) );
  AND U1021 ( .A(n62), .B(n1032), .Z(n55) );
  XOR U1022 ( .A(n56), .B(n1031), .Z(n1032) );
  XOR U1023 ( .A(n1033), .B(n1034), .Z(n1031) );
  AND U1024 ( .A(n82), .B(n1035), .Z(n1034) );
  XOR U1025 ( .A(n1036), .B(n19), .Z(n56) );
  AND U1026 ( .A(n65), .B(n1037), .Z(n19) );
  XOR U1027 ( .A(n20), .B(n1036), .Z(n1037) );
  XOR U1028 ( .A(n1038), .B(n1039), .Z(n20) );
  AND U1029 ( .A(n70), .B(n1040), .Z(n1039) );
  XOR U1030 ( .A(p_input[12]), .B(n1038), .Z(n1040) );
  XNOR U1031 ( .A(n1041), .B(n1042), .Z(n1038) );
  AND U1032 ( .A(n74), .B(n1043), .Z(n1042) );
  XOR U1033 ( .A(n1044), .B(n1045), .Z(n1036) );
  AND U1034 ( .A(n78), .B(n1035), .Z(n1045) );
  XNOR U1035 ( .A(n1046), .B(n1033), .Z(n1035) );
  XOR U1036 ( .A(n1047), .B(n1048), .Z(n1033) );
  AND U1037 ( .A(n102), .B(n1049), .Z(n1048) );
  IV U1038 ( .A(n1044), .Z(n1046) );
  XOR U1039 ( .A(n1050), .B(n1051), .Z(n1044) );
  AND U1040 ( .A(n86), .B(n1043), .Z(n1051) );
  XNOR U1041 ( .A(n1041), .B(n1050), .Z(n1043) );
  XNOR U1042 ( .A(n1052), .B(n1053), .Z(n1041) );
  AND U1043 ( .A(n90), .B(n1054), .Z(n1053) );
  XOR U1044 ( .A(p_input[28]), .B(n1052), .Z(n1054) );
  XNOR U1045 ( .A(n1055), .B(n1056), .Z(n1052) );
  AND U1046 ( .A(n94), .B(n1057), .Z(n1056) );
  XOR U1047 ( .A(n1058), .B(n1059), .Z(n1050) );
  AND U1048 ( .A(n98), .B(n1049), .Z(n1059) );
  XNOR U1049 ( .A(n1060), .B(n1047), .Z(n1049) );
  XOR U1050 ( .A(n1061), .B(n1062), .Z(n1047) );
  AND U1051 ( .A(n121), .B(n1063), .Z(n1062) );
  IV U1052 ( .A(n1058), .Z(n1060) );
  XOR U1053 ( .A(n1064), .B(n1065), .Z(n1058) );
  AND U1054 ( .A(n105), .B(n1057), .Z(n1065) );
  XNOR U1055 ( .A(n1055), .B(n1064), .Z(n1057) );
  XNOR U1056 ( .A(n1066), .B(n1067), .Z(n1055) );
  AND U1057 ( .A(n109), .B(n1068), .Z(n1067) );
  XOR U1058 ( .A(p_input[44]), .B(n1066), .Z(n1068) );
  XNOR U1059 ( .A(n1069), .B(n1070), .Z(n1066) );
  AND U1060 ( .A(n113), .B(n1071), .Z(n1070) );
  XOR U1061 ( .A(n1072), .B(n1073), .Z(n1064) );
  AND U1062 ( .A(n117), .B(n1063), .Z(n1073) );
  XNOR U1063 ( .A(n1074), .B(n1061), .Z(n1063) );
  XOR U1064 ( .A(n1075), .B(n1076), .Z(n1061) );
  AND U1065 ( .A(n140), .B(n1077), .Z(n1076) );
  IV U1066 ( .A(n1072), .Z(n1074) );
  XOR U1067 ( .A(n1078), .B(n1079), .Z(n1072) );
  AND U1068 ( .A(n124), .B(n1071), .Z(n1079) );
  XNOR U1069 ( .A(n1069), .B(n1078), .Z(n1071) );
  XNOR U1070 ( .A(n1080), .B(n1081), .Z(n1069) );
  AND U1071 ( .A(n128), .B(n1082), .Z(n1081) );
  XOR U1072 ( .A(p_input[60]), .B(n1080), .Z(n1082) );
  XNOR U1073 ( .A(n1083), .B(n1084), .Z(n1080) );
  AND U1074 ( .A(n132), .B(n1085), .Z(n1084) );
  XOR U1075 ( .A(n1086), .B(n1087), .Z(n1078) );
  AND U1076 ( .A(n136), .B(n1077), .Z(n1087) );
  XNOR U1077 ( .A(n1088), .B(n1075), .Z(n1077) );
  XOR U1078 ( .A(n1089), .B(n1090), .Z(n1075) );
  AND U1079 ( .A(n158), .B(n1091), .Z(n1090) );
  IV U1080 ( .A(n1086), .Z(n1088) );
  XOR U1081 ( .A(n1092), .B(n1093), .Z(n1086) );
  AND U1082 ( .A(n143), .B(n1085), .Z(n1093) );
  XNOR U1083 ( .A(n1083), .B(n1092), .Z(n1085) );
  XNOR U1084 ( .A(n1094), .B(n1095), .Z(n1083) );
  AND U1085 ( .A(n147), .B(n1096), .Z(n1095) );
  XOR U1086 ( .A(p_input[76]), .B(n1094), .Z(n1096) );
  XOR U1087 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n1097), 
        .Z(n1094) );
  AND U1088 ( .A(n150), .B(n1098), .Z(n1097) );
  XOR U1089 ( .A(n1099), .B(n1100), .Z(n1092) );
  AND U1090 ( .A(n154), .B(n1091), .Z(n1100) );
  XNOR U1091 ( .A(n1101), .B(n1089), .Z(n1091) );
  XOR U1092 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n1102), .Z(n1089) );
  AND U1093 ( .A(n166), .B(n1103), .Z(n1102) );
  IV U1094 ( .A(n1099), .Z(n1101) );
  XOR U1095 ( .A(n1104), .B(n1105), .Z(n1099) );
  AND U1096 ( .A(n161), .B(n1098), .Z(n1105) );
  XOR U1097 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n1104), 
        .Z(n1098) );
  XOR U1098 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n1106), 
        .Z(n1104) );
  AND U1099 ( .A(n163), .B(n1103), .Z(n1106) );
  XOR U1100 ( .A(\knn_comb_/min_val_out[0][12] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n1103) );
  XOR U1101 ( .A(n57), .B(n1107), .Z(o[11]) );
  AND U1102 ( .A(n62), .B(n1108), .Z(n57) );
  XOR U1103 ( .A(n58), .B(n1107), .Z(n1108) );
  XOR U1104 ( .A(n1109), .B(n1110), .Z(n1107) );
  AND U1105 ( .A(n82), .B(n1111), .Z(n1110) );
  XOR U1106 ( .A(n1112), .B(n21), .Z(n58) );
  AND U1107 ( .A(n65), .B(n1113), .Z(n21) );
  XOR U1108 ( .A(n22), .B(n1112), .Z(n1113) );
  XOR U1109 ( .A(n1114), .B(n1115), .Z(n22) );
  AND U1110 ( .A(n70), .B(n1116), .Z(n1115) );
  XOR U1111 ( .A(p_input[11]), .B(n1114), .Z(n1116) );
  XNOR U1112 ( .A(n1117), .B(n1118), .Z(n1114) );
  AND U1113 ( .A(n74), .B(n1119), .Z(n1118) );
  XOR U1114 ( .A(n1120), .B(n1121), .Z(n1112) );
  AND U1115 ( .A(n78), .B(n1111), .Z(n1121) );
  XNOR U1116 ( .A(n1122), .B(n1109), .Z(n1111) );
  XOR U1117 ( .A(n1123), .B(n1124), .Z(n1109) );
  AND U1118 ( .A(n102), .B(n1125), .Z(n1124) );
  IV U1119 ( .A(n1120), .Z(n1122) );
  XOR U1120 ( .A(n1126), .B(n1127), .Z(n1120) );
  AND U1121 ( .A(n86), .B(n1119), .Z(n1127) );
  XNOR U1122 ( .A(n1117), .B(n1126), .Z(n1119) );
  XNOR U1123 ( .A(n1128), .B(n1129), .Z(n1117) );
  AND U1124 ( .A(n90), .B(n1130), .Z(n1129) );
  XOR U1125 ( .A(p_input[27]), .B(n1128), .Z(n1130) );
  XNOR U1126 ( .A(n1131), .B(n1132), .Z(n1128) );
  AND U1127 ( .A(n94), .B(n1133), .Z(n1132) );
  XOR U1128 ( .A(n1134), .B(n1135), .Z(n1126) );
  AND U1129 ( .A(n98), .B(n1125), .Z(n1135) );
  XNOR U1130 ( .A(n1136), .B(n1123), .Z(n1125) );
  XOR U1131 ( .A(n1137), .B(n1138), .Z(n1123) );
  AND U1132 ( .A(n121), .B(n1139), .Z(n1138) );
  IV U1133 ( .A(n1134), .Z(n1136) );
  XOR U1134 ( .A(n1140), .B(n1141), .Z(n1134) );
  AND U1135 ( .A(n105), .B(n1133), .Z(n1141) );
  XNOR U1136 ( .A(n1131), .B(n1140), .Z(n1133) );
  XNOR U1137 ( .A(n1142), .B(n1143), .Z(n1131) );
  AND U1138 ( .A(n109), .B(n1144), .Z(n1143) );
  XOR U1139 ( .A(p_input[43]), .B(n1142), .Z(n1144) );
  XNOR U1140 ( .A(n1145), .B(n1146), .Z(n1142) );
  AND U1141 ( .A(n113), .B(n1147), .Z(n1146) );
  XOR U1142 ( .A(n1148), .B(n1149), .Z(n1140) );
  AND U1143 ( .A(n117), .B(n1139), .Z(n1149) );
  XNOR U1144 ( .A(n1150), .B(n1137), .Z(n1139) );
  XOR U1145 ( .A(n1151), .B(n1152), .Z(n1137) );
  AND U1146 ( .A(n140), .B(n1153), .Z(n1152) );
  IV U1147 ( .A(n1148), .Z(n1150) );
  XOR U1148 ( .A(n1154), .B(n1155), .Z(n1148) );
  AND U1149 ( .A(n124), .B(n1147), .Z(n1155) );
  XNOR U1150 ( .A(n1145), .B(n1154), .Z(n1147) );
  XNOR U1151 ( .A(n1156), .B(n1157), .Z(n1145) );
  AND U1152 ( .A(n128), .B(n1158), .Z(n1157) );
  XOR U1153 ( .A(p_input[59]), .B(n1156), .Z(n1158) );
  XNOR U1154 ( .A(n1159), .B(n1160), .Z(n1156) );
  AND U1155 ( .A(n132), .B(n1161), .Z(n1160) );
  XOR U1156 ( .A(n1162), .B(n1163), .Z(n1154) );
  AND U1157 ( .A(n136), .B(n1153), .Z(n1163) );
  XNOR U1158 ( .A(n1164), .B(n1151), .Z(n1153) );
  XOR U1159 ( .A(n1165), .B(n1166), .Z(n1151) );
  AND U1160 ( .A(n158), .B(n1167), .Z(n1166) );
  IV U1161 ( .A(n1162), .Z(n1164) );
  XOR U1162 ( .A(n1168), .B(n1169), .Z(n1162) );
  AND U1163 ( .A(n143), .B(n1161), .Z(n1169) );
  XNOR U1164 ( .A(n1159), .B(n1168), .Z(n1161) );
  XNOR U1165 ( .A(n1170), .B(n1171), .Z(n1159) );
  AND U1166 ( .A(n147), .B(n1172), .Z(n1171) );
  XOR U1167 ( .A(p_input[75]), .B(n1170), .Z(n1172) );
  XOR U1168 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n1173), 
        .Z(n1170) );
  AND U1169 ( .A(n150), .B(n1174), .Z(n1173) );
  XOR U1170 ( .A(n1175), .B(n1176), .Z(n1168) );
  AND U1171 ( .A(n154), .B(n1167), .Z(n1176) );
  XNOR U1172 ( .A(n1177), .B(n1165), .Z(n1167) );
  XOR U1173 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n1178), .Z(n1165) );
  AND U1174 ( .A(n166), .B(n1179), .Z(n1178) );
  IV U1175 ( .A(n1175), .Z(n1177) );
  XOR U1176 ( .A(n1180), .B(n1181), .Z(n1175) );
  AND U1177 ( .A(n161), .B(n1174), .Z(n1181) );
  XOR U1178 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n1180), 
        .Z(n1174) );
  XOR U1179 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n1182), 
        .Z(n1180) );
  AND U1180 ( .A(n163), .B(n1179), .Z(n1182) );
  XOR U1181 ( .A(n1183), .B(n1184), .Z(n1179) );
  IV U1182 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n1184) );
  IV U1183 ( .A(\knn_comb_/min_val_out[0][11] ), .Z(n1183) );
  XOR U1184 ( .A(n59), .B(n1185), .Z(o[10]) );
  AND U1185 ( .A(n62), .B(n1186), .Z(n59) );
  XOR U1186 ( .A(n60), .B(n1185), .Z(n1186) );
  XOR U1187 ( .A(n1187), .B(n1188), .Z(n1185) );
  AND U1188 ( .A(n82), .B(n1189), .Z(n1188) );
  XOR U1189 ( .A(n1190), .B(n23), .Z(n60) );
  AND U1190 ( .A(n65), .B(n1191), .Z(n23) );
  XOR U1191 ( .A(n24), .B(n1190), .Z(n1191) );
  XOR U1192 ( .A(n1192), .B(n1193), .Z(n24) );
  AND U1193 ( .A(n70), .B(n1194), .Z(n1193) );
  XOR U1194 ( .A(p_input[10]), .B(n1192), .Z(n1194) );
  XNOR U1195 ( .A(n1195), .B(n1196), .Z(n1192) );
  AND U1196 ( .A(n74), .B(n1197), .Z(n1196) );
  XOR U1197 ( .A(n1198), .B(n1199), .Z(n1190) );
  AND U1198 ( .A(n78), .B(n1189), .Z(n1199) );
  XNOR U1199 ( .A(n1200), .B(n1187), .Z(n1189) );
  XOR U1200 ( .A(n1201), .B(n1202), .Z(n1187) );
  AND U1201 ( .A(n102), .B(n1203), .Z(n1202) );
  IV U1202 ( .A(n1198), .Z(n1200) );
  XOR U1203 ( .A(n1204), .B(n1205), .Z(n1198) );
  AND U1204 ( .A(n86), .B(n1197), .Z(n1205) );
  XNOR U1205 ( .A(n1195), .B(n1204), .Z(n1197) );
  XNOR U1206 ( .A(n1206), .B(n1207), .Z(n1195) );
  AND U1207 ( .A(n90), .B(n1208), .Z(n1207) );
  XOR U1208 ( .A(p_input[26]), .B(n1206), .Z(n1208) );
  XNOR U1209 ( .A(n1209), .B(n1210), .Z(n1206) );
  AND U1210 ( .A(n94), .B(n1211), .Z(n1210) );
  XOR U1211 ( .A(n1212), .B(n1213), .Z(n1204) );
  AND U1212 ( .A(n98), .B(n1203), .Z(n1213) );
  XNOR U1213 ( .A(n1214), .B(n1201), .Z(n1203) );
  XOR U1214 ( .A(n1215), .B(n1216), .Z(n1201) );
  AND U1215 ( .A(n121), .B(n1217), .Z(n1216) );
  IV U1216 ( .A(n1212), .Z(n1214) );
  XOR U1217 ( .A(n1218), .B(n1219), .Z(n1212) );
  AND U1218 ( .A(n105), .B(n1211), .Z(n1219) );
  XNOR U1219 ( .A(n1209), .B(n1218), .Z(n1211) );
  XNOR U1220 ( .A(n1220), .B(n1221), .Z(n1209) );
  AND U1221 ( .A(n109), .B(n1222), .Z(n1221) );
  XOR U1222 ( .A(p_input[42]), .B(n1220), .Z(n1222) );
  XNOR U1223 ( .A(n1223), .B(n1224), .Z(n1220) );
  AND U1224 ( .A(n113), .B(n1225), .Z(n1224) );
  XOR U1225 ( .A(n1226), .B(n1227), .Z(n1218) );
  AND U1226 ( .A(n117), .B(n1217), .Z(n1227) );
  XNOR U1227 ( .A(n1228), .B(n1215), .Z(n1217) );
  XOR U1228 ( .A(n1229), .B(n1230), .Z(n1215) );
  AND U1229 ( .A(n140), .B(n1231), .Z(n1230) );
  IV U1230 ( .A(n1226), .Z(n1228) );
  XOR U1231 ( .A(n1232), .B(n1233), .Z(n1226) );
  AND U1232 ( .A(n124), .B(n1225), .Z(n1233) );
  XNOR U1233 ( .A(n1223), .B(n1232), .Z(n1225) );
  XNOR U1234 ( .A(n1234), .B(n1235), .Z(n1223) );
  AND U1235 ( .A(n128), .B(n1236), .Z(n1235) );
  XOR U1236 ( .A(p_input[58]), .B(n1234), .Z(n1236) );
  XNOR U1237 ( .A(n1237), .B(n1238), .Z(n1234) );
  AND U1238 ( .A(n132), .B(n1239), .Z(n1238) );
  XOR U1239 ( .A(n1240), .B(n1241), .Z(n1232) );
  AND U1240 ( .A(n136), .B(n1231), .Z(n1241) );
  XNOR U1241 ( .A(n1242), .B(n1229), .Z(n1231) );
  XOR U1242 ( .A(n1243), .B(n1244), .Z(n1229) );
  AND U1243 ( .A(n158), .B(n1245), .Z(n1244) );
  IV U1244 ( .A(n1240), .Z(n1242) );
  XOR U1245 ( .A(n1246), .B(n1247), .Z(n1240) );
  AND U1246 ( .A(n143), .B(n1239), .Z(n1247) );
  XNOR U1247 ( .A(n1237), .B(n1246), .Z(n1239) );
  XNOR U1248 ( .A(n1248), .B(n1249), .Z(n1237) );
  AND U1249 ( .A(n147), .B(n1250), .Z(n1249) );
  XOR U1250 ( .A(p_input[74]), .B(n1248), .Z(n1250) );
  XOR U1251 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n1251), 
        .Z(n1248) );
  AND U1252 ( .A(n150), .B(n1252), .Z(n1251) );
  XOR U1253 ( .A(n1253), .B(n1254), .Z(n1246) );
  AND U1254 ( .A(n154), .B(n1245), .Z(n1254) );
  XNOR U1255 ( .A(n1255), .B(n1243), .Z(n1245) );
  XOR U1256 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n1256), .Z(n1243) );
  AND U1257 ( .A(n166), .B(n1257), .Z(n1256) );
  IV U1258 ( .A(n1253), .Z(n1255) );
  XOR U1259 ( .A(n1258), .B(n1259), .Z(n1253) );
  AND U1260 ( .A(n161), .B(n1252), .Z(n1259) );
  XOR U1261 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n1258), 
        .Z(n1252) );
  XOR U1262 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(n1260), 
        .Z(n1258) );
  AND U1263 ( .A(n163), .B(n1257), .Z(n1260) );
  XOR U1264 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n1257) );
  XOR U1265 ( .A(n797), .B(n1261), .Z(o[0]) );
  AND U1266 ( .A(n62), .B(n1262), .Z(n797) );
  XOR U1267 ( .A(n798), .B(n1261), .Z(n1262) );
  XOR U1268 ( .A(n1263), .B(n1264), .Z(n1261) );
  AND U1269 ( .A(n82), .B(n1265), .Z(n1264) );
  XOR U1270 ( .A(n1266), .B(n45), .Z(n798) );
  AND U1271 ( .A(n65), .B(n1267), .Z(n45) );
  XOR U1272 ( .A(n46), .B(n1266), .Z(n1267) );
  XOR U1273 ( .A(n1268), .B(n1269), .Z(n46) );
  AND U1274 ( .A(n70), .B(n1270), .Z(n1269) );
  XOR U1275 ( .A(p_input[0]), .B(n1268), .Z(n1270) );
  XNOR U1276 ( .A(n1271), .B(n1272), .Z(n1268) );
  AND U1277 ( .A(n74), .B(n1273), .Z(n1272) );
  XOR U1278 ( .A(n1274), .B(n1275), .Z(n1266) );
  AND U1279 ( .A(n78), .B(n1265), .Z(n1275) );
  XNOR U1280 ( .A(n1276), .B(n1263), .Z(n1265) );
  XOR U1281 ( .A(n1277), .B(n1278), .Z(n1263) );
  AND U1282 ( .A(n102), .B(n1279), .Z(n1278) );
  IV U1283 ( .A(n1274), .Z(n1276) );
  XOR U1284 ( .A(n1280), .B(n1281), .Z(n1274) );
  AND U1285 ( .A(n86), .B(n1273), .Z(n1281) );
  XNOR U1286 ( .A(n1271), .B(n1280), .Z(n1273) );
  XNOR U1287 ( .A(n1282), .B(n1283), .Z(n1271) );
  AND U1288 ( .A(n90), .B(n1284), .Z(n1283) );
  XOR U1289 ( .A(p_input[16]), .B(n1282), .Z(n1284) );
  XNOR U1290 ( .A(n1285), .B(n1286), .Z(n1282) );
  AND U1291 ( .A(n94), .B(n1287), .Z(n1286) );
  XOR U1292 ( .A(n1288), .B(n1289), .Z(n1280) );
  AND U1293 ( .A(n98), .B(n1279), .Z(n1289) );
  XNOR U1294 ( .A(n1290), .B(n1277), .Z(n1279) );
  XOR U1295 ( .A(n1291), .B(n1292), .Z(n1277) );
  AND U1296 ( .A(n121), .B(n1293), .Z(n1292) );
  IV U1297 ( .A(n1288), .Z(n1290) );
  XOR U1298 ( .A(n1294), .B(n1295), .Z(n1288) );
  AND U1299 ( .A(n105), .B(n1287), .Z(n1295) );
  XNOR U1300 ( .A(n1285), .B(n1294), .Z(n1287) );
  XNOR U1301 ( .A(n1296), .B(n1297), .Z(n1285) );
  AND U1302 ( .A(n109), .B(n1298), .Z(n1297) );
  XOR U1303 ( .A(p_input[32]), .B(n1296), .Z(n1298) );
  XNOR U1304 ( .A(n1299), .B(n1300), .Z(n1296) );
  AND U1305 ( .A(n113), .B(n1301), .Z(n1300) );
  XOR U1306 ( .A(n1302), .B(n1303), .Z(n1294) );
  AND U1307 ( .A(n117), .B(n1293), .Z(n1303) );
  XNOR U1308 ( .A(n1304), .B(n1291), .Z(n1293) );
  XOR U1309 ( .A(n1305), .B(n1306), .Z(n1291) );
  AND U1310 ( .A(n140), .B(n1307), .Z(n1306) );
  IV U1311 ( .A(n1302), .Z(n1304) );
  XOR U1312 ( .A(n1308), .B(n1309), .Z(n1302) );
  AND U1313 ( .A(n124), .B(n1301), .Z(n1309) );
  XNOR U1314 ( .A(n1299), .B(n1308), .Z(n1301) );
  XNOR U1315 ( .A(n1310), .B(n1311), .Z(n1299) );
  AND U1316 ( .A(n128), .B(n1312), .Z(n1311) );
  XOR U1317 ( .A(p_input[48]), .B(n1310), .Z(n1312) );
  XNOR U1318 ( .A(n1313), .B(n1314), .Z(n1310) );
  AND U1319 ( .A(n132), .B(n1315), .Z(n1314) );
  XOR U1320 ( .A(n1316), .B(n1317), .Z(n1308) );
  AND U1321 ( .A(n136), .B(n1307), .Z(n1317) );
  XNOR U1322 ( .A(n1318), .B(n1305), .Z(n1307) );
  XOR U1323 ( .A(n1319), .B(n1320), .Z(n1305) );
  AND U1324 ( .A(n158), .B(n1321), .Z(n1320) );
  IV U1325 ( .A(n1316), .Z(n1318) );
  XOR U1326 ( .A(n1322), .B(n1323), .Z(n1316) );
  AND U1327 ( .A(n143), .B(n1315), .Z(n1323) );
  XNOR U1328 ( .A(n1313), .B(n1322), .Z(n1315) );
  XNOR U1329 ( .A(n1324), .B(n1325), .Z(n1313) );
  AND U1330 ( .A(n147), .B(n1326), .Z(n1325) );
  XOR U1331 ( .A(p_input[64]), .B(n1324), .Z(n1326) );
  XOR U1332 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n1327), 
        .Z(n1324) );
  AND U1333 ( .A(n150), .B(n1328), .Z(n1327) );
  XOR U1334 ( .A(n1329), .B(n1330), .Z(n1322) );
  AND U1335 ( .A(n154), .B(n1321), .Z(n1330) );
  XNOR U1336 ( .A(n1331), .B(n1319), .Z(n1321) );
  XOR U1337 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n1332), .Z(n1319) );
  AND U1338 ( .A(n166), .B(n1333), .Z(n1332) );
  IV U1339 ( .A(n1329), .Z(n1331) );
  XOR U1340 ( .A(n1334), .B(n1335), .Z(n1329) );
  AND U1341 ( .A(n161), .B(n1328), .Z(n1335) );
  XOR U1342 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n1334), 
        .Z(n1328) );
  XOR U1343 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(n1336), 
        .Z(n1334) );
  AND U1344 ( .A(n163), .B(n1333), .Z(n1336) );
  XOR U1345 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n1333) );
  XNOR U1346 ( .A(n1337), .B(n1338), .Z(n62) );
  AND U1347 ( .A(n1339), .B(n1340), .Z(n1338) );
  XNOR U1348 ( .A(n1337), .B(n1341), .Z(n1340) );
  XOR U1349 ( .A(n1342), .B(n1343), .Z(n1341) );
  AND U1350 ( .A(n65), .B(n1344), .Z(n1343) );
  XNOR U1351 ( .A(n1342), .B(n1345), .Z(n1344) );
  XNOR U1352 ( .A(n1337), .B(n1346), .Z(n1339) );
  XOR U1353 ( .A(n1347), .B(n1348), .Z(n1346) );
  AND U1354 ( .A(n82), .B(n1349), .Z(n1348) );
  XOR U1355 ( .A(n1350), .B(n1351), .Z(n1337) );
  AND U1356 ( .A(n1352), .B(n1353), .Z(n1351) );
  XOR U1357 ( .A(n1354), .B(n1350), .Z(n1353) );
  XNOR U1358 ( .A(n1355), .B(n1356), .Z(n1354) );
  AND U1359 ( .A(n65), .B(n1357), .Z(n1356) );
  XNOR U1360 ( .A(n1358), .B(n1355), .Z(n1357) );
  XNOR U1361 ( .A(n1350), .B(n1359), .Z(n1352) );
  XOR U1362 ( .A(n1360), .B(n1361), .Z(n1359) );
  AND U1363 ( .A(n82), .B(n1362), .Z(n1361) );
  XOR U1364 ( .A(n1363), .B(n1364), .Z(n1350) );
  AND U1365 ( .A(n1365), .B(n1366), .Z(n1364) );
  XOR U1366 ( .A(n1367), .B(n1363), .Z(n1366) );
  XNOR U1367 ( .A(n1368), .B(n1369), .Z(n1367) );
  AND U1368 ( .A(n65), .B(n1370), .Z(n1369) );
  XNOR U1369 ( .A(n1371), .B(n1368), .Z(n1370) );
  XNOR U1370 ( .A(n1363), .B(n1372), .Z(n1365) );
  XOR U1371 ( .A(n1373), .B(n1374), .Z(n1372) );
  AND U1372 ( .A(n82), .B(n1375), .Z(n1374) );
  XOR U1373 ( .A(n1376), .B(n1377), .Z(n1363) );
  AND U1374 ( .A(n1378), .B(n1379), .Z(n1377) );
  XOR U1375 ( .A(n1376), .B(n1380), .Z(n1379) );
  XOR U1376 ( .A(n1381), .B(n1382), .Z(n1380) );
  AND U1377 ( .A(n65), .B(n1383), .Z(n1382) );
  XOR U1378 ( .A(n1384), .B(n1381), .Z(n1383) );
  XNOR U1379 ( .A(n1385), .B(n1376), .Z(n1378) );
  XNOR U1380 ( .A(n1386), .B(n1387), .Z(n1385) );
  AND U1381 ( .A(n82), .B(n1388), .Z(n1387) );
  AND U1382 ( .A(n1389), .B(n1390), .Z(n1376) );
  XNOR U1383 ( .A(n1391), .B(n1392), .Z(n1390) );
  AND U1384 ( .A(n65), .B(n1393), .Z(n1392) );
  XNOR U1385 ( .A(n1394), .B(n1391), .Z(n1393) );
  XNOR U1386 ( .A(n1395), .B(n1396), .Z(n65) );
  AND U1387 ( .A(n1397), .B(n1398), .Z(n1396) );
  XOR U1388 ( .A(n1345), .B(n1395), .Z(n1398) );
  XOR U1389 ( .A(n1399), .B(n1400), .Z(n1345) );
  AND U1390 ( .A(n70), .B(n1401), .Z(n1400) );
  XOR U1391 ( .A(n1402), .B(n1399), .Z(n1401) );
  XNOR U1392 ( .A(n1403), .B(n1395), .Z(n1397) );
  IV U1393 ( .A(n1342), .Z(n1403) );
  XOR U1394 ( .A(n1404), .B(n1405), .Z(n1342) );
  AND U1395 ( .A(n78), .B(n1349), .Z(n1405) );
  XNOR U1396 ( .A(n1404), .B(n1347), .Z(n1349) );
  XOR U1397 ( .A(n1406), .B(n1407), .Z(n1395) );
  AND U1398 ( .A(n1408), .B(n1409), .Z(n1407) );
  XOR U1399 ( .A(n1358), .B(n1406), .Z(n1409) );
  XOR U1400 ( .A(n1410), .B(n1411), .Z(n1358) );
  AND U1401 ( .A(n70), .B(n1412), .Z(n1411) );
  XOR U1402 ( .A(n1413), .B(n1410), .Z(n1412) );
  XOR U1403 ( .A(n1406), .B(n1355), .Z(n1408) );
  XOR U1404 ( .A(n1414), .B(n1415), .Z(n1355) );
  AND U1405 ( .A(n78), .B(n1362), .Z(n1415) );
  XOR U1406 ( .A(n1414), .B(n1416), .Z(n1362) );
  XOR U1407 ( .A(n1417), .B(n1418), .Z(n1406) );
  AND U1408 ( .A(n1419), .B(n1420), .Z(n1418) );
  XOR U1409 ( .A(n1371), .B(n1417), .Z(n1420) );
  XOR U1410 ( .A(n1421), .B(n1422), .Z(n1371) );
  AND U1411 ( .A(n70), .B(n1423), .Z(n1422) );
  XNOR U1412 ( .A(n1424), .B(n1421), .Z(n1423) );
  XOR U1413 ( .A(n1417), .B(n1368), .Z(n1419) );
  XOR U1414 ( .A(n1425), .B(n1426), .Z(n1368) );
  AND U1415 ( .A(n78), .B(n1375), .Z(n1426) );
  XOR U1416 ( .A(n1425), .B(n1427), .Z(n1375) );
  XOR U1417 ( .A(n1428), .B(n1429), .Z(n1417) );
  AND U1418 ( .A(n1430), .B(n1431), .Z(n1429) );
  XOR U1419 ( .A(n1428), .B(n1384), .Z(n1431) );
  XOR U1420 ( .A(n1432), .B(n1433), .Z(n1384) );
  AND U1421 ( .A(n70), .B(n1434), .Z(n1433) );
  XOR U1422 ( .A(n1435), .B(n1432), .Z(n1434) );
  XNOR U1423 ( .A(n1381), .B(n1428), .Z(n1430) );
  XNOR U1424 ( .A(n1436), .B(n1437), .Z(n1381) );
  AND U1425 ( .A(n78), .B(n1388), .Z(n1437) );
  XOR U1426 ( .A(n1436), .B(n1386), .Z(n1388) );
  AND U1427 ( .A(n1391), .B(n1394), .Z(n1428) );
  XOR U1428 ( .A(n1438), .B(n1439), .Z(n1394) );
  AND U1429 ( .A(n70), .B(n1440), .Z(n1439) );
  XNOR U1430 ( .A(n1441), .B(n1442), .Z(n1440) );
  XNOR U1431 ( .A(n1443), .B(n1444), .Z(n70) );
  AND U1432 ( .A(n1445), .B(n1446), .Z(n1444) );
  XOR U1433 ( .A(n1402), .B(n1443), .Z(n1446) );
  AND U1434 ( .A(n1447), .B(n1448), .Z(n1402) );
  XNOR U1435 ( .A(n1399), .B(n1443), .Z(n1445) );
  XNOR U1436 ( .A(n1449), .B(n1450), .Z(n1399) );
  AND U1437 ( .A(n1451), .B(n74), .Z(n1450) );
  AND U1438 ( .A(n1449), .B(n1452), .Z(n1451) );
  XOR U1439 ( .A(n1453), .B(n1454), .Z(n1443) );
  AND U1440 ( .A(n1455), .B(n1456), .Z(n1454) );
  XNOR U1441 ( .A(n1453), .B(n1447), .Z(n1456) );
  IV U1442 ( .A(n1413), .Z(n1447) );
  XOR U1443 ( .A(n1457), .B(n1458), .Z(n1413) );
  XOR U1444 ( .A(n1459), .B(n1448), .Z(n1458) );
  AND U1445 ( .A(n1424), .B(n1460), .Z(n1448) );
  AND U1446 ( .A(n1461), .B(n1462), .Z(n1459) );
  XOR U1447 ( .A(n1463), .B(n1457), .Z(n1461) );
  XNOR U1448 ( .A(n1410), .B(n1453), .Z(n1455) );
  XNOR U1449 ( .A(n1464), .B(n1465), .Z(n1410) );
  AND U1450 ( .A(n74), .B(n1466), .Z(n1465) );
  XNOR U1451 ( .A(n1467), .B(n1468), .Z(n1466) );
  XOR U1452 ( .A(n1469), .B(n1470), .Z(n1453) );
  AND U1453 ( .A(n1471), .B(n1472), .Z(n1470) );
  XNOR U1454 ( .A(n1469), .B(n1424), .Z(n1472) );
  XOR U1455 ( .A(n1473), .B(n1462), .Z(n1424) );
  XNOR U1456 ( .A(n1474), .B(n1457), .Z(n1462) );
  XOR U1457 ( .A(n1475), .B(n1476), .Z(n1457) );
  AND U1458 ( .A(n1477), .B(n1478), .Z(n1476) );
  XOR U1459 ( .A(n1479), .B(n1475), .Z(n1477) );
  XNOR U1460 ( .A(n1480), .B(n1481), .Z(n1474) );
  AND U1461 ( .A(n1482), .B(n1483), .Z(n1481) );
  XOR U1462 ( .A(n1480), .B(n1484), .Z(n1482) );
  XNOR U1463 ( .A(n1463), .B(n1460), .Z(n1473) );
  AND U1464 ( .A(n1485), .B(n1486), .Z(n1460) );
  XOR U1465 ( .A(n1487), .B(n1488), .Z(n1463) );
  AND U1466 ( .A(n1489), .B(n1490), .Z(n1488) );
  XOR U1467 ( .A(n1487), .B(n1491), .Z(n1489) );
  XNOR U1468 ( .A(n1421), .B(n1469), .Z(n1471) );
  XNOR U1469 ( .A(n1492), .B(n1493), .Z(n1421) );
  AND U1470 ( .A(n74), .B(n1494), .Z(n1493) );
  XNOR U1471 ( .A(n1495), .B(n1496), .Z(n1494) );
  XOR U1472 ( .A(n1497), .B(n1498), .Z(n1469) );
  AND U1473 ( .A(n1499), .B(n1500), .Z(n1498) );
  XNOR U1474 ( .A(n1497), .B(n1485), .Z(n1500) );
  IV U1475 ( .A(n1435), .Z(n1485) );
  XNOR U1476 ( .A(n1501), .B(n1478), .Z(n1435) );
  XNOR U1477 ( .A(n1502), .B(n1484), .Z(n1478) );
  XNOR U1478 ( .A(n1503), .B(n1504), .Z(n1484) );
  NOR U1479 ( .A(n1505), .B(n1506), .Z(n1504) );
  XOR U1480 ( .A(n1503), .B(n1507), .Z(n1505) );
  XNOR U1481 ( .A(n1483), .B(n1475), .Z(n1502) );
  XOR U1482 ( .A(n1508), .B(n1509), .Z(n1475) );
  AND U1483 ( .A(n1510), .B(n1511), .Z(n1509) );
  XNOR U1484 ( .A(n1508), .B(n1512), .Z(n1510) );
  XNOR U1485 ( .A(n1513), .B(n1480), .Z(n1483) );
  XOR U1486 ( .A(n1514), .B(n1515), .Z(n1480) );
  AND U1487 ( .A(n1516), .B(n1517), .Z(n1515) );
  XOR U1488 ( .A(n1514), .B(n1518), .Z(n1516) );
  XNOR U1489 ( .A(n1519), .B(n1520), .Z(n1513) );
  NOR U1490 ( .A(n1521), .B(n1522), .Z(n1520) );
  XOR U1491 ( .A(n1519), .B(n1523), .Z(n1521) );
  XNOR U1492 ( .A(n1479), .B(n1486), .Z(n1501) );
  NOR U1493 ( .A(n1441), .B(n1524), .Z(n1486) );
  XOR U1494 ( .A(n1491), .B(n1490), .Z(n1479) );
  XNOR U1495 ( .A(n1525), .B(n1487), .Z(n1490) );
  XOR U1496 ( .A(n1526), .B(n1527), .Z(n1487) );
  AND U1497 ( .A(n1528), .B(n1529), .Z(n1527) );
  XOR U1498 ( .A(n1526), .B(n1530), .Z(n1528) );
  XNOR U1499 ( .A(n1531), .B(n1532), .Z(n1525) );
  NOR U1500 ( .A(n1533), .B(n1534), .Z(n1532) );
  XNOR U1501 ( .A(n1531), .B(n1535), .Z(n1533) );
  XOR U1502 ( .A(n1536), .B(n1537), .Z(n1491) );
  NOR U1503 ( .A(n1538), .B(n1539), .Z(n1537) );
  XNOR U1504 ( .A(n1536), .B(n1540), .Z(n1538) );
  XNOR U1505 ( .A(n1432), .B(n1497), .Z(n1499) );
  XNOR U1506 ( .A(n1541), .B(n1542), .Z(n1432) );
  AND U1507 ( .A(n74), .B(n1543), .Z(n1542) );
  XNOR U1508 ( .A(n1544), .B(n1545), .Z(n1543) );
  AND U1509 ( .A(n1442), .B(n1441), .Z(n1497) );
  XOR U1510 ( .A(n1546), .B(n1524), .Z(n1441) );
  XNOR U1511 ( .A(p_input[0]), .B(p_input[128]), .Z(n1524) );
  XOR U1512 ( .A(n1512), .B(n1511), .Z(n1546) );
  XNOR U1513 ( .A(n1547), .B(n1518), .Z(n1511) );
  XNOR U1514 ( .A(n1507), .B(n1506), .Z(n1518) );
  XOR U1515 ( .A(n1548), .B(n1549), .Z(n1506) );
  IV U1516 ( .A(n1503), .Z(n1549) );
  XNOR U1517 ( .A(p_input[10]), .B(p_input[138]), .Z(n1503) );
  XOR U1518 ( .A(p_input[11]), .B(n1550), .Z(n1548) );
  XOR U1519 ( .A(p_input[12]), .B(p_input[140]), .Z(n1507) );
  XNOR U1520 ( .A(n1517), .B(n1508), .Z(n1547) );
  XOR U1521 ( .A(p_input[129]), .B(p_input[1]), .Z(n1508) );
  XOR U1522 ( .A(n1551), .B(n1523), .Z(n1517) );
  XNOR U1523 ( .A(p_input[143]), .B(p_input[15]), .Z(n1523) );
  XOR U1524 ( .A(n1514), .B(n1522), .Z(n1551) );
  XOR U1525 ( .A(n1552), .B(n1519), .Z(n1522) );
  XOR U1526 ( .A(p_input[13]), .B(p_input[141]), .Z(n1519) );
  XNOR U1527 ( .A(p_input[142]), .B(p_input[14]), .Z(n1552) );
  XOR U1528 ( .A(p_input[137]), .B(p_input[9]), .Z(n1514) );
  XNOR U1529 ( .A(n1530), .B(n1529), .Z(n1512) );
  XNOR U1530 ( .A(n1553), .B(n1535), .Z(n1529) );
  XOR U1531 ( .A(p_input[136]), .B(p_input[8]), .Z(n1535) );
  XOR U1532 ( .A(n1526), .B(n1534), .Z(n1553) );
  XOR U1533 ( .A(n1554), .B(n1531), .Z(n1534) );
  XOR U1534 ( .A(p_input[134]), .B(p_input[6]), .Z(n1531) );
  XNOR U1535 ( .A(p_input[135]), .B(p_input[7]), .Z(n1554) );
  XOR U1536 ( .A(p_input[130]), .B(p_input[2]), .Z(n1526) );
  XNOR U1537 ( .A(n1540), .B(n1539), .Z(n1530) );
  XOR U1538 ( .A(n1555), .B(n1536), .Z(n1539) );
  XOR U1539 ( .A(p_input[131]), .B(p_input[3]), .Z(n1536) );
  XNOR U1540 ( .A(p_input[132]), .B(p_input[4]), .Z(n1555) );
  XOR U1541 ( .A(p_input[133]), .B(p_input[5]), .Z(n1540) );
  IV U1542 ( .A(n1438), .Z(n1442) );
  XOR U1543 ( .A(n1556), .B(n1557), .Z(n1438) );
  AND U1544 ( .A(n74), .B(n1558), .Z(n1557) );
  XNOR U1545 ( .A(n1559), .B(n1560), .Z(n74) );
  AND U1546 ( .A(n1561), .B(n1562), .Z(n1560) );
  XNOR U1547 ( .A(n1449), .B(n1559), .Z(n1562) );
  XNOR U1548 ( .A(n1452), .B(n1559), .Z(n1561) );
  XOR U1549 ( .A(n1563), .B(n1564), .Z(n1559) );
  AND U1550 ( .A(n1565), .B(n1566), .Z(n1564) );
  XOR U1551 ( .A(n1467), .B(n1563), .Z(n1566) );
  XOR U1552 ( .A(n1563), .B(n1468), .Z(n1565) );
  XOR U1553 ( .A(n1567), .B(n1568), .Z(n1563) );
  AND U1554 ( .A(n1569), .B(n1570), .Z(n1568) );
  XOR U1555 ( .A(n1495), .B(n1567), .Z(n1570) );
  XOR U1556 ( .A(n1567), .B(n1496), .Z(n1569) );
  XOR U1557 ( .A(n1571), .B(n1572), .Z(n1567) );
  AND U1558 ( .A(n1573), .B(n1574), .Z(n1572) );
  XOR U1559 ( .A(n1571), .B(n1544), .Z(n1574) );
  XNOR U1560 ( .A(n1575), .B(n1576), .Z(n1391) );
  AND U1561 ( .A(n78), .B(n1577), .Z(n1576) );
  XNOR U1562 ( .A(n1578), .B(n1579), .Z(n78) );
  AND U1563 ( .A(n1580), .B(n1581), .Z(n1579) );
  XNOR U1564 ( .A(n1578), .B(n1404), .Z(n1581) );
  XNOR U1565 ( .A(n1578), .B(n1347), .Z(n1580) );
  XOR U1566 ( .A(n1582), .B(n1583), .Z(n1578) );
  AND U1567 ( .A(n1584), .B(n1585), .Z(n1583) );
  XNOR U1568 ( .A(n1414), .B(n1582), .Z(n1585) );
  XOR U1569 ( .A(n1582), .B(n1416), .Z(n1584) );
  XOR U1570 ( .A(n1586), .B(n1587), .Z(n1582) );
  AND U1571 ( .A(n1588), .B(n1589), .Z(n1587) );
  XOR U1572 ( .A(n1586), .B(n1427), .Z(n1588) );
  IV U1573 ( .A(n1373), .Z(n1427) );
  XOR U1574 ( .A(n1590), .B(n1591), .Z(n1389) );
  AND U1575 ( .A(n82), .B(n1577), .Z(n1591) );
  XNOR U1576 ( .A(n1575), .B(n1590), .Z(n1577) );
  XNOR U1577 ( .A(n1592), .B(n1593), .Z(n82) );
  AND U1578 ( .A(n1594), .B(n1595), .Z(n1593) );
  XNOR U1579 ( .A(n1404), .B(n1592), .Z(n1595) );
  XNOR U1580 ( .A(n1452), .B(n1596), .Z(n1404) );
  AND U1581 ( .A(n1597), .B(n86), .Z(n1596) );
  NOR U1582 ( .A(n1598), .B(n1599), .Z(n1597) );
  XNOR U1583 ( .A(n1592), .B(n1347), .Z(n1594) );
  AND U1584 ( .A(n1600), .B(n1601), .Z(n1347) );
  XOR U1585 ( .A(n1602), .B(n1603), .Z(n1592) );
  AND U1586 ( .A(n1604), .B(n1605), .Z(n1603) );
  XNOR U1587 ( .A(n1602), .B(n1414), .Z(n1605) );
  XOR U1588 ( .A(n1468), .B(n1606), .Z(n1414) );
  AND U1589 ( .A(n86), .B(n1607), .Z(n1606) );
  XOR U1590 ( .A(n1464), .B(n1468), .Z(n1607) );
  XNOR U1591 ( .A(n1360), .B(n1602), .Z(n1604) );
  IV U1592 ( .A(n1416), .Z(n1360) );
  XOR U1593 ( .A(n1608), .B(n1609), .Z(n1416) );
  AND U1594 ( .A(n102), .B(n1610), .Z(n1609) );
  XOR U1595 ( .A(n1586), .B(n1611), .Z(n1602) );
  AND U1596 ( .A(n1612), .B(n1589), .Z(n1611) );
  XNOR U1597 ( .A(n1425), .B(n1586), .Z(n1589) );
  XOR U1598 ( .A(n1496), .B(n1613), .Z(n1425) );
  AND U1599 ( .A(n86), .B(n1614), .Z(n1613) );
  XOR U1600 ( .A(n1492), .B(n1496), .Z(n1614) );
  XNOR U1601 ( .A(n1373), .B(n1586), .Z(n1612) );
  XNOR U1602 ( .A(n1615), .B(n1616), .Z(n1373) );
  AND U1603 ( .A(n102), .B(n1617), .Z(n1616) );
  XOR U1604 ( .A(n1618), .B(n1619), .Z(n1586) );
  AND U1605 ( .A(n1620), .B(n1621), .Z(n1619) );
  XNOR U1606 ( .A(n1618), .B(n1436), .Z(n1621) );
  XOR U1607 ( .A(n1545), .B(n1622), .Z(n1436) );
  AND U1608 ( .A(n86), .B(n1623), .Z(n1622) );
  XOR U1609 ( .A(n1541), .B(n1545), .Z(n1623) );
  XNOR U1610 ( .A(n1624), .B(n1618), .Z(n1620) );
  IV U1611 ( .A(n1386), .Z(n1624) );
  XOR U1612 ( .A(n1625), .B(n1626), .Z(n1386) );
  AND U1613 ( .A(n102), .B(n1627), .Z(n1626) );
  AND U1614 ( .A(n1590), .B(n1575), .Z(n1618) );
  XNOR U1615 ( .A(n1628), .B(n1629), .Z(n1575) );
  AND U1616 ( .A(n86), .B(n1558), .Z(n1629) );
  XNOR U1617 ( .A(n1556), .B(n1628), .Z(n1558) );
  XNOR U1618 ( .A(n1630), .B(n1631), .Z(n86) );
  AND U1619 ( .A(n1632), .B(n1633), .Z(n1631) );
  XNOR U1620 ( .A(n1449), .B(n1630), .Z(n1633) );
  IV U1621 ( .A(n1598), .Z(n1449) );
  AND U1622 ( .A(n1634), .B(n1635), .Z(n1598) );
  IV U1623 ( .A(n1636), .Z(n1634) );
  XNOR U1624 ( .A(n1452), .B(n1630), .Z(n1632) );
  IV U1625 ( .A(n1599), .Z(n1452) );
  NOR U1626 ( .A(n1600), .B(n1601), .Z(n1599) );
  XOR U1627 ( .A(n1637), .B(n1638), .Z(n1630) );
  AND U1628 ( .A(n1639), .B(n1640), .Z(n1638) );
  XNOR U1629 ( .A(n1637), .B(n1464), .Z(n1640) );
  IV U1630 ( .A(n1467), .Z(n1464) );
  XOR U1631 ( .A(n1641), .B(n1642), .Z(n1467) );
  AND U1632 ( .A(n90), .B(n1643), .Z(n1642) );
  XOR U1633 ( .A(n1644), .B(n1641), .Z(n1643) );
  XOR U1634 ( .A(n1468), .B(n1637), .Z(n1639) );
  XOR U1635 ( .A(n1645), .B(n1646), .Z(n1468) );
  AND U1636 ( .A(n98), .B(n1610), .Z(n1646) );
  XOR U1637 ( .A(n1645), .B(n1608), .Z(n1610) );
  XOR U1638 ( .A(n1647), .B(n1648), .Z(n1637) );
  AND U1639 ( .A(n1649), .B(n1650), .Z(n1648) );
  XNOR U1640 ( .A(n1647), .B(n1492), .Z(n1650) );
  IV U1641 ( .A(n1495), .Z(n1492) );
  XOR U1642 ( .A(n1651), .B(n1652), .Z(n1495) );
  AND U1643 ( .A(n90), .B(n1653), .Z(n1652) );
  XNOR U1644 ( .A(n1654), .B(n1651), .Z(n1653) );
  XOR U1645 ( .A(n1496), .B(n1647), .Z(n1649) );
  XOR U1646 ( .A(n1655), .B(n1656), .Z(n1496) );
  AND U1647 ( .A(n98), .B(n1617), .Z(n1656) );
  XOR U1648 ( .A(n1655), .B(n1615), .Z(n1617) );
  XOR U1649 ( .A(n1571), .B(n1657), .Z(n1647) );
  AND U1650 ( .A(n1573), .B(n1658), .Z(n1657) );
  XNOR U1651 ( .A(n1571), .B(n1541), .Z(n1658) );
  IV U1652 ( .A(n1544), .Z(n1541) );
  XOR U1653 ( .A(n1659), .B(n1660), .Z(n1544) );
  AND U1654 ( .A(n90), .B(n1661), .Z(n1660) );
  XOR U1655 ( .A(n1662), .B(n1659), .Z(n1661) );
  XOR U1656 ( .A(n1545), .B(n1571), .Z(n1573) );
  XOR U1657 ( .A(n1663), .B(n1664), .Z(n1545) );
  AND U1658 ( .A(n98), .B(n1627), .Z(n1664) );
  XOR U1659 ( .A(n1663), .B(n1625), .Z(n1627) );
  AND U1660 ( .A(n1628), .B(n1556), .Z(n1571) );
  XNOR U1661 ( .A(n1665), .B(n1666), .Z(n1556) );
  AND U1662 ( .A(n90), .B(n1667), .Z(n1666) );
  XNOR U1663 ( .A(n1668), .B(n1665), .Z(n1667) );
  XNOR U1664 ( .A(n1669), .B(n1670), .Z(n90) );
  NOR U1665 ( .A(n1671), .B(n1672), .Z(n1670) );
  XNOR U1666 ( .A(n1669), .B(n1636), .Z(n1672) );
  NOR U1667 ( .A(n1673), .B(n1674), .Z(n1636) );
  NOR U1668 ( .A(n1669), .B(n1635), .Z(n1671) );
  AND U1669 ( .A(n1675), .B(n1676), .Z(n1635) );
  XOR U1670 ( .A(n1677), .B(n1678), .Z(n1669) );
  AND U1671 ( .A(n1679), .B(n1680), .Z(n1678) );
  XNOR U1672 ( .A(n1677), .B(n1675), .Z(n1680) );
  IV U1673 ( .A(n1644), .Z(n1675) );
  XOR U1674 ( .A(n1681), .B(n1682), .Z(n1644) );
  XOR U1675 ( .A(n1683), .B(n1676), .Z(n1682) );
  AND U1676 ( .A(n1654), .B(n1684), .Z(n1676) );
  AND U1677 ( .A(n1685), .B(n1686), .Z(n1683) );
  XOR U1678 ( .A(n1687), .B(n1681), .Z(n1685) );
  XNOR U1679 ( .A(n1641), .B(n1677), .Z(n1679) );
  XNOR U1680 ( .A(n1688), .B(n1689), .Z(n1641) );
  AND U1681 ( .A(n94), .B(n1690), .Z(n1689) );
  XNOR U1682 ( .A(n1691), .B(n1692), .Z(n1690) );
  XOR U1683 ( .A(n1693), .B(n1694), .Z(n1677) );
  AND U1684 ( .A(n1695), .B(n1696), .Z(n1694) );
  XNOR U1685 ( .A(n1693), .B(n1654), .Z(n1696) );
  XOR U1686 ( .A(n1697), .B(n1686), .Z(n1654) );
  XNOR U1687 ( .A(n1698), .B(n1681), .Z(n1686) );
  XOR U1688 ( .A(n1699), .B(n1700), .Z(n1681) );
  AND U1689 ( .A(n1701), .B(n1702), .Z(n1700) );
  XOR U1690 ( .A(n1703), .B(n1699), .Z(n1701) );
  XNOR U1691 ( .A(n1704), .B(n1705), .Z(n1698) );
  AND U1692 ( .A(n1706), .B(n1707), .Z(n1705) );
  XOR U1693 ( .A(n1704), .B(n1708), .Z(n1706) );
  XNOR U1694 ( .A(n1687), .B(n1684), .Z(n1697) );
  AND U1695 ( .A(n1709), .B(n1710), .Z(n1684) );
  XOR U1696 ( .A(n1711), .B(n1712), .Z(n1687) );
  AND U1697 ( .A(n1713), .B(n1714), .Z(n1712) );
  XOR U1698 ( .A(n1711), .B(n1715), .Z(n1713) );
  XNOR U1699 ( .A(n1651), .B(n1693), .Z(n1695) );
  XNOR U1700 ( .A(n1716), .B(n1717), .Z(n1651) );
  AND U1701 ( .A(n94), .B(n1718), .Z(n1717) );
  XNOR U1702 ( .A(n1719), .B(n1720), .Z(n1718) );
  XOR U1703 ( .A(n1721), .B(n1722), .Z(n1693) );
  AND U1704 ( .A(n1723), .B(n1724), .Z(n1722) );
  XNOR U1705 ( .A(n1721), .B(n1709), .Z(n1724) );
  IV U1706 ( .A(n1662), .Z(n1709) );
  XNOR U1707 ( .A(n1725), .B(n1702), .Z(n1662) );
  XNOR U1708 ( .A(n1726), .B(n1708), .Z(n1702) );
  XOR U1709 ( .A(n1727), .B(n1728), .Z(n1708) );
  NOR U1710 ( .A(n1729), .B(n1730), .Z(n1728) );
  XNOR U1711 ( .A(n1727), .B(n1731), .Z(n1729) );
  XNOR U1712 ( .A(n1707), .B(n1699), .Z(n1726) );
  XOR U1713 ( .A(n1732), .B(n1733), .Z(n1699) );
  AND U1714 ( .A(n1734), .B(n1735), .Z(n1733) );
  XNOR U1715 ( .A(n1732), .B(n1736), .Z(n1734) );
  XNOR U1716 ( .A(n1737), .B(n1704), .Z(n1707) );
  XOR U1717 ( .A(n1738), .B(n1739), .Z(n1704) );
  AND U1718 ( .A(n1740), .B(n1741), .Z(n1739) );
  XOR U1719 ( .A(n1738), .B(n1742), .Z(n1740) );
  XNOR U1720 ( .A(n1743), .B(n1744), .Z(n1737) );
  NOR U1721 ( .A(n1745), .B(n1746), .Z(n1744) );
  XOR U1722 ( .A(n1743), .B(n1747), .Z(n1745) );
  XNOR U1723 ( .A(n1703), .B(n1710), .Z(n1725) );
  NOR U1724 ( .A(n1668), .B(n1748), .Z(n1710) );
  XOR U1725 ( .A(n1715), .B(n1714), .Z(n1703) );
  XNOR U1726 ( .A(n1749), .B(n1711), .Z(n1714) );
  XOR U1727 ( .A(n1750), .B(n1751), .Z(n1711) );
  AND U1728 ( .A(n1752), .B(n1753), .Z(n1751) );
  XOR U1729 ( .A(n1750), .B(n1754), .Z(n1752) );
  XNOR U1730 ( .A(n1755), .B(n1756), .Z(n1749) );
  NOR U1731 ( .A(n1757), .B(n1758), .Z(n1756) );
  XNOR U1732 ( .A(n1755), .B(n1759), .Z(n1757) );
  XOR U1733 ( .A(n1760), .B(n1761), .Z(n1715) );
  NOR U1734 ( .A(n1762), .B(n1763), .Z(n1761) );
  XNOR U1735 ( .A(n1760), .B(n1764), .Z(n1762) );
  XNOR U1736 ( .A(n1659), .B(n1721), .Z(n1723) );
  XNOR U1737 ( .A(n1765), .B(n1766), .Z(n1659) );
  AND U1738 ( .A(n94), .B(n1767), .Z(n1766) );
  XNOR U1739 ( .A(n1768), .B(n1769), .Z(n1767) );
  AND U1740 ( .A(n1665), .B(n1668), .Z(n1721) );
  XOR U1741 ( .A(n1770), .B(n1748), .Z(n1668) );
  XNOR U1742 ( .A(p_input[128]), .B(p_input[16]), .Z(n1748) );
  XOR U1743 ( .A(n1736), .B(n1735), .Z(n1770) );
  XNOR U1744 ( .A(n1771), .B(n1742), .Z(n1735) );
  XNOR U1745 ( .A(n1731), .B(n1730), .Z(n1742) );
  XOR U1746 ( .A(n1772), .B(n1727), .Z(n1730) );
  XOR U1747 ( .A(p_input[138]), .B(p_input[26]), .Z(n1727) );
  XNOR U1748 ( .A(p_input[139]), .B(p_input[27]), .Z(n1772) );
  XOR U1749 ( .A(p_input[140]), .B(p_input[28]), .Z(n1731) );
  XNOR U1750 ( .A(n1741), .B(n1732), .Z(n1771) );
  XOR U1751 ( .A(p_input[129]), .B(p_input[17]), .Z(n1732) );
  XOR U1752 ( .A(n1773), .B(n1747), .Z(n1741) );
  XNOR U1753 ( .A(p_input[143]), .B(p_input[31]), .Z(n1747) );
  XOR U1754 ( .A(n1738), .B(n1746), .Z(n1773) );
  XOR U1755 ( .A(n1774), .B(n1743), .Z(n1746) );
  XOR U1756 ( .A(p_input[141]), .B(p_input[29]), .Z(n1743) );
  XNOR U1757 ( .A(p_input[142]), .B(p_input[30]), .Z(n1774) );
  XOR U1758 ( .A(p_input[137]), .B(p_input[25]), .Z(n1738) );
  XNOR U1759 ( .A(n1754), .B(n1753), .Z(n1736) );
  XNOR U1760 ( .A(n1775), .B(n1759), .Z(n1753) );
  XOR U1761 ( .A(p_input[136]), .B(p_input[24]), .Z(n1759) );
  XOR U1762 ( .A(n1750), .B(n1758), .Z(n1775) );
  XOR U1763 ( .A(n1776), .B(n1755), .Z(n1758) );
  XOR U1764 ( .A(p_input[134]), .B(p_input[22]), .Z(n1755) );
  XNOR U1765 ( .A(p_input[135]), .B(p_input[23]), .Z(n1776) );
  XOR U1766 ( .A(p_input[130]), .B(p_input[18]), .Z(n1750) );
  XNOR U1767 ( .A(n1764), .B(n1763), .Z(n1754) );
  XOR U1768 ( .A(n1777), .B(n1760), .Z(n1763) );
  XOR U1769 ( .A(p_input[131]), .B(p_input[19]), .Z(n1760) );
  XNOR U1770 ( .A(p_input[132]), .B(p_input[20]), .Z(n1777) );
  XOR U1771 ( .A(p_input[133]), .B(p_input[21]), .Z(n1764) );
  XNOR U1772 ( .A(n1778), .B(n1779), .Z(n1665) );
  AND U1773 ( .A(n94), .B(n1780), .Z(n1779) );
  XNOR U1774 ( .A(n1781), .B(n1782), .Z(n94) );
  NOR U1775 ( .A(n1783), .B(n1784), .Z(n1782) );
  XNOR U1776 ( .A(n1781), .B(n1785), .Z(n1784) );
  NOR U1777 ( .A(n1781), .B(n1674), .Z(n1783) );
  XOR U1778 ( .A(n1786), .B(n1787), .Z(n1781) );
  AND U1779 ( .A(n1788), .B(n1789), .Z(n1787) );
  XOR U1780 ( .A(n1691), .B(n1786), .Z(n1789) );
  XOR U1781 ( .A(n1786), .B(n1692), .Z(n1788) );
  XOR U1782 ( .A(n1790), .B(n1791), .Z(n1786) );
  AND U1783 ( .A(n1792), .B(n1793), .Z(n1791) );
  XOR U1784 ( .A(n1719), .B(n1790), .Z(n1793) );
  XOR U1785 ( .A(n1790), .B(n1720), .Z(n1792) );
  XOR U1786 ( .A(n1794), .B(n1795), .Z(n1790) );
  AND U1787 ( .A(n1796), .B(n1797), .Z(n1795) );
  XOR U1788 ( .A(n1794), .B(n1768), .Z(n1797) );
  XNOR U1789 ( .A(n1798), .B(n1799), .Z(n1628) );
  AND U1790 ( .A(n98), .B(n1800), .Z(n1799) );
  XNOR U1791 ( .A(n1801), .B(n1802), .Z(n98) );
  NOR U1792 ( .A(n1803), .B(n1804), .Z(n1802) );
  XOR U1793 ( .A(n1601), .B(n1801), .Z(n1804) );
  NOR U1794 ( .A(n1801), .B(n1600), .Z(n1803) );
  XOR U1795 ( .A(n1805), .B(n1806), .Z(n1801) );
  AND U1796 ( .A(n1807), .B(n1808), .Z(n1806) );
  XOR U1797 ( .A(n1805), .B(n1608), .Z(n1807) );
  XOR U1798 ( .A(n1809), .B(n1810), .Z(n1590) );
  AND U1799 ( .A(n102), .B(n1800), .Z(n1810) );
  XNOR U1800 ( .A(n1798), .B(n1809), .Z(n1800) );
  XNOR U1801 ( .A(n1811), .B(n1812), .Z(n102) );
  NOR U1802 ( .A(n1813), .B(n1814), .Z(n1812) );
  XNOR U1803 ( .A(n1601), .B(n1815), .Z(n1814) );
  IV U1804 ( .A(n1811), .Z(n1815) );
  AND U1805 ( .A(n1816), .B(n1817), .Z(n1601) );
  NOR U1806 ( .A(n1811), .B(n1600), .Z(n1813) );
  AND U1807 ( .A(n1674), .B(n1673), .Z(n1600) );
  IV U1808 ( .A(n1785), .Z(n1673) );
  XOR U1809 ( .A(n1805), .B(n1818), .Z(n1811) );
  AND U1810 ( .A(n1819), .B(n1808), .Z(n1818) );
  XNOR U1811 ( .A(n1645), .B(n1805), .Z(n1808) );
  XOR U1812 ( .A(n1692), .B(n1820), .Z(n1645) );
  AND U1813 ( .A(n105), .B(n1821), .Z(n1820) );
  XOR U1814 ( .A(n1688), .B(n1692), .Z(n1821) );
  XNOR U1815 ( .A(n1822), .B(n1805), .Z(n1819) );
  IV U1816 ( .A(n1608), .Z(n1822) );
  XOR U1817 ( .A(n1823), .B(n1824), .Z(n1608) );
  AND U1818 ( .A(n121), .B(n1825), .Z(n1824) );
  XOR U1819 ( .A(n1826), .B(n1827), .Z(n1805) );
  AND U1820 ( .A(n1828), .B(n1829), .Z(n1827) );
  XNOR U1821 ( .A(n1655), .B(n1826), .Z(n1829) );
  XOR U1822 ( .A(n1720), .B(n1830), .Z(n1655) );
  AND U1823 ( .A(n105), .B(n1831), .Z(n1830) );
  XOR U1824 ( .A(n1716), .B(n1720), .Z(n1831) );
  XOR U1825 ( .A(n1826), .B(n1615), .Z(n1828) );
  XOR U1826 ( .A(n1832), .B(n1833), .Z(n1615) );
  AND U1827 ( .A(n121), .B(n1834), .Z(n1833) );
  XOR U1828 ( .A(n1835), .B(n1836), .Z(n1826) );
  AND U1829 ( .A(n1837), .B(n1838), .Z(n1836) );
  XNOR U1830 ( .A(n1835), .B(n1663), .Z(n1838) );
  XOR U1831 ( .A(n1769), .B(n1839), .Z(n1663) );
  AND U1832 ( .A(n105), .B(n1840), .Z(n1839) );
  XOR U1833 ( .A(n1765), .B(n1769), .Z(n1840) );
  XNOR U1834 ( .A(n1841), .B(n1835), .Z(n1837) );
  IV U1835 ( .A(n1625), .Z(n1841) );
  XOR U1836 ( .A(n1842), .B(n1843), .Z(n1625) );
  AND U1837 ( .A(n121), .B(n1844), .Z(n1843) );
  AND U1838 ( .A(n1809), .B(n1798), .Z(n1835) );
  XNOR U1839 ( .A(n1845), .B(n1846), .Z(n1798) );
  AND U1840 ( .A(n105), .B(n1780), .Z(n1846) );
  XNOR U1841 ( .A(n1778), .B(n1845), .Z(n1780) );
  XNOR U1842 ( .A(n1847), .B(n1848), .Z(n105) );
  NOR U1843 ( .A(n1849), .B(n1850), .Z(n1848) );
  XNOR U1844 ( .A(n1847), .B(n1785), .Z(n1850) );
  NOR U1845 ( .A(n1816), .B(n1817), .Z(n1785) );
  NOR U1846 ( .A(n1847), .B(n1674), .Z(n1849) );
  AND U1847 ( .A(n1851), .B(n1852), .Z(n1674) );
  IV U1848 ( .A(n1853), .Z(n1851) );
  XOR U1849 ( .A(n1854), .B(n1855), .Z(n1847) );
  AND U1850 ( .A(n1856), .B(n1857), .Z(n1855) );
  XNOR U1851 ( .A(n1854), .B(n1688), .Z(n1857) );
  IV U1852 ( .A(n1691), .Z(n1688) );
  XOR U1853 ( .A(n1858), .B(n1859), .Z(n1691) );
  AND U1854 ( .A(n109), .B(n1860), .Z(n1859) );
  XOR U1855 ( .A(n1861), .B(n1858), .Z(n1860) );
  XOR U1856 ( .A(n1692), .B(n1854), .Z(n1856) );
  XOR U1857 ( .A(n1862), .B(n1863), .Z(n1692) );
  AND U1858 ( .A(n117), .B(n1825), .Z(n1863) );
  XOR U1859 ( .A(n1862), .B(n1823), .Z(n1825) );
  XOR U1860 ( .A(n1864), .B(n1865), .Z(n1854) );
  AND U1861 ( .A(n1866), .B(n1867), .Z(n1865) );
  XNOR U1862 ( .A(n1864), .B(n1716), .Z(n1867) );
  IV U1863 ( .A(n1719), .Z(n1716) );
  XOR U1864 ( .A(n1868), .B(n1869), .Z(n1719) );
  AND U1865 ( .A(n109), .B(n1870), .Z(n1869) );
  XNOR U1866 ( .A(n1871), .B(n1868), .Z(n1870) );
  XOR U1867 ( .A(n1720), .B(n1864), .Z(n1866) );
  XOR U1868 ( .A(n1872), .B(n1873), .Z(n1720) );
  AND U1869 ( .A(n117), .B(n1834), .Z(n1873) );
  XOR U1870 ( .A(n1872), .B(n1832), .Z(n1834) );
  XOR U1871 ( .A(n1794), .B(n1874), .Z(n1864) );
  AND U1872 ( .A(n1796), .B(n1875), .Z(n1874) );
  XNOR U1873 ( .A(n1794), .B(n1765), .Z(n1875) );
  IV U1874 ( .A(n1768), .Z(n1765) );
  XOR U1875 ( .A(n1876), .B(n1877), .Z(n1768) );
  AND U1876 ( .A(n109), .B(n1878), .Z(n1877) );
  XOR U1877 ( .A(n1879), .B(n1876), .Z(n1878) );
  XOR U1878 ( .A(n1769), .B(n1794), .Z(n1796) );
  XOR U1879 ( .A(n1880), .B(n1881), .Z(n1769) );
  AND U1880 ( .A(n117), .B(n1844), .Z(n1881) );
  XOR U1881 ( .A(n1880), .B(n1842), .Z(n1844) );
  AND U1882 ( .A(n1845), .B(n1778), .Z(n1794) );
  XNOR U1883 ( .A(n1882), .B(n1883), .Z(n1778) );
  AND U1884 ( .A(n109), .B(n1884), .Z(n1883) );
  XNOR U1885 ( .A(n1885), .B(n1882), .Z(n1884) );
  XNOR U1886 ( .A(n1886), .B(n1887), .Z(n109) );
  NOR U1887 ( .A(n1888), .B(n1889), .Z(n1887) );
  XNOR U1888 ( .A(n1886), .B(n1853), .Z(n1889) );
  NOR U1889 ( .A(n1890), .B(n1891), .Z(n1853) );
  NOR U1890 ( .A(n1886), .B(n1852), .Z(n1888) );
  AND U1891 ( .A(n1892), .B(n1893), .Z(n1852) );
  XOR U1892 ( .A(n1894), .B(n1895), .Z(n1886) );
  AND U1893 ( .A(n1896), .B(n1897), .Z(n1895) );
  XNOR U1894 ( .A(n1894), .B(n1892), .Z(n1897) );
  IV U1895 ( .A(n1861), .Z(n1892) );
  XOR U1896 ( .A(n1898), .B(n1899), .Z(n1861) );
  XOR U1897 ( .A(n1900), .B(n1893), .Z(n1899) );
  AND U1898 ( .A(n1871), .B(n1901), .Z(n1893) );
  AND U1899 ( .A(n1902), .B(n1903), .Z(n1900) );
  XOR U1900 ( .A(n1904), .B(n1898), .Z(n1902) );
  XNOR U1901 ( .A(n1858), .B(n1894), .Z(n1896) );
  XNOR U1902 ( .A(n1905), .B(n1906), .Z(n1858) );
  AND U1903 ( .A(n113), .B(n1907), .Z(n1906) );
  XNOR U1904 ( .A(n1908), .B(n1909), .Z(n1907) );
  XOR U1905 ( .A(n1910), .B(n1911), .Z(n1894) );
  AND U1906 ( .A(n1912), .B(n1913), .Z(n1911) );
  XNOR U1907 ( .A(n1910), .B(n1871), .Z(n1913) );
  XOR U1908 ( .A(n1914), .B(n1903), .Z(n1871) );
  XNOR U1909 ( .A(n1915), .B(n1898), .Z(n1903) );
  XOR U1910 ( .A(n1916), .B(n1917), .Z(n1898) );
  AND U1911 ( .A(n1918), .B(n1919), .Z(n1917) );
  XOR U1912 ( .A(n1920), .B(n1916), .Z(n1918) );
  XNOR U1913 ( .A(n1921), .B(n1922), .Z(n1915) );
  AND U1914 ( .A(n1923), .B(n1924), .Z(n1922) );
  XOR U1915 ( .A(n1921), .B(n1925), .Z(n1923) );
  XNOR U1916 ( .A(n1904), .B(n1901), .Z(n1914) );
  AND U1917 ( .A(n1926), .B(n1927), .Z(n1901) );
  XOR U1918 ( .A(n1928), .B(n1929), .Z(n1904) );
  AND U1919 ( .A(n1930), .B(n1931), .Z(n1929) );
  XOR U1920 ( .A(n1928), .B(n1932), .Z(n1930) );
  XNOR U1921 ( .A(n1868), .B(n1910), .Z(n1912) );
  XNOR U1922 ( .A(n1933), .B(n1934), .Z(n1868) );
  AND U1923 ( .A(n113), .B(n1935), .Z(n1934) );
  XNOR U1924 ( .A(n1936), .B(n1937), .Z(n1935) );
  XOR U1925 ( .A(n1938), .B(n1939), .Z(n1910) );
  AND U1926 ( .A(n1940), .B(n1941), .Z(n1939) );
  XNOR U1927 ( .A(n1938), .B(n1926), .Z(n1941) );
  IV U1928 ( .A(n1879), .Z(n1926) );
  XNOR U1929 ( .A(n1942), .B(n1919), .Z(n1879) );
  XNOR U1930 ( .A(n1943), .B(n1925), .Z(n1919) );
  XOR U1931 ( .A(n1944), .B(n1945), .Z(n1925) );
  NOR U1932 ( .A(n1946), .B(n1947), .Z(n1945) );
  XNOR U1933 ( .A(n1944), .B(n1948), .Z(n1946) );
  XNOR U1934 ( .A(n1924), .B(n1916), .Z(n1943) );
  XOR U1935 ( .A(n1949), .B(n1950), .Z(n1916) );
  AND U1936 ( .A(n1951), .B(n1952), .Z(n1950) );
  XNOR U1937 ( .A(n1949), .B(n1953), .Z(n1951) );
  XNOR U1938 ( .A(n1954), .B(n1921), .Z(n1924) );
  XOR U1939 ( .A(n1955), .B(n1956), .Z(n1921) );
  AND U1940 ( .A(n1957), .B(n1958), .Z(n1956) );
  XOR U1941 ( .A(n1955), .B(n1959), .Z(n1957) );
  XNOR U1942 ( .A(n1960), .B(n1961), .Z(n1954) );
  NOR U1943 ( .A(n1962), .B(n1963), .Z(n1961) );
  XOR U1944 ( .A(n1960), .B(n1964), .Z(n1962) );
  XNOR U1945 ( .A(n1920), .B(n1927), .Z(n1942) );
  NOR U1946 ( .A(n1885), .B(n1965), .Z(n1927) );
  XOR U1947 ( .A(n1932), .B(n1931), .Z(n1920) );
  XNOR U1948 ( .A(n1966), .B(n1928), .Z(n1931) );
  XOR U1949 ( .A(n1967), .B(n1968), .Z(n1928) );
  AND U1950 ( .A(n1969), .B(n1970), .Z(n1968) );
  XOR U1951 ( .A(n1967), .B(n1971), .Z(n1969) );
  XNOR U1952 ( .A(n1972), .B(n1973), .Z(n1966) );
  NOR U1953 ( .A(n1974), .B(n1975), .Z(n1973) );
  XNOR U1954 ( .A(n1972), .B(n1976), .Z(n1974) );
  XOR U1955 ( .A(n1977), .B(n1978), .Z(n1932) );
  NOR U1956 ( .A(n1979), .B(n1980), .Z(n1978) );
  XNOR U1957 ( .A(n1977), .B(n1981), .Z(n1979) );
  XNOR U1958 ( .A(n1876), .B(n1938), .Z(n1940) );
  XNOR U1959 ( .A(n1982), .B(n1983), .Z(n1876) );
  AND U1960 ( .A(n113), .B(n1984), .Z(n1983) );
  XNOR U1961 ( .A(n1985), .B(n1986), .Z(n1984) );
  AND U1962 ( .A(n1882), .B(n1885), .Z(n1938) );
  XOR U1963 ( .A(n1987), .B(n1965), .Z(n1885) );
  XNOR U1964 ( .A(p_input[128]), .B(p_input[32]), .Z(n1965) );
  XOR U1965 ( .A(n1953), .B(n1952), .Z(n1987) );
  XNOR U1966 ( .A(n1988), .B(n1959), .Z(n1952) );
  XNOR U1967 ( .A(n1948), .B(n1947), .Z(n1959) );
  XOR U1968 ( .A(n1989), .B(n1944), .Z(n1947) );
  XOR U1969 ( .A(p_input[138]), .B(p_input[42]), .Z(n1944) );
  XNOR U1970 ( .A(p_input[139]), .B(p_input[43]), .Z(n1989) );
  XOR U1971 ( .A(p_input[140]), .B(p_input[44]), .Z(n1948) );
  XNOR U1972 ( .A(n1958), .B(n1949), .Z(n1988) );
  XOR U1973 ( .A(p_input[129]), .B(p_input[33]), .Z(n1949) );
  XOR U1974 ( .A(n1990), .B(n1964), .Z(n1958) );
  XNOR U1975 ( .A(p_input[143]), .B(p_input[47]), .Z(n1964) );
  XOR U1976 ( .A(n1955), .B(n1963), .Z(n1990) );
  XOR U1977 ( .A(n1991), .B(n1960), .Z(n1963) );
  XOR U1978 ( .A(p_input[141]), .B(p_input[45]), .Z(n1960) );
  XNOR U1979 ( .A(p_input[142]), .B(p_input[46]), .Z(n1991) );
  XOR U1980 ( .A(p_input[137]), .B(p_input[41]), .Z(n1955) );
  XNOR U1981 ( .A(n1971), .B(n1970), .Z(n1953) );
  XNOR U1982 ( .A(n1992), .B(n1976), .Z(n1970) );
  XOR U1983 ( .A(p_input[136]), .B(p_input[40]), .Z(n1976) );
  XOR U1984 ( .A(n1967), .B(n1975), .Z(n1992) );
  XOR U1985 ( .A(n1993), .B(n1972), .Z(n1975) );
  XOR U1986 ( .A(p_input[134]), .B(p_input[38]), .Z(n1972) );
  XNOR U1987 ( .A(p_input[135]), .B(p_input[39]), .Z(n1993) );
  XOR U1988 ( .A(p_input[130]), .B(p_input[34]), .Z(n1967) );
  XNOR U1989 ( .A(n1981), .B(n1980), .Z(n1971) );
  XOR U1990 ( .A(n1994), .B(n1977), .Z(n1980) );
  XOR U1991 ( .A(p_input[131]), .B(p_input[35]), .Z(n1977) );
  XNOR U1992 ( .A(p_input[132]), .B(p_input[36]), .Z(n1994) );
  XOR U1993 ( .A(p_input[133]), .B(p_input[37]), .Z(n1981) );
  XNOR U1994 ( .A(n1995), .B(n1996), .Z(n1882) );
  AND U1995 ( .A(n113), .B(n1997), .Z(n1996) );
  XNOR U1996 ( .A(n1998), .B(n1999), .Z(n113) );
  NOR U1997 ( .A(n2000), .B(n2001), .Z(n1999) );
  XNOR U1998 ( .A(n1998), .B(n2002), .Z(n2001) );
  NOR U1999 ( .A(n1998), .B(n1891), .Z(n2000) );
  XOR U2000 ( .A(n2003), .B(n2004), .Z(n1998) );
  AND U2001 ( .A(n2005), .B(n2006), .Z(n2004) );
  XOR U2002 ( .A(n1908), .B(n2003), .Z(n2006) );
  XOR U2003 ( .A(n2003), .B(n1909), .Z(n2005) );
  XOR U2004 ( .A(n2007), .B(n2008), .Z(n2003) );
  AND U2005 ( .A(n2009), .B(n2010), .Z(n2008) );
  XOR U2006 ( .A(n1936), .B(n2007), .Z(n2010) );
  XOR U2007 ( .A(n2007), .B(n1937), .Z(n2009) );
  XOR U2008 ( .A(n2011), .B(n2012), .Z(n2007) );
  AND U2009 ( .A(n2013), .B(n2014), .Z(n2012) );
  XOR U2010 ( .A(n2011), .B(n1985), .Z(n2014) );
  XNOR U2011 ( .A(n2015), .B(n2016), .Z(n1845) );
  AND U2012 ( .A(n117), .B(n2017), .Z(n2016) );
  XNOR U2013 ( .A(n2018), .B(n2019), .Z(n117) );
  NOR U2014 ( .A(n2020), .B(n2021), .Z(n2019) );
  XOR U2015 ( .A(n1817), .B(n2018), .Z(n2021) );
  NOR U2016 ( .A(n2018), .B(n1816), .Z(n2020) );
  XOR U2017 ( .A(n2022), .B(n2023), .Z(n2018) );
  AND U2018 ( .A(n2024), .B(n2025), .Z(n2023) );
  XOR U2019 ( .A(n2022), .B(n1823), .Z(n2024) );
  XOR U2020 ( .A(n2026), .B(n2027), .Z(n1809) );
  AND U2021 ( .A(n121), .B(n2017), .Z(n2027) );
  XNOR U2022 ( .A(n2015), .B(n2026), .Z(n2017) );
  XNOR U2023 ( .A(n2028), .B(n2029), .Z(n121) );
  NOR U2024 ( .A(n2030), .B(n2031), .Z(n2029) );
  XNOR U2025 ( .A(n1817), .B(n2032), .Z(n2031) );
  IV U2026 ( .A(n2028), .Z(n2032) );
  AND U2027 ( .A(n2033), .B(n2034), .Z(n1817) );
  NOR U2028 ( .A(n2028), .B(n1816), .Z(n2030) );
  AND U2029 ( .A(n1891), .B(n1890), .Z(n1816) );
  IV U2030 ( .A(n2002), .Z(n1890) );
  XOR U2031 ( .A(n2022), .B(n2035), .Z(n2028) );
  AND U2032 ( .A(n2036), .B(n2025), .Z(n2035) );
  XNOR U2033 ( .A(n1862), .B(n2022), .Z(n2025) );
  XOR U2034 ( .A(n1909), .B(n2037), .Z(n1862) );
  AND U2035 ( .A(n124), .B(n2038), .Z(n2037) );
  XOR U2036 ( .A(n1905), .B(n1909), .Z(n2038) );
  XNOR U2037 ( .A(n2039), .B(n2022), .Z(n2036) );
  IV U2038 ( .A(n1823), .Z(n2039) );
  XOR U2039 ( .A(n2040), .B(n2041), .Z(n1823) );
  AND U2040 ( .A(n140), .B(n2042), .Z(n2041) );
  XOR U2041 ( .A(n2043), .B(n2044), .Z(n2022) );
  AND U2042 ( .A(n2045), .B(n2046), .Z(n2044) );
  XNOR U2043 ( .A(n1872), .B(n2043), .Z(n2046) );
  XOR U2044 ( .A(n1937), .B(n2047), .Z(n1872) );
  AND U2045 ( .A(n124), .B(n2048), .Z(n2047) );
  XOR U2046 ( .A(n1933), .B(n1937), .Z(n2048) );
  XOR U2047 ( .A(n2043), .B(n1832), .Z(n2045) );
  XOR U2048 ( .A(n2049), .B(n2050), .Z(n1832) );
  AND U2049 ( .A(n140), .B(n2051), .Z(n2050) );
  XOR U2050 ( .A(n2052), .B(n2053), .Z(n2043) );
  AND U2051 ( .A(n2054), .B(n2055), .Z(n2053) );
  XNOR U2052 ( .A(n2052), .B(n1880), .Z(n2055) );
  XOR U2053 ( .A(n1986), .B(n2056), .Z(n1880) );
  AND U2054 ( .A(n124), .B(n2057), .Z(n2056) );
  XOR U2055 ( .A(n1982), .B(n1986), .Z(n2057) );
  XNOR U2056 ( .A(n2058), .B(n2052), .Z(n2054) );
  IV U2057 ( .A(n1842), .Z(n2058) );
  XOR U2058 ( .A(n2059), .B(n2060), .Z(n1842) );
  AND U2059 ( .A(n140), .B(n2061), .Z(n2060) );
  AND U2060 ( .A(n2026), .B(n2015), .Z(n2052) );
  XNOR U2061 ( .A(n2062), .B(n2063), .Z(n2015) );
  AND U2062 ( .A(n124), .B(n1997), .Z(n2063) );
  XNOR U2063 ( .A(n1995), .B(n2062), .Z(n1997) );
  XNOR U2064 ( .A(n2064), .B(n2065), .Z(n124) );
  NOR U2065 ( .A(n2066), .B(n2067), .Z(n2065) );
  XNOR U2066 ( .A(n2064), .B(n2002), .Z(n2067) );
  NOR U2067 ( .A(n2033), .B(n2034), .Z(n2002) );
  NOR U2068 ( .A(n2064), .B(n1891), .Z(n2066) );
  AND U2069 ( .A(n2068), .B(n2069), .Z(n1891) );
  IV U2070 ( .A(n2070), .Z(n2068) );
  XOR U2071 ( .A(n2071), .B(n2072), .Z(n2064) );
  AND U2072 ( .A(n2073), .B(n2074), .Z(n2072) );
  XNOR U2073 ( .A(n2071), .B(n1905), .Z(n2074) );
  IV U2074 ( .A(n1908), .Z(n1905) );
  XOR U2075 ( .A(n2075), .B(n2076), .Z(n1908) );
  AND U2076 ( .A(n128), .B(n2077), .Z(n2076) );
  XOR U2077 ( .A(n2078), .B(n2075), .Z(n2077) );
  XOR U2078 ( .A(n1909), .B(n2071), .Z(n2073) );
  XOR U2079 ( .A(n2079), .B(n2080), .Z(n1909) );
  AND U2080 ( .A(n136), .B(n2042), .Z(n2080) );
  XOR U2081 ( .A(n2079), .B(n2040), .Z(n2042) );
  XOR U2082 ( .A(n2081), .B(n2082), .Z(n2071) );
  AND U2083 ( .A(n2083), .B(n2084), .Z(n2082) );
  XNOR U2084 ( .A(n2081), .B(n1933), .Z(n2084) );
  IV U2085 ( .A(n1936), .Z(n1933) );
  XOR U2086 ( .A(n2085), .B(n2086), .Z(n1936) );
  AND U2087 ( .A(n128), .B(n2087), .Z(n2086) );
  XNOR U2088 ( .A(n2088), .B(n2085), .Z(n2087) );
  XOR U2089 ( .A(n1937), .B(n2081), .Z(n2083) );
  XOR U2090 ( .A(n2089), .B(n2090), .Z(n1937) );
  AND U2091 ( .A(n136), .B(n2051), .Z(n2090) );
  XOR U2092 ( .A(n2089), .B(n2049), .Z(n2051) );
  XOR U2093 ( .A(n2011), .B(n2091), .Z(n2081) );
  AND U2094 ( .A(n2013), .B(n2092), .Z(n2091) );
  XNOR U2095 ( .A(n2011), .B(n1982), .Z(n2092) );
  IV U2096 ( .A(n1985), .Z(n1982) );
  XOR U2097 ( .A(n2093), .B(n2094), .Z(n1985) );
  AND U2098 ( .A(n128), .B(n2095), .Z(n2094) );
  XOR U2099 ( .A(n2096), .B(n2093), .Z(n2095) );
  XOR U2100 ( .A(n1986), .B(n2011), .Z(n2013) );
  XOR U2101 ( .A(n2097), .B(n2098), .Z(n1986) );
  AND U2102 ( .A(n136), .B(n2061), .Z(n2098) );
  XOR U2103 ( .A(n2097), .B(n2059), .Z(n2061) );
  AND U2104 ( .A(n2062), .B(n1995), .Z(n2011) );
  XNOR U2105 ( .A(n2099), .B(n2100), .Z(n1995) );
  AND U2106 ( .A(n128), .B(n2101), .Z(n2100) );
  XNOR U2107 ( .A(n2102), .B(n2099), .Z(n2101) );
  XNOR U2108 ( .A(n2103), .B(n2104), .Z(n128) );
  NOR U2109 ( .A(n2105), .B(n2106), .Z(n2104) );
  XNOR U2110 ( .A(n2103), .B(n2070), .Z(n2106) );
  NOR U2111 ( .A(n2107), .B(n2108), .Z(n2070) );
  NOR U2112 ( .A(n2103), .B(n2069), .Z(n2105) );
  AND U2113 ( .A(n2109), .B(n2110), .Z(n2069) );
  XOR U2114 ( .A(n2111), .B(n2112), .Z(n2103) );
  AND U2115 ( .A(n2113), .B(n2114), .Z(n2112) );
  XNOR U2116 ( .A(n2111), .B(n2109), .Z(n2114) );
  IV U2117 ( .A(n2078), .Z(n2109) );
  XOR U2118 ( .A(n2115), .B(n2116), .Z(n2078) );
  XOR U2119 ( .A(n2117), .B(n2110), .Z(n2116) );
  AND U2120 ( .A(n2088), .B(n2118), .Z(n2110) );
  AND U2121 ( .A(n2119), .B(n2120), .Z(n2117) );
  XOR U2122 ( .A(n2121), .B(n2115), .Z(n2119) );
  XNOR U2123 ( .A(n2075), .B(n2111), .Z(n2113) );
  XNOR U2124 ( .A(n2122), .B(n2123), .Z(n2075) );
  AND U2125 ( .A(n132), .B(n2124), .Z(n2123) );
  XNOR U2126 ( .A(n2125), .B(n2126), .Z(n2124) );
  XOR U2127 ( .A(n2127), .B(n2128), .Z(n2111) );
  AND U2128 ( .A(n2129), .B(n2130), .Z(n2128) );
  XNOR U2129 ( .A(n2127), .B(n2088), .Z(n2130) );
  XOR U2130 ( .A(n2131), .B(n2120), .Z(n2088) );
  XNOR U2131 ( .A(n2132), .B(n2115), .Z(n2120) );
  XOR U2132 ( .A(n2133), .B(n2134), .Z(n2115) );
  AND U2133 ( .A(n2135), .B(n2136), .Z(n2134) );
  XOR U2134 ( .A(n2137), .B(n2133), .Z(n2135) );
  XNOR U2135 ( .A(n2138), .B(n2139), .Z(n2132) );
  AND U2136 ( .A(n2140), .B(n2141), .Z(n2139) );
  XOR U2137 ( .A(n2138), .B(n2142), .Z(n2140) );
  XNOR U2138 ( .A(n2121), .B(n2118), .Z(n2131) );
  AND U2139 ( .A(n2143), .B(n2144), .Z(n2118) );
  XOR U2140 ( .A(n2145), .B(n2146), .Z(n2121) );
  AND U2141 ( .A(n2147), .B(n2148), .Z(n2146) );
  XOR U2142 ( .A(n2145), .B(n2149), .Z(n2147) );
  XNOR U2143 ( .A(n2085), .B(n2127), .Z(n2129) );
  XNOR U2144 ( .A(n2150), .B(n2151), .Z(n2085) );
  AND U2145 ( .A(n132), .B(n2152), .Z(n2151) );
  XNOR U2146 ( .A(n2153), .B(n2154), .Z(n2152) );
  XOR U2147 ( .A(n2155), .B(n2156), .Z(n2127) );
  AND U2148 ( .A(n2157), .B(n2158), .Z(n2156) );
  XNOR U2149 ( .A(n2155), .B(n2143), .Z(n2158) );
  IV U2150 ( .A(n2096), .Z(n2143) );
  XNOR U2151 ( .A(n2159), .B(n2136), .Z(n2096) );
  XNOR U2152 ( .A(n2160), .B(n2142), .Z(n2136) );
  XOR U2153 ( .A(n2161), .B(n2162), .Z(n2142) );
  NOR U2154 ( .A(n2163), .B(n2164), .Z(n2162) );
  XNOR U2155 ( .A(n2161), .B(n2165), .Z(n2163) );
  XNOR U2156 ( .A(n2141), .B(n2133), .Z(n2160) );
  XOR U2157 ( .A(n2166), .B(n2167), .Z(n2133) );
  AND U2158 ( .A(n2168), .B(n2169), .Z(n2167) );
  XNOR U2159 ( .A(n2166), .B(n2170), .Z(n2168) );
  XNOR U2160 ( .A(n2171), .B(n2138), .Z(n2141) );
  XOR U2161 ( .A(n2172), .B(n2173), .Z(n2138) );
  AND U2162 ( .A(n2174), .B(n2175), .Z(n2173) );
  XOR U2163 ( .A(n2172), .B(n2176), .Z(n2174) );
  XNOR U2164 ( .A(n2177), .B(n2178), .Z(n2171) );
  NOR U2165 ( .A(n2179), .B(n2180), .Z(n2178) );
  XOR U2166 ( .A(n2177), .B(n2181), .Z(n2179) );
  XNOR U2167 ( .A(n2137), .B(n2144), .Z(n2159) );
  NOR U2168 ( .A(n2102), .B(n2182), .Z(n2144) );
  XOR U2169 ( .A(n2149), .B(n2148), .Z(n2137) );
  XNOR U2170 ( .A(n2183), .B(n2145), .Z(n2148) );
  XOR U2171 ( .A(n2184), .B(n2185), .Z(n2145) );
  AND U2172 ( .A(n2186), .B(n2187), .Z(n2185) );
  XOR U2173 ( .A(n2184), .B(n2188), .Z(n2186) );
  XNOR U2174 ( .A(n2189), .B(n2190), .Z(n2183) );
  NOR U2175 ( .A(n2191), .B(n2192), .Z(n2190) );
  XNOR U2176 ( .A(n2189), .B(n2193), .Z(n2191) );
  XOR U2177 ( .A(n2194), .B(n2195), .Z(n2149) );
  NOR U2178 ( .A(n2196), .B(n2197), .Z(n2195) );
  XNOR U2179 ( .A(n2194), .B(n2198), .Z(n2196) );
  XNOR U2180 ( .A(n2093), .B(n2155), .Z(n2157) );
  XNOR U2181 ( .A(n2199), .B(n2200), .Z(n2093) );
  AND U2182 ( .A(n132), .B(n2201), .Z(n2200) );
  XNOR U2183 ( .A(n2202), .B(n2203), .Z(n2201) );
  AND U2184 ( .A(n2099), .B(n2102), .Z(n2155) );
  XOR U2185 ( .A(n2204), .B(n2182), .Z(n2102) );
  XNOR U2186 ( .A(p_input[128]), .B(p_input[48]), .Z(n2182) );
  XOR U2187 ( .A(n2170), .B(n2169), .Z(n2204) );
  XNOR U2188 ( .A(n2205), .B(n2176), .Z(n2169) );
  XNOR U2189 ( .A(n2165), .B(n2164), .Z(n2176) );
  XOR U2190 ( .A(n2206), .B(n2161), .Z(n2164) );
  XOR U2191 ( .A(p_input[138]), .B(p_input[58]), .Z(n2161) );
  XNOR U2192 ( .A(p_input[139]), .B(p_input[59]), .Z(n2206) );
  XOR U2193 ( .A(p_input[140]), .B(p_input[60]), .Z(n2165) );
  XNOR U2194 ( .A(n2175), .B(n2166), .Z(n2205) );
  XOR U2195 ( .A(p_input[129]), .B(p_input[49]), .Z(n2166) );
  XOR U2196 ( .A(n2207), .B(n2181), .Z(n2175) );
  XNOR U2197 ( .A(p_input[143]), .B(p_input[63]), .Z(n2181) );
  XOR U2198 ( .A(n2172), .B(n2180), .Z(n2207) );
  XOR U2199 ( .A(n2208), .B(n2177), .Z(n2180) );
  XOR U2200 ( .A(p_input[141]), .B(p_input[61]), .Z(n2177) );
  XNOR U2201 ( .A(p_input[142]), .B(p_input[62]), .Z(n2208) );
  XOR U2202 ( .A(p_input[137]), .B(p_input[57]), .Z(n2172) );
  XNOR U2203 ( .A(n2188), .B(n2187), .Z(n2170) );
  XNOR U2204 ( .A(n2209), .B(n2193), .Z(n2187) );
  XOR U2205 ( .A(p_input[136]), .B(p_input[56]), .Z(n2193) );
  XOR U2206 ( .A(n2184), .B(n2192), .Z(n2209) );
  XOR U2207 ( .A(n2210), .B(n2189), .Z(n2192) );
  XOR U2208 ( .A(p_input[134]), .B(p_input[54]), .Z(n2189) );
  XNOR U2209 ( .A(p_input[135]), .B(p_input[55]), .Z(n2210) );
  XOR U2210 ( .A(p_input[130]), .B(p_input[50]), .Z(n2184) );
  XNOR U2211 ( .A(n2198), .B(n2197), .Z(n2188) );
  XOR U2212 ( .A(n2211), .B(n2194), .Z(n2197) );
  XOR U2213 ( .A(p_input[131]), .B(p_input[51]), .Z(n2194) );
  XNOR U2214 ( .A(p_input[132]), .B(p_input[52]), .Z(n2211) );
  XOR U2215 ( .A(p_input[133]), .B(p_input[53]), .Z(n2198) );
  XNOR U2216 ( .A(n2212), .B(n2213), .Z(n2099) );
  AND U2217 ( .A(n132), .B(n2214), .Z(n2213) );
  XNOR U2218 ( .A(n2215), .B(n2216), .Z(n132) );
  NOR U2219 ( .A(n2217), .B(n2218), .Z(n2216) );
  XNOR U2220 ( .A(n2215), .B(n2219), .Z(n2218) );
  NOR U2221 ( .A(n2215), .B(n2108), .Z(n2217) );
  XOR U2222 ( .A(n2220), .B(n2221), .Z(n2215) );
  AND U2223 ( .A(n2222), .B(n2223), .Z(n2221) );
  XOR U2224 ( .A(n2125), .B(n2220), .Z(n2223) );
  XOR U2225 ( .A(n2220), .B(n2126), .Z(n2222) );
  XOR U2226 ( .A(n2224), .B(n2225), .Z(n2220) );
  AND U2227 ( .A(n2226), .B(n2227), .Z(n2225) );
  XOR U2228 ( .A(n2153), .B(n2224), .Z(n2227) );
  XOR U2229 ( .A(n2224), .B(n2154), .Z(n2226) );
  XOR U2230 ( .A(n2228), .B(n2229), .Z(n2224) );
  AND U2231 ( .A(n2230), .B(n2231), .Z(n2229) );
  XOR U2232 ( .A(n2228), .B(n2202), .Z(n2231) );
  XNOR U2233 ( .A(n2232), .B(n2233), .Z(n2062) );
  AND U2234 ( .A(n136), .B(n2234), .Z(n2233) );
  XNOR U2235 ( .A(n2235), .B(n2236), .Z(n136) );
  NOR U2236 ( .A(n2237), .B(n2238), .Z(n2236) );
  XOR U2237 ( .A(n2034), .B(n2235), .Z(n2238) );
  NOR U2238 ( .A(n2235), .B(n2033), .Z(n2237) );
  XOR U2239 ( .A(n2239), .B(n2240), .Z(n2235) );
  AND U2240 ( .A(n2241), .B(n2242), .Z(n2240) );
  XOR U2241 ( .A(n2239), .B(n2040), .Z(n2241) );
  XOR U2242 ( .A(n2243), .B(n2244), .Z(n2026) );
  AND U2243 ( .A(n140), .B(n2234), .Z(n2244) );
  XNOR U2244 ( .A(n2232), .B(n2243), .Z(n2234) );
  XNOR U2245 ( .A(n2245), .B(n2246), .Z(n140) );
  NOR U2246 ( .A(n2247), .B(n2248), .Z(n2246) );
  XNOR U2247 ( .A(n2034), .B(n2249), .Z(n2248) );
  IV U2248 ( .A(n2245), .Z(n2249) );
  AND U2249 ( .A(n2250), .B(n2251), .Z(n2034) );
  NOR U2250 ( .A(n2245), .B(n2033), .Z(n2247) );
  AND U2251 ( .A(n2108), .B(n2107), .Z(n2033) );
  IV U2252 ( .A(n2219), .Z(n2107) );
  XOR U2253 ( .A(n2239), .B(n2252), .Z(n2245) );
  AND U2254 ( .A(n2253), .B(n2242), .Z(n2252) );
  XNOR U2255 ( .A(n2079), .B(n2239), .Z(n2242) );
  XOR U2256 ( .A(n2126), .B(n2254), .Z(n2079) );
  AND U2257 ( .A(n143), .B(n2255), .Z(n2254) );
  XOR U2258 ( .A(n2122), .B(n2126), .Z(n2255) );
  XNOR U2259 ( .A(n2256), .B(n2239), .Z(n2253) );
  IV U2260 ( .A(n2040), .Z(n2256) );
  XOR U2261 ( .A(n2257), .B(n2258), .Z(n2040) );
  AND U2262 ( .A(n158), .B(n2259), .Z(n2258) );
  XOR U2263 ( .A(n2260), .B(n2261), .Z(n2239) );
  AND U2264 ( .A(n2262), .B(n2263), .Z(n2261) );
  XNOR U2265 ( .A(n2089), .B(n2260), .Z(n2263) );
  XOR U2266 ( .A(n2154), .B(n2264), .Z(n2089) );
  AND U2267 ( .A(n143), .B(n2265), .Z(n2264) );
  XOR U2268 ( .A(n2150), .B(n2154), .Z(n2265) );
  XOR U2269 ( .A(n2260), .B(n2049), .Z(n2262) );
  XOR U2270 ( .A(n2266), .B(n2267), .Z(n2049) );
  AND U2271 ( .A(n158), .B(n2268), .Z(n2267) );
  XOR U2272 ( .A(n2269), .B(n2270), .Z(n2260) );
  AND U2273 ( .A(n2271), .B(n2272), .Z(n2270) );
  XNOR U2274 ( .A(n2269), .B(n2097), .Z(n2272) );
  XOR U2275 ( .A(n2203), .B(n2273), .Z(n2097) );
  AND U2276 ( .A(n143), .B(n2274), .Z(n2273) );
  XOR U2277 ( .A(n2199), .B(n2203), .Z(n2274) );
  XNOR U2278 ( .A(n2275), .B(n2269), .Z(n2271) );
  IV U2279 ( .A(n2059), .Z(n2275) );
  XOR U2280 ( .A(n2276), .B(n2277), .Z(n2059) );
  AND U2281 ( .A(n158), .B(n2278), .Z(n2277) );
  AND U2282 ( .A(n2243), .B(n2232), .Z(n2269) );
  XNOR U2283 ( .A(n2279), .B(n2280), .Z(n2232) );
  AND U2284 ( .A(n143), .B(n2214), .Z(n2280) );
  XNOR U2285 ( .A(n2212), .B(n2279), .Z(n2214) );
  XNOR U2286 ( .A(n2281), .B(n2282), .Z(n143) );
  NOR U2287 ( .A(n2283), .B(n2284), .Z(n2282) );
  XNOR U2288 ( .A(n2281), .B(n2219), .Z(n2284) );
  NOR U2289 ( .A(n2250), .B(n2251), .Z(n2219) );
  NOR U2290 ( .A(n2281), .B(n2108), .Z(n2283) );
  AND U2291 ( .A(n2285), .B(n2286), .Z(n2108) );
  IV U2292 ( .A(n2287), .Z(n2285) );
  XOR U2293 ( .A(n2288), .B(n2289), .Z(n2281) );
  AND U2294 ( .A(n2290), .B(n2291), .Z(n2289) );
  XNOR U2295 ( .A(n2288), .B(n2122), .Z(n2291) );
  IV U2296 ( .A(n2125), .Z(n2122) );
  XOR U2297 ( .A(n2292), .B(n2293), .Z(n2125) );
  AND U2298 ( .A(n147), .B(n2294), .Z(n2293) );
  XOR U2299 ( .A(n2295), .B(n2292), .Z(n2294) );
  XOR U2300 ( .A(n2126), .B(n2288), .Z(n2290) );
  XOR U2301 ( .A(n2296), .B(n2297), .Z(n2126) );
  AND U2302 ( .A(n154), .B(n2259), .Z(n2297) );
  XOR U2303 ( .A(n2296), .B(n2257), .Z(n2259) );
  XOR U2304 ( .A(n2298), .B(n2299), .Z(n2288) );
  AND U2305 ( .A(n2300), .B(n2301), .Z(n2299) );
  XNOR U2306 ( .A(n2298), .B(n2150), .Z(n2301) );
  IV U2307 ( .A(n2153), .Z(n2150) );
  XOR U2308 ( .A(n2302), .B(n2303), .Z(n2153) );
  AND U2309 ( .A(n147), .B(n2304), .Z(n2303) );
  XNOR U2310 ( .A(n2305), .B(n2302), .Z(n2304) );
  XOR U2311 ( .A(n2154), .B(n2298), .Z(n2300) );
  XOR U2312 ( .A(n2306), .B(n2307), .Z(n2154) );
  AND U2313 ( .A(n154), .B(n2268), .Z(n2307) );
  XOR U2314 ( .A(n2306), .B(n2266), .Z(n2268) );
  XOR U2315 ( .A(n2228), .B(n2308), .Z(n2298) );
  AND U2316 ( .A(n2230), .B(n2309), .Z(n2308) );
  XNOR U2317 ( .A(n2228), .B(n2199), .Z(n2309) );
  IV U2318 ( .A(n2202), .Z(n2199) );
  XOR U2319 ( .A(n2310), .B(n2311), .Z(n2202) );
  AND U2320 ( .A(n147), .B(n2312), .Z(n2311) );
  XOR U2321 ( .A(n2313), .B(n2310), .Z(n2312) );
  XOR U2322 ( .A(n2203), .B(n2228), .Z(n2230) );
  XOR U2323 ( .A(n2314), .B(n2315), .Z(n2203) );
  AND U2324 ( .A(n154), .B(n2278), .Z(n2315) );
  XOR U2325 ( .A(n2314), .B(n2276), .Z(n2278) );
  AND U2326 ( .A(n2279), .B(n2212), .Z(n2228) );
  XNOR U2327 ( .A(n2316), .B(n2317), .Z(n2212) );
  AND U2328 ( .A(n147), .B(n2318), .Z(n2317) );
  XNOR U2329 ( .A(n2319), .B(n2316), .Z(n2318) );
  XNOR U2330 ( .A(n2320), .B(n2321), .Z(n147) );
  NOR U2331 ( .A(n2322), .B(n2323), .Z(n2321) );
  XNOR U2332 ( .A(n2320), .B(n2287), .Z(n2323) );
  NOR U2333 ( .A(n2324), .B(n2325), .Z(n2287) );
  NOR U2334 ( .A(n2320), .B(n2286), .Z(n2322) );
  AND U2335 ( .A(n2326), .B(n2327), .Z(n2286) );
  XOR U2336 ( .A(n2328), .B(n2329), .Z(n2320) );
  AND U2337 ( .A(n2330), .B(n2331), .Z(n2329) );
  XNOR U2338 ( .A(n2328), .B(n2326), .Z(n2331) );
  IV U2339 ( .A(n2295), .Z(n2326) );
  XOR U2340 ( .A(n2332), .B(n2333), .Z(n2295) );
  XOR U2341 ( .A(n2334), .B(n2327), .Z(n2333) );
  AND U2342 ( .A(n2305), .B(n2335), .Z(n2327) );
  AND U2343 ( .A(n2336), .B(n2337), .Z(n2334) );
  XOR U2344 ( .A(n2338), .B(n2332), .Z(n2336) );
  XNOR U2345 ( .A(n2292), .B(n2328), .Z(n2330) );
  XNOR U2346 ( .A(n2339), .B(n2340), .Z(n2292) );
  AND U2347 ( .A(n150), .B(n2341), .Z(n2340) );
  XOR U2348 ( .A(n2342), .B(n2343), .Z(n2328) );
  AND U2349 ( .A(n2344), .B(n2345), .Z(n2343) );
  XNOR U2350 ( .A(n2342), .B(n2305), .Z(n2345) );
  XOR U2351 ( .A(n2346), .B(n2337), .Z(n2305) );
  XNOR U2352 ( .A(n2347), .B(n2332), .Z(n2337) );
  XOR U2353 ( .A(n2348), .B(n2349), .Z(n2332) );
  AND U2354 ( .A(n2350), .B(n2351), .Z(n2349) );
  XOR U2355 ( .A(n2352), .B(n2348), .Z(n2350) );
  XNOR U2356 ( .A(n2353), .B(n2354), .Z(n2347) );
  AND U2357 ( .A(n2355), .B(n2356), .Z(n2354) );
  XOR U2358 ( .A(n2353), .B(n2357), .Z(n2355) );
  XNOR U2359 ( .A(n2338), .B(n2335), .Z(n2346) );
  AND U2360 ( .A(n2358), .B(n2359), .Z(n2335) );
  XOR U2361 ( .A(n2360), .B(n2361), .Z(n2338) );
  AND U2362 ( .A(n2362), .B(n2363), .Z(n2361) );
  XOR U2363 ( .A(n2360), .B(n2364), .Z(n2362) );
  XNOR U2364 ( .A(n2302), .B(n2342), .Z(n2344) );
  XNOR U2365 ( .A(n2365), .B(n2366), .Z(n2302) );
  AND U2366 ( .A(n150), .B(n2367), .Z(n2366) );
  XOR U2367 ( .A(n2368), .B(n2369), .Z(n2342) );
  AND U2368 ( .A(n2370), .B(n2371), .Z(n2369) );
  XNOR U2369 ( .A(n2368), .B(n2358), .Z(n2371) );
  IV U2370 ( .A(n2313), .Z(n2358) );
  XNOR U2371 ( .A(n2372), .B(n2351), .Z(n2313) );
  XNOR U2372 ( .A(n2373), .B(n2357), .Z(n2351) );
  XOR U2373 ( .A(n2374), .B(n2375), .Z(n2357) );
  NOR U2374 ( .A(n2376), .B(n2377), .Z(n2375) );
  XNOR U2375 ( .A(n2374), .B(n2378), .Z(n2376) );
  XNOR U2376 ( .A(n2356), .B(n2348), .Z(n2373) );
  XOR U2377 ( .A(n2379), .B(n2380), .Z(n2348) );
  AND U2378 ( .A(n2381), .B(n2382), .Z(n2380) );
  XNOR U2379 ( .A(n2379), .B(n2383), .Z(n2381) );
  XNOR U2380 ( .A(n2384), .B(n2353), .Z(n2356) );
  XOR U2381 ( .A(n2385), .B(n2386), .Z(n2353) );
  AND U2382 ( .A(n2387), .B(n2388), .Z(n2386) );
  XOR U2383 ( .A(n2385), .B(n2389), .Z(n2387) );
  XNOR U2384 ( .A(n2390), .B(n2391), .Z(n2384) );
  NOR U2385 ( .A(n2392), .B(n2393), .Z(n2391) );
  XOR U2386 ( .A(n2390), .B(n2394), .Z(n2392) );
  XNOR U2387 ( .A(n2352), .B(n2359), .Z(n2372) );
  NOR U2388 ( .A(n2319), .B(n2395), .Z(n2359) );
  XOR U2389 ( .A(n2364), .B(n2363), .Z(n2352) );
  XNOR U2390 ( .A(n2396), .B(n2360), .Z(n2363) );
  XOR U2391 ( .A(n2397), .B(n2398), .Z(n2360) );
  AND U2392 ( .A(n2399), .B(n2400), .Z(n2398) );
  XOR U2393 ( .A(n2397), .B(n2401), .Z(n2399) );
  XNOR U2394 ( .A(n2402), .B(n2403), .Z(n2396) );
  NOR U2395 ( .A(n2404), .B(n2405), .Z(n2403) );
  XNOR U2396 ( .A(n2402), .B(n2406), .Z(n2404) );
  XOR U2397 ( .A(n2407), .B(n2408), .Z(n2364) );
  NOR U2398 ( .A(n2409), .B(n2410), .Z(n2408) );
  XNOR U2399 ( .A(n2407), .B(n2411), .Z(n2409) );
  XNOR U2400 ( .A(n2310), .B(n2368), .Z(n2370) );
  XNOR U2401 ( .A(n2412), .B(n2413), .Z(n2310) );
  AND U2402 ( .A(n150), .B(n2414), .Z(n2413) );
  XNOR U2403 ( .A(n2415), .B(n2416), .Z(n2414) );
  AND U2404 ( .A(n2316), .B(n2319), .Z(n2368) );
  XOR U2405 ( .A(n2417), .B(n2395), .Z(n2319) );
  XNOR U2406 ( .A(p_input[128]), .B(p_input[64]), .Z(n2395) );
  XOR U2407 ( .A(n2383), .B(n2382), .Z(n2417) );
  XNOR U2408 ( .A(n2418), .B(n2389), .Z(n2382) );
  XNOR U2409 ( .A(n2378), .B(n2377), .Z(n2389) );
  XOR U2410 ( .A(n2419), .B(n2374), .Z(n2377) );
  XOR U2411 ( .A(p_input[138]), .B(p_input[74]), .Z(n2374) );
  XNOR U2412 ( .A(p_input[139]), .B(p_input[75]), .Z(n2419) );
  XOR U2413 ( .A(p_input[140]), .B(p_input[76]), .Z(n2378) );
  XNOR U2414 ( .A(n2388), .B(n2379), .Z(n2418) );
  XOR U2415 ( .A(p_input[129]), .B(p_input[65]), .Z(n2379) );
  XOR U2416 ( .A(n2420), .B(n2394), .Z(n2388) );
  XNOR U2417 ( .A(p_input[143]), .B(p_input[79]), .Z(n2394) );
  XOR U2418 ( .A(n2385), .B(n2393), .Z(n2420) );
  XOR U2419 ( .A(n2421), .B(n2390), .Z(n2393) );
  XOR U2420 ( .A(p_input[141]), .B(p_input[77]), .Z(n2390) );
  XNOR U2421 ( .A(p_input[142]), .B(p_input[78]), .Z(n2421) );
  XOR U2422 ( .A(p_input[137]), .B(p_input[73]), .Z(n2385) );
  XNOR U2423 ( .A(n2401), .B(n2400), .Z(n2383) );
  XNOR U2424 ( .A(n2422), .B(n2406), .Z(n2400) );
  XOR U2425 ( .A(p_input[136]), .B(p_input[72]), .Z(n2406) );
  XOR U2426 ( .A(n2397), .B(n2405), .Z(n2422) );
  XOR U2427 ( .A(n2423), .B(n2402), .Z(n2405) );
  XOR U2428 ( .A(p_input[134]), .B(p_input[70]), .Z(n2402) );
  XNOR U2429 ( .A(p_input[135]), .B(p_input[71]), .Z(n2423) );
  XOR U2430 ( .A(p_input[130]), .B(p_input[66]), .Z(n2397) );
  XNOR U2431 ( .A(n2411), .B(n2410), .Z(n2401) );
  XOR U2432 ( .A(n2424), .B(n2407), .Z(n2410) );
  XOR U2433 ( .A(p_input[131]), .B(p_input[67]), .Z(n2407) );
  XNOR U2434 ( .A(p_input[132]), .B(p_input[68]), .Z(n2424) );
  XOR U2435 ( .A(p_input[133]), .B(p_input[69]), .Z(n2411) );
  XNOR U2436 ( .A(n2425), .B(n2426), .Z(n2316) );
  AND U2437 ( .A(n150), .B(n2427), .Z(n2426) );
  XNOR U2438 ( .A(n2428), .B(n2429), .Z(n150) );
  NOR U2439 ( .A(n2430), .B(n2431), .Z(n2429) );
  XOR U2440 ( .A(n2428), .B(n2324), .Z(n2431) );
  XNOR U2441 ( .A(n2432), .B(n2433), .Z(n2279) );
  AND U2442 ( .A(n154), .B(n2434), .Z(n2433) );
  XNOR U2443 ( .A(n2435), .B(n2436), .Z(n154) );
  NOR U2444 ( .A(n2437), .B(n2438), .Z(n2436) );
  XOR U2445 ( .A(n2251), .B(n2435), .Z(n2438) );
  NOR U2446 ( .A(n2435), .B(n2250), .Z(n2437) );
  XOR U2447 ( .A(n2439), .B(n2440), .Z(n2435) );
  AND U2448 ( .A(n2441), .B(n2442), .Z(n2440) );
  XOR U2449 ( .A(n2439), .B(n2257), .Z(n2441) );
  XOR U2450 ( .A(n2443), .B(n2444), .Z(n2243) );
  AND U2451 ( .A(n158), .B(n2434), .Z(n2444) );
  XNOR U2452 ( .A(n2432), .B(n2443), .Z(n2434) );
  XNOR U2453 ( .A(n2445), .B(n2446), .Z(n158) );
  NOR U2454 ( .A(n2447), .B(n2448), .Z(n2446) );
  XNOR U2455 ( .A(n2251), .B(n2449), .Z(n2448) );
  IV U2456 ( .A(n2445), .Z(n2449) );
  AND U2457 ( .A(n2450), .B(n2451), .Z(n2251) );
  NOR U2458 ( .A(n2445), .B(n2250), .Z(n2447) );
  AND U2459 ( .A(n2324), .B(n2325), .Z(n2250) );
  IV U2460 ( .A(n2452), .Z(n2324) );
  XOR U2461 ( .A(n2439), .B(n2453), .Z(n2445) );
  AND U2462 ( .A(n2454), .B(n2442), .Z(n2453) );
  XNOR U2463 ( .A(n2296), .B(n2439), .Z(n2442) );
  XOR U2464 ( .A(n2455), .B(n2456), .Z(n2296) );
  AND U2465 ( .A(n161), .B(n2341), .Z(n2456) );
  XOR U2466 ( .A(n2339), .B(n2455), .Z(n2341) );
  XNOR U2467 ( .A(n2457), .B(n2439), .Z(n2454) );
  IV U2468 ( .A(n2257), .Z(n2457) );
  XOR U2469 ( .A(n2458), .B(n2459), .Z(n2257) );
  AND U2470 ( .A(n166), .B(n2460), .Z(n2459) );
  XOR U2471 ( .A(n2461), .B(n2462), .Z(n2439) );
  AND U2472 ( .A(n2463), .B(n2464), .Z(n2462) );
  XNOR U2473 ( .A(n2306), .B(n2461), .Z(n2464) );
  XOR U2474 ( .A(n2465), .B(n2466), .Z(n2306) );
  AND U2475 ( .A(n161), .B(n2367), .Z(n2466) );
  XOR U2476 ( .A(n2365), .B(n2465), .Z(n2367) );
  XOR U2477 ( .A(n2461), .B(n2266), .Z(n2463) );
  XOR U2478 ( .A(n2467), .B(n2468), .Z(n2266) );
  AND U2479 ( .A(n166), .B(n2469), .Z(n2468) );
  XOR U2480 ( .A(n2470), .B(n2471), .Z(n2461) );
  AND U2481 ( .A(n2472), .B(n2473), .Z(n2471) );
  XNOR U2482 ( .A(n2470), .B(n2314), .Z(n2473) );
  XOR U2483 ( .A(n2416), .B(n2474), .Z(n2314) );
  AND U2484 ( .A(n161), .B(n2475), .Z(n2474) );
  XOR U2485 ( .A(n2412), .B(n2416), .Z(n2475) );
  XNOR U2486 ( .A(n2476), .B(n2470), .Z(n2472) );
  IV U2487 ( .A(n2276), .Z(n2476) );
  XOR U2488 ( .A(n2477), .B(n2478), .Z(n2276) );
  AND U2489 ( .A(n166), .B(n2479), .Z(n2478) );
  AND U2490 ( .A(n2443), .B(n2432), .Z(n2470) );
  XNOR U2491 ( .A(n2480), .B(n2481), .Z(n2432) );
  AND U2492 ( .A(n161), .B(n2427), .Z(n2481) );
  XOR U2493 ( .A(n2482), .B(n2480), .Z(n2427) );
  XNOR U2494 ( .A(n2428), .B(n2483), .Z(n161) );
  NOR U2495 ( .A(n2430), .B(n2484), .Z(n2483) );
  XNOR U2496 ( .A(n2428), .B(n2452), .Z(n2484) );
  NOR U2497 ( .A(n2450), .B(n2451), .Z(n2452) );
  NOR U2498 ( .A(n2428), .B(n2325), .Z(n2430) );
  AND U2499 ( .A(n2339), .B(n2485), .Z(n2325) );
  XOR U2500 ( .A(n2486), .B(n2487), .Z(n2428) );
  AND U2501 ( .A(n2488), .B(n2489), .Z(n2487) );
  XNOR U2502 ( .A(n2339), .B(n2486), .Z(n2489) );
  XNOR U2503 ( .A(n2490), .B(n2491), .Z(n2339) );
  XOR U2504 ( .A(n2492), .B(n2485), .Z(n2491) );
  AND U2505 ( .A(n2365), .B(n2493), .Z(n2485) );
  AND U2506 ( .A(n2494), .B(n2495), .Z(n2492) );
  XOR U2507 ( .A(n2496), .B(n2490), .Z(n2494) );
  XOR U2508 ( .A(n2486), .B(n2455), .Z(n2488) );
  XOR U2509 ( .A(n2497), .B(n2498), .Z(n2455) );
  AND U2510 ( .A(n163), .B(n2460), .Z(n2498) );
  XOR U2511 ( .A(n2497), .B(n2458), .Z(n2460) );
  XOR U2512 ( .A(n2499), .B(n2500), .Z(n2486) );
  AND U2513 ( .A(n2501), .B(n2502), .Z(n2500) );
  XNOR U2514 ( .A(n2365), .B(n2499), .Z(n2502) );
  XOR U2515 ( .A(n2503), .B(n2495), .Z(n2365) );
  XNOR U2516 ( .A(n2504), .B(n2490), .Z(n2495) );
  XOR U2517 ( .A(n2505), .B(n2506), .Z(n2490) );
  AND U2518 ( .A(n2507), .B(n2508), .Z(n2506) );
  XOR U2519 ( .A(n2509), .B(n2505), .Z(n2507) );
  XNOR U2520 ( .A(n2510), .B(n2511), .Z(n2504) );
  AND U2521 ( .A(n2512), .B(n2513), .Z(n2511) );
  XOR U2522 ( .A(n2510), .B(n2514), .Z(n2512) );
  XNOR U2523 ( .A(n2496), .B(n2493), .Z(n2503) );
  AND U2524 ( .A(n2412), .B(n2515), .Z(n2493) );
  XOR U2525 ( .A(n2516), .B(n2517), .Z(n2496) );
  AND U2526 ( .A(n2518), .B(n2519), .Z(n2517) );
  XOR U2527 ( .A(n2516), .B(n2520), .Z(n2518) );
  XOR U2528 ( .A(n2499), .B(n2465), .Z(n2501) );
  XOR U2529 ( .A(n2521), .B(n2522), .Z(n2465) );
  AND U2530 ( .A(n163), .B(n2469), .Z(n2522) );
  XOR U2531 ( .A(n2521), .B(n2467), .Z(n2469) );
  XOR U2532 ( .A(n2523), .B(n2524), .Z(n2499) );
  AND U2533 ( .A(n2525), .B(n2526), .Z(n2524) );
  XNOR U2534 ( .A(n2523), .B(n2412), .Z(n2526) );
  IV U2535 ( .A(n2415), .Z(n2412) );
  XNOR U2536 ( .A(n2527), .B(n2508), .Z(n2415) );
  XNOR U2537 ( .A(n2528), .B(n2514), .Z(n2508) );
  XOR U2538 ( .A(n2529), .B(n2530), .Z(n2514) );
  NOR U2539 ( .A(n2531), .B(n2532), .Z(n2530) );
  XNOR U2540 ( .A(n2529), .B(n2533), .Z(n2531) );
  XNOR U2541 ( .A(n2513), .B(n2505), .Z(n2528) );
  XOR U2542 ( .A(n2534), .B(n2535), .Z(n2505) );
  AND U2543 ( .A(n2536), .B(n2537), .Z(n2535) );
  XNOR U2544 ( .A(n2534), .B(n2538), .Z(n2536) );
  XNOR U2545 ( .A(n2539), .B(n2510), .Z(n2513) );
  XOR U2546 ( .A(n2540), .B(n2541), .Z(n2510) );
  AND U2547 ( .A(n2542), .B(n2543), .Z(n2541) );
  XNOR U2548 ( .A(n2544), .B(n2545), .Z(n2542) );
  XNOR U2549 ( .A(n2546), .B(n2547), .Z(n2539) );
  NOR U2550 ( .A(n2548), .B(n2549), .Z(n2547) );
  XOR U2551 ( .A(n2546), .B(n2550), .Z(n2548) );
  XNOR U2552 ( .A(n2509), .B(n2515), .Z(n2527) );
  AND U2553 ( .A(n2482), .B(n2551), .Z(n2515) );
  IV U2554 ( .A(n2425), .Z(n2482) );
  XOR U2555 ( .A(n2520), .B(n2519), .Z(n2509) );
  XNOR U2556 ( .A(n2552), .B(n2516), .Z(n2519) );
  XOR U2557 ( .A(n2553), .B(n2554), .Z(n2516) );
  AND U2558 ( .A(n2555), .B(n2556), .Z(n2554) );
  XNOR U2559 ( .A(n2557), .B(n2558), .Z(n2555) );
  XNOR U2560 ( .A(n2559), .B(n2560), .Z(n2552) );
  AND U2561 ( .A(n2561), .B(n2562), .Z(n2560) );
  XNOR U2562 ( .A(n2559), .B(n2563), .Z(n2561) );
  XOR U2563 ( .A(n2564), .B(n2565), .Z(n2520) );
  AND U2564 ( .A(n2566), .B(n2567), .Z(n2565) );
  XOR U2565 ( .A(n2564), .B(n2568), .Z(n2566) );
  XOR U2566 ( .A(n2416), .B(n2523), .Z(n2525) );
  XOR U2567 ( .A(n2569), .B(n2570), .Z(n2416) );
  AND U2568 ( .A(n163), .B(n2479), .Z(n2570) );
  XOR U2569 ( .A(n2569), .B(n2477), .Z(n2479) );
  AND U2570 ( .A(n2480), .B(n2425), .Z(n2523) );
  XNOR U2571 ( .A(n2571), .B(n2551), .Z(n2425) );
  XOR U2572 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(
        p_input[128]), .Z(n2551) );
  XOR U2573 ( .A(n2538), .B(n2537), .Z(n2571) );
  XNOR U2574 ( .A(n2572), .B(n2545), .Z(n2537) );
  XNOR U2575 ( .A(n2533), .B(n2532), .Z(n2545) );
  XOR U2576 ( .A(n2573), .B(n2529), .Z(n2532) );
  XOR U2577 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(
        p_input[138]), .Z(n2529) );
  XOR U2578 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n1550), 
        .Z(n2573) );
  XOR U2579 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(
        p_input[140]), .Z(n2533) );
  XNOR U2580 ( .A(n2543), .B(n2534), .Z(n2572) );
  XOR U2581 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(
        p_input[129]), .Z(n2534) );
  XOR U2582 ( .A(n2574), .B(n2550), .Z(n2543) );
  XNOR U2583 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(
        p_input[143]), .Z(n2550) );
  XOR U2584 ( .A(n2540), .B(n2549), .Z(n2574) );
  XOR U2585 ( .A(n2575), .B(n2546), .Z(n2549) );
  XOR U2586 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(
        p_input[141]), .Z(n2546) );
  XNOR U2587 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(
        p_input[142]), .Z(n2575) );
  IV U2588 ( .A(n2544), .Z(n2540) );
  XNOR U2589 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(
        p_input[137]), .Z(n2544) );
  XNOR U2590 ( .A(n2558), .B(n2556), .Z(n2538) );
  XOR U2591 ( .A(n2576), .B(n2563), .Z(n2556) );
  XNOR U2592 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(
        p_input[136]), .Z(n2563) );
  XNOR U2593 ( .A(n2553), .B(n2562), .Z(n2576) );
  XNOR U2594 ( .A(n2577), .B(n2559), .Z(n2562) );
  XOR U2595 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(
        p_input[134]), .Z(n2559) );
  XNOR U2596 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(
        p_input[135]), .Z(n2577) );
  IV U2597 ( .A(n2557), .Z(n2553) );
  XNOR U2598 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(
        p_input[130]), .Z(n2557) );
  XOR U2599 ( .A(n2568), .B(n2567), .Z(n2558) );
  XNOR U2600 ( .A(n2578), .B(n2564), .Z(n2567) );
  XOR U2601 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(
        p_input[131]), .Z(n2564) );
  XNOR U2602 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(
        p_input[132]), .Z(n2578) );
  XOR U2603 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(
        p_input[133]), .Z(n2568) );
  XNOR U2604 ( .A(n2579), .B(n2580), .Z(n2480) );
  AND U2605 ( .A(n163), .B(n2581), .Z(n2580) );
  XNOR U2606 ( .A(n2582), .B(n2583), .Z(n163) );
  NOR U2607 ( .A(n2584), .B(n2585), .Z(n2583) );
  XOR U2608 ( .A(n2451), .B(n2582), .Z(n2585) );
  NOR U2609 ( .A(n2582), .B(n2450), .Z(n2584) );
  XOR U2610 ( .A(n2586), .B(n2587), .Z(n2582) );
  AND U2611 ( .A(n2588), .B(n2589), .Z(n2587) );
  XOR U2612 ( .A(n2586), .B(n2458), .Z(n2588) );
  XOR U2613 ( .A(n2590), .B(n2591), .Z(n2443) );
  AND U2614 ( .A(n166), .B(n2581), .Z(n2591) );
  XOR U2615 ( .A(n2592), .B(n2590), .Z(n2581) );
  XNOR U2616 ( .A(n2593), .B(n2594), .Z(n166) );
  NOR U2617 ( .A(n2595), .B(n2596), .Z(n2594) );
  XNOR U2618 ( .A(n2451), .B(n2597), .Z(n2596) );
  IV U2619 ( .A(n2593), .Z(n2597) );
  AND U2620 ( .A(n2458), .B(n2598), .Z(n2451) );
  NOR U2621 ( .A(n2593), .B(n2450), .Z(n2595) );
  AND U2622 ( .A(n2497), .B(n2599), .Z(n2450) );
  XOR U2623 ( .A(n2586), .B(n2600), .Z(n2593) );
  AND U2624 ( .A(n2601), .B(n2589), .Z(n2600) );
  XNOR U2625 ( .A(n2497), .B(n2586), .Z(n2589) );
  XNOR U2626 ( .A(n2602), .B(n2603), .Z(n2497) );
  XOR U2627 ( .A(n2604), .B(n2599), .Z(n2603) );
  AND U2628 ( .A(n2521), .B(n2605), .Z(n2599) );
  AND U2629 ( .A(n2606), .B(n2607), .Z(n2604) );
  XOR U2630 ( .A(n2608), .B(n2602), .Z(n2606) );
  XNOR U2631 ( .A(n2609), .B(n2586), .Z(n2601) );
  IV U2632 ( .A(n2458), .Z(n2609) );
  XNOR U2633 ( .A(n2610), .B(n2611), .Z(n2458) );
  XOR U2634 ( .A(n2612), .B(n2598), .Z(n2611) );
  AND U2635 ( .A(n2467), .B(n2613), .Z(n2598) );
  AND U2636 ( .A(n2614), .B(n2615), .Z(n2612) );
  XNOR U2637 ( .A(n2610), .B(n2616), .Z(n2614) );
  XOR U2638 ( .A(n2617), .B(n2618), .Z(n2586) );
  AND U2639 ( .A(n2619), .B(n2620), .Z(n2618) );
  XNOR U2640 ( .A(n2521), .B(n2617), .Z(n2620) );
  XOR U2641 ( .A(n2621), .B(n2607), .Z(n2521) );
  XNOR U2642 ( .A(n2622), .B(n2602), .Z(n2607) );
  XOR U2643 ( .A(n2623), .B(n2624), .Z(n2602) );
  AND U2644 ( .A(n2625), .B(n2626), .Z(n2624) );
  XOR U2645 ( .A(n2627), .B(n2623), .Z(n2625) );
  XNOR U2646 ( .A(n2628), .B(n2629), .Z(n2622) );
  AND U2647 ( .A(n2630), .B(n2631), .Z(n2629) );
  XOR U2648 ( .A(n2628), .B(n2632), .Z(n2630) );
  XNOR U2649 ( .A(n2608), .B(n2605), .Z(n2621) );
  AND U2650 ( .A(n2569), .B(n2633), .Z(n2605) );
  XOR U2651 ( .A(n2634), .B(n2635), .Z(n2608) );
  AND U2652 ( .A(n2636), .B(n2637), .Z(n2635) );
  XOR U2653 ( .A(n2634), .B(n2638), .Z(n2636) );
  XOR U2654 ( .A(n2617), .B(n2467), .Z(n2619) );
  XNOR U2655 ( .A(n2639), .B(n2616), .Z(n2467) );
  XNOR U2656 ( .A(n2640), .B(n2641), .Z(n2616) );
  AND U2657 ( .A(n2642), .B(n2643), .Z(n2641) );
  XOR U2658 ( .A(n2640), .B(n2644), .Z(n2642) );
  XNOR U2659 ( .A(n2615), .B(n2613), .Z(n2639) );
  AND U2660 ( .A(n2477), .B(n2645), .Z(n2613) );
  XNOR U2661 ( .A(n2646), .B(n2610), .Z(n2615) );
  XOR U2662 ( .A(n2647), .B(n2648), .Z(n2610) );
  AND U2663 ( .A(n2649), .B(n2650), .Z(n2648) );
  XOR U2664 ( .A(n2647), .B(n2651), .Z(n2649) );
  XNOR U2665 ( .A(n2652), .B(n2653), .Z(n2646) );
  AND U2666 ( .A(n2654), .B(n2655), .Z(n2653) );
  XNOR U2667 ( .A(n2652), .B(n2656), .Z(n2654) );
  XOR U2668 ( .A(n2657), .B(n2658), .Z(n2617) );
  AND U2669 ( .A(n2659), .B(n2660), .Z(n2658) );
  XNOR U2670 ( .A(n2657), .B(n2569), .Z(n2660) );
  XOR U2671 ( .A(n2661), .B(n2626), .Z(n2569) );
  XNOR U2672 ( .A(n2662), .B(n2632), .Z(n2626) );
  XOR U2673 ( .A(n2663), .B(n2664), .Z(n2632) );
  NOR U2674 ( .A(n2665), .B(n2666), .Z(n2664) );
  XNOR U2675 ( .A(n2663), .B(n2667), .Z(n2665) );
  XNOR U2676 ( .A(n2631), .B(n2623), .Z(n2662) );
  XOR U2677 ( .A(n2668), .B(n2669), .Z(n2623) );
  AND U2678 ( .A(n2670), .B(n2671), .Z(n2669) );
  XNOR U2679 ( .A(n2668), .B(n2672), .Z(n2670) );
  XNOR U2680 ( .A(n2673), .B(n2628), .Z(n2631) );
  XOR U2681 ( .A(n2674), .B(n2675), .Z(n2628) );
  AND U2682 ( .A(n2676), .B(n2677), .Z(n2675) );
  XOR U2683 ( .A(n2674), .B(n2678), .Z(n2676) );
  XNOR U2684 ( .A(n2679), .B(n2680), .Z(n2673) );
  NOR U2685 ( .A(n2681), .B(n2682), .Z(n2680) );
  XOR U2686 ( .A(n2679), .B(n2683), .Z(n2681) );
  XNOR U2687 ( .A(n2627), .B(n2633), .Z(n2661) );
  AND U2688 ( .A(n2592), .B(n2684), .Z(n2633) );
  IV U2689 ( .A(n2579), .Z(n2592) );
  XOR U2690 ( .A(n2638), .B(n2637), .Z(n2627) );
  XNOR U2691 ( .A(n2685), .B(n2634), .Z(n2637) );
  XOR U2692 ( .A(n2686), .B(n2687), .Z(n2634) );
  AND U2693 ( .A(n2688), .B(n2689), .Z(n2687) );
  XOR U2694 ( .A(n2686), .B(n2690), .Z(n2688) );
  XNOR U2695 ( .A(n2691), .B(n2692), .Z(n2685) );
  NOR U2696 ( .A(n2693), .B(n2694), .Z(n2692) );
  XNOR U2697 ( .A(n2691), .B(n2695), .Z(n2693) );
  XOR U2698 ( .A(n2696), .B(n2697), .Z(n2638) );
  NOR U2699 ( .A(n2698), .B(n2699), .Z(n2697) );
  XNOR U2700 ( .A(n2696), .B(n2700), .Z(n2698) );
  XNOR U2701 ( .A(n2701), .B(n2657), .Z(n2659) );
  IV U2702 ( .A(n2477), .Z(n2701) );
  XOR U2703 ( .A(n2702), .B(n2651), .Z(n2477) );
  XOR U2704 ( .A(n2644), .B(n2643), .Z(n2651) );
  XNOR U2705 ( .A(n2703), .B(n2640), .Z(n2643) );
  XOR U2706 ( .A(n2704), .B(n2705), .Z(n2640) );
  AND U2707 ( .A(n2706), .B(n2707), .Z(n2705) );
  XOR U2708 ( .A(n2704), .B(n2708), .Z(n2706) );
  XNOR U2709 ( .A(n2709), .B(n2710), .Z(n2703) );
  NOR U2710 ( .A(n2711), .B(n2712), .Z(n2710) );
  XNOR U2711 ( .A(n2709), .B(n2713), .Z(n2711) );
  XOR U2712 ( .A(n2714), .B(n2715), .Z(n2644) );
  NOR U2713 ( .A(n2716), .B(n2717), .Z(n2715) );
  XNOR U2714 ( .A(n2714), .B(n2718), .Z(n2716) );
  XNOR U2715 ( .A(n2650), .B(n2645), .Z(n2702) );
  AND U2716 ( .A(n2590), .B(n2719), .Z(n2645) );
  XOR U2717 ( .A(n2720), .B(n2656), .Z(n2650) );
  XNOR U2718 ( .A(n2721), .B(n2722), .Z(n2656) );
  NOR U2719 ( .A(n2723), .B(n2724), .Z(n2722) );
  XNOR U2720 ( .A(n2721), .B(n2725), .Z(n2723) );
  XNOR U2721 ( .A(n2655), .B(n2647), .Z(n2720) );
  XOR U2722 ( .A(n2726), .B(n2727), .Z(n2647) );
  AND U2723 ( .A(n2728), .B(n2729), .Z(n2727) );
  XOR U2724 ( .A(n2726), .B(n2730), .Z(n2728) );
  XNOR U2725 ( .A(n2731), .B(n2652), .Z(n2655) );
  XOR U2726 ( .A(n2732), .B(n2733), .Z(n2652) );
  AND U2727 ( .A(n2734), .B(n2735), .Z(n2733) );
  XOR U2728 ( .A(n2732), .B(n2736), .Z(n2734) );
  XNOR U2729 ( .A(n2737), .B(n2738), .Z(n2731) );
  NOR U2730 ( .A(n2739), .B(n2740), .Z(n2738) );
  XOR U2731 ( .A(n2737), .B(n2741), .Z(n2739) );
  AND U2732 ( .A(n2590), .B(n2579), .Z(n2657) );
  XNOR U2733 ( .A(n2742), .B(n2684), .Z(n2579) );
  XOR U2734 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(
        p_input[128]), .Z(n2684) );
  XOR U2735 ( .A(n2672), .B(n2671), .Z(n2742) );
  XNOR U2736 ( .A(n2743), .B(n2678), .Z(n2671) );
  XNOR U2737 ( .A(n2667), .B(n2666), .Z(n2678) );
  XOR U2738 ( .A(n2744), .B(n2663), .Z(n2666) );
  XOR U2739 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(
        p_input[138]), .Z(n2663) );
  XOR U2740 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n1550), 
        .Z(n2744) );
  XOR U2741 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(
        p_input[140]), .Z(n2667) );
  XNOR U2742 ( .A(n2677), .B(n2668), .Z(n2743) );
  XOR U2743 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(
        p_input[129]), .Z(n2668) );
  XOR U2744 ( .A(n2745), .B(n2683), .Z(n2677) );
  XNOR U2745 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(
        p_input[143]), .Z(n2683) );
  XOR U2746 ( .A(n2674), .B(n2682), .Z(n2745) );
  XOR U2747 ( .A(n2746), .B(n2679), .Z(n2682) );
  XOR U2748 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(
        p_input[141]), .Z(n2679) );
  XOR U2749 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n2747), 
        .Z(n2746) );
  XNOR U2750 ( .A(n168), .B(p_input[137]), .Z(n2674) );
  IV U2751 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n168) );
  XNOR U2752 ( .A(n2690), .B(n2689), .Z(n2672) );
  XNOR U2753 ( .A(n2748), .B(n2695), .Z(n2689) );
  XNOR U2754 ( .A(n247), .B(p_input[136]), .Z(n2695) );
  IV U2755 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n247) );
  XOR U2756 ( .A(n2686), .B(n2694), .Z(n2748) );
  XOR U2757 ( .A(n2749), .B(n2691), .Z(n2694) );
  XNOR U2758 ( .A(n405), .B(p_input[134]), .Z(n2691) );
  IV U2759 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n405) );
  XOR U2760 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(n2750), 
        .Z(n2749) );
  XOR U2761 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(
        p_input[130]), .Z(n2686) );
  XNOR U2762 ( .A(n2700), .B(n2699), .Z(n2690) );
  XOR U2763 ( .A(n2751), .B(n2696), .Z(n2699) );
  XNOR U2764 ( .A(n644), .B(p_input[131]), .Z(n2696) );
  IV U2765 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n644) );
  XOR U2766 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n2752), 
        .Z(n2751) );
  XNOR U2767 ( .A(n484), .B(p_input[133]), .Z(n2700) );
  IV U2768 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n484) );
  XOR U2769 ( .A(n2753), .B(n2730), .Z(n2590) );
  XOR U2770 ( .A(n2708), .B(n2707), .Z(n2730) );
  XNOR U2771 ( .A(n2754), .B(n2713), .Z(n2707) );
  XNOR U2772 ( .A(n246), .B(p_input[136]), .Z(n2713) );
  IV U2773 ( .A(\knn_comb_/min_val_out[0][8] ), .Z(n246) );
  XOR U2774 ( .A(n2704), .B(n2712), .Z(n2754) );
  XOR U2775 ( .A(n2755), .B(n2709), .Z(n2712) );
  XNOR U2776 ( .A(n404), .B(p_input[134]), .Z(n2709) );
  IV U2777 ( .A(\knn_comb_/min_val_out[0][6] ), .Z(n404) );
  XOR U2778 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n2750), .Z(n2755) );
  IV U2779 ( .A(p_input[135]), .Z(n2750) );
  XOR U2780 ( .A(\knn_comb_/min_val_out[0][2] ), .B(p_input[130]), .Z(n2704)
         );
  XNOR U2781 ( .A(n2718), .B(n2717), .Z(n2708) );
  XOR U2782 ( .A(n2756), .B(n2714), .Z(n2717) );
  XNOR U2783 ( .A(n643), .B(p_input[131]), .Z(n2714) );
  IV U2784 ( .A(\knn_comb_/min_val_out[0][3] ), .Z(n643) );
  XOR U2785 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n2752), .Z(n2756) );
  IV U2786 ( .A(p_input[132]), .Z(n2752) );
  XNOR U2787 ( .A(n483), .B(p_input[133]), .Z(n2718) );
  IV U2788 ( .A(\knn_comb_/min_val_out[0][5] ), .Z(n483) );
  XNOR U2789 ( .A(n2729), .B(n2719), .Z(n2753) );
  XOR U2790 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[128]), .Z(n2719)
         );
  XNOR U2791 ( .A(n2757), .B(n2736), .Z(n2729) );
  XNOR U2792 ( .A(n2725), .B(n2724), .Z(n2736) );
  XOR U2793 ( .A(n2758), .B(n2721), .Z(n2724) );
  XOR U2794 ( .A(\knn_comb_/min_val_out[0][10] ), .B(p_input[138]), .Z(n2721)
         );
  XOR U2795 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n1550), .Z(n2758) );
  IV U2796 ( .A(p_input[139]), .Z(n1550) );
  XOR U2797 ( .A(\knn_comb_/min_val_out[0][12] ), .B(p_input[140]), .Z(n2725)
         );
  XNOR U2798 ( .A(n2735), .B(n2726), .Z(n2757) );
  XOR U2799 ( .A(\knn_comb_/min_val_out[0][1] ), .B(p_input[129]), .Z(n2726)
         );
  XOR U2800 ( .A(n2759), .B(n2741), .Z(n2735) );
  XNOR U2801 ( .A(\knn_comb_/min_val_out[0][15] ), .B(p_input[143]), .Z(n2741)
         );
  XOR U2802 ( .A(n2732), .B(n2740), .Z(n2759) );
  XOR U2803 ( .A(n2760), .B(n2737), .Z(n2740) );
  XOR U2804 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[141]), .Z(n2737)
         );
  XOR U2805 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n2747), .Z(n2760) );
  IV U2806 ( .A(p_input[142]), .Z(n2747) );
  XNOR U2807 ( .A(n167), .B(p_input[137]), .Z(n2732) );
  IV U2808 ( .A(\knn_comb_/min_val_out[0][9] ), .Z(n167) );
endmodule

