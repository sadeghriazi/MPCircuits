
module voting_N2_M3 ( p_input, o );
  input [15:0] p_input;
  output [1:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221;

  XOR U2 ( .A(n1), .B(n2), .Z(o[0]) );
  AND U3 ( .A(o[1]), .B(n3), .Z(n1) );
  XOR U4 ( .A(n4), .B(n2), .Z(n3) );
  XOR U5 ( .A(n5), .B(n6), .Z(o[1]) );
  MUX U6 ( .IN0(n7), .IN1(n8), .SEL(n6), .F(n5) );
  XNOR U7 ( .A(n9), .B(n10), .Z(n6) );
  AND U8 ( .A(n11), .B(n12), .Z(n10) );
  XNOR U9 ( .A(n13), .B(n14), .Z(n12) );
  XOR U10 ( .A(n9), .B(n15), .Z(n14) );
  AND U11 ( .A(n4), .B(n16), .Z(n15) );
  XNOR U12 ( .A(n17), .B(n18), .Z(n16) );
  XNOR U13 ( .A(n19), .B(n20), .Z(n11) );
  XOR U14 ( .A(n9), .B(n21), .Z(n20) );
  AND U15 ( .A(n22), .B(n19), .Z(n21) );
  AND U16 ( .A(n23), .B(n24), .Z(n9) );
  XNOR U17 ( .A(n25), .B(n26), .Z(n24) );
  AND U18 ( .A(n4), .B(n27), .Z(n25) );
  XNOR U19 ( .A(n28), .B(n26), .Z(n27) );
  XOR U20 ( .A(n29), .B(n30), .Z(n4) );
  MUX U21 ( .IN0(n31), .IN1(n32), .SEL(n29), .F(n30) );
  XNOR U22 ( .A(n33), .B(n34), .Z(n29) );
  AND U23 ( .A(n35), .B(n36), .Z(n34) );
  XNOR U24 ( .A(n18), .B(n33), .Z(n36) );
  XNOR U25 ( .A(n33), .B(n17), .Z(n35) );
  IV U26 ( .A(n13), .Z(n17) );
  AND U27 ( .A(n26), .B(n28), .Z(n33) );
  XOR U28 ( .A(n37), .B(n38), .Z(n28) );
  XNOR U29 ( .A(n39), .B(n40), .Z(n26) );
  XOR U30 ( .A(n41), .B(n42), .Z(n23) );
  AND U31 ( .A(n2), .B(n43), .Z(n42) );
  XNOR U32 ( .A(n41), .B(n44), .Z(n43) );
  XOR U33 ( .A(n45), .B(n46), .Z(n2) );
  MUX U34 ( .IN0(n47), .IN1(n48), .SEL(n45), .F(n46) );
  XNOR U35 ( .A(n49), .B(n50), .Z(n45) );
  AND U36 ( .A(n51), .B(n52), .Z(n50) );
  XNOR U37 ( .A(n22), .B(n49), .Z(n52) );
  XNOR U38 ( .A(n49), .B(n19), .Z(n51) );
  AND U39 ( .A(n41), .B(n44), .Z(n49) );
  XOR U40 ( .A(n53), .B(n54), .Z(n44) );
  XNOR U41 ( .A(n55), .B(n56), .Z(n41) );
  AND U42 ( .A(n31), .B(n32), .Z(n8) );
  XOR U43 ( .A(n57), .B(n58), .Z(n32) );
  XOR U44 ( .A(n59), .B(n60), .Z(n58) );
  NOR U45 ( .A(n61), .B(n62), .Z(n60) );
  AND U46 ( .A(n63), .B(n64), .Z(n62) );
  NOR U47 ( .A(n63), .B(n65), .Z(n59) );
  XNOR U48 ( .A(n66), .B(n67), .Z(n57) );
  AND U49 ( .A(n18), .B(n68), .Z(n67) );
  XNOR U50 ( .A(n64), .B(n68), .Z(n18) );
  AND U51 ( .A(n38), .B(n37), .Z(n68) );
  XOR U52 ( .A(n69), .B(n70), .Z(n37) );
  AND U53 ( .A(p_input[15]), .B(p_input[14]), .Z(n38) );
  XOR U54 ( .A(n71), .B(n63), .Z(n64) );
  AND U55 ( .A(n70), .B(n69), .Z(n63) );
  XOR U56 ( .A(n72), .B(n73), .Z(n69) );
  AND U57 ( .A(p_input[13]), .B(p_input[12]), .Z(n70) );
  AND U58 ( .A(n74), .B(n75), .Z(n66) );
  IV U59 ( .A(n76), .Z(n75) );
  NOR U60 ( .A(n77), .B(n78), .Z(n76) );
  NOR U61 ( .A(n61), .B(n79), .Z(n74) );
  AND U62 ( .A(n65), .B(n71), .Z(n79) );
  XOR U63 ( .A(n80), .B(n77), .Z(n71) );
  XOR U64 ( .A(n78), .B(n81), .Z(n77) );
  AND U65 ( .A(n82), .B(n83), .Z(n81) );
  XNOR U66 ( .A(n84), .B(n85), .Z(n78) );
  NOR U67 ( .A(n86), .B(n87), .Z(n85) );
  AND U68 ( .A(n88), .B(n89), .Z(n87) );
  AND U69 ( .A(n90), .B(n91), .Z(n86) );
  XNOR U70 ( .A(n88), .B(n89), .Z(n84) );
  XNOR U71 ( .A(n61), .B(n65), .Z(n80) );
  AND U72 ( .A(n73), .B(n72), .Z(n65) );
  XOR U73 ( .A(n92), .B(n93), .Z(n72) );
  AND U74 ( .A(p_input[11]), .B(p_input[10]), .Z(n73) );
  AND U75 ( .A(n93), .B(n92), .Z(n61) );
  XOR U76 ( .A(n83), .B(n82), .Z(n92) );
  AND U77 ( .A(p_input[7]), .B(p_input[6]), .Z(n82) );
  XOR U78 ( .A(n90), .B(n91), .Z(n83) );
  XOR U79 ( .A(n88), .B(n89), .Z(n91) );
  AND U80 ( .A(p_input[3]), .B(p_input[2]), .Z(n89) );
  AND U81 ( .A(p_input[1]), .B(p_input[0]), .Z(n88) );
  AND U82 ( .A(p_input[5]), .B(p_input[4]), .Z(n90) );
  AND U83 ( .A(p_input[9]), .B(p_input[8]), .Z(n93) );
  XOR U84 ( .A(n94), .B(n95), .Z(n31) );
  XOR U85 ( .A(n96), .B(n97), .Z(n95) );
  NOR U86 ( .A(n98), .B(n99), .Z(n97) );
  AND U87 ( .A(n100), .B(n101), .Z(n99) );
  NOR U88 ( .A(n100), .B(n102), .Z(n96) );
  XNOR U89 ( .A(n103), .B(n104), .Z(n94) );
  AND U90 ( .A(n13), .B(n105), .Z(n104) );
  XNOR U91 ( .A(n101), .B(n105), .Z(n13) );
  AND U92 ( .A(n40), .B(n39), .Z(n105) );
  XOR U93 ( .A(n106), .B(n107), .Z(n39) );
  NOR U94 ( .A(n108), .B(p_input[14]), .Z(n40) );
  IV U95 ( .A(p_input[15]), .Z(n108) );
  XOR U96 ( .A(n109), .B(n100), .Z(n101) );
  AND U97 ( .A(n107), .B(n106), .Z(n100) );
  XOR U98 ( .A(n110), .B(n111), .Z(n106) );
  NOR U99 ( .A(n112), .B(p_input[12]), .Z(n107) );
  IV U100 ( .A(p_input[13]), .Z(n112) );
  AND U101 ( .A(n113), .B(n114), .Z(n103) );
  IV U102 ( .A(n115), .Z(n114) );
  NOR U103 ( .A(n116), .B(n117), .Z(n115) );
  NOR U104 ( .A(n98), .B(n118), .Z(n113) );
  AND U105 ( .A(n102), .B(n109), .Z(n118) );
  XOR U106 ( .A(n119), .B(n116), .Z(n109) );
  XOR U107 ( .A(n117), .B(n120), .Z(n116) );
  AND U108 ( .A(n121), .B(n122), .Z(n120) );
  XNOR U109 ( .A(n123), .B(n124), .Z(n117) );
  NOR U110 ( .A(n125), .B(n126), .Z(n124) );
  AND U111 ( .A(n127), .B(n128), .Z(n126) );
  AND U112 ( .A(n129), .B(n130), .Z(n125) );
  XNOR U113 ( .A(n127), .B(n128), .Z(n123) );
  XNOR U114 ( .A(n98), .B(n102), .Z(n119) );
  AND U115 ( .A(n111), .B(n110), .Z(n102) );
  XOR U116 ( .A(n131), .B(n132), .Z(n110) );
  NOR U117 ( .A(n133), .B(p_input[10]), .Z(n111) );
  IV U118 ( .A(p_input[11]), .Z(n133) );
  AND U119 ( .A(n132), .B(n131), .Z(n98) );
  XOR U120 ( .A(n122), .B(n121), .Z(n131) );
  NOR U121 ( .A(n134), .B(p_input[6]), .Z(n121) );
  IV U122 ( .A(p_input[7]), .Z(n134) );
  XOR U123 ( .A(n129), .B(n130), .Z(n122) );
  XOR U124 ( .A(n127), .B(n128), .Z(n130) );
  NOR U125 ( .A(n135), .B(p_input[2]), .Z(n128) );
  IV U126 ( .A(p_input[3]), .Z(n135) );
  NOR U127 ( .A(n136), .B(p_input[0]), .Z(n127) );
  IV U128 ( .A(p_input[1]), .Z(n136) );
  NOR U129 ( .A(n137), .B(p_input[4]), .Z(n129) );
  IV U130 ( .A(p_input[5]), .Z(n137) );
  NOR U131 ( .A(n138), .B(p_input[8]), .Z(n132) );
  IV U132 ( .A(p_input[9]), .Z(n138) );
  AND U133 ( .A(n47), .B(n48), .Z(n7) );
  XOR U134 ( .A(n139), .B(n140), .Z(n48) );
  XOR U135 ( .A(n141), .B(n142), .Z(n140) );
  NOR U136 ( .A(n143), .B(n144), .Z(n142) );
  AND U137 ( .A(n145), .B(n146), .Z(n144) );
  NOR U138 ( .A(n145), .B(n147), .Z(n141) );
  XNOR U139 ( .A(n148), .B(n149), .Z(n139) );
  AND U140 ( .A(n22), .B(n150), .Z(n149) );
  XNOR U141 ( .A(n146), .B(n150), .Z(n22) );
  AND U142 ( .A(n54), .B(n53), .Z(n150) );
  XOR U143 ( .A(n151), .B(n152), .Z(n53) );
  NOR U144 ( .A(n153), .B(p_input[15]), .Z(n54) );
  IV U145 ( .A(p_input[14]), .Z(n153) );
  XOR U146 ( .A(n154), .B(n145), .Z(n146) );
  AND U147 ( .A(n152), .B(n151), .Z(n145) );
  XOR U148 ( .A(n155), .B(n156), .Z(n151) );
  NOR U149 ( .A(n157), .B(p_input[13]), .Z(n152) );
  IV U150 ( .A(p_input[12]), .Z(n157) );
  AND U151 ( .A(n158), .B(n159), .Z(n148) );
  IV U152 ( .A(n160), .Z(n159) );
  NOR U153 ( .A(n161), .B(n162), .Z(n160) );
  NOR U154 ( .A(n143), .B(n163), .Z(n158) );
  AND U155 ( .A(n147), .B(n154), .Z(n163) );
  XOR U156 ( .A(n164), .B(n161), .Z(n154) );
  XOR U157 ( .A(n162), .B(n165), .Z(n161) );
  AND U158 ( .A(n166), .B(n167), .Z(n165) );
  XNOR U159 ( .A(n168), .B(n169), .Z(n162) );
  NOR U160 ( .A(n170), .B(n171), .Z(n169) );
  AND U161 ( .A(n172), .B(n173), .Z(n171) );
  AND U162 ( .A(n174), .B(n175), .Z(n170) );
  XNOR U163 ( .A(n172), .B(n173), .Z(n168) );
  XNOR U164 ( .A(n143), .B(n147), .Z(n164) );
  AND U165 ( .A(n156), .B(n155), .Z(n147) );
  XOR U166 ( .A(n176), .B(n177), .Z(n155) );
  NOR U167 ( .A(n178), .B(p_input[11]), .Z(n156) );
  IV U168 ( .A(p_input[10]), .Z(n178) );
  AND U169 ( .A(n177), .B(n176), .Z(n143) );
  XOR U170 ( .A(n167), .B(n166), .Z(n176) );
  NOR U171 ( .A(n179), .B(p_input[7]), .Z(n166) );
  IV U172 ( .A(p_input[6]), .Z(n179) );
  XOR U173 ( .A(n174), .B(n175), .Z(n167) );
  XOR U174 ( .A(n172), .B(n173), .Z(n175) );
  NOR U175 ( .A(n180), .B(p_input[3]), .Z(n173) );
  IV U176 ( .A(p_input[2]), .Z(n180) );
  NOR U177 ( .A(n181), .B(p_input[1]), .Z(n172) );
  IV U178 ( .A(p_input[0]), .Z(n181) );
  NOR U179 ( .A(n182), .B(p_input[5]), .Z(n174) );
  IV U180 ( .A(p_input[4]), .Z(n182) );
  NOR U181 ( .A(n183), .B(p_input[9]), .Z(n177) );
  IV U182 ( .A(p_input[8]), .Z(n183) );
  XOR U183 ( .A(n184), .B(n185), .Z(n47) );
  XOR U184 ( .A(n186), .B(n187), .Z(n185) );
  NOR U185 ( .A(n188), .B(n189), .Z(n187) );
  AND U186 ( .A(n190), .B(n191), .Z(n189) );
  NOR U187 ( .A(n190), .B(n192), .Z(n186) );
  XNOR U188 ( .A(n193), .B(n194), .Z(n184) );
  NOR U189 ( .A(n19), .B(n195), .Z(n194) );
  XNOR U190 ( .A(n191), .B(n195), .Z(n19) );
  IV U191 ( .A(n196), .Z(n195) );
  AND U192 ( .A(n56), .B(n55), .Z(n196) );
  XOR U193 ( .A(n197), .B(n198), .Z(n55) );
  NOR U194 ( .A(p_input[15]), .B(p_input[14]), .Z(n56) );
  XOR U195 ( .A(n199), .B(n190), .Z(n191) );
  AND U196 ( .A(n198), .B(n197), .Z(n190) );
  XOR U197 ( .A(n200), .B(n201), .Z(n197) );
  NOR U198 ( .A(p_input[13]), .B(p_input[12]), .Z(n198) );
  AND U199 ( .A(n202), .B(n203), .Z(n193) );
  IV U200 ( .A(n204), .Z(n203) );
  NOR U201 ( .A(n205), .B(n206), .Z(n204) );
  NOR U202 ( .A(n188), .B(n207), .Z(n202) );
  AND U203 ( .A(n192), .B(n199), .Z(n207) );
  XOR U204 ( .A(n208), .B(n205), .Z(n199) );
  XOR U205 ( .A(n206), .B(n209), .Z(n205) );
  AND U206 ( .A(n210), .B(n211), .Z(n209) );
  XNOR U207 ( .A(n212), .B(n213), .Z(n206) );
  NOR U208 ( .A(n214), .B(n215), .Z(n213) );
  AND U209 ( .A(n216), .B(n217), .Z(n215) );
  AND U210 ( .A(n218), .B(n219), .Z(n214) );
  XNOR U211 ( .A(n216), .B(n217), .Z(n212) );
  XNOR U212 ( .A(n188), .B(n192), .Z(n208) );
  AND U213 ( .A(n201), .B(n200), .Z(n192) );
  XOR U214 ( .A(n220), .B(n221), .Z(n200) );
  NOR U215 ( .A(p_input[11]), .B(p_input[10]), .Z(n201) );
  AND U216 ( .A(n221), .B(n220), .Z(n188) );
  XOR U217 ( .A(n211), .B(n210), .Z(n220) );
  NOR U218 ( .A(p_input[7]), .B(p_input[6]), .Z(n210) );
  XOR U219 ( .A(n218), .B(n219), .Z(n211) );
  XOR U220 ( .A(n216), .B(n217), .Z(n219) );
  NOR U221 ( .A(p_input[3]), .B(p_input[2]), .Z(n217) );
  NOR U222 ( .A(p_input[1]), .B(p_input[0]), .Z(n216) );
  NOR U223 ( .A(p_input[5]), .B(p_input[4]), .Z(n218) );
  NOR U224 ( .A(p_input[9]), .B(p_input[8]), .Z(n221) );
endmodule

