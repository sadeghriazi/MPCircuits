
module voting_N3_M4 ( p_input, o );
  input [47:0] p_input;
  output [2:0] o;
  wire   \one_vote[1].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[1].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[1].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[1].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[1].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[1].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[1].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[1].decoder_/sll_39/ML_int[2][3] ,
         \one_vote[2].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[2].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[2].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[2].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[2].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[2].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[2].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[2].decoder_/sll_39/ML_int[2][3] ,
         \one_vote[3].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[3].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[3].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[3].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[3].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[3].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[3].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[3].decoder_/sll_39/ML_int[2][3] ,
         \one_vote[4].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[4].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[4].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[4].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[4].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[4].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[4].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[4].decoder_/sll_39/ML_int[2][3] ,
         \one_vote[5].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[5].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[5].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[5].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[5].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[5].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[5].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[5].decoder_/sll_39/ML_int[2][3] ,
         \one_vote[6].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[6].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[6].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[6].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[6].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[6].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[6].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[6].decoder_/sll_39/ML_int[2][3] ,
         \one_vote[7].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[7].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[7].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[7].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[7].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[7].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[7].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[7].decoder_/sll_39/ML_int[2][3] ,
         \one_vote[8].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[8].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[8].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[8].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[8].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[8].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[8].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[8].decoder_/sll_39/ML_int[2][3] ,
         \one_vote[9].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[9].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[9].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[9].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[9].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[9].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[9].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[9].decoder_/sll_39/ML_int[2][3] ,
         \one_vote[10].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[10].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[10].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[10].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[10].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[10].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[10].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[10].decoder_/sll_39/ML_int[2][3] ,
         \one_vote[11].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[11].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[11].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[11].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[11].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[11].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[11].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[11].decoder_/sll_39/ML_int[2][3] ,
         \one_vote[12].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[12].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[12].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[12].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[12].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[12].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[12].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[12].decoder_/sll_39/ML_int[2][3] ,
         \one_vote[13].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[13].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[13].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[13].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[13].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[13].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[13].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[13].decoder_/sll_39/ML_int[2][3] ,
         \one_vote[14].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[14].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[14].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[14].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[14].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[14].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[14].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[14].decoder_/sll_39/ML_int[2][3] ,
         \one_vote[15].decoder_/sll_39/ML_int[3][4] ,
         \one_vote[15].decoder_/sll_39/ML_int[3][5] ,
         \one_vote[15].decoder_/sll_39/ML_int[3][6] ,
         \one_vote[15].decoder_/sll_39/ML_int[3][7] ,
         \one_vote[15].decoder_/sll_39/ML_int[2][0] ,
         \one_vote[15].decoder_/sll_39/ML_int[2][1] ,
         \one_vote[15].decoder_/sll_39/ML_int[2][2] ,
         \one_vote[15].decoder_/sll_39/ML_int[2][3] ,
         \decoder_/sll_39/ML_int[3][4] , \decoder_/sll_39/ML_int[3][5] ,
         \decoder_/sll_39/ML_int[3][6] , \decoder_/sll_39/ML_int[3][7] ,
         \decoder_/sll_39/ML_int[2][0] , \decoder_/sll_39/ML_int[2][1] ,
         \decoder_/sll_39/ML_int[2][2] , \decoder_/sll_39/ML_int[2][3] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;

  AND U2 ( .A(p_input[4]), .B(n1020), .Z(
        \one_vote[1].decoder_/sll_39/ML_int[2][2] ) );
  AND U3 ( .A(p_input[4]), .B(p_input[3]), .Z(
        \one_vote[1].decoder_/sll_39/ML_int[2][3] ) );
  AND U4 ( .A(p_input[7]), .B(n1019), .Z(
        \one_vote[2].decoder_/sll_39/ML_int[2][2] ) );
  AND U5 ( .A(p_input[7]), .B(p_input[6]), .Z(
        \one_vote[2].decoder_/sll_39/ML_int[2][3] ) );
  AND U6 ( .A(p_input[10]), .B(n1018), .Z(
        \one_vote[3].decoder_/sll_39/ML_int[2][2] ) );
  AND U7 ( .A(p_input[10]), .B(p_input[9]), .Z(
        \one_vote[3].decoder_/sll_39/ML_int[2][3] ) );
  AND U8 ( .A(p_input[13]), .B(n1017), .Z(
        \one_vote[4].decoder_/sll_39/ML_int[2][2] ) );
  AND U9 ( .A(p_input[13]), .B(p_input[12]), .Z(
        \one_vote[4].decoder_/sll_39/ML_int[2][3] ) );
  AND U10 ( .A(p_input[16]), .B(n1016), .Z(
        \one_vote[5].decoder_/sll_39/ML_int[2][2] ) );
  AND U11 ( .A(p_input[16]), .B(p_input[15]), .Z(
        \one_vote[5].decoder_/sll_39/ML_int[2][3] ) );
  AND U12 ( .A(p_input[19]), .B(n1015), .Z(
        \one_vote[6].decoder_/sll_39/ML_int[2][2] ) );
  AND U13 ( .A(p_input[19]), .B(p_input[18]), .Z(
        \one_vote[6].decoder_/sll_39/ML_int[2][3] ) );
  AND U14 ( .A(p_input[22]), .B(n1014), .Z(
        \one_vote[7].decoder_/sll_39/ML_int[2][2] ) );
  AND U15 ( .A(p_input[22]), .B(p_input[21]), .Z(
        \one_vote[7].decoder_/sll_39/ML_int[2][3] ) );
  AND U16 ( .A(p_input[25]), .B(n1013), .Z(
        \one_vote[8].decoder_/sll_39/ML_int[2][2] ) );
  AND U17 ( .A(p_input[25]), .B(p_input[24]), .Z(
        \one_vote[8].decoder_/sll_39/ML_int[2][3] ) );
  AND U18 ( .A(p_input[28]), .B(n1012), .Z(
        \one_vote[9].decoder_/sll_39/ML_int[2][2] ) );
  AND U19 ( .A(p_input[28]), .B(p_input[27]), .Z(
        \one_vote[9].decoder_/sll_39/ML_int[2][3] ) );
  AND U20 ( .A(p_input[31]), .B(n1011), .Z(
        \one_vote[10].decoder_/sll_39/ML_int[2][2] ) );
  AND U21 ( .A(p_input[31]), .B(p_input[30]), .Z(
        \one_vote[10].decoder_/sll_39/ML_int[2][3] ) );
  AND U22 ( .A(p_input[34]), .B(n1010), .Z(
        \one_vote[11].decoder_/sll_39/ML_int[2][2] ) );
  AND U23 ( .A(p_input[34]), .B(p_input[33]), .Z(
        \one_vote[11].decoder_/sll_39/ML_int[2][3] ) );
  AND U24 ( .A(p_input[37]), .B(n1009), .Z(
        \one_vote[12].decoder_/sll_39/ML_int[2][2] ) );
  AND U25 ( .A(p_input[37]), .B(p_input[36]), .Z(
        \one_vote[12].decoder_/sll_39/ML_int[2][3] ) );
  AND U26 ( .A(p_input[40]), .B(n1008), .Z(
        \one_vote[13].decoder_/sll_39/ML_int[2][2] ) );
  AND U27 ( .A(p_input[40]), .B(p_input[39]), .Z(
        \one_vote[13].decoder_/sll_39/ML_int[2][3] ) );
  AND U28 ( .A(p_input[43]), .B(n1007), .Z(
        \one_vote[14].decoder_/sll_39/ML_int[2][2] ) );
  AND U29 ( .A(p_input[43]), .B(p_input[42]), .Z(
        \one_vote[14].decoder_/sll_39/ML_int[2][3] ) );
  AND U30 ( .A(p_input[46]), .B(n1006), .Z(
        \one_vote[15].decoder_/sll_39/ML_int[2][2] ) );
  AND U31 ( .A(p_input[46]), .B(p_input[45]), .Z(
        \one_vote[15].decoder_/sll_39/ML_int[2][3] ) );
  AND U32 ( .A(p_input[1]), .B(n1021), .Z(\decoder_/sll_39/ML_int[2][2] ) );
  AND U33 ( .A(p_input[1]), .B(p_input[0]), .Z(\decoder_/sll_39/ML_int[2][3] )
         );
  AND U34 ( .A(p_input[2]), .B(\decoder_/sll_39/ML_int[2][0] ), .Z(
        \decoder_/sll_39/ML_int[3][4] ) );
  AND U35 ( .A(p_input[2]), .B(\decoder_/sll_39/ML_int[2][1] ), .Z(
        \decoder_/sll_39/ML_int[3][5] ) );
  AND U36 ( .A(p_input[2]), .B(\decoder_/sll_39/ML_int[2][2] ), .Z(
        \decoder_/sll_39/ML_int[3][6] ) );
  AND U37 ( .A(p_input[2]), .B(\decoder_/sll_39/ML_int[2][3] ), .Z(
        \decoder_/sll_39/ML_int[3][7] ) );
  AND U38 ( .A(p_input[5]), .B(\one_vote[1].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[1].decoder_/sll_39/ML_int[3][4] ) );
  AND U39 ( .A(p_input[5]), .B(\one_vote[1].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[1].decoder_/sll_39/ML_int[3][5] ) );
  AND U40 ( .A(p_input[5]), .B(\one_vote[1].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[1].decoder_/sll_39/ML_int[3][6] ) );
  AND U41 ( .A(p_input[5]), .B(\one_vote[1].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[1].decoder_/sll_39/ML_int[3][7] ) );
  AND U42 ( .A(p_input[8]), .B(\one_vote[2].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[2].decoder_/sll_39/ML_int[3][4] ) );
  AND U43 ( .A(p_input[8]), .B(\one_vote[2].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[2].decoder_/sll_39/ML_int[3][5] ) );
  AND U44 ( .A(p_input[8]), .B(\one_vote[2].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[2].decoder_/sll_39/ML_int[3][6] ) );
  AND U45 ( .A(p_input[8]), .B(\one_vote[2].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[2].decoder_/sll_39/ML_int[3][7] ) );
  AND U46 ( .A(p_input[11]), .B(\one_vote[3].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[3].decoder_/sll_39/ML_int[3][4] ) );
  AND U47 ( .A(p_input[11]), .B(\one_vote[3].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[3].decoder_/sll_39/ML_int[3][5] ) );
  AND U48 ( .A(p_input[11]), .B(\one_vote[3].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[3].decoder_/sll_39/ML_int[3][6] ) );
  AND U49 ( .A(p_input[11]), .B(\one_vote[3].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[3].decoder_/sll_39/ML_int[3][7] ) );
  AND U50 ( .A(p_input[14]), .B(\one_vote[4].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[4].decoder_/sll_39/ML_int[3][4] ) );
  AND U51 ( .A(p_input[14]), .B(\one_vote[4].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[4].decoder_/sll_39/ML_int[3][5] ) );
  AND U52 ( .A(p_input[14]), .B(\one_vote[4].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[4].decoder_/sll_39/ML_int[3][6] ) );
  AND U53 ( .A(p_input[14]), .B(\one_vote[4].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[4].decoder_/sll_39/ML_int[3][7] ) );
  AND U54 ( .A(p_input[17]), .B(\one_vote[5].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[5].decoder_/sll_39/ML_int[3][4] ) );
  AND U55 ( .A(p_input[17]), .B(\one_vote[5].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[5].decoder_/sll_39/ML_int[3][5] ) );
  AND U56 ( .A(p_input[17]), .B(\one_vote[5].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[5].decoder_/sll_39/ML_int[3][6] ) );
  AND U57 ( .A(p_input[17]), .B(\one_vote[5].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[5].decoder_/sll_39/ML_int[3][7] ) );
  AND U58 ( .A(p_input[20]), .B(\one_vote[6].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[6].decoder_/sll_39/ML_int[3][4] ) );
  AND U59 ( .A(p_input[20]), .B(\one_vote[6].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[6].decoder_/sll_39/ML_int[3][5] ) );
  AND U60 ( .A(p_input[20]), .B(\one_vote[6].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[6].decoder_/sll_39/ML_int[3][6] ) );
  AND U61 ( .A(p_input[20]), .B(\one_vote[6].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[6].decoder_/sll_39/ML_int[3][7] ) );
  AND U62 ( .A(p_input[23]), .B(\one_vote[7].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[7].decoder_/sll_39/ML_int[3][4] ) );
  AND U63 ( .A(p_input[23]), .B(\one_vote[7].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[7].decoder_/sll_39/ML_int[3][5] ) );
  AND U64 ( .A(p_input[23]), .B(\one_vote[7].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[7].decoder_/sll_39/ML_int[3][6] ) );
  AND U65 ( .A(p_input[23]), .B(\one_vote[7].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[7].decoder_/sll_39/ML_int[3][7] ) );
  AND U66 ( .A(p_input[26]), .B(\one_vote[8].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[8].decoder_/sll_39/ML_int[3][4] ) );
  AND U67 ( .A(p_input[26]), .B(\one_vote[8].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[8].decoder_/sll_39/ML_int[3][5] ) );
  AND U68 ( .A(p_input[26]), .B(\one_vote[8].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[8].decoder_/sll_39/ML_int[3][6] ) );
  AND U69 ( .A(p_input[26]), .B(\one_vote[8].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[8].decoder_/sll_39/ML_int[3][7] ) );
  AND U70 ( .A(p_input[29]), .B(\one_vote[9].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[9].decoder_/sll_39/ML_int[3][4] ) );
  AND U71 ( .A(p_input[29]), .B(\one_vote[9].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[9].decoder_/sll_39/ML_int[3][5] ) );
  AND U72 ( .A(p_input[29]), .B(\one_vote[9].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[9].decoder_/sll_39/ML_int[3][6] ) );
  AND U73 ( .A(p_input[29]), .B(\one_vote[9].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[9].decoder_/sll_39/ML_int[3][7] ) );
  AND U74 ( .A(p_input[32]), .B(\one_vote[10].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[10].decoder_/sll_39/ML_int[3][4] ) );
  AND U75 ( .A(p_input[32]), .B(\one_vote[10].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[10].decoder_/sll_39/ML_int[3][5] ) );
  AND U76 ( .A(p_input[32]), .B(\one_vote[10].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[10].decoder_/sll_39/ML_int[3][6] ) );
  AND U77 ( .A(p_input[32]), .B(\one_vote[10].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[10].decoder_/sll_39/ML_int[3][7] ) );
  AND U78 ( .A(p_input[35]), .B(\one_vote[11].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[11].decoder_/sll_39/ML_int[3][4] ) );
  AND U79 ( .A(p_input[35]), .B(\one_vote[11].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[11].decoder_/sll_39/ML_int[3][5] ) );
  AND U80 ( .A(p_input[35]), .B(\one_vote[11].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[11].decoder_/sll_39/ML_int[3][6] ) );
  AND U81 ( .A(p_input[35]), .B(\one_vote[11].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[11].decoder_/sll_39/ML_int[3][7] ) );
  AND U82 ( .A(p_input[38]), .B(\one_vote[12].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[12].decoder_/sll_39/ML_int[3][4] ) );
  AND U83 ( .A(p_input[38]), .B(\one_vote[12].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[12].decoder_/sll_39/ML_int[3][5] ) );
  AND U84 ( .A(p_input[38]), .B(\one_vote[12].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[12].decoder_/sll_39/ML_int[3][6] ) );
  AND U85 ( .A(p_input[38]), .B(\one_vote[12].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[12].decoder_/sll_39/ML_int[3][7] ) );
  AND U86 ( .A(p_input[41]), .B(\one_vote[13].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[13].decoder_/sll_39/ML_int[3][4] ) );
  AND U87 ( .A(p_input[41]), .B(\one_vote[13].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[13].decoder_/sll_39/ML_int[3][5] ) );
  AND U88 ( .A(p_input[41]), .B(\one_vote[13].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[13].decoder_/sll_39/ML_int[3][6] ) );
  AND U89 ( .A(p_input[41]), .B(\one_vote[13].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[13].decoder_/sll_39/ML_int[3][7] ) );
  AND U90 ( .A(p_input[44]), .B(\one_vote[14].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[14].decoder_/sll_39/ML_int[3][4] ) );
  AND U91 ( .A(p_input[44]), .B(\one_vote[14].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[14].decoder_/sll_39/ML_int[3][5] ) );
  AND U92 ( .A(p_input[44]), .B(\one_vote[14].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[14].decoder_/sll_39/ML_int[3][6] ) );
  AND U93 ( .A(p_input[44]), .B(\one_vote[14].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[14].decoder_/sll_39/ML_int[3][7] ) );
  AND U94 ( .A(p_input[47]), .B(\one_vote[15].decoder_/sll_39/ML_int[2][0] ), 
        .Z(\one_vote[15].decoder_/sll_39/ML_int[3][4] ) );
  AND U95 ( .A(p_input[47]), .B(\one_vote[15].decoder_/sll_39/ML_int[2][1] ), 
        .Z(\one_vote[15].decoder_/sll_39/ML_int[3][5] ) );
  AND U96 ( .A(p_input[47]), .B(\one_vote[15].decoder_/sll_39/ML_int[2][2] ), 
        .Z(\one_vote[15].decoder_/sll_39/ML_int[3][6] ) );
  AND U97 ( .A(p_input[47]), .B(\one_vote[15].decoder_/sll_39/ML_int[2][3] ), 
        .Z(\one_vote[15].decoder_/sll_39/ML_int[3][7] ) );
  XNOR U98 ( .A(n1), .B(n2), .Z(o[0]) );
  AND U99 ( .A(o[1]), .B(n3), .Z(n2) );
  XOR U100 ( .A(n4), .B(n1), .Z(n3) );
  XNOR U101 ( .A(n5), .B(n6), .Z(n4) );
  AND U102 ( .A(o[2]), .B(n7), .Z(n6) );
  XOR U103 ( .A(n8), .B(n5), .Z(n7) );
  XOR U104 ( .A(n9), .B(n10), .Z(o[1]) );
  AND U105 ( .A(o[2]), .B(n11), .Z(n10) );
  XOR U106 ( .A(n12), .B(n9), .Z(n11) );
  XNOR U107 ( .A(n13), .B(n14), .Z(n1) );
  AND U108 ( .A(o[2]), .B(n15), .Z(n14) );
  XOR U109 ( .A(n13), .B(n16), .Z(n15) );
  NOR U110 ( .A(n17), .B(n18), .Z(o[2]) );
  XOR U111 ( .A(n19), .B(n20), .Z(n18) );
  AND U112 ( .A(n21), .B(n22), .Z(n19) );
  XOR U113 ( .A(n23), .B(n20), .Z(n22) );
  AND U114 ( .A(n24), .B(n25), .Z(n23) );
  XNOR U115 ( .A(n20), .B(n26), .Z(n21) );
  AND U116 ( .A(n27), .B(n28), .Z(n26) );
  XOR U117 ( .A(n29), .B(n30), .Z(n20) );
  AND U118 ( .A(n31), .B(n32), .Z(n30) );
  XOR U119 ( .A(n29), .B(n33), .Z(n32) );
  XOR U120 ( .A(n34), .B(n35), .Z(n33) );
  AND U121 ( .A(n12), .B(n36), .Z(n34) );
  XOR U122 ( .A(n37), .B(n35), .Z(n36) );
  XOR U123 ( .A(n38), .B(n29), .Z(n31) );
  XNOR U124 ( .A(n39), .B(n40), .Z(n38) );
  AND U125 ( .A(n9), .B(n41), .Z(n40) );
  XOR U126 ( .A(n42), .B(n39), .Z(n41) );
  XOR U127 ( .A(n43), .B(n44), .Z(n29) );
  AND U128 ( .A(n45), .B(n46), .Z(n44) );
  XNOR U129 ( .A(n47), .B(n48), .Z(n46) );
  XOR U130 ( .A(n43), .B(n49), .Z(n48) );
  AND U131 ( .A(n12), .B(n50), .Z(n49) );
  XOR U132 ( .A(n47), .B(n51), .Z(n50) );
  XOR U133 ( .A(n52), .B(n53), .Z(n45) );
  XOR U134 ( .A(n43), .B(n54), .Z(n53) );
  AND U135 ( .A(n9), .B(n55), .Z(n54) );
  XOR U136 ( .A(n56), .B(n52), .Z(n55) );
  AND U137 ( .A(n57), .B(n58), .Z(n43) );
  XOR U138 ( .A(n59), .B(n60), .Z(n58) );
  AND U139 ( .A(n12), .B(n61), .Z(n59) );
  XNOR U140 ( .A(n62), .B(n60), .Z(n61) );
  NOR U141 ( .A(n63), .B(n64), .Z(n12) );
  XOR U142 ( .A(n65), .B(n66), .Z(n64) );
  AND U143 ( .A(n67), .B(n68), .Z(n65) );
  XOR U144 ( .A(n25), .B(n66), .Z(n68) );
  NOR U145 ( .A(n69), .B(n70), .Z(n25) );
  XNOR U146 ( .A(n66), .B(n24), .Z(n67) );
  NOR U147 ( .A(n71), .B(n72), .Z(n24) );
  XOR U148 ( .A(n73), .B(n74), .Z(n66) );
  AND U149 ( .A(n75), .B(n76), .Z(n74) );
  XOR U150 ( .A(n73), .B(n37), .Z(n76) );
  XNOR U151 ( .A(n77), .B(n78), .Z(n37) );
  AND U152 ( .A(n8), .B(n79), .Z(n78) );
  XOR U153 ( .A(n77), .B(n80), .Z(n79) );
  XNOR U154 ( .A(n35), .B(n73), .Z(n75) );
  XNOR U155 ( .A(n81), .B(n82), .Z(n35) );
  AND U156 ( .A(n5), .B(n83), .Z(n82) );
  XOR U157 ( .A(n81), .B(n84), .Z(n83) );
  XOR U158 ( .A(n85), .B(n86), .Z(n73) );
  AND U159 ( .A(n87), .B(n88), .Z(n86) );
  XNOR U160 ( .A(n51), .B(n85), .Z(n88) );
  XOR U161 ( .A(n89), .B(n90), .Z(n51) );
  AND U162 ( .A(n8), .B(n91), .Z(n90) );
  XOR U163 ( .A(n89), .B(n92), .Z(n91) );
  XOR U164 ( .A(n85), .B(n47), .Z(n87) );
  XOR U165 ( .A(n93), .B(n94), .Z(n47) );
  AND U166 ( .A(n5), .B(n95), .Z(n94) );
  XOR U167 ( .A(n93), .B(n96), .Z(n95) );
  NOR U168 ( .A(n60), .B(n62), .Z(n85) );
  XNOR U169 ( .A(n97), .B(n98), .Z(n62) );
  AND U170 ( .A(n8), .B(n99), .Z(n98) );
  XNOR U171 ( .A(n100), .B(n97), .Z(n99) );
  NOR U172 ( .A(n101), .B(n102), .Z(n8) );
  XOR U173 ( .A(n103), .B(n104), .Z(n102) );
  AND U174 ( .A(n105), .B(n106), .Z(n103) );
  XNOR U175 ( .A(n104), .B(n70), .Z(n106) );
  XOR U176 ( .A(n107), .B(n108), .Z(n70) );
  XOR U177 ( .A(n69), .B(n104), .Z(n105) );
  XOR U178 ( .A(n109), .B(n110), .Z(n104) );
  AND U179 ( .A(n111), .B(n112), .Z(n110) );
  XNOR U180 ( .A(n80), .B(n109), .Z(n112) );
  XOR U181 ( .A(n109), .B(n77), .Z(n111) );
  XOR U182 ( .A(n113), .B(n114), .Z(n109) );
  AND U183 ( .A(n115), .B(n116), .Z(n114) );
  XNOR U184 ( .A(n92), .B(n113), .Z(n116) );
  XOR U185 ( .A(n113), .B(n89), .Z(n115) );
  NOR U186 ( .A(n97), .B(n100), .Z(n113) );
  XNOR U187 ( .A(n117), .B(\one_vote[15].decoder_/sll_39/ML_int[3][7] ), .Z(
        n100) );
  XOR U188 ( .A(n118), .B(n119), .Z(n69) );
  NOR U189 ( .A(n120), .B(n121), .Z(n101) );
  IV U190 ( .A(n122), .Z(n120) );
  XOR U191 ( .A(n123), .B(\one_vote[15].decoder_/sll_39/ML_int[3][6] ), .Z(n97) );
  XOR U192 ( .A(n124), .B(n125), .Z(n60) );
  AND U193 ( .A(n5), .B(n126), .Z(n125) );
  XNOR U194 ( .A(n127), .B(n124), .Z(n126) );
  NOR U195 ( .A(n128), .B(n129), .Z(n5) );
  XOR U196 ( .A(n130), .B(n131), .Z(n129) );
  AND U197 ( .A(n132), .B(n133), .Z(n130) );
  XNOR U198 ( .A(n131), .B(n72), .Z(n133) );
  XOR U199 ( .A(n134), .B(n135), .Z(n72) );
  XOR U200 ( .A(n71), .B(n131), .Z(n132) );
  XOR U201 ( .A(n136), .B(n137), .Z(n131) );
  AND U202 ( .A(n138), .B(n139), .Z(n137) );
  XNOR U203 ( .A(n84), .B(n136), .Z(n139) );
  XOR U204 ( .A(n136), .B(n81), .Z(n138) );
  XOR U205 ( .A(n140), .B(n141), .Z(n136) );
  AND U206 ( .A(n142), .B(n143), .Z(n141) );
  XNOR U207 ( .A(n96), .B(n140), .Z(n143) );
  XOR U208 ( .A(n140), .B(n93), .Z(n142) );
  NOR U209 ( .A(n124), .B(n127), .Z(n140) );
  XNOR U210 ( .A(n144), .B(\one_vote[15].decoder_/sll_39/ML_int[3][5] ), .Z(
        n127) );
  XOR U211 ( .A(n145), .B(n146), .Z(n71) );
  NOR U212 ( .A(n147), .B(n148), .Z(n128) );
  IV U213 ( .A(n149), .Z(n147) );
  XOR U214 ( .A(n150), .B(\one_vote[15].decoder_/sll_39/ML_int[3][4] ), .Z(
        n124) );
  AND U215 ( .A(n151), .B(n152), .Z(n63) );
  XOR U216 ( .A(n153), .B(n154), .Z(n57) );
  AND U217 ( .A(n9), .B(n155), .Z(n154) );
  XNOR U218 ( .A(n153), .B(n156), .Z(n155) );
  NOR U219 ( .A(n157), .B(n158), .Z(n9) );
  XOR U220 ( .A(n159), .B(n160), .Z(n158) );
  AND U221 ( .A(n161), .B(n162), .Z(n159) );
  XOR U222 ( .A(n28), .B(n160), .Z(n162) );
  NOR U223 ( .A(n163), .B(n164), .Z(n28) );
  XNOR U224 ( .A(n160), .B(n27), .Z(n161) );
  AND U225 ( .A(n165), .B(n166), .Z(n27) );
  XOR U226 ( .A(n167), .B(n168), .Z(n160) );
  AND U227 ( .A(n169), .B(n170), .Z(n168) );
  XOR U228 ( .A(n167), .B(n42), .Z(n170) );
  XNOR U229 ( .A(n171), .B(n172), .Z(n42) );
  AND U230 ( .A(n16), .B(n173), .Z(n172) );
  XOR U231 ( .A(n171), .B(n174), .Z(n173) );
  XNOR U232 ( .A(n39), .B(n167), .Z(n169) );
  XNOR U233 ( .A(n175), .B(n176), .Z(n39) );
  AND U234 ( .A(n13), .B(n177), .Z(n176) );
  XOR U235 ( .A(n178), .B(n175), .Z(n177) );
  XOR U236 ( .A(n179), .B(n180), .Z(n167) );
  AND U237 ( .A(n181), .B(n182), .Z(n180) );
  XNOR U238 ( .A(n56), .B(n179), .Z(n182) );
  XOR U239 ( .A(n183), .B(n184), .Z(n56) );
  AND U240 ( .A(n16), .B(n185), .Z(n184) );
  XOR U241 ( .A(n183), .B(n186), .Z(n185) );
  XOR U242 ( .A(n179), .B(n52), .Z(n181) );
  XOR U243 ( .A(n187), .B(n188), .Z(n52) );
  AND U244 ( .A(n13), .B(n189), .Z(n188) );
  XOR U245 ( .A(n190), .B(n187), .Z(n189) );
  AND U246 ( .A(n153), .B(n156), .Z(n179) );
  XOR U247 ( .A(n191), .B(n192), .Z(n156) );
  AND U248 ( .A(n16), .B(n193), .Z(n192) );
  XNOR U249 ( .A(n191), .B(n194), .Z(n193) );
  NOR U250 ( .A(n195), .B(n196), .Z(n16) );
  XOR U251 ( .A(n197), .B(n198), .Z(n196) );
  AND U252 ( .A(n199), .B(n200), .Z(n197) );
  XNOR U253 ( .A(n198), .B(n164), .Z(n200) );
  XOR U254 ( .A(n201), .B(n202), .Z(n164) );
  XOR U255 ( .A(n163), .B(n198), .Z(n199) );
  XOR U256 ( .A(n203), .B(n204), .Z(n198) );
  AND U257 ( .A(n205), .B(n206), .Z(n204) );
  XNOR U258 ( .A(n174), .B(n203), .Z(n206) );
  XOR U259 ( .A(n203), .B(n171), .Z(n205) );
  XOR U260 ( .A(n207), .B(n208), .Z(n203) );
  AND U261 ( .A(n209), .B(n210), .Z(n208) );
  XNOR U262 ( .A(n186), .B(n207), .Z(n210) );
  XOR U263 ( .A(n207), .B(n183), .Z(n209) );
  NOR U264 ( .A(n191), .B(n194), .Z(n207) );
  XNOR U265 ( .A(n211), .B(n212), .Z(n194) );
  XOR U266 ( .A(n213), .B(n214), .Z(n163) );
  NOR U267 ( .A(n215), .B(n216), .Z(n195) );
  IV U268 ( .A(n217), .Z(n215) );
  XOR U269 ( .A(n218), .B(n219), .Z(n191) );
  NOR U270 ( .A(n220), .B(n221), .Z(n157) );
  IV U271 ( .A(n222), .Z(n220) );
  XNOR U272 ( .A(n223), .B(n224), .Z(n153) );
  AND U273 ( .A(n13), .B(n225), .Z(n224) );
  XNOR U274 ( .A(n223), .B(n226), .Z(n225) );
  AND U275 ( .A(n227), .B(n151), .Z(n17) );
  AND U276 ( .A(n122), .B(n121), .Z(n151) );
  NOR U277 ( .A(n119), .B(n118), .Z(n121) );
  XOR U278 ( .A(n228), .B(n229), .Z(n118) );
  XOR U279 ( .A(n230), .B(n231), .Z(n229) );
  NOR U280 ( .A(n232), .B(n233), .Z(n231) );
  NOR U281 ( .A(n234), .B(n235), .Z(n230) );
  AND U282 ( .A(n236), .B(n237), .Z(n235) );
  IV U283 ( .A(n238), .Z(n234) );
  NOR U284 ( .A(n239), .B(n240), .Z(n238) );
  AND U285 ( .A(n232), .B(n241), .Z(n240) );
  AND U286 ( .A(n233), .B(n242), .Z(n239) );
  XNOR U287 ( .A(n243), .B(n244), .Z(n228) );
  AND U288 ( .A(n245), .B(n246), .Z(n244) );
  AND U289 ( .A(n247), .B(n248), .Z(n243) );
  AND U290 ( .A(n249), .B(n250), .Z(n248) );
  IV U291 ( .A(n251), .Z(n250) );
  NOR U292 ( .A(n252), .B(n253), .Z(n249) );
  NOR U293 ( .A(n254), .B(n255), .Z(n247) );
  AND U294 ( .A(n77), .B(n256), .Z(n119) );
  XOR U295 ( .A(n245), .B(n256), .Z(n77) );
  AND U296 ( .A(n89), .B(n257), .Z(n256) );
  XOR U297 ( .A(n258), .B(n257), .Z(n89) );
  AND U298 ( .A(\one_vote[15].decoder_/sll_39/ML_int[3][6] ), .B(n123), .Z(
        n257) );
  XOR U299 ( .A(n259), .B(\one_vote[14].decoder_/sll_39/ML_int[3][6] ), .Z(
        n123) );
  XNOR U300 ( .A(n242), .B(n246), .Z(n245) );
  AND U301 ( .A(n258), .B(n260), .Z(n246) );
  XOR U302 ( .A(n261), .B(n260), .Z(n258) );
  AND U303 ( .A(\one_vote[14].decoder_/sll_39/ML_int[3][6] ), .B(n259), .Z(
        n260) );
  XOR U304 ( .A(n262), .B(\one_vote[13].decoder_/sll_39/ML_int[3][6] ), .Z(
        n259) );
  XOR U305 ( .A(n241), .B(n233), .Z(n242) );
  AND U306 ( .A(n261), .B(n263), .Z(n233) );
  XOR U307 ( .A(n264), .B(n263), .Z(n261) );
  AND U308 ( .A(\one_vote[13].decoder_/sll_39/ML_int[3][6] ), .B(n262), .Z(
        n263) );
  XOR U309 ( .A(n265), .B(\one_vote[12].decoder_/sll_39/ML_int[3][6] ), .Z(
        n262) );
  XNOR U310 ( .A(n236), .B(n232), .Z(n241) );
  AND U311 ( .A(n264), .B(n266), .Z(n232) );
  XOR U312 ( .A(n267), .B(n266), .Z(n264) );
  AND U313 ( .A(\one_vote[12].decoder_/sll_39/ML_int[3][6] ), .B(n265), .Z(
        n266) );
  XOR U314 ( .A(n268), .B(\one_vote[11].decoder_/sll_39/ML_int[3][6] ), .Z(
        n265) );
  XOR U315 ( .A(n269), .B(n270), .Z(n236) );
  XOR U316 ( .A(n254), .B(n271), .Z(n270) );
  XOR U317 ( .A(n252), .B(n251), .Z(n271) );
  AND U318 ( .A(n272), .B(n273), .Z(n251) );
  AND U319 ( .A(n274), .B(n275), .Z(n252) );
  AND U320 ( .A(n276), .B(n277), .Z(n254) );
  XNOR U321 ( .A(n278), .B(n253), .Z(n269) );
  XOR U322 ( .A(n279), .B(n280), .Z(n253) );
  XOR U323 ( .A(n281), .B(n282), .Z(n280) );
  AND U324 ( .A(n283), .B(n284), .Z(n282) );
  XNOR U325 ( .A(n285), .B(n286), .Z(n279) );
  NOR U326 ( .A(n287), .B(n288), .Z(n286) );
  AND U327 ( .A(n289), .B(n290), .Z(n288) );
  IV U328 ( .A(n291), .Z(n287) );
  NOR U329 ( .A(n281), .B(n292), .Z(n291) );
  AND U330 ( .A(n293), .B(n294), .Z(n292) );
  NOR U331 ( .A(n283), .B(n293), .Z(n285) );
  XNOR U332 ( .A(n255), .B(n237), .Z(n278) );
  AND U333 ( .A(n267), .B(n295), .Z(n237) );
  XOR U334 ( .A(n296), .B(n295), .Z(n267) );
  AND U335 ( .A(\one_vote[11].decoder_/sll_39/ML_int[3][6] ), .B(n268), .Z(
        n295) );
  XOR U336 ( .A(n297), .B(\one_vote[10].decoder_/sll_39/ML_int[3][6] ), .Z(
        n268) );
  AND U337 ( .A(n296), .B(n298), .Z(n255) );
  XOR U338 ( .A(n276), .B(n298), .Z(n296) );
  AND U339 ( .A(\one_vote[10].decoder_/sll_39/ML_int[3][6] ), .B(n297), .Z(
        n298) );
  XOR U340 ( .A(n299), .B(\one_vote[9].decoder_/sll_39/ML_int[3][6] ), .Z(n297) );
  XOR U341 ( .A(n272), .B(n277), .Z(n276) );
  AND U342 ( .A(\one_vote[9].decoder_/sll_39/ML_int[3][6] ), .B(n299), .Z(n277) );
  XOR U343 ( .A(n300), .B(\one_vote[8].decoder_/sll_39/ML_int[3][6] ), .Z(n299) );
  XOR U344 ( .A(n274), .B(n273), .Z(n272) );
  AND U345 ( .A(\one_vote[8].decoder_/sll_39/ML_int[3][6] ), .B(n300), .Z(n273) );
  XOR U346 ( .A(n301), .B(\one_vote[7].decoder_/sll_39/ML_int[3][6] ), .Z(n300) );
  XNOR U347 ( .A(n284), .B(n275), .Z(n274) );
  AND U348 ( .A(\one_vote[7].decoder_/sll_39/ML_int[3][6] ), .B(n301), .Z(n275) );
  XOR U349 ( .A(n302), .B(\one_vote[6].decoder_/sll_39/ML_int[3][6] ), .Z(n301) );
  XOR U350 ( .A(n294), .B(n283), .Z(n284) );
  AND U351 ( .A(\one_vote[6].decoder_/sll_39/ML_int[3][6] ), .B(n302), .Z(n283) );
  XOR U352 ( .A(n303), .B(\one_vote[5].decoder_/sll_39/ML_int[3][6] ), .Z(n302) );
  XNOR U353 ( .A(n304), .B(n289), .Z(n294) );
  XOR U354 ( .A(n290), .B(n305), .Z(n289) );
  AND U355 ( .A(\one_vote[3].decoder_/sll_39/ML_int[3][6] ), .B(n306), .Z(n305) );
  XOR U356 ( .A(n307), .B(n308), .Z(n290) );
  NOR U357 ( .A(n309), .B(n310), .Z(n308) );
  AND U358 ( .A(\decoder_/sll_39/ML_int[3][6] ), .B(
        \one_vote[1].decoder_/sll_39/ML_int[3][6] ), .Z(n310) );
  AND U359 ( .A(\one_vote[2].decoder_/sll_39/ML_int[3][6] ), .B(n311), .Z(n309) );
  XNOR U360 ( .A(\decoder_/sll_39/ML_int[3][6] ), .B(
        \one_vote[1].decoder_/sll_39/ML_int[3][6] ), .Z(n307) );
  XNOR U361 ( .A(n281), .B(n293), .Z(n304) );
  AND U362 ( .A(\one_vote[5].decoder_/sll_39/ML_int[3][6] ), .B(n303), .Z(n293) );
  XOR U363 ( .A(n312), .B(\one_vote[4].decoder_/sll_39/ML_int[3][6] ), .Z(n303) );
  AND U364 ( .A(\one_vote[4].decoder_/sll_39/ML_int[3][6] ), .B(n312), .Z(n281) );
  XOR U365 ( .A(n306), .B(\one_vote[3].decoder_/sll_39/ML_int[3][6] ), .Z(n312) );
  XOR U366 ( .A(\one_vote[2].decoder_/sll_39/ML_int[3][6] ), .B(n311), .Z(n306) );
  XOR U367 ( .A(\decoder_/sll_39/ML_int[3][6] ), .B(
        \one_vote[1].decoder_/sll_39/ML_int[3][6] ), .Z(n311) );
  NOR U368 ( .A(n108), .B(n107), .Z(n122) );
  XNOR U369 ( .A(n313), .B(n314), .Z(n107) );
  AND U370 ( .A(n315), .B(n316), .Z(n314) );
  NOR U371 ( .A(n317), .B(n318), .Z(n316) );
  NOR U372 ( .A(n319), .B(n320), .Z(n315) );
  AND U373 ( .A(n321), .B(n322), .Z(n320) );
  AND U374 ( .A(n323), .B(n324), .Z(n313) );
  NOR U375 ( .A(n325), .B(n326), .Z(n324) );
  AND U376 ( .A(n319), .B(n327), .Z(n326) );
  AND U377 ( .A(n317), .B(n328), .Z(n325) );
  NOR U378 ( .A(n329), .B(n330), .Z(n323) );
  AND U379 ( .A(n331), .B(n332), .Z(n330) );
  AND U380 ( .A(n333), .B(n334), .Z(n332) );
  IV U381 ( .A(n335), .Z(n334) );
  NOR U382 ( .A(n336), .B(n337), .Z(n333) );
  NOR U383 ( .A(n338), .B(n339), .Z(n331) );
  AND U384 ( .A(n318), .B(n340), .Z(n329) );
  AND U385 ( .A(n80), .B(n341), .Z(n108) );
  XOR U386 ( .A(n321), .B(n341), .Z(n80) );
  AND U387 ( .A(n92), .B(n342), .Z(n341) );
  XOR U388 ( .A(n343), .B(n342), .Z(n92) );
  AND U389 ( .A(\one_vote[15].decoder_/sll_39/ML_int[3][7] ), .B(n117), .Z(
        n342) );
  XOR U390 ( .A(n344), .B(\one_vote[14].decoder_/sll_39/ML_int[3][7] ), .Z(
        n117) );
  XNOR U391 ( .A(n328), .B(n322), .Z(n321) );
  AND U392 ( .A(n343), .B(n345), .Z(n322) );
  XOR U393 ( .A(n346), .B(n345), .Z(n343) );
  AND U394 ( .A(\one_vote[14].decoder_/sll_39/ML_int[3][7] ), .B(n344), .Z(
        n345) );
  XOR U395 ( .A(n347), .B(\one_vote[13].decoder_/sll_39/ML_int[3][7] ), .Z(
        n344) );
  XOR U396 ( .A(n327), .B(n317), .Z(n328) );
  AND U397 ( .A(n346), .B(n348), .Z(n317) );
  XOR U398 ( .A(n349), .B(n348), .Z(n346) );
  AND U399 ( .A(\one_vote[13].decoder_/sll_39/ML_int[3][7] ), .B(n347), .Z(
        n348) );
  XOR U400 ( .A(n350), .B(\one_vote[12].decoder_/sll_39/ML_int[3][7] ), .Z(
        n347) );
  XOR U401 ( .A(n340), .B(n319), .Z(n327) );
  AND U402 ( .A(n349), .B(n351), .Z(n319) );
  XOR U403 ( .A(n352), .B(n351), .Z(n349) );
  AND U404 ( .A(\one_vote[12].decoder_/sll_39/ML_int[3][7] ), .B(n350), .Z(
        n351) );
  XOR U405 ( .A(n353), .B(\one_vote[11].decoder_/sll_39/ML_int[3][7] ), .Z(
        n350) );
  XNOR U406 ( .A(n354), .B(n355), .Z(n340) );
  XOR U407 ( .A(n338), .B(n356), .Z(n355) );
  XOR U408 ( .A(n336), .B(n335), .Z(n356) );
  AND U409 ( .A(n357), .B(n358), .Z(n335) );
  AND U410 ( .A(n359), .B(n360), .Z(n336) );
  AND U411 ( .A(n361), .B(n362), .Z(n338) );
  XNOR U412 ( .A(n363), .B(n337), .Z(n354) );
  XOR U413 ( .A(n364), .B(n365), .Z(n337) );
  XOR U414 ( .A(n366), .B(n367), .Z(n365) );
  AND U415 ( .A(n368), .B(n369), .Z(n367) );
  XNOR U416 ( .A(n370), .B(n371), .Z(n364) );
  NOR U417 ( .A(n372), .B(n373), .Z(n371) );
  AND U418 ( .A(n374), .B(n375), .Z(n373) );
  IV U419 ( .A(n376), .Z(n372) );
  NOR U420 ( .A(n366), .B(n377), .Z(n376) );
  AND U421 ( .A(n378), .B(n379), .Z(n377) );
  NOR U422 ( .A(n368), .B(n378), .Z(n370) );
  XNOR U423 ( .A(n339), .B(n318), .Z(n363) );
  AND U424 ( .A(n352), .B(n380), .Z(n318) );
  XOR U425 ( .A(n381), .B(n380), .Z(n352) );
  AND U426 ( .A(\one_vote[11].decoder_/sll_39/ML_int[3][7] ), .B(n353), .Z(
        n380) );
  XOR U427 ( .A(n382), .B(\one_vote[10].decoder_/sll_39/ML_int[3][7] ), .Z(
        n353) );
  AND U428 ( .A(n381), .B(n383), .Z(n339) );
  XOR U429 ( .A(n361), .B(n383), .Z(n381) );
  AND U430 ( .A(\one_vote[10].decoder_/sll_39/ML_int[3][7] ), .B(n382), .Z(
        n383) );
  XOR U431 ( .A(n384), .B(\one_vote[9].decoder_/sll_39/ML_int[3][7] ), .Z(n382) );
  XOR U432 ( .A(n357), .B(n362), .Z(n361) );
  AND U433 ( .A(\one_vote[9].decoder_/sll_39/ML_int[3][7] ), .B(n384), .Z(n362) );
  XOR U434 ( .A(n385), .B(\one_vote[8].decoder_/sll_39/ML_int[3][7] ), .Z(n384) );
  XOR U435 ( .A(n359), .B(n358), .Z(n357) );
  AND U436 ( .A(\one_vote[8].decoder_/sll_39/ML_int[3][7] ), .B(n385), .Z(n358) );
  XOR U437 ( .A(n386), .B(\one_vote[7].decoder_/sll_39/ML_int[3][7] ), .Z(n385) );
  XNOR U438 ( .A(n369), .B(n360), .Z(n359) );
  AND U439 ( .A(\one_vote[7].decoder_/sll_39/ML_int[3][7] ), .B(n386), .Z(n360) );
  XOR U440 ( .A(n387), .B(\one_vote[6].decoder_/sll_39/ML_int[3][7] ), .Z(n386) );
  XOR U441 ( .A(n379), .B(n368), .Z(n369) );
  AND U442 ( .A(\one_vote[6].decoder_/sll_39/ML_int[3][7] ), .B(n387), .Z(n368) );
  XOR U443 ( .A(n388), .B(\one_vote[5].decoder_/sll_39/ML_int[3][7] ), .Z(n387) );
  XNOR U444 ( .A(n389), .B(n374), .Z(n379) );
  XOR U445 ( .A(n375), .B(n390), .Z(n374) );
  AND U446 ( .A(\one_vote[3].decoder_/sll_39/ML_int[3][7] ), .B(n391), .Z(n390) );
  XOR U447 ( .A(n392), .B(n393), .Z(n375) );
  NOR U448 ( .A(n394), .B(n395), .Z(n393) );
  AND U449 ( .A(\decoder_/sll_39/ML_int[3][7] ), .B(
        \one_vote[1].decoder_/sll_39/ML_int[3][7] ), .Z(n395) );
  AND U450 ( .A(\one_vote[2].decoder_/sll_39/ML_int[3][7] ), .B(n396), .Z(n394) );
  XNOR U451 ( .A(\decoder_/sll_39/ML_int[3][7] ), .B(
        \one_vote[1].decoder_/sll_39/ML_int[3][7] ), .Z(n392) );
  XNOR U452 ( .A(n366), .B(n378), .Z(n389) );
  AND U453 ( .A(\one_vote[5].decoder_/sll_39/ML_int[3][7] ), .B(n388), .Z(n378) );
  XOR U454 ( .A(n397), .B(\one_vote[4].decoder_/sll_39/ML_int[3][7] ), .Z(n388) );
  AND U455 ( .A(\one_vote[4].decoder_/sll_39/ML_int[3][7] ), .B(n397), .Z(n366) );
  XOR U456 ( .A(n391), .B(\one_vote[3].decoder_/sll_39/ML_int[3][7] ), .Z(n397) );
  XOR U457 ( .A(\one_vote[2].decoder_/sll_39/ML_int[3][7] ), .B(n396), .Z(n391) );
  XOR U458 ( .A(\decoder_/sll_39/ML_int[3][7] ), .B(
        \one_vote[1].decoder_/sll_39/ML_int[3][7] ), .Z(n396) );
  NOR U459 ( .A(n398), .B(n152), .Z(n227) );
  IV U460 ( .A(n399), .Z(n152) );
  AND U461 ( .A(n149), .B(n148), .Z(n399) );
  NOR U462 ( .A(n146), .B(n145), .Z(n148) );
  XOR U463 ( .A(n400), .B(n401), .Z(n145) );
  XOR U464 ( .A(n402), .B(n403), .Z(n401) );
  NOR U465 ( .A(n404), .B(n405), .Z(n403) );
  NOR U466 ( .A(n406), .B(n407), .Z(n402) );
  AND U467 ( .A(n408), .B(n409), .Z(n407) );
  IV U468 ( .A(n410), .Z(n406) );
  NOR U469 ( .A(n411), .B(n412), .Z(n410) );
  AND U470 ( .A(n404), .B(n413), .Z(n412) );
  AND U471 ( .A(n405), .B(n414), .Z(n411) );
  XNOR U472 ( .A(n415), .B(n416), .Z(n400) );
  AND U473 ( .A(n417), .B(n418), .Z(n416) );
  AND U474 ( .A(n419), .B(n420), .Z(n415) );
  AND U475 ( .A(n421), .B(n422), .Z(n420) );
  IV U476 ( .A(n423), .Z(n422) );
  NOR U477 ( .A(n424), .B(n425), .Z(n421) );
  NOR U478 ( .A(n426), .B(n427), .Z(n419) );
  AND U479 ( .A(n81), .B(n428), .Z(n146) );
  XOR U480 ( .A(n417), .B(n428), .Z(n81) );
  AND U481 ( .A(n93), .B(n429), .Z(n428) );
  XOR U482 ( .A(n430), .B(n429), .Z(n93) );
  AND U483 ( .A(\one_vote[15].decoder_/sll_39/ML_int[3][4] ), .B(n150), .Z(
        n429) );
  XOR U484 ( .A(n431), .B(\one_vote[14].decoder_/sll_39/ML_int[3][4] ), .Z(
        n150) );
  XNOR U485 ( .A(n414), .B(n418), .Z(n417) );
  AND U486 ( .A(n430), .B(n432), .Z(n418) );
  XOR U487 ( .A(n433), .B(n432), .Z(n430) );
  AND U488 ( .A(\one_vote[14].decoder_/sll_39/ML_int[3][4] ), .B(n431), .Z(
        n432) );
  XOR U489 ( .A(n434), .B(\one_vote[13].decoder_/sll_39/ML_int[3][4] ), .Z(
        n431) );
  XOR U490 ( .A(n413), .B(n405), .Z(n414) );
  AND U491 ( .A(n433), .B(n435), .Z(n405) );
  XOR U492 ( .A(n436), .B(n435), .Z(n433) );
  AND U493 ( .A(\one_vote[13].decoder_/sll_39/ML_int[3][4] ), .B(n434), .Z(
        n435) );
  XOR U494 ( .A(n437), .B(\one_vote[12].decoder_/sll_39/ML_int[3][4] ), .Z(
        n434) );
  XNOR U495 ( .A(n408), .B(n404), .Z(n413) );
  AND U496 ( .A(n436), .B(n438), .Z(n404) );
  XOR U497 ( .A(n439), .B(n438), .Z(n436) );
  AND U498 ( .A(\one_vote[12].decoder_/sll_39/ML_int[3][4] ), .B(n437), .Z(
        n438) );
  XOR U499 ( .A(n440), .B(\one_vote[11].decoder_/sll_39/ML_int[3][4] ), .Z(
        n437) );
  XOR U500 ( .A(n441), .B(n442), .Z(n408) );
  XOR U501 ( .A(n426), .B(n443), .Z(n442) );
  XOR U502 ( .A(n424), .B(n423), .Z(n443) );
  AND U503 ( .A(n444), .B(n445), .Z(n423) );
  AND U504 ( .A(n446), .B(n447), .Z(n424) );
  AND U505 ( .A(n448), .B(n449), .Z(n426) );
  XNOR U506 ( .A(n450), .B(n425), .Z(n441) );
  XOR U507 ( .A(n451), .B(n452), .Z(n425) );
  XOR U508 ( .A(n453), .B(n454), .Z(n452) );
  AND U509 ( .A(n455), .B(n456), .Z(n454) );
  XNOR U510 ( .A(n457), .B(n458), .Z(n451) );
  NOR U511 ( .A(n459), .B(n460), .Z(n458) );
  AND U512 ( .A(n461), .B(n462), .Z(n460) );
  IV U513 ( .A(n463), .Z(n459) );
  NOR U514 ( .A(n453), .B(n464), .Z(n463) );
  AND U515 ( .A(n465), .B(n466), .Z(n464) );
  NOR U516 ( .A(n455), .B(n465), .Z(n457) );
  XNOR U517 ( .A(n427), .B(n409), .Z(n450) );
  AND U518 ( .A(n439), .B(n467), .Z(n409) );
  XOR U519 ( .A(n468), .B(n467), .Z(n439) );
  AND U520 ( .A(\one_vote[11].decoder_/sll_39/ML_int[3][4] ), .B(n440), .Z(
        n467) );
  XOR U521 ( .A(n469), .B(\one_vote[10].decoder_/sll_39/ML_int[3][4] ), .Z(
        n440) );
  AND U522 ( .A(n468), .B(n470), .Z(n427) );
  XOR U523 ( .A(n448), .B(n470), .Z(n468) );
  AND U524 ( .A(\one_vote[10].decoder_/sll_39/ML_int[3][4] ), .B(n469), .Z(
        n470) );
  XOR U525 ( .A(n471), .B(\one_vote[9].decoder_/sll_39/ML_int[3][4] ), .Z(n469) );
  XOR U526 ( .A(n444), .B(n449), .Z(n448) );
  AND U527 ( .A(\one_vote[9].decoder_/sll_39/ML_int[3][4] ), .B(n471), .Z(n449) );
  XOR U528 ( .A(n472), .B(\one_vote[8].decoder_/sll_39/ML_int[3][4] ), .Z(n471) );
  XOR U529 ( .A(n446), .B(n445), .Z(n444) );
  AND U530 ( .A(\one_vote[8].decoder_/sll_39/ML_int[3][4] ), .B(n472), .Z(n445) );
  XOR U531 ( .A(n473), .B(\one_vote[7].decoder_/sll_39/ML_int[3][4] ), .Z(n472) );
  XNOR U532 ( .A(n456), .B(n447), .Z(n446) );
  AND U533 ( .A(\one_vote[7].decoder_/sll_39/ML_int[3][4] ), .B(n473), .Z(n447) );
  XOR U534 ( .A(n474), .B(\one_vote[6].decoder_/sll_39/ML_int[3][4] ), .Z(n473) );
  XOR U535 ( .A(n466), .B(n455), .Z(n456) );
  AND U536 ( .A(\one_vote[6].decoder_/sll_39/ML_int[3][4] ), .B(n474), .Z(n455) );
  XOR U537 ( .A(n475), .B(\one_vote[5].decoder_/sll_39/ML_int[3][4] ), .Z(n474) );
  XNOR U538 ( .A(n476), .B(n461), .Z(n466) );
  XOR U539 ( .A(n462), .B(n477), .Z(n461) );
  AND U540 ( .A(\one_vote[3].decoder_/sll_39/ML_int[3][4] ), .B(n478), .Z(n477) );
  XOR U541 ( .A(n479), .B(n480), .Z(n462) );
  NOR U542 ( .A(n481), .B(n482), .Z(n480) );
  AND U543 ( .A(\decoder_/sll_39/ML_int[3][4] ), .B(
        \one_vote[1].decoder_/sll_39/ML_int[3][4] ), .Z(n482) );
  AND U544 ( .A(\one_vote[2].decoder_/sll_39/ML_int[3][4] ), .B(n483), .Z(n481) );
  XNOR U545 ( .A(\decoder_/sll_39/ML_int[3][4] ), .B(
        \one_vote[1].decoder_/sll_39/ML_int[3][4] ), .Z(n479) );
  XNOR U546 ( .A(n453), .B(n465), .Z(n476) );
  AND U547 ( .A(\one_vote[5].decoder_/sll_39/ML_int[3][4] ), .B(n475), .Z(n465) );
  XOR U548 ( .A(n484), .B(\one_vote[4].decoder_/sll_39/ML_int[3][4] ), .Z(n475) );
  AND U549 ( .A(\one_vote[4].decoder_/sll_39/ML_int[3][4] ), .B(n484), .Z(n453) );
  XOR U550 ( .A(n478), .B(\one_vote[3].decoder_/sll_39/ML_int[3][4] ), .Z(n484) );
  XOR U551 ( .A(\one_vote[2].decoder_/sll_39/ML_int[3][4] ), .B(n483), .Z(n478) );
  XOR U552 ( .A(\decoder_/sll_39/ML_int[3][4] ), .B(
        \one_vote[1].decoder_/sll_39/ML_int[3][4] ), .Z(n483) );
  NOR U553 ( .A(n135), .B(n134), .Z(n149) );
  XNOR U554 ( .A(n485), .B(n486), .Z(n134) );
  AND U555 ( .A(n487), .B(n488), .Z(n486) );
  NOR U556 ( .A(n489), .B(n490), .Z(n488) );
  NOR U557 ( .A(n491), .B(n492), .Z(n487) );
  AND U558 ( .A(n493), .B(n494), .Z(n492) );
  AND U559 ( .A(n495), .B(n496), .Z(n485) );
  NOR U560 ( .A(n497), .B(n498), .Z(n496) );
  AND U561 ( .A(n491), .B(n499), .Z(n498) );
  AND U562 ( .A(n489), .B(n500), .Z(n497) );
  NOR U563 ( .A(n501), .B(n502), .Z(n495) );
  AND U564 ( .A(n503), .B(n504), .Z(n502) );
  AND U565 ( .A(n505), .B(n506), .Z(n504) );
  IV U566 ( .A(n507), .Z(n506) );
  NOR U567 ( .A(n508), .B(n509), .Z(n505) );
  NOR U568 ( .A(n510), .B(n511), .Z(n503) );
  AND U569 ( .A(n490), .B(n512), .Z(n501) );
  AND U570 ( .A(n84), .B(n513), .Z(n135) );
  XOR U571 ( .A(n493), .B(n513), .Z(n84) );
  AND U572 ( .A(n96), .B(n514), .Z(n513) );
  XOR U573 ( .A(n515), .B(n514), .Z(n96) );
  AND U574 ( .A(\one_vote[15].decoder_/sll_39/ML_int[3][5] ), .B(n144), .Z(
        n514) );
  XOR U575 ( .A(n516), .B(\one_vote[14].decoder_/sll_39/ML_int[3][5] ), .Z(
        n144) );
  XNOR U576 ( .A(n500), .B(n494), .Z(n493) );
  AND U577 ( .A(n515), .B(n517), .Z(n494) );
  XOR U578 ( .A(n518), .B(n517), .Z(n515) );
  AND U579 ( .A(\one_vote[14].decoder_/sll_39/ML_int[3][5] ), .B(n516), .Z(
        n517) );
  XOR U580 ( .A(n519), .B(\one_vote[13].decoder_/sll_39/ML_int[3][5] ), .Z(
        n516) );
  XOR U581 ( .A(n499), .B(n489), .Z(n500) );
  AND U582 ( .A(n518), .B(n520), .Z(n489) );
  XOR U583 ( .A(n521), .B(n520), .Z(n518) );
  AND U584 ( .A(\one_vote[13].decoder_/sll_39/ML_int[3][5] ), .B(n519), .Z(
        n520) );
  XOR U585 ( .A(n522), .B(\one_vote[12].decoder_/sll_39/ML_int[3][5] ), .Z(
        n519) );
  XOR U586 ( .A(n512), .B(n491), .Z(n499) );
  AND U587 ( .A(n521), .B(n523), .Z(n491) );
  XOR U588 ( .A(n524), .B(n523), .Z(n521) );
  AND U589 ( .A(\one_vote[12].decoder_/sll_39/ML_int[3][5] ), .B(n522), .Z(
        n523) );
  XOR U590 ( .A(n525), .B(\one_vote[11].decoder_/sll_39/ML_int[3][5] ), .Z(
        n522) );
  XNOR U591 ( .A(n526), .B(n527), .Z(n512) );
  XOR U592 ( .A(n510), .B(n528), .Z(n527) );
  XOR U593 ( .A(n508), .B(n507), .Z(n528) );
  AND U594 ( .A(n529), .B(n530), .Z(n507) );
  AND U595 ( .A(n531), .B(n532), .Z(n508) );
  AND U596 ( .A(n533), .B(n534), .Z(n510) );
  XNOR U597 ( .A(n535), .B(n509), .Z(n526) );
  XOR U598 ( .A(n536), .B(n537), .Z(n509) );
  XOR U599 ( .A(n538), .B(n539), .Z(n537) );
  AND U600 ( .A(n540), .B(n541), .Z(n539) );
  XNOR U601 ( .A(n542), .B(n543), .Z(n536) );
  NOR U602 ( .A(n544), .B(n545), .Z(n543) );
  AND U603 ( .A(n546), .B(n547), .Z(n545) );
  IV U604 ( .A(n548), .Z(n544) );
  NOR U605 ( .A(n538), .B(n549), .Z(n548) );
  AND U606 ( .A(n550), .B(n551), .Z(n549) );
  NOR U607 ( .A(n540), .B(n550), .Z(n542) );
  XNOR U608 ( .A(n511), .B(n490), .Z(n535) );
  AND U609 ( .A(n524), .B(n552), .Z(n490) );
  XOR U610 ( .A(n553), .B(n552), .Z(n524) );
  AND U611 ( .A(\one_vote[11].decoder_/sll_39/ML_int[3][5] ), .B(n525), .Z(
        n552) );
  XOR U612 ( .A(n554), .B(\one_vote[10].decoder_/sll_39/ML_int[3][5] ), .Z(
        n525) );
  AND U613 ( .A(n553), .B(n555), .Z(n511) );
  XOR U614 ( .A(n533), .B(n555), .Z(n553) );
  AND U615 ( .A(\one_vote[10].decoder_/sll_39/ML_int[3][5] ), .B(n554), .Z(
        n555) );
  XOR U616 ( .A(n556), .B(\one_vote[9].decoder_/sll_39/ML_int[3][5] ), .Z(n554) );
  XOR U617 ( .A(n529), .B(n534), .Z(n533) );
  AND U618 ( .A(\one_vote[9].decoder_/sll_39/ML_int[3][5] ), .B(n556), .Z(n534) );
  XOR U619 ( .A(n557), .B(\one_vote[8].decoder_/sll_39/ML_int[3][5] ), .Z(n556) );
  XOR U620 ( .A(n531), .B(n530), .Z(n529) );
  AND U621 ( .A(\one_vote[8].decoder_/sll_39/ML_int[3][5] ), .B(n557), .Z(n530) );
  XOR U622 ( .A(n558), .B(\one_vote[7].decoder_/sll_39/ML_int[3][5] ), .Z(n557) );
  XNOR U623 ( .A(n541), .B(n532), .Z(n531) );
  AND U624 ( .A(\one_vote[7].decoder_/sll_39/ML_int[3][5] ), .B(n558), .Z(n532) );
  XOR U625 ( .A(n559), .B(\one_vote[6].decoder_/sll_39/ML_int[3][5] ), .Z(n558) );
  XOR U626 ( .A(n551), .B(n540), .Z(n541) );
  AND U627 ( .A(\one_vote[6].decoder_/sll_39/ML_int[3][5] ), .B(n559), .Z(n540) );
  XOR U628 ( .A(n560), .B(\one_vote[5].decoder_/sll_39/ML_int[3][5] ), .Z(n559) );
  XNOR U629 ( .A(n561), .B(n546), .Z(n551) );
  XOR U630 ( .A(n547), .B(n562), .Z(n546) );
  AND U631 ( .A(\one_vote[3].decoder_/sll_39/ML_int[3][5] ), .B(n563), .Z(n562) );
  XOR U632 ( .A(n564), .B(n565), .Z(n547) );
  NOR U633 ( .A(n566), .B(n567), .Z(n565) );
  AND U634 ( .A(\decoder_/sll_39/ML_int[3][5] ), .B(
        \one_vote[1].decoder_/sll_39/ML_int[3][5] ), .Z(n567) );
  AND U635 ( .A(\one_vote[2].decoder_/sll_39/ML_int[3][5] ), .B(n568), .Z(n566) );
  XNOR U636 ( .A(\decoder_/sll_39/ML_int[3][5] ), .B(
        \one_vote[1].decoder_/sll_39/ML_int[3][5] ), .Z(n564) );
  XNOR U637 ( .A(n538), .B(n550), .Z(n561) );
  AND U638 ( .A(\one_vote[5].decoder_/sll_39/ML_int[3][5] ), .B(n560), .Z(n550) );
  XOR U639 ( .A(n569), .B(\one_vote[4].decoder_/sll_39/ML_int[3][5] ), .Z(n560) );
  AND U640 ( .A(\one_vote[4].decoder_/sll_39/ML_int[3][5] ), .B(n569), .Z(n538) );
  XOR U641 ( .A(n563), .B(\one_vote[3].decoder_/sll_39/ML_int[3][5] ), .Z(n569) );
  XOR U642 ( .A(\one_vote[2].decoder_/sll_39/ML_int[3][5] ), .B(n568), .Z(n563) );
  XOR U643 ( .A(\decoder_/sll_39/ML_int[3][5] ), .B(
        \one_vote[1].decoder_/sll_39/ML_int[3][5] ), .Z(n568) );
  AND U644 ( .A(n222), .B(n221), .Z(n398) );
  AND U645 ( .A(n570), .B(n571), .Z(n221) );
  AND U646 ( .A(n217), .B(n216), .Z(n222) );
  NOR U647 ( .A(n214), .B(n213), .Z(n216) );
  XOR U648 ( .A(n572), .B(n573), .Z(n213) );
  XOR U649 ( .A(n574), .B(n575), .Z(n573) );
  NOR U650 ( .A(n576), .B(n577), .Z(n575) );
  NOR U651 ( .A(n578), .B(n579), .Z(n574) );
  AND U652 ( .A(n580), .B(n581), .Z(n579) );
  IV U653 ( .A(n582), .Z(n578) );
  NOR U654 ( .A(n583), .B(n584), .Z(n582) );
  AND U655 ( .A(n576), .B(n585), .Z(n584) );
  AND U656 ( .A(n577), .B(n586), .Z(n583) );
  XNOR U657 ( .A(n587), .B(n588), .Z(n572) );
  AND U658 ( .A(n589), .B(n590), .Z(n588) );
  AND U659 ( .A(n591), .B(n592), .Z(n587) );
  AND U660 ( .A(n593), .B(n594), .Z(n592) );
  IV U661 ( .A(n595), .Z(n594) );
  NOR U662 ( .A(n596), .B(n597), .Z(n593) );
  NOR U663 ( .A(n598), .B(n599), .Z(n591) );
  AND U664 ( .A(n171), .B(n600), .Z(n214) );
  XOR U665 ( .A(n589), .B(n600), .Z(n171) );
  AND U666 ( .A(n183), .B(n601), .Z(n600) );
  XOR U667 ( .A(n602), .B(n601), .Z(n183) );
  AND U668 ( .A(n219), .B(n218), .Z(n601) );
  XOR U669 ( .A(n603), .B(n604), .Z(n218) );
  AND U670 ( .A(\one_vote[15].decoder_/sll_39/ML_int[2][2] ), .B(n605), .Z(
        n219) );
  XNOR U671 ( .A(n586), .B(n590), .Z(n589) );
  AND U672 ( .A(n602), .B(n606), .Z(n590) );
  XOR U673 ( .A(n607), .B(n606), .Z(n602) );
  AND U674 ( .A(n604), .B(n603), .Z(n606) );
  XOR U675 ( .A(n608), .B(n609), .Z(n603) );
  AND U676 ( .A(\one_vote[14].decoder_/sll_39/ML_int[2][2] ), .B(n610), .Z(
        n604) );
  XOR U677 ( .A(n585), .B(n577), .Z(n586) );
  AND U678 ( .A(n607), .B(n611), .Z(n577) );
  XOR U679 ( .A(n612), .B(n611), .Z(n607) );
  AND U680 ( .A(n609), .B(n608), .Z(n611) );
  XOR U681 ( .A(n613), .B(n614), .Z(n608) );
  AND U682 ( .A(\one_vote[13].decoder_/sll_39/ML_int[2][2] ), .B(n615), .Z(
        n609) );
  XNOR U683 ( .A(n580), .B(n576), .Z(n585) );
  AND U684 ( .A(n612), .B(n616), .Z(n576) );
  XOR U685 ( .A(n617), .B(n616), .Z(n612) );
  AND U686 ( .A(n614), .B(n613), .Z(n616) );
  XOR U687 ( .A(n618), .B(n619), .Z(n613) );
  AND U688 ( .A(\one_vote[12].decoder_/sll_39/ML_int[2][2] ), .B(n620), .Z(
        n614) );
  XOR U689 ( .A(n621), .B(n622), .Z(n580) );
  XOR U690 ( .A(n598), .B(n623), .Z(n622) );
  XOR U691 ( .A(n596), .B(n595), .Z(n623) );
  AND U692 ( .A(n624), .B(n625), .Z(n595) );
  AND U693 ( .A(n626), .B(n627), .Z(n596) );
  AND U694 ( .A(n628), .B(n629), .Z(n598) );
  XNOR U695 ( .A(n630), .B(n597), .Z(n621) );
  XOR U696 ( .A(n631), .B(n632), .Z(n597) );
  XOR U697 ( .A(n633), .B(n634), .Z(n632) );
  AND U698 ( .A(n635), .B(n636), .Z(n634) );
  XNOR U699 ( .A(n637), .B(n638), .Z(n631) );
  NOR U700 ( .A(n639), .B(n640), .Z(n638) );
  AND U701 ( .A(n641), .B(n642), .Z(n640) );
  IV U702 ( .A(n643), .Z(n639) );
  NOR U703 ( .A(n633), .B(n644), .Z(n643) );
  AND U704 ( .A(n645), .B(n646), .Z(n644) );
  NOR U705 ( .A(n635), .B(n645), .Z(n637) );
  XNOR U706 ( .A(n599), .B(n581), .Z(n630) );
  AND U707 ( .A(n617), .B(n647), .Z(n581) );
  XOR U708 ( .A(n648), .B(n647), .Z(n617) );
  AND U709 ( .A(n619), .B(n618), .Z(n647) );
  XOR U710 ( .A(n649), .B(n650), .Z(n618) );
  AND U711 ( .A(\one_vote[11].decoder_/sll_39/ML_int[2][2] ), .B(n651), .Z(
        n619) );
  AND U712 ( .A(n648), .B(n652), .Z(n599) );
  XOR U713 ( .A(n628), .B(n652), .Z(n648) );
  AND U714 ( .A(n650), .B(n649), .Z(n652) );
  XOR U715 ( .A(n653), .B(n654), .Z(n649) );
  AND U716 ( .A(\one_vote[10].decoder_/sll_39/ML_int[2][2] ), .B(n655), .Z(
        n650) );
  XOR U717 ( .A(n624), .B(n629), .Z(n628) );
  AND U718 ( .A(n654), .B(n653), .Z(n629) );
  XOR U719 ( .A(n656), .B(n657), .Z(n653) );
  AND U720 ( .A(\one_vote[9].decoder_/sll_39/ML_int[2][2] ), .B(n658), .Z(n654) );
  XOR U721 ( .A(n626), .B(n625), .Z(n624) );
  AND U722 ( .A(n657), .B(n656), .Z(n625) );
  XOR U723 ( .A(n659), .B(n660), .Z(n656) );
  AND U724 ( .A(\one_vote[8].decoder_/sll_39/ML_int[2][2] ), .B(n661), .Z(n657) );
  XNOR U725 ( .A(n636), .B(n627), .Z(n626) );
  AND U726 ( .A(n660), .B(n659), .Z(n627) );
  XOR U727 ( .A(n662), .B(n663), .Z(n659) );
  AND U728 ( .A(\one_vote[7].decoder_/sll_39/ML_int[2][2] ), .B(n664), .Z(n660) );
  XOR U729 ( .A(n646), .B(n635), .Z(n636) );
  AND U730 ( .A(n663), .B(n662), .Z(n635) );
  XOR U731 ( .A(n665), .B(n666), .Z(n662) );
  AND U732 ( .A(\one_vote[6].decoder_/sll_39/ML_int[2][2] ), .B(n667), .Z(n663) );
  XNOR U733 ( .A(n668), .B(n641), .Z(n646) );
  XOR U734 ( .A(n642), .B(n669), .Z(n641) );
  AND U735 ( .A(n670), .B(n671), .Z(n669) );
  XOR U736 ( .A(n672), .B(n673), .Z(n642) );
  NOR U737 ( .A(n674), .B(n675), .Z(n673) );
  AND U738 ( .A(n676), .B(n677), .Z(n675) );
  AND U739 ( .A(n678), .B(n679), .Z(n674) );
  XNOR U740 ( .A(n676), .B(n677), .Z(n672) );
  XNOR U741 ( .A(n633), .B(n645), .Z(n668) );
  AND U742 ( .A(n666), .B(n665), .Z(n645) );
  XOR U743 ( .A(n680), .B(n681), .Z(n665) );
  AND U744 ( .A(\one_vote[5].decoder_/sll_39/ML_int[2][2] ), .B(n682), .Z(n666) );
  AND U745 ( .A(n681), .B(n680), .Z(n633) );
  XOR U746 ( .A(n671), .B(n670), .Z(n680) );
  AND U747 ( .A(\one_vote[3].decoder_/sll_39/ML_int[2][2] ), .B(n683), .Z(n670) );
  XOR U748 ( .A(n678), .B(n679), .Z(n671) );
  XOR U749 ( .A(n676), .B(n677), .Z(n679) );
  AND U750 ( .A(\one_vote[1].decoder_/sll_39/ML_int[2][2] ), .B(n684), .Z(n677) );
  AND U751 ( .A(\decoder_/sll_39/ML_int[2][2] ), .B(n685), .Z(n676) );
  AND U752 ( .A(\one_vote[2].decoder_/sll_39/ML_int[2][2] ), .B(n686), .Z(n678) );
  AND U753 ( .A(\one_vote[4].decoder_/sll_39/ML_int[2][2] ), .B(n687), .Z(n681) );
  NOR U754 ( .A(n202), .B(n201), .Z(n217) );
  XNOR U755 ( .A(n688), .B(n689), .Z(n201) );
  AND U756 ( .A(n690), .B(n691), .Z(n689) );
  NOR U757 ( .A(n692), .B(n693), .Z(n691) );
  NOR U758 ( .A(n694), .B(n695), .Z(n690) );
  AND U759 ( .A(n696), .B(n697), .Z(n695) );
  AND U760 ( .A(n698), .B(n699), .Z(n688) );
  NOR U761 ( .A(n700), .B(n701), .Z(n699) );
  AND U762 ( .A(n694), .B(n702), .Z(n701) );
  AND U763 ( .A(n692), .B(n703), .Z(n700) );
  NOR U764 ( .A(n704), .B(n705), .Z(n698) );
  AND U765 ( .A(n706), .B(n707), .Z(n705) );
  AND U766 ( .A(n708), .B(n709), .Z(n707) );
  IV U767 ( .A(n710), .Z(n709) );
  NOR U768 ( .A(n711), .B(n712), .Z(n708) );
  NOR U769 ( .A(n713), .B(n714), .Z(n706) );
  AND U770 ( .A(n693), .B(n715), .Z(n704) );
  AND U771 ( .A(n174), .B(n716), .Z(n202) );
  XOR U772 ( .A(n696), .B(n716), .Z(n174) );
  AND U773 ( .A(n186), .B(n717), .Z(n716) );
  XOR U774 ( .A(n718), .B(n717), .Z(n186) );
  AND U775 ( .A(n212), .B(n211), .Z(n717) );
  XOR U776 ( .A(n719), .B(n720), .Z(n211) );
  AND U777 ( .A(\one_vote[15].decoder_/sll_39/ML_int[2][3] ), .B(n605), .Z(
        n212) );
  XNOR U778 ( .A(n703), .B(n697), .Z(n696) );
  AND U779 ( .A(n718), .B(n721), .Z(n697) );
  XOR U780 ( .A(n722), .B(n721), .Z(n718) );
  AND U781 ( .A(n720), .B(n719), .Z(n721) );
  XOR U782 ( .A(n723), .B(n724), .Z(n719) );
  AND U783 ( .A(\one_vote[14].decoder_/sll_39/ML_int[2][3] ), .B(n610), .Z(
        n720) );
  XOR U784 ( .A(n702), .B(n692), .Z(n703) );
  AND U785 ( .A(n722), .B(n725), .Z(n692) );
  XOR U786 ( .A(n726), .B(n725), .Z(n722) );
  AND U787 ( .A(n724), .B(n723), .Z(n725) );
  XOR U788 ( .A(n727), .B(n728), .Z(n723) );
  AND U789 ( .A(\one_vote[13].decoder_/sll_39/ML_int[2][3] ), .B(n615), .Z(
        n724) );
  XOR U790 ( .A(n715), .B(n694), .Z(n702) );
  AND U791 ( .A(n726), .B(n729), .Z(n694) );
  XOR U792 ( .A(n730), .B(n729), .Z(n726) );
  AND U793 ( .A(n728), .B(n727), .Z(n729) );
  XOR U794 ( .A(n731), .B(n732), .Z(n727) );
  AND U795 ( .A(\one_vote[12].decoder_/sll_39/ML_int[2][3] ), .B(n620), .Z(
        n728) );
  XNOR U796 ( .A(n733), .B(n734), .Z(n715) );
  XOR U797 ( .A(n713), .B(n735), .Z(n734) );
  XOR U798 ( .A(n711), .B(n710), .Z(n735) );
  AND U799 ( .A(n736), .B(n737), .Z(n710) );
  AND U800 ( .A(n738), .B(n739), .Z(n711) );
  AND U801 ( .A(n740), .B(n741), .Z(n713) );
  XNOR U802 ( .A(n742), .B(n712), .Z(n733) );
  XOR U803 ( .A(n743), .B(n744), .Z(n712) );
  XOR U804 ( .A(n745), .B(n746), .Z(n744) );
  AND U805 ( .A(n747), .B(n748), .Z(n746) );
  XNOR U806 ( .A(n749), .B(n750), .Z(n743) );
  NOR U807 ( .A(n751), .B(n752), .Z(n750) );
  AND U808 ( .A(n753), .B(n754), .Z(n752) );
  IV U809 ( .A(n755), .Z(n751) );
  NOR U810 ( .A(n745), .B(n756), .Z(n755) );
  AND U811 ( .A(n757), .B(n758), .Z(n756) );
  NOR U812 ( .A(n747), .B(n757), .Z(n749) );
  XNOR U813 ( .A(n714), .B(n693), .Z(n742) );
  AND U814 ( .A(n730), .B(n759), .Z(n693) );
  XOR U815 ( .A(n760), .B(n759), .Z(n730) );
  AND U816 ( .A(n732), .B(n731), .Z(n759) );
  XOR U817 ( .A(n761), .B(n762), .Z(n731) );
  AND U818 ( .A(\one_vote[11].decoder_/sll_39/ML_int[2][3] ), .B(n651), .Z(
        n732) );
  AND U819 ( .A(n760), .B(n763), .Z(n714) );
  XOR U820 ( .A(n740), .B(n763), .Z(n760) );
  AND U821 ( .A(n762), .B(n761), .Z(n763) );
  XOR U822 ( .A(n764), .B(n765), .Z(n761) );
  AND U823 ( .A(\one_vote[10].decoder_/sll_39/ML_int[2][3] ), .B(n655), .Z(
        n762) );
  XOR U824 ( .A(n736), .B(n741), .Z(n740) );
  AND U825 ( .A(n765), .B(n764), .Z(n741) );
  XOR U826 ( .A(n766), .B(n767), .Z(n764) );
  AND U827 ( .A(\one_vote[9].decoder_/sll_39/ML_int[2][3] ), .B(n658), .Z(n765) );
  XOR U828 ( .A(n738), .B(n737), .Z(n736) );
  AND U829 ( .A(n767), .B(n766), .Z(n737) );
  XOR U830 ( .A(n768), .B(n769), .Z(n766) );
  AND U831 ( .A(\one_vote[8].decoder_/sll_39/ML_int[2][3] ), .B(n661), .Z(n767) );
  XNOR U832 ( .A(n748), .B(n739), .Z(n738) );
  AND U833 ( .A(n769), .B(n768), .Z(n739) );
  XOR U834 ( .A(n770), .B(n771), .Z(n768) );
  AND U835 ( .A(\one_vote[7].decoder_/sll_39/ML_int[2][3] ), .B(n664), .Z(n769) );
  XOR U836 ( .A(n758), .B(n747), .Z(n748) );
  AND U837 ( .A(n771), .B(n770), .Z(n747) );
  XOR U838 ( .A(n772), .B(n773), .Z(n770) );
  AND U839 ( .A(\one_vote[6].decoder_/sll_39/ML_int[2][3] ), .B(n667), .Z(n771) );
  XNOR U840 ( .A(n774), .B(n753), .Z(n758) );
  XOR U841 ( .A(n754), .B(n775), .Z(n753) );
  AND U842 ( .A(n776), .B(n777), .Z(n775) );
  XOR U843 ( .A(n778), .B(n779), .Z(n754) );
  NOR U844 ( .A(n780), .B(n781), .Z(n779) );
  AND U845 ( .A(n782), .B(n783), .Z(n781) );
  AND U846 ( .A(n784), .B(n785), .Z(n780) );
  XNOR U847 ( .A(n782), .B(n783), .Z(n778) );
  XNOR U848 ( .A(n745), .B(n757), .Z(n774) );
  AND U849 ( .A(n773), .B(n772), .Z(n757) );
  XOR U850 ( .A(n786), .B(n787), .Z(n772) );
  AND U851 ( .A(\one_vote[5].decoder_/sll_39/ML_int[2][3] ), .B(n682), .Z(n773) );
  AND U852 ( .A(n787), .B(n786), .Z(n745) );
  XOR U853 ( .A(n777), .B(n776), .Z(n786) );
  AND U854 ( .A(\one_vote[3].decoder_/sll_39/ML_int[2][3] ), .B(n683), .Z(n776) );
  XOR U855 ( .A(n784), .B(n785), .Z(n777) );
  XOR U856 ( .A(n782), .B(n783), .Z(n785) );
  AND U857 ( .A(\one_vote[1].decoder_/sll_39/ML_int[2][3] ), .B(n684), .Z(n783) );
  AND U858 ( .A(\decoder_/sll_39/ML_int[2][3] ), .B(n685), .Z(n782) );
  AND U859 ( .A(\one_vote[2].decoder_/sll_39/ML_int[2][3] ), .B(n686), .Z(n784) );
  AND U860 ( .A(\one_vote[4].decoder_/sll_39/ML_int[2][3] ), .B(n687), .Z(n787) );
  XNOR U861 ( .A(n788), .B(n789), .Z(n13) );
  AND U862 ( .A(n790), .B(n791), .Z(n789) );
  XOR U863 ( .A(n788), .B(n166), .Z(n791) );
  XOR U864 ( .A(n571), .B(n792), .Z(n166) );
  AND U865 ( .A(n178), .B(n793), .Z(n792) );
  XOR U866 ( .A(n794), .B(n795), .Z(n571) );
  AND U867 ( .A(n796), .B(n797), .Z(n795) );
  NOR U868 ( .A(n798), .B(n799), .Z(n797) );
  NOR U869 ( .A(n800), .B(n801), .Z(n796) );
  AND U870 ( .A(n802), .B(n803), .Z(n801) );
  AND U871 ( .A(n804), .B(n805), .Z(n794) );
  NOR U872 ( .A(n806), .B(n807), .Z(n805) );
  AND U873 ( .A(n800), .B(n808), .Z(n807) );
  AND U874 ( .A(n798), .B(n809), .Z(n806) );
  NOR U875 ( .A(n810), .B(n811), .Z(n804) );
  AND U876 ( .A(n812), .B(n813), .Z(n811) );
  AND U877 ( .A(n814), .B(n815), .Z(n813) );
  IV U878 ( .A(n816), .Z(n815) );
  NOR U879 ( .A(n817), .B(n818), .Z(n814) );
  NOR U880 ( .A(n819), .B(n820), .Z(n812) );
  AND U881 ( .A(n799), .B(n821), .Z(n810) );
  XNOR U882 ( .A(n165), .B(n788), .Z(n790) );
  XOR U883 ( .A(n570), .B(n822), .Z(n165) );
  AND U884 ( .A(n175), .B(n823), .Z(n822) );
  XNOR U885 ( .A(n824), .B(n825), .Z(n570) );
  XOR U886 ( .A(n826), .B(n827), .Z(n825) );
  NOR U887 ( .A(n828), .B(n829), .Z(n827) );
  NOR U888 ( .A(n830), .B(n831), .Z(n826) );
  AND U889 ( .A(n832), .B(n833), .Z(n831) );
  IV U890 ( .A(n834), .Z(n830) );
  NOR U891 ( .A(n835), .B(n836), .Z(n834) );
  AND U892 ( .A(n828), .B(n837), .Z(n836) );
  AND U893 ( .A(n829), .B(n838), .Z(n835) );
  XNOR U894 ( .A(n839), .B(n840), .Z(n824) );
  AND U895 ( .A(n841), .B(n842), .Z(n840) );
  AND U896 ( .A(n843), .B(n844), .Z(n839) );
  NOR U897 ( .A(n845), .B(n846), .Z(n844) );
  IV U898 ( .A(n847), .Z(n845) );
  NOR U899 ( .A(n848), .B(n849), .Z(n847) );
  NOR U900 ( .A(n850), .B(n851), .Z(n843) );
  XOR U901 ( .A(n852), .B(n853), .Z(n788) );
  AND U902 ( .A(n854), .B(n855), .Z(n853) );
  XNOR U903 ( .A(n852), .B(n178), .Z(n855) );
  XOR U904 ( .A(n802), .B(n793), .Z(n178) );
  AND U905 ( .A(n190), .B(n856), .Z(n793) );
  XNOR U906 ( .A(n809), .B(n803), .Z(n802) );
  AND U907 ( .A(n857), .B(n858), .Z(n803) );
  XOR U908 ( .A(n808), .B(n798), .Z(n809) );
  AND U909 ( .A(n859), .B(n860), .Z(n798) );
  XOR U910 ( .A(n821), .B(n800), .Z(n808) );
  AND U911 ( .A(n861), .B(n862), .Z(n800) );
  XNOR U912 ( .A(n863), .B(n864), .Z(n821) );
  XOR U913 ( .A(n819), .B(n865), .Z(n864) );
  XOR U914 ( .A(n817), .B(n816), .Z(n865) );
  AND U915 ( .A(n866), .B(n867), .Z(n816) );
  AND U916 ( .A(n868), .B(n869), .Z(n817) );
  AND U917 ( .A(n870), .B(n871), .Z(n819) );
  XNOR U918 ( .A(n872), .B(n818), .Z(n863) );
  XOR U919 ( .A(n873), .B(n874), .Z(n818) );
  XOR U920 ( .A(n875), .B(n876), .Z(n874) );
  AND U921 ( .A(n877), .B(n878), .Z(n876) );
  XNOR U922 ( .A(n879), .B(n880), .Z(n873) );
  NOR U923 ( .A(n881), .B(n882), .Z(n880) );
  AND U924 ( .A(n883), .B(n884), .Z(n882) );
  IV U925 ( .A(n885), .Z(n881) );
  NOR U926 ( .A(n875), .B(n886), .Z(n885) );
  AND U927 ( .A(n887), .B(n888), .Z(n886) );
  NOR U928 ( .A(n877), .B(n887), .Z(n879) );
  XNOR U929 ( .A(n820), .B(n799), .Z(n872) );
  AND U930 ( .A(n889), .B(n890), .Z(n799) );
  AND U931 ( .A(n891), .B(n892), .Z(n820) );
  XOR U932 ( .A(n175), .B(n852), .Z(n854) );
  XOR U933 ( .A(n841), .B(n823), .Z(n175) );
  AND U934 ( .A(n187), .B(n893), .Z(n823) );
  XNOR U935 ( .A(n838), .B(n842), .Z(n841) );
  AND U936 ( .A(n894), .B(n895), .Z(n842) );
  XOR U937 ( .A(n837), .B(n829), .Z(n838) );
  AND U938 ( .A(n896), .B(n897), .Z(n829) );
  XNOR U939 ( .A(n832), .B(n828), .Z(n837) );
  AND U940 ( .A(n898), .B(n899), .Z(n828) );
  XOR U941 ( .A(n900), .B(n901), .Z(n832) );
  XOR U942 ( .A(n850), .B(n902), .Z(n901) );
  XOR U943 ( .A(n848), .B(n846), .Z(n902) );
  AND U944 ( .A(n903), .B(n904), .Z(n846) );
  AND U945 ( .A(n905), .B(n906), .Z(n848) );
  AND U946 ( .A(n907), .B(n908), .Z(n850) );
  XNOR U947 ( .A(n909), .B(n849), .Z(n900) );
  XOR U948 ( .A(n910), .B(n911), .Z(n849) );
  XOR U949 ( .A(n912), .B(n913), .Z(n911) );
  AND U950 ( .A(n914), .B(n915), .Z(n913) );
  XNOR U951 ( .A(n916), .B(n917), .Z(n910) );
  NOR U952 ( .A(n918), .B(n919), .Z(n917) );
  AND U953 ( .A(n920), .B(n921), .Z(n919) );
  IV U954 ( .A(n922), .Z(n918) );
  NOR U955 ( .A(n912), .B(n923), .Z(n922) );
  AND U956 ( .A(n924), .B(n925), .Z(n923) );
  NOR U957 ( .A(n914), .B(n924), .Z(n916) );
  XNOR U958 ( .A(n851), .B(n833), .Z(n909) );
  AND U959 ( .A(n926), .B(n927), .Z(n833) );
  AND U960 ( .A(n928), .B(n929), .Z(n851) );
  XOR U961 ( .A(n930), .B(n931), .Z(n852) );
  AND U962 ( .A(n932), .B(n933), .Z(n931) );
  XNOR U963 ( .A(n190), .B(n930), .Z(n933) );
  XOR U964 ( .A(n857), .B(n856), .Z(n190) );
  AND U965 ( .A(n934), .B(n935), .Z(n856) );
  XOR U966 ( .A(n859), .B(n858), .Z(n857) );
  AND U967 ( .A(n936), .B(n937), .Z(n858) );
  XOR U968 ( .A(n861), .B(n860), .Z(n859) );
  AND U969 ( .A(n938), .B(n939), .Z(n860) );
  XOR U970 ( .A(n889), .B(n862), .Z(n861) );
  AND U971 ( .A(n940), .B(n941), .Z(n862) );
  XOR U972 ( .A(n891), .B(n890), .Z(n889) );
  AND U973 ( .A(n942), .B(n943), .Z(n890) );
  XOR U974 ( .A(n870), .B(n892), .Z(n891) );
  AND U975 ( .A(n944), .B(n945), .Z(n892) );
  XOR U976 ( .A(n866), .B(n871), .Z(n870) );
  AND U977 ( .A(n946), .B(n947), .Z(n871) );
  XOR U978 ( .A(n868), .B(n867), .Z(n866) );
  AND U979 ( .A(n948), .B(n949), .Z(n867) );
  XNOR U980 ( .A(n878), .B(n869), .Z(n868) );
  AND U981 ( .A(n950), .B(n951), .Z(n869) );
  XOR U982 ( .A(n888), .B(n877), .Z(n878) );
  AND U983 ( .A(n952), .B(n953), .Z(n877) );
  XNOR U984 ( .A(n954), .B(n883), .Z(n888) );
  XOR U985 ( .A(n884), .B(n955), .Z(n883) );
  AND U986 ( .A(n956), .B(n957), .Z(n955) );
  XOR U987 ( .A(n958), .B(n959), .Z(n884) );
  NOR U988 ( .A(n960), .B(n961), .Z(n959) );
  AND U989 ( .A(n962), .B(n963), .Z(n961) );
  AND U990 ( .A(n964), .B(n965), .Z(n960) );
  XNOR U991 ( .A(n962), .B(n963), .Z(n958) );
  XNOR U992 ( .A(n875), .B(n887), .Z(n954) );
  AND U993 ( .A(n966), .B(n967), .Z(n887) );
  AND U994 ( .A(n968), .B(n969), .Z(n875) );
  XOR U995 ( .A(n930), .B(n187), .Z(n932) );
  XOR U996 ( .A(n894), .B(n893), .Z(n187) );
  AND U997 ( .A(n970), .B(n971), .Z(n893) );
  XOR U998 ( .A(n896), .B(n895), .Z(n894) );
  AND U999 ( .A(n972), .B(n973), .Z(n895) );
  XOR U1000 ( .A(n898), .B(n897), .Z(n896) );
  AND U1001 ( .A(n974), .B(n975), .Z(n897) );
  XOR U1002 ( .A(n926), .B(n899), .Z(n898) );
  AND U1003 ( .A(n976), .B(n977), .Z(n899) );
  XOR U1004 ( .A(n928), .B(n927), .Z(n926) );
  AND U1005 ( .A(n978), .B(n979), .Z(n927) );
  XOR U1006 ( .A(n907), .B(n929), .Z(n928) );
  AND U1007 ( .A(n980), .B(n981), .Z(n929) );
  XOR U1008 ( .A(n903), .B(n908), .Z(n907) );
  AND U1009 ( .A(n982), .B(n983), .Z(n908) );
  XOR U1010 ( .A(n905), .B(n904), .Z(n903) );
  AND U1011 ( .A(n984), .B(n985), .Z(n904) );
  XNOR U1012 ( .A(n915), .B(n906), .Z(n905) );
  AND U1013 ( .A(n986), .B(n987), .Z(n906) );
  XOR U1014 ( .A(n925), .B(n914), .Z(n915) );
  AND U1015 ( .A(n988), .B(n989), .Z(n914) );
  XNOR U1016 ( .A(n990), .B(n920), .Z(n925) );
  XOR U1017 ( .A(n921), .B(n991), .Z(n920) );
  AND U1018 ( .A(n992), .B(n993), .Z(n991) );
  XOR U1019 ( .A(n994), .B(n995), .Z(n921) );
  NOR U1020 ( .A(n996), .B(n997), .Z(n995) );
  AND U1021 ( .A(n998), .B(n999), .Z(n997) );
  AND U1022 ( .A(n1000), .B(n1001), .Z(n996) );
  XNOR U1023 ( .A(n998), .B(n999), .Z(n994) );
  XNOR U1024 ( .A(n912), .B(n924), .Z(n990) );
  AND U1025 ( .A(n1002), .B(n1003), .Z(n924) );
  AND U1026 ( .A(n1004), .B(n1005), .Z(n912) );
  NOR U1027 ( .A(n223), .B(n226), .Z(n930) );
  XNOR U1028 ( .A(n935), .B(n934), .Z(n226) );
  AND U1029 ( .A(\one_vote[15].decoder_/sll_39/ML_int[2][1] ), .B(n605), .Z(
        n934) );
  NOR U1030 ( .A(n1006), .B(p_input[46]), .Z(
        \one_vote[15].decoder_/sll_39/ML_int[2][1] ) );
  XOR U1031 ( .A(n937), .B(n936), .Z(n935) );
  AND U1032 ( .A(\one_vote[14].decoder_/sll_39/ML_int[2][1] ), .B(n610), .Z(
        n936) );
  NOR U1033 ( .A(n1007), .B(p_input[43]), .Z(
        \one_vote[14].decoder_/sll_39/ML_int[2][1] ) );
  XOR U1034 ( .A(n939), .B(n938), .Z(n937) );
  AND U1035 ( .A(\one_vote[13].decoder_/sll_39/ML_int[2][1] ), .B(n615), .Z(
        n938) );
  NOR U1036 ( .A(n1008), .B(p_input[40]), .Z(
        \one_vote[13].decoder_/sll_39/ML_int[2][1] ) );
  XOR U1037 ( .A(n941), .B(n940), .Z(n939) );
  AND U1038 ( .A(\one_vote[12].decoder_/sll_39/ML_int[2][1] ), .B(n620), .Z(
        n940) );
  NOR U1039 ( .A(n1009), .B(p_input[37]), .Z(
        \one_vote[12].decoder_/sll_39/ML_int[2][1] ) );
  XOR U1040 ( .A(n943), .B(n942), .Z(n941) );
  AND U1041 ( .A(\one_vote[11].decoder_/sll_39/ML_int[2][1] ), .B(n651), .Z(
        n942) );
  NOR U1042 ( .A(n1010), .B(p_input[34]), .Z(
        \one_vote[11].decoder_/sll_39/ML_int[2][1] ) );
  XOR U1043 ( .A(n945), .B(n944), .Z(n943) );
  AND U1044 ( .A(\one_vote[10].decoder_/sll_39/ML_int[2][1] ), .B(n655), .Z(
        n944) );
  NOR U1045 ( .A(n1011), .B(p_input[31]), .Z(
        \one_vote[10].decoder_/sll_39/ML_int[2][1] ) );
  XOR U1046 ( .A(n947), .B(n946), .Z(n945) );
  AND U1047 ( .A(\one_vote[9].decoder_/sll_39/ML_int[2][1] ), .B(n658), .Z(
        n946) );
  NOR U1048 ( .A(n1012), .B(p_input[28]), .Z(
        \one_vote[9].decoder_/sll_39/ML_int[2][1] ) );
  XOR U1049 ( .A(n949), .B(n948), .Z(n947) );
  AND U1050 ( .A(\one_vote[8].decoder_/sll_39/ML_int[2][1] ), .B(n661), .Z(
        n948) );
  NOR U1051 ( .A(n1013), .B(p_input[25]), .Z(
        \one_vote[8].decoder_/sll_39/ML_int[2][1] ) );
  XOR U1052 ( .A(n951), .B(n950), .Z(n949) );
  AND U1053 ( .A(\one_vote[7].decoder_/sll_39/ML_int[2][1] ), .B(n664), .Z(
        n950) );
  NOR U1054 ( .A(n1014), .B(p_input[22]), .Z(
        \one_vote[7].decoder_/sll_39/ML_int[2][1] ) );
  XOR U1055 ( .A(n953), .B(n952), .Z(n951) );
  AND U1056 ( .A(\one_vote[6].decoder_/sll_39/ML_int[2][1] ), .B(n667), .Z(
        n952) );
  NOR U1057 ( .A(n1015), .B(p_input[19]), .Z(
        \one_vote[6].decoder_/sll_39/ML_int[2][1] ) );
  XOR U1058 ( .A(n967), .B(n966), .Z(n953) );
  AND U1059 ( .A(\one_vote[5].decoder_/sll_39/ML_int[2][1] ), .B(n682), .Z(
        n966) );
  NOR U1060 ( .A(n1016), .B(p_input[16]), .Z(
        \one_vote[5].decoder_/sll_39/ML_int[2][1] ) );
  XOR U1061 ( .A(n969), .B(n968), .Z(n967) );
  AND U1062 ( .A(\one_vote[4].decoder_/sll_39/ML_int[2][1] ), .B(n687), .Z(
        n968) );
  NOR U1063 ( .A(n1017), .B(p_input[13]), .Z(
        \one_vote[4].decoder_/sll_39/ML_int[2][1] ) );
  XOR U1064 ( .A(n957), .B(n956), .Z(n969) );
  AND U1065 ( .A(\one_vote[3].decoder_/sll_39/ML_int[2][1] ), .B(n683), .Z(
        n956) );
  NOR U1066 ( .A(n1018), .B(p_input[10]), .Z(
        \one_vote[3].decoder_/sll_39/ML_int[2][1] ) );
  XOR U1067 ( .A(n964), .B(n965), .Z(n957) );
  XOR U1068 ( .A(n962), .B(n963), .Z(n965) );
  AND U1069 ( .A(\one_vote[1].decoder_/sll_39/ML_int[2][1] ), .B(n684), .Z(
        n963) );
  NOR U1070 ( .A(n1020), .B(p_input[4]), .Z(
        \one_vote[1].decoder_/sll_39/ML_int[2][1] ) );
  AND U1071 ( .A(\decoder_/sll_39/ML_int[2][1] ), .B(n685), .Z(n962) );
  AND U1072 ( .A(\one_vote[2].decoder_/sll_39/ML_int[2][1] ), .B(n686), .Z(
        n964) );
  NOR U1073 ( .A(n1019), .B(p_input[7]), .Z(
        \one_vote[2].decoder_/sll_39/ML_int[2][1] ) );
  XOR U1074 ( .A(n971), .B(n970), .Z(n223) );
  AND U1075 ( .A(\one_vote[15].decoder_/sll_39/ML_int[2][0] ), .B(n605), .Z(
        n970) );
  IV U1076 ( .A(p_input[47]), .Z(n605) );
  NOR U1077 ( .A(p_input[46]), .B(p_input[45]), .Z(
        \one_vote[15].decoder_/sll_39/ML_int[2][0] ) );
  XOR U1078 ( .A(n973), .B(n972), .Z(n971) );
  AND U1079 ( .A(\one_vote[14].decoder_/sll_39/ML_int[2][0] ), .B(n610), .Z(
        n972) );
  IV U1080 ( .A(p_input[44]), .Z(n610) );
  NOR U1081 ( .A(p_input[43]), .B(p_input[42]), .Z(
        \one_vote[14].decoder_/sll_39/ML_int[2][0] ) );
  XOR U1082 ( .A(n975), .B(n974), .Z(n973) );
  AND U1083 ( .A(\one_vote[13].decoder_/sll_39/ML_int[2][0] ), .B(n615), .Z(
        n974) );
  IV U1084 ( .A(p_input[41]), .Z(n615) );
  NOR U1085 ( .A(p_input[40]), .B(p_input[39]), .Z(
        \one_vote[13].decoder_/sll_39/ML_int[2][0] ) );
  XOR U1086 ( .A(n977), .B(n976), .Z(n975) );
  AND U1087 ( .A(\one_vote[12].decoder_/sll_39/ML_int[2][0] ), .B(n620), .Z(
        n976) );
  IV U1088 ( .A(p_input[38]), .Z(n620) );
  NOR U1089 ( .A(p_input[37]), .B(p_input[36]), .Z(
        \one_vote[12].decoder_/sll_39/ML_int[2][0] ) );
  XOR U1090 ( .A(n979), .B(n978), .Z(n977) );
  AND U1091 ( .A(\one_vote[11].decoder_/sll_39/ML_int[2][0] ), .B(n651), .Z(
        n978) );
  IV U1092 ( .A(p_input[35]), .Z(n651) );
  NOR U1093 ( .A(p_input[34]), .B(p_input[33]), .Z(
        \one_vote[11].decoder_/sll_39/ML_int[2][0] ) );
  XOR U1094 ( .A(n981), .B(n980), .Z(n979) );
  AND U1095 ( .A(\one_vote[10].decoder_/sll_39/ML_int[2][0] ), .B(n655), .Z(
        n980) );
  IV U1096 ( .A(p_input[32]), .Z(n655) );
  NOR U1097 ( .A(p_input[31]), .B(p_input[30]), .Z(
        \one_vote[10].decoder_/sll_39/ML_int[2][0] ) );
  XOR U1098 ( .A(n983), .B(n982), .Z(n981) );
  AND U1099 ( .A(\one_vote[9].decoder_/sll_39/ML_int[2][0] ), .B(n658), .Z(
        n982) );
  IV U1100 ( .A(p_input[29]), .Z(n658) );
  NOR U1101 ( .A(p_input[28]), .B(p_input[27]), .Z(
        \one_vote[9].decoder_/sll_39/ML_int[2][0] ) );
  XOR U1102 ( .A(n985), .B(n984), .Z(n983) );
  AND U1103 ( .A(\one_vote[8].decoder_/sll_39/ML_int[2][0] ), .B(n661), .Z(
        n984) );
  IV U1104 ( .A(p_input[26]), .Z(n661) );
  NOR U1105 ( .A(p_input[25]), .B(p_input[24]), .Z(
        \one_vote[8].decoder_/sll_39/ML_int[2][0] ) );
  XOR U1106 ( .A(n987), .B(n986), .Z(n985) );
  AND U1107 ( .A(\one_vote[7].decoder_/sll_39/ML_int[2][0] ), .B(n664), .Z(
        n986) );
  IV U1108 ( .A(p_input[23]), .Z(n664) );
  NOR U1109 ( .A(p_input[22]), .B(p_input[21]), .Z(
        \one_vote[7].decoder_/sll_39/ML_int[2][0] ) );
  XOR U1110 ( .A(n989), .B(n988), .Z(n987) );
  AND U1111 ( .A(\one_vote[6].decoder_/sll_39/ML_int[2][0] ), .B(n667), .Z(
        n988) );
  IV U1112 ( .A(p_input[20]), .Z(n667) );
  NOR U1113 ( .A(p_input[19]), .B(p_input[18]), .Z(
        \one_vote[6].decoder_/sll_39/ML_int[2][0] ) );
  XOR U1114 ( .A(n1003), .B(n1002), .Z(n989) );
  AND U1115 ( .A(\one_vote[5].decoder_/sll_39/ML_int[2][0] ), .B(n682), .Z(
        n1002) );
  IV U1116 ( .A(p_input[17]), .Z(n682) );
  NOR U1117 ( .A(p_input[16]), .B(p_input[15]), .Z(
        \one_vote[5].decoder_/sll_39/ML_int[2][0] ) );
  XOR U1118 ( .A(n1005), .B(n1004), .Z(n1003) );
  AND U1119 ( .A(\one_vote[4].decoder_/sll_39/ML_int[2][0] ), .B(n687), .Z(
        n1004) );
  IV U1120 ( .A(p_input[14]), .Z(n687) );
  NOR U1121 ( .A(p_input[13]), .B(p_input[12]), .Z(
        \one_vote[4].decoder_/sll_39/ML_int[2][0] ) );
  XOR U1122 ( .A(n993), .B(n992), .Z(n1005) );
  AND U1123 ( .A(\one_vote[3].decoder_/sll_39/ML_int[2][0] ), .B(n683), .Z(
        n992) );
  IV U1124 ( .A(p_input[11]), .Z(n683) );
  NOR U1125 ( .A(p_input[9]), .B(p_input[10]), .Z(
        \one_vote[3].decoder_/sll_39/ML_int[2][0] ) );
  XOR U1126 ( .A(n1000), .B(n1001), .Z(n993) );
  XOR U1127 ( .A(n998), .B(n999), .Z(n1001) );
  AND U1128 ( .A(\one_vote[1].decoder_/sll_39/ML_int[2][0] ), .B(n684), .Z(
        n999) );
  IV U1129 ( .A(p_input[5]), .Z(n684) );
  NOR U1130 ( .A(p_input[4]), .B(p_input[3]), .Z(
        \one_vote[1].decoder_/sll_39/ML_int[2][0] ) );
  AND U1131 ( .A(\decoder_/sll_39/ML_int[2][0] ), .B(n685), .Z(n998) );
  IV U1132 ( .A(p_input[2]), .Z(n685) );
  AND U1133 ( .A(\one_vote[2].decoder_/sll_39/ML_int[2][0] ), .B(n686), .Z(
        n1000) );
  IV U1134 ( .A(p_input[8]), .Z(n686) );
  NOR U1135 ( .A(p_input[7]), .B(p_input[6]), .Z(
        \one_vote[2].decoder_/sll_39/ML_int[2][0] ) );
  IV U1136 ( .A(p_input[45]), .Z(n1006) );
  IV U1137 ( .A(p_input[42]), .Z(n1007) );
  IV U1138 ( .A(p_input[39]), .Z(n1008) );
  IV U1139 ( .A(p_input[36]), .Z(n1009) );
  IV U1140 ( .A(p_input[33]), .Z(n1010) );
  IV U1141 ( .A(p_input[30]), .Z(n1011) );
  IV U1142 ( .A(p_input[27]), .Z(n1012) );
  IV U1143 ( .A(p_input[24]), .Z(n1013) );
  IV U1144 ( .A(p_input[21]), .Z(n1014) );
  IV U1145 ( .A(p_input[18]), .Z(n1015) );
  IV U1146 ( .A(p_input[15]), .Z(n1016) );
  IV U1147 ( .A(p_input[12]), .Z(n1017) );
  IV U1148 ( .A(p_input[9]), .Z(n1018) );
  IV U1149 ( .A(p_input[6]), .Z(n1019) );
  IV U1150 ( .A(p_input[3]), .Z(n1020) );
  NOR U1151 ( .A(n1021), .B(p_input[1]), .Z(\decoder_/sll_39/ML_int[2][1] ) );
  IV U1152 ( .A(p_input[0]), .Z(n1021) );
  NOR U1153 ( .A(p_input[1]), .B(p_input[0]), .Z(
        \decoder_/sll_39/ML_int[2][0] ) );
endmodule

