
module auction_BMR_N8_W16 ( p_input, o );
  input [4095:0] p_input;
  output [23:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245;

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(o[7]), .B(n3), .Z(n1) );
  XOR U3 ( .A(n4), .B(n5), .Z(n3) );
  XNOR U4 ( .A(n6), .B(n7), .Z(o[8]) );
  AND U5 ( .A(o[7]), .B(n8), .Z(n6) );
  XNOR U6 ( .A(n9), .B(n7), .Z(n8) );
  XOR U7 ( .A(n10), .B(n11), .Z(o[23]) );
  AND U8 ( .A(o[7]), .B(n12), .Z(n10) );
  XOR U9 ( .A(n13), .B(n14), .Z(n12) );
  XOR U10 ( .A(n15), .B(n16), .Z(o[22]) );
  AND U11 ( .A(o[7]), .B(n17), .Z(n15) );
  XOR U12 ( .A(n18), .B(n19), .Z(n17) );
  XOR U13 ( .A(n20), .B(n21), .Z(o[21]) );
  AND U14 ( .A(o[7]), .B(n22), .Z(n20) );
  XOR U15 ( .A(n23), .B(n24), .Z(n22) );
  XOR U16 ( .A(n25), .B(n26), .Z(o[20]) );
  AND U17 ( .A(o[7]), .B(n27), .Z(n25) );
  XOR U18 ( .A(n28), .B(n29), .Z(n27) );
  XOR U19 ( .A(n30), .B(n31), .Z(o[19]) );
  AND U20 ( .A(o[7]), .B(n32), .Z(n30) );
  XOR U21 ( .A(n33), .B(n34), .Z(n32) );
  XOR U22 ( .A(n35), .B(n36), .Z(o[18]) );
  AND U23 ( .A(o[7]), .B(n37), .Z(n35) );
  XOR U24 ( .A(n38), .B(n39), .Z(n37) );
  XOR U25 ( .A(n40), .B(n41), .Z(o[17]) );
  AND U26 ( .A(o[7]), .B(n42), .Z(n40) );
  XOR U27 ( .A(n43), .B(n44), .Z(n42) );
  XOR U28 ( .A(n45), .B(n46), .Z(o[16]) );
  AND U29 ( .A(o[7]), .B(n47), .Z(n45) );
  XOR U30 ( .A(n48), .B(n49), .Z(n47) );
  XOR U31 ( .A(n50), .B(n51), .Z(o[15]) );
  AND U32 ( .A(o[7]), .B(n52), .Z(n50) );
  XOR U33 ( .A(n53), .B(n54), .Z(n52) );
  XOR U34 ( .A(n55), .B(n56), .Z(o[14]) );
  AND U35 ( .A(o[7]), .B(n57), .Z(n55) );
  XOR U36 ( .A(n58), .B(n59), .Z(n57) );
  XOR U37 ( .A(n60), .B(n61), .Z(o[13]) );
  AND U38 ( .A(o[7]), .B(n62), .Z(n60) );
  XOR U39 ( .A(n63), .B(n64), .Z(n62) );
  XOR U40 ( .A(n65), .B(n66), .Z(o[12]) );
  AND U41 ( .A(o[7]), .B(n67), .Z(n65) );
  XOR U42 ( .A(n68), .B(n69), .Z(n67) );
  XOR U43 ( .A(n70), .B(n71), .Z(o[11]) );
  AND U44 ( .A(o[7]), .B(n72), .Z(n70) );
  XOR U45 ( .A(n73), .B(n74), .Z(n72) );
  XOR U46 ( .A(n75), .B(n76), .Z(o[10]) );
  AND U47 ( .A(o[7]), .B(n77), .Z(n75) );
  XOR U48 ( .A(n78), .B(n79), .Z(n77) );
  XOR U49 ( .A(n80), .B(n81), .Z(o[0]) );
  AND U50 ( .A(o[1]), .B(n82), .Z(n81) );
  XNOR U51 ( .A(n83), .B(n84), .Z(n82) );
  XNOR U52 ( .A(n85), .B(n80), .Z(n84) );
  AND U53 ( .A(o[2]), .B(n86), .Z(n85) );
  XNOR U54 ( .A(n87), .B(n88), .Z(n86) );
  XNOR U55 ( .A(n89), .B(n83), .Z(n88) );
  AND U56 ( .A(o[3]), .B(n90), .Z(n89) );
  XNOR U57 ( .A(n91), .B(n92), .Z(n90) );
  XNOR U58 ( .A(n93), .B(n87), .Z(n92) );
  AND U59 ( .A(o[4]), .B(n94), .Z(n93) );
  XNOR U60 ( .A(n95), .B(n96), .Z(n94) );
  XNOR U61 ( .A(n97), .B(n91), .Z(n96) );
  AND U62 ( .A(o[5]), .B(n98), .Z(n97) );
  XNOR U63 ( .A(n99), .B(n100), .Z(n98) );
  XNOR U64 ( .A(n101), .B(n95), .Z(n100) );
  AND U65 ( .A(o[6]), .B(n102), .Z(n101) );
  XNOR U66 ( .A(n99), .B(n103), .Z(n102) );
  XNOR U67 ( .A(n104), .B(n105), .Z(n103) );
  AND U68 ( .A(o[7]), .B(n106), .Z(n104) );
  XOR U69 ( .A(n105), .B(n107), .Z(n106) );
  XOR U70 ( .A(n108), .B(n109), .Z(n99) );
  AND U71 ( .A(o[7]), .B(n110), .Z(n109) );
  XOR U72 ( .A(n108), .B(n111), .Z(n110) );
  XOR U73 ( .A(n112), .B(n113), .Z(n95) );
  AND U74 ( .A(o[6]), .B(n114), .Z(n113) );
  XNOR U75 ( .A(n112), .B(n115), .Z(n114) );
  XNOR U76 ( .A(n116), .B(n117), .Z(n115) );
  AND U77 ( .A(o[7]), .B(n118), .Z(n116) );
  XOR U78 ( .A(n117), .B(n119), .Z(n118) );
  XOR U79 ( .A(n120), .B(n121), .Z(n112) );
  AND U80 ( .A(o[7]), .B(n122), .Z(n121) );
  XOR U81 ( .A(n120), .B(n123), .Z(n122) );
  XOR U82 ( .A(n124), .B(n125), .Z(n91) );
  AND U83 ( .A(o[5]), .B(n126), .Z(n125) );
  XNOR U84 ( .A(n127), .B(n128), .Z(n126) );
  XNOR U85 ( .A(n129), .B(n124), .Z(n128) );
  AND U86 ( .A(o[6]), .B(n130), .Z(n129) );
  XNOR U87 ( .A(n127), .B(n131), .Z(n130) );
  XNOR U88 ( .A(n132), .B(n133), .Z(n131) );
  AND U89 ( .A(o[7]), .B(n134), .Z(n132) );
  XOR U90 ( .A(n133), .B(n135), .Z(n134) );
  XOR U91 ( .A(n136), .B(n137), .Z(n127) );
  AND U92 ( .A(o[7]), .B(n138), .Z(n137) );
  XOR U93 ( .A(n136), .B(n139), .Z(n138) );
  XOR U94 ( .A(n140), .B(n141), .Z(n124) );
  AND U95 ( .A(o[6]), .B(n142), .Z(n141) );
  XNOR U96 ( .A(n140), .B(n143), .Z(n142) );
  XNOR U97 ( .A(n144), .B(n145), .Z(n143) );
  AND U98 ( .A(o[7]), .B(n146), .Z(n144) );
  XOR U99 ( .A(n145), .B(n147), .Z(n146) );
  XOR U100 ( .A(n148), .B(n149), .Z(n140) );
  AND U101 ( .A(o[7]), .B(n150), .Z(n149) );
  XOR U102 ( .A(n148), .B(n151), .Z(n150) );
  XOR U103 ( .A(n152), .B(n153), .Z(n87) );
  AND U104 ( .A(o[4]), .B(n154), .Z(n153) );
  XNOR U105 ( .A(n155), .B(n156), .Z(n154) );
  XNOR U106 ( .A(n157), .B(n152), .Z(n156) );
  AND U107 ( .A(o[5]), .B(n158), .Z(n157) );
  XNOR U108 ( .A(n159), .B(n160), .Z(n158) );
  XNOR U109 ( .A(n161), .B(n155), .Z(n160) );
  AND U110 ( .A(o[6]), .B(n162), .Z(n161) );
  XNOR U111 ( .A(n159), .B(n163), .Z(n162) );
  XNOR U112 ( .A(n164), .B(n165), .Z(n163) );
  AND U113 ( .A(o[7]), .B(n166), .Z(n164) );
  XOR U114 ( .A(n165), .B(n167), .Z(n166) );
  XOR U115 ( .A(n168), .B(n169), .Z(n159) );
  AND U116 ( .A(o[7]), .B(n170), .Z(n169) );
  XOR U117 ( .A(n168), .B(n171), .Z(n170) );
  XOR U118 ( .A(n172), .B(n173), .Z(n155) );
  AND U119 ( .A(o[6]), .B(n174), .Z(n173) );
  XNOR U120 ( .A(n172), .B(n175), .Z(n174) );
  XNOR U121 ( .A(n176), .B(n177), .Z(n175) );
  AND U122 ( .A(o[7]), .B(n178), .Z(n176) );
  XOR U123 ( .A(n177), .B(n179), .Z(n178) );
  XOR U124 ( .A(n180), .B(n181), .Z(n172) );
  AND U125 ( .A(o[7]), .B(n182), .Z(n181) );
  XOR U126 ( .A(n180), .B(n183), .Z(n182) );
  XOR U127 ( .A(n184), .B(n185), .Z(n152) );
  AND U128 ( .A(o[5]), .B(n186), .Z(n185) );
  XNOR U129 ( .A(n187), .B(n188), .Z(n186) );
  XNOR U130 ( .A(n189), .B(n184), .Z(n188) );
  AND U131 ( .A(o[6]), .B(n190), .Z(n189) );
  XNOR U132 ( .A(n187), .B(n191), .Z(n190) );
  XNOR U133 ( .A(n192), .B(n193), .Z(n191) );
  AND U134 ( .A(o[7]), .B(n194), .Z(n192) );
  XOR U135 ( .A(n193), .B(n195), .Z(n194) );
  XOR U136 ( .A(n196), .B(n197), .Z(n187) );
  AND U137 ( .A(o[7]), .B(n198), .Z(n197) );
  XOR U138 ( .A(n196), .B(n199), .Z(n198) );
  XOR U139 ( .A(n200), .B(n201), .Z(n184) );
  AND U140 ( .A(o[6]), .B(n202), .Z(n201) );
  XNOR U141 ( .A(n200), .B(n203), .Z(n202) );
  XNOR U142 ( .A(n204), .B(n205), .Z(n203) );
  AND U143 ( .A(o[7]), .B(n206), .Z(n204) );
  XOR U144 ( .A(n205), .B(n207), .Z(n206) );
  XOR U145 ( .A(n208), .B(n209), .Z(n200) );
  AND U146 ( .A(o[7]), .B(n210), .Z(n209) );
  XOR U147 ( .A(n208), .B(n211), .Z(n210) );
  XOR U148 ( .A(n212), .B(n213), .Z(n83) );
  AND U149 ( .A(o[3]), .B(n214), .Z(n213) );
  XNOR U150 ( .A(n215), .B(n216), .Z(n214) );
  XNOR U151 ( .A(n217), .B(n212), .Z(n216) );
  AND U152 ( .A(o[4]), .B(n218), .Z(n217) );
  XNOR U153 ( .A(n219), .B(n220), .Z(n218) );
  XNOR U154 ( .A(n221), .B(n215), .Z(n220) );
  AND U155 ( .A(o[5]), .B(n222), .Z(n221) );
  XNOR U156 ( .A(n223), .B(n224), .Z(n222) );
  XNOR U157 ( .A(n225), .B(n219), .Z(n224) );
  AND U158 ( .A(o[6]), .B(n226), .Z(n225) );
  XNOR U159 ( .A(n223), .B(n227), .Z(n226) );
  XNOR U160 ( .A(n228), .B(n229), .Z(n227) );
  AND U161 ( .A(o[7]), .B(n230), .Z(n228) );
  XOR U162 ( .A(n229), .B(n231), .Z(n230) );
  XOR U163 ( .A(n232), .B(n233), .Z(n223) );
  AND U164 ( .A(o[7]), .B(n234), .Z(n233) );
  XOR U165 ( .A(n232), .B(n235), .Z(n234) );
  XOR U166 ( .A(n236), .B(n237), .Z(n219) );
  AND U167 ( .A(o[6]), .B(n238), .Z(n237) );
  XNOR U168 ( .A(n236), .B(n239), .Z(n238) );
  XNOR U169 ( .A(n240), .B(n241), .Z(n239) );
  AND U170 ( .A(o[7]), .B(n242), .Z(n240) );
  XOR U171 ( .A(n241), .B(n243), .Z(n242) );
  XOR U172 ( .A(n244), .B(n245), .Z(n236) );
  AND U173 ( .A(o[7]), .B(n246), .Z(n245) );
  XOR U174 ( .A(n244), .B(n247), .Z(n246) );
  XOR U175 ( .A(n248), .B(n249), .Z(n215) );
  AND U176 ( .A(o[5]), .B(n250), .Z(n249) );
  XNOR U177 ( .A(n251), .B(n252), .Z(n250) );
  XNOR U178 ( .A(n253), .B(n248), .Z(n252) );
  AND U179 ( .A(o[6]), .B(n254), .Z(n253) );
  XNOR U180 ( .A(n251), .B(n255), .Z(n254) );
  XNOR U181 ( .A(n256), .B(n257), .Z(n255) );
  AND U182 ( .A(o[7]), .B(n258), .Z(n256) );
  XOR U183 ( .A(n257), .B(n259), .Z(n258) );
  XOR U184 ( .A(n260), .B(n261), .Z(n251) );
  AND U185 ( .A(o[7]), .B(n262), .Z(n261) );
  XOR U186 ( .A(n260), .B(n263), .Z(n262) );
  XOR U187 ( .A(n264), .B(n265), .Z(n248) );
  AND U188 ( .A(o[6]), .B(n266), .Z(n265) );
  XNOR U189 ( .A(n264), .B(n267), .Z(n266) );
  XNOR U190 ( .A(n268), .B(n269), .Z(n267) );
  AND U191 ( .A(o[7]), .B(n270), .Z(n268) );
  XOR U192 ( .A(n269), .B(n271), .Z(n270) );
  XOR U193 ( .A(n272), .B(n273), .Z(n264) );
  AND U194 ( .A(o[7]), .B(n274), .Z(n273) );
  XOR U195 ( .A(n272), .B(n275), .Z(n274) );
  XOR U196 ( .A(n276), .B(n277), .Z(n212) );
  AND U197 ( .A(o[4]), .B(n278), .Z(n277) );
  XNOR U198 ( .A(n279), .B(n280), .Z(n278) );
  XNOR U199 ( .A(n281), .B(n276), .Z(n280) );
  AND U200 ( .A(o[5]), .B(n282), .Z(n281) );
  XNOR U201 ( .A(n283), .B(n284), .Z(n282) );
  XNOR U202 ( .A(n285), .B(n279), .Z(n284) );
  AND U203 ( .A(o[6]), .B(n286), .Z(n285) );
  XNOR U204 ( .A(n283), .B(n287), .Z(n286) );
  XNOR U205 ( .A(n288), .B(n289), .Z(n287) );
  AND U206 ( .A(o[7]), .B(n290), .Z(n288) );
  XOR U207 ( .A(n289), .B(n291), .Z(n290) );
  XOR U208 ( .A(n292), .B(n293), .Z(n283) );
  AND U209 ( .A(o[7]), .B(n294), .Z(n293) );
  XOR U210 ( .A(n292), .B(n295), .Z(n294) );
  XOR U211 ( .A(n296), .B(n297), .Z(n279) );
  AND U212 ( .A(o[6]), .B(n298), .Z(n297) );
  XNOR U213 ( .A(n296), .B(n299), .Z(n298) );
  XNOR U214 ( .A(n300), .B(n301), .Z(n299) );
  AND U215 ( .A(o[7]), .B(n302), .Z(n300) );
  XOR U216 ( .A(n301), .B(n303), .Z(n302) );
  XOR U217 ( .A(n304), .B(n305), .Z(n296) );
  AND U218 ( .A(o[7]), .B(n306), .Z(n305) );
  XOR U219 ( .A(n304), .B(n307), .Z(n306) );
  XOR U220 ( .A(n308), .B(n309), .Z(n276) );
  AND U221 ( .A(o[5]), .B(n310), .Z(n309) );
  XNOR U222 ( .A(n311), .B(n312), .Z(n310) );
  XNOR U223 ( .A(n313), .B(n308), .Z(n312) );
  AND U224 ( .A(o[6]), .B(n314), .Z(n313) );
  XNOR U225 ( .A(n311), .B(n315), .Z(n314) );
  XNOR U226 ( .A(n316), .B(n317), .Z(n315) );
  AND U227 ( .A(o[7]), .B(n318), .Z(n316) );
  XOR U228 ( .A(n317), .B(n319), .Z(n318) );
  XOR U229 ( .A(n320), .B(n321), .Z(n311) );
  AND U230 ( .A(o[7]), .B(n322), .Z(n321) );
  XOR U231 ( .A(n320), .B(n323), .Z(n322) );
  XOR U232 ( .A(n324), .B(n325), .Z(n308) );
  AND U233 ( .A(o[6]), .B(n326), .Z(n325) );
  XNOR U234 ( .A(n324), .B(n327), .Z(n326) );
  XNOR U235 ( .A(n328), .B(n329), .Z(n327) );
  AND U236 ( .A(o[7]), .B(n330), .Z(n328) );
  XOR U237 ( .A(n329), .B(n331), .Z(n330) );
  XOR U238 ( .A(n332), .B(n333), .Z(n324) );
  AND U239 ( .A(o[7]), .B(n334), .Z(n333) );
  XOR U240 ( .A(n332), .B(n335), .Z(n334) );
  XOR U241 ( .A(n336), .B(n337), .Z(o[1]) );
  AND U242 ( .A(o[2]), .B(n338), .Z(n337) );
  XNOR U243 ( .A(n339), .B(n340), .Z(n338) );
  XNOR U244 ( .A(n341), .B(n336), .Z(n340) );
  AND U245 ( .A(o[3]), .B(n342), .Z(n341) );
  XNOR U246 ( .A(n343), .B(n344), .Z(n342) );
  XNOR U247 ( .A(n345), .B(n339), .Z(n344) );
  AND U248 ( .A(o[4]), .B(n346), .Z(n345) );
  XNOR U249 ( .A(n347), .B(n348), .Z(n346) );
  XNOR U250 ( .A(n349), .B(n343), .Z(n348) );
  AND U251 ( .A(o[5]), .B(n350), .Z(n349) );
  XNOR U252 ( .A(n351), .B(n352), .Z(n350) );
  XNOR U253 ( .A(n353), .B(n347), .Z(n352) );
  AND U254 ( .A(o[6]), .B(n354), .Z(n353) );
  XNOR U255 ( .A(n351), .B(n355), .Z(n354) );
  XNOR U256 ( .A(n356), .B(n357), .Z(n355) );
  AND U257 ( .A(o[7]), .B(n358), .Z(n356) );
  XOR U258 ( .A(n357), .B(n359), .Z(n358) );
  XOR U259 ( .A(n360), .B(n361), .Z(n351) );
  AND U260 ( .A(o[7]), .B(n362), .Z(n361) );
  XOR U261 ( .A(n360), .B(n363), .Z(n362) );
  XOR U262 ( .A(n364), .B(n365), .Z(n347) );
  AND U263 ( .A(o[6]), .B(n366), .Z(n365) );
  XNOR U264 ( .A(n364), .B(n367), .Z(n366) );
  XNOR U265 ( .A(n368), .B(n369), .Z(n367) );
  AND U266 ( .A(o[7]), .B(n370), .Z(n368) );
  XOR U267 ( .A(n369), .B(n371), .Z(n370) );
  XOR U268 ( .A(n372), .B(n373), .Z(n364) );
  AND U269 ( .A(o[7]), .B(n374), .Z(n373) );
  XOR U270 ( .A(n372), .B(n375), .Z(n374) );
  XOR U271 ( .A(n376), .B(n377), .Z(n343) );
  AND U272 ( .A(o[5]), .B(n378), .Z(n377) );
  XNOR U273 ( .A(n379), .B(n380), .Z(n378) );
  XNOR U274 ( .A(n381), .B(n376), .Z(n380) );
  AND U275 ( .A(o[6]), .B(n382), .Z(n381) );
  XNOR U276 ( .A(n379), .B(n383), .Z(n382) );
  XNOR U277 ( .A(n384), .B(n385), .Z(n383) );
  AND U278 ( .A(o[7]), .B(n386), .Z(n384) );
  XOR U279 ( .A(n385), .B(n387), .Z(n386) );
  XOR U280 ( .A(n388), .B(n389), .Z(n379) );
  AND U281 ( .A(o[7]), .B(n390), .Z(n389) );
  XOR U282 ( .A(n388), .B(n391), .Z(n390) );
  XOR U283 ( .A(n392), .B(n393), .Z(n376) );
  AND U284 ( .A(o[6]), .B(n394), .Z(n393) );
  XNOR U285 ( .A(n392), .B(n395), .Z(n394) );
  XNOR U286 ( .A(n396), .B(n397), .Z(n395) );
  AND U287 ( .A(o[7]), .B(n398), .Z(n396) );
  XOR U288 ( .A(n397), .B(n399), .Z(n398) );
  XOR U289 ( .A(n400), .B(n401), .Z(n392) );
  AND U290 ( .A(o[7]), .B(n402), .Z(n401) );
  XOR U291 ( .A(n400), .B(n403), .Z(n402) );
  XOR U292 ( .A(n404), .B(n405), .Z(n339) );
  AND U293 ( .A(o[4]), .B(n406), .Z(n405) );
  XNOR U294 ( .A(n407), .B(n408), .Z(n406) );
  XNOR U295 ( .A(n409), .B(n404), .Z(n408) );
  AND U296 ( .A(o[5]), .B(n410), .Z(n409) );
  XNOR U297 ( .A(n411), .B(n412), .Z(n410) );
  XNOR U298 ( .A(n413), .B(n407), .Z(n412) );
  AND U299 ( .A(o[6]), .B(n414), .Z(n413) );
  XNOR U300 ( .A(n411), .B(n415), .Z(n414) );
  XNOR U301 ( .A(n416), .B(n417), .Z(n415) );
  AND U302 ( .A(o[7]), .B(n418), .Z(n416) );
  XOR U303 ( .A(n417), .B(n419), .Z(n418) );
  XOR U304 ( .A(n420), .B(n421), .Z(n411) );
  AND U305 ( .A(o[7]), .B(n422), .Z(n421) );
  XOR U306 ( .A(n420), .B(n423), .Z(n422) );
  XOR U307 ( .A(n424), .B(n425), .Z(n407) );
  AND U308 ( .A(o[6]), .B(n426), .Z(n425) );
  XNOR U309 ( .A(n424), .B(n427), .Z(n426) );
  XNOR U310 ( .A(n428), .B(n429), .Z(n427) );
  AND U311 ( .A(o[7]), .B(n430), .Z(n428) );
  XOR U312 ( .A(n429), .B(n431), .Z(n430) );
  XOR U313 ( .A(n432), .B(n433), .Z(n424) );
  AND U314 ( .A(o[7]), .B(n434), .Z(n433) );
  XOR U315 ( .A(n432), .B(n435), .Z(n434) );
  XOR U316 ( .A(n436), .B(n437), .Z(n404) );
  AND U317 ( .A(o[5]), .B(n438), .Z(n437) );
  XNOR U318 ( .A(n439), .B(n440), .Z(n438) );
  XNOR U319 ( .A(n441), .B(n436), .Z(n440) );
  AND U320 ( .A(o[6]), .B(n442), .Z(n441) );
  XNOR U321 ( .A(n439), .B(n443), .Z(n442) );
  XNOR U322 ( .A(n444), .B(n445), .Z(n443) );
  AND U323 ( .A(o[7]), .B(n446), .Z(n444) );
  XOR U324 ( .A(n445), .B(n447), .Z(n446) );
  XOR U325 ( .A(n448), .B(n449), .Z(n439) );
  AND U326 ( .A(o[7]), .B(n450), .Z(n449) );
  XOR U327 ( .A(n448), .B(n451), .Z(n450) );
  XOR U328 ( .A(n452), .B(n453), .Z(n436) );
  AND U329 ( .A(o[6]), .B(n454), .Z(n453) );
  XNOR U330 ( .A(n452), .B(n455), .Z(n454) );
  XNOR U331 ( .A(n456), .B(n457), .Z(n455) );
  AND U332 ( .A(o[7]), .B(n458), .Z(n456) );
  XOR U333 ( .A(n457), .B(n459), .Z(n458) );
  XOR U334 ( .A(n460), .B(n461), .Z(n452) );
  AND U335 ( .A(o[7]), .B(n462), .Z(n461) );
  XOR U336 ( .A(n460), .B(n463), .Z(n462) );
  XOR U337 ( .A(n464), .B(n465), .Z(n336) );
  AND U338 ( .A(o[3]), .B(n466), .Z(n465) );
  XNOR U339 ( .A(n467), .B(n468), .Z(n466) );
  XNOR U340 ( .A(n469), .B(n464), .Z(n468) );
  AND U341 ( .A(o[4]), .B(n470), .Z(n469) );
  XNOR U342 ( .A(n471), .B(n472), .Z(n470) );
  XNOR U343 ( .A(n473), .B(n467), .Z(n472) );
  AND U344 ( .A(o[5]), .B(n474), .Z(n473) );
  XNOR U345 ( .A(n475), .B(n476), .Z(n474) );
  XNOR U346 ( .A(n477), .B(n471), .Z(n476) );
  AND U347 ( .A(o[6]), .B(n478), .Z(n477) );
  XNOR U348 ( .A(n475), .B(n479), .Z(n478) );
  XNOR U349 ( .A(n480), .B(n481), .Z(n479) );
  AND U350 ( .A(o[7]), .B(n482), .Z(n480) );
  XOR U351 ( .A(n481), .B(n483), .Z(n482) );
  XOR U352 ( .A(n484), .B(n485), .Z(n475) );
  AND U353 ( .A(o[7]), .B(n486), .Z(n485) );
  XOR U354 ( .A(n484), .B(n487), .Z(n486) );
  XOR U355 ( .A(n488), .B(n489), .Z(n471) );
  AND U356 ( .A(o[6]), .B(n490), .Z(n489) );
  XNOR U357 ( .A(n488), .B(n491), .Z(n490) );
  XNOR U358 ( .A(n492), .B(n493), .Z(n491) );
  AND U359 ( .A(o[7]), .B(n494), .Z(n492) );
  XOR U360 ( .A(n493), .B(n495), .Z(n494) );
  XOR U361 ( .A(n496), .B(n497), .Z(n488) );
  AND U362 ( .A(o[7]), .B(n498), .Z(n497) );
  XOR U363 ( .A(n496), .B(n499), .Z(n498) );
  XOR U364 ( .A(n500), .B(n501), .Z(n467) );
  AND U365 ( .A(o[5]), .B(n502), .Z(n501) );
  XNOR U366 ( .A(n503), .B(n504), .Z(n502) );
  XNOR U367 ( .A(n505), .B(n500), .Z(n504) );
  AND U368 ( .A(o[6]), .B(n506), .Z(n505) );
  XNOR U369 ( .A(n503), .B(n507), .Z(n506) );
  XNOR U370 ( .A(n508), .B(n509), .Z(n507) );
  AND U371 ( .A(o[7]), .B(n510), .Z(n508) );
  XOR U372 ( .A(n509), .B(n511), .Z(n510) );
  XOR U373 ( .A(n512), .B(n513), .Z(n503) );
  AND U374 ( .A(o[7]), .B(n514), .Z(n513) );
  XOR U375 ( .A(n512), .B(n515), .Z(n514) );
  XOR U376 ( .A(n516), .B(n517), .Z(n500) );
  AND U377 ( .A(o[6]), .B(n518), .Z(n517) );
  XNOR U378 ( .A(n516), .B(n519), .Z(n518) );
  XNOR U379 ( .A(n520), .B(n521), .Z(n519) );
  AND U380 ( .A(o[7]), .B(n522), .Z(n520) );
  XOR U381 ( .A(n521), .B(n523), .Z(n522) );
  XOR U382 ( .A(n524), .B(n525), .Z(n516) );
  AND U383 ( .A(o[7]), .B(n526), .Z(n525) );
  XOR U384 ( .A(n524), .B(n527), .Z(n526) );
  XOR U385 ( .A(n528), .B(n529), .Z(n464) );
  AND U386 ( .A(o[4]), .B(n530), .Z(n529) );
  XNOR U387 ( .A(n531), .B(n532), .Z(n530) );
  XNOR U388 ( .A(n533), .B(n528), .Z(n532) );
  AND U389 ( .A(o[5]), .B(n534), .Z(n533) );
  XNOR U390 ( .A(n535), .B(n536), .Z(n534) );
  XNOR U391 ( .A(n537), .B(n531), .Z(n536) );
  AND U392 ( .A(o[6]), .B(n538), .Z(n537) );
  XNOR U393 ( .A(n535), .B(n539), .Z(n538) );
  XNOR U394 ( .A(n540), .B(n541), .Z(n539) );
  AND U395 ( .A(o[7]), .B(n542), .Z(n540) );
  XOR U396 ( .A(n541), .B(n543), .Z(n542) );
  XOR U397 ( .A(n544), .B(n545), .Z(n535) );
  AND U398 ( .A(o[7]), .B(n546), .Z(n545) );
  XOR U399 ( .A(n544), .B(n547), .Z(n546) );
  XOR U400 ( .A(n548), .B(n549), .Z(n531) );
  AND U401 ( .A(o[6]), .B(n550), .Z(n549) );
  XNOR U402 ( .A(n548), .B(n551), .Z(n550) );
  XNOR U403 ( .A(n552), .B(n553), .Z(n551) );
  AND U404 ( .A(o[7]), .B(n554), .Z(n552) );
  XOR U405 ( .A(n553), .B(n555), .Z(n554) );
  XOR U406 ( .A(n556), .B(n557), .Z(n548) );
  AND U407 ( .A(o[7]), .B(n558), .Z(n557) );
  XOR U408 ( .A(n556), .B(n559), .Z(n558) );
  XOR U409 ( .A(n560), .B(n561), .Z(n528) );
  AND U410 ( .A(o[5]), .B(n562), .Z(n561) );
  XNOR U411 ( .A(n563), .B(n564), .Z(n562) );
  XNOR U412 ( .A(n565), .B(n560), .Z(n564) );
  AND U413 ( .A(o[6]), .B(n566), .Z(n565) );
  XNOR U414 ( .A(n563), .B(n567), .Z(n566) );
  XNOR U415 ( .A(n568), .B(n569), .Z(n567) );
  AND U416 ( .A(o[7]), .B(n570), .Z(n568) );
  XOR U417 ( .A(n569), .B(n571), .Z(n570) );
  XOR U418 ( .A(n572), .B(n573), .Z(n563) );
  AND U419 ( .A(o[7]), .B(n574), .Z(n573) );
  XOR U420 ( .A(n572), .B(n575), .Z(n574) );
  XOR U421 ( .A(n576), .B(n577), .Z(n560) );
  AND U422 ( .A(o[6]), .B(n578), .Z(n577) );
  XNOR U423 ( .A(n576), .B(n579), .Z(n578) );
  XNOR U424 ( .A(n580), .B(n581), .Z(n579) );
  AND U425 ( .A(o[7]), .B(n582), .Z(n580) );
  XOR U426 ( .A(n581), .B(n583), .Z(n582) );
  XOR U427 ( .A(n584), .B(n585), .Z(n576) );
  AND U428 ( .A(o[7]), .B(n586), .Z(n585) );
  XOR U429 ( .A(n584), .B(n587), .Z(n586) );
  XOR U430 ( .A(n588), .B(n589), .Z(n80) );
  AND U431 ( .A(o[2]), .B(n590), .Z(n589) );
  XNOR U432 ( .A(n591), .B(n592), .Z(n590) );
  XNOR U433 ( .A(n593), .B(n588), .Z(n592) );
  AND U434 ( .A(o[3]), .B(n594), .Z(n593) );
  XNOR U435 ( .A(n595), .B(n596), .Z(n594) );
  XNOR U436 ( .A(n597), .B(n591), .Z(n596) );
  AND U437 ( .A(o[4]), .B(n598), .Z(n597) );
  XNOR U438 ( .A(n599), .B(n600), .Z(n598) );
  XNOR U439 ( .A(n601), .B(n595), .Z(n600) );
  AND U440 ( .A(o[5]), .B(n602), .Z(n601) );
  XNOR U441 ( .A(n603), .B(n604), .Z(n602) );
  XNOR U442 ( .A(n605), .B(n599), .Z(n604) );
  AND U443 ( .A(o[6]), .B(n606), .Z(n605) );
  XNOR U444 ( .A(n603), .B(n607), .Z(n606) );
  XNOR U445 ( .A(n608), .B(n609), .Z(n607) );
  AND U446 ( .A(o[7]), .B(n610), .Z(n608) );
  XOR U447 ( .A(n609), .B(n611), .Z(n610) );
  XOR U448 ( .A(n612), .B(n613), .Z(n603) );
  AND U449 ( .A(o[7]), .B(n614), .Z(n613) );
  XOR U450 ( .A(n612), .B(n615), .Z(n614) );
  XOR U451 ( .A(n616), .B(n617), .Z(n599) );
  AND U452 ( .A(o[6]), .B(n618), .Z(n617) );
  XNOR U453 ( .A(n616), .B(n619), .Z(n618) );
  XNOR U454 ( .A(n620), .B(n621), .Z(n619) );
  AND U455 ( .A(o[7]), .B(n622), .Z(n620) );
  XOR U456 ( .A(n621), .B(n623), .Z(n622) );
  XOR U457 ( .A(n624), .B(n625), .Z(n616) );
  AND U458 ( .A(o[7]), .B(n626), .Z(n625) );
  XOR U459 ( .A(n624), .B(n627), .Z(n626) );
  XOR U460 ( .A(n628), .B(n629), .Z(n595) );
  AND U461 ( .A(o[5]), .B(n630), .Z(n629) );
  XNOR U462 ( .A(n631), .B(n632), .Z(n630) );
  XNOR U463 ( .A(n633), .B(n628), .Z(n632) );
  AND U464 ( .A(o[6]), .B(n634), .Z(n633) );
  XNOR U465 ( .A(n631), .B(n635), .Z(n634) );
  XNOR U466 ( .A(n636), .B(n637), .Z(n635) );
  AND U467 ( .A(o[7]), .B(n638), .Z(n636) );
  XOR U468 ( .A(n637), .B(n639), .Z(n638) );
  XOR U469 ( .A(n640), .B(n641), .Z(n631) );
  AND U470 ( .A(o[7]), .B(n642), .Z(n641) );
  XOR U471 ( .A(n640), .B(n643), .Z(n642) );
  XOR U472 ( .A(n644), .B(n645), .Z(n628) );
  AND U473 ( .A(o[6]), .B(n646), .Z(n645) );
  XNOR U474 ( .A(n644), .B(n647), .Z(n646) );
  XNOR U475 ( .A(n648), .B(n649), .Z(n647) );
  AND U476 ( .A(o[7]), .B(n650), .Z(n648) );
  XOR U477 ( .A(n649), .B(n651), .Z(n650) );
  XOR U478 ( .A(n652), .B(n653), .Z(n644) );
  AND U479 ( .A(o[7]), .B(n654), .Z(n653) );
  XOR U480 ( .A(n652), .B(n655), .Z(n654) );
  XOR U481 ( .A(n656), .B(n657), .Z(n591) );
  AND U482 ( .A(o[4]), .B(n658), .Z(n657) );
  XNOR U483 ( .A(n659), .B(n660), .Z(n658) );
  XNOR U484 ( .A(n661), .B(n656), .Z(n660) );
  AND U485 ( .A(o[5]), .B(n662), .Z(n661) );
  XNOR U486 ( .A(n663), .B(n664), .Z(n662) );
  XNOR U487 ( .A(n665), .B(n659), .Z(n664) );
  AND U488 ( .A(o[6]), .B(n666), .Z(n665) );
  XNOR U489 ( .A(n663), .B(n667), .Z(n666) );
  XNOR U490 ( .A(n668), .B(n669), .Z(n667) );
  AND U491 ( .A(o[7]), .B(n670), .Z(n668) );
  XOR U492 ( .A(n669), .B(n671), .Z(n670) );
  XOR U493 ( .A(n672), .B(n673), .Z(n663) );
  AND U494 ( .A(o[7]), .B(n674), .Z(n673) );
  XOR U495 ( .A(n672), .B(n675), .Z(n674) );
  XOR U496 ( .A(n676), .B(n677), .Z(n659) );
  AND U497 ( .A(o[6]), .B(n678), .Z(n677) );
  XNOR U498 ( .A(n676), .B(n679), .Z(n678) );
  XNOR U499 ( .A(n680), .B(n681), .Z(n679) );
  AND U500 ( .A(o[7]), .B(n682), .Z(n680) );
  XOR U501 ( .A(n681), .B(n683), .Z(n682) );
  XOR U502 ( .A(n684), .B(n685), .Z(n676) );
  AND U503 ( .A(o[7]), .B(n686), .Z(n685) );
  XOR U504 ( .A(n684), .B(n687), .Z(n686) );
  XOR U505 ( .A(n688), .B(n689), .Z(n656) );
  AND U506 ( .A(o[5]), .B(n690), .Z(n689) );
  XNOR U507 ( .A(n691), .B(n692), .Z(n690) );
  XNOR U508 ( .A(n693), .B(n688), .Z(n692) );
  AND U509 ( .A(o[6]), .B(n694), .Z(n693) );
  XNOR U510 ( .A(n691), .B(n695), .Z(n694) );
  XNOR U511 ( .A(n696), .B(n697), .Z(n695) );
  AND U512 ( .A(o[7]), .B(n698), .Z(n696) );
  XOR U513 ( .A(n697), .B(n699), .Z(n698) );
  XOR U514 ( .A(n700), .B(n701), .Z(n691) );
  AND U515 ( .A(o[7]), .B(n702), .Z(n701) );
  XOR U516 ( .A(n700), .B(n703), .Z(n702) );
  XOR U517 ( .A(n704), .B(n705), .Z(n688) );
  AND U518 ( .A(o[6]), .B(n706), .Z(n705) );
  XNOR U519 ( .A(n704), .B(n707), .Z(n706) );
  XNOR U520 ( .A(n708), .B(n709), .Z(n707) );
  AND U521 ( .A(o[7]), .B(n710), .Z(n708) );
  XOR U522 ( .A(n709), .B(n711), .Z(n710) );
  XOR U523 ( .A(n712), .B(n713), .Z(n704) );
  AND U524 ( .A(o[7]), .B(n714), .Z(n713) );
  XOR U525 ( .A(n712), .B(n715), .Z(n714) );
  XOR U526 ( .A(n716), .B(n717), .Z(o[2]) );
  AND U527 ( .A(o[3]), .B(n718), .Z(n717) );
  XNOR U528 ( .A(n719), .B(n720), .Z(n718) );
  XNOR U529 ( .A(n721), .B(n716), .Z(n720) );
  AND U530 ( .A(o[4]), .B(n722), .Z(n721) );
  XNOR U531 ( .A(n723), .B(n724), .Z(n722) );
  XNOR U532 ( .A(n725), .B(n719), .Z(n724) );
  AND U533 ( .A(o[5]), .B(n726), .Z(n725) );
  XNOR U534 ( .A(n727), .B(n728), .Z(n726) );
  XNOR U535 ( .A(n729), .B(n723), .Z(n728) );
  AND U536 ( .A(o[6]), .B(n730), .Z(n729) );
  XNOR U537 ( .A(n727), .B(n731), .Z(n730) );
  XNOR U538 ( .A(n732), .B(n733), .Z(n731) );
  AND U539 ( .A(o[7]), .B(n734), .Z(n732) );
  XOR U540 ( .A(n733), .B(n735), .Z(n734) );
  XOR U541 ( .A(n736), .B(n737), .Z(n727) );
  AND U542 ( .A(o[7]), .B(n738), .Z(n737) );
  XOR U543 ( .A(n736), .B(n739), .Z(n738) );
  XOR U544 ( .A(n740), .B(n741), .Z(n723) );
  AND U545 ( .A(o[6]), .B(n742), .Z(n741) );
  XNOR U546 ( .A(n740), .B(n743), .Z(n742) );
  XNOR U547 ( .A(n744), .B(n745), .Z(n743) );
  AND U548 ( .A(o[7]), .B(n746), .Z(n744) );
  XOR U549 ( .A(n745), .B(n747), .Z(n746) );
  XOR U550 ( .A(n748), .B(n749), .Z(n740) );
  AND U551 ( .A(o[7]), .B(n750), .Z(n749) );
  XOR U552 ( .A(n748), .B(n751), .Z(n750) );
  XOR U553 ( .A(n752), .B(n753), .Z(n719) );
  AND U554 ( .A(o[5]), .B(n754), .Z(n753) );
  XNOR U555 ( .A(n755), .B(n756), .Z(n754) );
  XNOR U556 ( .A(n757), .B(n752), .Z(n756) );
  AND U557 ( .A(o[6]), .B(n758), .Z(n757) );
  XNOR U558 ( .A(n755), .B(n759), .Z(n758) );
  XNOR U559 ( .A(n760), .B(n761), .Z(n759) );
  AND U560 ( .A(o[7]), .B(n762), .Z(n760) );
  XOR U561 ( .A(n761), .B(n763), .Z(n762) );
  XOR U562 ( .A(n764), .B(n765), .Z(n755) );
  AND U563 ( .A(o[7]), .B(n766), .Z(n765) );
  XOR U564 ( .A(n764), .B(n767), .Z(n766) );
  XOR U565 ( .A(n768), .B(n769), .Z(n752) );
  AND U566 ( .A(o[6]), .B(n770), .Z(n769) );
  XNOR U567 ( .A(n768), .B(n771), .Z(n770) );
  XNOR U568 ( .A(n772), .B(n773), .Z(n771) );
  AND U569 ( .A(o[7]), .B(n774), .Z(n772) );
  XOR U570 ( .A(n773), .B(n775), .Z(n774) );
  XOR U571 ( .A(n776), .B(n777), .Z(n768) );
  AND U572 ( .A(o[7]), .B(n778), .Z(n777) );
  XOR U573 ( .A(n776), .B(n779), .Z(n778) );
  XOR U574 ( .A(n780), .B(n781), .Z(n716) );
  AND U575 ( .A(o[4]), .B(n782), .Z(n781) );
  XNOR U576 ( .A(n783), .B(n784), .Z(n782) );
  XNOR U577 ( .A(n785), .B(n780), .Z(n784) );
  AND U578 ( .A(o[5]), .B(n786), .Z(n785) );
  XNOR U579 ( .A(n787), .B(n788), .Z(n786) );
  XNOR U580 ( .A(n789), .B(n783), .Z(n788) );
  AND U581 ( .A(o[6]), .B(n790), .Z(n789) );
  XNOR U582 ( .A(n787), .B(n791), .Z(n790) );
  XNOR U583 ( .A(n792), .B(n793), .Z(n791) );
  AND U584 ( .A(o[7]), .B(n794), .Z(n792) );
  XOR U585 ( .A(n793), .B(n795), .Z(n794) );
  XOR U586 ( .A(n796), .B(n797), .Z(n787) );
  AND U587 ( .A(o[7]), .B(n798), .Z(n797) );
  XOR U588 ( .A(n796), .B(n799), .Z(n798) );
  XOR U589 ( .A(n800), .B(n801), .Z(n783) );
  AND U590 ( .A(o[6]), .B(n802), .Z(n801) );
  XNOR U591 ( .A(n800), .B(n803), .Z(n802) );
  XNOR U592 ( .A(n804), .B(n805), .Z(n803) );
  AND U593 ( .A(o[7]), .B(n806), .Z(n804) );
  XOR U594 ( .A(n805), .B(n807), .Z(n806) );
  XOR U595 ( .A(n808), .B(n809), .Z(n800) );
  AND U596 ( .A(o[7]), .B(n810), .Z(n809) );
  XOR U597 ( .A(n808), .B(n811), .Z(n810) );
  XOR U598 ( .A(n812), .B(n813), .Z(n780) );
  AND U599 ( .A(o[5]), .B(n814), .Z(n813) );
  XNOR U600 ( .A(n815), .B(n816), .Z(n814) );
  XNOR U601 ( .A(n817), .B(n812), .Z(n816) );
  AND U602 ( .A(o[6]), .B(n818), .Z(n817) );
  XNOR U603 ( .A(n815), .B(n819), .Z(n818) );
  XNOR U604 ( .A(n820), .B(n821), .Z(n819) );
  AND U605 ( .A(o[7]), .B(n822), .Z(n820) );
  XOR U606 ( .A(n821), .B(n823), .Z(n822) );
  XOR U607 ( .A(n824), .B(n825), .Z(n815) );
  AND U608 ( .A(o[7]), .B(n826), .Z(n825) );
  XOR U609 ( .A(n824), .B(n827), .Z(n826) );
  XOR U610 ( .A(n828), .B(n829), .Z(n812) );
  AND U611 ( .A(o[6]), .B(n830), .Z(n829) );
  XNOR U612 ( .A(n828), .B(n831), .Z(n830) );
  XNOR U613 ( .A(n832), .B(n833), .Z(n831) );
  AND U614 ( .A(o[7]), .B(n834), .Z(n832) );
  XOR U615 ( .A(n833), .B(n835), .Z(n834) );
  XOR U616 ( .A(n836), .B(n837), .Z(n828) );
  AND U617 ( .A(o[7]), .B(n838), .Z(n837) );
  XOR U618 ( .A(n836), .B(n839), .Z(n838) );
  XOR U619 ( .A(n840), .B(n841), .Z(n588) );
  AND U620 ( .A(o[3]), .B(n842), .Z(n841) );
  XNOR U621 ( .A(n843), .B(n844), .Z(n842) );
  XNOR U622 ( .A(n845), .B(n840), .Z(n844) );
  AND U623 ( .A(o[4]), .B(n846), .Z(n845) );
  XNOR U624 ( .A(n847), .B(n848), .Z(n846) );
  XNOR U625 ( .A(n849), .B(n843), .Z(n848) );
  AND U626 ( .A(o[5]), .B(n850), .Z(n849) );
  XNOR U627 ( .A(n851), .B(n852), .Z(n850) );
  XNOR U628 ( .A(n853), .B(n847), .Z(n852) );
  AND U629 ( .A(o[6]), .B(n854), .Z(n853) );
  XNOR U630 ( .A(n851), .B(n855), .Z(n854) );
  XNOR U631 ( .A(n856), .B(n857), .Z(n855) );
  AND U632 ( .A(o[7]), .B(n858), .Z(n856) );
  XOR U633 ( .A(n857), .B(n859), .Z(n858) );
  XOR U634 ( .A(n860), .B(n861), .Z(n851) );
  AND U635 ( .A(o[7]), .B(n862), .Z(n861) );
  XOR U636 ( .A(n860), .B(n863), .Z(n862) );
  XOR U637 ( .A(n864), .B(n865), .Z(n847) );
  AND U638 ( .A(o[6]), .B(n866), .Z(n865) );
  XNOR U639 ( .A(n864), .B(n867), .Z(n866) );
  XNOR U640 ( .A(n868), .B(n869), .Z(n867) );
  AND U641 ( .A(o[7]), .B(n870), .Z(n868) );
  XOR U642 ( .A(n869), .B(n871), .Z(n870) );
  XOR U643 ( .A(n872), .B(n873), .Z(n864) );
  AND U644 ( .A(o[7]), .B(n874), .Z(n873) );
  XOR U645 ( .A(n872), .B(n875), .Z(n874) );
  XOR U646 ( .A(n876), .B(n877), .Z(n843) );
  AND U647 ( .A(o[5]), .B(n878), .Z(n877) );
  XNOR U648 ( .A(n879), .B(n880), .Z(n878) );
  XNOR U649 ( .A(n881), .B(n876), .Z(n880) );
  AND U650 ( .A(o[6]), .B(n882), .Z(n881) );
  XNOR U651 ( .A(n879), .B(n883), .Z(n882) );
  XNOR U652 ( .A(n884), .B(n885), .Z(n883) );
  AND U653 ( .A(o[7]), .B(n886), .Z(n884) );
  XOR U654 ( .A(n885), .B(n887), .Z(n886) );
  XOR U655 ( .A(n888), .B(n889), .Z(n879) );
  AND U656 ( .A(o[7]), .B(n890), .Z(n889) );
  XOR U657 ( .A(n888), .B(n891), .Z(n890) );
  XOR U658 ( .A(n892), .B(n893), .Z(n876) );
  AND U659 ( .A(o[6]), .B(n894), .Z(n893) );
  XNOR U660 ( .A(n892), .B(n895), .Z(n894) );
  XNOR U661 ( .A(n896), .B(n897), .Z(n895) );
  AND U662 ( .A(o[7]), .B(n898), .Z(n896) );
  XOR U663 ( .A(n897), .B(n899), .Z(n898) );
  XOR U664 ( .A(n900), .B(n901), .Z(n892) );
  AND U665 ( .A(o[7]), .B(n902), .Z(n901) );
  XOR U666 ( .A(n900), .B(n903), .Z(n902) );
  XOR U667 ( .A(n904), .B(n905), .Z(o[3]) );
  AND U668 ( .A(o[4]), .B(n906), .Z(n905) );
  XNOR U669 ( .A(n907), .B(n908), .Z(n906) );
  XNOR U670 ( .A(n909), .B(n904), .Z(n908) );
  AND U671 ( .A(o[5]), .B(n910), .Z(n909) );
  XNOR U672 ( .A(n911), .B(n912), .Z(n910) );
  XNOR U673 ( .A(n913), .B(n907), .Z(n912) );
  AND U674 ( .A(o[6]), .B(n914), .Z(n913) );
  XNOR U675 ( .A(n911), .B(n915), .Z(n914) );
  XNOR U676 ( .A(n916), .B(n917), .Z(n915) );
  AND U677 ( .A(o[7]), .B(n918), .Z(n916) );
  XOR U678 ( .A(n917), .B(n919), .Z(n918) );
  XOR U679 ( .A(n920), .B(n921), .Z(n911) );
  AND U680 ( .A(o[7]), .B(n922), .Z(n921) );
  XOR U681 ( .A(n920), .B(n923), .Z(n922) );
  XOR U682 ( .A(n924), .B(n925), .Z(n907) );
  AND U683 ( .A(o[6]), .B(n926), .Z(n925) );
  XNOR U684 ( .A(n924), .B(n927), .Z(n926) );
  XNOR U685 ( .A(n928), .B(n929), .Z(n927) );
  AND U686 ( .A(o[7]), .B(n930), .Z(n928) );
  XOR U687 ( .A(n929), .B(n931), .Z(n930) );
  XOR U688 ( .A(n932), .B(n933), .Z(n924) );
  AND U689 ( .A(o[7]), .B(n934), .Z(n933) );
  XOR U690 ( .A(n932), .B(n935), .Z(n934) );
  XOR U691 ( .A(n936), .B(n937), .Z(n904) );
  AND U692 ( .A(o[5]), .B(n938), .Z(n937) );
  XNOR U693 ( .A(n939), .B(n940), .Z(n938) );
  XNOR U694 ( .A(n941), .B(n936), .Z(n940) );
  AND U695 ( .A(o[6]), .B(n942), .Z(n941) );
  XNOR U696 ( .A(n939), .B(n943), .Z(n942) );
  XNOR U697 ( .A(n944), .B(n945), .Z(n943) );
  AND U698 ( .A(o[7]), .B(n946), .Z(n944) );
  XOR U699 ( .A(n945), .B(n947), .Z(n946) );
  XOR U700 ( .A(n948), .B(n949), .Z(n939) );
  AND U701 ( .A(o[7]), .B(n950), .Z(n949) );
  XOR U702 ( .A(n948), .B(n951), .Z(n950) );
  XOR U703 ( .A(n952), .B(n953), .Z(n936) );
  AND U704 ( .A(o[6]), .B(n954), .Z(n953) );
  XNOR U705 ( .A(n952), .B(n955), .Z(n954) );
  XNOR U706 ( .A(n956), .B(n957), .Z(n955) );
  AND U707 ( .A(o[7]), .B(n958), .Z(n956) );
  XOR U708 ( .A(n957), .B(n959), .Z(n958) );
  XOR U709 ( .A(n960), .B(n961), .Z(n952) );
  AND U710 ( .A(o[7]), .B(n962), .Z(n961) );
  XOR U711 ( .A(n960), .B(n963), .Z(n962) );
  XOR U712 ( .A(n964), .B(n965), .Z(n840) );
  AND U713 ( .A(o[4]), .B(n966), .Z(n965) );
  XNOR U714 ( .A(n967), .B(n968), .Z(n966) );
  XNOR U715 ( .A(n969), .B(n964), .Z(n968) );
  AND U716 ( .A(o[5]), .B(n970), .Z(n969) );
  XNOR U717 ( .A(n971), .B(n972), .Z(n970) );
  XNOR U718 ( .A(n973), .B(n967), .Z(n972) );
  AND U719 ( .A(o[6]), .B(n974), .Z(n973) );
  XNOR U720 ( .A(n971), .B(n975), .Z(n974) );
  XNOR U721 ( .A(n976), .B(n977), .Z(n975) );
  AND U722 ( .A(o[7]), .B(n978), .Z(n976) );
  XOR U723 ( .A(n977), .B(n979), .Z(n978) );
  XOR U724 ( .A(n980), .B(n981), .Z(n971) );
  AND U725 ( .A(o[7]), .B(n982), .Z(n981) );
  XOR U726 ( .A(n980), .B(n983), .Z(n982) );
  XOR U727 ( .A(n984), .B(n985), .Z(n967) );
  AND U728 ( .A(o[6]), .B(n986), .Z(n985) );
  XNOR U729 ( .A(n984), .B(n987), .Z(n986) );
  XNOR U730 ( .A(n988), .B(n989), .Z(n987) );
  AND U731 ( .A(o[7]), .B(n990), .Z(n988) );
  XOR U732 ( .A(n989), .B(n991), .Z(n990) );
  XOR U733 ( .A(n992), .B(n993), .Z(n984) );
  AND U734 ( .A(o[7]), .B(n994), .Z(n993) );
  XOR U735 ( .A(n992), .B(n995), .Z(n994) );
  XOR U736 ( .A(n996), .B(n997), .Z(o[4]) );
  AND U737 ( .A(o[5]), .B(n998), .Z(n997) );
  XNOR U738 ( .A(n999), .B(n1000), .Z(n998) );
  XNOR U739 ( .A(n1001), .B(n996), .Z(n1000) );
  AND U740 ( .A(o[6]), .B(n1002), .Z(n1001) );
  XNOR U741 ( .A(n999), .B(n1003), .Z(n1002) );
  XNOR U742 ( .A(n1004), .B(n1005), .Z(n1003) );
  AND U743 ( .A(o[7]), .B(n1006), .Z(n1004) );
  XOR U744 ( .A(n1005), .B(n1007), .Z(n1006) );
  XOR U745 ( .A(n1008), .B(n1009), .Z(n999) );
  AND U746 ( .A(o[7]), .B(n1010), .Z(n1009) );
  XOR U747 ( .A(n1008), .B(n1011), .Z(n1010) );
  XOR U748 ( .A(n1012), .B(n1013), .Z(n996) );
  AND U749 ( .A(o[6]), .B(n1014), .Z(n1013) );
  XNOR U750 ( .A(n1012), .B(n1015), .Z(n1014) );
  XNOR U751 ( .A(n1016), .B(n1017), .Z(n1015) );
  AND U752 ( .A(o[7]), .B(n1018), .Z(n1016) );
  XOR U753 ( .A(n1017), .B(n1019), .Z(n1018) );
  XOR U754 ( .A(n1020), .B(n1021), .Z(n1012) );
  AND U755 ( .A(o[7]), .B(n1022), .Z(n1021) );
  XOR U756 ( .A(n1020), .B(n1023), .Z(n1022) );
  XOR U757 ( .A(n1024), .B(n1025), .Z(n964) );
  AND U758 ( .A(o[5]), .B(n1026), .Z(n1025) );
  XNOR U759 ( .A(n1027), .B(n1028), .Z(n1026) );
  XNOR U760 ( .A(n1029), .B(n1024), .Z(n1028) );
  AND U761 ( .A(o[6]), .B(n1030), .Z(n1029) );
  XNOR U762 ( .A(n1027), .B(n1031), .Z(n1030) );
  XNOR U763 ( .A(n1032), .B(n1033), .Z(n1031) );
  AND U764 ( .A(o[7]), .B(n1034), .Z(n1032) );
  XOR U765 ( .A(n1033), .B(n1035), .Z(n1034) );
  XOR U766 ( .A(n1036), .B(n1037), .Z(n1027) );
  AND U767 ( .A(o[7]), .B(n1038), .Z(n1037) );
  XOR U768 ( .A(n1036), .B(n1039), .Z(n1038) );
  XOR U769 ( .A(n1040), .B(n1041), .Z(o[5]) );
  AND U770 ( .A(o[6]), .B(n1042), .Z(n1041) );
  XNOR U771 ( .A(n1040), .B(n1043), .Z(n1042) );
  XNOR U772 ( .A(n1044), .B(n1045), .Z(n1043) );
  AND U773 ( .A(o[7]), .B(n1046), .Z(n1044) );
  XOR U774 ( .A(n1045), .B(n1047), .Z(n1046) );
  XOR U775 ( .A(n1048), .B(n1049), .Z(n1040) );
  AND U776 ( .A(o[7]), .B(n1050), .Z(n1049) );
  XOR U777 ( .A(n1048), .B(n1051), .Z(n1050) );
  XOR U778 ( .A(n1052), .B(n1053), .Z(n1024) );
  AND U779 ( .A(o[6]), .B(n1054), .Z(n1053) );
  XNOR U780 ( .A(n1052), .B(n1055), .Z(n1054) );
  XNOR U781 ( .A(n1056), .B(n1057), .Z(n1055) );
  AND U782 ( .A(o[7]), .B(n1058), .Z(n1056) );
  XOR U783 ( .A(n1057), .B(n1059), .Z(n1058) );
  XOR U784 ( .A(n1060), .B(n1061), .Z(o[6]) );
  AND U785 ( .A(o[7]), .B(n1062), .Z(n1061) );
  XOR U786 ( .A(n1060), .B(n1063), .Z(n1062) );
  XOR U787 ( .A(n1064), .B(n1065), .Z(n1052) );
  AND U788 ( .A(o[7]), .B(n1066), .Z(n1065) );
  XOR U789 ( .A(n1064), .B(n1067), .Z(n1066) );
  XOR U790 ( .A(n1068), .B(n1069), .Z(o[7]) );
  AND U791 ( .A(n1070), .B(n1071), .Z(n1069) );
  XOR U792 ( .A(n1068), .B(n13), .Z(n1071) );
  XOR U793 ( .A(n1072), .B(n1073), .Z(n13) );
  AND U794 ( .A(n1063), .B(n1074), .Z(n1073) );
  XOR U795 ( .A(n1075), .B(n1072), .Z(n1074) );
  XNOR U796 ( .A(n14), .B(n1068), .Z(n1070) );
  IV U797 ( .A(n11), .Z(n14) );
  XNOR U798 ( .A(n1076), .B(n1077), .Z(n11) );
  AND U799 ( .A(n1060), .B(n1078), .Z(n1077) );
  XOR U800 ( .A(n1079), .B(n1076), .Z(n1078) );
  XOR U801 ( .A(n1080), .B(n1081), .Z(n1068) );
  AND U802 ( .A(n1082), .B(n1083), .Z(n1081) );
  XOR U803 ( .A(n1080), .B(n18), .Z(n1083) );
  XOR U804 ( .A(n1084), .B(n1085), .Z(n18) );
  AND U805 ( .A(n1063), .B(n1086), .Z(n1085) );
  XOR U806 ( .A(n1087), .B(n1084), .Z(n1086) );
  XNOR U807 ( .A(n19), .B(n1080), .Z(n1082) );
  IV U808 ( .A(n16), .Z(n19) );
  XNOR U809 ( .A(n1088), .B(n1089), .Z(n16) );
  AND U810 ( .A(n1060), .B(n1090), .Z(n1089) );
  XOR U811 ( .A(n1091), .B(n1088), .Z(n1090) );
  XOR U812 ( .A(n1092), .B(n1093), .Z(n1080) );
  AND U813 ( .A(n1094), .B(n1095), .Z(n1093) );
  XOR U814 ( .A(n1092), .B(n23), .Z(n1095) );
  XOR U815 ( .A(n1096), .B(n1097), .Z(n23) );
  AND U816 ( .A(n1063), .B(n1098), .Z(n1097) );
  XOR U817 ( .A(n1099), .B(n1096), .Z(n1098) );
  XNOR U818 ( .A(n24), .B(n1092), .Z(n1094) );
  IV U819 ( .A(n21), .Z(n24) );
  XNOR U820 ( .A(n1100), .B(n1101), .Z(n21) );
  AND U821 ( .A(n1060), .B(n1102), .Z(n1101) );
  XOR U822 ( .A(n1103), .B(n1100), .Z(n1102) );
  XOR U823 ( .A(n1104), .B(n1105), .Z(n1092) );
  AND U824 ( .A(n1106), .B(n1107), .Z(n1105) );
  XOR U825 ( .A(n1104), .B(n28), .Z(n1107) );
  XOR U826 ( .A(n1108), .B(n1109), .Z(n28) );
  AND U827 ( .A(n1063), .B(n1110), .Z(n1109) );
  XOR U828 ( .A(n1111), .B(n1108), .Z(n1110) );
  XNOR U829 ( .A(n29), .B(n1104), .Z(n1106) );
  IV U830 ( .A(n26), .Z(n29) );
  XNOR U831 ( .A(n1112), .B(n1113), .Z(n26) );
  AND U832 ( .A(n1060), .B(n1114), .Z(n1113) );
  XOR U833 ( .A(n1115), .B(n1112), .Z(n1114) );
  XOR U834 ( .A(n1116), .B(n1117), .Z(n1104) );
  AND U835 ( .A(n1118), .B(n1119), .Z(n1117) );
  XOR U836 ( .A(n1116), .B(n33), .Z(n1119) );
  XOR U837 ( .A(n1120), .B(n1121), .Z(n33) );
  AND U838 ( .A(n1063), .B(n1122), .Z(n1121) );
  XOR U839 ( .A(n1123), .B(n1120), .Z(n1122) );
  XNOR U840 ( .A(n34), .B(n1116), .Z(n1118) );
  IV U841 ( .A(n31), .Z(n34) );
  XNOR U842 ( .A(n1124), .B(n1125), .Z(n31) );
  AND U843 ( .A(n1060), .B(n1126), .Z(n1125) );
  XOR U844 ( .A(n1127), .B(n1124), .Z(n1126) );
  XOR U845 ( .A(n1128), .B(n1129), .Z(n1116) );
  AND U846 ( .A(n1130), .B(n1131), .Z(n1129) );
  XOR U847 ( .A(n1128), .B(n38), .Z(n1131) );
  XOR U848 ( .A(n1132), .B(n1133), .Z(n38) );
  AND U849 ( .A(n1063), .B(n1134), .Z(n1133) );
  XOR U850 ( .A(n1135), .B(n1132), .Z(n1134) );
  XNOR U851 ( .A(n39), .B(n1128), .Z(n1130) );
  IV U852 ( .A(n36), .Z(n39) );
  XNOR U853 ( .A(n1136), .B(n1137), .Z(n36) );
  AND U854 ( .A(n1060), .B(n1138), .Z(n1137) );
  XOR U855 ( .A(n1139), .B(n1136), .Z(n1138) );
  XOR U856 ( .A(n1140), .B(n1141), .Z(n1128) );
  AND U857 ( .A(n1142), .B(n1143), .Z(n1141) );
  XOR U858 ( .A(n1140), .B(n43), .Z(n1143) );
  XOR U859 ( .A(n1144), .B(n1145), .Z(n43) );
  AND U860 ( .A(n1063), .B(n1146), .Z(n1145) );
  XOR U861 ( .A(n1147), .B(n1144), .Z(n1146) );
  XNOR U862 ( .A(n44), .B(n1140), .Z(n1142) );
  IV U863 ( .A(n41), .Z(n44) );
  XNOR U864 ( .A(n1148), .B(n1149), .Z(n41) );
  AND U865 ( .A(n1060), .B(n1150), .Z(n1149) );
  XOR U866 ( .A(n1151), .B(n1148), .Z(n1150) );
  XOR U867 ( .A(n1152), .B(n1153), .Z(n1140) );
  AND U868 ( .A(n1154), .B(n1155), .Z(n1153) );
  XOR U869 ( .A(n1152), .B(n48), .Z(n1155) );
  XOR U870 ( .A(n1156), .B(n1157), .Z(n48) );
  AND U871 ( .A(n1063), .B(n1158), .Z(n1157) );
  XOR U872 ( .A(n1159), .B(n1156), .Z(n1158) );
  XNOR U873 ( .A(n49), .B(n1152), .Z(n1154) );
  IV U874 ( .A(n46), .Z(n49) );
  XNOR U875 ( .A(n1160), .B(n1161), .Z(n46) );
  AND U876 ( .A(n1060), .B(n1162), .Z(n1161) );
  XOR U877 ( .A(n1163), .B(n1160), .Z(n1162) );
  XOR U878 ( .A(n1164), .B(n1165), .Z(n1152) );
  AND U879 ( .A(n1166), .B(n1167), .Z(n1165) );
  XOR U880 ( .A(n1164), .B(n53), .Z(n1167) );
  XOR U881 ( .A(n1168), .B(n1169), .Z(n53) );
  AND U882 ( .A(n1063), .B(n1170), .Z(n1169) );
  XOR U883 ( .A(n1171), .B(n1168), .Z(n1170) );
  XNOR U884 ( .A(n54), .B(n1164), .Z(n1166) );
  IV U885 ( .A(n51), .Z(n54) );
  XNOR U886 ( .A(n1172), .B(n1173), .Z(n51) );
  AND U887 ( .A(n1060), .B(n1174), .Z(n1173) );
  XOR U888 ( .A(n1175), .B(n1172), .Z(n1174) );
  XOR U889 ( .A(n1176), .B(n1177), .Z(n1164) );
  AND U890 ( .A(n1178), .B(n1179), .Z(n1177) );
  XOR U891 ( .A(n1176), .B(n58), .Z(n1179) );
  XOR U892 ( .A(n1180), .B(n1181), .Z(n58) );
  AND U893 ( .A(n1063), .B(n1182), .Z(n1181) );
  XOR U894 ( .A(n1183), .B(n1180), .Z(n1182) );
  XNOR U895 ( .A(n59), .B(n1176), .Z(n1178) );
  IV U896 ( .A(n56), .Z(n59) );
  XNOR U897 ( .A(n1184), .B(n1185), .Z(n56) );
  AND U898 ( .A(n1060), .B(n1186), .Z(n1185) );
  XOR U899 ( .A(n1187), .B(n1184), .Z(n1186) );
  XOR U900 ( .A(n1188), .B(n1189), .Z(n1176) );
  AND U901 ( .A(n1190), .B(n1191), .Z(n1189) );
  XOR U902 ( .A(n1188), .B(n63), .Z(n1191) );
  XOR U903 ( .A(n1192), .B(n1193), .Z(n63) );
  AND U904 ( .A(n1063), .B(n1194), .Z(n1193) );
  XOR U905 ( .A(n1195), .B(n1192), .Z(n1194) );
  XNOR U906 ( .A(n64), .B(n1188), .Z(n1190) );
  IV U907 ( .A(n61), .Z(n64) );
  XNOR U908 ( .A(n1196), .B(n1197), .Z(n61) );
  AND U909 ( .A(n1060), .B(n1198), .Z(n1197) );
  XOR U910 ( .A(n1199), .B(n1196), .Z(n1198) );
  XOR U911 ( .A(n1200), .B(n1201), .Z(n1188) );
  AND U912 ( .A(n1202), .B(n1203), .Z(n1201) );
  XOR U913 ( .A(n1200), .B(n68), .Z(n1203) );
  XOR U914 ( .A(n1204), .B(n1205), .Z(n68) );
  AND U915 ( .A(n1063), .B(n1206), .Z(n1205) );
  XOR U916 ( .A(n1207), .B(n1204), .Z(n1206) );
  XNOR U917 ( .A(n69), .B(n1200), .Z(n1202) );
  IV U918 ( .A(n66), .Z(n69) );
  XNOR U919 ( .A(n1208), .B(n1209), .Z(n66) );
  AND U920 ( .A(n1060), .B(n1210), .Z(n1209) );
  XOR U921 ( .A(n1211), .B(n1208), .Z(n1210) );
  XOR U922 ( .A(n1212), .B(n1213), .Z(n1200) );
  AND U923 ( .A(n1214), .B(n1215), .Z(n1213) );
  XOR U924 ( .A(n1212), .B(n73), .Z(n1215) );
  XOR U925 ( .A(n1216), .B(n1217), .Z(n73) );
  AND U926 ( .A(n1063), .B(n1218), .Z(n1217) );
  XOR U927 ( .A(n1219), .B(n1216), .Z(n1218) );
  XNOR U928 ( .A(n74), .B(n1212), .Z(n1214) );
  IV U929 ( .A(n71), .Z(n74) );
  XNOR U930 ( .A(n1220), .B(n1221), .Z(n71) );
  AND U931 ( .A(n1060), .B(n1222), .Z(n1221) );
  XOR U932 ( .A(n1223), .B(n1220), .Z(n1222) );
  XOR U933 ( .A(n1224), .B(n1225), .Z(n1212) );
  AND U934 ( .A(n1226), .B(n1227), .Z(n1225) );
  XOR U935 ( .A(n1224), .B(n78), .Z(n1227) );
  XOR U936 ( .A(n1228), .B(n1229), .Z(n78) );
  AND U937 ( .A(n1063), .B(n1230), .Z(n1229) );
  XOR U938 ( .A(n1231), .B(n1228), .Z(n1230) );
  XNOR U939 ( .A(n79), .B(n1224), .Z(n1226) );
  IV U940 ( .A(n76), .Z(n79) );
  XNOR U941 ( .A(n1232), .B(n1233), .Z(n76) );
  AND U942 ( .A(n1060), .B(n1234), .Z(n1233) );
  XOR U943 ( .A(n1235), .B(n1232), .Z(n1234) );
  XNOR U944 ( .A(n1236), .B(n1237), .Z(n1224) );
  AND U945 ( .A(n1238), .B(n1239), .Z(n1237) );
  XNOR U946 ( .A(n1236), .B(n5), .Z(n1239) );
  XOR U947 ( .A(n1240), .B(n1241), .Z(n5) );
  AND U948 ( .A(n1063), .B(n1242), .Z(n1241) );
  XOR U949 ( .A(n1240), .B(n1243), .Z(n1242) );
  XOR U950 ( .A(n4), .B(n1236), .Z(n1238) );
  IV U951 ( .A(n2), .Z(n4) );
  XNOR U952 ( .A(n1244), .B(n1245), .Z(n2) );
  AND U953 ( .A(n1060), .B(n1246), .Z(n1245) );
  XOR U954 ( .A(n1244), .B(n1247), .Z(n1246) );
  AND U955 ( .A(n7), .B(n9), .Z(n1236) );
  XNOR U956 ( .A(n1248), .B(n1249), .Z(n9) );
  AND U957 ( .A(n1063), .B(n1250), .Z(n1249) );
  XNOR U958 ( .A(n1251), .B(n1248), .Z(n1250) );
  XOR U959 ( .A(n1252), .B(n1253), .Z(n1063) );
  AND U960 ( .A(n1254), .B(n1255), .Z(n1253) );
  XOR U961 ( .A(n1252), .B(n1075), .Z(n1255) );
  XOR U962 ( .A(n1256), .B(n1257), .Z(n1075) );
  AND U963 ( .A(n1047), .B(n1258), .Z(n1257) );
  XOR U964 ( .A(n1259), .B(n1256), .Z(n1258) );
  XNOR U965 ( .A(n1072), .B(n1252), .Z(n1254) );
  XOR U966 ( .A(n1260), .B(n1261), .Z(n1072) );
  AND U967 ( .A(n1045), .B(n1262), .Z(n1261) );
  XOR U968 ( .A(n1263), .B(n1260), .Z(n1262) );
  XOR U969 ( .A(n1264), .B(n1265), .Z(n1252) );
  AND U970 ( .A(n1266), .B(n1267), .Z(n1265) );
  XOR U971 ( .A(n1264), .B(n1087), .Z(n1267) );
  XOR U972 ( .A(n1268), .B(n1269), .Z(n1087) );
  AND U973 ( .A(n1047), .B(n1270), .Z(n1269) );
  XOR U974 ( .A(n1271), .B(n1268), .Z(n1270) );
  XNOR U975 ( .A(n1084), .B(n1264), .Z(n1266) );
  XOR U976 ( .A(n1272), .B(n1273), .Z(n1084) );
  AND U977 ( .A(n1045), .B(n1274), .Z(n1273) );
  XOR U978 ( .A(n1275), .B(n1272), .Z(n1274) );
  XOR U979 ( .A(n1276), .B(n1277), .Z(n1264) );
  AND U980 ( .A(n1278), .B(n1279), .Z(n1277) );
  XOR U981 ( .A(n1276), .B(n1099), .Z(n1279) );
  XOR U982 ( .A(n1280), .B(n1281), .Z(n1099) );
  AND U983 ( .A(n1047), .B(n1282), .Z(n1281) );
  XOR U984 ( .A(n1283), .B(n1280), .Z(n1282) );
  XNOR U985 ( .A(n1096), .B(n1276), .Z(n1278) );
  XOR U986 ( .A(n1284), .B(n1285), .Z(n1096) );
  AND U987 ( .A(n1045), .B(n1286), .Z(n1285) );
  XOR U988 ( .A(n1287), .B(n1284), .Z(n1286) );
  XOR U989 ( .A(n1288), .B(n1289), .Z(n1276) );
  AND U990 ( .A(n1290), .B(n1291), .Z(n1289) );
  XOR U991 ( .A(n1288), .B(n1111), .Z(n1291) );
  XOR U992 ( .A(n1292), .B(n1293), .Z(n1111) );
  AND U993 ( .A(n1047), .B(n1294), .Z(n1293) );
  XOR U994 ( .A(n1295), .B(n1292), .Z(n1294) );
  XNOR U995 ( .A(n1108), .B(n1288), .Z(n1290) );
  XOR U996 ( .A(n1296), .B(n1297), .Z(n1108) );
  AND U997 ( .A(n1045), .B(n1298), .Z(n1297) );
  XOR U998 ( .A(n1299), .B(n1296), .Z(n1298) );
  XOR U999 ( .A(n1300), .B(n1301), .Z(n1288) );
  AND U1000 ( .A(n1302), .B(n1303), .Z(n1301) );
  XOR U1001 ( .A(n1300), .B(n1123), .Z(n1303) );
  XOR U1002 ( .A(n1304), .B(n1305), .Z(n1123) );
  AND U1003 ( .A(n1047), .B(n1306), .Z(n1305) );
  XOR U1004 ( .A(n1307), .B(n1304), .Z(n1306) );
  XNOR U1005 ( .A(n1120), .B(n1300), .Z(n1302) );
  XOR U1006 ( .A(n1308), .B(n1309), .Z(n1120) );
  AND U1007 ( .A(n1045), .B(n1310), .Z(n1309) );
  XOR U1008 ( .A(n1311), .B(n1308), .Z(n1310) );
  XOR U1009 ( .A(n1312), .B(n1313), .Z(n1300) );
  AND U1010 ( .A(n1314), .B(n1315), .Z(n1313) );
  XOR U1011 ( .A(n1312), .B(n1135), .Z(n1315) );
  XOR U1012 ( .A(n1316), .B(n1317), .Z(n1135) );
  AND U1013 ( .A(n1047), .B(n1318), .Z(n1317) );
  XOR U1014 ( .A(n1319), .B(n1316), .Z(n1318) );
  XNOR U1015 ( .A(n1132), .B(n1312), .Z(n1314) );
  XOR U1016 ( .A(n1320), .B(n1321), .Z(n1132) );
  AND U1017 ( .A(n1045), .B(n1322), .Z(n1321) );
  XOR U1018 ( .A(n1323), .B(n1320), .Z(n1322) );
  XOR U1019 ( .A(n1324), .B(n1325), .Z(n1312) );
  AND U1020 ( .A(n1326), .B(n1327), .Z(n1325) );
  XOR U1021 ( .A(n1324), .B(n1147), .Z(n1327) );
  XOR U1022 ( .A(n1328), .B(n1329), .Z(n1147) );
  AND U1023 ( .A(n1047), .B(n1330), .Z(n1329) );
  XOR U1024 ( .A(n1331), .B(n1328), .Z(n1330) );
  XNOR U1025 ( .A(n1144), .B(n1324), .Z(n1326) );
  XOR U1026 ( .A(n1332), .B(n1333), .Z(n1144) );
  AND U1027 ( .A(n1045), .B(n1334), .Z(n1333) );
  XOR U1028 ( .A(n1335), .B(n1332), .Z(n1334) );
  XOR U1029 ( .A(n1336), .B(n1337), .Z(n1324) );
  AND U1030 ( .A(n1338), .B(n1339), .Z(n1337) );
  XOR U1031 ( .A(n1336), .B(n1159), .Z(n1339) );
  XOR U1032 ( .A(n1340), .B(n1341), .Z(n1159) );
  AND U1033 ( .A(n1047), .B(n1342), .Z(n1341) );
  XOR U1034 ( .A(n1343), .B(n1340), .Z(n1342) );
  XNOR U1035 ( .A(n1156), .B(n1336), .Z(n1338) );
  XOR U1036 ( .A(n1344), .B(n1345), .Z(n1156) );
  AND U1037 ( .A(n1045), .B(n1346), .Z(n1345) );
  XOR U1038 ( .A(n1347), .B(n1344), .Z(n1346) );
  XOR U1039 ( .A(n1348), .B(n1349), .Z(n1336) );
  AND U1040 ( .A(n1350), .B(n1351), .Z(n1349) );
  XOR U1041 ( .A(n1348), .B(n1171), .Z(n1351) );
  XOR U1042 ( .A(n1352), .B(n1353), .Z(n1171) );
  AND U1043 ( .A(n1047), .B(n1354), .Z(n1353) );
  XOR U1044 ( .A(n1355), .B(n1352), .Z(n1354) );
  XNOR U1045 ( .A(n1168), .B(n1348), .Z(n1350) );
  XOR U1046 ( .A(n1356), .B(n1357), .Z(n1168) );
  AND U1047 ( .A(n1045), .B(n1358), .Z(n1357) );
  XOR U1048 ( .A(n1359), .B(n1356), .Z(n1358) );
  XOR U1049 ( .A(n1360), .B(n1361), .Z(n1348) );
  AND U1050 ( .A(n1362), .B(n1363), .Z(n1361) );
  XOR U1051 ( .A(n1360), .B(n1183), .Z(n1363) );
  XOR U1052 ( .A(n1364), .B(n1365), .Z(n1183) );
  AND U1053 ( .A(n1047), .B(n1366), .Z(n1365) );
  XOR U1054 ( .A(n1367), .B(n1364), .Z(n1366) );
  XNOR U1055 ( .A(n1180), .B(n1360), .Z(n1362) );
  XOR U1056 ( .A(n1368), .B(n1369), .Z(n1180) );
  AND U1057 ( .A(n1045), .B(n1370), .Z(n1369) );
  XOR U1058 ( .A(n1371), .B(n1368), .Z(n1370) );
  XOR U1059 ( .A(n1372), .B(n1373), .Z(n1360) );
  AND U1060 ( .A(n1374), .B(n1375), .Z(n1373) );
  XOR U1061 ( .A(n1372), .B(n1195), .Z(n1375) );
  XOR U1062 ( .A(n1376), .B(n1377), .Z(n1195) );
  AND U1063 ( .A(n1047), .B(n1378), .Z(n1377) );
  XOR U1064 ( .A(n1379), .B(n1376), .Z(n1378) );
  XNOR U1065 ( .A(n1192), .B(n1372), .Z(n1374) );
  XOR U1066 ( .A(n1380), .B(n1381), .Z(n1192) );
  AND U1067 ( .A(n1045), .B(n1382), .Z(n1381) );
  XOR U1068 ( .A(n1383), .B(n1380), .Z(n1382) );
  XOR U1069 ( .A(n1384), .B(n1385), .Z(n1372) );
  AND U1070 ( .A(n1386), .B(n1387), .Z(n1385) );
  XOR U1071 ( .A(n1384), .B(n1207), .Z(n1387) );
  XOR U1072 ( .A(n1388), .B(n1389), .Z(n1207) );
  AND U1073 ( .A(n1047), .B(n1390), .Z(n1389) );
  XOR U1074 ( .A(n1391), .B(n1388), .Z(n1390) );
  XNOR U1075 ( .A(n1204), .B(n1384), .Z(n1386) );
  XOR U1076 ( .A(n1392), .B(n1393), .Z(n1204) );
  AND U1077 ( .A(n1045), .B(n1394), .Z(n1393) );
  XOR U1078 ( .A(n1395), .B(n1392), .Z(n1394) );
  XOR U1079 ( .A(n1396), .B(n1397), .Z(n1384) );
  AND U1080 ( .A(n1398), .B(n1399), .Z(n1397) );
  XOR U1081 ( .A(n1396), .B(n1219), .Z(n1399) );
  XOR U1082 ( .A(n1400), .B(n1401), .Z(n1219) );
  AND U1083 ( .A(n1047), .B(n1402), .Z(n1401) );
  XOR U1084 ( .A(n1403), .B(n1400), .Z(n1402) );
  XNOR U1085 ( .A(n1216), .B(n1396), .Z(n1398) );
  XOR U1086 ( .A(n1404), .B(n1405), .Z(n1216) );
  AND U1087 ( .A(n1045), .B(n1406), .Z(n1405) );
  XOR U1088 ( .A(n1407), .B(n1404), .Z(n1406) );
  XOR U1089 ( .A(n1408), .B(n1409), .Z(n1396) );
  AND U1090 ( .A(n1410), .B(n1411), .Z(n1409) );
  XOR U1091 ( .A(n1408), .B(n1231), .Z(n1411) );
  XOR U1092 ( .A(n1412), .B(n1413), .Z(n1231) );
  AND U1093 ( .A(n1047), .B(n1414), .Z(n1413) );
  XOR U1094 ( .A(n1415), .B(n1412), .Z(n1414) );
  XNOR U1095 ( .A(n1228), .B(n1408), .Z(n1410) );
  XOR U1096 ( .A(n1416), .B(n1417), .Z(n1228) );
  AND U1097 ( .A(n1045), .B(n1418), .Z(n1417) );
  XOR U1098 ( .A(n1419), .B(n1416), .Z(n1418) );
  XOR U1099 ( .A(n1420), .B(n1421), .Z(n1408) );
  AND U1100 ( .A(n1422), .B(n1423), .Z(n1421) );
  XNOR U1101 ( .A(n1424), .B(n1243), .Z(n1423) );
  XOR U1102 ( .A(n1425), .B(n1426), .Z(n1243) );
  AND U1103 ( .A(n1047), .B(n1427), .Z(n1426) );
  XOR U1104 ( .A(n1425), .B(n1428), .Z(n1427) );
  XNOR U1105 ( .A(n1240), .B(n1420), .Z(n1422) );
  XOR U1106 ( .A(n1429), .B(n1430), .Z(n1240) );
  AND U1107 ( .A(n1045), .B(n1431), .Z(n1430) );
  XOR U1108 ( .A(n1429), .B(n1432), .Z(n1431) );
  IV U1109 ( .A(n1424), .Z(n1420) );
  AND U1110 ( .A(n1248), .B(n1251), .Z(n1424) );
  XNOR U1111 ( .A(n1433), .B(n1434), .Z(n1251) );
  AND U1112 ( .A(n1047), .B(n1435), .Z(n1434) );
  XNOR U1113 ( .A(n1436), .B(n1433), .Z(n1435) );
  XOR U1114 ( .A(n1437), .B(n1438), .Z(n1047) );
  AND U1115 ( .A(n1439), .B(n1440), .Z(n1438) );
  XOR U1116 ( .A(n1437), .B(n1259), .Z(n1440) );
  XOR U1117 ( .A(n1441), .B(n1442), .Z(n1259) );
  AND U1118 ( .A(n1007), .B(n1443), .Z(n1442) );
  XOR U1119 ( .A(n1444), .B(n1441), .Z(n1443) );
  XNOR U1120 ( .A(n1256), .B(n1437), .Z(n1439) );
  XOR U1121 ( .A(n1445), .B(n1446), .Z(n1256) );
  AND U1122 ( .A(n1005), .B(n1447), .Z(n1446) );
  XOR U1123 ( .A(n1448), .B(n1445), .Z(n1447) );
  XOR U1124 ( .A(n1449), .B(n1450), .Z(n1437) );
  AND U1125 ( .A(n1451), .B(n1452), .Z(n1450) );
  XOR U1126 ( .A(n1449), .B(n1271), .Z(n1452) );
  XOR U1127 ( .A(n1453), .B(n1454), .Z(n1271) );
  AND U1128 ( .A(n1007), .B(n1455), .Z(n1454) );
  XOR U1129 ( .A(n1456), .B(n1453), .Z(n1455) );
  XNOR U1130 ( .A(n1268), .B(n1449), .Z(n1451) );
  XOR U1131 ( .A(n1457), .B(n1458), .Z(n1268) );
  AND U1132 ( .A(n1005), .B(n1459), .Z(n1458) );
  XOR U1133 ( .A(n1460), .B(n1457), .Z(n1459) );
  XOR U1134 ( .A(n1461), .B(n1462), .Z(n1449) );
  AND U1135 ( .A(n1463), .B(n1464), .Z(n1462) );
  XOR U1136 ( .A(n1461), .B(n1283), .Z(n1464) );
  XOR U1137 ( .A(n1465), .B(n1466), .Z(n1283) );
  AND U1138 ( .A(n1007), .B(n1467), .Z(n1466) );
  XOR U1139 ( .A(n1468), .B(n1465), .Z(n1467) );
  XNOR U1140 ( .A(n1280), .B(n1461), .Z(n1463) );
  XOR U1141 ( .A(n1469), .B(n1470), .Z(n1280) );
  AND U1142 ( .A(n1005), .B(n1471), .Z(n1470) );
  XOR U1143 ( .A(n1472), .B(n1469), .Z(n1471) );
  XOR U1144 ( .A(n1473), .B(n1474), .Z(n1461) );
  AND U1145 ( .A(n1475), .B(n1476), .Z(n1474) );
  XOR U1146 ( .A(n1473), .B(n1295), .Z(n1476) );
  XOR U1147 ( .A(n1477), .B(n1478), .Z(n1295) );
  AND U1148 ( .A(n1007), .B(n1479), .Z(n1478) );
  XOR U1149 ( .A(n1480), .B(n1477), .Z(n1479) );
  XNOR U1150 ( .A(n1292), .B(n1473), .Z(n1475) );
  XOR U1151 ( .A(n1481), .B(n1482), .Z(n1292) );
  AND U1152 ( .A(n1005), .B(n1483), .Z(n1482) );
  XOR U1153 ( .A(n1484), .B(n1481), .Z(n1483) );
  XOR U1154 ( .A(n1485), .B(n1486), .Z(n1473) );
  AND U1155 ( .A(n1487), .B(n1488), .Z(n1486) );
  XOR U1156 ( .A(n1485), .B(n1307), .Z(n1488) );
  XOR U1157 ( .A(n1489), .B(n1490), .Z(n1307) );
  AND U1158 ( .A(n1007), .B(n1491), .Z(n1490) );
  XOR U1159 ( .A(n1492), .B(n1489), .Z(n1491) );
  XNOR U1160 ( .A(n1304), .B(n1485), .Z(n1487) );
  XOR U1161 ( .A(n1493), .B(n1494), .Z(n1304) );
  AND U1162 ( .A(n1005), .B(n1495), .Z(n1494) );
  XOR U1163 ( .A(n1496), .B(n1493), .Z(n1495) );
  XOR U1164 ( .A(n1497), .B(n1498), .Z(n1485) );
  AND U1165 ( .A(n1499), .B(n1500), .Z(n1498) );
  XOR U1166 ( .A(n1497), .B(n1319), .Z(n1500) );
  XOR U1167 ( .A(n1501), .B(n1502), .Z(n1319) );
  AND U1168 ( .A(n1007), .B(n1503), .Z(n1502) );
  XOR U1169 ( .A(n1504), .B(n1501), .Z(n1503) );
  XNOR U1170 ( .A(n1316), .B(n1497), .Z(n1499) );
  XOR U1171 ( .A(n1505), .B(n1506), .Z(n1316) );
  AND U1172 ( .A(n1005), .B(n1507), .Z(n1506) );
  XOR U1173 ( .A(n1508), .B(n1505), .Z(n1507) );
  XOR U1174 ( .A(n1509), .B(n1510), .Z(n1497) );
  AND U1175 ( .A(n1511), .B(n1512), .Z(n1510) );
  XOR U1176 ( .A(n1509), .B(n1331), .Z(n1512) );
  XOR U1177 ( .A(n1513), .B(n1514), .Z(n1331) );
  AND U1178 ( .A(n1007), .B(n1515), .Z(n1514) );
  XOR U1179 ( .A(n1516), .B(n1513), .Z(n1515) );
  XNOR U1180 ( .A(n1328), .B(n1509), .Z(n1511) );
  XOR U1181 ( .A(n1517), .B(n1518), .Z(n1328) );
  AND U1182 ( .A(n1005), .B(n1519), .Z(n1518) );
  XOR U1183 ( .A(n1520), .B(n1517), .Z(n1519) );
  XOR U1184 ( .A(n1521), .B(n1522), .Z(n1509) );
  AND U1185 ( .A(n1523), .B(n1524), .Z(n1522) );
  XOR U1186 ( .A(n1521), .B(n1343), .Z(n1524) );
  XOR U1187 ( .A(n1525), .B(n1526), .Z(n1343) );
  AND U1188 ( .A(n1007), .B(n1527), .Z(n1526) );
  XOR U1189 ( .A(n1528), .B(n1525), .Z(n1527) );
  XNOR U1190 ( .A(n1340), .B(n1521), .Z(n1523) );
  XOR U1191 ( .A(n1529), .B(n1530), .Z(n1340) );
  AND U1192 ( .A(n1005), .B(n1531), .Z(n1530) );
  XOR U1193 ( .A(n1532), .B(n1529), .Z(n1531) );
  XOR U1194 ( .A(n1533), .B(n1534), .Z(n1521) );
  AND U1195 ( .A(n1535), .B(n1536), .Z(n1534) );
  XOR U1196 ( .A(n1533), .B(n1355), .Z(n1536) );
  XOR U1197 ( .A(n1537), .B(n1538), .Z(n1355) );
  AND U1198 ( .A(n1007), .B(n1539), .Z(n1538) );
  XOR U1199 ( .A(n1540), .B(n1537), .Z(n1539) );
  XNOR U1200 ( .A(n1352), .B(n1533), .Z(n1535) );
  XOR U1201 ( .A(n1541), .B(n1542), .Z(n1352) );
  AND U1202 ( .A(n1005), .B(n1543), .Z(n1542) );
  XOR U1203 ( .A(n1544), .B(n1541), .Z(n1543) );
  XOR U1204 ( .A(n1545), .B(n1546), .Z(n1533) );
  AND U1205 ( .A(n1547), .B(n1548), .Z(n1546) );
  XOR U1206 ( .A(n1545), .B(n1367), .Z(n1548) );
  XOR U1207 ( .A(n1549), .B(n1550), .Z(n1367) );
  AND U1208 ( .A(n1007), .B(n1551), .Z(n1550) );
  XOR U1209 ( .A(n1552), .B(n1549), .Z(n1551) );
  XNOR U1210 ( .A(n1364), .B(n1545), .Z(n1547) );
  XOR U1211 ( .A(n1553), .B(n1554), .Z(n1364) );
  AND U1212 ( .A(n1005), .B(n1555), .Z(n1554) );
  XOR U1213 ( .A(n1556), .B(n1553), .Z(n1555) );
  XOR U1214 ( .A(n1557), .B(n1558), .Z(n1545) );
  AND U1215 ( .A(n1559), .B(n1560), .Z(n1558) );
  XOR U1216 ( .A(n1557), .B(n1379), .Z(n1560) );
  XOR U1217 ( .A(n1561), .B(n1562), .Z(n1379) );
  AND U1218 ( .A(n1007), .B(n1563), .Z(n1562) );
  XOR U1219 ( .A(n1564), .B(n1561), .Z(n1563) );
  XNOR U1220 ( .A(n1376), .B(n1557), .Z(n1559) );
  XOR U1221 ( .A(n1565), .B(n1566), .Z(n1376) );
  AND U1222 ( .A(n1005), .B(n1567), .Z(n1566) );
  XOR U1223 ( .A(n1568), .B(n1565), .Z(n1567) );
  XOR U1224 ( .A(n1569), .B(n1570), .Z(n1557) );
  AND U1225 ( .A(n1571), .B(n1572), .Z(n1570) );
  XOR U1226 ( .A(n1569), .B(n1391), .Z(n1572) );
  XOR U1227 ( .A(n1573), .B(n1574), .Z(n1391) );
  AND U1228 ( .A(n1007), .B(n1575), .Z(n1574) );
  XOR U1229 ( .A(n1576), .B(n1573), .Z(n1575) );
  XNOR U1230 ( .A(n1388), .B(n1569), .Z(n1571) );
  XOR U1231 ( .A(n1577), .B(n1578), .Z(n1388) );
  AND U1232 ( .A(n1005), .B(n1579), .Z(n1578) );
  XOR U1233 ( .A(n1580), .B(n1577), .Z(n1579) );
  XOR U1234 ( .A(n1581), .B(n1582), .Z(n1569) );
  AND U1235 ( .A(n1583), .B(n1584), .Z(n1582) );
  XOR U1236 ( .A(n1581), .B(n1403), .Z(n1584) );
  XOR U1237 ( .A(n1585), .B(n1586), .Z(n1403) );
  AND U1238 ( .A(n1007), .B(n1587), .Z(n1586) );
  XOR U1239 ( .A(n1588), .B(n1585), .Z(n1587) );
  XNOR U1240 ( .A(n1400), .B(n1581), .Z(n1583) );
  XOR U1241 ( .A(n1589), .B(n1590), .Z(n1400) );
  AND U1242 ( .A(n1005), .B(n1591), .Z(n1590) );
  XOR U1243 ( .A(n1592), .B(n1589), .Z(n1591) );
  XOR U1244 ( .A(n1593), .B(n1594), .Z(n1581) );
  AND U1245 ( .A(n1595), .B(n1596), .Z(n1594) );
  XOR U1246 ( .A(n1593), .B(n1415), .Z(n1596) );
  XOR U1247 ( .A(n1597), .B(n1598), .Z(n1415) );
  AND U1248 ( .A(n1007), .B(n1599), .Z(n1598) );
  XOR U1249 ( .A(n1600), .B(n1597), .Z(n1599) );
  XNOR U1250 ( .A(n1412), .B(n1593), .Z(n1595) );
  XOR U1251 ( .A(n1601), .B(n1602), .Z(n1412) );
  AND U1252 ( .A(n1005), .B(n1603), .Z(n1602) );
  XOR U1253 ( .A(n1604), .B(n1601), .Z(n1603) );
  XOR U1254 ( .A(n1605), .B(n1606), .Z(n1593) );
  AND U1255 ( .A(n1607), .B(n1608), .Z(n1606) );
  XNOR U1256 ( .A(n1609), .B(n1428), .Z(n1608) );
  XOR U1257 ( .A(n1610), .B(n1611), .Z(n1428) );
  AND U1258 ( .A(n1007), .B(n1612), .Z(n1611) );
  XOR U1259 ( .A(n1610), .B(n1613), .Z(n1612) );
  XNOR U1260 ( .A(n1425), .B(n1605), .Z(n1607) );
  XOR U1261 ( .A(n1614), .B(n1615), .Z(n1425) );
  AND U1262 ( .A(n1005), .B(n1616), .Z(n1615) );
  XOR U1263 ( .A(n1614), .B(n1617), .Z(n1616) );
  IV U1264 ( .A(n1609), .Z(n1605) );
  AND U1265 ( .A(n1433), .B(n1436), .Z(n1609) );
  XNOR U1266 ( .A(n1618), .B(n1619), .Z(n1436) );
  AND U1267 ( .A(n1007), .B(n1620), .Z(n1619) );
  XNOR U1268 ( .A(n1621), .B(n1618), .Z(n1620) );
  XOR U1269 ( .A(n1622), .B(n1623), .Z(n1007) );
  AND U1270 ( .A(n1624), .B(n1625), .Z(n1623) );
  XOR U1271 ( .A(n1622), .B(n1444), .Z(n1625) );
  XNOR U1272 ( .A(n1626), .B(n1627), .Z(n1444) );
  AND U1273 ( .A(n1628), .B(n919), .Z(n1627) );
  AND U1274 ( .A(n1626), .B(n1629), .Z(n1628) );
  XNOR U1275 ( .A(n1441), .B(n1622), .Z(n1624) );
  XOR U1276 ( .A(n1630), .B(n1631), .Z(n1441) );
  AND U1277 ( .A(n1632), .B(n917), .Z(n1631) );
  NOR U1278 ( .A(n1630), .B(n1633), .Z(n1632) );
  XOR U1279 ( .A(n1634), .B(n1635), .Z(n1622) );
  AND U1280 ( .A(n1636), .B(n1637), .Z(n1635) );
  XOR U1281 ( .A(n1634), .B(n1456), .Z(n1637) );
  XOR U1282 ( .A(n1638), .B(n1639), .Z(n1456) );
  AND U1283 ( .A(n919), .B(n1640), .Z(n1639) );
  XOR U1284 ( .A(n1641), .B(n1638), .Z(n1640) );
  XNOR U1285 ( .A(n1453), .B(n1634), .Z(n1636) );
  XOR U1286 ( .A(n1642), .B(n1643), .Z(n1453) );
  AND U1287 ( .A(n917), .B(n1644), .Z(n1643) );
  XOR U1288 ( .A(n1645), .B(n1642), .Z(n1644) );
  XOR U1289 ( .A(n1646), .B(n1647), .Z(n1634) );
  AND U1290 ( .A(n1648), .B(n1649), .Z(n1647) );
  XOR U1291 ( .A(n1646), .B(n1468), .Z(n1649) );
  XOR U1292 ( .A(n1650), .B(n1651), .Z(n1468) );
  AND U1293 ( .A(n919), .B(n1652), .Z(n1651) );
  XOR U1294 ( .A(n1653), .B(n1650), .Z(n1652) );
  XNOR U1295 ( .A(n1465), .B(n1646), .Z(n1648) );
  XOR U1296 ( .A(n1654), .B(n1655), .Z(n1465) );
  AND U1297 ( .A(n917), .B(n1656), .Z(n1655) );
  XOR U1298 ( .A(n1657), .B(n1654), .Z(n1656) );
  XOR U1299 ( .A(n1658), .B(n1659), .Z(n1646) );
  AND U1300 ( .A(n1660), .B(n1661), .Z(n1659) );
  XOR U1301 ( .A(n1658), .B(n1480), .Z(n1661) );
  XOR U1302 ( .A(n1662), .B(n1663), .Z(n1480) );
  AND U1303 ( .A(n919), .B(n1664), .Z(n1663) );
  XOR U1304 ( .A(n1665), .B(n1662), .Z(n1664) );
  XNOR U1305 ( .A(n1477), .B(n1658), .Z(n1660) );
  XOR U1306 ( .A(n1666), .B(n1667), .Z(n1477) );
  AND U1307 ( .A(n917), .B(n1668), .Z(n1667) );
  XOR U1308 ( .A(n1669), .B(n1666), .Z(n1668) );
  XOR U1309 ( .A(n1670), .B(n1671), .Z(n1658) );
  AND U1310 ( .A(n1672), .B(n1673), .Z(n1671) );
  XOR U1311 ( .A(n1670), .B(n1492), .Z(n1673) );
  XOR U1312 ( .A(n1674), .B(n1675), .Z(n1492) );
  AND U1313 ( .A(n919), .B(n1676), .Z(n1675) );
  XOR U1314 ( .A(n1677), .B(n1674), .Z(n1676) );
  XNOR U1315 ( .A(n1489), .B(n1670), .Z(n1672) );
  XOR U1316 ( .A(n1678), .B(n1679), .Z(n1489) );
  AND U1317 ( .A(n917), .B(n1680), .Z(n1679) );
  XOR U1318 ( .A(n1681), .B(n1678), .Z(n1680) );
  XOR U1319 ( .A(n1682), .B(n1683), .Z(n1670) );
  AND U1320 ( .A(n1684), .B(n1685), .Z(n1683) );
  XOR U1321 ( .A(n1682), .B(n1504), .Z(n1685) );
  XOR U1322 ( .A(n1686), .B(n1687), .Z(n1504) );
  AND U1323 ( .A(n919), .B(n1688), .Z(n1687) );
  XOR U1324 ( .A(n1689), .B(n1686), .Z(n1688) );
  XNOR U1325 ( .A(n1501), .B(n1682), .Z(n1684) );
  XOR U1326 ( .A(n1690), .B(n1691), .Z(n1501) );
  AND U1327 ( .A(n917), .B(n1692), .Z(n1691) );
  XOR U1328 ( .A(n1693), .B(n1690), .Z(n1692) );
  XOR U1329 ( .A(n1694), .B(n1695), .Z(n1682) );
  AND U1330 ( .A(n1696), .B(n1697), .Z(n1695) );
  XOR U1331 ( .A(n1694), .B(n1516), .Z(n1697) );
  XOR U1332 ( .A(n1698), .B(n1699), .Z(n1516) );
  AND U1333 ( .A(n919), .B(n1700), .Z(n1699) );
  XOR U1334 ( .A(n1701), .B(n1698), .Z(n1700) );
  XNOR U1335 ( .A(n1513), .B(n1694), .Z(n1696) );
  XOR U1336 ( .A(n1702), .B(n1703), .Z(n1513) );
  AND U1337 ( .A(n917), .B(n1704), .Z(n1703) );
  XOR U1338 ( .A(n1705), .B(n1702), .Z(n1704) );
  XOR U1339 ( .A(n1706), .B(n1707), .Z(n1694) );
  AND U1340 ( .A(n1708), .B(n1709), .Z(n1707) );
  XOR U1341 ( .A(n1706), .B(n1528), .Z(n1709) );
  XOR U1342 ( .A(n1710), .B(n1711), .Z(n1528) );
  AND U1343 ( .A(n919), .B(n1712), .Z(n1711) );
  XOR U1344 ( .A(n1713), .B(n1710), .Z(n1712) );
  XNOR U1345 ( .A(n1525), .B(n1706), .Z(n1708) );
  XOR U1346 ( .A(n1714), .B(n1715), .Z(n1525) );
  AND U1347 ( .A(n917), .B(n1716), .Z(n1715) );
  XOR U1348 ( .A(n1717), .B(n1714), .Z(n1716) );
  XOR U1349 ( .A(n1718), .B(n1719), .Z(n1706) );
  AND U1350 ( .A(n1720), .B(n1721), .Z(n1719) );
  XOR U1351 ( .A(n1718), .B(n1540), .Z(n1721) );
  XOR U1352 ( .A(n1722), .B(n1723), .Z(n1540) );
  AND U1353 ( .A(n919), .B(n1724), .Z(n1723) );
  XOR U1354 ( .A(n1725), .B(n1722), .Z(n1724) );
  XNOR U1355 ( .A(n1537), .B(n1718), .Z(n1720) );
  XOR U1356 ( .A(n1726), .B(n1727), .Z(n1537) );
  AND U1357 ( .A(n917), .B(n1728), .Z(n1727) );
  XOR U1358 ( .A(n1729), .B(n1726), .Z(n1728) );
  XOR U1359 ( .A(n1730), .B(n1731), .Z(n1718) );
  AND U1360 ( .A(n1732), .B(n1733), .Z(n1731) );
  XOR U1361 ( .A(n1730), .B(n1552), .Z(n1733) );
  XOR U1362 ( .A(n1734), .B(n1735), .Z(n1552) );
  AND U1363 ( .A(n919), .B(n1736), .Z(n1735) );
  XOR U1364 ( .A(n1737), .B(n1734), .Z(n1736) );
  XNOR U1365 ( .A(n1549), .B(n1730), .Z(n1732) );
  XOR U1366 ( .A(n1738), .B(n1739), .Z(n1549) );
  AND U1367 ( .A(n917), .B(n1740), .Z(n1739) );
  XOR U1368 ( .A(n1741), .B(n1738), .Z(n1740) );
  XOR U1369 ( .A(n1742), .B(n1743), .Z(n1730) );
  AND U1370 ( .A(n1744), .B(n1745), .Z(n1743) );
  XOR U1371 ( .A(n1742), .B(n1564), .Z(n1745) );
  XOR U1372 ( .A(n1746), .B(n1747), .Z(n1564) );
  AND U1373 ( .A(n919), .B(n1748), .Z(n1747) );
  XOR U1374 ( .A(n1749), .B(n1746), .Z(n1748) );
  XNOR U1375 ( .A(n1561), .B(n1742), .Z(n1744) );
  XOR U1376 ( .A(n1750), .B(n1751), .Z(n1561) );
  AND U1377 ( .A(n917), .B(n1752), .Z(n1751) );
  XOR U1378 ( .A(n1753), .B(n1750), .Z(n1752) );
  XOR U1379 ( .A(n1754), .B(n1755), .Z(n1742) );
  AND U1380 ( .A(n1756), .B(n1757), .Z(n1755) );
  XOR U1381 ( .A(n1754), .B(n1576), .Z(n1757) );
  XOR U1382 ( .A(n1758), .B(n1759), .Z(n1576) );
  AND U1383 ( .A(n919), .B(n1760), .Z(n1759) );
  XOR U1384 ( .A(n1761), .B(n1758), .Z(n1760) );
  XNOR U1385 ( .A(n1573), .B(n1754), .Z(n1756) );
  XOR U1386 ( .A(n1762), .B(n1763), .Z(n1573) );
  AND U1387 ( .A(n917), .B(n1764), .Z(n1763) );
  XOR U1388 ( .A(n1765), .B(n1762), .Z(n1764) );
  XOR U1389 ( .A(n1766), .B(n1767), .Z(n1754) );
  AND U1390 ( .A(n1768), .B(n1769), .Z(n1767) );
  XOR U1391 ( .A(n1766), .B(n1588), .Z(n1769) );
  XOR U1392 ( .A(n1770), .B(n1771), .Z(n1588) );
  AND U1393 ( .A(n919), .B(n1772), .Z(n1771) );
  XOR U1394 ( .A(n1773), .B(n1770), .Z(n1772) );
  XNOR U1395 ( .A(n1585), .B(n1766), .Z(n1768) );
  XOR U1396 ( .A(n1774), .B(n1775), .Z(n1585) );
  AND U1397 ( .A(n917), .B(n1776), .Z(n1775) );
  XOR U1398 ( .A(n1777), .B(n1774), .Z(n1776) );
  XOR U1399 ( .A(n1778), .B(n1779), .Z(n1766) );
  AND U1400 ( .A(n1780), .B(n1781), .Z(n1779) );
  XOR U1401 ( .A(n1778), .B(n1600), .Z(n1781) );
  XOR U1402 ( .A(n1782), .B(n1783), .Z(n1600) );
  AND U1403 ( .A(n919), .B(n1784), .Z(n1783) );
  XOR U1404 ( .A(n1785), .B(n1782), .Z(n1784) );
  XNOR U1405 ( .A(n1597), .B(n1778), .Z(n1780) );
  XOR U1406 ( .A(n1786), .B(n1787), .Z(n1597) );
  AND U1407 ( .A(n917), .B(n1788), .Z(n1787) );
  XOR U1408 ( .A(n1789), .B(n1786), .Z(n1788) );
  XOR U1409 ( .A(n1790), .B(n1791), .Z(n1778) );
  AND U1410 ( .A(n1792), .B(n1793), .Z(n1791) );
  XNOR U1411 ( .A(n1794), .B(n1613), .Z(n1793) );
  XOR U1412 ( .A(n1795), .B(n1796), .Z(n1613) );
  AND U1413 ( .A(n919), .B(n1797), .Z(n1796) );
  XOR U1414 ( .A(n1795), .B(n1798), .Z(n1797) );
  XNOR U1415 ( .A(n1610), .B(n1790), .Z(n1792) );
  XOR U1416 ( .A(n1799), .B(n1800), .Z(n1610) );
  AND U1417 ( .A(n917), .B(n1801), .Z(n1800) );
  XOR U1418 ( .A(n1799), .B(n1802), .Z(n1801) );
  IV U1419 ( .A(n1794), .Z(n1790) );
  AND U1420 ( .A(n1618), .B(n1621), .Z(n1794) );
  XNOR U1421 ( .A(n1803), .B(n1804), .Z(n1621) );
  AND U1422 ( .A(n919), .B(n1805), .Z(n1804) );
  XNOR U1423 ( .A(n1806), .B(n1803), .Z(n1805) );
  XOR U1424 ( .A(n1807), .B(n1808), .Z(n919) );
  AND U1425 ( .A(n1809), .B(n1810), .Z(n1808) );
  XOR U1426 ( .A(n1629), .B(n1807), .Z(n1810) );
  IV U1427 ( .A(n1811), .Z(n1629) );
  AND U1428 ( .A(n1812), .B(n1813), .Z(n1811) );
  XOR U1429 ( .A(n1807), .B(n1626), .Z(n1809) );
  AND U1430 ( .A(n1814), .B(n1815), .Z(n1626) );
  XOR U1431 ( .A(n1816), .B(n1817), .Z(n1807) );
  AND U1432 ( .A(n1818), .B(n1819), .Z(n1817) );
  XOR U1433 ( .A(n1816), .B(n1641), .Z(n1819) );
  XOR U1434 ( .A(n1820), .B(n1821), .Z(n1641) );
  AND U1435 ( .A(n735), .B(n1822), .Z(n1821) );
  XOR U1436 ( .A(n1823), .B(n1820), .Z(n1822) );
  XNOR U1437 ( .A(n1638), .B(n1816), .Z(n1818) );
  XOR U1438 ( .A(n1824), .B(n1825), .Z(n1638) );
  AND U1439 ( .A(n733), .B(n1826), .Z(n1825) );
  XOR U1440 ( .A(n1827), .B(n1824), .Z(n1826) );
  XOR U1441 ( .A(n1828), .B(n1829), .Z(n1816) );
  AND U1442 ( .A(n1830), .B(n1831), .Z(n1829) );
  XOR U1443 ( .A(n1828), .B(n1653), .Z(n1831) );
  XOR U1444 ( .A(n1832), .B(n1833), .Z(n1653) );
  AND U1445 ( .A(n735), .B(n1834), .Z(n1833) );
  XOR U1446 ( .A(n1835), .B(n1832), .Z(n1834) );
  XNOR U1447 ( .A(n1650), .B(n1828), .Z(n1830) );
  XOR U1448 ( .A(n1836), .B(n1837), .Z(n1650) );
  AND U1449 ( .A(n733), .B(n1838), .Z(n1837) );
  XOR U1450 ( .A(n1839), .B(n1836), .Z(n1838) );
  XOR U1451 ( .A(n1840), .B(n1841), .Z(n1828) );
  AND U1452 ( .A(n1842), .B(n1843), .Z(n1841) );
  XOR U1453 ( .A(n1840), .B(n1665), .Z(n1843) );
  XOR U1454 ( .A(n1844), .B(n1845), .Z(n1665) );
  AND U1455 ( .A(n735), .B(n1846), .Z(n1845) );
  XOR U1456 ( .A(n1847), .B(n1844), .Z(n1846) );
  XNOR U1457 ( .A(n1662), .B(n1840), .Z(n1842) );
  XOR U1458 ( .A(n1848), .B(n1849), .Z(n1662) );
  AND U1459 ( .A(n733), .B(n1850), .Z(n1849) );
  XOR U1460 ( .A(n1851), .B(n1848), .Z(n1850) );
  XOR U1461 ( .A(n1852), .B(n1853), .Z(n1840) );
  AND U1462 ( .A(n1854), .B(n1855), .Z(n1853) );
  XOR U1463 ( .A(n1852), .B(n1677), .Z(n1855) );
  XOR U1464 ( .A(n1856), .B(n1857), .Z(n1677) );
  AND U1465 ( .A(n735), .B(n1858), .Z(n1857) );
  XOR U1466 ( .A(n1859), .B(n1856), .Z(n1858) );
  XNOR U1467 ( .A(n1674), .B(n1852), .Z(n1854) );
  XOR U1468 ( .A(n1860), .B(n1861), .Z(n1674) );
  AND U1469 ( .A(n733), .B(n1862), .Z(n1861) );
  XOR U1470 ( .A(n1863), .B(n1860), .Z(n1862) );
  XOR U1471 ( .A(n1864), .B(n1865), .Z(n1852) );
  AND U1472 ( .A(n1866), .B(n1867), .Z(n1865) );
  XOR U1473 ( .A(n1864), .B(n1689), .Z(n1867) );
  XOR U1474 ( .A(n1868), .B(n1869), .Z(n1689) );
  AND U1475 ( .A(n735), .B(n1870), .Z(n1869) );
  XOR U1476 ( .A(n1871), .B(n1868), .Z(n1870) );
  XNOR U1477 ( .A(n1686), .B(n1864), .Z(n1866) );
  XOR U1478 ( .A(n1872), .B(n1873), .Z(n1686) );
  AND U1479 ( .A(n733), .B(n1874), .Z(n1873) );
  XOR U1480 ( .A(n1875), .B(n1872), .Z(n1874) );
  XOR U1481 ( .A(n1876), .B(n1877), .Z(n1864) );
  AND U1482 ( .A(n1878), .B(n1879), .Z(n1877) );
  XOR U1483 ( .A(n1876), .B(n1701), .Z(n1879) );
  XOR U1484 ( .A(n1880), .B(n1881), .Z(n1701) );
  AND U1485 ( .A(n735), .B(n1882), .Z(n1881) );
  XOR U1486 ( .A(n1883), .B(n1880), .Z(n1882) );
  XNOR U1487 ( .A(n1698), .B(n1876), .Z(n1878) );
  XOR U1488 ( .A(n1884), .B(n1885), .Z(n1698) );
  AND U1489 ( .A(n733), .B(n1886), .Z(n1885) );
  XOR U1490 ( .A(n1887), .B(n1884), .Z(n1886) );
  XOR U1491 ( .A(n1888), .B(n1889), .Z(n1876) );
  AND U1492 ( .A(n1890), .B(n1891), .Z(n1889) );
  XOR U1493 ( .A(n1888), .B(n1713), .Z(n1891) );
  XOR U1494 ( .A(n1892), .B(n1893), .Z(n1713) );
  AND U1495 ( .A(n735), .B(n1894), .Z(n1893) );
  XOR U1496 ( .A(n1895), .B(n1892), .Z(n1894) );
  XNOR U1497 ( .A(n1710), .B(n1888), .Z(n1890) );
  XOR U1498 ( .A(n1896), .B(n1897), .Z(n1710) );
  AND U1499 ( .A(n733), .B(n1898), .Z(n1897) );
  XOR U1500 ( .A(n1899), .B(n1896), .Z(n1898) );
  XOR U1501 ( .A(n1900), .B(n1901), .Z(n1888) );
  AND U1502 ( .A(n1902), .B(n1903), .Z(n1901) );
  XOR U1503 ( .A(n1900), .B(n1725), .Z(n1903) );
  XOR U1504 ( .A(n1904), .B(n1905), .Z(n1725) );
  AND U1505 ( .A(n735), .B(n1906), .Z(n1905) );
  XOR U1506 ( .A(n1907), .B(n1904), .Z(n1906) );
  XNOR U1507 ( .A(n1722), .B(n1900), .Z(n1902) );
  XOR U1508 ( .A(n1908), .B(n1909), .Z(n1722) );
  AND U1509 ( .A(n733), .B(n1910), .Z(n1909) );
  XOR U1510 ( .A(n1911), .B(n1908), .Z(n1910) );
  XOR U1511 ( .A(n1912), .B(n1913), .Z(n1900) );
  AND U1512 ( .A(n1914), .B(n1915), .Z(n1913) );
  XOR U1513 ( .A(n1912), .B(n1737), .Z(n1915) );
  XOR U1514 ( .A(n1916), .B(n1917), .Z(n1737) );
  AND U1515 ( .A(n735), .B(n1918), .Z(n1917) );
  XOR U1516 ( .A(n1919), .B(n1916), .Z(n1918) );
  XNOR U1517 ( .A(n1734), .B(n1912), .Z(n1914) );
  XOR U1518 ( .A(n1920), .B(n1921), .Z(n1734) );
  AND U1519 ( .A(n733), .B(n1922), .Z(n1921) );
  XOR U1520 ( .A(n1923), .B(n1920), .Z(n1922) );
  XOR U1521 ( .A(n1924), .B(n1925), .Z(n1912) );
  AND U1522 ( .A(n1926), .B(n1927), .Z(n1925) );
  XOR U1523 ( .A(n1924), .B(n1749), .Z(n1927) );
  XOR U1524 ( .A(n1928), .B(n1929), .Z(n1749) );
  AND U1525 ( .A(n735), .B(n1930), .Z(n1929) );
  XOR U1526 ( .A(n1931), .B(n1928), .Z(n1930) );
  XNOR U1527 ( .A(n1746), .B(n1924), .Z(n1926) );
  XOR U1528 ( .A(n1932), .B(n1933), .Z(n1746) );
  AND U1529 ( .A(n733), .B(n1934), .Z(n1933) );
  XOR U1530 ( .A(n1935), .B(n1932), .Z(n1934) );
  XOR U1531 ( .A(n1936), .B(n1937), .Z(n1924) );
  AND U1532 ( .A(n1938), .B(n1939), .Z(n1937) );
  XOR U1533 ( .A(n1936), .B(n1761), .Z(n1939) );
  XOR U1534 ( .A(n1940), .B(n1941), .Z(n1761) );
  AND U1535 ( .A(n735), .B(n1942), .Z(n1941) );
  XOR U1536 ( .A(n1943), .B(n1940), .Z(n1942) );
  XNOR U1537 ( .A(n1758), .B(n1936), .Z(n1938) );
  XOR U1538 ( .A(n1944), .B(n1945), .Z(n1758) );
  AND U1539 ( .A(n733), .B(n1946), .Z(n1945) );
  XOR U1540 ( .A(n1947), .B(n1944), .Z(n1946) );
  XOR U1541 ( .A(n1948), .B(n1949), .Z(n1936) );
  AND U1542 ( .A(n1950), .B(n1951), .Z(n1949) );
  XOR U1543 ( .A(n1948), .B(n1773), .Z(n1951) );
  XOR U1544 ( .A(n1952), .B(n1953), .Z(n1773) );
  AND U1545 ( .A(n735), .B(n1954), .Z(n1953) );
  XOR U1546 ( .A(n1955), .B(n1952), .Z(n1954) );
  XNOR U1547 ( .A(n1770), .B(n1948), .Z(n1950) );
  XOR U1548 ( .A(n1956), .B(n1957), .Z(n1770) );
  AND U1549 ( .A(n733), .B(n1958), .Z(n1957) );
  XOR U1550 ( .A(n1959), .B(n1956), .Z(n1958) );
  XOR U1551 ( .A(n1960), .B(n1961), .Z(n1948) );
  AND U1552 ( .A(n1962), .B(n1963), .Z(n1961) );
  XOR U1553 ( .A(n1960), .B(n1785), .Z(n1963) );
  XOR U1554 ( .A(n1964), .B(n1965), .Z(n1785) );
  AND U1555 ( .A(n735), .B(n1966), .Z(n1965) );
  XOR U1556 ( .A(n1967), .B(n1964), .Z(n1966) );
  XNOR U1557 ( .A(n1782), .B(n1960), .Z(n1962) );
  XOR U1558 ( .A(n1968), .B(n1969), .Z(n1782) );
  AND U1559 ( .A(n733), .B(n1970), .Z(n1969) );
  XOR U1560 ( .A(n1971), .B(n1968), .Z(n1970) );
  XOR U1561 ( .A(n1972), .B(n1973), .Z(n1960) );
  AND U1562 ( .A(n1974), .B(n1975), .Z(n1973) );
  XNOR U1563 ( .A(n1976), .B(n1798), .Z(n1975) );
  XOR U1564 ( .A(n1977), .B(n1978), .Z(n1798) );
  AND U1565 ( .A(n735), .B(n1979), .Z(n1978) );
  XOR U1566 ( .A(n1977), .B(n1980), .Z(n1979) );
  XNOR U1567 ( .A(n1795), .B(n1972), .Z(n1974) );
  XOR U1568 ( .A(n1981), .B(n1982), .Z(n1795) );
  AND U1569 ( .A(n733), .B(n1983), .Z(n1982) );
  XOR U1570 ( .A(n1981), .B(n1984), .Z(n1983) );
  IV U1571 ( .A(n1976), .Z(n1972) );
  AND U1572 ( .A(n1803), .B(n1806), .Z(n1976) );
  XNOR U1573 ( .A(n1985), .B(n1986), .Z(n1806) );
  AND U1574 ( .A(n735), .B(n1987), .Z(n1986) );
  XNOR U1575 ( .A(n1988), .B(n1985), .Z(n1987) );
  XOR U1576 ( .A(n1989), .B(n1990), .Z(n735) );
  AND U1577 ( .A(n1991), .B(n1992), .Z(n1990) );
  XNOR U1578 ( .A(n1812), .B(n1989), .Z(n1992) );
  AND U1579 ( .A(n1993), .B(n1994), .Z(n1812) );
  XOR U1580 ( .A(n1989), .B(n1813), .Z(n1991) );
  AND U1581 ( .A(n1995), .B(n1996), .Z(n1813) );
  XOR U1582 ( .A(n1997), .B(n1998), .Z(n1989) );
  AND U1583 ( .A(n1999), .B(n2000), .Z(n1998) );
  XOR U1584 ( .A(n1997), .B(n1823), .Z(n2000) );
  XOR U1585 ( .A(n2001), .B(n2002), .Z(n1823) );
  AND U1586 ( .A(n359), .B(n2003), .Z(n2002) );
  XOR U1587 ( .A(n2004), .B(n2001), .Z(n2003) );
  XNOR U1588 ( .A(n1820), .B(n1997), .Z(n1999) );
  XOR U1589 ( .A(n2005), .B(n2006), .Z(n1820) );
  AND U1590 ( .A(n357), .B(n2007), .Z(n2006) );
  XOR U1591 ( .A(n2008), .B(n2005), .Z(n2007) );
  XOR U1592 ( .A(n2009), .B(n2010), .Z(n1997) );
  AND U1593 ( .A(n2011), .B(n2012), .Z(n2010) );
  XOR U1594 ( .A(n2009), .B(n1835), .Z(n2012) );
  XOR U1595 ( .A(n2013), .B(n2014), .Z(n1835) );
  AND U1596 ( .A(n359), .B(n2015), .Z(n2014) );
  XOR U1597 ( .A(n2016), .B(n2013), .Z(n2015) );
  XNOR U1598 ( .A(n1832), .B(n2009), .Z(n2011) );
  XOR U1599 ( .A(n2017), .B(n2018), .Z(n1832) );
  AND U1600 ( .A(n357), .B(n2019), .Z(n2018) );
  XOR U1601 ( .A(n2020), .B(n2017), .Z(n2019) );
  XOR U1602 ( .A(n2021), .B(n2022), .Z(n2009) );
  AND U1603 ( .A(n2023), .B(n2024), .Z(n2022) );
  XOR U1604 ( .A(n2021), .B(n1847), .Z(n2024) );
  XOR U1605 ( .A(n2025), .B(n2026), .Z(n1847) );
  AND U1606 ( .A(n359), .B(n2027), .Z(n2026) );
  XOR U1607 ( .A(n2028), .B(n2025), .Z(n2027) );
  XNOR U1608 ( .A(n1844), .B(n2021), .Z(n2023) );
  XOR U1609 ( .A(n2029), .B(n2030), .Z(n1844) );
  AND U1610 ( .A(n357), .B(n2031), .Z(n2030) );
  XOR U1611 ( .A(n2032), .B(n2029), .Z(n2031) );
  XOR U1612 ( .A(n2033), .B(n2034), .Z(n2021) );
  AND U1613 ( .A(n2035), .B(n2036), .Z(n2034) );
  XOR U1614 ( .A(n2033), .B(n1859), .Z(n2036) );
  XOR U1615 ( .A(n2037), .B(n2038), .Z(n1859) );
  AND U1616 ( .A(n359), .B(n2039), .Z(n2038) );
  XOR U1617 ( .A(n2040), .B(n2037), .Z(n2039) );
  XNOR U1618 ( .A(n1856), .B(n2033), .Z(n2035) );
  XOR U1619 ( .A(n2041), .B(n2042), .Z(n1856) );
  AND U1620 ( .A(n357), .B(n2043), .Z(n2042) );
  XOR U1621 ( .A(n2044), .B(n2041), .Z(n2043) );
  XOR U1622 ( .A(n2045), .B(n2046), .Z(n2033) );
  AND U1623 ( .A(n2047), .B(n2048), .Z(n2046) );
  XOR U1624 ( .A(n2045), .B(n1871), .Z(n2048) );
  XOR U1625 ( .A(n2049), .B(n2050), .Z(n1871) );
  AND U1626 ( .A(n359), .B(n2051), .Z(n2050) );
  XOR U1627 ( .A(n2052), .B(n2049), .Z(n2051) );
  XNOR U1628 ( .A(n1868), .B(n2045), .Z(n2047) );
  XOR U1629 ( .A(n2053), .B(n2054), .Z(n1868) );
  AND U1630 ( .A(n357), .B(n2055), .Z(n2054) );
  XOR U1631 ( .A(n2056), .B(n2053), .Z(n2055) );
  XOR U1632 ( .A(n2057), .B(n2058), .Z(n2045) );
  AND U1633 ( .A(n2059), .B(n2060), .Z(n2058) );
  XOR U1634 ( .A(n2057), .B(n1883), .Z(n2060) );
  XOR U1635 ( .A(n2061), .B(n2062), .Z(n1883) );
  AND U1636 ( .A(n359), .B(n2063), .Z(n2062) );
  XOR U1637 ( .A(n2064), .B(n2061), .Z(n2063) );
  XNOR U1638 ( .A(n1880), .B(n2057), .Z(n2059) );
  XOR U1639 ( .A(n2065), .B(n2066), .Z(n1880) );
  AND U1640 ( .A(n357), .B(n2067), .Z(n2066) );
  XOR U1641 ( .A(n2068), .B(n2065), .Z(n2067) );
  XOR U1642 ( .A(n2069), .B(n2070), .Z(n2057) );
  AND U1643 ( .A(n2071), .B(n2072), .Z(n2070) );
  XOR U1644 ( .A(n2069), .B(n1895), .Z(n2072) );
  XOR U1645 ( .A(n2073), .B(n2074), .Z(n1895) );
  AND U1646 ( .A(n359), .B(n2075), .Z(n2074) );
  XOR U1647 ( .A(n2076), .B(n2073), .Z(n2075) );
  XNOR U1648 ( .A(n1892), .B(n2069), .Z(n2071) );
  XOR U1649 ( .A(n2077), .B(n2078), .Z(n1892) );
  AND U1650 ( .A(n357), .B(n2079), .Z(n2078) );
  XOR U1651 ( .A(n2080), .B(n2077), .Z(n2079) );
  XOR U1652 ( .A(n2081), .B(n2082), .Z(n2069) );
  AND U1653 ( .A(n2083), .B(n2084), .Z(n2082) );
  XOR U1654 ( .A(n2081), .B(n1907), .Z(n2084) );
  XOR U1655 ( .A(n2085), .B(n2086), .Z(n1907) );
  AND U1656 ( .A(n359), .B(n2087), .Z(n2086) );
  XOR U1657 ( .A(n2088), .B(n2085), .Z(n2087) );
  XNOR U1658 ( .A(n1904), .B(n2081), .Z(n2083) );
  XOR U1659 ( .A(n2089), .B(n2090), .Z(n1904) );
  AND U1660 ( .A(n357), .B(n2091), .Z(n2090) );
  XOR U1661 ( .A(n2092), .B(n2089), .Z(n2091) );
  XOR U1662 ( .A(n2093), .B(n2094), .Z(n2081) );
  AND U1663 ( .A(n2095), .B(n2096), .Z(n2094) );
  XOR U1664 ( .A(n2093), .B(n1919), .Z(n2096) );
  XOR U1665 ( .A(n2097), .B(n2098), .Z(n1919) );
  AND U1666 ( .A(n359), .B(n2099), .Z(n2098) );
  XOR U1667 ( .A(n2100), .B(n2097), .Z(n2099) );
  XNOR U1668 ( .A(n1916), .B(n2093), .Z(n2095) );
  XOR U1669 ( .A(n2101), .B(n2102), .Z(n1916) );
  AND U1670 ( .A(n357), .B(n2103), .Z(n2102) );
  XOR U1671 ( .A(n2104), .B(n2101), .Z(n2103) );
  XOR U1672 ( .A(n2105), .B(n2106), .Z(n2093) );
  AND U1673 ( .A(n2107), .B(n2108), .Z(n2106) );
  XOR U1674 ( .A(n2105), .B(n1931), .Z(n2108) );
  XOR U1675 ( .A(n2109), .B(n2110), .Z(n1931) );
  AND U1676 ( .A(n359), .B(n2111), .Z(n2110) );
  XOR U1677 ( .A(n2112), .B(n2109), .Z(n2111) );
  XNOR U1678 ( .A(n1928), .B(n2105), .Z(n2107) );
  XOR U1679 ( .A(n2113), .B(n2114), .Z(n1928) );
  AND U1680 ( .A(n357), .B(n2115), .Z(n2114) );
  XOR U1681 ( .A(n2116), .B(n2113), .Z(n2115) );
  XOR U1682 ( .A(n2117), .B(n2118), .Z(n2105) );
  AND U1683 ( .A(n2119), .B(n2120), .Z(n2118) );
  XOR U1684 ( .A(n2117), .B(n1943), .Z(n2120) );
  XOR U1685 ( .A(n2121), .B(n2122), .Z(n1943) );
  AND U1686 ( .A(n359), .B(n2123), .Z(n2122) );
  XOR U1687 ( .A(n2124), .B(n2121), .Z(n2123) );
  XNOR U1688 ( .A(n1940), .B(n2117), .Z(n2119) );
  XOR U1689 ( .A(n2125), .B(n2126), .Z(n1940) );
  AND U1690 ( .A(n357), .B(n2127), .Z(n2126) );
  XOR U1691 ( .A(n2128), .B(n2125), .Z(n2127) );
  XOR U1692 ( .A(n2129), .B(n2130), .Z(n2117) );
  AND U1693 ( .A(n2131), .B(n2132), .Z(n2130) );
  XOR U1694 ( .A(n2129), .B(n1955), .Z(n2132) );
  XOR U1695 ( .A(n2133), .B(n2134), .Z(n1955) );
  AND U1696 ( .A(n359), .B(n2135), .Z(n2134) );
  XOR U1697 ( .A(n2136), .B(n2133), .Z(n2135) );
  XNOR U1698 ( .A(n1952), .B(n2129), .Z(n2131) );
  XOR U1699 ( .A(n2137), .B(n2138), .Z(n1952) );
  AND U1700 ( .A(n357), .B(n2139), .Z(n2138) );
  XOR U1701 ( .A(n2140), .B(n2137), .Z(n2139) );
  XOR U1702 ( .A(n2141), .B(n2142), .Z(n2129) );
  AND U1703 ( .A(n2143), .B(n2144), .Z(n2142) );
  XOR U1704 ( .A(n2141), .B(n1967), .Z(n2144) );
  XOR U1705 ( .A(n2145), .B(n2146), .Z(n1967) );
  AND U1706 ( .A(n359), .B(n2147), .Z(n2146) );
  XOR U1707 ( .A(n2148), .B(n2145), .Z(n2147) );
  XNOR U1708 ( .A(n1964), .B(n2141), .Z(n2143) );
  XOR U1709 ( .A(n2149), .B(n2150), .Z(n1964) );
  AND U1710 ( .A(n357), .B(n2151), .Z(n2150) );
  XOR U1711 ( .A(n2152), .B(n2149), .Z(n2151) );
  XOR U1712 ( .A(n2153), .B(n2154), .Z(n2141) );
  AND U1713 ( .A(n2155), .B(n2156), .Z(n2154) );
  XNOR U1714 ( .A(n2157), .B(n1980), .Z(n2156) );
  XOR U1715 ( .A(n2158), .B(n2159), .Z(n1980) );
  AND U1716 ( .A(n359), .B(n2160), .Z(n2159) );
  XOR U1717 ( .A(n2158), .B(n2161), .Z(n2160) );
  XNOR U1718 ( .A(n1977), .B(n2153), .Z(n2155) );
  XOR U1719 ( .A(n2162), .B(n2163), .Z(n1977) );
  AND U1720 ( .A(n357), .B(n2164), .Z(n2163) );
  XOR U1721 ( .A(n2162), .B(n2165), .Z(n2164) );
  IV U1722 ( .A(n2157), .Z(n2153) );
  AND U1723 ( .A(n1985), .B(n1988), .Z(n2157) );
  XNOR U1724 ( .A(n2166), .B(n2167), .Z(n1988) );
  AND U1725 ( .A(n359), .B(n2168), .Z(n2167) );
  XNOR U1726 ( .A(n2169), .B(n2166), .Z(n2168) );
  XOR U1727 ( .A(n2170), .B(n2171), .Z(n359) );
  AND U1728 ( .A(n2172), .B(n2173), .Z(n2171) );
  XNOR U1729 ( .A(n1993), .B(n2170), .Z(n2173) );
  AND U1730 ( .A(p_input[4095]), .B(p_input[4079]), .Z(n1993) );
  XOR U1731 ( .A(n2170), .B(n1994), .Z(n2172) );
  AND U1732 ( .A(p_input[4063]), .B(p_input[4047]), .Z(n1994) );
  XOR U1733 ( .A(n2174), .B(n2175), .Z(n2170) );
  AND U1734 ( .A(n2176), .B(n2177), .Z(n2175) );
  XOR U1735 ( .A(n2174), .B(n2004), .Z(n2177) );
  XNOR U1736 ( .A(p_input[4078]), .B(n2178), .Z(n2004) );
  AND U1737 ( .A(n107), .B(n2179), .Z(n2178) );
  XOR U1738 ( .A(p_input[4094]), .B(p_input[4078]), .Z(n2179) );
  XNOR U1739 ( .A(n2001), .B(n2174), .Z(n2176) );
  XOR U1740 ( .A(n2180), .B(n2181), .Z(n2001) );
  AND U1741 ( .A(n105), .B(n2182), .Z(n2181) );
  XOR U1742 ( .A(p_input[4062]), .B(p_input[4046]), .Z(n2182) );
  XOR U1743 ( .A(n2183), .B(n2184), .Z(n2174) );
  AND U1744 ( .A(n2185), .B(n2186), .Z(n2184) );
  XOR U1745 ( .A(n2183), .B(n2016), .Z(n2186) );
  XNOR U1746 ( .A(p_input[4077]), .B(n2187), .Z(n2016) );
  AND U1747 ( .A(n107), .B(n2188), .Z(n2187) );
  XOR U1748 ( .A(p_input[4093]), .B(p_input[4077]), .Z(n2188) );
  XNOR U1749 ( .A(n2013), .B(n2183), .Z(n2185) );
  XOR U1750 ( .A(n2189), .B(n2190), .Z(n2013) );
  AND U1751 ( .A(n105), .B(n2191), .Z(n2190) );
  XOR U1752 ( .A(p_input[4061]), .B(p_input[4045]), .Z(n2191) );
  XOR U1753 ( .A(n2192), .B(n2193), .Z(n2183) );
  AND U1754 ( .A(n2194), .B(n2195), .Z(n2193) );
  XOR U1755 ( .A(n2192), .B(n2028), .Z(n2195) );
  XNOR U1756 ( .A(p_input[4076]), .B(n2196), .Z(n2028) );
  AND U1757 ( .A(n107), .B(n2197), .Z(n2196) );
  XOR U1758 ( .A(p_input[4092]), .B(p_input[4076]), .Z(n2197) );
  XNOR U1759 ( .A(n2025), .B(n2192), .Z(n2194) );
  XOR U1760 ( .A(n2198), .B(n2199), .Z(n2025) );
  AND U1761 ( .A(n105), .B(n2200), .Z(n2199) );
  XOR U1762 ( .A(p_input[4060]), .B(p_input[4044]), .Z(n2200) );
  XOR U1763 ( .A(n2201), .B(n2202), .Z(n2192) );
  AND U1764 ( .A(n2203), .B(n2204), .Z(n2202) );
  XOR U1765 ( .A(n2201), .B(n2040), .Z(n2204) );
  XNOR U1766 ( .A(p_input[4075]), .B(n2205), .Z(n2040) );
  AND U1767 ( .A(n107), .B(n2206), .Z(n2205) );
  XOR U1768 ( .A(p_input[4091]), .B(p_input[4075]), .Z(n2206) );
  XNOR U1769 ( .A(n2037), .B(n2201), .Z(n2203) );
  XOR U1770 ( .A(n2207), .B(n2208), .Z(n2037) );
  AND U1771 ( .A(n105), .B(n2209), .Z(n2208) );
  XOR U1772 ( .A(p_input[4059]), .B(p_input[4043]), .Z(n2209) );
  XOR U1773 ( .A(n2210), .B(n2211), .Z(n2201) );
  AND U1774 ( .A(n2212), .B(n2213), .Z(n2211) );
  XOR U1775 ( .A(n2210), .B(n2052), .Z(n2213) );
  XNOR U1776 ( .A(p_input[4074]), .B(n2214), .Z(n2052) );
  AND U1777 ( .A(n107), .B(n2215), .Z(n2214) );
  XOR U1778 ( .A(p_input[4090]), .B(p_input[4074]), .Z(n2215) );
  XNOR U1779 ( .A(n2049), .B(n2210), .Z(n2212) );
  XOR U1780 ( .A(n2216), .B(n2217), .Z(n2049) );
  AND U1781 ( .A(n105), .B(n2218), .Z(n2217) );
  XOR U1782 ( .A(p_input[4058]), .B(p_input[4042]), .Z(n2218) );
  XOR U1783 ( .A(n2219), .B(n2220), .Z(n2210) );
  AND U1784 ( .A(n2221), .B(n2222), .Z(n2220) );
  XOR U1785 ( .A(n2219), .B(n2064), .Z(n2222) );
  XNOR U1786 ( .A(p_input[4073]), .B(n2223), .Z(n2064) );
  AND U1787 ( .A(n107), .B(n2224), .Z(n2223) );
  XOR U1788 ( .A(p_input[4089]), .B(p_input[4073]), .Z(n2224) );
  XNOR U1789 ( .A(n2061), .B(n2219), .Z(n2221) );
  XOR U1790 ( .A(n2225), .B(n2226), .Z(n2061) );
  AND U1791 ( .A(n105), .B(n2227), .Z(n2226) );
  XOR U1792 ( .A(p_input[4057]), .B(p_input[4041]), .Z(n2227) );
  XOR U1793 ( .A(n2228), .B(n2229), .Z(n2219) );
  AND U1794 ( .A(n2230), .B(n2231), .Z(n2229) );
  XOR U1795 ( .A(n2228), .B(n2076), .Z(n2231) );
  XNOR U1796 ( .A(p_input[4072]), .B(n2232), .Z(n2076) );
  AND U1797 ( .A(n107), .B(n2233), .Z(n2232) );
  XOR U1798 ( .A(p_input[4088]), .B(p_input[4072]), .Z(n2233) );
  XNOR U1799 ( .A(n2073), .B(n2228), .Z(n2230) );
  XOR U1800 ( .A(n2234), .B(n2235), .Z(n2073) );
  AND U1801 ( .A(n105), .B(n2236), .Z(n2235) );
  XOR U1802 ( .A(p_input[4056]), .B(p_input[4040]), .Z(n2236) );
  XOR U1803 ( .A(n2237), .B(n2238), .Z(n2228) );
  AND U1804 ( .A(n2239), .B(n2240), .Z(n2238) );
  XOR U1805 ( .A(n2237), .B(n2088), .Z(n2240) );
  XNOR U1806 ( .A(p_input[4071]), .B(n2241), .Z(n2088) );
  AND U1807 ( .A(n107), .B(n2242), .Z(n2241) );
  XOR U1808 ( .A(p_input[4087]), .B(p_input[4071]), .Z(n2242) );
  XNOR U1809 ( .A(n2085), .B(n2237), .Z(n2239) );
  XOR U1810 ( .A(n2243), .B(n2244), .Z(n2085) );
  AND U1811 ( .A(n105), .B(n2245), .Z(n2244) );
  XOR U1812 ( .A(p_input[4055]), .B(p_input[4039]), .Z(n2245) );
  XOR U1813 ( .A(n2246), .B(n2247), .Z(n2237) );
  AND U1814 ( .A(n2248), .B(n2249), .Z(n2247) );
  XOR U1815 ( .A(n2246), .B(n2100), .Z(n2249) );
  XNOR U1816 ( .A(p_input[4070]), .B(n2250), .Z(n2100) );
  AND U1817 ( .A(n107), .B(n2251), .Z(n2250) );
  XOR U1818 ( .A(p_input[4086]), .B(p_input[4070]), .Z(n2251) );
  XNOR U1819 ( .A(n2097), .B(n2246), .Z(n2248) );
  XOR U1820 ( .A(n2252), .B(n2253), .Z(n2097) );
  AND U1821 ( .A(n105), .B(n2254), .Z(n2253) );
  XOR U1822 ( .A(p_input[4054]), .B(p_input[4038]), .Z(n2254) );
  XOR U1823 ( .A(n2255), .B(n2256), .Z(n2246) );
  AND U1824 ( .A(n2257), .B(n2258), .Z(n2256) );
  XOR U1825 ( .A(n2255), .B(n2112), .Z(n2258) );
  XNOR U1826 ( .A(p_input[4069]), .B(n2259), .Z(n2112) );
  AND U1827 ( .A(n107), .B(n2260), .Z(n2259) );
  XOR U1828 ( .A(p_input[4085]), .B(p_input[4069]), .Z(n2260) );
  XNOR U1829 ( .A(n2109), .B(n2255), .Z(n2257) );
  XOR U1830 ( .A(n2261), .B(n2262), .Z(n2109) );
  AND U1831 ( .A(n105), .B(n2263), .Z(n2262) );
  XOR U1832 ( .A(p_input[4053]), .B(p_input[4037]), .Z(n2263) );
  XOR U1833 ( .A(n2264), .B(n2265), .Z(n2255) );
  AND U1834 ( .A(n2266), .B(n2267), .Z(n2265) );
  XOR U1835 ( .A(n2264), .B(n2124), .Z(n2267) );
  XNOR U1836 ( .A(p_input[4068]), .B(n2268), .Z(n2124) );
  AND U1837 ( .A(n107), .B(n2269), .Z(n2268) );
  XOR U1838 ( .A(p_input[4084]), .B(p_input[4068]), .Z(n2269) );
  XNOR U1839 ( .A(n2121), .B(n2264), .Z(n2266) );
  XOR U1840 ( .A(n2270), .B(n2271), .Z(n2121) );
  AND U1841 ( .A(n105), .B(n2272), .Z(n2271) );
  XOR U1842 ( .A(p_input[4052]), .B(p_input[4036]), .Z(n2272) );
  XOR U1843 ( .A(n2273), .B(n2274), .Z(n2264) );
  AND U1844 ( .A(n2275), .B(n2276), .Z(n2274) );
  XOR U1845 ( .A(n2273), .B(n2136), .Z(n2276) );
  XNOR U1846 ( .A(p_input[4067]), .B(n2277), .Z(n2136) );
  AND U1847 ( .A(n107), .B(n2278), .Z(n2277) );
  XOR U1848 ( .A(p_input[4083]), .B(p_input[4067]), .Z(n2278) );
  XNOR U1849 ( .A(n2133), .B(n2273), .Z(n2275) );
  XOR U1850 ( .A(n2279), .B(n2280), .Z(n2133) );
  AND U1851 ( .A(n105), .B(n2281), .Z(n2280) );
  XOR U1852 ( .A(p_input[4051]), .B(p_input[4035]), .Z(n2281) );
  XOR U1853 ( .A(n2282), .B(n2283), .Z(n2273) );
  AND U1854 ( .A(n2284), .B(n2285), .Z(n2283) );
  XOR U1855 ( .A(n2282), .B(n2148), .Z(n2285) );
  XNOR U1856 ( .A(p_input[4066]), .B(n2286), .Z(n2148) );
  AND U1857 ( .A(n107), .B(n2287), .Z(n2286) );
  XOR U1858 ( .A(p_input[4082]), .B(p_input[4066]), .Z(n2287) );
  XNOR U1859 ( .A(n2145), .B(n2282), .Z(n2284) );
  XOR U1860 ( .A(n2288), .B(n2289), .Z(n2145) );
  AND U1861 ( .A(n105), .B(n2290), .Z(n2289) );
  XOR U1862 ( .A(p_input[4050]), .B(p_input[4034]), .Z(n2290) );
  XOR U1863 ( .A(n2291), .B(n2292), .Z(n2282) );
  AND U1864 ( .A(n2293), .B(n2294), .Z(n2292) );
  XNOR U1865 ( .A(n2295), .B(n2161), .Z(n2294) );
  XNOR U1866 ( .A(p_input[4065]), .B(n2296), .Z(n2161) );
  AND U1867 ( .A(n107), .B(n2297), .Z(n2296) );
  XNOR U1868 ( .A(p_input[4081]), .B(n2298), .Z(n2297) );
  IV U1869 ( .A(p_input[4065]), .Z(n2298) );
  XNOR U1870 ( .A(n2158), .B(n2291), .Z(n2293) );
  XNOR U1871 ( .A(p_input[4033]), .B(n2299), .Z(n2158) );
  AND U1872 ( .A(n105), .B(n2300), .Z(n2299) );
  XOR U1873 ( .A(p_input[4049]), .B(p_input[4033]), .Z(n2300) );
  IV U1874 ( .A(n2295), .Z(n2291) );
  AND U1875 ( .A(n2166), .B(n2169), .Z(n2295) );
  XOR U1876 ( .A(p_input[4064]), .B(n2301), .Z(n2169) );
  AND U1877 ( .A(n107), .B(n2302), .Z(n2301) );
  XOR U1878 ( .A(p_input[4080]), .B(p_input[4064]), .Z(n2302) );
  XOR U1879 ( .A(n2303), .B(n2304), .Z(n107) );
  AND U1880 ( .A(n2305), .B(n2306), .Z(n2304) );
  XNOR U1881 ( .A(p_input[4095]), .B(n2303), .Z(n2306) );
  XOR U1882 ( .A(n2303), .B(p_input[4079]), .Z(n2305) );
  XOR U1883 ( .A(n2307), .B(n2308), .Z(n2303) );
  AND U1884 ( .A(n2309), .B(n2310), .Z(n2308) );
  XNOR U1885 ( .A(p_input[4094]), .B(n2307), .Z(n2310) );
  XOR U1886 ( .A(n2307), .B(p_input[4078]), .Z(n2309) );
  XOR U1887 ( .A(n2311), .B(n2312), .Z(n2307) );
  AND U1888 ( .A(n2313), .B(n2314), .Z(n2312) );
  XNOR U1889 ( .A(p_input[4093]), .B(n2311), .Z(n2314) );
  XOR U1890 ( .A(n2311), .B(p_input[4077]), .Z(n2313) );
  XOR U1891 ( .A(n2315), .B(n2316), .Z(n2311) );
  AND U1892 ( .A(n2317), .B(n2318), .Z(n2316) );
  XNOR U1893 ( .A(p_input[4092]), .B(n2315), .Z(n2318) );
  XOR U1894 ( .A(n2315), .B(p_input[4076]), .Z(n2317) );
  XOR U1895 ( .A(n2319), .B(n2320), .Z(n2315) );
  AND U1896 ( .A(n2321), .B(n2322), .Z(n2320) );
  XNOR U1897 ( .A(p_input[4091]), .B(n2319), .Z(n2322) );
  XOR U1898 ( .A(n2319), .B(p_input[4075]), .Z(n2321) );
  XOR U1899 ( .A(n2323), .B(n2324), .Z(n2319) );
  AND U1900 ( .A(n2325), .B(n2326), .Z(n2324) );
  XNOR U1901 ( .A(p_input[4090]), .B(n2323), .Z(n2326) );
  XOR U1902 ( .A(n2323), .B(p_input[4074]), .Z(n2325) );
  XOR U1903 ( .A(n2327), .B(n2328), .Z(n2323) );
  AND U1904 ( .A(n2329), .B(n2330), .Z(n2328) );
  XNOR U1905 ( .A(p_input[4089]), .B(n2327), .Z(n2330) );
  XOR U1906 ( .A(n2327), .B(p_input[4073]), .Z(n2329) );
  XOR U1907 ( .A(n2331), .B(n2332), .Z(n2327) );
  AND U1908 ( .A(n2333), .B(n2334), .Z(n2332) );
  XNOR U1909 ( .A(p_input[4088]), .B(n2331), .Z(n2334) );
  XOR U1910 ( .A(n2331), .B(p_input[4072]), .Z(n2333) );
  XOR U1911 ( .A(n2335), .B(n2336), .Z(n2331) );
  AND U1912 ( .A(n2337), .B(n2338), .Z(n2336) );
  XNOR U1913 ( .A(p_input[4087]), .B(n2335), .Z(n2338) );
  XOR U1914 ( .A(n2335), .B(p_input[4071]), .Z(n2337) );
  XOR U1915 ( .A(n2339), .B(n2340), .Z(n2335) );
  AND U1916 ( .A(n2341), .B(n2342), .Z(n2340) );
  XNOR U1917 ( .A(p_input[4086]), .B(n2339), .Z(n2342) );
  XOR U1918 ( .A(n2339), .B(p_input[4070]), .Z(n2341) );
  XOR U1919 ( .A(n2343), .B(n2344), .Z(n2339) );
  AND U1920 ( .A(n2345), .B(n2346), .Z(n2344) );
  XNOR U1921 ( .A(p_input[4085]), .B(n2343), .Z(n2346) );
  XOR U1922 ( .A(n2343), .B(p_input[4069]), .Z(n2345) );
  XOR U1923 ( .A(n2347), .B(n2348), .Z(n2343) );
  AND U1924 ( .A(n2349), .B(n2350), .Z(n2348) );
  XNOR U1925 ( .A(p_input[4084]), .B(n2347), .Z(n2350) );
  XOR U1926 ( .A(n2347), .B(p_input[4068]), .Z(n2349) );
  XOR U1927 ( .A(n2351), .B(n2352), .Z(n2347) );
  AND U1928 ( .A(n2353), .B(n2354), .Z(n2352) );
  XNOR U1929 ( .A(p_input[4083]), .B(n2351), .Z(n2354) );
  XOR U1930 ( .A(n2351), .B(p_input[4067]), .Z(n2353) );
  XOR U1931 ( .A(n2355), .B(n2356), .Z(n2351) );
  AND U1932 ( .A(n2357), .B(n2358), .Z(n2356) );
  XNOR U1933 ( .A(p_input[4082]), .B(n2355), .Z(n2358) );
  XOR U1934 ( .A(n2355), .B(p_input[4066]), .Z(n2357) );
  XNOR U1935 ( .A(n2359), .B(n2360), .Z(n2355) );
  AND U1936 ( .A(n2361), .B(n2362), .Z(n2360) );
  XOR U1937 ( .A(p_input[4081]), .B(n2359), .Z(n2362) );
  XNOR U1938 ( .A(p_input[4065]), .B(n2359), .Z(n2361) );
  AND U1939 ( .A(p_input[4080]), .B(n2363), .Z(n2359) );
  IV U1940 ( .A(p_input[4064]), .Z(n2363) );
  XNOR U1941 ( .A(p_input[4032]), .B(n2364), .Z(n2166) );
  AND U1942 ( .A(n105), .B(n2365), .Z(n2364) );
  XOR U1943 ( .A(p_input[4048]), .B(p_input[4032]), .Z(n2365) );
  XOR U1944 ( .A(n2366), .B(n2367), .Z(n105) );
  AND U1945 ( .A(n2368), .B(n2369), .Z(n2367) );
  XNOR U1946 ( .A(p_input[4063]), .B(n2366), .Z(n2369) );
  XOR U1947 ( .A(n2366), .B(p_input[4047]), .Z(n2368) );
  XOR U1948 ( .A(n2370), .B(n2371), .Z(n2366) );
  AND U1949 ( .A(n2372), .B(n2373), .Z(n2371) );
  XNOR U1950 ( .A(p_input[4062]), .B(n2370), .Z(n2373) );
  XNOR U1951 ( .A(n2370), .B(n2180), .Z(n2372) );
  IV U1952 ( .A(p_input[4046]), .Z(n2180) );
  XOR U1953 ( .A(n2374), .B(n2375), .Z(n2370) );
  AND U1954 ( .A(n2376), .B(n2377), .Z(n2375) );
  XNOR U1955 ( .A(p_input[4061]), .B(n2374), .Z(n2377) );
  XNOR U1956 ( .A(n2374), .B(n2189), .Z(n2376) );
  IV U1957 ( .A(p_input[4045]), .Z(n2189) );
  XOR U1958 ( .A(n2378), .B(n2379), .Z(n2374) );
  AND U1959 ( .A(n2380), .B(n2381), .Z(n2379) );
  XNOR U1960 ( .A(p_input[4060]), .B(n2378), .Z(n2381) );
  XNOR U1961 ( .A(n2378), .B(n2198), .Z(n2380) );
  IV U1962 ( .A(p_input[4044]), .Z(n2198) );
  XOR U1963 ( .A(n2382), .B(n2383), .Z(n2378) );
  AND U1964 ( .A(n2384), .B(n2385), .Z(n2383) );
  XNOR U1965 ( .A(p_input[4059]), .B(n2382), .Z(n2385) );
  XNOR U1966 ( .A(n2382), .B(n2207), .Z(n2384) );
  IV U1967 ( .A(p_input[4043]), .Z(n2207) );
  XOR U1968 ( .A(n2386), .B(n2387), .Z(n2382) );
  AND U1969 ( .A(n2388), .B(n2389), .Z(n2387) );
  XNOR U1970 ( .A(p_input[4058]), .B(n2386), .Z(n2389) );
  XNOR U1971 ( .A(n2386), .B(n2216), .Z(n2388) );
  IV U1972 ( .A(p_input[4042]), .Z(n2216) );
  XOR U1973 ( .A(n2390), .B(n2391), .Z(n2386) );
  AND U1974 ( .A(n2392), .B(n2393), .Z(n2391) );
  XNOR U1975 ( .A(p_input[4057]), .B(n2390), .Z(n2393) );
  XNOR U1976 ( .A(n2390), .B(n2225), .Z(n2392) );
  IV U1977 ( .A(p_input[4041]), .Z(n2225) );
  XOR U1978 ( .A(n2394), .B(n2395), .Z(n2390) );
  AND U1979 ( .A(n2396), .B(n2397), .Z(n2395) );
  XNOR U1980 ( .A(p_input[4056]), .B(n2394), .Z(n2397) );
  XNOR U1981 ( .A(n2394), .B(n2234), .Z(n2396) );
  IV U1982 ( .A(p_input[4040]), .Z(n2234) );
  XOR U1983 ( .A(n2398), .B(n2399), .Z(n2394) );
  AND U1984 ( .A(n2400), .B(n2401), .Z(n2399) );
  XNOR U1985 ( .A(p_input[4055]), .B(n2398), .Z(n2401) );
  XNOR U1986 ( .A(n2398), .B(n2243), .Z(n2400) );
  IV U1987 ( .A(p_input[4039]), .Z(n2243) );
  XOR U1988 ( .A(n2402), .B(n2403), .Z(n2398) );
  AND U1989 ( .A(n2404), .B(n2405), .Z(n2403) );
  XNOR U1990 ( .A(p_input[4054]), .B(n2402), .Z(n2405) );
  XNOR U1991 ( .A(n2402), .B(n2252), .Z(n2404) );
  IV U1992 ( .A(p_input[4038]), .Z(n2252) );
  XOR U1993 ( .A(n2406), .B(n2407), .Z(n2402) );
  AND U1994 ( .A(n2408), .B(n2409), .Z(n2407) );
  XNOR U1995 ( .A(p_input[4053]), .B(n2406), .Z(n2409) );
  XNOR U1996 ( .A(n2406), .B(n2261), .Z(n2408) );
  IV U1997 ( .A(p_input[4037]), .Z(n2261) );
  XOR U1998 ( .A(n2410), .B(n2411), .Z(n2406) );
  AND U1999 ( .A(n2412), .B(n2413), .Z(n2411) );
  XNOR U2000 ( .A(p_input[4052]), .B(n2410), .Z(n2413) );
  XNOR U2001 ( .A(n2410), .B(n2270), .Z(n2412) );
  IV U2002 ( .A(p_input[4036]), .Z(n2270) );
  XOR U2003 ( .A(n2414), .B(n2415), .Z(n2410) );
  AND U2004 ( .A(n2416), .B(n2417), .Z(n2415) );
  XNOR U2005 ( .A(p_input[4051]), .B(n2414), .Z(n2417) );
  XNOR U2006 ( .A(n2414), .B(n2279), .Z(n2416) );
  IV U2007 ( .A(p_input[4035]), .Z(n2279) );
  XOR U2008 ( .A(n2418), .B(n2419), .Z(n2414) );
  AND U2009 ( .A(n2420), .B(n2421), .Z(n2419) );
  XNOR U2010 ( .A(p_input[4050]), .B(n2418), .Z(n2421) );
  XNOR U2011 ( .A(n2418), .B(n2288), .Z(n2420) );
  IV U2012 ( .A(p_input[4034]), .Z(n2288) );
  XNOR U2013 ( .A(n2422), .B(n2423), .Z(n2418) );
  AND U2014 ( .A(n2424), .B(n2425), .Z(n2423) );
  XOR U2015 ( .A(p_input[4049]), .B(n2422), .Z(n2425) );
  XNOR U2016 ( .A(p_input[4033]), .B(n2422), .Z(n2424) );
  AND U2017 ( .A(p_input[4048]), .B(n2426), .Z(n2422) );
  IV U2018 ( .A(p_input[4032]), .Z(n2426) );
  XOR U2019 ( .A(n2427), .B(n2428), .Z(n1985) );
  AND U2020 ( .A(n357), .B(n2429), .Z(n2428) );
  XNOR U2021 ( .A(n2430), .B(n2427), .Z(n2429) );
  XOR U2022 ( .A(n2431), .B(n2432), .Z(n357) );
  AND U2023 ( .A(n2433), .B(n2434), .Z(n2432) );
  XNOR U2024 ( .A(n1995), .B(n2431), .Z(n2434) );
  AND U2025 ( .A(p_input[4031]), .B(p_input[4015]), .Z(n1995) );
  XOR U2026 ( .A(n2431), .B(n1996), .Z(n2433) );
  AND U2027 ( .A(p_input[3999]), .B(p_input[3983]), .Z(n1996) );
  XOR U2028 ( .A(n2435), .B(n2436), .Z(n2431) );
  AND U2029 ( .A(n2437), .B(n2438), .Z(n2436) );
  XOR U2030 ( .A(n2435), .B(n2008), .Z(n2438) );
  XNOR U2031 ( .A(p_input[4014]), .B(n2439), .Z(n2008) );
  AND U2032 ( .A(n111), .B(n2440), .Z(n2439) );
  XOR U2033 ( .A(p_input[4030]), .B(p_input[4014]), .Z(n2440) );
  XNOR U2034 ( .A(n2005), .B(n2435), .Z(n2437) );
  XOR U2035 ( .A(n2441), .B(n2442), .Z(n2005) );
  AND U2036 ( .A(n108), .B(n2443), .Z(n2442) );
  XOR U2037 ( .A(p_input[3998]), .B(p_input[3982]), .Z(n2443) );
  XOR U2038 ( .A(n2444), .B(n2445), .Z(n2435) );
  AND U2039 ( .A(n2446), .B(n2447), .Z(n2445) );
  XOR U2040 ( .A(n2444), .B(n2020), .Z(n2447) );
  XNOR U2041 ( .A(p_input[4013]), .B(n2448), .Z(n2020) );
  AND U2042 ( .A(n111), .B(n2449), .Z(n2448) );
  XOR U2043 ( .A(p_input[4029]), .B(p_input[4013]), .Z(n2449) );
  XNOR U2044 ( .A(n2017), .B(n2444), .Z(n2446) );
  XOR U2045 ( .A(n2450), .B(n2451), .Z(n2017) );
  AND U2046 ( .A(n108), .B(n2452), .Z(n2451) );
  XOR U2047 ( .A(p_input[3997]), .B(p_input[3981]), .Z(n2452) );
  XOR U2048 ( .A(n2453), .B(n2454), .Z(n2444) );
  AND U2049 ( .A(n2455), .B(n2456), .Z(n2454) );
  XOR U2050 ( .A(n2453), .B(n2032), .Z(n2456) );
  XNOR U2051 ( .A(p_input[4012]), .B(n2457), .Z(n2032) );
  AND U2052 ( .A(n111), .B(n2458), .Z(n2457) );
  XOR U2053 ( .A(p_input[4028]), .B(p_input[4012]), .Z(n2458) );
  XNOR U2054 ( .A(n2029), .B(n2453), .Z(n2455) );
  XOR U2055 ( .A(n2459), .B(n2460), .Z(n2029) );
  AND U2056 ( .A(n108), .B(n2461), .Z(n2460) );
  XOR U2057 ( .A(p_input[3996]), .B(p_input[3980]), .Z(n2461) );
  XOR U2058 ( .A(n2462), .B(n2463), .Z(n2453) );
  AND U2059 ( .A(n2464), .B(n2465), .Z(n2463) );
  XOR U2060 ( .A(n2462), .B(n2044), .Z(n2465) );
  XNOR U2061 ( .A(p_input[4011]), .B(n2466), .Z(n2044) );
  AND U2062 ( .A(n111), .B(n2467), .Z(n2466) );
  XOR U2063 ( .A(p_input[4027]), .B(p_input[4011]), .Z(n2467) );
  XNOR U2064 ( .A(n2041), .B(n2462), .Z(n2464) );
  XOR U2065 ( .A(n2468), .B(n2469), .Z(n2041) );
  AND U2066 ( .A(n108), .B(n2470), .Z(n2469) );
  XOR U2067 ( .A(p_input[3995]), .B(p_input[3979]), .Z(n2470) );
  XOR U2068 ( .A(n2471), .B(n2472), .Z(n2462) );
  AND U2069 ( .A(n2473), .B(n2474), .Z(n2472) );
  XOR U2070 ( .A(n2471), .B(n2056), .Z(n2474) );
  XNOR U2071 ( .A(p_input[4010]), .B(n2475), .Z(n2056) );
  AND U2072 ( .A(n111), .B(n2476), .Z(n2475) );
  XOR U2073 ( .A(p_input[4026]), .B(p_input[4010]), .Z(n2476) );
  XNOR U2074 ( .A(n2053), .B(n2471), .Z(n2473) );
  XOR U2075 ( .A(n2477), .B(n2478), .Z(n2053) );
  AND U2076 ( .A(n108), .B(n2479), .Z(n2478) );
  XOR U2077 ( .A(p_input[3994]), .B(p_input[3978]), .Z(n2479) );
  XOR U2078 ( .A(n2480), .B(n2481), .Z(n2471) );
  AND U2079 ( .A(n2482), .B(n2483), .Z(n2481) );
  XOR U2080 ( .A(n2480), .B(n2068), .Z(n2483) );
  XNOR U2081 ( .A(p_input[4009]), .B(n2484), .Z(n2068) );
  AND U2082 ( .A(n111), .B(n2485), .Z(n2484) );
  XOR U2083 ( .A(p_input[4025]), .B(p_input[4009]), .Z(n2485) );
  XNOR U2084 ( .A(n2065), .B(n2480), .Z(n2482) );
  XOR U2085 ( .A(n2486), .B(n2487), .Z(n2065) );
  AND U2086 ( .A(n108), .B(n2488), .Z(n2487) );
  XOR U2087 ( .A(p_input[3993]), .B(p_input[3977]), .Z(n2488) );
  XOR U2088 ( .A(n2489), .B(n2490), .Z(n2480) );
  AND U2089 ( .A(n2491), .B(n2492), .Z(n2490) );
  XOR U2090 ( .A(n2489), .B(n2080), .Z(n2492) );
  XNOR U2091 ( .A(p_input[4008]), .B(n2493), .Z(n2080) );
  AND U2092 ( .A(n111), .B(n2494), .Z(n2493) );
  XOR U2093 ( .A(p_input[4024]), .B(p_input[4008]), .Z(n2494) );
  XNOR U2094 ( .A(n2077), .B(n2489), .Z(n2491) );
  XOR U2095 ( .A(n2495), .B(n2496), .Z(n2077) );
  AND U2096 ( .A(n108), .B(n2497), .Z(n2496) );
  XOR U2097 ( .A(p_input[3992]), .B(p_input[3976]), .Z(n2497) );
  XOR U2098 ( .A(n2498), .B(n2499), .Z(n2489) );
  AND U2099 ( .A(n2500), .B(n2501), .Z(n2499) );
  XOR U2100 ( .A(n2498), .B(n2092), .Z(n2501) );
  XNOR U2101 ( .A(p_input[4007]), .B(n2502), .Z(n2092) );
  AND U2102 ( .A(n111), .B(n2503), .Z(n2502) );
  XOR U2103 ( .A(p_input[4023]), .B(p_input[4007]), .Z(n2503) );
  XNOR U2104 ( .A(n2089), .B(n2498), .Z(n2500) );
  XOR U2105 ( .A(n2504), .B(n2505), .Z(n2089) );
  AND U2106 ( .A(n108), .B(n2506), .Z(n2505) );
  XOR U2107 ( .A(p_input[3991]), .B(p_input[3975]), .Z(n2506) );
  XOR U2108 ( .A(n2507), .B(n2508), .Z(n2498) );
  AND U2109 ( .A(n2509), .B(n2510), .Z(n2508) );
  XOR U2110 ( .A(n2507), .B(n2104), .Z(n2510) );
  XNOR U2111 ( .A(p_input[4006]), .B(n2511), .Z(n2104) );
  AND U2112 ( .A(n111), .B(n2512), .Z(n2511) );
  XOR U2113 ( .A(p_input[4022]), .B(p_input[4006]), .Z(n2512) );
  XNOR U2114 ( .A(n2101), .B(n2507), .Z(n2509) );
  XOR U2115 ( .A(n2513), .B(n2514), .Z(n2101) );
  AND U2116 ( .A(n108), .B(n2515), .Z(n2514) );
  XOR U2117 ( .A(p_input[3990]), .B(p_input[3974]), .Z(n2515) );
  XOR U2118 ( .A(n2516), .B(n2517), .Z(n2507) );
  AND U2119 ( .A(n2518), .B(n2519), .Z(n2517) );
  XOR U2120 ( .A(n2516), .B(n2116), .Z(n2519) );
  XNOR U2121 ( .A(p_input[4005]), .B(n2520), .Z(n2116) );
  AND U2122 ( .A(n111), .B(n2521), .Z(n2520) );
  XOR U2123 ( .A(p_input[4021]), .B(p_input[4005]), .Z(n2521) );
  XNOR U2124 ( .A(n2113), .B(n2516), .Z(n2518) );
  XOR U2125 ( .A(n2522), .B(n2523), .Z(n2113) );
  AND U2126 ( .A(n108), .B(n2524), .Z(n2523) );
  XOR U2127 ( .A(p_input[3989]), .B(p_input[3973]), .Z(n2524) );
  XOR U2128 ( .A(n2525), .B(n2526), .Z(n2516) );
  AND U2129 ( .A(n2527), .B(n2528), .Z(n2526) );
  XOR U2130 ( .A(n2525), .B(n2128), .Z(n2528) );
  XNOR U2131 ( .A(p_input[4004]), .B(n2529), .Z(n2128) );
  AND U2132 ( .A(n111), .B(n2530), .Z(n2529) );
  XOR U2133 ( .A(p_input[4020]), .B(p_input[4004]), .Z(n2530) );
  XNOR U2134 ( .A(n2125), .B(n2525), .Z(n2527) );
  XOR U2135 ( .A(n2531), .B(n2532), .Z(n2125) );
  AND U2136 ( .A(n108), .B(n2533), .Z(n2532) );
  XOR U2137 ( .A(p_input[3988]), .B(p_input[3972]), .Z(n2533) );
  XOR U2138 ( .A(n2534), .B(n2535), .Z(n2525) );
  AND U2139 ( .A(n2536), .B(n2537), .Z(n2535) );
  XOR U2140 ( .A(n2534), .B(n2140), .Z(n2537) );
  XNOR U2141 ( .A(p_input[4003]), .B(n2538), .Z(n2140) );
  AND U2142 ( .A(n111), .B(n2539), .Z(n2538) );
  XOR U2143 ( .A(p_input[4019]), .B(p_input[4003]), .Z(n2539) );
  XNOR U2144 ( .A(n2137), .B(n2534), .Z(n2536) );
  XOR U2145 ( .A(n2540), .B(n2541), .Z(n2137) );
  AND U2146 ( .A(n108), .B(n2542), .Z(n2541) );
  XOR U2147 ( .A(p_input[3987]), .B(p_input[3971]), .Z(n2542) );
  XOR U2148 ( .A(n2543), .B(n2544), .Z(n2534) );
  AND U2149 ( .A(n2545), .B(n2546), .Z(n2544) );
  XOR U2150 ( .A(n2543), .B(n2152), .Z(n2546) );
  XNOR U2151 ( .A(p_input[4002]), .B(n2547), .Z(n2152) );
  AND U2152 ( .A(n111), .B(n2548), .Z(n2547) );
  XOR U2153 ( .A(p_input[4018]), .B(p_input[4002]), .Z(n2548) );
  XNOR U2154 ( .A(n2149), .B(n2543), .Z(n2545) );
  XOR U2155 ( .A(n2549), .B(n2550), .Z(n2149) );
  AND U2156 ( .A(n108), .B(n2551), .Z(n2550) );
  XOR U2157 ( .A(p_input[3986]), .B(p_input[3970]), .Z(n2551) );
  XOR U2158 ( .A(n2552), .B(n2553), .Z(n2543) );
  AND U2159 ( .A(n2554), .B(n2555), .Z(n2553) );
  XNOR U2160 ( .A(n2556), .B(n2165), .Z(n2555) );
  XNOR U2161 ( .A(p_input[4001]), .B(n2557), .Z(n2165) );
  AND U2162 ( .A(n111), .B(n2558), .Z(n2557) );
  XNOR U2163 ( .A(p_input[4017]), .B(n2559), .Z(n2558) );
  IV U2164 ( .A(p_input[4001]), .Z(n2559) );
  XNOR U2165 ( .A(n2162), .B(n2552), .Z(n2554) );
  XNOR U2166 ( .A(p_input[3969]), .B(n2560), .Z(n2162) );
  AND U2167 ( .A(n108), .B(n2561), .Z(n2560) );
  XOR U2168 ( .A(p_input[3985]), .B(p_input[3969]), .Z(n2561) );
  IV U2169 ( .A(n2556), .Z(n2552) );
  AND U2170 ( .A(n2427), .B(n2430), .Z(n2556) );
  XOR U2171 ( .A(p_input[4000]), .B(n2562), .Z(n2430) );
  AND U2172 ( .A(n111), .B(n2563), .Z(n2562) );
  XOR U2173 ( .A(p_input[4016]), .B(p_input[4000]), .Z(n2563) );
  XOR U2174 ( .A(n2564), .B(n2565), .Z(n111) );
  AND U2175 ( .A(n2566), .B(n2567), .Z(n2565) );
  XNOR U2176 ( .A(p_input[4031]), .B(n2564), .Z(n2567) );
  XOR U2177 ( .A(n2564), .B(p_input[4015]), .Z(n2566) );
  XOR U2178 ( .A(n2568), .B(n2569), .Z(n2564) );
  AND U2179 ( .A(n2570), .B(n2571), .Z(n2569) );
  XNOR U2180 ( .A(p_input[4030]), .B(n2568), .Z(n2571) );
  XOR U2181 ( .A(n2568), .B(p_input[4014]), .Z(n2570) );
  XOR U2182 ( .A(n2572), .B(n2573), .Z(n2568) );
  AND U2183 ( .A(n2574), .B(n2575), .Z(n2573) );
  XNOR U2184 ( .A(p_input[4029]), .B(n2572), .Z(n2575) );
  XOR U2185 ( .A(n2572), .B(p_input[4013]), .Z(n2574) );
  XOR U2186 ( .A(n2576), .B(n2577), .Z(n2572) );
  AND U2187 ( .A(n2578), .B(n2579), .Z(n2577) );
  XNOR U2188 ( .A(p_input[4028]), .B(n2576), .Z(n2579) );
  XOR U2189 ( .A(n2576), .B(p_input[4012]), .Z(n2578) );
  XOR U2190 ( .A(n2580), .B(n2581), .Z(n2576) );
  AND U2191 ( .A(n2582), .B(n2583), .Z(n2581) );
  XNOR U2192 ( .A(p_input[4027]), .B(n2580), .Z(n2583) );
  XOR U2193 ( .A(n2580), .B(p_input[4011]), .Z(n2582) );
  XOR U2194 ( .A(n2584), .B(n2585), .Z(n2580) );
  AND U2195 ( .A(n2586), .B(n2587), .Z(n2585) );
  XNOR U2196 ( .A(p_input[4026]), .B(n2584), .Z(n2587) );
  XOR U2197 ( .A(n2584), .B(p_input[4010]), .Z(n2586) );
  XOR U2198 ( .A(n2588), .B(n2589), .Z(n2584) );
  AND U2199 ( .A(n2590), .B(n2591), .Z(n2589) );
  XNOR U2200 ( .A(p_input[4025]), .B(n2588), .Z(n2591) );
  XOR U2201 ( .A(n2588), .B(p_input[4009]), .Z(n2590) );
  XOR U2202 ( .A(n2592), .B(n2593), .Z(n2588) );
  AND U2203 ( .A(n2594), .B(n2595), .Z(n2593) );
  XNOR U2204 ( .A(p_input[4024]), .B(n2592), .Z(n2595) );
  XOR U2205 ( .A(n2592), .B(p_input[4008]), .Z(n2594) );
  XOR U2206 ( .A(n2596), .B(n2597), .Z(n2592) );
  AND U2207 ( .A(n2598), .B(n2599), .Z(n2597) );
  XNOR U2208 ( .A(p_input[4023]), .B(n2596), .Z(n2599) );
  XOR U2209 ( .A(n2596), .B(p_input[4007]), .Z(n2598) );
  XOR U2210 ( .A(n2600), .B(n2601), .Z(n2596) );
  AND U2211 ( .A(n2602), .B(n2603), .Z(n2601) );
  XNOR U2212 ( .A(p_input[4022]), .B(n2600), .Z(n2603) );
  XOR U2213 ( .A(n2600), .B(p_input[4006]), .Z(n2602) );
  XOR U2214 ( .A(n2604), .B(n2605), .Z(n2600) );
  AND U2215 ( .A(n2606), .B(n2607), .Z(n2605) );
  XNOR U2216 ( .A(p_input[4021]), .B(n2604), .Z(n2607) );
  XOR U2217 ( .A(n2604), .B(p_input[4005]), .Z(n2606) );
  XOR U2218 ( .A(n2608), .B(n2609), .Z(n2604) );
  AND U2219 ( .A(n2610), .B(n2611), .Z(n2609) );
  XNOR U2220 ( .A(p_input[4020]), .B(n2608), .Z(n2611) );
  XOR U2221 ( .A(n2608), .B(p_input[4004]), .Z(n2610) );
  XOR U2222 ( .A(n2612), .B(n2613), .Z(n2608) );
  AND U2223 ( .A(n2614), .B(n2615), .Z(n2613) );
  XNOR U2224 ( .A(p_input[4019]), .B(n2612), .Z(n2615) );
  XOR U2225 ( .A(n2612), .B(p_input[4003]), .Z(n2614) );
  XOR U2226 ( .A(n2616), .B(n2617), .Z(n2612) );
  AND U2227 ( .A(n2618), .B(n2619), .Z(n2617) );
  XNOR U2228 ( .A(p_input[4018]), .B(n2616), .Z(n2619) );
  XOR U2229 ( .A(n2616), .B(p_input[4002]), .Z(n2618) );
  XNOR U2230 ( .A(n2620), .B(n2621), .Z(n2616) );
  AND U2231 ( .A(n2622), .B(n2623), .Z(n2621) );
  XOR U2232 ( .A(p_input[4017]), .B(n2620), .Z(n2623) );
  XNOR U2233 ( .A(p_input[4001]), .B(n2620), .Z(n2622) );
  AND U2234 ( .A(p_input[4016]), .B(n2624), .Z(n2620) );
  IV U2235 ( .A(p_input[4000]), .Z(n2624) );
  XNOR U2236 ( .A(p_input[3968]), .B(n2625), .Z(n2427) );
  AND U2237 ( .A(n108), .B(n2626), .Z(n2625) );
  XOR U2238 ( .A(p_input[3984]), .B(p_input[3968]), .Z(n2626) );
  XOR U2239 ( .A(n2627), .B(n2628), .Z(n108) );
  AND U2240 ( .A(n2629), .B(n2630), .Z(n2628) );
  XNOR U2241 ( .A(p_input[3999]), .B(n2627), .Z(n2630) );
  XOR U2242 ( .A(n2627), .B(p_input[3983]), .Z(n2629) );
  XOR U2243 ( .A(n2631), .B(n2632), .Z(n2627) );
  AND U2244 ( .A(n2633), .B(n2634), .Z(n2632) );
  XNOR U2245 ( .A(p_input[3998]), .B(n2631), .Z(n2634) );
  XNOR U2246 ( .A(n2631), .B(n2441), .Z(n2633) );
  IV U2247 ( .A(p_input[3982]), .Z(n2441) );
  XOR U2248 ( .A(n2635), .B(n2636), .Z(n2631) );
  AND U2249 ( .A(n2637), .B(n2638), .Z(n2636) );
  XNOR U2250 ( .A(p_input[3997]), .B(n2635), .Z(n2638) );
  XNOR U2251 ( .A(n2635), .B(n2450), .Z(n2637) );
  IV U2252 ( .A(p_input[3981]), .Z(n2450) );
  XOR U2253 ( .A(n2639), .B(n2640), .Z(n2635) );
  AND U2254 ( .A(n2641), .B(n2642), .Z(n2640) );
  XNOR U2255 ( .A(p_input[3996]), .B(n2639), .Z(n2642) );
  XNOR U2256 ( .A(n2639), .B(n2459), .Z(n2641) );
  IV U2257 ( .A(p_input[3980]), .Z(n2459) );
  XOR U2258 ( .A(n2643), .B(n2644), .Z(n2639) );
  AND U2259 ( .A(n2645), .B(n2646), .Z(n2644) );
  XNOR U2260 ( .A(p_input[3995]), .B(n2643), .Z(n2646) );
  XNOR U2261 ( .A(n2643), .B(n2468), .Z(n2645) );
  IV U2262 ( .A(p_input[3979]), .Z(n2468) );
  XOR U2263 ( .A(n2647), .B(n2648), .Z(n2643) );
  AND U2264 ( .A(n2649), .B(n2650), .Z(n2648) );
  XNOR U2265 ( .A(p_input[3994]), .B(n2647), .Z(n2650) );
  XNOR U2266 ( .A(n2647), .B(n2477), .Z(n2649) );
  IV U2267 ( .A(p_input[3978]), .Z(n2477) );
  XOR U2268 ( .A(n2651), .B(n2652), .Z(n2647) );
  AND U2269 ( .A(n2653), .B(n2654), .Z(n2652) );
  XNOR U2270 ( .A(p_input[3993]), .B(n2651), .Z(n2654) );
  XNOR U2271 ( .A(n2651), .B(n2486), .Z(n2653) );
  IV U2272 ( .A(p_input[3977]), .Z(n2486) );
  XOR U2273 ( .A(n2655), .B(n2656), .Z(n2651) );
  AND U2274 ( .A(n2657), .B(n2658), .Z(n2656) );
  XNOR U2275 ( .A(p_input[3992]), .B(n2655), .Z(n2658) );
  XNOR U2276 ( .A(n2655), .B(n2495), .Z(n2657) );
  IV U2277 ( .A(p_input[3976]), .Z(n2495) );
  XOR U2278 ( .A(n2659), .B(n2660), .Z(n2655) );
  AND U2279 ( .A(n2661), .B(n2662), .Z(n2660) );
  XNOR U2280 ( .A(p_input[3991]), .B(n2659), .Z(n2662) );
  XNOR U2281 ( .A(n2659), .B(n2504), .Z(n2661) );
  IV U2282 ( .A(p_input[3975]), .Z(n2504) );
  XOR U2283 ( .A(n2663), .B(n2664), .Z(n2659) );
  AND U2284 ( .A(n2665), .B(n2666), .Z(n2664) );
  XNOR U2285 ( .A(p_input[3990]), .B(n2663), .Z(n2666) );
  XNOR U2286 ( .A(n2663), .B(n2513), .Z(n2665) );
  IV U2287 ( .A(p_input[3974]), .Z(n2513) );
  XOR U2288 ( .A(n2667), .B(n2668), .Z(n2663) );
  AND U2289 ( .A(n2669), .B(n2670), .Z(n2668) );
  XNOR U2290 ( .A(p_input[3989]), .B(n2667), .Z(n2670) );
  XNOR U2291 ( .A(n2667), .B(n2522), .Z(n2669) );
  IV U2292 ( .A(p_input[3973]), .Z(n2522) );
  XOR U2293 ( .A(n2671), .B(n2672), .Z(n2667) );
  AND U2294 ( .A(n2673), .B(n2674), .Z(n2672) );
  XNOR U2295 ( .A(p_input[3988]), .B(n2671), .Z(n2674) );
  XNOR U2296 ( .A(n2671), .B(n2531), .Z(n2673) );
  IV U2297 ( .A(p_input[3972]), .Z(n2531) );
  XOR U2298 ( .A(n2675), .B(n2676), .Z(n2671) );
  AND U2299 ( .A(n2677), .B(n2678), .Z(n2676) );
  XNOR U2300 ( .A(p_input[3987]), .B(n2675), .Z(n2678) );
  XNOR U2301 ( .A(n2675), .B(n2540), .Z(n2677) );
  IV U2302 ( .A(p_input[3971]), .Z(n2540) );
  XOR U2303 ( .A(n2679), .B(n2680), .Z(n2675) );
  AND U2304 ( .A(n2681), .B(n2682), .Z(n2680) );
  XNOR U2305 ( .A(p_input[3986]), .B(n2679), .Z(n2682) );
  XNOR U2306 ( .A(n2679), .B(n2549), .Z(n2681) );
  IV U2307 ( .A(p_input[3970]), .Z(n2549) );
  XNOR U2308 ( .A(n2683), .B(n2684), .Z(n2679) );
  AND U2309 ( .A(n2685), .B(n2686), .Z(n2684) );
  XOR U2310 ( .A(p_input[3985]), .B(n2683), .Z(n2686) );
  XNOR U2311 ( .A(p_input[3969]), .B(n2683), .Z(n2685) );
  AND U2312 ( .A(p_input[3984]), .B(n2687), .Z(n2683) );
  IV U2313 ( .A(p_input[3968]), .Z(n2687) );
  XOR U2314 ( .A(n2688), .B(n2689), .Z(n1803) );
  AND U2315 ( .A(n733), .B(n2690), .Z(n2689) );
  XNOR U2316 ( .A(n2691), .B(n2688), .Z(n2690) );
  XOR U2317 ( .A(n2692), .B(n2693), .Z(n733) );
  AND U2318 ( .A(n2694), .B(n2695), .Z(n2693) );
  XNOR U2319 ( .A(n1815), .B(n2692), .Z(n2695) );
  AND U2320 ( .A(n2696), .B(n2697), .Z(n1815) );
  XOR U2321 ( .A(n2692), .B(n1814), .Z(n2694) );
  AND U2322 ( .A(n2698), .B(n2699), .Z(n1814) );
  XOR U2323 ( .A(n2700), .B(n2701), .Z(n2692) );
  AND U2324 ( .A(n2702), .B(n2703), .Z(n2701) );
  XOR U2325 ( .A(n2700), .B(n1827), .Z(n2703) );
  XOR U2326 ( .A(n2704), .B(n2705), .Z(n1827) );
  AND U2327 ( .A(n363), .B(n2706), .Z(n2705) );
  XOR U2328 ( .A(n2707), .B(n2704), .Z(n2706) );
  XNOR U2329 ( .A(n1824), .B(n2700), .Z(n2702) );
  XOR U2330 ( .A(n2708), .B(n2709), .Z(n1824) );
  AND U2331 ( .A(n360), .B(n2710), .Z(n2709) );
  XOR U2332 ( .A(n2711), .B(n2708), .Z(n2710) );
  XOR U2333 ( .A(n2712), .B(n2713), .Z(n2700) );
  AND U2334 ( .A(n2714), .B(n2715), .Z(n2713) );
  XOR U2335 ( .A(n2712), .B(n1839), .Z(n2715) );
  XOR U2336 ( .A(n2716), .B(n2717), .Z(n1839) );
  AND U2337 ( .A(n363), .B(n2718), .Z(n2717) );
  XOR U2338 ( .A(n2719), .B(n2716), .Z(n2718) );
  XNOR U2339 ( .A(n1836), .B(n2712), .Z(n2714) );
  XOR U2340 ( .A(n2720), .B(n2721), .Z(n1836) );
  AND U2341 ( .A(n360), .B(n2722), .Z(n2721) );
  XOR U2342 ( .A(n2723), .B(n2720), .Z(n2722) );
  XOR U2343 ( .A(n2724), .B(n2725), .Z(n2712) );
  AND U2344 ( .A(n2726), .B(n2727), .Z(n2725) );
  XOR U2345 ( .A(n2724), .B(n1851), .Z(n2727) );
  XOR U2346 ( .A(n2728), .B(n2729), .Z(n1851) );
  AND U2347 ( .A(n363), .B(n2730), .Z(n2729) );
  XOR U2348 ( .A(n2731), .B(n2728), .Z(n2730) );
  XNOR U2349 ( .A(n1848), .B(n2724), .Z(n2726) );
  XOR U2350 ( .A(n2732), .B(n2733), .Z(n1848) );
  AND U2351 ( .A(n360), .B(n2734), .Z(n2733) );
  XOR U2352 ( .A(n2735), .B(n2732), .Z(n2734) );
  XOR U2353 ( .A(n2736), .B(n2737), .Z(n2724) );
  AND U2354 ( .A(n2738), .B(n2739), .Z(n2737) );
  XOR U2355 ( .A(n2736), .B(n1863), .Z(n2739) );
  XOR U2356 ( .A(n2740), .B(n2741), .Z(n1863) );
  AND U2357 ( .A(n363), .B(n2742), .Z(n2741) );
  XOR U2358 ( .A(n2743), .B(n2740), .Z(n2742) );
  XNOR U2359 ( .A(n1860), .B(n2736), .Z(n2738) );
  XOR U2360 ( .A(n2744), .B(n2745), .Z(n1860) );
  AND U2361 ( .A(n360), .B(n2746), .Z(n2745) );
  XOR U2362 ( .A(n2747), .B(n2744), .Z(n2746) );
  XOR U2363 ( .A(n2748), .B(n2749), .Z(n2736) );
  AND U2364 ( .A(n2750), .B(n2751), .Z(n2749) );
  XOR U2365 ( .A(n2748), .B(n1875), .Z(n2751) );
  XOR U2366 ( .A(n2752), .B(n2753), .Z(n1875) );
  AND U2367 ( .A(n363), .B(n2754), .Z(n2753) );
  XOR U2368 ( .A(n2755), .B(n2752), .Z(n2754) );
  XNOR U2369 ( .A(n1872), .B(n2748), .Z(n2750) );
  XOR U2370 ( .A(n2756), .B(n2757), .Z(n1872) );
  AND U2371 ( .A(n360), .B(n2758), .Z(n2757) );
  XOR U2372 ( .A(n2759), .B(n2756), .Z(n2758) );
  XOR U2373 ( .A(n2760), .B(n2761), .Z(n2748) );
  AND U2374 ( .A(n2762), .B(n2763), .Z(n2761) );
  XOR U2375 ( .A(n2760), .B(n1887), .Z(n2763) );
  XOR U2376 ( .A(n2764), .B(n2765), .Z(n1887) );
  AND U2377 ( .A(n363), .B(n2766), .Z(n2765) );
  XOR U2378 ( .A(n2767), .B(n2764), .Z(n2766) );
  XNOR U2379 ( .A(n1884), .B(n2760), .Z(n2762) );
  XOR U2380 ( .A(n2768), .B(n2769), .Z(n1884) );
  AND U2381 ( .A(n360), .B(n2770), .Z(n2769) );
  XOR U2382 ( .A(n2771), .B(n2768), .Z(n2770) );
  XOR U2383 ( .A(n2772), .B(n2773), .Z(n2760) );
  AND U2384 ( .A(n2774), .B(n2775), .Z(n2773) );
  XOR U2385 ( .A(n2772), .B(n1899), .Z(n2775) );
  XOR U2386 ( .A(n2776), .B(n2777), .Z(n1899) );
  AND U2387 ( .A(n363), .B(n2778), .Z(n2777) );
  XOR U2388 ( .A(n2779), .B(n2776), .Z(n2778) );
  XNOR U2389 ( .A(n1896), .B(n2772), .Z(n2774) );
  XOR U2390 ( .A(n2780), .B(n2781), .Z(n1896) );
  AND U2391 ( .A(n360), .B(n2782), .Z(n2781) );
  XOR U2392 ( .A(n2783), .B(n2780), .Z(n2782) );
  XOR U2393 ( .A(n2784), .B(n2785), .Z(n2772) );
  AND U2394 ( .A(n2786), .B(n2787), .Z(n2785) );
  XOR U2395 ( .A(n2784), .B(n1911), .Z(n2787) );
  XOR U2396 ( .A(n2788), .B(n2789), .Z(n1911) );
  AND U2397 ( .A(n363), .B(n2790), .Z(n2789) );
  XOR U2398 ( .A(n2791), .B(n2788), .Z(n2790) );
  XNOR U2399 ( .A(n1908), .B(n2784), .Z(n2786) );
  XOR U2400 ( .A(n2792), .B(n2793), .Z(n1908) );
  AND U2401 ( .A(n360), .B(n2794), .Z(n2793) );
  XOR U2402 ( .A(n2795), .B(n2792), .Z(n2794) );
  XOR U2403 ( .A(n2796), .B(n2797), .Z(n2784) );
  AND U2404 ( .A(n2798), .B(n2799), .Z(n2797) );
  XOR U2405 ( .A(n2796), .B(n1923), .Z(n2799) );
  XOR U2406 ( .A(n2800), .B(n2801), .Z(n1923) );
  AND U2407 ( .A(n363), .B(n2802), .Z(n2801) );
  XOR U2408 ( .A(n2803), .B(n2800), .Z(n2802) );
  XNOR U2409 ( .A(n1920), .B(n2796), .Z(n2798) );
  XOR U2410 ( .A(n2804), .B(n2805), .Z(n1920) );
  AND U2411 ( .A(n360), .B(n2806), .Z(n2805) );
  XOR U2412 ( .A(n2807), .B(n2804), .Z(n2806) );
  XOR U2413 ( .A(n2808), .B(n2809), .Z(n2796) );
  AND U2414 ( .A(n2810), .B(n2811), .Z(n2809) );
  XOR U2415 ( .A(n2808), .B(n1935), .Z(n2811) );
  XOR U2416 ( .A(n2812), .B(n2813), .Z(n1935) );
  AND U2417 ( .A(n363), .B(n2814), .Z(n2813) );
  XOR U2418 ( .A(n2815), .B(n2812), .Z(n2814) );
  XNOR U2419 ( .A(n1932), .B(n2808), .Z(n2810) );
  XOR U2420 ( .A(n2816), .B(n2817), .Z(n1932) );
  AND U2421 ( .A(n360), .B(n2818), .Z(n2817) );
  XOR U2422 ( .A(n2819), .B(n2816), .Z(n2818) );
  XOR U2423 ( .A(n2820), .B(n2821), .Z(n2808) );
  AND U2424 ( .A(n2822), .B(n2823), .Z(n2821) );
  XOR U2425 ( .A(n2820), .B(n1947), .Z(n2823) );
  XOR U2426 ( .A(n2824), .B(n2825), .Z(n1947) );
  AND U2427 ( .A(n363), .B(n2826), .Z(n2825) );
  XOR U2428 ( .A(n2827), .B(n2824), .Z(n2826) );
  XNOR U2429 ( .A(n1944), .B(n2820), .Z(n2822) );
  XOR U2430 ( .A(n2828), .B(n2829), .Z(n1944) );
  AND U2431 ( .A(n360), .B(n2830), .Z(n2829) );
  XOR U2432 ( .A(n2831), .B(n2828), .Z(n2830) );
  XOR U2433 ( .A(n2832), .B(n2833), .Z(n2820) );
  AND U2434 ( .A(n2834), .B(n2835), .Z(n2833) );
  XOR U2435 ( .A(n2832), .B(n1959), .Z(n2835) );
  XOR U2436 ( .A(n2836), .B(n2837), .Z(n1959) );
  AND U2437 ( .A(n363), .B(n2838), .Z(n2837) );
  XOR U2438 ( .A(n2839), .B(n2836), .Z(n2838) );
  XNOR U2439 ( .A(n1956), .B(n2832), .Z(n2834) );
  XOR U2440 ( .A(n2840), .B(n2841), .Z(n1956) );
  AND U2441 ( .A(n360), .B(n2842), .Z(n2841) );
  XOR U2442 ( .A(n2843), .B(n2840), .Z(n2842) );
  XOR U2443 ( .A(n2844), .B(n2845), .Z(n2832) );
  AND U2444 ( .A(n2846), .B(n2847), .Z(n2845) );
  XOR U2445 ( .A(n2844), .B(n1971), .Z(n2847) );
  XOR U2446 ( .A(n2848), .B(n2849), .Z(n1971) );
  AND U2447 ( .A(n363), .B(n2850), .Z(n2849) );
  XOR U2448 ( .A(n2851), .B(n2848), .Z(n2850) );
  XNOR U2449 ( .A(n1968), .B(n2844), .Z(n2846) );
  XOR U2450 ( .A(n2852), .B(n2853), .Z(n1968) );
  AND U2451 ( .A(n360), .B(n2854), .Z(n2853) );
  XOR U2452 ( .A(n2855), .B(n2852), .Z(n2854) );
  XOR U2453 ( .A(n2856), .B(n2857), .Z(n2844) );
  AND U2454 ( .A(n2858), .B(n2859), .Z(n2857) );
  XNOR U2455 ( .A(n2860), .B(n1984), .Z(n2859) );
  XOR U2456 ( .A(n2861), .B(n2862), .Z(n1984) );
  AND U2457 ( .A(n363), .B(n2863), .Z(n2862) );
  XOR U2458 ( .A(n2861), .B(n2864), .Z(n2863) );
  XNOR U2459 ( .A(n1981), .B(n2856), .Z(n2858) );
  XOR U2460 ( .A(n2865), .B(n2866), .Z(n1981) );
  AND U2461 ( .A(n360), .B(n2867), .Z(n2866) );
  XOR U2462 ( .A(n2865), .B(n2868), .Z(n2867) );
  IV U2463 ( .A(n2860), .Z(n2856) );
  AND U2464 ( .A(n2688), .B(n2691), .Z(n2860) );
  XNOR U2465 ( .A(n2869), .B(n2870), .Z(n2691) );
  AND U2466 ( .A(n363), .B(n2871), .Z(n2870) );
  XNOR U2467 ( .A(n2872), .B(n2869), .Z(n2871) );
  XOR U2468 ( .A(n2873), .B(n2874), .Z(n363) );
  AND U2469 ( .A(n2875), .B(n2876), .Z(n2874) );
  XNOR U2470 ( .A(n2696), .B(n2873), .Z(n2876) );
  AND U2471 ( .A(p_input[3967]), .B(p_input[3951]), .Z(n2696) );
  XOR U2472 ( .A(n2873), .B(n2697), .Z(n2875) );
  AND U2473 ( .A(p_input[3935]), .B(p_input[3919]), .Z(n2697) );
  XOR U2474 ( .A(n2877), .B(n2878), .Z(n2873) );
  AND U2475 ( .A(n2879), .B(n2880), .Z(n2878) );
  XOR U2476 ( .A(n2877), .B(n2707), .Z(n2880) );
  XNOR U2477 ( .A(p_input[3950]), .B(n2881), .Z(n2707) );
  AND U2478 ( .A(n119), .B(n2882), .Z(n2881) );
  XOR U2479 ( .A(p_input[3966]), .B(p_input[3950]), .Z(n2882) );
  XNOR U2480 ( .A(n2704), .B(n2877), .Z(n2879) );
  XOR U2481 ( .A(n2883), .B(n2884), .Z(n2704) );
  AND U2482 ( .A(n117), .B(n2885), .Z(n2884) );
  XOR U2483 ( .A(p_input[3934]), .B(p_input[3918]), .Z(n2885) );
  XOR U2484 ( .A(n2886), .B(n2887), .Z(n2877) );
  AND U2485 ( .A(n2888), .B(n2889), .Z(n2887) );
  XOR U2486 ( .A(n2886), .B(n2719), .Z(n2889) );
  XNOR U2487 ( .A(p_input[3949]), .B(n2890), .Z(n2719) );
  AND U2488 ( .A(n119), .B(n2891), .Z(n2890) );
  XOR U2489 ( .A(p_input[3965]), .B(p_input[3949]), .Z(n2891) );
  XNOR U2490 ( .A(n2716), .B(n2886), .Z(n2888) );
  XOR U2491 ( .A(n2892), .B(n2893), .Z(n2716) );
  AND U2492 ( .A(n117), .B(n2894), .Z(n2893) );
  XOR U2493 ( .A(p_input[3933]), .B(p_input[3917]), .Z(n2894) );
  XOR U2494 ( .A(n2895), .B(n2896), .Z(n2886) );
  AND U2495 ( .A(n2897), .B(n2898), .Z(n2896) );
  XOR U2496 ( .A(n2895), .B(n2731), .Z(n2898) );
  XNOR U2497 ( .A(p_input[3948]), .B(n2899), .Z(n2731) );
  AND U2498 ( .A(n119), .B(n2900), .Z(n2899) );
  XOR U2499 ( .A(p_input[3964]), .B(p_input[3948]), .Z(n2900) );
  XNOR U2500 ( .A(n2728), .B(n2895), .Z(n2897) );
  XOR U2501 ( .A(n2901), .B(n2902), .Z(n2728) );
  AND U2502 ( .A(n117), .B(n2903), .Z(n2902) );
  XOR U2503 ( .A(p_input[3932]), .B(p_input[3916]), .Z(n2903) );
  XOR U2504 ( .A(n2904), .B(n2905), .Z(n2895) );
  AND U2505 ( .A(n2906), .B(n2907), .Z(n2905) );
  XOR U2506 ( .A(n2904), .B(n2743), .Z(n2907) );
  XNOR U2507 ( .A(p_input[3947]), .B(n2908), .Z(n2743) );
  AND U2508 ( .A(n119), .B(n2909), .Z(n2908) );
  XOR U2509 ( .A(p_input[3963]), .B(p_input[3947]), .Z(n2909) );
  XNOR U2510 ( .A(n2740), .B(n2904), .Z(n2906) );
  XOR U2511 ( .A(n2910), .B(n2911), .Z(n2740) );
  AND U2512 ( .A(n117), .B(n2912), .Z(n2911) );
  XOR U2513 ( .A(p_input[3931]), .B(p_input[3915]), .Z(n2912) );
  XOR U2514 ( .A(n2913), .B(n2914), .Z(n2904) );
  AND U2515 ( .A(n2915), .B(n2916), .Z(n2914) );
  XOR U2516 ( .A(n2913), .B(n2755), .Z(n2916) );
  XNOR U2517 ( .A(p_input[3946]), .B(n2917), .Z(n2755) );
  AND U2518 ( .A(n119), .B(n2918), .Z(n2917) );
  XOR U2519 ( .A(p_input[3962]), .B(p_input[3946]), .Z(n2918) );
  XNOR U2520 ( .A(n2752), .B(n2913), .Z(n2915) );
  XOR U2521 ( .A(n2919), .B(n2920), .Z(n2752) );
  AND U2522 ( .A(n117), .B(n2921), .Z(n2920) );
  XOR U2523 ( .A(p_input[3930]), .B(p_input[3914]), .Z(n2921) );
  XOR U2524 ( .A(n2922), .B(n2923), .Z(n2913) );
  AND U2525 ( .A(n2924), .B(n2925), .Z(n2923) );
  XOR U2526 ( .A(n2922), .B(n2767), .Z(n2925) );
  XNOR U2527 ( .A(p_input[3945]), .B(n2926), .Z(n2767) );
  AND U2528 ( .A(n119), .B(n2927), .Z(n2926) );
  XOR U2529 ( .A(p_input[3961]), .B(p_input[3945]), .Z(n2927) );
  XNOR U2530 ( .A(n2764), .B(n2922), .Z(n2924) );
  XOR U2531 ( .A(n2928), .B(n2929), .Z(n2764) );
  AND U2532 ( .A(n117), .B(n2930), .Z(n2929) );
  XOR U2533 ( .A(p_input[3929]), .B(p_input[3913]), .Z(n2930) );
  XOR U2534 ( .A(n2931), .B(n2932), .Z(n2922) );
  AND U2535 ( .A(n2933), .B(n2934), .Z(n2932) );
  XOR U2536 ( .A(n2931), .B(n2779), .Z(n2934) );
  XNOR U2537 ( .A(p_input[3944]), .B(n2935), .Z(n2779) );
  AND U2538 ( .A(n119), .B(n2936), .Z(n2935) );
  XOR U2539 ( .A(p_input[3960]), .B(p_input[3944]), .Z(n2936) );
  XNOR U2540 ( .A(n2776), .B(n2931), .Z(n2933) );
  XOR U2541 ( .A(n2937), .B(n2938), .Z(n2776) );
  AND U2542 ( .A(n117), .B(n2939), .Z(n2938) );
  XOR U2543 ( .A(p_input[3928]), .B(p_input[3912]), .Z(n2939) );
  XOR U2544 ( .A(n2940), .B(n2941), .Z(n2931) );
  AND U2545 ( .A(n2942), .B(n2943), .Z(n2941) );
  XOR U2546 ( .A(n2940), .B(n2791), .Z(n2943) );
  XNOR U2547 ( .A(p_input[3943]), .B(n2944), .Z(n2791) );
  AND U2548 ( .A(n119), .B(n2945), .Z(n2944) );
  XOR U2549 ( .A(p_input[3959]), .B(p_input[3943]), .Z(n2945) );
  XNOR U2550 ( .A(n2788), .B(n2940), .Z(n2942) );
  XOR U2551 ( .A(n2946), .B(n2947), .Z(n2788) );
  AND U2552 ( .A(n117), .B(n2948), .Z(n2947) );
  XOR U2553 ( .A(p_input[3927]), .B(p_input[3911]), .Z(n2948) );
  XOR U2554 ( .A(n2949), .B(n2950), .Z(n2940) );
  AND U2555 ( .A(n2951), .B(n2952), .Z(n2950) );
  XOR U2556 ( .A(n2949), .B(n2803), .Z(n2952) );
  XNOR U2557 ( .A(p_input[3942]), .B(n2953), .Z(n2803) );
  AND U2558 ( .A(n119), .B(n2954), .Z(n2953) );
  XOR U2559 ( .A(p_input[3958]), .B(p_input[3942]), .Z(n2954) );
  XNOR U2560 ( .A(n2800), .B(n2949), .Z(n2951) );
  XOR U2561 ( .A(n2955), .B(n2956), .Z(n2800) );
  AND U2562 ( .A(n117), .B(n2957), .Z(n2956) );
  XOR U2563 ( .A(p_input[3926]), .B(p_input[3910]), .Z(n2957) );
  XOR U2564 ( .A(n2958), .B(n2959), .Z(n2949) );
  AND U2565 ( .A(n2960), .B(n2961), .Z(n2959) );
  XOR U2566 ( .A(n2958), .B(n2815), .Z(n2961) );
  XNOR U2567 ( .A(p_input[3941]), .B(n2962), .Z(n2815) );
  AND U2568 ( .A(n119), .B(n2963), .Z(n2962) );
  XOR U2569 ( .A(p_input[3957]), .B(p_input[3941]), .Z(n2963) );
  XNOR U2570 ( .A(n2812), .B(n2958), .Z(n2960) );
  XOR U2571 ( .A(n2964), .B(n2965), .Z(n2812) );
  AND U2572 ( .A(n117), .B(n2966), .Z(n2965) );
  XOR U2573 ( .A(p_input[3925]), .B(p_input[3909]), .Z(n2966) );
  XOR U2574 ( .A(n2967), .B(n2968), .Z(n2958) );
  AND U2575 ( .A(n2969), .B(n2970), .Z(n2968) );
  XOR U2576 ( .A(n2967), .B(n2827), .Z(n2970) );
  XNOR U2577 ( .A(p_input[3940]), .B(n2971), .Z(n2827) );
  AND U2578 ( .A(n119), .B(n2972), .Z(n2971) );
  XOR U2579 ( .A(p_input[3956]), .B(p_input[3940]), .Z(n2972) );
  XNOR U2580 ( .A(n2824), .B(n2967), .Z(n2969) );
  XOR U2581 ( .A(n2973), .B(n2974), .Z(n2824) );
  AND U2582 ( .A(n117), .B(n2975), .Z(n2974) );
  XOR U2583 ( .A(p_input[3924]), .B(p_input[3908]), .Z(n2975) );
  XOR U2584 ( .A(n2976), .B(n2977), .Z(n2967) );
  AND U2585 ( .A(n2978), .B(n2979), .Z(n2977) );
  XOR U2586 ( .A(n2976), .B(n2839), .Z(n2979) );
  XNOR U2587 ( .A(p_input[3939]), .B(n2980), .Z(n2839) );
  AND U2588 ( .A(n119), .B(n2981), .Z(n2980) );
  XOR U2589 ( .A(p_input[3955]), .B(p_input[3939]), .Z(n2981) );
  XNOR U2590 ( .A(n2836), .B(n2976), .Z(n2978) );
  XOR U2591 ( .A(n2982), .B(n2983), .Z(n2836) );
  AND U2592 ( .A(n117), .B(n2984), .Z(n2983) );
  XOR U2593 ( .A(p_input[3923]), .B(p_input[3907]), .Z(n2984) );
  XOR U2594 ( .A(n2985), .B(n2986), .Z(n2976) );
  AND U2595 ( .A(n2987), .B(n2988), .Z(n2986) );
  XOR U2596 ( .A(n2985), .B(n2851), .Z(n2988) );
  XNOR U2597 ( .A(p_input[3938]), .B(n2989), .Z(n2851) );
  AND U2598 ( .A(n119), .B(n2990), .Z(n2989) );
  XOR U2599 ( .A(p_input[3954]), .B(p_input[3938]), .Z(n2990) );
  XNOR U2600 ( .A(n2848), .B(n2985), .Z(n2987) );
  XOR U2601 ( .A(n2991), .B(n2992), .Z(n2848) );
  AND U2602 ( .A(n117), .B(n2993), .Z(n2992) );
  XOR U2603 ( .A(p_input[3922]), .B(p_input[3906]), .Z(n2993) );
  XOR U2604 ( .A(n2994), .B(n2995), .Z(n2985) );
  AND U2605 ( .A(n2996), .B(n2997), .Z(n2995) );
  XNOR U2606 ( .A(n2998), .B(n2864), .Z(n2997) );
  XNOR U2607 ( .A(p_input[3937]), .B(n2999), .Z(n2864) );
  AND U2608 ( .A(n119), .B(n3000), .Z(n2999) );
  XNOR U2609 ( .A(p_input[3953]), .B(n3001), .Z(n3000) );
  IV U2610 ( .A(p_input[3937]), .Z(n3001) );
  XNOR U2611 ( .A(n2861), .B(n2994), .Z(n2996) );
  XNOR U2612 ( .A(p_input[3905]), .B(n3002), .Z(n2861) );
  AND U2613 ( .A(n117), .B(n3003), .Z(n3002) );
  XOR U2614 ( .A(p_input[3921]), .B(p_input[3905]), .Z(n3003) );
  IV U2615 ( .A(n2998), .Z(n2994) );
  AND U2616 ( .A(n2869), .B(n2872), .Z(n2998) );
  XOR U2617 ( .A(p_input[3936]), .B(n3004), .Z(n2872) );
  AND U2618 ( .A(n119), .B(n3005), .Z(n3004) );
  XOR U2619 ( .A(p_input[3952]), .B(p_input[3936]), .Z(n3005) );
  XOR U2620 ( .A(n3006), .B(n3007), .Z(n119) );
  AND U2621 ( .A(n3008), .B(n3009), .Z(n3007) );
  XNOR U2622 ( .A(p_input[3967]), .B(n3006), .Z(n3009) );
  XOR U2623 ( .A(n3006), .B(p_input[3951]), .Z(n3008) );
  XOR U2624 ( .A(n3010), .B(n3011), .Z(n3006) );
  AND U2625 ( .A(n3012), .B(n3013), .Z(n3011) );
  XNOR U2626 ( .A(p_input[3966]), .B(n3010), .Z(n3013) );
  XOR U2627 ( .A(n3010), .B(p_input[3950]), .Z(n3012) );
  XOR U2628 ( .A(n3014), .B(n3015), .Z(n3010) );
  AND U2629 ( .A(n3016), .B(n3017), .Z(n3015) );
  XNOR U2630 ( .A(p_input[3965]), .B(n3014), .Z(n3017) );
  XOR U2631 ( .A(n3014), .B(p_input[3949]), .Z(n3016) );
  XOR U2632 ( .A(n3018), .B(n3019), .Z(n3014) );
  AND U2633 ( .A(n3020), .B(n3021), .Z(n3019) );
  XNOR U2634 ( .A(p_input[3964]), .B(n3018), .Z(n3021) );
  XOR U2635 ( .A(n3018), .B(p_input[3948]), .Z(n3020) );
  XOR U2636 ( .A(n3022), .B(n3023), .Z(n3018) );
  AND U2637 ( .A(n3024), .B(n3025), .Z(n3023) );
  XNOR U2638 ( .A(p_input[3963]), .B(n3022), .Z(n3025) );
  XOR U2639 ( .A(n3022), .B(p_input[3947]), .Z(n3024) );
  XOR U2640 ( .A(n3026), .B(n3027), .Z(n3022) );
  AND U2641 ( .A(n3028), .B(n3029), .Z(n3027) );
  XNOR U2642 ( .A(p_input[3962]), .B(n3026), .Z(n3029) );
  XOR U2643 ( .A(n3026), .B(p_input[3946]), .Z(n3028) );
  XOR U2644 ( .A(n3030), .B(n3031), .Z(n3026) );
  AND U2645 ( .A(n3032), .B(n3033), .Z(n3031) );
  XNOR U2646 ( .A(p_input[3961]), .B(n3030), .Z(n3033) );
  XOR U2647 ( .A(n3030), .B(p_input[3945]), .Z(n3032) );
  XOR U2648 ( .A(n3034), .B(n3035), .Z(n3030) );
  AND U2649 ( .A(n3036), .B(n3037), .Z(n3035) );
  XNOR U2650 ( .A(p_input[3960]), .B(n3034), .Z(n3037) );
  XOR U2651 ( .A(n3034), .B(p_input[3944]), .Z(n3036) );
  XOR U2652 ( .A(n3038), .B(n3039), .Z(n3034) );
  AND U2653 ( .A(n3040), .B(n3041), .Z(n3039) );
  XNOR U2654 ( .A(p_input[3959]), .B(n3038), .Z(n3041) );
  XOR U2655 ( .A(n3038), .B(p_input[3943]), .Z(n3040) );
  XOR U2656 ( .A(n3042), .B(n3043), .Z(n3038) );
  AND U2657 ( .A(n3044), .B(n3045), .Z(n3043) );
  XNOR U2658 ( .A(p_input[3958]), .B(n3042), .Z(n3045) );
  XOR U2659 ( .A(n3042), .B(p_input[3942]), .Z(n3044) );
  XOR U2660 ( .A(n3046), .B(n3047), .Z(n3042) );
  AND U2661 ( .A(n3048), .B(n3049), .Z(n3047) );
  XNOR U2662 ( .A(p_input[3957]), .B(n3046), .Z(n3049) );
  XOR U2663 ( .A(n3046), .B(p_input[3941]), .Z(n3048) );
  XOR U2664 ( .A(n3050), .B(n3051), .Z(n3046) );
  AND U2665 ( .A(n3052), .B(n3053), .Z(n3051) );
  XNOR U2666 ( .A(p_input[3956]), .B(n3050), .Z(n3053) );
  XOR U2667 ( .A(n3050), .B(p_input[3940]), .Z(n3052) );
  XOR U2668 ( .A(n3054), .B(n3055), .Z(n3050) );
  AND U2669 ( .A(n3056), .B(n3057), .Z(n3055) );
  XNOR U2670 ( .A(p_input[3955]), .B(n3054), .Z(n3057) );
  XOR U2671 ( .A(n3054), .B(p_input[3939]), .Z(n3056) );
  XOR U2672 ( .A(n3058), .B(n3059), .Z(n3054) );
  AND U2673 ( .A(n3060), .B(n3061), .Z(n3059) );
  XNOR U2674 ( .A(p_input[3954]), .B(n3058), .Z(n3061) );
  XOR U2675 ( .A(n3058), .B(p_input[3938]), .Z(n3060) );
  XNOR U2676 ( .A(n3062), .B(n3063), .Z(n3058) );
  AND U2677 ( .A(n3064), .B(n3065), .Z(n3063) );
  XOR U2678 ( .A(p_input[3953]), .B(n3062), .Z(n3065) );
  XNOR U2679 ( .A(p_input[3937]), .B(n3062), .Z(n3064) );
  AND U2680 ( .A(p_input[3952]), .B(n3066), .Z(n3062) );
  IV U2681 ( .A(p_input[3936]), .Z(n3066) );
  XNOR U2682 ( .A(p_input[3904]), .B(n3067), .Z(n2869) );
  AND U2683 ( .A(n117), .B(n3068), .Z(n3067) );
  XOR U2684 ( .A(p_input[3920]), .B(p_input[3904]), .Z(n3068) );
  XOR U2685 ( .A(n3069), .B(n3070), .Z(n117) );
  AND U2686 ( .A(n3071), .B(n3072), .Z(n3070) );
  XNOR U2687 ( .A(p_input[3935]), .B(n3069), .Z(n3072) );
  XOR U2688 ( .A(n3069), .B(p_input[3919]), .Z(n3071) );
  XOR U2689 ( .A(n3073), .B(n3074), .Z(n3069) );
  AND U2690 ( .A(n3075), .B(n3076), .Z(n3074) );
  XNOR U2691 ( .A(p_input[3934]), .B(n3073), .Z(n3076) );
  XNOR U2692 ( .A(n3073), .B(n2883), .Z(n3075) );
  IV U2693 ( .A(p_input[3918]), .Z(n2883) );
  XOR U2694 ( .A(n3077), .B(n3078), .Z(n3073) );
  AND U2695 ( .A(n3079), .B(n3080), .Z(n3078) );
  XNOR U2696 ( .A(p_input[3933]), .B(n3077), .Z(n3080) );
  XNOR U2697 ( .A(n3077), .B(n2892), .Z(n3079) );
  IV U2698 ( .A(p_input[3917]), .Z(n2892) );
  XOR U2699 ( .A(n3081), .B(n3082), .Z(n3077) );
  AND U2700 ( .A(n3083), .B(n3084), .Z(n3082) );
  XNOR U2701 ( .A(p_input[3932]), .B(n3081), .Z(n3084) );
  XNOR U2702 ( .A(n3081), .B(n2901), .Z(n3083) );
  IV U2703 ( .A(p_input[3916]), .Z(n2901) );
  XOR U2704 ( .A(n3085), .B(n3086), .Z(n3081) );
  AND U2705 ( .A(n3087), .B(n3088), .Z(n3086) );
  XNOR U2706 ( .A(p_input[3931]), .B(n3085), .Z(n3088) );
  XNOR U2707 ( .A(n3085), .B(n2910), .Z(n3087) );
  IV U2708 ( .A(p_input[3915]), .Z(n2910) );
  XOR U2709 ( .A(n3089), .B(n3090), .Z(n3085) );
  AND U2710 ( .A(n3091), .B(n3092), .Z(n3090) );
  XNOR U2711 ( .A(p_input[3930]), .B(n3089), .Z(n3092) );
  XNOR U2712 ( .A(n3089), .B(n2919), .Z(n3091) );
  IV U2713 ( .A(p_input[3914]), .Z(n2919) );
  XOR U2714 ( .A(n3093), .B(n3094), .Z(n3089) );
  AND U2715 ( .A(n3095), .B(n3096), .Z(n3094) );
  XNOR U2716 ( .A(p_input[3929]), .B(n3093), .Z(n3096) );
  XNOR U2717 ( .A(n3093), .B(n2928), .Z(n3095) );
  IV U2718 ( .A(p_input[3913]), .Z(n2928) );
  XOR U2719 ( .A(n3097), .B(n3098), .Z(n3093) );
  AND U2720 ( .A(n3099), .B(n3100), .Z(n3098) );
  XNOR U2721 ( .A(p_input[3928]), .B(n3097), .Z(n3100) );
  XNOR U2722 ( .A(n3097), .B(n2937), .Z(n3099) );
  IV U2723 ( .A(p_input[3912]), .Z(n2937) );
  XOR U2724 ( .A(n3101), .B(n3102), .Z(n3097) );
  AND U2725 ( .A(n3103), .B(n3104), .Z(n3102) );
  XNOR U2726 ( .A(p_input[3927]), .B(n3101), .Z(n3104) );
  XNOR U2727 ( .A(n3101), .B(n2946), .Z(n3103) );
  IV U2728 ( .A(p_input[3911]), .Z(n2946) );
  XOR U2729 ( .A(n3105), .B(n3106), .Z(n3101) );
  AND U2730 ( .A(n3107), .B(n3108), .Z(n3106) );
  XNOR U2731 ( .A(p_input[3926]), .B(n3105), .Z(n3108) );
  XNOR U2732 ( .A(n3105), .B(n2955), .Z(n3107) );
  IV U2733 ( .A(p_input[3910]), .Z(n2955) );
  XOR U2734 ( .A(n3109), .B(n3110), .Z(n3105) );
  AND U2735 ( .A(n3111), .B(n3112), .Z(n3110) );
  XNOR U2736 ( .A(p_input[3925]), .B(n3109), .Z(n3112) );
  XNOR U2737 ( .A(n3109), .B(n2964), .Z(n3111) );
  IV U2738 ( .A(p_input[3909]), .Z(n2964) );
  XOR U2739 ( .A(n3113), .B(n3114), .Z(n3109) );
  AND U2740 ( .A(n3115), .B(n3116), .Z(n3114) );
  XNOR U2741 ( .A(p_input[3924]), .B(n3113), .Z(n3116) );
  XNOR U2742 ( .A(n3113), .B(n2973), .Z(n3115) );
  IV U2743 ( .A(p_input[3908]), .Z(n2973) );
  XOR U2744 ( .A(n3117), .B(n3118), .Z(n3113) );
  AND U2745 ( .A(n3119), .B(n3120), .Z(n3118) );
  XNOR U2746 ( .A(p_input[3923]), .B(n3117), .Z(n3120) );
  XNOR U2747 ( .A(n3117), .B(n2982), .Z(n3119) );
  IV U2748 ( .A(p_input[3907]), .Z(n2982) );
  XOR U2749 ( .A(n3121), .B(n3122), .Z(n3117) );
  AND U2750 ( .A(n3123), .B(n3124), .Z(n3122) );
  XNOR U2751 ( .A(p_input[3922]), .B(n3121), .Z(n3124) );
  XNOR U2752 ( .A(n3121), .B(n2991), .Z(n3123) );
  IV U2753 ( .A(p_input[3906]), .Z(n2991) );
  XNOR U2754 ( .A(n3125), .B(n3126), .Z(n3121) );
  AND U2755 ( .A(n3127), .B(n3128), .Z(n3126) );
  XOR U2756 ( .A(p_input[3921]), .B(n3125), .Z(n3128) );
  XNOR U2757 ( .A(p_input[3905]), .B(n3125), .Z(n3127) );
  AND U2758 ( .A(p_input[3920]), .B(n3129), .Z(n3125) );
  IV U2759 ( .A(p_input[3904]), .Z(n3129) );
  XOR U2760 ( .A(n3130), .B(n3131), .Z(n2688) );
  AND U2761 ( .A(n360), .B(n3132), .Z(n3131) );
  XNOR U2762 ( .A(n3133), .B(n3130), .Z(n3132) );
  XOR U2763 ( .A(n3134), .B(n3135), .Z(n360) );
  AND U2764 ( .A(n3136), .B(n3137), .Z(n3135) );
  XNOR U2765 ( .A(n2699), .B(n3134), .Z(n3137) );
  AND U2766 ( .A(p_input[3903]), .B(p_input[3887]), .Z(n2699) );
  XOR U2767 ( .A(n3134), .B(n2698), .Z(n3136) );
  AND U2768 ( .A(p_input[3855]), .B(p_input[3871]), .Z(n2698) );
  XOR U2769 ( .A(n3138), .B(n3139), .Z(n3134) );
  AND U2770 ( .A(n3140), .B(n3141), .Z(n3139) );
  XOR U2771 ( .A(n3138), .B(n2711), .Z(n3141) );
  XNOR U2772 ( .A(p_input[3886]), .B(n3142), .Z(n2711) );
  AND U2773 ( .A(n123), .B(n3143), .Z(n3142) );
  XOR U2774 ( .A(p_input[3902]), .B(p_input[3886]), .Z(n3143) );
  XNOR U2775 ( .A(n2708), .B(n3138), .Z(n3140) );
  XOR U2776 ( .A(n3144), .B(n3145), .Z(n2708) );
  AND U2777 ( .A(n120), .B(n3146), .Z(n3145) );
  XOR U2778 ( .A(p_input[3870]), .B(p_input[3854]), .Z(n3146) );
  XOR U2779 ( .A(n3147), .B(n3148), .Z(n3138) );
  AND U2780 ( .A(n3149), .B(n3150), .Z(n3148) );
  XOR U2781 ( .A(n3147), .B(n2723), .Z(n3150) );
  XNOR U2782 ( .A(p_input[3885]), .B(n3151), .Z(n2723) );
  AND U2783 ( .A(n123), .B(n3152), .Z(n3151) );
  XOR U2784 ( .A(p_input[3901]), .B(p_input[3885]), .Z(n3152) );
  XNOR U2785 ( .A(n2720), .B(n3147), .Z(n3149) );
  XOR U2786 ( .A(n3153), .B(n3154), .Z(n2720) );
  AND U2787 ( .A(n120), .B(n3155), .Z(n3154) );
  XOR U2788 ( .A(p_input[3869]), .B(p_input[3853]), .Z(n3155) );
  XOR U2789 ( .A(n3156), .B(n3157), .Z(n3147) );
  AND U2790 ( .A(n3158), .B(n3159), .Z(n3157) );
  XOR U2791 ( .A(n3156), .B(n2735), .Z(n3159) );
  XNOR U2792 ( .A(p_input[3884]), .B(n3160), .Z(n2735) );
  AND U2793 ( .A(n123), .B(n3161), .Z(n3160) );
  XOR U2794 ( .A(p_input[3900]), .B(p_input[3884]), .Z(n3161) );
  XNOR U2795 ( .A(n2732), .B(n3156), .Z(n3158) );
  XOR U2796 ( .A(n3162), .B(n3163), .Z(n2732) );
  AND U2797 ( .A(n120), .B(n3164), .Z(n3163) );
  XOR U2798 ( .A(p_input[3868]), .B(p_input[3852]), .Z(n3164) );
  XOR U2799 ( .A(n3165), .B(n3166), .Z(n3156) );
  AND U2800 ( .A(n3167), .B(n3168), .Z(n3166) );
  XOR U2801 ( .A(n3165), .B(n2747), .Z(n3168) );
  XNOR U2802 ( .A(p_input[3883]), .B(n3169), .Z(n2747) );
  AND U2803 ( .A(n123), .B(n3170), .Z(n3169) );
  XOR U2804 ( .A(p_input[3899]), .B(p_input[3883]), .Z(n3170) );
  XNOR U2805 ( .A(n2744), .B(n3165), .Z(n3167) );
  XOR U2806 ( .A(n3171), .B(n3172), .Z(n2744) );
  AND U2807 ( .A(n120), .B(n3173), .Z(n3172) );
  XOR U2808 ( .A(p_input[3867]), .B(p_input[3851]), .Z(n3173) );
  XOR U2809 ( .A(n3174), .B(n3175), .Z(n3165) );
  AND U2810 ( .A(n3176), .B(n3177), .Z(n3175) );
  XOR U2811 ( .A(n3174), .B(n2759), .Z(n3177) );
  XNOR U2812 ( .A(p_input[3882]), .B(n3178), .Z(n2759) );
  AND U2813 ( .A(n123), .B(n3179), .Z(n3178) );
  XOR U2814 ( .A(p_input[3898]), .B(p_input[3882]), .Z(n3179) );
  XNOR U2815 ( .A(n2756), .B(n3174), .Z(n3176) );
  XOR U2816 ( .A(n3180), .B(n3181), .Z(n2756) );
  AND U2817 ( .A(n120), .B(n3182), .Z(n3181) );
  XOR U2818 ( .A(p_input[3866]), .B(p_input[3850]), .Z(n3182) );
  XOR U2819 ( .A(n3183), .B(n3184), .Z(n3174) );
  AND U2820 ( .A(n3185), .B(n3186), .Z(n3184) );
  XOR U2821 ( .A(n3183), .B(n2771), .Z(n3186) );
  XNOR U2822 ( .A(p_input[3881]), .B(n3187), .Z(n2771) );
  AND U2823 ( .A(n123), .B(n3188), .Z(n3187) );
  XOR U2824 ( .A(p_input[3897]), .B(p_input[3881]), .Z(n3188) );
  XNOR U2825 ( .A(n2768), .B(n3183), .Z(n3185) );
  XOR U2826 ( .A(n3189), .B(n3190), .Z(n2768) );
  AND U2827 ( .A(n120), .B(n3191), .Z(n3190) );
  XOR U2828 ( .A(p_input[3865]), .B(p_input[3849]), .Z(n3191) );
  XOR U2829 ( .A(n3192), .B(n3193), .Z(n3183) );
  AND U2830 ( .A(n3194), .B(n3195), .Z(n3193) );
  XOR U2831 ( .A(n3192), .B(n2783), .Z(n3195) );
  XNOR U2832 ( .A(p_input[3880]), .B(n3196), .Z(n2783) );
  AND U2833 ( .A(n123), .B(n3197), .Z(n3196) );
  XOR U2834 ( .A(p_input[3896]), .B(p_input[3880]), .Z(n3197) );
  XNOR U2835 ( .A(n2780), .B(n3192), .Z(n3194) );
  XOR U2836 ( .A(n3198), .B(n3199), .Z(n2780) );
  AND U2837 ( .A(n120), .B(n3200), .Z(n3199) );
  XOR U2838 ( .A(p_input[3864]), .B(p_input[3848]), .Z(n3200) );
  XOR U2839 ( .A(n3201), .B(n3202), .Z(n3192) );
  AND U2840 ( .A(n3203), .B(n3204), .Z(n3202) );
  XOR U2841 ( .A(n3201), .B(n2795), .Z(n3204) );
  XNOR U2842 ( .A(p_input[3879]), .B(n3205), .Z(n2795) );
  AND U2843 ( .A(n123), .B(n3206), .Z(n3205) );
  XOR U2844 ( .A(p_input[3895]), .B(p_input[3879]), .Z(n3206) );
  XNOR U2845 ( .A(n2792), .B(n3201), .Z(n3203) );
  XOR U2846 ( .A(n3207), .B(n3208), .Z(n2792) );
  AND U2847 ( .A(n120), .B(n3209), .Z(n3208) );
  XOR U2848 ( .A(p_input[3863]), .B(p_input[3847]), .Z(n3209) );
  XOR U2849 ( .A(n3210), .B(n3211), .Z(n3201) );
  AND U2850 ( .A(n3212), .B(n3213), .Z(n3211) );
  XOR U2851 ( .A(n3210), .B(n2807), .Z(n3213) );
  XNOR U2852 ( .A(p_input[3878]), .B(n3214), .Z(n2807) );
  AND U2853 ( .A(n123), .B(n3215), .Z(n3214) );
  XOR U2854 ( .A(p_input[3894]), .B(p_input[3878]), .Z(n3215) );
  XNOR U2855 ( .A(n2804), .B(n3210), .Z(n3212) );
  XOR U2856 ( .A(n3216), .B(n3217), .Z(n2804) );
  AND U2857 ( .A(n120), .B(n3218), .Z(n3217) );
  XOR U2858 ( .A(p_input[3862]), .B(p_input[3846]), .Z(n3218) );
  XOR U2859 ( .A(n3219), .B(n3220), .Z(n3210) );
  AND U2860 ( .A(n3221), .B(n3222), .Z(n3220) );
  XOR U2861 ( .A(n3219), .B(n2819), .Z(n3222) );
  XNOR U2862 ( .A(p_input[3877]), .B(n3223), .Z(n2819) );
  AND U2863 ( .A(n123), .B(n3224), .Z(n3223) );
  XOR U2864 ( .A(p_input[3893]), .B(p_input[3877]), .Z(n3224) );
  XNOR U2865 ( .A(n2816), .B(n3219), .Z(n3221) );
  XOR U2866 ( .A(n3225), .B(n3226), .Z(n2816) );
  AND U2867 ( .A(n120), .B(n3227), .Z(n3226) );
  XOR U2868 ( .A(p_input[3861]), .B(p_input[3845]), .Z(n3227) );
  XOR U2869 ( .A(n3228), .B(n3229), .Z(n3219) );
  AND U2870 ( .A(n3230), .B(n3231), .Z(n3229) );
  XOR U2871 ( .A(n3228), .B(n2831), .Z(n3231) );
  XNOR U2872 ( .A(p_input[3876]), .B(n3232), .Z(n2831) );
  AND U2873 ( .A(n123), .B(n3233), .Z(n3232) );
  XOR U2874 ( .A(p_input[3892]), .B(p_input[3876]), .Z(n3233) );
  XNOR U2875 ( .A(n2828), .B(n3228), .Z(n3230) );
  XOR U2876 ( .A(n3234), .B(n3235), .Z(n2828) );
  AND U2877 ( .A(n120), .B(n3236), .Z(n3235) );
  XOR U2878 ( .A(p_input[3860]), .B(p_input[3844]), .Z(n3236) );
  XOR U2879 ( .A(n3237), .B(n3238), .Z(n3228) );
  AND U2880 ( .A(n3239), .B(n3240), .Z(n3238) );
  XOR U2881 ( .A(n3237), .B(n2843), .Z(n3240) );
  XNOR U2882 ( .A(p_input[3875]), .B(n3241), .Z(n2843) );
  AND U2883 ( .A(n123), .B(n3242), .Z(n3241) );
  XOR U2884 ( .A(p_input[3891]), .B(p_input[3875]), .Z(n3242) );
  XNOR U2885 ( .A(n2840), .B(n3237), .Z(n3239) );
  XOR U2886 ( .A(n3243), .B(n3244), .Z(n2840) );
  AND U2887 ( .A(n120), .B(n3245), .Z(n3244) );
  XOR U2888 ( .A(p_input[3859]), .B(p_input[3843]), .Z(n3245) );
  XOR U2889 ( .A(n3246), .B(n3247), .Z(n3237) );
  AND U2890 ( .A(n3248), .B(n3249), .Z(n3247) );
  XOR U2891 ( .A(n3246), .B(n2855), .Z(n3249) );
  XNOR U2892 ( .A(p_input[3874]), .B(n3250), .Z(n2855) );
  AND U2893 ( .A(n123), .B(n3251), .Z(n3250) );
  XOR U2894 ( .A(p_input[3890]), .B(p_input[3874]), .Z(n3251) );
  XNOR U2895 ( .A(n2852), .B(n3246), .Z(n3248) );
  XOR U2896 ( .A(n3252), .B(n3253), .Z(n2852) );
  AND U2897 ( .A(n120), .B(n3254), .Z(n3253) );
  XOR U2898 ( .A(p_input[3858]), .B(p_input[3842]), .Z(n3254) );
  XOR U2899 ( .A(n3255), .B(n3256), .Z(n3246) );
  AND U2900 ( .A(n3257), .B(n3258), .Z(n3256) );
  XNOR U2901 ( .A(n3259), .B(n2868), .Z(n3258) );
  XNOR U2902 ( .A(p_input[3873]), .B(n3260), .Z(n2868) );
  AND U2903 ( .A(n123), .B(n3261), .Z(n3260) );
  XNOR U2904 ( .A(p_input[3889]), .B(n3262), .Z(n3261) );
  IV U2905 ( .A(p_input[3873]), .Z(n3262) );
  XNOR U2906 ( .A(n2865), .B(n3255), .Z(n3257) );
  XNOR U2907 ( .A(p_input[3841]), .B(n3263), .Z(n2865) );
  AND U2908 ( .A(n120), .B(n3264), .Z(n3263) );
  XOR U2909 ( .A(p_input[3857]), .B(p_input[3841]), .Z(n3264) );
  IV U2910 ( .A(n3259), .Z(n3255) );
  AND U2911 ( .A(n3130), .B(n3133), .Z(n3259) );
  XOR U2912 ( .A(p_input[3872]), .B(n3265), .Z(n3133) );
  AND U2913 ( .A(n123), .B(n3266), .Z(n3265) );
  XOR U2914 ( .A(p_input[3888]), .B(p_input[3872]), .Z(n3266) );
  XOR U2915 ( .A(n3267), .B(n3268), .Z(n123) );
  AND U2916 ( .A(n3269), .B(n3270), .Z(n3268) );
  XNOR U2917 ( .A(p_input[3903]), .B(n3267), .Z(n3270) );
  XOR U2918 ( .A(n3267), .B(p_input[3887]), .Z(n3269) );
  XOR U2919 ( .A(n3271), .B(n3272), .Z(n3267) );
  AND U2920 ( .A(n3273), .B(n3274), .Z(n3272) );
  XNOR U2921 ( .A(p_input[3902]), .B(n3271), .Z(n3274) );
  XOR U2922 ( .A(n3271), .B(p_input[3886]), .Z(n3273) );
  XOR U2923 ( .A(n3275), .B(n3276), .Z(n3271) );
  AND U2924 ( .A(n3277), .B(n3278), .Z(n3276) );
  XNOR U2925 ( .A(p_input[3901]), .B(n3275), .Z(n3278) );
  XOR U2926 ( .A(n3275), .B(p_input[3885]), .Z(n3277) );
  XOR U2927 ( .A(n3279), .B(n3280), .Z(n3275) );
  AND U2928 ( .A(n3281), .B(n3282), .Z(n3280) );
  XNOR U2929 ( .A(p_input[3900]), .B(n3279), .Z(n3282) );
  XOR U2930 ( .A(n3279), .B(p_input[3884]), .Z(n3281) );
  XOR U2931 ( .A(n3283), .B(n3284), .Z(n3279) );
  AND U2932 ( .A(n3285), .B(n3286), .Z(n3284) );
  XNOR U2933 ( .A(p_input[3899]), .B(n3283), .Z(n3286) );
  XOR U2934 ( .A(n3283), .B(p_input[3883]), .Z(n3285) );
  XOR U2935 ( .A(n3287), .B(n3288), .Z(n3283) );
  AND U2936 ( .A(n3289), .B(n3290), .Z(n3288) );
  XNOR U2937 ( .A(p_input[3898]), .B(n3287), .Z(n3290) );
  XOR U2938 ( .A(n3287), .B(p_input[3882]), .Z(n3289) );
  XOR U2939 ( .A(n3291), .B(n3292), .Z(n3287) );
  AND U2940 ( .A(n3293), .B(n3294), .Z(n3292) );
  XNOR U2941 ( .A(p_input[3897]), .B(n3291), .Z(n3294) );
  XOR U2942 ( .A(n3291), .B(p_input[3881]), .Z(n3293) );
  XOR U2943 ( .A(n3295), .B(n3296), .Z(n3291) );
  AND U2944 ( .A(n3297), .B(n3298), .Z(n3296) );
  XNOR U2945 ( .A(p_input[3896]), .B(n3295), .Z(n3298) );
  XOR U2946 ( .A(n3295), .B(p_input[3880]), .Z(n3297) );
  XOR U2947 ( .A(n3299), .B(n3300), .Z(n3295) );
  AND U2948 ( .A(n3301), .B(n3302), .Z(n3300) );
  XNOR U2949 ( .A(p_input[3895]), .B(n3299), .Z(n3302) );
  XOR U2950 ( .A(n3299), .B(p_input[3879]), .Z(n3301) );
  XOR U2951 ( .A(n3303), .B(n3304), .Z(n3299) );
  AND U2952 ( .A(n3305), .B(n3306), .Z(n3304) );
  XNOR U2953 ( .A(p_input[3894]), .B(n3303), .Z(n3306) );
  XOR U2954 ( .A(n3303), .B(p_input[3878]), .Z(n3305) );
  XOR U2955 ( .A(n3307), .B(n3308), .Z(n3303) );
  AND U2956 ( .A(n3309), .B(n3310), .Z(n3308) );
  XNOR U2957 ( .A(p_input[3893]), .B(n3307), .Z(n3310) );
  XOR U2958 ( .A(n3307), .B(p_input[3877]), .Z(n3309) );
  XOR U2959 ( .A(n3311), .B(n3312), .Z(n3307) );
  AND U2960 ( .A(n3313), .B(n3314), .Z(n3312) );
  XNOR U2961 ( .A(p_input[3892]), .B(n3311), .Z(n3314) );
  XOR U2962 ( .A(n3311), .B(p_input[3876]), .Z(n3313) );
  XOR U2963 ( .A(n3315), .B(n3316), .Z(n3311) );
  AND U2964 ( .A(n3317), .B(n3318), .Z(n3316) );
  XNOR U2965 ( .A(p_input[3891]), .B(n3315), .Z(n3318) );
  XOR U2966 ( .A(n3315), .B(p_input[3875]), .Z(n3317) );
  XOR U2967 ( .A(n3319), .B(n3320), .Z(n3315) );
  AND U2968 ( .A(n3321), .B(n3322), .Z(n3320) );
  XNOR U2969 ( .A(p_input[3890]), .B(n3319), .Z(n3322) );
  XOR U2970 ( .A(n3319), .B(p_input[3874]), .Z(n3321) );
  XNOR U2971 ( .A(n3323), .B(n3324), .Z(n3319) );
  AND U2972 ( .A(n3325), .B(n3326), .Z(n3324) );
  XOR U2973 ( .A(p_input[3889]), .B(n3323), .Z(n3326) );
  XNOR U2974 ( .A(p_input[3873]), .B(n3323), .Z(n3325) );
  AND U2975 ( .A(p_input[3888]), .B(n3327), .Z(n3323) );
  IV U2976 ( .A(p_input[3872]), .Z(n3327) );
  XNOR U2977 ( .A(p_input[3840]), .B(n3328), .Z(n3130) );
  AND U2978 ( .A(n120), .B(n3329), .Z(n3328) );
  XOR U2979 ( .A(p_input[3856]), .B(p_input[3840]), .Z(n3329) );
  XOR U2980 ( .A(n3330), .B(n3331), .Z(n120) );
  AND U2981 ( .A(n3332), .B(n3333), .Z(n3331) );
  XNOR U2982 ( .A(p_input[3871]), .B(n3330), .Z(n3333) );
  XOR U2983 ( .A(n3330), .B(p_input[3855]), .Z(n3332) );
  XOR U2984 ( .A(n3334), .B(n3335), .Z(n3330) );
  AND U2985 ( .A(n3336), .B(n3337), .Z(n3335) );
  XNOR U2986 ( .A(p_input[3870]), .B(n3334), .Z(n3337) );
  XNOR U2987 ( .A(n3334), .B(n3144), .Z(n3336) );
  IV U2988 ( .A(p_input[3854]), .Z(n3144) );
  XOR U2989 ( .A(n3338), .B(n3339), .Z(n3334) );
  AND U2990 ( .A(n3340), .B(n3341), .Z(n3339) );
  XNOR U2991 ( .A(p_input[3869]), .B(n3338), .Z(n3341) );
  XNOR U2992 ( .A(n3338), .B(n3153), .Z(n3340) );
  IV U2993 ( .A(p_input[3853]), .Z(n3153) );
  XOR U2994 ( .A(n3342), .B(n3343), .Z(n3338) );
  AND U2995 ( .A(n3344), .B(n3345), .Z(n3343) );
  XNOR U2996 ( .A(p_input[3868]), .B(n3342), .Z(n3345) );
  XNOR U2997 ( .A(n3342), .B(n3162), .Z(n3344) );
  IV U2998 ( .A(p_input[3852]), .Z(n3162) );
  XOR U2999 ( .A(n3346), .B(n3347), .Z(n3342) );
  AND U3000 ( .A(n3348), .B(n3349), .Z(n3347) );
  XNOR U3001 ( .A(p_input[3867]), .B(n3346), .Z(n3349) );
  XNOR U3002 ( .A(n3346), .B(n3171), .Z(n3348) );
  IV U3003 ( .A(p_input[3851]), .Z(n3171) );
  XOR U3004 ( .A(n3350), .B(n3351), .Z(n3346) );
  AND U3005 ( .A(n3352), .B(n3353), .Z(n3351) );
  XNOR U3006 ( .A(p_input[3866]), .B(n3350), .Z(n3353) );
  XNOR U3007 ( .A(n3350), .B(n3180), .Z(n3352) );
  IV U3008 ( .A(p_input[3850]), .Z(n3180) );
  XOR U3009 ( .A(n3354), .B(n3355), .Z(n3350) );
  AND U3010 ( .A(n3356), .B(n3357), .Z(n3355) );
  XNOR U3011 ( .A(p_input[3865]), .B(n3354), .Z(n3357) );
  XNOR U3012 ( .A(n3354), .B(n3189), .Z(n3356) );
  IV U3013 ( .A(p_input[3849]), .Z(n3189) );
  XOR U3014 ( .A(n3358), .B(n3359), .Z(n3354) );
  AND U3015 ( .A(n3360), .B(n3361), .Z(n3359) );
  XNOR U3016 ( .A(p_input[3864]), .B(n3358), .Z(n3361) );
  XNOR U3017 ( .A(n3358), .B(n3198), .Z(n3360) );
  IV U3018 ( .A(p_input[3848]), .Z(n3198) );
  XOR U3019 ( .A(n3362), .B(n3363), .Z(n3358) );
  AND U3020 ( .A(n3364), .B(n3365), .Z(n3363) );
  XNOR U3021 ( .A(p_input[3863]), .B(n3362), .Z(n3365) );
  XNOR U3022 ( .A(n3362), .B(n3207), .Z(n3364) );
  IV U3023 ( .A(p_input[3847]), .Z(n3207) );
  XOR U3024 ( .A(n3366), .B(n3367), .Z(n3362) );
  AND U3025 ( .A(n3368), .B(n3369), .Z(n3367) );
  XNOR U3026 ( .A(p_input[3862]), .B(n3366), .Z(n3369) );
  XNOR U3027 ( .A(n3366), .B(n3216), .Z(n3368) );
  IV U3028 ( .A(p_input[3846]), .Z(n3216) );
  XOR U3029 ( .A(n3370), .B(n3371), .Z(n3366) );
  AND U3030 ( .A(n3372), .B(n3373), .Z(n3371) );
  XNOR U3031 ( .A(p_input[3861]), .B(n3370), .Z(n3373) );
  XNOR U3032 ( .A(n3370), .B(n3225), .Z(n3372) );
  IV U3033 ( .A(p_input[3845]), .Z(n3225) );
  XOR U3034 ( .A(n3374), .B(n3375), .Z(n3370) );
  AND U3035 ( .A(n3376), .B(n3377), .Z(n3375) );
  XNOR U3036 ( .A(p_input[3860]), .B(n3374), .Z(n3377) );
  XNOR U3037 ( .A(n3374), .B(n3234), .Z(n3376) );
  IV U3038 ( .A(p_input[3844]), .Z(n3234) );
  XOR U3039 ( .A(n3378), .B(n3379), .Z(n3374) );
  AND U3040 ( .A(n3380), .B(n3381), .Z(n3379) );
  XNOR U3041 ( .A(p_input[3859]), .B(n3378), .Z(n3381) );
  XNOR U3042 ( .A(n3378), .B(n3243), .Z(n3380) );
  IV U3043 ( .A(p_input[3843]), .Z(n3243) );
  XOR U3044 ( .A(n3382), .B(n3383), .Z(n3378) );
  AND U3045 ( .A(n3384), .B(n3385), .Z(n3383) );
  XNOR U3046 ( .A(p_input[3858]), .B(n3382), .Z(n3385) );
  XNOR U3047 ( .A(n3382), .B(n3252), .Z(n3384) );
  IV U3048 ( .A(p_input[3842]), .Z(n3252) );
  XNOR U3049 ( .A(n3386), .B(n3387), .Z(n3382) );
  AND U3050 ( .A(n3388), .B(n3389), .Z(n3387) );
  XOR U3051 ( .A(p_input[3857]), .B(n3386), .Z(n3389) );
  XNOR U3052 ( .A(p_input[3841]), .B(n3386), .Z(n3388) );
  AND U3053 ( .A(p_input[3856]), .B(n3390), .Z(n3386) );
  IV U3054 ( .A(p_input[3840]), .Z(n3390) );
  XOR U3055 ( .A(n3391), .B(n3392), .Z(n1618) );
  AND U3056 ( .A(n917), .B(n3393), .Z(n3392) );
  XNOR U3057 ( .A(n3394), .B(n3391), .Z(n3393) );
  XOR U3058 ( .A(n3395), .B(n3396), .Z(n917) );
  AND U3059 ( .A(n3397), .B(n3398), .Z(n3396) );
  XNOR U3060 ( .A(n1633), .B(n3395), .Z(n3398) );
  AND U3061 ( .A(n3399), .B(n3400), .Z(n1633) );
  XNOR U3062 ( .A(n3395), .B(n1630), .Z(n3397) );
  IV U3063 ( .A(n3401), .Z(n1630) );
  AND U3064 ( .A(n3402), .B(n3403), .Z(n3401) );
  XOR U3065 ( .A(n3404), .B(n3405), .Z(n3395) );
  AND U3066 ( .A(n3406), .B(n3407), .Z(n3405) );
  XOR U3067 ( .A(n3404), .B(n1645), .Z(n3407) );
  XOR U3068 ( .A(n3408), .B(n3409), .Z(n1645) );
  AND U3069 ( .A(n739), .B(n3410), .Z(n3409) );
  XOR U3070 ( .A(n3411), .B(n3408), .Z(n3410) );
  XNOR U3071 ( .A(n1642), .B(n3404), .Z(n3406) );
  XOR U3072 ( .A(n3412), .B(n3413), .Z(n1642) );
  AND U3073 ( .A(n736), .B(n3414), .Z(n3413) );
  XOR U3074 ( .A(n3415), .B(n3412), .Z(n3414) );
  XOR U3075 ( .A(n3416), .B(n3417), .Z(n3404) );
  AND U3076 ( .A(n3418), .B(n3419), .Z(n3417) );
  XOR U3077 ( .A(n3416), .B(n1657), .Z(n3419) );
  XOR U3078 ( .A(n3420), .B(n3421), .Z(n1657) );
  AND U3079 ( .A(n739), .B(n3422), .Z(n3421) );
  XOR U3080 ( .A(n3423), .B(n3420), .Z(n3422) );
  XNOR U3081 ( .A(n1654), .B(n3416), .Z(n3418) );
  XOR U3082 ( .A(n3424), .B(n3425), .Z(n1654) );
  AND U3083 ( .A(n736), .B(n3426), .Z(n3425) );
  XOR U3084 ( .A(n3427), .B(n3424), .Z(n3426) );
  XOR U3085 ( .A(n3428), .B(n3429), .Z(n3416) );
  AND U3086 ( .A(n3430), .B(n3431), .Z(n3429) );
  XOR U3087 ( .A(n3428), .B(n1669), .Z(n3431) );
  XOR U3088 ( .A(n3432), .B(n3433), .Z(n1669) );
  AND U3089 ( .A(n739), .B(n3434), .Z(n3433) );
  XOR U3090 ( .A(n3435), .B(n3432), .Z(n3434) );
  XNOR U3091 ( .A(n1666), .B(n3428), .Z(n3430) );
  XOR U3092 ( .A(n3436), .B(n3437), .Z(n1666) );
  AND U3093 ( .A(n736), .B(n3438), .Z(n3437) );
  XOR U3094 ( .A(n3439), .B(n3436), .Z(n3438) );
  XOR U3095 ( .A(n3440), .B(n3441), .Z(n3428) );
  AND U3096 ( .A(n3442), .B(n3443), .Z(n3441) );
  XOR U3097 ( .A(n3440), .B(n1681), .Z(n3443) );
  XOR U3098 ( .A(n3444), .B(n3445), .Z(n1681) );
  AND U3099 ( .A(n739), .B(n3446), .Z(n3445) );
  XOR U3100 ( .A(n3447), .B(n3444), .Z(n3446) );
  XNOR U3101 ( .A(n1678), .B(n3440), .Z(n3442) );
  XOR U3102 ( .A(n3448), .B(n3449), .Z(n1678) );
  AND U3103 ( .A(n736), .B(n3450), .Z(n3449) );
  XOR U3104 ( .A(n3451), .B(n3448), .Z(n3450) );
  XOR U3105 ( .A(n3452), .B(n3453), .Z(n3440) );
  AND U3106 ( .A(n3454), .B(n3455), .Z(n3453) );
  XOR U3107 ( .A(n3452), .B(n1693), .Z(n3455) );
  XOR U3108 ( .A(n3456), .B(n3457), .Z(n1693) );
  AND U3109 ( .A(n739), .B(n3458), .Z(n3457) );
  XOR U3110 ( .A(n3459), .B(n3456), .Z(n3458) );
  XNOR U3111 ( .A(n1690), .B(n3452), .Z(n3454) );
  XOR U3112 ( .A(n3460), .B(n3461), .Z(n1690) );
  AND U3113 ( .A(n736), .B(n3462), .Z(n3461) );
  XOR U3114 ( .A(n3463), .B(n3460), .Z(n3462) );
  XOR U3115 ( .A(n3464), .B(n3465), .Z(n3452) );
  AND U3116 ( .A(n3466), .B(n3467), .Z(n3465) );
  XOR U3117 ( .A(n3464), .B(n1705), .Z(n3467) );
  XOR U3118 ( .A(n3468), .B(n3469), .Z(n1705) );
  AND U3119 ( .A(n739), .B(n3470), .Z(n3469) );
  XOR U3120 ( .A(n3471), .B(n3468), .Z(n3470) );
  XNOR U3121 ( .A(n1702), .B(n3464), .Z(n3466) );
  XOR U3122 ( .A(n3472), .B(n3473), .Z(n1702) );
  AND U3123 ( .A(n736), .B(n3474), .Z(n3473) );
  XOR U3124 ( .A(n3475), .B(n3472), .Z(n3474) );
  XOR U3125 ( .A(n3476), .B(n3477), .Z(n3464) );
  AND U3126 ( .A(n3478), .B(n3479), .Z(n3477) );
  XOR U3127 ( .A(n3476), .B(n1717), .Z(n3479) );
  XOR U3128 ( .A(n3480), .B(n3481), .Z(n1717) );
  AND U3129 ( .A(n739), .B(n3482), .Z(n3481) );
  XOR U3130 ( .A(n3483), .B(n3480), .Z(n3482) );
  XNOR U3131 ( .A(n1714), .B(n3476), .Z(n3478) );
  XOR U3132 ( .A(n3484), .B(n3485), .Z(n1714) );
  AND U3133 ( .A(n736), .B(n3486), .Z(n3485) );
  XOR U3134 ( .A(n3487), .B(n3484), .Z(n3486) );
  XOR U3135 ( .A(n3488), .B(n3489), .Z(n3476) );
  AND U3136 ( .A(n3490), .B(n3491), .Z(n3489) );
  XOR U3137 ( .A(n3488), .B(n1729), .Z(n3491) );
  XOR U3138 ( .A(n3492), .B(n3493), .Z(n1729) );
  AND U3139 ( .A(n739), .B(n3494), .Z(n3493) );
  XOR U3140 ( .A(n3495), .B(n3492), .Z(n3494) );
  XNOR U3141 ( .A(n1726), .B(n3488), .Z(n3490) );
  XOR U3142 ( .A(n3496), .B(n3497), .Z(n1726) );
  AND U3143 ( .A(n736), .B(n3498), .Z(n3497) );
  XOR U3144 ( .A(n3499), .B(n3496), .Z(n3498) );
  XOR U3145 ( .A(n3500), .B(n3501), .Z(n3488) );
  AND U3146 ( .A(n3502), .B(n3503), .Z(n3501) );
  XOR U3147 ( .A(n3500), .B(n1741), .Z(n3503) );
  XOR U3148 ( .A(n3504), .B(n3505), .Z(n1741) );
  AND U3149 ( .A(n739), .B(n3506), .Z(n3505) );
  XOR U3150 ( .A(n3507), .B(n3504), .Z(n3506) );
  XNOR U3151 ( .A(n1738), .B(n3500), .Z(n3502) );
  XOR U3152 ( .A(n3508), .B(n3509), .Z(n1738) );
  AND U3153 ( .A(n736), .B(n3510), .Z(n3509) );
  XOR U3154 ( .A(n3511), .B(n3508), .Z(n3510) );
  XOR U3155 ( .A(n3512), .B(n3513), .Z(n3500) );
  AND U3156 ( .A(n3514), .B(n3515), .Z(n3513) );
  XOR U3157 ( .A(n3512), .B(n1753), .Z(n3515) );
  XOR U3158 ( .A(n3516), .B(n3517), .Z(n1753) );
  AND U3159 ( .A(n739), .B(n3518), .Z(n3517) );
  XOR U3160 ( .A(n3519), .B(n3516), .Z(n3518) );
  XNOR U3161 ( .A(n1750), .B(n3512), .Z(n3514) );
  XOR U3162 ( .A(n3520), .B(n3521), .Z(n1750) );
  AND U3163 ( .A(n736), .B(n3522), .Z(n3521) );
  XOR U3164 ( .A(n3523), .B(n3520), .Z(n3522) );
  XOR U3165 ( .A(n3524), .B(n3525), .Z(n3512) );
  AND U3166 ( .A(n3526), .B(n3527), .Z(n3525) );
  XOR U3167 ( .A(n3524), .B(n1765), .Z(n3527) );
  XOR U3168 ( .A(n3528), .B(n3529), .Z(n1765) );
  AND U3169 ( .A(n739), .B(n3530), .Z(n3529) );
  XOR U3170 ( .A(n3531), .B(n3528), .Z(n3530) );
  XNOR U3171 ( .A(n1762), .B(n3524), .Z(n3526) );
  XOR U3172 ( .A(n3532), .B(n3533), .Z(n1762) );
  AND U3173 ( .A(n736), .B(n3534), .Z(n3533) );
  XOR U3174 ( .A(n3535), .B(n3532), .Z(n3534) );
  XOR U3175 ( .A(n3536), .B(n3537), .Z(n3524) );
  AND U3176 ( .A(n3538), .B(n3539), .Z(n3537) );
  XOR U3177 ( .A(n3536), .B(n1777), .Z(n3539) );
  XOR U3178 ( .A(n3540), .B(n3541), .Z(n1777) );
  AND U3179 ( .A(n739), .B(n3542), .Z(n3541) );
  XOR U3180 ( .A(n3543), .B(n3540), .Z(n3542) );
  XNOR U3181 ( .A(n1774), .B(n3536), .Z(n3538) );
  XOR U3182 ( .A(n3544), .B(n3545), .Z(n1774) );
  AND U3183 ( .A(n736), .B(n3546), .Z(n3545) );
  XOR U3184 ( .A(n3547), .B(n3544), .Z(n3546) );
  XOR U3185 ( .A(n3548), .B(n3549), .Z(n3536) );
  AND U3186 ( .A(n3550), .B(n3551), .Z(n3549) );
  XOR U3187 ( .A(n3548), .B(n1789), .Z(n3551) );
  XOR U3188 ( .A(n3552), .B(n3553), .Z(n1789) );
  AND U3189 ( .A(n739), .B(n3554), .Z(n3553) );
  XOR U3190 ( .A(n3555), .B(n3552), .Z(n3554) );
  XNOR U3191 ( .A(n1786), .B(n3548), .Z(n3550) );
  XOR U3192 ( .A(n3556), .B(n3557), .Z(n1786) );
  AND U3193 ( .A(n736), .B(n3558), .Z(n3557) );
  XOR U3194 ( .A(n3559), .B(n3556), .Z(n3558) );
  XOR U3195 ( .A(n3560), .B(n3561), .Z(n3548) );
  AND U3196 ( .A(n3562), .B(n3563), .Z(n3561) );
  XNOR U3197 ( .A(n3564), .B(n1802), .Z(n3563) );
  XOR U3198 ( .A(n3565), .B(n3566), .Z(n1802) );
  AND U3199 ( .A(n739), .B(n3567), .Z(n3566) );
  XOR U3200 ( .A(n3565), .B(n3568), .Z(n3567) );
  XNOR U3201 ( .A(n1799), .B(n3560), .Z(n3562) );
  XOR U3202 ( .A(n3569), .B(n3570), .Z(n1799) );
  AND U3203 ( .A(n736), .B(n3571), .Z(n3570) );
  XOR U3204 ( .A(n3569), .B(n3572), .Z(n3571) );
  IV U3205 ( .A(n3564), .Z(n3560) );
  AND U3206 ( .A(n3391), .B(n3394), .Z(n3564) );
  XNOR U3207 ( .A(n3573), .B(n3574), .Z(n3394) );
  AND U3208 ( .A(n739), .B(n3575), .Z(n3574) );
  XNOR U3209 ( .A(n3576), .B(n3573), .Z(n3575) );
  XOR U3210 ( .A(n3577), .B(n3578), .Z(n739) );
  AND U3211 ( .A(n3579), .B(n3580), .Z(n3578) );
  XNOR U3212 ( .A(n3399), .B(n3577), .Z(n3580) );
  AND U3213 ( .A(n3581), .B(n3582), .Z(n3399) );
  XOR U3214 ( .A(n3577), .B(n3400), .Z(n3579) );
  AND U3215 ( .A(n3583), .B(n3584), .Z(n3400) );
  XOR U3216 ( .A(n3585), .B(n3586), .Z(n3577) );
  AND U3217 ( .A(n3587), .B(n3588), .Z(n3586) );
  XOR U3218 ( .A(n3585), .B(n3411), .Z(n3588) );
  XOR U3219 ( .A(n3589), .B(n3590), .Z(n3411) );
  AND U3220 ( .A(n371), .B(n3591), .Z(n3590) );
  XOR U3221 ( .A(n3592), .B(n3589), .Z(n3591) );
  XNOR U3222 ( .A(n3408), .B(n3585), .Z(n3587) );
  XOR U3223 ( .A(n3593), .B(n3594), .Z(n3408) );
  AND U3224 ( .A(n369), .B(n3595), .Z(n3594) );
  XOR U3225 ( .A(n3596), .B(n3593), .Z(n3595) );
  XOR U3226 ( .A(n3597), .B(n3598), .Z(n3585) );
  AND U3227 ( .A(n3599), .B(n3600), .Z(n3598) );
  XOR U3228 ( .A(n3597), .B(n3423), .Z(n3600) );
  XOR U3229 ( .A(n3601), .B(n3602), .Z(n3423) );
  AND U3230 ( .A(n371), .B(n3603), .Z(n3602) );
  XOR U3231 ( .A(n3604), .B(n3601), .Z(n3603) );
  XNOR U3232 ( .A(n3420), .B(n3597), .Z(n3599) );
  XOR U3233 ( .A(n3605), .B(n3606), .Z(n3420) );
  AND U3234 ( .A(n369), .B(n3607), .Z(n3606) );
  XOR U3235 ( .A(n3608), .B(n3605), .Z(n3607) );
  XOR U3236 ( .A(n3609), .B(n3610), .Z(n3597) );
  AND U3237 ( .A(n3611), .B(n3612), .Z(n3610) );
  XOR U3238 ( .A(n3609), .B(n3435), .Z(n3612) );
  XOR U3239 ( .A(n3613), .B(n3614), .Z(n3435) );
  AND U3240 ( .A(n371), .B(n3615), .Z(n3614) );
  XOR U3241 ( .A(n3616), .B(n3613), .Z(n3615) );
  XNOR U3242 ( .A(n3432), .B(n3609), .Z(n3611) );
  XOR U3243 ( .A(n3617), .B(n3618), .Z(n3432) );
  AND U3244 ( .A(n369), .B(n3619), .Z(n3618) );
  XOR U3245 ( .A(n3620), .B(n3617), .Z(n3619) );
  XOR U3246 ( .A(n3621), .B(n3622), .Z(n3609) );
  AND U3247 ( .A(n3623), .B(n3624), .Z(n3622) );
  XOR U3248 ( .A(n3621), .B(n3447), .Z(n3624) );
  XOR U3249 ( .A(n3625), .B(n3626), .Z(n3447) );
  AND U3250 ( .A(n371), .B(n3627), .Z(n3626) );
  XOR U3251 ( .A(n3628), .B(n3625), .Z(n3627) );
  XNOR U3252 ( .A(n3444), .B(n3621), .Z(n3623) );
  XOR U3253 ( .A(n3629), .B(n3630), .Z(n3444) );
  AND U3254 ( .A(n369), .B(n3631), .Z(n3630) );
  XOR U3255 ( .A(n3632), .B(n3629), .Z(n3631) );
  XOR U3256 ( .A(n3633), .B(n3634), .Z(n3621) );
  AND U3257 ( .A(n3635), .B(n3636), .Z(n3634) );
  XOR U3258 ( .A(n3633), .B(n3459), .Z(n3636) );
  XOR U3259 ( .A(n3637), .B(n3638), .Z(n3459) );
  AND U3260 ( .A(n371), .B(n3639), .Z(n3638) );
  XOR U3261 ( .A(n3640), .B(n3637), .Z(n3639) );
  XNOR U3262 ( .A(n3456), .B(n3633), .Z(n3635) );
  XOR U3263 ( .A(n3641), .B(n3642), .Z(n3456) );
  AND U3264 ( .A(n369), .B(n3643), .Z(n3642) );
  XOR U3265 ( .A(n3644), .B(n3641), .Z(n3643) );
  XOR U3266 ( .A(n3645), .B(n3646), .Z(n3633) );
  AND U3267 ( .A(n3647), .B(n3648), .Z(n3646) );
  XOR U3268 ( .A(n3645), .B(n3471), .Z(n3648) );
  XOR U3269 ( .A(n3649), .B(n3650), .Z(n3471) );
  AND U3270 ( .A(n371), .B(n3651), .Z(n3650) );
  XOR U3271 ( .A(n3652), .B(n3649), .Z(n3651) );
  XNOR U3272 ( .A(n3468), .B(n3645), .Z(n3647) );
  XOR U3273 ( .A(n3653), .B(n3654), .Z(n3468) );
  AND U3274 ( .A(n369), .B(n3655), .Z(n3654) );
  XOR U3275 ( .A(n3656), .B(n3653), .Z(n3655) );
  XOR U3276 ( .A(n3657), .B(n3658), .Z(n3645) );
  AND U3277 ( .A(n3659), .B(n3660), .Z(n3658) );
  XOR U3278 ( .A(n3657), .B(n3483), .Z(n3660) );
  XOR U3279 ( .A(n3661), .B(n3662), .Z(n3483) );
  AND U3280 ( .A(n371), .B(n3663), .Z(n3662) );
  XOR U3281 ( .A(n3664), .B(n3661), .Z(n3663) );
  XNOR U3282 ( .A(n3480), .B(n3657), .Z(n3659) );
  XOR U3283 ( .A(n3665), .B(n3666), .Z(n3480) );
  AND U3284 ( .A(n369), .B(n3667), .Z(n3666) );
  XOR U3285 ( .A(n3668), .B(n3665), .Z(n3667) );
  XOR U3286 ( .A(n3669), .B(n3670), .Z(n3657) );
  AND U3287 ( .A(n3671), .B(n3672), .Z(n3670) );
  XOR U3288 ( .A(n3669), .B(n3495), .Z(n3672) );
  XOR U3289 ( .A(n3673), .B(n3674), .Z(n3495) );
  AND U3290 ( .A(n371), .B(n3675), .Z(n3674) );
  XOR U3291 ( .A(n3676), .B(n3673), .Z(n3675) );
  XNOR U3292 ( .A(n3492), .B(n3669), .Z(n3671) );
  XOR U3293 ( .A(n3677), .B(n3678), .Z(n3492) );
  AND U3294 ( .A(n369), .B(n3679), .Z(n3678) );
  XOR U3295 ( .A(n3680), .B(n3677), .Z(n3679) );
  XOR U3296 ( .A(n3681), .B(n3682), .Z(n3669) );
  AND U3297 ( .A(n3683), .B(n3684), .Z(n3682) );
  XOR U3298 ( .A(n3681), .B(n3507), .Z(n3684) );
  XOR U3299 ( .A(n3685), .B(n3686), .Z(n3507) );
  AND U3300 ( .A(n371), .B(n3687), .Z(n3686) );
  XOR U3301 ( .A(n3688), .B(n3685), .Z(n3687) );
  XNOR U3302 ( .A(n3504), .B(n3681), .Z(n3683) );
  XOR U3303 ( .A(n3689), .B(n3690), .Z(n3504) );
  AND U3304 ( .A(n369), .B(n3691), .Z(n3690) );
  XOR U3305 ( .A(n3692), .B(n3689), .Z(n3691) );
  XOR U3306 ( .A(n3693), .B(n3694), .Z(n3681) );
  AND U3307 ( .A(n3695), .B(n3696), .Z(n3694) );
  XOR U3308 ( .A(n3693), .B(n3519), .Z(n3696) );
  XOR U3309 ( .A(n3697), .B(n3698), .Z(n3519) );
  AND U3310 ( .A(n371), .B(n3699), .Z(n3698) );
  XOR U3311 ( .A(n3700), .B(n3697), .Z(n3699) );
  XNOR U3312 ( .A(n3516), .B(n3693), .Z(n3695) );
  XOR U3313 ( .A(n3701), .B(n3702), .Z(n3516) );
  AND U3314 ( .A(n369), .B(n3703), .Z(n3702) );
  XOR U3315 ( .A(n3704), .B(n3701), .Z(n3703) );
  XOR U3316 ( .A(n3705), .B(n3706), .Z(n3693) );
  AND U3317 ( .A(n3707), .B(n3708), .Z(n3706) );
  XOR U3318 ( .A(n3705), .B(n3531), .Z(n3708) );
  XOR U3319 ( .A(n3709), .B(n3710), .Z(n3531) );
  AND U3320 ( .A(n371), .B(n3711), .Z(n3710) );
  XOR U3321 ( .A(n3712), .B(n3709), .Z(n3711) );
  XNOR U3322 ( .A(n3528), .B(n3705), .Z(n3707) );
  XOR U3323 ( .A(n3713), .B(n3714), .Z(n3528) );
  AND U3324 ( .A(n369), .B(n3715), .Z(n3714) );
  XOR U3325 ( .A(n3716), .B(n3713), .Z(n3715) );
  XOR U3326 ( .A(n3717), .B(n3718), .Z(n3705) );
  AND U3327 ( .A(n3719), .B(n3720), .Z(n3718) );
  XOR U3328 ( .A(n3717), .B(n3543), .Z(n3720) );
  XOR U3329 ( .A(n3721), .B(n3722), .Z(n3543) );
  AND U3330 ( .A(n371), .B(n3723), .Z(n3722) );
  XOR U3331 ( .A(n3724), .B(n3721), .Z(n3723) );
  XNOR U3332 ( .A(n3540), .B(n3717), .Z(n3719) );
  XOR U3333 ( .A(n3725), .B(n3726), .Z(n3540) );
  AND U3334 ( .A(n369), .B(n3727), .Z(n3726) );
  XOR U3335 ( .A(n3728), .B(n3725), .Z(n3727) );
  XOR U3336 ( .A(n3729), .B(n3730), .Z(n3717) );
  AND U3337 ( .A(n3731), .B(n3732), .Z(n3730) );
  XOR U3338 ( .A(n3729), .B(n3555), .Z(n3732) );
  XOR U3339 ( .A(n3733), .B(n3734), .Z(n3555) );
  AND U3340 ( .A(n371), .B(n3735), .Z(n3734) );
  XOR U3341 ( .A(n3736), .B(n3733), .Z(n3735) );
  XNOR U3342 ( .A(n3552), .B(n3729), .Z(n3731) );
  XOR U3343 ( .A(n3737), .B(n3738), .Z(n3552) );
  AND U3344 ( .A(n369), .B(n3739), .Z(n3738) );
  XOR U3345 ( .A(n3740), .B(n3737), .Z(n3739) );
  XOR U3346 ( .A(n3741), .B(n3742), .Z(n3729) );
  AND U3347 ( .A(n3743), .B(n3744), .Z(n3742) );
  XNOR U3348 ( .A(n3745), .B(n3568), .Z(n3744) );
  XOR U3349 ( .A(n3746), .B(n3747), .Z(n3568) );
  AND U3350 ( .A(n371), .B(n3748), .Z(n3747) );
  XOR U3351 ( .A(n3746), .B(n3749), .Z(n3748) );
  XNOR U3352 ( .A(n3565), .B(n3741), .Z(n3743) );
  XOR U3353 ( .A(n3750), .B(n3751), .Z(n3565) );
  AND U3354 ( .A(n369), .B(n3752), .Z(n3751) );
  XOR U3355 ( .A(n3750), .B(n3753), .Z(n3752) );
  IV U3356 ( .A(n3745), .Z(n3741) );
  AND U3357 ( .A(n3573), .B(n3576), .Z(n3745) );
  XNOR U3358 ( .A(n3754), .B(n3755), .Z(n3576) );
  AND U3359 ( .A(n371), .B(n3756), .Z(n3755) );
  XNOR U3360 ( .A(n3757), .B(n3754), .Z(n3756) );
  XOR U3361 ( .A(n3758), .B(n3759), .Z(n371) );
  AND U3362 ( .A(n3760), .B(n3761), .Z(n3759) );
  XNOR U3363 ( .A(n3581), .B(n3758), .Z(n3761) );
  AND U3364 ( .A(p_input[3839]), .B(p_input[3823]), .Z(n3581) );
  XOR U3365 ( .A(n3758), .B(n3582), .Z(n3760) );
  AND U3366 ( .A(p_input[3807]), .B(p_input[3791]), .Z(n3582) );
  XOR U3367 ( .A(n3762), .B(n3763), .Z(n3758) );
  AND U3368 ( .A(n3764), .B(n3765), .Z(n3763) );
  XOR U3369 ( .A(n3762), .B(n3592), .Z(n3765) );
  XNOR U3370 ( .A(p_input[3822]), .B(n3766), .Z(n3592) );
  AND U3371 ( .A(n135), .B(n3767), .Z(n3766) );
  XOR U3372 ( .A(p_input[3838]), .B(p_input[3822]), .Z(n3767) );
  XNOR U3373 ( .A(n3589), .B(n3762), .Z(n3764) );
  XOR U3374 ( .A(n3768), .B(n3769), .Z(n3589) );
  AND U3375 ( .A(n133), .B(n3770), .Z(n3769) );
  XOR U3376 ( .A(p_input[3806]), .B(p_input[3790]), .Z(n3770) );
  XOR U3377 ( .A(n3771), .B(n3772), .Z(n3762) );
  AND U3378 ( .A(n3773), .B(n3774), .Z(n3772) );
  XOR U3379 ( .A(n3771), .B(n3604), .Z(n3774) );
  XNOR U3380 ( .A(p_input[3821]), .B(n3775), .Z(n3604) );
  AND U3381 ( .A(n135), .B(n3776), .Z(n3775) );
  XOR U3382 ( .A(p_input[3837]), .B(p_input[3821]), .Z(n3776) );
  XNOR U3383 ( .A(n3601), .B(n3771), .Z(n3773) );
  XOR U3384 ( .A(n3777), .B(n3778), .Z(n3601) );
  AND U3385 ( .A(n133), .B(n3779), .Z(n3778) );
  XOR U3386 ( .A(p_input[3805]), .B(p_input[3789]), .Z(n3779) );
  XOR U3387 ( .A(n3780), .B(n3781), .Z(n3771) );
  AND U3388 ( .A(n3782), .B(n3783), .Z(n3781) );
  XOR U3389 ( .A(n3780), .B(n3616), .Z(n3783) );
  XNOR U3390 ( .A(p_input[3820]), .B(n3784), .Z(n3616) );
  AND U3391 ( .A(n135), .B(n3785), .Z(n3784) );
  XOR U3392 ( .A(p_input[3836]), .B(p_input[3820]), .Z(n3785) );
  XNOR U3393 ( .A(n3613), .B(n3780), .Z(n3782) );
  XOR U3394 ( .A(n3786), .B(n3787), .Z(n3613) );
  AND U3395 ( .A(n133), .B(n3788), .Z(n3787) );
  XOR U3396 ( .A(p_input[3804]), .B(p_input[3788]), .Z(n3788) );
  XOR U3397 ( .A(n3789), .B(n3790), .Z(n3780) );
  AND U3398 ( .A(n3791), .B(n3792), .Z(n3790) );
  XOR U3399 ( .A(n3789), .B(n3628), .Z(n3792) );
  XNOR U3400 ( .A(p_input[3819]), .B(n3793), .Z(n3628) );
  AND U3401 ( .A(n135), .B(n3794), .Z(n3793) );
  XOR U3402 ( .A(p_input[3835]), .B(p_input[3819]), .Z(n3794) );
  XNOR U3403 ( .A(n3625), .B(n3789), .Z(n3791) );
  XOR U3404 ( .A(n3795), .B(n3796), .Z(n3625) );
  AND U3405 ( .A(n133), .B(n3797), .Z(n3796) );
  XOR U3406 ( .A(p_input[3803]), .B(p_input[3787]), .Z(n3797) );
  XOR U3407 ( .A(n3798), .B(n3799), .Z(n3789) );
  AND U3408 ( .A(n3800), .B(n3801), .Z(n3799) );
  XOR U3409 ( .A(n3798), .B(n3640), .Z(n3801) );
  XNOR U3410 ( .A(p_input[3818]), .B(n3802), .Z(n3640) );
  AND U3411 ( .A(n135), .B(n3803), .Z(n3802) );
  XOR U3412 ( .A(p_input[3834]), .B(p_input[3818]), .Z(n3803) );
  XNOR U3413 ( .A(n3637), .B(n3798), .Z(n3800) );
  XOR U3414 ( .A(n3804), .B(n3805), .Z(n3637) );
  AND U3415 ( .A(n133), .B(n3806), .Z(n3805) );
  XOR U3416 ( .A(p_input[3802]), .B(p_input[3786]), .Z(n3806) );
  XOR U3417 ( .A(n3807), .B(n3808), .Z(n3798) );
  AND U3418 ( .A(n3809), .B(n3810), .Z(n3808) );
  XOR U3419 ( .A(n3807), .B(n3652), .Z(n3810) );
  XNOR U3420 ( .A(p_input[3817]), .B(n3811), .Z(n3652) );
  AND U3421 ( .A(n135), .B(n3812), .Z(n3811) );
  XOR U3422 ( .A(p_input[3833]), .B(p_input[3817]), .Z(n3812) );
  XNOR U3423 ( .A(n3649), .B(n3807), .Z(n3809) );
  XOR U3424 ( .A(n3813), .B(n3814), .Z(n3649) );
  AND U3425 ( .A(n133), .B(n3815), .Z(n3814) );
  XOR U3426 ( .A(p_input[3801]), .B(p_input[3785]), .Z(n3815) );
  XOR U3427 ( .A(n3816), .B(n3817), .Z(n3807) );
  AND U3428 ( .A(n3818), .B(n3819), .Z(n3817) );
  XOR U3429 ( .A(n3816), .B(n3664), .Z(n3819) );
  XNOR U3430 ( .A(p_input[3816]), .B(n3820), .Z(n3664) );
  AND U3431 ( .A(n135), .B(n3821), .Z(n3820) );
  XOR U3432 ( .A(p_input[3832]), .B(p_input[3816]), .Z(n3821) );
  XNOR U3433 ( .A(n3661), .B(n3816), .Z(n3818) );
  XOR U3434 ( .A(n3822), .B(n3823), .Z(n3661) );
  AND U3435 ( .A(n133), .B(n3824), .Z(n3823) );
  XOR U3436 ( .A(p_input[3800]), .B(p_input[3784]), .Z(n3824) );
  XOR U3437 ( .A(n3825), .B(n3826), .Z(n3816) );
  AND U3438 ( .A(n3827), .B(n3828), .Z(n3826) );
  XOR U3439 ( .A(n3825), .B(n3676), .Z(n3828) );
  XNOR U3440 ( .A(p_input[3815]), .B(n3829), .Z(n3676) );
  AND U3441 ( .A(n135), .B(n3830), .Z(n3829) );
  XOR U3442 ( .A(p_input[3831]), .B(p_input[3815]), .Z(n3830) );
  XNOR U3443 ( .A(n3673), .B(n3825), .Z(n3827) );
  XOR U3444 ( .A(n3831), .B(n3832), .Z(n3673) );
  AND U3445 ( .A(n133), .B(n3833), .Z(n3832) );
  XOR U3446 ( .A(p_input[3799]), .B(p_input[3783]), .Z(n3833) );
  XOR U3447 ( .A(n3834), .B(n3835), .Z(n3825) );
  AND U3448 ( .A(n3836), .B(n3837), .Z(n3835) );
  XOR U3449 ( .A(n3834), .B(n3688), .Z(n3837) );
  XNOR U3450 ( .A(p_input[3814]), .B(n3838), .Z(n3688) );
  AND U3451 ( .A(n135), .B(n3839), .Z(n3838) );
  XOR U3452 ( .A(p_input[3830]), .B(p_input[3814]), .Z(n3839) );
  XNOR U3453 ( .A(n3685), .B(n3834), .Z(n3836) );
  XOR U3454 ( .A(n3840), .B(n3841), .Z(n3685) );
  AND U3455 ( .A(n133), .B(n3842), .Z(n3841) );
  XOR U3456 ( .A(p_input[3798]), .B(p_input[3782]), .Z(n3842) );
  XOR U3457 ( .A(n3843), .B(n3844), .Z(n3834) );
  AND U3458 ( .A(n3845), .B(n3846), .Z(n3844) );
  XOR U3459 ( .A(n3843), .B(n3700), .Z(n3846) );
  XNOR U3460 ( .A(p_input[3813]), .B(n3847), .Z(n3700) );
  AND U3461 ( .A(n135), .B(n3848), .Z(n3847) );
  XOR U3462 ( .A(p_input[3829]), .B(p_input[3813]), .Z(n3848) );
  XNOR U3463 ( .A(n3697), .B(n3843), .Z(n3845) );
  XOR U3464 ( .A(n3849), .B(n3850), .Z(n3697) );
  AND U3465 ( .A(n133), .B(n3851), .Z(n3850) );
  XOR U3466 ( .A(p_input[3797]), .B(p_input[3781]), .Z(n3851) );
  XOR U3467 ( .A(n3852), .B(n3853), .Z(n3843) );
  AND U3468 ( .A(n3854), .B(n3855), .Z(n3853) );
  XOR U3469 ( .A(n3852), .B(n3712), .Z(n3855) );
  XNOR U3470 ( .A(p_input[3812]), .B(n3856), .Z(n3712) );
  AND U3471 ( .A(n135), .B(n3857), .Z(n3856) );
  XOR U3472 ( .A(p_input[3828]), .B(p_input[3812]), .Z(n3857) );
  XNOR U3473 ( .A(n3709), .B(n3852), .Z(n3854) );
  XOR U3474 ( .A(n3858), .B(n3859), .Z(n3709) );
  AND U3475 ( .A(n133), .B(n3860), .Z(n3859) );
  XOR U3476 ( .A(p_input[3796]), .B(p_input[3780]), .Z(n3860) );
  XOR U3477 ( .A(n3861), .B(n3862), .Z(n3852) );
  AND U3478 ( .A(n3863), .B(n3864), .Z(n3862) );
  XOR U3479 ( .A(n3861), .B(n3724), .Z(n3864) );
  XNOR U3480 ( .A(p_input[3811]), .B(n3865), .Z(n3724) );
  AND U3481 ( .A(n135), .B(n3866), .Z(n3865) );
  XOR U3482 ( .A(p_input[3827]), .B(p_input[3811]), .Z(n3866) );
  XNOR U3483 ( .A(n3721), .B(n3861), .Z(n3863) );
  XOR U3484 ( .A(n3867), .B(n3868), .Z(n3721) );
  AND U3485 ( .A(n133), .B(n3869), .Z(n3868) );
  XOR U3486 ( .A(p_input[3795]), .B(p_input[3779]), .Z(n3869) );
  XOR U3487 ( .A(n3870), .B(n3871), .Z(n3861) );
  AND U3488 ( .A(n3872), .B(n3873), .Z(n3871) );
  XOR U3489 ( .A(n3870), .B(n3736), .Z(n3873) );
  XNOR U3490 ( .A(p_input[3810]), .B(n3874), .Z(n3736) );
  AND U3491 ( .A(n135), .B(n3875), .Z(n3874) );
  XOR U3492 ( .A(p_input[3826]), .B(p_input[3810]), .Z(n3875) );
  XNOR U3493 ( .A(n3733), .B(n3870), .Z(n3872) );
  XOR U3494 ( .A(n3876), .B(n3877), .Z(n3733) );
  AND U3495 ( .A(n133), .B(n3878), .Z(n3877) );
  XOR U3496 ( .A(p_input[3794]), .B(p_input[3778]), .Z(n3878) );
  XOR U3497 ( .A(n3879), .B(n3880), .Z(n3870) );
  AND U3498 ( .A(n3881), .B(n3882), .Z(n3880) );
  XNOR U3499 ( .A(n3883), .B(n3749), .Z(n3882) );
  XNOR U3500 ( .A(p_input[3809]), .B(n3884), .Z(n3749) );
  AND U3501 ( .A(n135), .B(n3885), .Z(n3884) );
  XNOR U3502 ( .A(p_input[3825]), .B(n3886), .Z(n3885) );
  IV U3503 ( .A(p_input[3809]), .Z(n3886) );
  XNOR U3504 ( .A(n3746), .B(n3879), .Z(n3881) );
  XNOR U3505 ( .A(p_input[3777]), .B(n3887), .Z(n3746) );
  AND U3506 ( .A(n133), .B(n3888), .Z(n3887) );
  XOR U3507 ( .A(p_input[3793]), .B(p_input[3777]), .Z(n3888) );
  IV U3508 ( .A(n3883), .Z(n3879) );
  AND U3509 ( .A(n3754), .B(n3757), .Z(n3883) );
  XOR U3510 ( .A(p_input[3808]), .B(n3889), .Z(n3757) );
  AND U3511 ( .A(n135), .B(n3890), .Z(n3889) );
  XOR U3512 ( .A(p_input[3824]), .B(p_input[3808]), .Z(n3890) );
  XOR U3513 ( .A(n3891), .B(n3892), .Z(n135) );
  AND U3514 ( .A(n3893), .B(n3894), .Z(n3892) );
  XNOR U3515 ( .A(p_input[3839]), .B(n3891), .Z(n3894) );
  XOR U3516 ( .A(n3891), .B(p_input[3823]), .Z(n3893) );
  XOR U3517 ( .A(n3895), .B(n3896), .Z(n3891) );
  AND U3518 ( .A(n3897), .B(n3898), .Z(n3896) );
  XNOR U3519 ( .A(p_input[3838]), .B(n3895), .Z(n3898) );
  XOR U3520 ( .A(n3895), .B(p_input[3822]), .Z(n3897) );
  XOR U3521 ( .A(n3899), .B(n3900), .Z(n3895) );
  AND U3522 ( .A(n3901), .B(n3902), .Z(n3900) );
  XNOR U3523 ( .A(p_input[3837]), .B(n3899), .Z(n3902) );
  XOR U3524 ( .A(n3899), .B(p_input[3821]), .Z(n3901) );
  XOR U3525 ( .A(n3903), .B(n3904), .Z(n3899) );
  AND U3526 ( .A(n3905), .B(n3906), .Z(n3904) );
  XNOR U3527 ( .A(p_input[3836]), .B(n3903), .Z(n3906) );
  XOR U3528 ( .A(n3903), .B(p_input[3820]), .Z(n3905) );
  XOR U3529 ( .A(n3907), .B(n3908), .Z(n3903) );
  AND U3530 ( .A(n3909), .B(n3910), .Z(n3908) );
  XNOR U3531 ( .A(p_input[3835]), .B(n3907), .Z(n3910) );
  XOR U3532 ( .A(n3907), .B(p_input[3819]), .Z(n3909) );
  XOR U3533 ( .A(n3911), .B(n3912), .Z(n3907) );
  AND U3534 ( .A(n3913), .B(n3914), .Z(n3912) );
  XNOR U3535 ( .A(p_input[3834]), .B(n3911), .Z(n3914) );
  XOR U3536 ( .A(n3911), .B(p_input[3818]), .Z(n3913) );
  XOR U3537 ( .A(n3915), .B(n3916), .Z(n3911) );
  AND U3538 ( .A(n3917), .B(n3918), .Z(n3916) );
  XNOR U3539 ( .A(p_input[3833]), .B(n3915), .Z(n3918) );
  XOR U3540 ( .A(n3915), .B(p_input[3817]), .Z(n3917) );
  XOR U3541 ( .A(n3919), .B(n3920), .Z(n3915) );
  AND U3542 ( .A(n3921), .B(n3922), .Z(n3920) );
  XNOR U3543 ( .A(p_input[3832]), .B(n3919), .Z(n3922) );
  XOR U3544 ( .A(n3919), .B(p_input[3816]), .Z(n3921) );
  XOR U3545 ( .A(n3923), .B(n3924), .Z(n3919) );
  AND U3546 ( .A(n3925), .B(n3926), .Z(n3924) );
  XNOR U3547 ( .A(p_input[3831]), .B(n3923), .Z(n3926) );
  XOR U3548 ( .A(n3923), .B(p_input[3815]), .Z(n3925) );
  XOR U3549 ( .A(n3927), .B(n3928), .Z(n3923) );
  AND U3550 ( .A(n3929), .B(n3930), .Z(n3928) );
  XNOR U3551 ( .A(p_input[3830]), .B(n3927), .Z(n3930) );
  XOR U3552 ( .A(n3927), .B(p_input[3814]), .Z(n3929) );
  XOR U3553 ( .A(n3931), .B(n3932), .Z(n3927) );
  AND U3554 ( .A(n3933), .B(n3934), .Z(n3932) );
  XNOR U3555 ( .A(p_input[3829]), .B(n3931), .Z(n3934) );
  XOR U3556 ( .A(n3931), .B(p_input[3813]), .Z(n3933) );
  XOR U3557 ( .A(n3935), .B(n3936), .Z(n3931) );
  AND U3558 ( .A(n3937), .B(n3938), .Z(n3936) );
  XNOR U3559 ( .A(p_input[3828]), .B(n3935), .Z(n3938) );
  XOR U3560 ( .A(n3935), .B(p_input[3812]), .Z(n3937) );
  XOR U3561 ( .A(n3939), .B(n3940), .Z(n3935) );
  AND U3562 ( .A(n3941), .B(n3942), .Z(n3940) );
  XNOR U3563 ( .A(p_input[3827]), .B(n3939), .Z(n3942) );
  XOR U3564 ( .A(n3939), .B(p_input[3811]), .Z(n3941) );
  XOR U3565 ( .A(n3943), .B(n3944), .Z(n3939) );
  AND U3566 ( .A(n3945), .B(n3946), .Z(n3944) );
  XNOR U3567 ( .A(p_input[3826]), .B(n3943), .Z(n3946) );
  XOR U3568 ( .A(n3943), .B(p_input[3810]), .Z(n3945) );
  XNOR U3569 ( .A(n3947), .B(n3948), .Z(n3943) );
  AND U3570 ( .A(n3949), .B(n3950), .Z(n3948) );
  XOR U3571 ( .A(p_input[3825]), .B(n3947), .Z(n3950) );
  XNOR U3572 ( .A(p_input[3809]), .B(n3947), .Z(n3949) );
  AND U3573 ( .A(p_input[3824]), .B(n3951), .Z(n3947) );
  IV U3574 ( .A(p_input[3808]), .Z(n3951) );
  XNOR U3575 ( .A(p_input[3776]), .B(n3952), .Z(n3754) );
  AND U3576 ( .A(n133), .B(n3953), .Z(n3952) );
  XOR U3577 ( .A(p_input[3792]), .B(p_input[3776]), .Z(n3953) );
  XOR U3578 ( .A(n3954), .B(n3955), .Z(n133) );
  AND U3579 ( .A(n3956), .B(n3957), .Z(n3955) );
  XNOR U3580 ( .A(p_input[3807]), .B(n3954), .Z(n3957) );
  XOR U3581 ( .A(n3954), .B(p_input[3791]), .Z(n3956) );
  XOR U3582 ( .A(n3958), .B(n3959), .Z(n3954) );
  AND U3583 ( .A(n3960), .B(n3961), .Z(n3959) );
  XNOR U3584 ( .A(p_input[3806]), .B(n3958), .Z(n3961) );
  XNOR U3585 ( .A(n3958), .B(n3768), .Z(n3960) );
  IV U3586 ( .A(p_input[3790]), .Z(n3768) );
  XOR U3587 ( .A(n3962), .B(n3963), .Z(n3958) );
  AND U3588 ( .A(n3964), .B(n3965), .Z(n3963) );
  XNOR U3589 ( .A(p_input[3805]), .B(n3962), .Z(n3965) );
  XNOR U3590 ( .A(n3962), .B(n3777), .Z(n3964) );
  IV U3591 ( .A(p_input[3789]), .Z(n3777) );
  XOR U3592 ( .A(n3966), .B(n3967), .Z(n3962) );
  AND U3593 ( .A(n3968), .B(n3969), .Z(n3967) );
  XNOR U3594 ( .A(p_input[3804]), .B(n3966), .Z(n3969) );
  XNOR U3595 ( .A(n3966), .B(n3786), .Z(n3968) );
  IV U3596 ( .A(p_input[3788]), .Z(n3786) );
  XOR U3597 ( .A(n3970), .B(n3971), .Z(n3966) );
  AND U3598 ( .A(n3972), .B(n3973), .Z(n3971) );
  XNOR U3599 ( .A(p_input[3803]), .B(n3970), .Z(n3973) );
  XNOR U3600 ( .A(n3970), .B(n3795), .Z(n3972) );
  IV U3601 ( .A(p_input[3787]), .Z(n3795) );
  XOR U3602 ( .A(n3974), .B(n3975), .Z(n3970) );
  AND U3603 ( .A(n3976), .B(n3977), .Z(n3975) );
  XNOR U3604 ( .A(p_input[3802]), .B(n3974), .Z(n3977) );
  XNOR U3605 ( .A(n3974), .B(n3804), .Z(n3976) );
  IV U3606 ( .A(p_input[3786]), .Z(n3804) );
  XOR U3607 ( .A(n3978), .B(n3979), .Z(n3974) );
  AND U3608 ( .A(n3980), .B(n3981), .Z(n3979) );
  XNOR U3609 ( .A(p_input[3801]), .B(n3978), .Z(n3981) );
  XNOR U3610 ( .A(n3978), .B(n3813), .Z(n3980) );
  IV U3611 ( .A(p_input[3785]), .Z(n3813) );
  XOR U3612 ( .A(n3982), .B(n3983), .Z(n3978) );
  AND U3613 ( .A(n3984), .B(n3985), .Z(n3983) );
  XNOR U3614 ( .A(p_input[3800]), .B(n3982), .Z(n3985) );
  XNOR U3615 ( .A(n3982), .B(n3822), .Z(n3984) );
  IV U3616 ( .A(p_input[3784]), .Z(n3822) );
  XOR U3617 ( .A(n3986), .B(n3987), .Z(n3982) );
  AND U3618 ( .A(n3988), .B(n3989), .Z(n3987) );
  XNOR U3619 ( .A(p_input[3799]), .B(n3986), .Z(n3989) );
  XNOR U3620 ( .A(n3986), .B(n3831), .Z(n3988) );
  IV U3621 ( .A(p_input[3783]), .Z(n3831) );
  XOR U3622 ( .A(n3990), .B(n3991), .Z(n3986) );
  AND U3623 ( .A(n3992), .B(n3993), .Z(n3991) );
  XNOR U3624 ( .A(p_input[3798]), .B(n3990), .Z(n3993) );
  XNOR U3625 ( .A(n3990), .B(n3840), .Z(n3992) );
  IV U3626 ( .A(p_input[3782]), .Z(n3840) );
  XOR U3627 ( .A(n3994), .B(n3995), .Z(n3990) );
  AND U3628 ( .A(n3996), .B(n3997), .Z(n3995) );
  XNOR U3629 ( .A(p_input[3797]), .B(n3994), .Z(n3997) );
  XNOR U3630 ( .A(n3994), .B(n3849), .Z(n3996) );
  IV U3631 ( .A(p_input[3781]), .Z(n3849) );
  XOR U3632 ( .A(n3998), .B(n3999), .Z(n3994) );
  AND U3633 ( .A(n4000), .B(n4001), .Z(n3999) );
  XNOR U3634 ( .A(p_input[3796]), .B(n3998), .Z(n4001) );
  XNOR U3635 ( .A(n3998), .B(n3858), .Z(n4000) );
  IV U3636 ( .A(p_input[3780]), .Z(n3858) );
  XOR U3637 ( .A(n4002), .B(n4003), .Z(n3998) );
  AND U3638 ( .A(n4004), .B(n4005), .Z(n4003) );
  XNOR U3639 ( .A(p_input[3795]), .B(n4002), .Z(n4005) );
  XNOR U3640 ( .A(n4002), .B(n3867), .Z(n4004) );
  IV U3641 ( .A(p_input[3779]), .Z(n3867) );
  XOR U3642 ( .A(n4006), .B(n4007), .Z(n4002) );
  AND U3643 ( .A(n4008), .B(n4009), .Z(n4007) );
  XNOR U3644 ( .A(p_input[3794]), .B(n4006), .Z(n4009) );
  XNOR U3645 ( .A(n4006), .B(n3876), .Z(n4008) );
  IV U3646 ( .A(p_input[3778]), .Z(n3876) );
  XNOR U3647 ( .A(n4010), .B(n4011), .Z(n4006) );
  AND U3648 ( .A(n4012), .B(n4013), .Z(n4011) );
  XOR U3649 ( .A(p_input[3793]), .B(n4010), .Z(n4013) );
  XNOR U3650 ( .A(p_input[3777]), .B(n4010), .Z(n4012) );
  AND U3651 ( .A(p_input[3792]), .B(n4014), .Z(n4010) );
  IV U3652 ( .A(p_input[3776]), .Z(n4014) );
  XOR U3653 ( .A(n4015), .B(n4016), .Z(n3573) );
  AND U3654 ( .A(n369), .B(n4017), .Z(n4016) );
  XNOR U3655 ( .A(n4018), .B(n4015), .Z(n4017) );
  XOR U3656 ( .A(n4019), .B(n4020), .Z(n369) );
  AND U3657 ( .A(n4021), .B(n4022), .Z(n4020) );
  XNOR U3658 ( .A(n3583), .B(n4019), .Z(n4022) );
  AND U3659 ( .A(p_input[3775]), .B(p_input[3759]), .Z(n3583) );
  XOR U3660 ( .A(n4019), .B(n3584), .Z(n4021) );
  AND U3661 ( .A(p_input[3743]), .B(p_input[3727]), .Z(n3584) );
  XOR U3662 ( .A(n4023), .B(n4024), .Z(n4019) );
  AND U3663 ( .A(n4025), .B(n4026), .Z(n4024) );
  XOR U3664 ( .A(n4023), .B(n3596), .Z(n4026) );
  XNOR U3665 ( .A(p_input[3758]), .B(n4027), .Z(n3596) );
  AND U3666 ( .A(n139), .B(n4028), .Z(n4027) );
  XOR U3667 ( .A(p_input[3774]), .B(p_input[3758]), .Z(n4028) );
  XNOR U3668 ( .A(n3593), .B(n4023), .Z(n4025) );
  XOR U3669 ( .A(n4029), .B(n4030), .Z(n3593) );
  AND U3670 ( .A(n136), .B(n4031), .Z(n4030) );
  XOR U3671 ( .A(p_input[3742]), .B(p_input[3726]), .Z(n4031) );
  XOR U3672 ( .A(n4032), .B(n4033), .Z(n4023) );
  AND U3673 ( .A(n4034), .B(n4035), .Z(n4033) );
  XOR U3674 ( .A(n4032), .B(n3608), .Z(n4035) );
  XNOR U3675 ( .A(p_input[3757]), .B(n4036), .Z(n3608) );
  AND U3676 ( .A(n139), .B(n4037), .Z(n4036) );
  XOR U3677 ( .A(p_input[3773]), .B(p_input[3757]), .Z(n4037) );
  XNOR U3678 ( .A(n3605), .B(n4032), .Z(n4034) );
  XOR U3679 ( .A(n4038), .B(n4039), .Z(n3605) );
  AND U3680 ( .A(n136), .B(n4040), .Z(n4039) );
  XOR U3681 ( .A(p_input[3741]), .B(p_input[3725]), .Z(n4040) );
  XOR U3682 ( .A(n4041), .B(n4042), .Z(n4032) );
  AND U3683 ( .A(n4043), .B(n4044), .Z(n4042) );
  XOR U3684 ( .A(n4041), .B(n3620), .Z(n4044) );
  XNOR U3685 ( .A(p_input[3756]), .B(n4045), .Z(n3620) );
  AND U3686 ( .A(n139), .B(n4046), .Z(n4045) );
  XOR U3687 ( .A(p_input[3772]), .B(p_input[3756]), .Z(n4046) );
  XNOR U3688 ( .A(n3617), .B(n4041), .Z(n4043) );
  XOR U3689 ( .A(n4047), .B(n4048), .Z(n3617) );
  AND U3690 ( .A(n136), .B(n4049), .Z(n4048) );
  XOR U3691 ( .A(p_input[3740]), .B(p_input[3724]), .Z(n4049) );
  XOR U3692 ( .A(n4050), .B(n4051), .Z(n4041) );
  AND U3693 ( .A(n4052), .B(n4053), .Z(n4051) );
  XOR U3694 ( .A(n4050), .B(n3632), .Z(n4053) );
  XNOR U3695 ( .A(p_input[3755]), .B(n4054), .Z(n3632) );
  AND U3696 ( .A(n139), .B(n4055), .Z(n4054) );
  XOR U3697 ( .A(p_input[3771]), .B(p_input[3755]), .Z(n4055) );
  XNOR U3698 ( .A(n3629), .B(n4050), .Z(n4052) );
  XOR U3699 ( .A(n4056), .B(n4057), .Z(n3629) );
  AND U3700 ( .A(n136), .B(n4058), .Z(n4057) );
  XOR U3701 ( .A(p_input[3739]), .B(p_input[3723]), .Z(n4058) );
  XOR U3702 ( .A(n4059), .B(n4060), .Z(n4050) );
  AND U3703 ( .A(n4061), .B(n4062), .Z(n4060) );
  XOR U3704 ( .A(n4059), .B(n3644), .Z(n4062) );
  XNOR U3705 ( .A(p_input[3754]), .B(n4063), .Z(n3644) );
  AND U3706 ( .A(n139), .B(n4064), .Z(n4063) );
  XOR U3707 ( .A(p_input[3770]), .B(p_input[3754]), .Z(n4064) );
  XNOR U3708 ( .A(n3641), .B(n4059), .Z(n4061) );
  XOR U3709 ( .A(n4065), .B(n4066), .Z(n3641) );
  AND U3710 ( .A(n136), .B(n4067), .Z(n4066) );
  XOR U3711 ( .A(p_input[3738]), .B(p_input[3722]), .Z(n4067) );
  XOR U3712 ( .A(n4068), .B(n4069), .Z(n4059) );
  AND U3713 ( .A(n4070), .B(n4071), .Z(n4069) );
  XOR U3714 ( .A(n4068), .B(n3656), .Z(n4071) );
  XNOR U3715 ( .A(p_input[3753]), .B(n4072), .Z(n3656) );
  AND U3716 ( .A(n139), .B(n4073), .Z(n4072) );
  XOR U3717 ( .A(p_input[3769]), .B(p_input[3753]), .Z(n4073) );
  XNOR U3718 ( .A(n3653), .B(n4068), .Z(n4070) );
  XOR U3719 ( .A(n4074), .B(n4075), .Z(n3653) );
  AND U3720 ( .A(n136), .B(n4076), .Z(n4075) );
  XOR U3721 ( .A(p_input[3737]), .B(p_input[3721]), .Z(n4076) );
  XOR U3722 ( .A(n4077), .B(n4078), .Z(n4068) );
  AND U3723 ( .A(n4079), .B(n4080), .Z(n4078) );
  XOR U3724 ( .A(n4077), .B(n3668), .Z(n4080) );
  XNOR U3725 ( .A(p_input[3752]), .B(n4081), .Z(n3668) );
  AND U3726 ( .A(n139), .B(n4082), .Z(n4081) );
  XOR U3727 ( .A(p_input[3768]), .B(p_input[3752]), .Z(n4082) );
  XNOR U3728 ( .A(n3665), .B(n4077), .Z(n4079) );
  XOR U3729 ( .A(n4083), .B(n4084), .Z(n3665) );
  AND U3730 ( .A(n136), .B(n4085), .Z(n4084) );
  XOR U3731 ( .A(p_input[3736]), .B(p_input[3720]), .Z(n4085) );
  XOR U3732 ( .A(n4086), .B(n4087), .Z(n4077) );
  AND U3733 ( .A(n4088), .B(n4089), .Z(n4087) );
  XOR U3734 ( .A(n4086), .B(n3680), .Z(n4089) );
  XNOR U3735 ( .A(p_input[3751]), .B(n4090), .Z(n3680) );
  AND U3736 ( .A(n139), .B(n4091), .Z(n4090) );
  XOR U3737 ( .A(p_input[3767]), .B(p_input[3751]), .Z(n4091) );
  XNOR U3738 ( .A(n3677), .B(n4086), .Z(n4088) );
  XOR U3739 ( .A(n4092), .B(n4093), .Z(n3677) );
  AND U3740 ( .A(n136), .B(n4094), .Z(n4093) );
  XOR U3741 ( .A(p_input[3735]), .B(p_input[3719]), .Z(n4094) );
  XOR U3742 ( .A(n4095), .B(n4096), .Z(n4086) );
  AND U3743 ( .A(n4097), .B(n4098), .Z(n4096) );
  XOR U3744 ( .A(n4095), .B(n3692), .Z(n4098) );
  XNOR U3745 ( .A(p_input[3750]), .B(n4099), .Z(n3692) );
  AND U3746 ( .A(n139), .B(n4100), .Z(n4099) );
  XOR U3747 ( .A(p_input[3766]), .B(p_input[3750]), .Z(n4100) );
  XNOR U3748 ( .A(n3689), .B(n4095), .Z(n4097) );
  XOR U3749 ( .A(n4101), .B(n4102), .Z(n3689) );
  AND U3750 ( .A(n136), .B(n4103), .Z(n4102) );
  XOR U3751 ( .A(p_input[3734]), .B(p_input[3718]), .Z(n4103) );
  XOR U3752 ( .A(n4104), .B(n4105), .Z(n4095) );
  AND U3753 ( .A(n4106), .B(n4107), .Z(n4105) );
  XOR U3754 ( .A(n4104), .B(n3704), .Z(n4107) );
  XNOR U3755 ( .A(p_input[3749]), .B(n4108), .Z(n3704) );
  AND U3756 ( .A(n139), .B(n4109), .Z(n4108) );
  XOR U3757 ( .A(p_input[3765]), .B(p_input[3749]), .Z(n4109) );
  XNOR U3758 ( .A(n3701), .B(n4104), .Z(n4106) );
  XOR U3759 ( .A(n4110), .B(n4111), .Z(n3701) );
  AND U3760 ( .A(n136), .B(n4112), .Z(n4111) );
  XOR U3761 ( .A(p_input[3733]), .B(p_input[3717]), .Z(n4112) );
  XOR U3762 ( .A(n4113), .B(n4114), .Z(n4104) );
  AND U3763 ( .A(n4115), .B(n4116), .Z(n4114) );
  XOR U3764 ( .A(n4113), .B(n3716), .Z(n4116) );
  XNOR U3765 ( .A(p_input[3748]), .B(n4117), .Z(n3716) );
  AND U3766 ( .A(n139), .B(n4118), .Z(n4117) );
  XOR U3767 ( .A(p_input[3764]), .B(p_input[3748]), .Z(n4118) );
  XNOR U3768 ( .A(n3713), .B(n4113), .Z(n4115) );
  XOR U3769 ( .A(n4119), .B(n4120), .Z(n3713) );
  AND U3770 ( .A(n136), .B(n4121), .Z(n4120) );
  XOR U3771 ( .A(p_input[3732]), .B(p_input[3716]), .Z(n4121) );
  XOR U3772 ( .A(n4122), .B(n4123), .Z(n4113) );
  AND U3773 ( .A(n4124), .B(n4125), .Z(n4123) );
  XOR U3774 ( .A(n4122), .B(n3728), .Z(n4125) );
  XNOR U3775 ( .A(p_input[3747]), .B(n4126), .Z(n3728) );
  AND U3776 ( .A(n139), .B(n4127), .Z(n4126) );
  XOR U3777 ( .A(p_input[3763]), .B(p_input[3747]), .Z(n4127) );
  XNOR U3778 ( .A(n3725), .B(n4122), .Z(n4124) );
  XOR U3779 ( .A(n4128), .B(n4129), .Z(n3725) );
  AND U3780 ( .A(n136), .B(n4130), .Z(n4129) );
  XOR U3781 ( .A(p_input[3731]), .B(p_input[3715]), .Z(n4130) );
  XOR U3782 ( .A(n4131), .B(n4132), .Z(n4122) );
  AND U3783 ( .A(n4133), .B(n4134), .Z(n4132) );
  XOR U3784 ( .A(n4131), .B(n3740), .Z(n4134) );
  XNOR U3785 ( .A(p_input[3746]), .B(n4135), .Z(n3740) );
  AND U3786 ( .A(n139), .B(n4136), .Z(n4135) );
  XOR U3787 ( .A(p_input[3762]), .B(p_input[3746]), .Z(n4136) );
  XNOR U3788 ( .A(n3737), .B(n4131), .Z(n4133) );
  XOR U3789 ( .A(n4137), .B(n4138), .Z(n3737) );
  AND U3790 ( .A(n136), .B(n4139), .Z(n4138) );
  XOR U3791 ( .A(p_input[3730]), .B(p_input[3714]), .Z(n4139) );
  XOR U3792 ( .A(n4140), .B(n4141), .Z(n4131) );
  AND U3793 ( .A(n4142), .B(n4143), .Z(n4141) );
  XNOR U3794 ( .A(n4144), .B(n3753), .Z(n4143) );
  XNOR U3795 ( .A(p_input[3745]), .B(n4145), .Z(n3753) );
  AND U3796 ( .A(n139), .B(n4146), .Z(n4145) );
  XNOR U3797 ( .A(p_input[3761]), .B(n4147), .Z(n4146) );
  IV U3798 ( .A(p_input[3745]), .Z(n4147) );
  XNOR U3799 ( .A(n3750), .B(n4140), .Z(n4142) );
  XNOR U3800 ( .A(p_input[3713]), .B(n4148), .Z(n3750) );
  AND U3801 ( .A(n136), .B(n4149), .Z(n4148) );
  XOR U3802 ( .A(p_input[3729]), .B(p_input[3713]), .Z(n4149) );
  IV U3803 ( .A(n4144), .Z(n4140) );
  AND U3804 ( .A(n4015), .B(n4018), .Z(n4144) );
  XOR U3805 ( .A(p_input[3744]), .B(n4150), .Z(n4018) );
  AND U3806 ( .A(n139), .B(n4151), .Z(n4150) );
  XOR U3807 ( .A(p_input[3760]), .B(p_input[3744]), .Z(n4151) );
  XOR U3808 ( .A(n4152), .B(n4153), .Z(n139) );
  AND U3809 ( .A(n4154), .B(n4155), .Z(n4153) );
  XNOR U3810 ( .A(p_input[3775]), .B(n4152), .Z(n4155) );
  XOR U3811 ( .A(n4152), .B(p_input[3759]), .Z(n4154) );
  XOR U3812 ( .A(n4156), .B(n4157), .Z(n4152) );
  AND U3813 ( .A(n4158), .B(n4159), .Z(n4157) );
  XNOR U3814 ( .A(p_input[3774]), .B(n4156), .Z(n4159) );
  XOR U3815 ( .A(n4156), .B(p_input[3758]), .Z(n4158) );
  XOR U3816 ( .A(n4160), .B(n4161), .Z(n4156) );
  AND U3817 ( .A(n4162), .B(n4163), .Z(n4161) );
  XNOR U3818 ( .A(p_input[3773]), .B(n4160), .Z(n4163) );
  XOR U3819 ( .A(n4160), .B(p_input[3757]), .Z(n4162) );
  XOR U3820 ( .A(n4164), .B(n4165), .Z(n4160) );
  AND U3821 ( .A(n4166), .B(n4167), .Z(n4165) );
  XNOR U3822 ( .A(p_input[3772]), .B(n4164), .Z(n4167) );
  XOR U3823 ( .A(n4164), .B(p_input[3756]), .Z(n4166) );
  XOR U3824 ( .A(n4168), .B(n4169), .Z(n4164) );
  AND U3825 ( .A(n4170), .B(n4171), .Z(n4169) );
  XNOR U3826 ( .A(p_input[3771]), .B(n4168), .Z(n4171) );
  XOR U3827 ( .A(n4168), .B(p_input[3755]), .Z(n4170) );
  XOR U3828 ( .A(n4172), .B(n4173), .Z(n4168) );
  AND U3829 ( .A(n4174), .B(n4175), .Z(n4173) );
  XNOR U3830 ( .A(p_input[3770]), .B(n4172), .Z(n4175) );
  XOR U3831 ( .A(n4172), .B(p_input[3754]), .Z(n4174) );
  XOR U3832 ( .A(n4176), .B(n4177), .Z(n4172) );
  AND U3833 ( .A(n4178), .B(n4179), .Z(n4177) );
  XNOR U3834 ( .A(p_input[3769]), .B(n4176), .Z(n4179) );
  XOR U3835 ( .A(n4176), .B(p_input[3753]), .Z(n4178) );
  XOR U3836 ( .A(n4180), .B(n4181), .Z(n4176) );
  AND U3837 ( .A(n4182), .B(n4183), .Z(n4181) );
  XNOR U3838 ( .A(p_input[3768]), .B(n4180), .Z(n4183) );
  XOR U3839 ( .A(n4180), .B(p_input[3752]), .Z(n4182) );
  XOR U3840 ( .A(n4184), .B(n4185), .Z(n4180) );
  AND U3841 ( .A(n4186), .B(n4187), .Z(n4185) );
  XNOR U3842 ( .A(p_input[3767]), .B(n4184), .Z(n4187) );
  XOR U3843 ( .A(n4184), .B(p_input[3751]), .Z(n4186) );
  XOR U3844 ( .A(n4188), .B(n4189), .Z(n4184) );
  AND U3845 ( .A(n4190), .B(n4191), .Z(n4189) );
  XNOR U3846 ( .A(p_input[3766]), .B(n4188), .Z(n4191) );
  XOR U3847 ( .A(n4188), .B(p_input[3750]), .Z(n4190) );
  XOR U3848 ( .A(n4192), .B(n4193), .Z(n4188) );
  AND U3849 ( .A(n4194), .B(n4195), .Z(n4193) );
  XNOR U3850 ( .A(p_input[3765]), .B(n4192), .Z(n4195) );
  XOR U3851 ( .A(n4192), .B(p_input[3749]), .Z(n4194) );
  XOR U3852 ( .A(n4196), .B(n4197), .Z(n4192) );
  AND U3853 ( .A(n4198), .B(n4199), .Z(n4197) );
  XNOR U3854 ( .A(p_input[3764]), .B(n4196), .Z(n4199) );
  XOR U3855 ( .A(n4196), .B(p_input[3748]), .Z(n4198) );
  XOR U3856 ( .A(n4200), .B(n4201), .Z(n4196) );
  AND U3857 ( .A(n4202), .B(n4203), .Z(n4201) );
  XNOR U3858 ( .A(p_input[3763]), .B(n4200), .Z(n4203) );
  XOR U3859 ( .A(n4200), .B(p_input[3747]), .Z(n4202) );
  XOR U3860 ( .A(n4204), .B(n4205), .Z(n4200) );
  AND U3861 ( .A(n4206), .B(n4207), .Z(n4205) );
  XNOR U3862 ( .A(p_input[3762]), .B(n4204), .Z(n4207) );
  XOR U3863 ( .A(n4204), .B(p_input[3746]), .Z(n4206) );
  XNOR U3864 ( .A(n4208), .B(n4209), .Z(n4204) );
  AND U3865 ( .A(n4210), .B(n4211), .Z(n4209) );
  XOR U3866 ( .A(p_input[3761]), .B(n4208), .Z(n4211) );
  XNOR U3867 ( .A(p_input[3745]), .B(n4208), .Z(n4210) );
  AND U3868 ( .A(p_input[3760]), .B(n4212), .Z(n4208) );
  IV U3869 ( .A(p_input[3744]), .Z(n4212) );
  XNOR U3870 ( .A(p_input[3712]), .B(n4213), .Z(n4015) );
  AND U3871 ( .A(n136), .B(n4214), .Z(n4213) );
  XOR U3872 ( .A(p_input[3728]), .B(p_input[3712]), .Z(n4214) );
  XOR U3873 ( .A(n4215), .B(n4216), .Z(n136) );
  AND U3874 ( .A(n4217), .B(n4218), .Z(n4216) );
  XNOR U3875 ( .A(p_input[3743]), .B(n4215), .Z(n4218) );
  XOR U3876 ( .A(n4215), .B(p_input[3727]), .Z(n4217) );
  XOR U3877 ( .A(n4219), .B(n4220), .Z(n4215) );
  AND U3878 ( .A(n4221), .B(n4222), .Z(n4220) );
  XNOR U3879 ( .A(p_input[3742]), .B(n4219), .Z(n4222) );
  XNOR U3880 ( .A(n4219), .B(n4029), .Z(n4221) );
  IV U3881 ( .A(p_input[3726]), .Z(n4029) );
  XOR U3882 ( .A(n4223), .B(n4224), .Z(n4219) );
  AND U3883 ( .A(n4225), .B(n4226), .Z(n4224) );
  XNOR U3884 ( .A(p_input[3741]), .B(n4223), .Z(n4226) );
  XNOR U3885 ( .A(n4223), .B(n4038), .Z(n4225) );
  IV U3886 ( .A(p_input[3725]), .Z(n4038) );
  XOR U3887 ( .A(n4227), .B(n4228), .Z(n4223) );
  AND U3888 ( .A(n4229), .B(n4230), .Z(n4228) );
  XNOR U3889 ( .A(p_input[3740]), .B(n4227), .Z(n4230) );
  XNOR U3890 ( .A(n4227), .B(n4047), .Z(n4229) );
  IV U3891 ( .A(p_input[3724]), .Z(n4047) );
  XOR U3892 ( .A(n4231), .B(n4232), .Z(n4227) );
  AND U3893 ( .A(n4233), .B(n4234), .Z(n4232) );
  XNOR U3894 ( .A(p_input[3739]), .B(n4231), .Z(n4234) );
  XNOR U3895 ( .A(n4231), .B(n4056), .Z(n4233) );
  IV U3896 ( .A(p_input[3723]), .Z(n4056) );
  XOR U3897 ( .A(n4235), .B(n4236), .Z(n4231) );
  AND U3898 ( .A(n4237), .B(n4238), .Z(n4236) );
  XNOR U3899 ( .A(p_input[3738]), .B(n4235), .Z(n4238) );
  XNOR U3900 ( .A(n4235), .B(n4065), .Z(n4237) );
  IV U3901 ( .A(p_input[3722]), .Z(n4065) );
  XOR U3902 ( .A(n4239), .B(n4240), .Z(n4235) );
  AND U3903 ( .A(n4241), .B(n4242), .Z(n4240) );
  XNOR U3904 ( .A(p_input[3737]), .B(n4239), .Z(n4242) );
  XNOR U3905 ( .A(n4239), .B(n4074), .Z(n4241) );
  IV U3906 ( .A(p_input[3721]), .Z(n4074) );
  XOR U3907 ( .A(n4243), .B(n4244), .Z(n4239) );
  AND U3908 ( .A(n4245), .B(n4246), .Z(n4244) );
  XNOR U3909 ( .A(p_input[3736]), .B(n4243), .Z(n4246) );
  XNOR U3910 ( .A(n4243), .B(n4083), .Z(n4245) );
  IV U3911 ( .A(p_input[3720]), .Z(n4083) );
  XOR U3912 ( .A(n4247), .B(n4248), .Z(n4243) );
  AND U3913 ( .A(n4249), .B(n4250), .Z(n4248) );
  XNOR U3914 ( .A(p_input[3735]), .B(n4247), .Z(n4250) );
  XNOR U3915 ( .A(n4247), .B(n4092), .Z(n4249) );
  IV U3916 ( .A(p_input[3719]), .Z(n4092) );
  XOR U3917 ( .A(n4251), .B(n4252), .Z(n4247) );
  AND U3918 ( .A(n4253), .B(n4254), .Z(n4252) );
  XNOR U3919 ( .A(p_input[3734]), .B(n4251), .Z(n4254) );
  XNOR U3920 ( .A(n4251), .B(n4101), .Z(n4253) );
  IV U3921 ( .A(p_input[3718]), .Z(n4101) );
  XOR U3922 ( .A(n4255), .B(n4256), .Z(n4251) );
  AND U3923 ( .A(n4257), .B(n4258), .Z(n4256) );
  XNOR U3924 ( .A(p_input[3733]), .B(n4255), .Z(n4258) );
  XNOR U3925 ( .A(n4255), .B(n4110), .Z(n4257) );
  IV U3926 ( .A(p_input[3717]), .Z(n4110) );
  XOR U3927 ( .A(n4259), .B(n4260), .Z(n4255) );
  AND U3928 ( .A(n4261), .B(n4262), .Z(n4260) );
  XNOR U3929 ( .A(p_input[3732]), .B(n4259), .Z(n4262) );
  XNOR U3930 ( .A(n4259), .B(n4119), .Z(n4261) );
  IV U3931 ( .A(p_input[3716]), .Z(n4119) );
  XOR U3932 ( .A(n4263), .B(n4264), .Z(n4259) );
  AND U3933 ( .A(n4265), .B(n4266), .Z(n4264) );
  XNOR U3934 ( .A(p_input[3731]), .B(n4263), .Z(n4266) );
  XNOR U3935 ( .A(n4263), .B(n4128), .Z(n4265) );
  IV U3936 ( .A(p_input[3715]), .Z(n4128) );
  XOR U3937 ( .A(n4267), .B(n4268), .Z(n4263) );
  AND U3938 ( .A(n4269), .B(n4270), .Z(n4268) );
  XNOR U3939 ( .A(p_input[3730]), .B(n4267), .Z(n4270) );
  XNOR U3940 ( .A(n4267), .B(n4137), .Z(n4269) );
  IV U3941 ( .A(p_input[3714]), .Z(n4137) );
  XNOR U3942 ( .A(n4271), .B(n4272), .Z(n4267) );
  AND U3943 ( .A(n4273), .B(n4274), .Z(n4272) );
  XOR U3944 ( .A(p_input[3729]), .B(n4271), .Z(n4274) );
  XNOR U3945 ( .A(p_input[3713]), .B(n4271), .Z(n4273) );
  AND U3946 ( .A(p_input[3728]), .B(n4275), .Z(n4271) );
  IV U3947 ( .A(p_input[3712]), .Z(n4275) );
  XOR U3948 ( .A(n4276), .B(n4277), .Z(n3391) );
  AND U3949 ( .A(n736), .B(n4278), .Z(n4277) );
  XNOR U3950 ( .A(n4279), .B(n4276), .Z(n4278) );
  XOR U3951 ( .A(n4280), .B(n4281), .Z(n736) );
  AND U3952 ( .A(n4282), .B(n4283), .Z(n4281) );
  XNOR U3953 ( .A(n3403), .B(n4280), .Z(n4283) );
  AND U3954 ( .A(n4284), .B(n4285), .Z(n3403) );
  XOR U3955 ( .A(n4280), .B(n3402), .Z(n4282) );
  AND U3956 ( .A(n4286), .B(n4287), .Z(n3402) );
  XOR U3957 ( .A(n4288), .B(n4289), .Z(n4280) );
  AND U3958 ( .A(n4290), .B(n4291), .Z(n4289) );
  XOR U3959 ( .A(n4288), .B(n3415), .Z(n4291) );
  XOR U3960 ( .A(n4292), .B(n4293), .Z(n3415) );
  AND U3961 ( .A(n375), .B(n4294), .Z(n4293) );
  XOR U3962 ( .A(n4295), .B(n4292), .Z(n4294) );
  XNOR U3963 ( .A(n3412), .B(n4288), .Z(n4290) );
  XOR U3964 ( .A(n4296), .B(n4297), .Z(n3412) );
  AND U3965 ( .A(n372), .B(n4298), .Z(n4297) );
  XOR U3966 ( .A(n4299), .B(n4296), .Z(n4298) );
  XOR U3967 ( .A(n4300), .B(n4301), .Z(n4288) );
  AND U3968 ( .A(n4302), .B(n4303), .Z(n4301) );
  XOR U3969 ( .A(n4300), .B(n3427), .Z(n4303) );
  XOR U3970 ( .A(n4304), .B(n4305), .Z(n3427) );
  AND U3971 ( .A(n375), .B(n4306), .Z(n4305) );
  XOR U3972 ( .A(n4307), .B(n4304), .Z(n4306) );
  XNOR U3973 ( .A(n3424), .B(n4300), .Z(n4302) );
  XOR U3974 ( .A(n4308), .B(n4309), .Z(n3424) );
  AND U3975 ( .A(n372), .B(n4310), .Z(n4309) );
  XOR U3976 ( .A(n4311), .B(n4308), .Z(n4310) );
  XOR U3977 ( .A(n4312), .B(n4313), .Z(n4300) );
  AND U3978 ( .A(n4314), .B(n4315), .Z(n4313) );
  XOR U3979 ( .A(n4312), .B(n3439), .Z(n4315) );
  XOR U3980 ( .A(n4316), .B(n4317), .Z(n3439) );
  AND U3981 ( .A(n375), .B(n4318), .Z(n4317) );
  XOR U3982 ( .A(n4319), .B(n4316), .Z(n4318) );
  XNOR U3983 ( .A(n3436), .B(n4312), .Z(n4314) );
  XOR U3984 ( .A(n4320), .B(n4321), .Z(n3436) );
  AND U3985 ( .A(n372), .B(n4322), .Z(n4321) );
  XOR U3986 ( .A(n4323), .B(n4320), .Z(n4322) );
  XOR U3987 ( .A(n4324), .B(n4325), .Z(n4312) );
  AND U3988 ( .A(n4326), .B(n4327), .Z(n4325) );
  XOR U3989 ( .A(n4324), .B(n3451), .Z(n4327) );
  XOR U3990 ( .A(n4328), .B(n4329), .Z(n3451) );
  AND U3991 ( .A(n375), .B(n4330), .Z(n4329) );
  XOR U3992 ( .A(n4331), .B(n4328), .Z(n4330) );
  XNOR U3993 ( .A(n3448), .B(n4324), .Z(n4326) );
  XOR U3994 ( .A(n4332), .B(n4333), .Z(n3448) );
  AND U3995 ( .A(n372), .B(n4334), .Z(n4333) );
  XOR U3996 ( .A(n4335), .B(n4332), .Z(n4334) );
  XOR U3997 ( .A(n4336), .B(n4337), .Z(n4324) );
  AND U3998 ( .A(n4338), .B(n4339), .Z(n4337) );
  XOR U3999 ( .A(n4336), .B(n3463), .Z(n4339) );
  XOR U4000 ( .A(n4340), .B(n4341), .Z(n3463) );
  AND U4001 ( .A(n375), .B(n4342), .Z(n4341) );
  XOR U4002 ( .A(n4343), .B(n4340), .Z(n4342) );
  XNOR U4003 ( .A(n3460), .B(n4336), .Z(n4338) );
  XOR U4004 ( .A(n4344), .B(n4345), .Z(n3460) );
  AND U4005 ( .A(n372), .B(n4346), .Z(n4345) );
  XOR U4006 ( .A(n4347), .B(n4344), .Z(n4346) );
  XOR U4007 ( .A(n4348), .B(n4349), .Z(n4336) );
  AND U4008 ( .A(n4350), .B(n4351), .Z(n4349) );
  XOR U4009 ( .A(n4348), .B(n3475), .Z(n4351) );
  XOR U4010 ( .A(n4352), .B(n4353), .Z(n3475) );
  AND U4011 ( .A(n375), .B(n4354), .Z(n4353) );
  XOR U4012 ( .A(n4355), .B(n4352), .Z(n4354) );
  XNOR U4013 ( .A(n3472), .B(n4348), .Z(n4350) );
  XOR U4014 ( .A(n4356), .B(n4357), .Z(n3472) );
  AND U4015 ( .A(n372), .B(n4358), .Z(n4357) );
  XOR U4016 ( .A(n4359), .B(n4356), .Z(n4358) );
  XOR U4017 ( .A(n4360), .B(n4361), .Z(n4348) );
  AND U4018 ( .A(n4362), .B(n4363), .Z(n4361) );
  XOR U4019 ( .A(n4360), .B(n3487), .Z(n4363) );
  XOR U4020 ( .A(n4364), .B(n4365), .Z(n3487) );
  AND U4021 ( .A(n375), .B(n4366), .Z(n4365) );
  XOR U4022 ( .A(n4367), .B(n4364), .Z(n4366) );
  XNOR U4023 ( .A(n3484), .B(n4360), .Z(n4362) );
  XOR U4024 ( .A(n4368), .B(n4369), .Z(n3484) );
  AND U4025 ( .A(n372), .B(n4370), .Z(n4369) );
  XOR U4026 ( .A(n4371), .B(n4368), .Z(n4370) );
  XOR U4027 ( .A(n4372), .B(n4373), .Z(n4360) );
  AND U4028 ( .A(n4374), .B(n4375), .Z(n4373) );
  XOR U4029 ( .A(n4372), .B(n3499), .Z(n4375) );
  XOR U4030 ( .A(n4376), .B(n4377), .Z(n3499) );
  AND U4031 ( .A(n375), .B(n4378), .Z(n4377) );
  XOR U4032 ( .A(n4379), .B(n4376), .Z(n4378) );
  XNOR U4033 ( .A(n3496), .B(n4372), .Z(n4374) );
  XOR U4034 ( .A(n4380), .B(n4381), .Z(n3496) );
  AND U4035 ( .A(n372), .B(n4382), .Z(n4381) );
  XOR U4036 ( .A(n4383), .B(n4380), .Z(n4382) );
  XOR U4037 ( .A(n4384), .B(n4385), .Z(n4372) );
  AND U4038 ( .A(n4386), .B(n4387), .Z(n4385) );
  XOR U4039 ( .A(n4384), .B(n3511), .Z(n4387) );
  XOR U4040 ( .A(n4388), .B(n4389), .Z(n3511) );
  AND U4041 ( .A(n375), .B(n4390), .Z(n4389) );
  XOR U4042 ( .A(n4391), .B(n4388), .Z(n4390) );
  XNOR U4043 ( .A(n3508), .B(n4384), .Z(n4386) );
  XOR U4044 ( .A(n4392), .B(n4393), .Z(n3508) );
  AND U4045 ( .A(n372), .B(n4394), .Z(n4393) );
  XOR U4046 ( .A(n4395), .B(n4392), .Z(n4394) );
  XOR U4047 ( .A(n4396), .B(n4397), .Z(n4384) );
  AND U4048 ( .A(n4398), .B(n4399), .Z(n4397) );
  XOR U4049 ( .A(n4396), .B(n3523), .Z(n4399) );
  XOR U4050 ( .A(n4400), .B(n4401), .Z(n3523) );
  AND U4051 ( .A(n375), .B(n4402), .Z(n4401) );
  XOR U4052 ( .A(n4403), .B(n4400), .Z(n4402) );
  XNOR U4053 ( .A(n3520), .B(n4396), .Z(n4398) );
  XOR U4054 ( .A(n4404), .B(n4405), .Z(n3520) );
  AND U4055 ( .A(n372), .B(n4406), .Z(n4405) );
  XOR U4056 ( .A(n4407), .B(n4404), .Z(n4406) );
  XOR U4057 ( .A(n4408), .B(n4409), .Z(n4396) );
  AND U4058 ( .A(n4410), .B(n4411), .Z(n4409) );
  XOR U4059 ( .A(n4408), .B(n3535), .Z(n4411) );
  XOR U4060 ( .A(n4412), .B(n4413), .Z(n3535) );
  AND U4061 ( .A(n375), .B(n4414), .Z(n4413) );
  XOR U4062 ( .A(n4415), .B(n4412), .Z(n4414) );
  XNOR U4063 ( .A(n3532), .B(n4408), .Z(n4410) );
  XOR U4064 ( .A(n4416), .B(n4417), .Z(n3532) );
  AND U4065 ( .A(n372), .B(n4418), .Z(n4417) );
  XOR U4066 ( .A(n4419), .B(n4416), .Z(n4418) );
  XOR U4067 ( .A(n4420), .B(n4421), .Z(n4408) );
  AND U4068 ( .A(n4422), .B(n4423), .Z(n4421) );
  XOR U4069 ( .A(n4420), .B(n3547), .Z(n4423) );
  XOR U4070 ( .A(n4424), .B(n4425), .Z(n3547) );
  AND U4071 ( .A(n375), .B(n4426), .Z(n4425) );
  XOR U4072 ( .A(n4427), .B(n4424), .Z(n4426) );
  XNOR U4073 ( .A(n3544), .B(n4420), .Z(n4422) );
  XOR U4074 ( .A(n4428), .B(n4429), .Z(n3544) );
  AND U4075 ( .A(n372), .B(n4430), .Z(n4429) );
  XOR U4076 ( .A(n4431), .B(n4428), .Z(n4430) );
  XOR U4077 ( .A(n4432), .B(n4433), .Z(n4420) );
  AND U4078 ( .A(n4434), .B(n4435), .Z(n4433) );
  XOR U4079 ( .A(n4432), .B(n3559), .Z(n4435) );
  XOR U4080 ( .A(n4436), .B(n4437), .Z(n3559) );
  AND U4081 ( .A(n375), .B(n4438), .Z(n4437) );
  XOR U4082 ( .A(n4439), .B(n4436), .Z(n4438) );
  XNOR U4083 ( .A(n3556), .B(n4432), .Z(n4434) );
  XOR U4084 ( .A(n4440), .B(n4441), .Z(n3556) );
  AND U4085 ( .A(n372), .B(n4442), .Z(n4441) );
  XOR U4086 ( .A(n4443), .B(n4440), .Z(n4442) );
  XOR U4087 ( .A(n4444), .B(n4445), .Z(n4432) );
  AND U4088 ( .A(n4446), .B(n4447), .Z(n4445) );
  XNOR U4089 ( .A(n4448), .B(n3572), .Z(n4447) );
  XOR U4090 ( .A(n4449), .B(n4450), .Z(n3572) );
  AND U4091 ( .A(n375), .B(n4451), .Z(n4450) );
  XOR U4092 ( .A(n4449), .B(n4452), .Z(n4451) );
  XNOR U4093 ( .A(n3569), .B(n4444), .Z(n4446) );
  XOR U4094 ( .A(n4453), .B(n4454), .Z(n3569) );
  AND U4095 ( .A(n372), .B(n4455), .Z(n4454) );
  XOR U4096 ( .A(n4453), .B(n4456), .Z(n4455) );
  IV U4097 ( .A(n4448), .Z(n4444) );
  AND U4098 ( .A(n4276), .B(n4279), .Z(n4448) );
  XNOR U4099 ( .A(n4457), .B(n4458), .Z(n4279) );
  AND U4100 ( .A(n375), .B(n4459), .Z(n4458) );
  XNOR U4101 ( .A(n4460), .B(n4457), .Z(n4459) );
  XOR U4102 ( .A(n4461), .B(n4462), .Z(n375) );
  AND U4103 ( .A(n4463), .B(n4464), .Z(n4462) );
  XNOR U4104 ( .A(n4284), .B(n4461), .Z(n4464) );
  AND U4105 ( .A(p_input[3711]), .B(p_input[3695]), .Z(n4284) );
  XOR U4106 ( .A(n4461), .B(n4285), .Z(n4463) );
  AND U4107 ( .A(p_input[3679]), .B(p_input[3663]), .Z(n4285) );
  XOR U4108 ( .A(n4465), .B(n4466), .Z(n4461) );
  AND U4109 ( .A(n4467), .B(n4468), .Z(n4466) );
  XOR U4110 ( .A(n4465), .B(n4295), .Z(n4468) );
  XNOR U4111 ( .A(p_input[3694]), .B(n4469), .Z(n4295) );
  AND U4112 ( .A(n147), .B(n4470), .Z(n4469) );
  XOR U4113 ( .A(p_input[3710]), .B(p_input[3694]), .Z(n4470) );
  XNOR U4114 ( .A(n4292), .B(n4465), .Z(n4467) );
  XOR U4115 ( .A(n4471), .B(n4472), .Z(n4292) );
  AND U4116 ( .A(n145), .B(n4473), .Z(n4472) );
  XOR U4117 ( .A(p_input[3678]), .B(p_input[3662]), .Z(n4473) );
  XOR U4118 ( .A(n4474), .B(n4475), .Z(n4465) );
  AND U4119 ( .A(n4476), .B(n4477), .Z(n4475) );
  XOR U4120 ( .A(n4474), .B(n4307), .Z(n4477) );
  XNOR U4121 ( .A(p_input[3693]), .B(n4478), .Z(n4307) );
  AND U4122 ( .A(n147), .B(n4479), .Z(n4478) );
  XOR U4123 ( .A(p_input[3709]), .B(p_input[3693]), .Z(n4479) );
  XNOR U4124 ( .A(n4304), .B(n4474), .Z(n4476) );
  XOR U4125 ( .A(n4480), .B(n4481), .Z(n4304) );
  AND U4126 ( .A(n145), .B(n4482), .Z(n4481) );
  XOR U4127 ( .A(p_input[3677]), .B(p_input[3661]), .Z(n4482) );
  XOR U4128 ( .A(n4483), .B(n4484), .Z(n4474) );
  AND U4129 ( .A(n4485), .B(n4486), .Z(n4484) );
  XOR U4130 ( .A(n4483), .B(n4319), .Z(n4486) );
  XNOR U4131 ( .A(p_input[3692]), .B(n4487), .Z(n4319) );
  AND U4132 ( .A(n147), .B(n4488), .Z(n4487) );
  XOR U4133 ( .A(p_input[3708]), .B(p_input[3692]), .Z(n4488) );
  XNOR U4134 ( .A(n4316), .B(n4483), .Z(n4485) );
  XOR U4135 ( .A(n4489), .B(n4490), .Z(n4316) );
  AND U4136 ( .A(n145), .B(n4491), .Z(n4490) );
  XOR U4137 ( .A(p_input[3676]), .B(p_input[3660]), .Z(n4491) );
  XOR U4138 ( .A(n4492), .B(n4493), .Z(n4483) );
  AND U4139 ( .A(n4494), .B(n4495), .Z(n4493) );
  XOR U4140 ( .A(n4492), .B(n4331), .Z(n4495) );
  XNOR U4141 ( .A(p_input[3691]), .B(n4496), .Z(n4331) );
  AND U4142 ( .A(n147), .B(n4497), .Z(n4496) );
  XOR U4143 ( .A(p_input[3707]), .B(p_input[3691]), .Z(n4497) );
  XNOR U4144 ( .A(n4328), .B(n4492), .Z(n4494) );
  XOR U4145 ( .A(n4498), .B(n4499), .Z(n4328) );
  AND U4146 ( .A(n145), .B(n4500), .Z(n4499) );
  XOR U4147 ( .A(p_input[3675]), .B(p_input[3659]), .Z(n4500) );
  XOR U4148 ( .A(n4501), .B(n4502), .Z(n4492) );
  AND U4149 ( .A(n4503), .B(n4504), .Z(n4502) );
  XOR U4150 ( .A(n4501), .B(n4343), .Z(n4504) );
  XNOR U4151 ( .A(p_input[3690]), .B(n4505), .Z(n4343) );
  AND U4152 ( .A(n147), .B(n4506), .Z(n4505) );
  XOR U4153 ( .A(p_input[3706]), .B(p_input[3690]), .Z(n4506) );
  XNOR U4154 ( .A(n4340), .B(n4501), .Z(n4503) );
  XOR U4155 ( .A(n4507), .B(n4508), .Z(n4340) );
  AND U4156 ( .A(n145), .B(n4509), .Z(n4508) );
  XOR U4157 ( .A(p_input[3674]), .B(p_input[3658]), .Z(n4509) );
  XOR U4158 ( .A(n4510), .B(n4511), .Z(n4501) );
  AND U4159 ( .A(n4512), .B(n4513), .Z(n4511) );
  XOR U4160 ( .A(n4510), .B(n4355), .Z(n4513) );
  XNOR U4161 ( .A(p_input[3689]), .B(n4514), .Z(n4355) );
  AND U4162 ( .A(n147), .B(n4515), .Z(n4514) );
  XOR U4163 ( .A(p_input[3705]), .B(p_input[3689]), .Z(n4515) );
  XNOR U4164 ( .A(n4352), .B(n4510), .Z(n4512) );
  XOR U4165 ( .A(n4516), .B(n4517), .Z(n4352) );
  AND U4166 ( .A(n145), .B(n4518), .Z(n4517) );
  XOR U4167 ( .A(p_input[3673]), .B(p_input[3657]), .Z(n4518) );
  XOR U4168 ( .A(n4519), .B(n4520), .Z(n4510) );
  AND U4169 ( .A(n4521), .B(n4522), .Z(n4520) );
  XOR U4170 ( .A(n4519), .B(n4367), .Z(n4522) );
  XNOR U4171 ( .A(p_input[3688]), .B(n4523), .Z(n4367) );
  AND U4172 ( .A(n147), .B(n4524), .Z(n4523) );
  XOR U4173 ( .A(p_input[3704]), .B(p_input[3688]), .Z(n4524) );
  XNOR U4174 ( .A(n4364), .B(n4519), .Z(n4521) );
  XOR U4175 ( .A(n4525), .B(n4526), .Z(n4364) );
  AND U4176 ( .A(n145), .B(n4527), .Z(n4526) );
  XOR U4177 ( .A(p_input[3672]), .B(p_input[3656]), .Z(n4527) );
  XOR U4178 ( .A(n4528), .B(n4529), .Z(n4519) );
  AND U4179 ( .A(n4530), .B(n4531), .Z(n4529) );
  XOR U4180 ( .A(n4528), .B(n4379), .Z(n4531) );
  XNOR U4181 ( .A(p_input[3687]), .B(n4532), .Z(n4379) );
  AND U4182 ( .A(n147), .B(n4533), .Z(n4532) );
  XOR U4183 ( .A(p_input[3703]), .B(p_input[3687]), .Z(n4533) );
  XNOR U4184 ( .A(n4376), .B(n4528), .Z(n4530) );
  XOR U4185 ( .A(n4534), .B(n4535), .Z(n4376) );
  AND U4186 ( .A(n145), .B(n4536), .Z(n4535) );
  XOR U4187 ( .A(p_input[3671]), .B(p_input[3655]), .Z(n4536) );
  XOR U4188 ( .A(n4537), .B(n4538), .Z(n4528) );
  AND U4189 ( .A(n4539), .B(n4540), .Z(n4538) );
  XOR U4190 ( .A(n4537), .B(n4391), .Z(n4540) );
  XNOR U4191 ( .A(p_input[3686]), .B(n4541), .Z(n4391) );
  AND U4192 ( .A(n147), .B(n4542), .Z(n4541) );
  XOR U4193 ( .A(p_input[3702]), .B(p_input[3686]), .Z(n4542) );
  XNOR U4194 ( .A(n4388), .B(n4537), .Z(n4539) );
  XOR U4195 ( .A(n4543), .B(n4544), .Z(n4388) );
  AND U4196 ( .A(n145), .B(n4545), .Z(n4544) );
  XOR U4197 ( .A(p_input[3670]), .B(p_input[3654]), .Z(n4545) );
  XOR U4198 ( .A(n4546), .B(n4547), .Z(n4537) );
  AND U4199 ( .A(n4548), .B(n4549), .Z(n4547) );
  XOR U4200 ( .A(n4546), .B(n4403), .Z(n4549) );
  XNOR U4201 ( .A(p_input[3685]), .B(n4550), .Z(n4403) );
  AND U4202 ( .A(n147), .B(n4551), .Z(n4550) );
  XOR U4203 ( .A(p_input[3701]), .B(p_input[3685]), .Z(n4551) );
  XNOR U4204 ( .A(n4400), .B(n4546), .Z(n4548) );
  XOR U4205 ( .A(n4552), .B(n4553), .Z(n4400) );
  AND U4206 ( .A(n145), .B(n4554), .Z(n4553) );
  XOR U4207 ( .A(p_input[3669]), .B(p_input[3653]), .Z(n4554) );
  XOR U4208 ( .A(n4555), .B(n4556), .Z(n4546) );
  AND U4209 ( .A(n4557), .B(n4558), .Z(n4556) );
  XOR U4210 ( .A(n4555), .B(n4415), .Z(n4558) );
  XNOR U4211 ( .A(p_input[3684]), .B(n4559), .Z(n4415) );
  AND U4212 ( .A(n147), .B(n4560), .Z(n4559) );
  XOR U4213 ( .A(p_input[3700]), .B(p_input[3684]), .Z(n4560) );
  XNOR U4214 ( .A(n4412), .B(n4555), .Z(n4557) );
  XOR U4215 ( .A(n4561), .B(n4562), .Z(n4412) );
  AND U4216 ( .A(n145), .B(n4563), .Z(n4562) );
  XOR U4217 ( .A(p_input[3668]), .B(p_input[3652]), .Z(n4563) );
  XOR U4218 ( .A(n4564), .B(n4565), .Z(n4555) );
  AND U4219 ( .A(n4566), .B(n4567), .Z(n4565) );
  XOR U4220 ( .A(n4564), .B(n4427), .Z(n4567) );
  XNOR U4221 ( .A(p_input[3683]), .B(n4568), .Z(n4427) );
  AND U4222 ( .A(n147), .B(n4569), .Z(n4568) );
  XOR U4223 ( .A(p_input[3699]), .B(p_input[3683]), .Z(n4569) );
  XNOR U4224 ( .A(n4424), .B(n4564), .Z(n4566) );
  XOR U4225 ( .A(n4570), .B(n4571), .Z(n4424) );
  AND U4226 ( .A(n145), .B(n4572), .Z(n4571) );
  XOR U4227 ( .A(p_input[3667]), .B(p_input[3651]), .Z(n4572) );
  XOR U4228 ( .A(n4573), .B(n4574), .Z(n4564) );
  AND U4229 ( .A(n4575), .B(n4576), .Z(n4574) );
  XOR U4230 ( .A(n4573), .B(n4439), .Z(n4576) );
  XNOR U4231 ( .A(p_input[3682]), .B(n4577), .Z(n4439) );
  AND U4232 ( .A(n147), .B(n4578), .Z(n4577) );
  XOR U4233 ( .A(p_input[3698]), .B(p_input[3682]), .Z(n4578) );
  XNOR U4234 ( .A(n4436), .B(n4573), .Z(n4575) );
  XOR U4235 ( .A(n4579), .B(n4580), .Z(n4436) );
  AND U4236 ( .A(n145), .B(n4581), .Z(n4580) );
  XOR U4237 ( .A(p_input[3666]), .B(p_input[3650]), .Z(n4581) );
  XOR U4238 ( .A(n4582), .B(n4583), .Z(n4573) );
  AND U4239 ( .A(n4584), .B(n4585), .Z(n4583) );
  XNOR U4240 ( .A(n4586), .B(n4452), .Z(n4585) );
  XNOR U4241 ( .A(p_input[3681]), .B(n4587), .Z(n4452) );
  AND U4242 ( .A(n147), .B(n4588), .Z(n4587) );
  XNOR U4243 ( .A(p_input[3697]), .B(n4589), .Z(n4588) );
  IV U4244 ( .A(p_input[3681]), .Z(n4589) );
  XNOR U4245 ( .A(n4449), .B(n4582), .Z(n4584) );
  XNOR U4246 ( .A(p_input[3649]), .B(n4590), .Z(n4449) );
  AND U4247 ( .A(n145), .B(n4591), .Z(n4590) );
  XOR U4248 ( .A(p_input[3665]), .B(p_input[3649]), .Z(n4591) );
  IV U4249 ( .A(n4586), .Z(n4582) );
  AND U4250 ( .A(n4457), .B(n4460), .Z(n4586) );
  XOR U4251 ( .A(p_input[3680]), .B(n4592), .Z(n4460) );
  AND U4252 ( .A(n147), .B(n4593), .Z(n4592) );
  XOR U4253 ( .A(p_input[3696]), .B(p_input[3680]), .Z(n4593) );
  XOR U4254 ( .A(n4594), .B(n4595), .Z(n147) );
  AND U4255 ( .A(n4596), .B(n4597), .Z(n4595) );
  XNOR U4256 ( .A(p_input[3711]), .B(n4594), .Z(n4597) );
  XOR U4257 ( .A(n4594), .B(p_input[3695]), .Z(n4596) );
  XOR U4258 ( .A(n4598), .B(n4599), .Z(n4594) );
  AND U4259 ( .A(n4600), .B(n4601), .Z(n4599) );
  XNOR U4260 ( .A(p_input[3710]), .B(n4598), .Z(n4601) );
  XOR U4261 ( .A(n4598), .B(p_input[3694]), .Z(n4600) );
  XOR U4262 ( .A(n4602), .B(n4603), .Z(n4598) );
  AND U4263 ( .A(n4604), .B(n4605), .Z(n4603) );
  XNOR U4264 ( .A(p_input[3709]), .B(n4602), .Z(n4605) );
  XOR U4265 ( .A(n4602), .B(p_input[3693]), .Z(n4604) );
  XOR U4266 ( .A(n4606), .B(n4607), .Z(n4602) );
  AND U4267 ( .A(n4608), .B(n4609), .Z(n4607) );
  XNOR U4268 ( .A(p_input[3708]), .B(n4606), .Z(n4609) );
  XOR U4269 ( .A(n4606), .B(p_input[3692]), .Z(n4608) );
  XOR U4270 ( .A(n4610), .B(n4611), .Z(n4606) );
  AND U4271 ( .A(n4612), .B(n4613), .Z(n4611) );
  XNOR U4272 ( .A(p_input[3707]), .B(n4610), .Z(n4613) );
  XOR U4273 ( .A(n4610), .B(p_input[3691]), .Z(n4612) );
  XOR U4274 ( .A(n4614), .B(n4615), .Z(n4610) );
  AND U4275 ( .A(n4616), .B(n4617), .Z(n4615) );
  XNOR U4276 ( .A(p_input[3706]), .B(n4614), .Z(n4617) );
  XOR U4277 ( .A(n4614), .B(p_input[3690]), .Z(n4616) );
  XOR U4278 ( .A(n4618), .B(n4619), .Z(n4614) );
  AND U4279 ( .A(n4620), .B(n4621), .Z(n4619) );
  XNOR U4280 ( .A(p_input[3705]), .B(n4618), .Z(n4621) );
  XOR U4281 ( .A(n4618), .B(p_input[3689]), .Z(n4620) );
  XOR U4282 ( .A(n4622), .B(n4623), .Z(n4618) );
  AND U4283 ( .A(n4624), .B(n4625), .Z(n4623) );
  XNOR U4284 ( .A(p_input[3704]), .B(n4622), .Z(n4625) );
  XOR U4285 ( .A(n4622), .B(p_input[3688]), .Z(n4624) );
  XOR U4286 ( .A(n4626), .B(n4627), .Z(n4622) );
  AND U4287 ( .A(n4628), .B(n4629), .Z(n4627) );
  XNOR U4288 ( .A(p_input[3703]), .B(n4626), .Z(n4629) );
  XOR U4289 ( .A(n4626), .B(p_input[3687]), .Z(n4628) );
  XOR U4290 ( .A(n4630), .B(n4631), .Z(n4626) );
  AND U4291 ( .A(n4632), .B(n4633), .Z(n4631) );
  XNOR U4292 ( .A(p_input[3702]), .B(n4630), .Z(n4633) );
  XOR U4293 ( .A(n4630), .B(p_input[3686]), .Z(n4632) );
  XOR U4294 ( .A(n4634), .B(n4635), .Z(n4630) );
  AND U4295 ( .A(n4636), .B(n4637), .Z(n4635) );
  XNOR U4296 ( .A(p_input[3701]), .B(n4634), .Z(n4637) );
  XOR U4297 ( .A(n4634), .B(p_input[3685]), .Z(n4636) );
  XOR U4298 ( .A(n4638), .B(n4639), .Z(n4634) );
  AND U4299 ( .A(n4640), .B(n4641), .Z(n4639) );
  XNOR U4300 ( .A(p_input[3700]), .B(n4638), .Z(n4641) );
  XOR U4301 ( .A(n4638), .B(p_input[3684]), .Z(n4640) );
  XOR U4302 ( .A(n4642), .B(n4643), .Z(n4638) );
  AND U4303 ( .A(n4644), .B(n4645), .Z(n4643) );
  XNOR U4304 ( .A(p_input[3699]), .B(n4642), .Z(n4645) );
  XOR U4305 ( .A(n4642), .B(p_input[3683]), .Z(n4644) );
  XOR U4306 ( .A(n4646), .B(n4647), .Z(n4642) );
  AND U4307 ( .A(n4648), .B(n4649), .Z(n4647) );
  XNOR U4308 ( .A(p_input[3698]), .B(n4646), .Z(n4649) );
  XOR U4309 ( .A(n4646), .B(p_input[3682]), .Z(n4648) );
  XNOR U4310 ( .A(n4650), .B(n4651), .Z(n4646) );
  AND U4311 ( .A(n4652), .B(n4653), .Z(n4651) );
  XOR U4312 ( .A(p_input[3697]), .B(n4650), .Z(n4653) );
  XNOR U4313 ( .A(p_input[3681]), .B(n4650), .Z(n4652) );
  AND U4314 ( .A(p_input[3696]), .B(n4654), .Z(n4650) );
  IV U4315 ( .A(p_input[3680]), .Z(n4654) );
  XNOR U4316 ( .A(p_input[3648]), .B(n4655), .Z(n4457) );
  AND U4317 ( .A(n145), .B(n4656), .Z(n4655) );
  XOR U4318 ( .A(p_input[3664]), .B(p_input[3648]), .Z(n4656) );
  XOR U4319 ( .A(n4657), .B(n4658), .Z(n145) );
  AND U4320 ( .A(n4659), .B(n4660), .Z(n4658) );
  XNOR U4321 ( .A(p_input[3679]), .B(n4657), .Z(n4660) );
  XOR U4322 ( .A(n4657), .B(p_input[3663]), .Z(n4659) );
  XOR U4323 ( .A(n4661), .B(n4662), .Z(n4657) );
  AND U4324 ( .A(n4663), .B(n4664), .Z(n4662) );
  XNOR U4325 ( .A(p_input[3678]), .B(n4661), .Z(n4664) );
  XNOR U4326 ( .A(n4661), .B(n4471), .Z(n4663) );
  IV U4327 ( .A(p_input[3662]), .Z(n4471) );
  XOR U4328 ( .A(n4665), .B(n4666), .Z(n4661) );
  AND U4329 ( .A(n4667), .B(n4668), .Z(n4666) );
  XNOR U4330 ( .A(p_input[3677]), .B(n4665), .Z(n4668) );
  XNOR U4331 ( .A(n4665), .B(n4480), .Z(n4667) );
  IV U4332 ( .A(p_input[3661]), .Z(n4480) );
  XOR U4333 ( .A(n4669), .B(n4670), .Z(n4665) );
  AND U4334 ( .A(n4671), .B(n4672), .Z(n4670) );
  XNOR U4335 ( .A(p_input[3676]), .B(n4669), .Z(n4672) );
  XNOR U4336 ( .A(n4669), .B(n4489), .Z(n4671) );
  IV U4337 ( .A(p_input[3660]), .Z(n4489) );
  XOR U4338 ( .A(n4673), .B(n4674), .Z(n4669) );
  AND U4339 ( .A(n4675), .B(n4676), .Z(n4674) );
  XNOR U4340 ( .A(p_input[3675]), .B(n4673), .Z(n4676) );
  XNOR U4341 ( .A(n4673), .B(n4498), .Z(n4675) );
  IV U4342 ( .A(p_input[3659]), .Z(n4498) );
  XOR U4343 ( .A(n4677), .B(n4678), .Z(n4673) );
  AND U4344 ( .A(n4679), .B(n4680), .Z(n4678) );
  XNOR U4345 ( .A(p_input[3674]), .B(n4677), .Z(n4680) );
  XNOR U4346 ( .A(n4677), .B(n4507), .Z(n4679) );
  IV U4347 ( .A(p_input[3658]), .Z(n4507) );
  XOR U4348 ( .A(n4681), .B(n4682), .Z(n4677) );
  AND U4349 ( .A(n4683), .B(n4684), .Z(n4682) );
  XNOR U4350 ( .A(p_input[3673]), .B(n4681), .Z(n4684) );
  XNOR U4351 ( .A(n4681), .B(n4516), .Z(n4683) );
  IV U4352 ( .A(p_input[3657]), .Z(n4516) );
  XOR U4353 ( .A(n4685), .B(n4686), .Z(n4681) );
  AND U4354 ( .A(n4687), .B(n4688), .Z(n4686) );
  XNOR U4355 ( .A(p_input[3672]), .B(n4685), .Z(n4688) );
  XNOR U4356 ( .A(n4685), .B(n4525), .Z(n4687) );
  IV U4357 ( .A(p_input[3656]), .Z(n4525) );
  XOR U4358 ( .A(n4689), .B(n4690), .Z(n4685) );
  AND U4359 ( .A(n4691), .B(n4692), .Z(n4690) );
  XNOR U4360 ( .A(p_input[3671]), .B(n4689), .Z(n4692) );
  XNOR U4361 ( .A(n4689), .B(n4534), .Z(n4691) );
  IV U4362 ( .A(p_input[3655]), .Z(n4534) );
  XOR U4363 ( .A(n4693), .B(n4694), .Z(n4689) );
  AND U4364 ( .A(n4695), .B(n4696), .Z(n4694) );
  XNOR U4365 ( .A(p_input[3670]), .B(n4693), .Z(n4696) );
  XNOR U4366 ( .A(n4693), .B(n4543), .Z(n4695) );
  IV U4367 ( .A(p_input[3654]), .Z(n4543) );
  XOR U4368 ( .A(n4697), .B(n4698), .Z(n4693) );
  AND U4369 ( .A(n4699), .B(n4700), .Z(n4698) );
  XNOR U4370 ( .A(p_input[3669]), .B(n4697), .Z(n4700) );
  XNOR U4371 ( .A(n4697), .B(n4552), .Z(n4699) );
  IV U4372 ( .A(p_input[3653]), .Z(n4552) );
  XOR U4373 ( .A(n4701), .B(n4702), .Z(n4697) );
  AND U4374 ( .A(n4703), .B(n4704), .Z(n4702) );
  XNOR U4375 ( .A(p_input[3668]), .B(n4701), .Z(n4704) );
  XNOR U4376 ( .A(n4701), .B(n4561), .Z(n4703) );
  IV U4377 ( .A(p_input[3652]), .Z(n4561) );
  XOR U4378 ( .A(n4705), .B(n4706), .Z(n4701) );
  AND U4379 ( .A(n4707), .B(n4708), .Z(n4706) );
  XNOR U4380 ( .A(p_input[3667]), .B(n4705), .Z(n4708) );
  XNOR U4381 ( .A(n4705), .B(n4570), .Z(n4707) );
  IV U4382 ( .A(p_input[3651]), .Z(n4570) );
  XOR U4383 ( .A(n4709), .B(n4710), .Z(n4705) );
  AND U4384 ( .A(n4711), .B(n4712), .Z(n4710) );
  XNOR U4385 ( .A(p_input[3666]), .B(n4709), .Z(n4712) );
  XNOR U4386 ( .A(n4709), .B(n4579), .Z(n4711) );
  IV U4387 ( .A(p_input[3650]), .Z(n4579) );
  XNOR U4388 ( .A(n4713), .B(n4714), .Z(n4709) );
  AND U4389 ( .A(n4715), .B(n4716), .Z(n4714) );
  XOR U4390 ( .A(p_input[3665]), .B(n4713), .Z(n4716) );
  XNOR U4391 ( .A(p_input[3649]), .B(n4713), .Z(n4715) );
  AND U4392 ( .A(p_input[3664]), .B(n4717), .Z(n4713) );
  IV U4393 ( .A(p_input[3648]), .Z(n4717) );
  XOR U4394 ( .A(n4718), .B(n4719), .Z(n4276) );
  AND U4395 ( .A(n372), .B(n4720), .Z(n4719) );
  XNOR U4396 ( .A(n4721), .B(n4718), .Z(n4720) );
  XOR U4397 ( .A(n4722), .B(n4723), .Z(n372) );
  AND U4398 ( .A(n4724), .B(n4725), .Z(n4723) );
  XNOR U4399 ( .A(n4287), .B(n4722), .Z(n4725) );
  AND U4400 ( .A(p_input[3647]), .B(p_input[3631]), .Z(n4287) );
  XOR U4401 ( .A(n4722), .B(n4286), .Z(n4724) );
  AND U4402 ( .A(p_input[3599]), .B(p_input[3615]), .Z(n4286) );
  XOR U4403 ( .A(n4726), .B(n4727), .Z(n4722) );
  AND U4404 ( .A(n4728), .B(n4729), .Z(n4727) );
  XOR U4405 ( .A(n4726), .B(n4299), .Z(n4729) );
  XNOR U4406 ( .A(p_input[3630]), .B(n4730), .Z(n4299) );
  AND U4407 ( .A(n151), .B(n4731), .Z(n4730) );
  XOR U4408 ( .A(p_input[3646]), .B(p_input[3630]), .Z(n4731) );
  XNOR U4409 ( .A(n4296), .B(n4726), .Z(n4728) );
  XOR U4410 ( .A(n4732), .B(n4733), .Z(n4296) );
  AND U4411 ( .A(n148), .B(n4734), .Z(n4733) );
  XOR U4412 ( .A(p_input[3614]), .B(p_input[3598]), .Z(n4734) );
  XOR U4413 ( .A(n4735), .B(n4736), .Z(n4726) );
  AND U4414 ( .A(n4737), .B(n4738), .Z(n4736) );
  XOR U4415 ( .A(n4735), .B(n4311), .Z(n4738) );
  XNOR U4416 ( .A(p_input[3629]), .B(n4739), .Z(n4311) );
  AND U4417 ( .A(n151), .B(n4740), .Z(n4739) );
  XOR U4418 ( .A(p_input[3645]), .B(p_input[3629]), .Z(n4740) );
  XNOR U4419 ( .A(n4308), .B(n4735), .Z(n4737) );
  XOR U4420 ( .A(n4741), .B(n4742), .Z(n4308) );
  AND U4421 ( .A(n148), .B(n4743), .Z(n4742) );
  XOR U4422 ( .A(p_input[3613]), .B(p_input[3597]), .Z(n4743) );
  XOR U4423 ( .A(n4744), .B(n4745), .Z(n4735) );
  AND U4424 ( .A(n4746), .B(n4747), .Z(n4745) );
  XOR U4425 ( .A(n4744), .B(n4323), .Z(n4747) );
  XNOR U4426 ( .A(p_input[3628]), .B(n4748), .Z(n4323) );
  AND U4427 ( .A(n151), .B(n4749), .Z(n4748) );
  XOR U4428 ( .A(p_input[3644]), .B(p_input[3628]), .Z(n4749) );
  XNOR U4429 ( .A(n4320), .B(n4744), .Z(n4746) );
  XOR U4430 ( .A(n4750), .B(n4751), .Z(n4320) );
  AND U4431 ( .A(n148), .B(n4752), .Z(n4751) );
  XOR U4432 ( .A(p_input[3612]), .B(p_input[3596]), .Z(n4752) );
  XOR U4433 ( .A(n4753), .B(n4754), .Z(n4744) );
  AND U4434 ( .A(n4755), .B(n4756), .Z(n4754) );
  XOR U4435 ( .A(n4753), .B(n4335), .Z(n4756) );
  XNOR U4436 ( .A(p_input[3627]), .B(n4757), .Z(n4335) );
  AND U4437 ( .A(n151), .B(n4758), .Z(n4757) );
  XOR U4438 ( .A(p_input[3643]), .B(p_input[3627]), .Z(n4758) );
  XNOR U4439 ( .A(n4332), .B(n4753), .Z(n4755) );
  XOR U4440 ( .A(n4759), .B(n4760), .Z(n4332) );
  AND U4441 ( .A(n148), .B(n4761), .Z(n4760) );
  XOR U4442 ( .A(p_input[3611]), .B(p_input[3595]), .Z(n4761) );
  XOR U4443 ( .A(n4762), .B(n4763), .Z(n4753) );
  AND U4444 ( .A(n4764), .B(n4765), .Z(n4763) );
  XOR U4445 ( .A(n4762), .B(n4347), .Z(n4765) );
  XNOR U4446 ( .A(p_input[3626]), .B(n4766), .Z(n4347) );
  AND U4447 ( .A(n151), .B(n4767), .Z(n4766) );
  XOR U4448 ( .A(p_input[3642]), .B(p_input[3626]), .Z(n4767) );
  XNOR U4449 ( .A(n4344), .B(n4762), .Z(n4764) );
  XOR U4450 ( .A(n4768), .B(n4769), .Z(n4344) );
  AND U4451 ( .A(n148), .B(n4770), .Z(n4769) );
  XOR U4452 ( .A(p_input[3610]), .B(p_input[3594]), .Z(n4770) );
  XOR U4453 ( .A(n4771), .B(n4772), .Z(n4762) );
  AND U4454 ( .A(n4773), .B(n4774), .Z(n4772) );
  XOR U4455 ( .A(n4771), .B(n4359), .Z(n4774) );
  XNOR U4456 ( .A(p_input[3625]), .B(n4775), .Z(n4359) );
  AND U4457 ( .A(n151), .B(n4776), .Z(n4775) );
  XOR U4458 ( .A(p_input[3641]), .B(p_input[3625]), .Z(n4776) );
  XNOR U4459 ( .A(n4356), .B(n4771), .Z(n4773) );
  XOR U4460 ( .A(n4777), .B(n4778), .Z(n4356) );
  AND U4461 ( .A(n148), .B(n4779), .Z(n4778) );
  XOR U4462 ( .A(p_input[3609]), .B(p_input[3593]), .Z(n4779) );
  XOR U4463 ( .A(n4780), .B(n4781), .Z(n4771) );
  AND U4464 ( .A(n4782), .B(n4783), .Z(n4781) );
  XOR U4465 ( .A(n4780), .B(n4371), .Z(n4783) );
  XNOR U4466 ( .A(p_input[3624]), .B(n4784), .Z(n4371) );
  AND U4467 ( .A(n151), .B(n4785), .Z(n4784) );
  XOR U4468 ( .A(p_input[3640]), .B(p_input[3624]), .Z(n4785) );
  XNOR U4469 ( .A(n4368), .B(n4780), .Z(n4782) );
  XOR U4470 ( .A(n4786), .B(n4787), .Z(n4368) );
  AND U4471 ( .A(n148), .B(n4788), .Z(n4787) );
  XOR U4472 ( .A(p_input[3608]), .B(p_input[3592]), .Z(n4788) );
  XOR U4473 ( .A(n4789), .B(n4790), .Z(n4780) );
  AND U4474 ( .A(n4791), .B(n4792), .Z(n4790) );
  XOR U4475 ( .A(n4789), .B(n4383), .Z(n4792) );
  XNOR U4476 ( .A(p_input[3623]), .B(n4793), .Z(n4383) );
  AND U4477 ( .A(n151), .B(n4794), .Z(n4793) );
  XOR U4478 ( .A(p_input[3639]), .B(p_input[3623]), .Z(n4794) );
  XNOR U4479 ( .A(n4380), .B(n4789), .Z(n4791) );
  XOR U4480 ( .A(n4795), .B(n4796), .Z(n4380) );
  AND U4481 ( .A(n148), .B(n4797), .Z(n4796) );
  XOR U4482 ( .A(p_input[3607]), .B(p_input[3591]), .Z(n4797) );
  XOR U4483 ( .A(n4798), .B(n4799), .Z(n4789) );
  AND U4484 ( .A(n4800), .B(n4801), .Z(n4799) );
  XOR U4485 ( .A(n4798), .B(n4395), .Z(n4801) );
  XNOR U4486 ( .A(p_input[3622]), .B(n4802), .Z(n4395) );
  AND U4487 ( .A(n151), .B(n4803), .Z(n4802) );
  XOR U4488 ( .A(p_input[3638]), .B(p_input[3622]), .Z(n4803) );
  XNOR U4489 ( .A(n4392), .B(n4798), .Z(n4800) );
  XOR U4490 ( .A(n4804), .B(n4805), .Z(n4392) );
  AND U4491 ( .A(n148), .B(n4806), .Z(n4805) );
  XOR U4492 ( .A(p_input[3606]), .B(p_input[3590]), .Z(n4806) );
  XOR U4493 ( .A(n4807), .B(n4808), .Z(n4798) );
  AND U4494 ( .A(n4809), .B(n4810), .Z(n4808) );
  XOR U4495 ( .A(n4807), .B(n4407), .Z(n4810) );
  XNOR U4496 ( .A(p_input[3621]), .B(n4811), .Z(n4407) );
  AND U4497 ( .A(n151), .B(n4812), .Z(n4811) );
  XOR U4498 ( .A(p_input[3637]), .B(p_input[3621]), .Z(n4812) );
  XNOR U4499 ( .A(n4404), .B(n4807), .Z(n4809) );
  XOR U4500 ( .A(n4813), .B(n4814), .Z(n4404) );
  AND U4501 ( .A(n148), .B(n4815), .Z(n4814) );
  XOR U4502 ( .A(p_input[3605]), .B(p_input[3589]), .Z(n4815) );
  XOR U4503 ( .A(n4816), .B(n4817), .Z(n4807) );
  AND U4504 ( .A(n4818), .B(n4819), .Z(n4817) );
  XOR U4505 ( .A(n4816), .B(n4419), .Z(n4819) );
  XNOR U4506 ( .A(p_input[3620]), .B(n4820), .Z(n4419) );
  AND U4507 ( .A(n151), .B(n4821), .Z(n4820) );
  XOR U4508 ( .A(p_input[3636]), .B(p_input[3620]), .Z(n4821) );
  XNOR U4509 ( .A(n4416), .B(n4816), .Z(n4818) );
  XOR U4510 ( .A(n4822), .B(n4823), .Z(n4416) );
  AND U4511 ( .A(n148), .B(n4824), .Z(n4823) );
  XOR U4512 ( .A(p_input[3604]), .B(p_input[3588]), .Z(n4824) );
  XOR U4513 ( .A(n4825), .B(n4826), .Z(n4816) );
  AND U4514 ( .A(n4827), .B(n4828), .Z(n4826) );
  XOR U4515 ( .A(n4825), .B(n4431), .Z(n4828) );
  XNOR U4516 ( .A(p_input[3619]), .B(n4829), .Z(n4431) );
  AND U4517 ( .A(n151), .B(n4830), .Z(n4829) );
  XOR U4518 ( .A(p_input[3635]), .B(p_input[3619]), .Z(n4830) );
  XNOR U4519 ( .A(n4428), .B(n4825), .Z(n4827) );
  XOR U4520 ( .A(n4831), .B(n4832), .Z(n4428) );
  AND U4521 ( .A(n148), .B(n4833), .Z(n4832) );
  XOR U4522 ( .A(p_input[3603]), .B(p_input[3587]), .Z(n4833) );
  XOR U4523 ( .A(n4834), .B(n4835), .Z(n4825) );
  AND U4524 ( .A(n4836), .B(n4837), .Z(n4835) );
  XOR U4525 ( .A(n4834), .B(n4443), .Z(n4837) );
  XNOR U4526 ( .A(p_input[3618]), .B(n4838), .Z(n4443) );
  AND U4527 ( .A(n151), .B(n4839), .Z(n4838) );
  XOR U4528 ( .A(p_input[3634]), .B(p_input[3618]), .Z(n4839) );
  XNOR U4529 ( .A(n4440), .B(n4834), .Z(n4836) );
  XOR U4530 ( .A(n4840), .B(n4841), .Z(n4440) );
  AND U4531 ( .A(n148), .B(n4842), .Z(n4841) );
  XOR U4532 ( .A(p_input[3602]), .B(p_input[3586]), .Z(n4842) );
  XOR U4533 ( .A(n4843), .B(n4844), .Z(n4834) );
  AND U4534 ( .A(n4845), .B(n4846), .Z(n4844) );
  XNOR U4535 ( .A(n4847), .B(n4456), .Z(n4846) );
  XNOR U4536 ( .A(p_input[3617]), .B(n4848), .Z(n4456) );
  AND U4537 ( .A(n151), .B(n4849), .Z(n4848) );
  XNOR U4538 ( .A(p_input[3633]), .B(n4850), .Z(n4849) );
  IV U4539 ( .A(p_input[3617]), .Z(n4850) );
  XNOR U4540 ( .A(n4453), .B(n4843), .Z(n4845) );
  XNOR U4541 ( .A(p_input[3585]), .B(n4851), .Z(n4453) );
  AND U4542 ( .A(n148), .B(n4852), .Z(n4851) );
  XOR U4543 ( .A(p_input[3601]), .B(p_input[3585]), .Z(n4852) );
  IV U4544 ( .A(n4847), .Z(n4843) );
  AND U4545 ( .A(n4718), .B(n4721), .Z(n4847) );
  XOR U4546 ( .A(p_input[3616]), .B(n4853), .Z(n4721) );
  AND U4547 ( .A(n151), .B(n4854), .Z(n4853) );
  XOR U4548 ( .A(p_input[3632]), .B(p_input[3616]), .Z(n4854) );
  XOR U4549 ( .A(n4855), .B(n4856), .Z(n151) );
  AND U4550 ( .A(n4857), .B(n4858), .Z(n4856) );
  XNOR U4551 ( .A(p_input[3647]), .B(n4855), .Z(n4858) );
  XOR U4552 ( .A(n4855), .B(p_input[3631]), .Z(n4857) );
  XOR U4553 ( .A(n4859), .B(n4860), .Z(n4855) );
  AND U4554 ( .A(n4861), .B(n4862), .Z(n4860) );
  XNOR U4555 ( .A(p_input[3646]), .B(n4859), .Z(n4862) );
  XOR U4556 ( .A(n4859), .B(p_input[3630]), .Z(n4861) );
  XOR U4557 ( .A(n4863), .B(n4864), .Z(n4859) );
  AND U4558 ( .A(n4865), .B(n4866), .Z(n4864) );
  XNOR U4559 ( .A(p_input[3645]), .B(n4863), .Z(n4866) );
  XOR U4560 ( .A(n4863), .B(p_input[3629]), .Z(n4865) );
  XOR U4561 ( .A(n4867), .B(n4868), .Z(n4863) );
  AND U4562 ( .A(n4869), .B(n4870), .Z(n4868) );
  XNOR U4563 ( .A(p_input[3644]), .B(n4867), .Z(n4870) );
  XOR U4564 ( .A(n4867), .B(p_input[3628]), .Z(n4869) );
  XOR U4565 ( .A(n4871), .B(n4872), .Z(n4867) );
  AND U4566 ( .A(n4873), .B(n4874), .Z(n4872) );
  XNOR U4567 ( .A(p_input[3643]), .B(n4871), .Z(n4874) );
  XOR U4568 ( .A(n4871), .B(p_input[3627]), .Z(n4873) );
  XOR U4569 ( .A(n4875), .B(n4876), .Z(n4871) );
  AND U4570 ( .A(n4877), .B(n4878), .Z(n4876) );
  XNOR U4571 ( .A(p_input[3642]), .B(n4875), .Z(n4878) );
  XOR U4572 ( .A(n4875), .B(p_input[3626]), .Z(n4877) );
  XOR U4573 ( .A(n4879), .B(n4880), .Z(n4875) );
  AND U4574 ( .A(n4881), .B(n4882), .Z(n4880) );
  XNOR U4575 ( .A(p_input[3641]), .B(n4879), .Z(n4882) );
  XOR U4576 ( .A(n4879), .B(p_input[3625]), .Z(n4881) );
  XOR U4577 ( .A(n4883), .B(n4884), .Z(n4879) );
  AND U4578 ( .A(n4885), .B(n4886), .Z(n4884) );
  XNOR U4579 ( .A(p_input[3640]), .B(n4883), .Z(n4886) );
  XOR U4580 ( .A(n4883), .B(p_input[3624]), .Z(n4885) );
  XOR U4581 ( .A(n4887), .B(n4888), .Z(n4883) );
  AND U4582 ( .A(n4889), .B(n4890), .Z(n4888) );
  XNOR U4583 ( .A(p_input[3639]), .B(n4887), .Z(n4890) );
  XOR U4584 ( .A(n4887), .B(p_input[3623]), .Z(n4889) );
  XOR U4585 ( .A(n4891), .B(n4892), .Z(n4887) );
  AND U4586 ( .A(n4893), .B(n4894), .Z(n4892) );
  XNOR U4587 ( .A(p_input[3638]), .B(n4891), .Z(n4894) );
  XOR U4588 ( .A(n4891), .B(p_input[3622]), .Z(n4893) );
  XOR U4589 ( .A(n4895), .B(n4896), .Z(n4891) );
  AND U4590 ( .A(n4897), .B(n4898), .Z(n4896) );
  XNOR U4591 ( .A(p_input[3637]), .B(n4895), .Z(n4898) );
  XOR U4592 ( .A(n4895), .B(p_input[3621]), .Z(n4897) );
  XOR U4593 ( .A(n4899), .B(n4900), .Z(n4895) );
  AND U4594 ( .A(n4901), .B(n4902), .Z(n4900) );
  XNOR U4595 ( .A(p_input[3636]), .B(n4899), .Z(n4902) );
  XOR U4596 ( .A(n4899), .B(p_input[3620]), .Z(n4901) );
  XOR U4597 ( .A(n4903), .B(n4904), .Z(n4899) );
  AND U4598 ( .A(n4905), .B(n4906), .Z(n4904) );
  XNOR U4599 ( .A(p_input[3635]), .B(n4903), .Z(n4906) );
  XOR U4600 ( .A(n4903), .B(p_input[3619]), .Z(n4905) );
  XOR U4601 ( .A(n4907), .B(n4908), .Z(n4903) );
  AND U4602 ( .A(n4909), .B(n4910), .Z(n4908) );
  XNOR U4603 ( .A(p_input[3634]), .B(n4907), .Z(n4910) );
  XOR U4604 ( .A(n4907), .B(p_input[3618]), .Z(n4909) );
  XNOR U4605 ( .A(n4911), .B(n4912), .Z(n4907) );
  AND U4606 ( .A(n4913), .B(n4914), .Z(n4912) );
  XOR U4607 ( .A(p_input[3633]), .B(n4911), .Z(n4914) );
  XNOR U4608 ( .A(p_input[3617]), .B(n4911), .Z(n4913) );
  AND U4609 ( .A(p_input[3632]), .B(n4915), .Z(n4911) );
  IV U4610 ( .A(p_input[3616]), .Z(n4915) );
  XNOR U4611 ( .A(p_input[3584]), .B(n4916), .Z(n4718) );
  AND U4612 ( .A(n148), .B(n4917), .Z(n4916) );
  XOR U4613 ( .A(p_input[3600]), .B(p_input[3584]), .Z(n4917) );
  XOR U4614 ( .A(n4918), .B(n4919), .Z(n148) );
  AND U4615 ( .A(n4920), .B(n4921), .Z(n4919) );
  XNOR U4616 ( .A(p_input[3615]), .B(n4918), .Z(n4921) );
  XOR U4617 ( .A(n4918), .B(p_input[3599]), .Z(n4920) );
  XOR U4618 ( .A(n4922), .B(n4923), .Z(n4918) );
  AND U4619 ( .A(n4924), .B(n4925), .Z(n4923) );
  XNOR U4620 ( .A(p_input[3614]), .B(n4922), .Z(n4925) );
  XNOR U4621 ( .A(n4922), .B(n4732), .Z(n4924) );
  IV U4622 ( .A(p_input[3598]), .Z(n4732) );
  XOR U4623 ( .A(n4926), .B(n4927), .Z(n4922) );
  AND U4624 ( .A(n4928), .B(n4929), .Z(n4927) );
  XNOR U4625 ( .A(p_input[3613]), .B(n4926), .Z(n4929) );
  XNOR U4626 ( .A(n4926), .B(n4741), .Z(n4928) );
  IV U4627 ( .A(p_input[3597]), .Z(n4741) );
  XOR U4628 ( .A(n4930), .B(n4931), .Z(n4926) );
  AND U4629 ( .A(n4932), .B(n4933), .Z(n4931) );
  XNOR U4630 ( .A(p_input[3612]), .B(n4930), .Z(n4933) );
  XNOR U4631 ( .A(n4930), .B(n4750), .Z(n4932) );
  IV U4632 ( .A(p_input[3596]), .Z(n4750) );
  XOR U4633 ( .A(n4934), .B(n4935), .Z(n4930) );
  AND U4634 ( .A(n4936), .B(n4937), .Z(n4935) );
  XNOR U4635 ( .A(p_input[3611]), .B(n4934), .Z(n4937) );
  XNOR U4636 ( .A(n4934), .B(n4759), .Z(n4936) );
  IV U4637 ( .A(p_input[3595]), .Z(n4759) );
  XOR U4638 ( .A(n4938), .B(n4939), .Z(n4934) );
  AND U4639 ( .A(n4940), .B(n4941), .Z(n4939) );
  XNOR U4640 ( .A(p_input[3610]), .B(n4938), .Z(n4941) );
  XNOR U4641 ( .A(n4938), .B(n4768), .Z(n4940) );
  IV U4642 ( .A(p_input[3594]), .Z(n4768) );
  XOR U4643 ( .A(n4942), .B(n4943), .Z(n4938) );
  AND U4644 ( .A(n4944), .B(n4945), .Z(n4943) );
  XNOR U4645 ( .A(p_input[3609]), .B(n4942), .Z(n4945) );
  XNOR U4646 ( .A(n4942), .B(n4777), .Z(n4944) );
  IV U4647 ( .A(p_input[3593]), .Z(n4777) );
  XOR U4648 ( .A(n4946), .B(n4947), .Z(n4942) );
  AND U4649 ( .A(n4948), .B(n4949), .Z(n4947) );
  XNOR U4650 ( .A(p_input[3608]), .B(n4946), .Z(n4949) );
  XNOR U4651 ( .A(n4946), .B(n4786), .Z(n4948) );
  IV U4652 ( .A(p_input[3592]), .Z(n4786) );
  XOR U4653 ( .A(n4950), .B(n4951), .Z(n4946) );
  AND U4654 ( .A(n4952), .B(n4953), .Z(n4951) );
  XNOR U4655 ( .A(p_input[3607]), .B(n4950), .Z(n4953) );
  XNOR U4656 ( .A(n4950), .B(n4795), .Z(n4952) );
  IV U4657 ( .A(p_input[3591]), .Z(n4795) );
  XOR U4658 ( .A(n4954), .B(n4955), .Z(n4950) );
  AND U4659 ( .A(n4956), .B(n4957), .Z(n4955) );
  XNOR U4660 ( .A(p_input[3606]), .B(n4954), .Z(n4957) );
  XNOR U4661 ( .A(n4954), .B(n4804), .Z(n4956) );
  IV U4662 ( .A(p_input[3590]), .Z(n4804) );
  XOR U4663 ( .A(n4958), .B(n4959), .Z(n4954) );
  AND U4664 ( .A(n4960), .B(n4961), .Z(n4959) );
  XNOR U4665 ( .A(p_input[3605]), .B(n4958), .Z(n4961) );
  XNOR U4666 ( .A(n4958), .B(n4813), .Z(n4960) );
  IV U4667 ( .A(p_input[3589]), .Z(n4813) );
  XOR U4668 ( .A(n4962), .B(n4963), .Z(n4958) );
  AND U4669 ( .A(n4964), .B(n4965), .Z(n4963) );
  XNOR U4670 ( .A(p_input[3604]), .B(n4962), .Z(n4965) );
  XNOR U4671 ( .A(n4962), .B(n4822), .Z(n4964) );
  IV U4672 ( .A(p_input[3588]), .Z(n4822) );
  XOR U4673 ( .A(n4966), .B(n4967), .Z(n4962) );
  AND U4674 ( .A(n4968), .B(n4969), .Z(n4967) );
  XNOR U4675 ( .A(p_input[3603]), .B(n4966), .Z(n4969) );
  XNOR U4676 ( .A(n4966), .B(n4831), .Z(n4968) );
  IV U4677 ( .A(p_input[3587]), .Z(n4831) );
  XOR U4678 ( .A(n4970), .B(n4971), .Z(n4966) );
  AND U4679 ( .A(n4972), .B(n4973), .Z(n4971) );
  XNOR U4680 ( .A(p_input[3602]), .B(n4970), .Z(n4973) );
  XNOR U4681 ( .A(n4970), .B(n4840), .Z(n4972) );
  IV U4682 ( .A(p_input[3586]), .Z(n4840) );
  XNOR U4683 ( .A(n4974), .B(n4975), .Z(n4970) );
  AND U4684 ( .A(n4976), .B(n4977), .Z(n4975) );
  XOR U4685 ( .A(p_input[3601]), .B(n4974), .Z(n4977) );
  XNOR U4686 ( .A(p_input[3585]), .B(n4974), .Z(n4976) );
  AND U4687 ( .A(p_input[3600]), .B(n4978), .Z(n4974) );
  IV U4688 ( .A(p_input[3584]), .Z(n4978) );
  XOR U4689 ( .A(n4979), .B(n4980), .Z(n1433) );
  AND U4690 ( .A(n1005), .B(n4981), .Z(n4980) );
  XNOR U4691 ( .A(n4982), .B(n4979), .Z(n4981) );
  XOR U4692 ( .A(n4983), .B(n4984), .Z(n1005) );
  AND U4693 ( .A(n4985), .B(n4986), .Z(n4984) );
  XOR U4694 ( .A(n4983), .B(n1448), .Z(n4986) );
  XNOR U4695 ( .A(n4987), .B(n4988), .Z(n1448) );
  AND U4696 ( .A(n4989), .B(n923), .Z(n4988) );
  AND U4697 ( .A(n4987), .B(n4990), .Z(n4989) );
  XNOR U4698 ( .A(n1445), .B(n4983), .Z(n4985) );
  XOR U4699 ( .A(n4991), .B(n4992), .Z(n1445) );
  AND U4700 ( .A(n4993), .B(n920), .Z(n4992) );
  NOR U4701 ( .A(n4991), .B(n4994), .Z(n4993) );
  XOR U4702 ( .A(n4995), .B(n4996), .Z(n4983) );
  AND U4703 ( .A(n4997), .B(n4998), .Z(n4996) );
  XOR U4704 ( .A(n4995), .B(n1460), .Z(n4998) );
  XOR U4705 ( .A(n4999), .B(n5000), .Z(n1460) );
  AND U4706 ( .A(n923), .B(n5001), .Z(n5000) );
  XOR U4707 ( .A(n5002), .B(n4999), .Z(n5001) );
  XNOR U4708 ( .A(n1457), .B(n4995), .Z(n4997) );
  XOR U4709 ( .A(n5003), .B(n5004), .Z(n1457) );
  AND U4710 ( .A(n920), .B(n5005), .Z(n5004) );
  XOR U4711 ( .A(n5006), .B(n5003), .Z(n5005) );
  XOR U4712 ( .A(n5007), .B(n5008), .Z(n4995) );
  AND U4713 ( .A(n5009), .B(n5010), .Z(n5008) );
  XOR U4714 ( .A(n5007), .B(n1472), .Z(n5010) );
  XOR U4715 ( .A(n5011), .B(n5012), .Z(n1472) );
  AND U4716 ( .A(n923), .B(n5013), .Z(n5012) );
  XOR U4717 ( .A(n5014), .B(n5011), .Z(n5013) );
  XNOR U4718 ( .A(n1469), .B(n5007), .Z(n5009) );
  XOR U4719 ( .A(n5015), .B(n5016), .Z(n1469) );
  AND U4720 ( .A(n920), .B(n5017), .Z(n5016) );
  XOR U4721 ( .A(n5018), .B(n5015), .Z(n5017) );
  XOR U4722 ( .A(n5019), .B(n5020), .Z(n5007) );
  AND U4723 ( .A(n5021), .B(n5022), .Z(n5020) );
  XOR U4724 ( .A(n5019), .B(n1484), .Z(n5022) );
  XOR U4725 ( .A(n5023), .B(n5024), .Z(n1484) );
  AND U4726 ( .A(n923), .B(n5025), .Z(n5024) );
  XOR U4727 ( .A(n5026), .B(n5023), .Z(n5025) );
  XNOR U4728 ( .A(n1481), .B(n5019), .Z(n5021) );
  XOR U4729 ( .A(n5027), .B(n5028), .Z(n1481) );
  AND U4730 ( .A(n920), .B(n5029), .Z(n5028) );
  XOR U4731 ( .A(n5030), .B(n5027), .Z(n5029) );
  XOR U4732 ( .A(n5031), .B(n5032), .Z(n5019) );
  AND U4733 ( .A(n5033), .B(n5034), .Z(n5032) );
  XOR U4734 ( .A(n5031), .B(n1496), .Z(n5034) );
  XOR U4735 ( .A(n5035), .B(n5036), .Z(n1496) );
  AND U4736 ( .A(n923), .B(n5037), .Z(n5036) );
  XOR U4737 ( .A(n5038), .B(n5035), .Z(n5037) );
  XNOR U4738 ( .A(n1493), .B(n5031), .Z(n5033) );
  XOR U4739 ( .A(n5039), .B(n5040), .Z(n1493) );
  AND U4740 ( .A(n920), .B(n5041), .Z(n5040) );
  XOR U4741 ( .A(n5042), .B(n5039), .Z(n5041) );
  XOR U4742 ( .A(n5043), .B(n5044), .Z(n5031) );
  AND U4743 ( .A(n5045), .B(n5046), .Z(n5044) );
  XOR U4744 ( .A(n5043), .B(n1508), .Z(n5046) );
  XOR U4745 ( .A(n5047), .B(n5048), .Z(n1508) );
  AND U4746 ( .A(n923), .B(n5049), .Z(n5048) );
  XOR U4747 ( .A(n5050), .B(n5047), .Z(n5049) );
  XNOR U4748 ( .A(n1505), .B(n5043), .Z(n5045) );
  XOR U4749 ( .A(n5051), .B(n5052), .Z(n1505) );
  AND U4750 ( .A(n920), .B(n5053), .Z(n5052) );
  XOR U4751 ( .A(n5054), .B(n5051), .Z(n5053) );
  XOR U4752 ( .A(n5055), .B(n5056), .Z(n5043) );
  AND U4753 ( .A(n5057), .B(n5058), .Z(n5056) );
  XOR U4754 ( .A(n5055), .B(n1520), .Z(n5058) );
  XOR U4755 ( .A(n5059), .B(n5060), .Z(n1520) );
  AND U4756 ( .A(n923), .B(n5061), .Z(n5060) );
  XOR U4757 ( .A(n5062), .B(n5059), .Z(n5061) );
  XNOR U4758 ( .A(n1517), .B(n5055), .Z(n5057) );
  XOR U4759 ( .A(n5063), .B(n5064), .Z(n1517) );
  AND U4760 ( .A(n920), .B(n5065), .Z(n5064) );
  XOR U4761 ( .A(n5066), .B(n5063), .Z(n5065) );
  XOR U4762 ( .A(n5067), .B(n5068), .Z(n5055) );
  AND U4763 ( .A(n5069), .B(n5070), .Z(n5068) );
  XOR U4764 ( .A(n5067), .B(n1532), .Z(n5070) );
  XOR U4765 ( .A(n5071), .B(n5072), .Z(n1532) );
  AND U4766 ( .A(n923), .B(n5073), .Z(n5072) );
  XOR U4767 ( .A(n5074), .B(n5071), .Z(n5073) );
  XNOR U4768 ( .A(n1529), .B(n5067), .Z(n5069) );
  XOR U4769 ( .A(n5075), .B(n5076), .Z(n1529) );
  AND U4770 ( .A(n920), .B(n5077), .Z(n5076) );
  XOR U4771 ( .A(n5078), .B(n5075), .Z(n5077) );
  XOR U4772 ( .A(n5079), .B(n5080), .Z(n5067) );
  AND U4773 ( .A(n5081), .B(n5082), .Z(n5080) );
  XOR U4774 ( .A(n5079), .B(n1544), .Z(n5082) );
  XOR U4775 ( .A(n5083), .B(n5084), .Z(n1544) );
  AND U4776 ( .A(n923), .B(n5085), .Z(n5084) );
  XOR U4777 ( .A(n5086), .B(n5083), .Z(n5085) );
  XNOR U4778 ( .A(n1541), .B(n5079), .Z(n5081) );
  XOR U4779 ( .A(n5087), .B(n5088), .Z(n1541) );
  AND U4780 ( .A(n920), .B(n5089), .Z(n5088) );
  XOR U4781 ( .A(n5090), .B(n5087), .Z(n5089) );
  XOR U4782 ( .A(n5091), .B(n5092), .Z(n5079) );
  AND U4783 ( .A(n5093), .B(n5094), .Z(n5092) );
  XOR U4784 ( .A(n5091), .B(n1556), .Z(n5094) );
  XOR U4785 ( .A(n5095), .B(n5096), .Z(n1556) );
  AND U4786 ( .A(n923), .B(n5097), .Z(n5096) );
  XOR U4787 ( .A(n5098), .B(n5095), .Z(n5097) );
  XNOR U4788 ( .A(n1553), .B(n5091), .Z(n5093) );
  XOR U4789 ( .A(n5099), .B(n5100), .Z(n1553) );
  AND U4790 ( .A(n920), .B(n5101), .Z(n5100) );
  XOR U4791 ( .A(n5102), .B(n5099), .Z(n5101) );
  XOR U4792 ( .A(n5103), .B(n5104), .Z(n5091) );
  AND U4793 ( .A(n5105), .B(n5106), .Z(n5104) );
  XOR U4794 ( .A(n5103), .B(n1568), .Z(n5106) );
  XOR U4795 ( .A(n5107), .B(n5108), .Z(n1568) );
  AND U4796 ( .A(n923), .B(n5109), .Z(n5108) );
  XOR U4797 ( .A(n5110), .B(n5107), .Z(n5109) );
  XNOR U4798 ( .A(n1565), .B(n5103), .Z(n5105) );
  XOR U4799 ( .A(n5111), .B(n5112), .Z(n1565) );
  AND U4800 ( .A(n920), .B(n5113), .Z(n5112) );
  XOR U4801 ( .A(n5114), .B(n5111), .Z(n5113) );
  XOR U4802 ( .A(n5115), .B(n5116), .Z(n5103) );
  AND U4803 ( .A(n5117), .B(n5118), .Z(n5116) );
  XOR U4804 ( .A(n5115), .B(n1580), .Z(n5118) );
  XOR U4805 ( .A(n5119), .B(n5120), .Z(n1580) );
  AND U4806 ( .A(n923), .B(n5121), .Z(n5120) );
  XOR U4807 ( .A(n5122), .B(n5119), .Z(n5121) );
  XNOR U4808 ( .A(n1577), .B(n5115), .Z(n5117) );
  XOR U4809 ( .A(n5123), .B(n5124), .Z(n1577) );
  AND U4810 ( .A(n920), .B(n5125), .Z(n5124) );
  XOR U4811 ( .A(n5126), .B(n5123), .Z(n5125) );
  XOR U4812 ( .A(n5127), .B(n5128), .Z(n5115) );
  AND U4813 ( .A(n5129), .B(n5130), .Z(n5128) );
  XOR U4814 ( .A(n5127), .B(n1592), .Z(n5130) );
  XOR U4815 ( .A(n5131), .B(n5132), .Z(n1592) );
  AND U4816 ( .A(n923), .B(n5133), .Z(n5132) );
  XOR U4817 ( .A(n5134), .B(n5131), .Z(n5133) );
  XNOR U4818 ( .A(n1589), .B(n5127), .Z(n5129) );
  XOR U4819 ( .A(n5135), .B(n5136), .Z(n1589) );
  AND U4820 ( .A(n920), .B(n5137), .Z(n5136) );
  XOR U4821 ( .A(n5138), .B(n5135), .Z(n5137) );
  XOR U4822 ( .A(n5139), .B(n5140), .Z(n5127) );
  AND U4823 ( .A(n5141), .B(n5142), .Z(n5140) );
  XOR U4824 ( .A(n5139), .B(n1604), .Z(n5142) );
  XOR U4825 ( .A(n5143), .B(n5144), .Z(n1604) );
  AND U4826 ( .A(n923), .B(n5145), .Z(n5144) );
  XOR U4827 ( .A(n5146), .B(n5143), .Z(n5145) );
  XNOR U4828 ( .A(n1601), .B(n5139), .Z(n5141) );
  XOR U4829 ( .A(n5147), .B(n5148), .Z(n1601) );
  AND U4830 ( .A(n920), .B(n5149), .Z(n5148) );
  XOR U4831 ( .A(n5150), .B(n5147), .Z(n5149) );
  XOR U4832 ( .A(n5151), .B(n5152), .Z(n5139) );
  AND U4833 ( .A(n5153), .B(n5154), .Z(n5152) );
  XNOR U4834 ( .A(n5155), .B(n1617), .Z(n5154) );
  XOR U4835 ( .A(n5156), .B(n5157), .Z(n1617) );
  AND U4836 ( .A(n923), .B(n5158), .Z(n5157) );
  XOR U4837 ( .A(n5156), .B(n5159), .Z(n5158) );
  XNOR U4838 ( .A(n1614), .B(n5151), .Z(n5153) );
  XOR U4839 ( .A(n5160), .B(n5161), .Z(n1614) );
  AND U4840 ( .A(n920), .B(n5162), .Z(n5161) );
  XOR U4841 ( .A(n5160), .B(n5163), .Z(n5162) );
  IV U4842 ( .A(n5155), .Z(n5151) );
  AND U4843 ( .A(n4979), .B(n4982), .Z(n5155) );
  XNOR U4844 ( .A(n5164), .B(n5165), .Z(n4982) );
  AND U4845 ( .A(n923), .B(n5166), .Z(n5165) );
  XNOR U4846 ( .A(n5167), .B(n5164), .Z(n5166) );
  XOR U4847 ( .A(n5168), .B(n5169), .Z(n923) );
  AND U4848 ( .A(n5170), .B(n5171), .Z(n5169) );
  XOR U4849 ( .A(n4990), .B(n5168), .Z(n5171) );
  IV U4850 ( .A(n5172), .Z(n4990) );
  AND U4851 ( .A(n5173), .B(n5174), .Z(n5172) );
  XOR U4852 ( .A(n5168), .B(n4987), .Z(n5170) );
  AND U4853 ( .A(n5175), .B(n5176), .Z(n4987) );
  XOR U4854 ( .A(n5177), .B(n5178), .Z(n5168) );
  AND U4855 ( .A(n5179), .B(n5180), .Z(n5178) );
  XOR U4856 ( .A(n5177), .B(n5002), .Z(n5180) );
  XOR U4857 ( .A(n5181), .B(n5182), .Z(n5002) );
  AND U4858 ( .A(n747), .B(n5183), .Z(n5182) );
  XOR U4859 ( .A(n5184), .B(n5181), .Z(n5183) );
  XNOR U4860 ( .A(n4999), .B(n5177), .Z(n5179) );
  XOR U4861 ( .A(n5185), .B(n5186), .Z(n4999) );
  AND U4862 ( .A(n745), .B(n5187), .Z(n5186) );
  XOR U4863 ( .A(n5188), .B(n5185), .Z(n5187) );
  XOR U4864 ( .A(n5189), .B(n5190), .Z(n5177) );
  AND U4865 ( .A(n5191), .B(n5192), .Z(n5190) );
  XOR U4866 ( .A(n5189), .B(n5014), .Z(n5192) );
  XOR U4867 ( .A(n5193), .B(n5194), .Z(n5014) );
  AND U4868 ( .A(n747), .B(n5195), .Z(n5194) );
  XOR U4869 ( .A(n5196), .B(n5193), .Z(n5195) );
  XNOR U4870 ( .A(n5011), .B(n5189), .Z(n5191) );
  XOR U4871 ( .A(n5197), .B(n5198), .Z(n5011) );
  AND U4872 ( .A(n745), .B(n5199), .Z(n5198) );
  XOR U4873 ( .A(n5200), .B(n5197), .Z(n5199) );
  XOR U4874 ( .A(n5201), .B(n5202), .Z(n5189) );
  AND U4875 ( .A(n5203), .B(n5204), .Z(n5202) );
  XOR U4876 ( .A(n5201), .B(n5026), .Z(n5204) );
  XOR U4877 ( .A(n5205), .B(n5206), .Z(n5026) );
  AND U4878 ( .A(n747), .B(n5207), .Z(n5206) );
  XOR U4879 ( .A(n5208), .B(n5205), .Z(n5207) );
  XNOR U4880 ( .A(n5023), .B(n5201), .Z(n5203) );
  XOR U4881 ( .A(n5209), .B(n5210), .Z(n5023) );
  AND U4882 ( .A(n745), .B(n5211), .Z(n5210) );
  XOR U4883 ( .A(n5212), .B(n5209), .Z(n5211) );
  XOR U4884 ( .A(n5213), .B(n5214), .Z(n5201) );
  AND U4885 ( .A(n5215), .B(n5216), .Z(n5214) );
  XOR U4886 ( .A(n5213), .B(n5038), .Z(n5216) );
  XOR U4887 ( .A(n5217), .B(n5218), .Z(n5038) );
  AND U4888 ( .A(n747), .B(n5219), .Z(n5218) );
  XOR U4889 ( .A(n5220), .B(n5217), .Z(n5219) );
  XNOR U4890 ( .A(n5035), .B(n5213), .Z(n5215) );
  XOR U4891 ( .A(n5221), .B(n5222), .Z(n5035) );
  AND U4892 ( .A(n745), .B(n5223), .Z(n5222) );
  XOR U4893 ( .A(n5224), .B(n5221), .Z(n5223) );
  XOR U4894 ( .A(n5225), .B(n5226), .Z(n5213) );
  AND U4895 ( .A(n5227), .B(n5228), .Z(n5226) );
  XOR U4896 ( .A(n5225), .B(n5050), .Z(n5228) );
  XOR U4897 ( .A(n5229), .B(n5230), .Z(n5050) );
  AND U4898 ( .A(n747), .B(n5231), .Z(n5230) );
  XOR U4899 ( .A(n5232), .B(n5229), .Z(n5231) );
  XNOR U4900 ( .A(n5047), .B(n5225), .Z(n5227) );
  XOR U4901 ( .A(n5233), .B(n5234), .Z(n5047) );
  AND U4902 ( .A(n745), .B(n5235), .Z(n5234) );
  XOR U4903 ( .A(n5236), .B(n5233), .Z(n5235) );
  XOR U4904 ( .A(n5237), .B(n5238), .Z(n5225) );
  AND U4905 ( .A(n5239), .B(n5240), .Z(n5238) );
  XOR U4906 ( .A(n5237), .B(n5062), .Z(n5240) );
  XOR U4907 ( .A(n5241), .B(n5242), .Z(n5062) );
  AND U4908 ( .A(n747), .B(n5243), .Z(n5242) );
  XOR U4909 ( .A(n5244), .B(n5241), .Z(n5243) );
  XNOR U4910 ( .A(n5059), .B(n5237), .Z(n5239) );
  XOR U4911 ( .A(n5245), .B(n5246), .Z(n5059) );
  AND U4912 ( .A(n745), .B(n5247), .Z(n5246) );
  XOR U4913 ( .A(n5248), .B(n5245), .Z(n5247) );
  XOR U4914 ( .A(n5249), .B(n5250), .Z(n5237) );
  AND U4915 ( .A(n5251), .B(n5252), .Z(n5250) );
  XOR U4916 ( .A(n5249), .B(n5074), .Z(n5252) );
  XOR U4917 ( .A(n5253), .B(n5254), .Z(n5074) );
  AND U4918 ( .A(n747), .B(n5255), .Z(n5254) );
  XOR U4919 ( .A(n5256), .B(n5253), .Z(n5255) );
  XNOR U4920 ( .A(n5071), .B(n5249), .Z(n5251) );
  XOR U4921 ( .A(n5257), .B(n5258), .Z(n5071) );
  AND U4922 ( .A(n745), .B(n5259), .Z(n5258) );
  XOR U4923 ( .A(n5260), .B(n5257), .Z(n5259) );
  XOR U4924 ( .A(n5261), .B(n5262), .Z(n5249) );
  AND U4925 ( .A(n5263), .B(n5264), .Z(n5262) );
  XOR U4926 ( .A(n5261), .B(n5086), .Z(n5264) );
  XOR U4927 ( .A(n5265), .B(n5266), .Z(n5086) );
  AND U4928 ( .A(n747), .B(n5267), .Z(n5266) );
  XOR U4929 ( .A(n5268), .B(n5265), .Z(n5267) );
  XNOR U4930 ( .A(n5083), .B(n5261), .Z(n5263) );
  XOR U4931 ( .A(n5269), .B(n5270), .Z(n5083) );
  AND U4932 ( .A(n745), .B(n5271), .Z(n5270) );
  XOR U4933 ( .A(n5272), .B(n5269), .Z(n5271) );
  XOR U4934 ( .A(n5273), .B(n5274), .Z(n5261) );
  AND U4935 ( .A(n5275), .B(n5276), .Z(n5274) );
  XOR U4936 ( .A(n5273), .B(n5098), .Z(n5276) );
  XOR U4937 ( .A(n5277), .B(n5278), .Z(n5098) );
  AND U4938 ( .A(n747), .B(n5279), .Z(n5278) );
  XOR U4939 ( .A(n5280), .B(n5277), .Z(n5279) );
  XNOR U4940 ( .A(n5095), .B(n5273), .Z(n5275) );
  XOR U4941 ( .A(n5281), .B(n5282), .Z(n5095) );
  AND U4942 ( .A(n745), .B(n5283), .Z(n5282) );
  XOR U4943 ( .A(n5284), .B(n5281), .Z(n5283) );
  XOR U4944 ( .A(n5285), .B(n5286), .Z(n5273) );
  AND U4945 ( .A(n5287), .B(n5288), .Z(n5286) );
  XOR U4946 ( .A(n5285), .B(n5110), .Z(n5288) );
  XOR U4947 ( .A(n5289), .B(n5290), .Z(n5110) );
  AND U4948 ( .A(n747), .B(n5291), .Z(n5290) );
  XOR U4949 ( .A(n5292), .B(n5289), .Z(n5291) );
  XNOR U4950 ( .A(n5107), .B(n5285), .Z(n5287) );
  XOR U4951 ( .A(n5293), .B(n5294), .Z(n5107) );
  AND U4952 ( .A(n745), .B(n5295), .Z(n5294) );
  XOR U4953 ( .A(n5296), .B(n5293), .Z(n5295) );
  XOR U4954 ( .A(n5297), .B(n5298), .Z(n5285) );
  AND U4955 ( .A(n5299), .B(n5300), .Z(n5298) );
  XOR U4956 ( .A(n5297), .B(n5122), .Z(n5300) );
  XOR U4957 ( .A(n5301), .B(n5302), .Z(n5122) );
  AND U4958 ( .A(n747), .B(n5303), .Z(n5302) );
  XOR U4959 ( .A(n5304), .B(n5301), .Z(n5303) );
  XNOR U4960 ( .A(n5119), .B(n5297), .Z(n5299) );
  XOR U4961 ( .A(n5305), .B(n5306), .Z(n5119) );
  AND U4962 ( .A(n745), .B(n5307), .Z(n5306) );
  XOR U4963 ( .A(n5308), .B(n5305), .Z(n5307) );
  XOR U4964 ( .A(n5309), .B(n5310), .Z(n5297) );
  AND U4965 ( .A(n5311), .B(n5312), .Z(n5310) );
  XOR U4966 ( .A(n5309), .B(n5134), .Z(n5312) );
  XOR U4967 ( .A(n5313), .B(n5314), .Z(n5134) );
  AND U4968 ( .A(n747), .B(n5315), .Z(n5314) );
  XOR U4969 ( .A(n5316), .B(n5313), .Z(n5315) );
  XNOR U4970 ( .A(n5131), .B(n5309), .Z(n5311) );
  XOR U4971 ( .A(n5317), .B(n5318), .Z(n5131) );
  AND U4972 ( .A(n745), .B(n5319), .Z(n5318) );
  XOR U4973 ( .A(n5320), .B(n5317), .Z(n5319) );
  XOR U4974 ( .A(n5321), .B(n5322), .Z(n5309) );
  AND U4975 ( .A(n5323), .B(n5324), .Z(n5322) );
  XOR U4976 ( .A(n5321), .B(n5146), .Z(n5324) );
  XOR U4977 ( .A(n5325), .B(n5326), .Z(n5146) );
  AND U4978 ( .A(n747), .B(n5327), .Z(n5326) );
  XOR U4979 ( .A(n5328), .B(n5325), .Z(n5327) );
  XNOR U4980 ( .A(n5143), .B(n5321), .Z(n5323) );
  XOR U4981 ( .A(n5329), .B(n5330), .Z(n5143) );
  AND U4982 ( .A(n745), .B(n5331), .Z(n5330) );
  XOR U4983 ( .A(n5332), .B(n5329), .Z(n5331) );
  XOR U4984 ( .A(n5333), .B(n5334), .Z(n5321) );
  AND U4985 ( .A(n5335), .B(n5336), .Z(n5334) );
  XNOR U4986 ( .A(n5337), .B(n5159), .Z(n5336) );
  XOR U4987 ( .A(n5338), .B(n5339), .Z(n5159) );
  AND U4988 ( .A(n747), .B(n5340), .Z(n5339) );
  XOR U4989 ( .A(n5338), .B(n5341), .Z(n5340) );
  XNOR U4990 ( .A(n5156), .B(n5333), .Z(n5335) );
  XOR U4991 ( .A(n5342), .B(n5343), .Z(n5156) );
  AND U4992 ( .A(n745), .B(n5344), .Z(n5343) );
  XOR U4993 ( .A(n5342), .B(n5345), .Z(n5344) );
  IV U4994 ( .A(n5337), .Z(n5333) );
  AND U4995 ( .A(n5164), .B(n5167), .Z(n5337) );
  XNOR U4996 ( .A(n5346), .B(n5347), .Z(n5167) );
  AND U4997 ( .A(n747), .B(n5348), .Z(n5347) );
  XNOR U4998 ( .A(n5349), .B(n5346), .Z(n5348) );
  XOR U4999 ( .A(n5350), .B(n5351), .Z(n747) );
  AND U5000 ( .A(n5352), .B(n5353), .Z(n5351) );
  XNOR U5001 ( .A(n5173), .B(n5350), .Z(n5353) );
  AND U5002 ( .A(n5354), .B(n5355), .Z(n5173) );
  XOR U5003 ( .A(n5350), .B(n5174), .Z(n5352) );
  AND U5004 ( .A(n5356), .B(n5357), .Z(n5174) );
  XOR U5005 ( .A(n5358), .B(n5359), .Z(n5350) );
  AND U5006 ( .A(n5360), .B(n5361), .Z(n5359) );
  XOR U5007 ( .A(n5358), .B(n5184), .Z(n5361) );
  XOR U5008 ( .A(n5362), .B(n5363), .Z(n5184) );
  AND U5009 ( .A(n387), .B(n5364), .Z(n5363) );
  XOR U5010 ( .A(n5365), .B(n5362), .Z(n5364) );
  XNOR U5011 ( .A(n5181), .B(n5358), .Z(n5360) );
  XOR U5012 ( .A(n5366), .B(n5367), .Z(n5181) );
  AND U5013 ( .A(n385), .B(n5368), .Z(n5367) );
  XOR U5014 ( .A(n5369), .B(n5366), .Z(n5368) );
  XOR U5015 ( .A(n5370), .B(n5371), .Z(n5358) );
  AND U5016 ( .A(n5372), .B(n5373), .Z(n5371) );
  XOR U5017 ( .A(n5370), .B(n5196), .Z(n5373) );
  XOR U5018 ( .A(n5374), .B(n5375), .Z(n5196) );
  AND U5019 ( .A(n387), .B(n5376), .Z(n5375) );
  XOR U5020 ( .A(n5377), .B(n5374), .Z(n5376) );
  XNOR U5021 ( .A(n5193), .B(n5370), .Z(n5372) );
  XOR U5022 ( .A(n5378), .B(n5379), .Z(n5193) );
  AND U5023 ( .A(n385), .B(n5380), .Z(n5379) );
  XOR U5024 ( .A(n5381), .B(n5378), .Z(n5380) );
  XOR U5025 ( .A(n5382), .B(n5383), .Z(n5370) );
  AND U5026 ( .A(n5384), .B(n5385), .Z(n5383) );
  XOR U5027 ( .A(n5382), .B(n5208), .Z(n5385) );
  XOR U5028 ( .A(n5386), .B(n5387), .Z(n5208) );
  AND U5029 ( .A(n387), .B(n5388), .Z(n5387) );
  XOR U5030 ( .A(n5389), .B(n5386), .Z(n5388) );
  XNOR U5031 ( .A(n5205), .B(n5382), .Z(n5384) );
  XOR U5032 ( .A(n5390), .B(n5391), .Z(n5205) );
  AND U5033 ( .A(n385), .B(n5392), .Z(n5391) );
  XOR U5034 ( .A(n5393), .B(n5390), .Z(n5392) );
  XOR U5035 ( .A(n5394), .B(n5395), .Z(n5382) );
  AND U5036 ( .A(n5396), .B(n5397), .Z(n5395) );
  XOR U5037 ( .A(n5394), .B(n5220), .Z(n5397) );
  XOR U5038 ( .A(n5398), .B(n5399), .Z(n5220) );
  AND U5039 ( .A(n387), .B(n5400), .Z(n5399) );
  XOR U5040 ( .A(n5401), .B(n5398), .Z(n5400) );
  XNOR U5041 ( .A(n5217), .B(n5394), .Z(n5396) );
  XOR U5042 ( .A(n5402), .B(n5403), .Z(n5217) );
  AND U5043 ( .A(n385), .B(n5404), .Z(n5403) );
  XOR U5044 ( .A(n5405), .B(n5402), .Z(n5404) );
  XOR U5045 ( .A(n5406), .B(n5407), .Z(n5394) );
  AND U5046 ( .A(n5408), .B(n5409), .Z(n5407) );
  XOR U5047 ( .A(n5406), .B(n5232), .Z(n5409) );
  XOR U5048 ( .A(n5410), .B(n5411), .Z(n5232) );
  AND U5049 ( .A(n387), .B(n5412), .Z(n5411) );
  XOR U5050 ( .A(n5413), .B(n5410), .Z(n5412) );
  XNOR U5051 ( .A(n5229), .B(n5406), .Z(n5408) );
  XOR U5052 ( .A(n5414), .B(n5415), .Z(n5229) );
  AND U5053 ( .A(n385), .B(n5416), .Z(n5415) );
  XOR U5054 ( .A(n5417), .B(n5414), .Z(n5416) );
  XOR U5055 ( .A(n5418), .B(n5419), .Z(n5406) );
  AND U5056 ( .A(n5420), .B(n5421), .Z(n5419) );
  XOR U5057 ( .A(n5418), .B(n5244), .Z(n5421) );
  XOR U5058 ( .A(n5422), .B(n5423), .Z(n5244) );
  AND U5059 ( .A(n387), .B(n5424), .Z(n5423) );
  XOR U5060 ( .A(n5425), .B(n5422), .Z(n5424) );
  XNOR U5061 ( .A(n5241), .B(n5418), .Z(n5420) );
  XOR U5062 ( .A(n5426), .B(n5427), .Z(n5241) );
  AND U5063 ( .A(n385), .B(n5428), .Z(n5427) );
  XOR U5064 ( .A(n5429), .B(n5426), .Z(n5428) );
  XOR U5065 ( .A(n5430), .B(n5431), .Z(n5418) );
  AND U5066 ( .A(n5432), .B(n5433), .Z(n5431) );
  XOR U5067 ( .A(n5430), .B(n5256), .Z(n5433) );
  XOR U5068 ( .A(n5434), .B(n5435), .Z(n5256) );
  AND U5069 ( .A(n387), .B(n5436), .Z(n5435) );
  XOR U5070 ( .A(n5437), .B(n5434), .Z(n5436) );
  XNOR U5071 ( .A(n5253), .B(n5430), .Z(n5432) );
  XOR U5072 ( .A(n5438), .B(n5439), .Z(n5253) );
  AND U5073 ( .A(n385), .B(n5440), .Z(n5439) );
  XOR U5074 ( .A(n5441), .B(n5438), .Z(n5440) );
  XOR U5075 ( .A(n5442), .B(n5443), .Z(n5430) );
  AND U5076 ( .A(n5444), .B(n5445), .Z(n5443) );
  XOR U5077 ( .A(n5442), .B(n5268), .Z(n5445) );
  XOR U5078 ( .A(n5446), .B(n5447), .Z(n5268) );
  AND U5079 ( .A(n387), .B(n5448), .Z(n5447) );
  XOR U5080 ( .A(n5449), .B(n5446), .Z(n5448) );
  XNOR U5081 ( .A(n5265), .B(n5442), .Z(n5444) );
  XOR U5082 ( .A(n5450), .B(n5451), .Z(n5265) );
  AND U5083 ( .A(n385), .B(n5452), .Z(n5451) );
  XOR U5084 ( .A(n5453), .B(n5450), .Z(n5452) );
  XOR U5085 ( .A(n5454), .B(n5455), .Z(n5442) );
  AND U5086 ( .A(n5456), .B(n5457), .Z(n5455) );
  XOR U5087 ( .A(n5454), .B(n5280), .Z(n5457) );
  XOR U5088 ( .A(n5458), .B(n5459), .Z(n5280) );
  AND U5089 ( .A(n387), .B(n5460), .Z(n5459) );
  XOR U5090 ( .A(n5461), .B(n5458), .Z(n5460) );
  XNOR U5091 ( .A(n5277), .B(n5454), .Z(n5456) );
  XOR U5092 ( .A(n5462), .B(n5463), .Z(n5277) );
  AND U5093 ( .A(n385), .B(n5464), .Z(n5463) );
  XOR U5094 ( .A(n5465), .B(n5462), .Z(n5464) );
  XOR U5095 ( .A(n5466), .B(n5467), .Z(n5454) );
  AND U5096 ( .A(n5468), .B(n5469), .Z(n5467) );
  XOR U5097 ( .A(n5466), .B(n5292), .Z(n5469) );
  XOR U5098 ( .A(n5470), .B(n5471), .Z(n5292) );
  AND U5099 ( .A(n387), .B(n5472), .Z(n5471) );
  XOR U5100 ( .A(n5473), .B(n5470), .Z(n5472) );
  XNOR U5101 ( .A(n5289), .B(n5466), .Z(n5468) );
  XOR U5102 ( .A(n5474), .B(n5475), .Z(n5289) );
  AND U5103 ( .A(n385), .B(n5476), .Z(n5475) );
  XOR U5104 ( .A(n5477), .B(n5474), .Z(n5476) );
  XOR U5105 ( .A(n5478), .B(n5479), .Z(n5466) );
  AND U5106 ( .A(n5480), .B(n5481), .Z(n5479) );
  XOR U5107 ( .A(n5478), .B(n5304), .Z(n5481) );
  XOR U5108 ( .A(n5482), .B(n5483), .Z(n5304) );
  AND U5109 ( .A(n387), .B(n5484), .Z(n5483) );
  XOR U5110 ( .A(n5485), .B(n5482), .Z(n5484) );
  XNOR U5111 ( .A(n5301), .B(n5478), .Z(n5480) );
  XOR U5112 ( .A(n5486), .B(n5487), .Z(n5301) );
  AND U5113 ( .A(n385), .B(n5488), .Z(n5487) );
  XOR U5114 ( .A(n5489), .B(n5486), .Z(n5488) );
  XOR U5115 ( .A(n5490), .B(n5491), .Z(n5478) );
  AND U5116 ( .A(n5492), .B(n5493), .Z(n5491) );
  XOR U5117 ( .A(n5490), .B(n5316), .Z(n5493) );
  XOR U5118 ( .A(n5494), .B(n5495), .Z(n5316) );
  AND U5119 ( .A(n387), .B(n5496), .Z(n5495) );
  XOR U5120 ( .A(n5497), .B(n5494), .Z(n5496) );
  XNOR U5121 ( .A(n5313), .B(n5490), .Z(n5492) );
  XOR U5122 ( .A(n5498), .B(n5499), .Z(n5313) );
  AND U5123 ( .A(n385), .B(n5500), .Z(n5499) );
  XOR U5124 ( .A(n5501), .B(n5498), .Z(n5500) );
  XOR U5125 ( .A(n5502), .B(n5503), .Z(n5490) );
  AND U5126 ( .A(n5504), .B(n5505), .Z(n5503) );
  XOR U5127 ( .A(n5502), .B(n5328), .Z(n5505) );
  XOR U5128 ( .A(n5506), .B(n5507), .Z(n5328) );
  AND U5129 ( .A(n387), .B(n5508), .Z(n5507) );
  XOR U5130 ( .A(n5509), .B(n5506), .Z(n5508) );
  XNOR U5131 ( .A(n5325), .B(n5502), .Z(n5504) );
  XOR U5132 ( .A(n5510), .B(n5511), .Z(n5325) );
  AND U5133 ( .A(n385), .B(n5512), .Z(n5511) );
  XOR U5134 ( .A(n5513), .B(n5510), .Z(n5512) );
  XOR U5135 ( .A(n5514), .B(n5515), .Z(n5502) );
  AND U5136 ( .A(n5516), .B(n5517), .Z(n5515) );
  XNOR U5137 ( .A(n5518), .B(n5341), .Z(n5517) );
  XOR U5138 ( .A(n5519), .B(n5520), .Z(n5341) );
  AND U5139 ( .A(n387), .B(n5521), .Z(n5520) );
  XOR U5140 ( .A(n5519), .B(n5522), .Z(n5521) );
  XNOR U5141 ( .A(n5338), .B(n5514), .Z(n5516) );
  XOR U5142 ( .A(n5523), .B(n5524), .Z(n5338) );
  AND U5143 ( .A(n385), .B(n5525), .Z(n5524) );
  XOR U5144 ( .A(n5523), .B(n5526), .Z(n5525) );
  IV U5145 ( .A(n5518), .Z(n5514) );
  AND U5146 ( .A(n5346), .B(n5349), .Z(n5518) );
  XNOR U5147 ( .A(n5527), .B(n5528), .Z(n5349) );
  AND U5148 ( .A(n387), .B(n5529), .Z(n5528) );
  XNOR U5149 ( .A(n5530), .B(n5527), .Z(n5529) );
  XOR U5150 ( .A(n5531), .B(n5532), .Z(n387) );
  AND U5151 ( .A(n5533), .B(n5534), .Z(n5532) );
  XNOR U5152 ( .A(n5354), .B(n5531), .Z(n5534) );
  AND U5153 ( .A(p_input[3583]), .B(p_input[3567]), .Z(n5354) );
  XOR U5154 ( .A(n5531), .B(n5355), .Z(n5533) );
  AND U5155 ( .A(p_input[3551]), .B(p_input[3535]), .Z(n5355) );
  XOR U5156 ( .A(n5535), .B(n5536), .Z(n5531) );
  AND U5157 ( .A(n5537), .B(n5538), .Z(n5536) );
  XOR U5158 ( .A(n5535), .B(n5365), .Z(n5538) );
  XNOR U5159 ( .A(p_input[3566]), .B(n5539), .Z(n5365) );
  AND U5160 ( .A(n167), .B(n5540), .Z(n5539) );
  XOR U5161 ( .A(p_input[3582]), .B(p_input[3566]), .Z(n5540) );
  XNOR U5162 ( .A(n5362), .B(n5535), .Z(n5537) );
  XOR U5163 ( .A(n5541), .B(n5542), .Z(n5362) );
  AND U5164 ( .A(n165), .B(n5543), .Z(n5542) );
  XOR U5165 ( .A(p_input[3550]), .B(p_input[3534]), .Z(n5543) );
  XOR U5166 ( .A(n5544), .B(n5545), .Z(n5535) );
  AND U5167 ( .A(n5546), .B(n5547), .Z(n5545) );
  XOR U5168 ( .A(n5544), .B(n5377), .Z(n5547) );
  XNOR U5169 ( .A(p_input[3565]), .B(n5548), .Z(n5377) );
  AND U5170 ( .A(n167), .B(n5549), .Z(n5548) );
  XOR U5171 ( .A(p_input[3581]), .B(p_input[3565]), .Z(n5549) );
  XNOR U5172 ( .A(n5374), .B(n5544), .Z(n5546) );
  XOR U5173 ( .A(n5550), .B(n5551), .Z(n5374) );
  AND U5174 ( .A(n165), .B(n5552), .Z(n5551) );
  XOR U5175 ( .A(p_input[3549]), .B(p_input[3533]), .Z(n5552) );
  XOR U5176 ( .A(n5553), .B(n5554), .Z(n5544) );
  AND U5177 ( .A(n5555), .B(n5556), .Z(n5554) );
  XOR U5178 ( .A(n5553), .B(n5389), .Z(n5556) );
  XNOR U5179 ( .A(p_input[3564]), .B(n5557), .Z(n5389) );
  AND U5180 ( .A(n167), .B(n5558), .Z(n5557) );
  XOR U5181 ( .A(p_input[3580]), .B(p_input[3564]), .Z(n5558) );
  XNOR U5182 ( .A(n5386), .B(n5553), .Z(n5555) );
  XOR U5183 ( .A(n5559), .B(n5560), .Z(n5386) );
  AND U5184 ( .A(n165), .B(n5561), .Z(n5560) );
  XOR U5185 ( .A(p_input[3548]), .B(p_input[3532]), .Z(n5561) );
  XOR U5186 ( .A(n5562), .B(n5563), .Z(n5553) );
  AND U5187 ( .A(n5564), .B(n5565), .Z(n5563) );
  XOR U5188 ( .A(n5562), .B(n5401), .Z(n5565) );
  XNOR U5189 ( .A(p_input[3563]), .B(n5566), .Z(n5401) );
  AND U5190 ( .A(n167), .B(n5567), .Z(n5566) );
  XOR U5191 ( .A(p_input[3579]), .B(p_input[3563]), .Z(n5567) );
  XNOR U5192 ( .A(n5398), .B(n5562), .Z(n5564) );
  XOR U5193 ( .A(n5568), .B(n5569), .Z(n5398) );
  AND U5194 ( .A(n165), .B(n5570), .Z(n5569) );
  XOR U5195 ( .A(p_input[3547]), .B(p_input[3531]), .Z(n5570) );
  XOR U5196 ( .A(n5571), .B(n5572), .Z(n5562) );
  AND U5197 ( .A(n5573), .B(n5574), .Z(n5572) );
  XOR U5198 ( .A(n5571), .B(n5413), .Z(n5574) );
  XNOR U5199 ( .A(p_input[3562]), .B(n5575), .Z(n5413) );
  AND U5200 ( .A(n167), .B(n5576), .Z(n5575) );
  XOR U5201 ( .A(p_input[3578]), .B(p_input[3562]), .Z(n5576) );
  XNOR U5202 ( .A(n5410), .B(n5571), .Z(n5573) );
  XOR U5203 ( .A(n5577), .B(n5578), .Z(n5410) );
  AND U5204 ( .A(n165), .B(n5579), .Z(n5578) );
  XOR U5205 ( .A(p_input[3546]), .B(p_input[3530]), .Z(n5579) );
  XOR U5206 ( .A(n5580), .B(n5581), .Z(n5571) );
  AND U5207 ( .A(n5582), .B(n5583), .Z(n5581) );
  XOR U5208 ( .A(n5580), .B(n5425), .Z(n5583) );
  XNOR U5209 ( .A(p_input[3561]), .B(n5584), .Z(n5425) );
  AND U5210 ( .A(n167), .B(n5585), .Z(n5584) );
  XOR U5211 ( .A(p_input[3577]), .B(p_input[3561]), .Z(n5585) );
  XNOR U5212 ( .A(n5422), .B(n5580), .Z(n5582) );
  XOR U5213 ( .A(n5586), .B(n5587), .Z(n5422) );
  AND U5214 ( .A(n165), .B(n5588), .Z(n5587) );
  XOR U5215 ( .A(p_input[3545]), .B(p_input[3529]), .Z(n5588) );
  XOR U5216 ( .A(n5589), .B(n5590), .Z(n5580) );
  AND U5217 ( .A(n5591), .B(n5592), .Z(n5590) );
  XOR U5218 ( .A(n5589), .B(n5437), .Z(n5592) );
  XNOR U5219 ( .A(p_input[3560]), .B(n5593), .Z(n5437) );
  AND U5220 ( .A(n167), .B(n5594), .Z(n5593) );
  XOR U5221 ( .A(p_input[3576]), .B(p_input[3560]), .Z(n5594) );
  XNOR U5222 ( .A(n5434), .B(n5589), .Z(n5591) );
  XOR U5223 ( .A(n5595), .B(n5596), .Z(n5434) );
  AND U5224 ( .A(n165), .B(n5597), .Z(n5596) );
  XOR U5225 ( .A(p_input[3544]), .B(p_input[3528]), .Z(n5597) );
  XOR U5226 ( .A(n5598), .B(n5599), .Z(n5589) );
  AND U5227 ( .A(n5600), .B(n5601), .Z(n5599) );
  XOR U5228 ( .A(n5598), .B(n5449), .Z(n5601) );
  XNOR U5229 ( .A(p_input[3559]), .B(n5602), .Z(n5449) );
  AND U5230 ( .A(n167), .B(n5603), .Z(n5602) );
  XOR U5231 ( .A(p_input[3575]), .B(p_input[3559]), .Z(n5603) );
  XNOR U5232 ( .A(n5446), .B(n5598), .Z(n5600) );
  XOR U5233 ( .A(n5604), .B(n5605), .Z(n5446) );
  AND U5234 ( .A(n165), .B(n5606), .Z(n5605) );
  XOR U5235 ( .A(p_input[3543]), .B(p_input[3527]), .Z(n5606) );
  XOR U5236 ( .A(n5607), .B(n5608), .Z(n5598) );
  AND U5237 ( .A(n5609), .B(n5610), .Z(n5608) );
  XOR U5238 ( .A(n5607), .B(n5461), .Z(n5610) );
  XNOR U5239 ( .A(p_input[3558]), .B(n5611), .Z(n5461) );
  AND U5240 ( .A(n167), .B(n5612), .Z(n5611) );
  XOR U5241 ( .A(p_input[3574]), .B(p_input[3558]), .Z(n5612) );
  XNOR U5242 ( .A(n5458), .B(n5607), .Z(n5609) );
  XOR U5243 ( .A(n5613), .B(n5614), .Z(n5458) );
  AND U5244 ( .A(n165), .B(n5615), .Z(n5614) );
  XOR U5245 ( .A(p_input[3542]), .B(p_input[3526]), .Z(n5615) );
  XOR U5246 ( .A(n5616), .B(n5617), .Z(n5607) );
  AND U5247 ( .A(n5618), .B(n5619), .Z(n5617) );
  XOR U5248 ( .A(n5616), .B(n5473), .Z(n5619) );
  XNOR U5249 ( .A(p_input[3557]), .B(n5620), .Z(n5473) );
  AND U5250 ( .A(n167), .B(n5621), .Z(n5620) );
  XOR U5251 ( .A(p_input[3573]), .B(p_input[3557]), .Z(n5621) );
  XNOR U5252 ( .A(n5470), .B(n5616), .Z(n5618) );
  XOR U5253 ( .A(n5622), .B(n5623), .Z(n5470) );
  AND U5254 ( .A(n165), .B(n5624), .Z(n5623) );
  XOR U5255 ( .A(p_input[3541]), .B(p_input[3525]), .Z(n5624) );
  XOR U5256 ( .A(n5625), .B(n5626), .Z(n5616) );
  AND U5257 ( .A(n5627), .B(n5628), .Z(n5626) );
  XOR U5258 ( .A(n5625), .B(n5485), .Z(n5628) );
  XNOR U5259 ( .A(p_input[3556]), .B(n5629), .Z(n5485) );
  AND U5260 ( .A(n167), .B(n5630), .Z(n5629) );
  XOR U5261 ( .A(p_input[3572]), .B(p_input[3556]), .Z(n5630) );
  XNOR U5262 ( .A(n5482), .B(n5625), .Z(n5627) );
  XOR U5263 ( .A(n5631), .B(n5632), .Z(n5482) );
  AND U5264 ( .A(n165), .B(n5633), .Z(n5632) );
  XOR U5265 ( .A(p_input[3540]), .B(p_input[3524]), .Z(n5633) );
  XOR U5266 ( .A(n5634), .B(n5635), .Z(n5625) );
  AND U5267 ( .A(n5636), .B(n5637), .Z(n5635) );
  XOR U5268 ( .A(n5634), .B(n5497), .Z(n5637) );
  XNOR U5269 ( .A(p_input[3555]), .B(n5638), .Z(n5497) );
  AND U5270 ( .A(n167), .B(n5639), .Z(n5638) );
  XOR U5271 ( .A(p_input[3571]), .B(p_input[3555]), .Z(n5639) );
  XNOR U5272 ( .A(n5494), .B(n5634), .Z(n5636) );
  XOR U5273 ( .A(n5640), .B(n5641), .Z(n5494) );
  AND U5274 ( .A(n165), .B(n5642), .Z(n5641) );
  XOR U5275 ( .A(p_input[3539]), .B(p_input[3523]), .Z(n5642) );
  XOR U5276 ( .A(n5643), .B(n5644), .Z(n5634) );
  AND U5277 ( .A(n5645), .B(n5646), .Z(n5644) );
  XOR U5278 ( .A(n5643), .B(n5509), .Z(n5646) );
  XNOR U5279 ( .A(p_input[3554]), .B(n5647), .Z(n5509) );
  AND U5280 ( .A(n167), .B(n5648), .Z(n5647) );
  XOR U5281 ( .A(p_input[3570]), .B(p_input[3554]), .Z(n5648) );
  XNOR U5282 ( .A(n5506), .B(n5643), .Z(n5645) );
  XOR U5283 ( .A(n5649), .B(n5650), .Z(n5506) );
  AND U5284 ( .A(n165), .B(n5651), .Z(n5650) );
  XOR U5285 ( .A(p_input[3538]), .B(p_input[3522]), .Z(n5651) );
  XOR U5286 ( .A(n5652), .B(n5653), .Z(n5643) );
  AND U5287 ( .A(n5654), .B(n5655), .Z(n5653) );
  XNOR U5288 ( .A(n5656), .B(n5522), .Z(n5655) );
  XNOR U5289 ( .A(p_input[3553]), .B(n5657), .Z(n5522) );
  AND U5290 ( .A(n167), .B(n5658), .Z(n5657) );
  XNOR U5291 ( .A(p_input[3569]), .B(n5659), .Z(n5658) );
  IV U5292 ( .A(p_input[3553]), .Z(n5659) );
  XNOR U5293 ( .A(n5519), .B(n5652), .Z(n5654) );
  XNOR U5294 ( .A(p_input[3521]), .B(n5660), .Z(n5519) );
  AND U5295 ( .A(n165), .B(n5661), .Z(n5660) );
  XOR U5296 ( .A(p_input[3537]), .B(p_input[3521]), .Z(n5661) );
  IV U5297 ( .A(n5656), .Z(n5652) );
  AND U5298 ( .A(n5527), .B(n5530), .Z(n5656) );
  XOR U5299 ( .A(p_input[3552]), .B(n5662), .Z(n5530) );
  AND U5300 ( .A(n167), .B(n5663), .Z(n5662) );
  XOR U5301 ( .A(p_input[3568]), .B(p_input[3552]), .Z(n5663) );
  XOR U5302 ( .A(n5664), .B(n5665), .Z(n167) );
  AND U5303 ( .A(n5666), .B(n5667), .Z(n5665) );
  XNOR U5304 ( .A(p_input[3583]), .B(n5664), .Z(n5667) );
  XOR U5305 ( .A(n5664), .B(p_input[3567]), .Z(n5666) );
  XOR U5306 ( .A(n5668), .B(n5669), .Z(n5664) );
  AND U5307 ( .A(n5670), .B(n5671), .Z(n5669) );
  XNOR U5308 ( .A(p_input[3582]), .B(n5668), .Z(n5671) );
  XOR U5309 ( .A(n5668), .B(p_input[3566]), .Z(n5670) );
  XOR U5310 ( .A(n5672), .B(n5673), .Z(n5668) );
  AND U5311 ( .A(n5674), .B(n5675), .Z(n5673) );
  XNOR U5312 ( .A(p_input[3581]), .B(n5672), .Z(n5675) );
  XOR U5313 ( .A(n5672), .B(p_input[3565]), .Z(n5674) );
  XOR U5314 ( .A(n5676), .B(n5677), .Z(n5672) );
  AND U5315 ( .A(n5678), .B(n5679), .Z(n5677) );
  XNOR U5316 ( .A(p_input[3580]), .B(n5676), .Z(n5679) );
  XOR U5317 ( .A(n5676), .B(p_input[3564]), .Z(n5678) );
  XOR U5318 ( .A(n5680), .B(n5681), .Z(n5676) );
  AND U5319 ( .A(n5682), .B(n5683), .Z(n5681) );
  XNOR U5320 ( .A(p_input[3579]), .B(n5680), .Z(n5683) );
  XOR U5321 ( .A(n5680), .B(p_input[3563]), .Z(n5682) );
  XOR U5322 ( .A(n5684), .B(n5685), .Z(n5680) );
  AND U5323 ( .A(n5686), .B(n5687), .Z(n5685) );
  XNOR U5324 ( .A(p_input[3578]), .B(n5684), .Z(n5687) );
  XOR U5325 ( .A(n5684), .B(p_input[3562]), .Z(n5686) );
  XOR U5326 ( .A(n5688), .B(n5689), .Z(n5684) );
  AND U5327 ( .A(n5690), .B(n5691), .Z(n5689) );
  XNOR U5328 ( .A(p_input[3577]), .B(n5688), .Z(n5691) );
  XOR U5329 ( .A(n5688), .B(p_input[3561]), .Z(n5690) );
  XOR U5330 ( .A(n5692), .B(n5693), .Z(n5688) );
  AND U5331 ( .A(n5694), .B(n5695), .Z(n5693) );
  XNOR U5332 ( .A(p_input[3576]), .B(n5692), .Z(n5695) );
  XOR U5333 ( .A(n5692), .B(p_input[3560]), .Z(n5694) );
  XOR U5334 ( .A(n5696), .B(n5697), .Z(n5692) );
  AND U5335 ( .A(n5698), .B(n5699), .Z(n5697) );
  XNOR U5336 ( .A(p_input[3575]), .B(n5696), .Z(n5699) );
  XOR U5337 ( .A(n5696), .B(p_input[3559]), .Z(n5698) );
  XOR U5338 ( .A(n5700), .B(n5701), .Z(n5696) );
  AND U5339 ( .A(n5702), .B(n5703), .Z(n5701) );
  XNOR U5340 ( .A(p_input[3574]), .B(n5700), .Z(n5703) );
  XOR U5341 ( .A(n5700), .B(p_input[3558]), .Z(n5702) );
  XOR U5342 ( .A(n5704), .B(n5705), .Z(n5700) );
  AND U5343 ( .A(n5706), .B(n5707), .Z(n5705) );
  XNOR U5344 ( .A(p_input[3573]), .B(n5704), .Z(n5707) );
  XOR U5345 ( .A(n5704), .B(p_input[3557]), .Z(n5706) );
  XOR U5346 ( .A(n5708), .B(n5709), .Z(n5704) );
  AND U5347 ( .A(n5710), .B(n5711), .Z(n5709) );
  XNOR U5348 ( .A(p_input[3572]), .B(n5708), .Z(n5711) );
  XOR U5349 ( .A(n5708), .B(p_input[3556]), .Z(n5710) );
  XOR U5350 ( .A(n5712), .B(n5713), .Z(n5708) );
  AND U5351 ( .A(n5714), .B(n5715), .Z(n5713) );
  XNOR U5352 ( .A(p_input[3571]), .B(n5712), .Z(n5715) );
  XOR U5353 ( .A(n5712), .B(p_input[3555]), .Z(n5714) );
  XOR U5354 ( .A(n5716), .B(n5717), .Z(n5712) );
  AND U5355 ( .A(n5718), .B(n5719), .Z(n5717) );
  XNOR U5356 ( .A(p_input[3570]), .B(n5716), .Z(n5719) );
  XOR U5357 ( .A(n5716), .B(p_input[3554]), .Z(n5718) );
  XNOR U5358 ( .A(n5720), .B(n5721), .Z(n5716) );
  AND U5359 ( .A(n5722), .B(n5723), .Z(n5721) );
  XOR U5360 ( .A(p_input[3569]), .B(n5720), .Z(n5723) );
  XNOR U5361 ( .A(p_input[3553]), .B(n5720), .Z(n5722) );
  AND U5362 ( .A(p_input[3568]), .B(n5724), .Z(n5720) );
  IV U5363 ( .A(p_input[3552]), .Z(n5724) );
  XNOR U5364 ( .A(p_input[3520]), .B(n5725), .Z(n5527) );
  AND U5365 ( .A(n165), .B(n5726), .Z(n5725) );
  XOR U5366 ( .A(p_input[3536]), .B(p_input[3520]), .Z(n5726) );
  XOR U5367 ( .A(n5727), .B(n5728), .Z(n165) );
  AND U5368 ( .A(n5729), .B(n5730), .Z(n5728) );
  XNOR U5369 ( .A(p_input[3551]), .B(n5727), .Z(n5730) );
  XOR U5370 ( .A(n5727), .B(p_input[3535]), .Z(n5729) );
  XOR U5371 ( .A(n5731), .B(n5732), .Z(n5727) );
  AND U5372 ( .A(n5733), .B(n5734), .Z(n5732) );
  XNOR U5373 ( .A(p_input[3550]), .B(n5731), .Z(n5734) );
  XNOR U5374 ( .A(n5731), .B(n5541), .Z(n5733) );
  IV U5375 ( .A(p_input[3534]), .Z(n5541) );
  XOR U5376 ( .A(n5735), .B(n5736), .Z(n5731) );
  AND U5377 ( .A(n5737), .B(n5738), .Z(n5736) );
  XNOR U5378 ( .A(p_input[3549]), .B(n5735), .Z(n5738) );
  XNOR U5379 ( .A(n5735), .B(n5550), .Z(n5737) );
  IV U5380 ( .A(p_input[3533]), .Z(n5550) );
  XOR U5381 ( .A(n5739), .B(n5740), .Z(n5735) );
  AND U5382 ( .A(n5741), .B(n5742), .Z(n5740) );
  XNOR U5383 ( .A(p_input[3548]), .B(n5739), .Z(n5742) );
  XNOR U5384 ( .A(n5739), .B(n5559), .Z(n5741) );
  IV U5385 ( .A(p_input[3532]), .Z(n5559) );
  XOR U5386 ( .A(n5743), .B(n5744), .Z(n5739) );
  AND U5387 ( .A(n5745), .B(n5746), .Z(n5744) );
  XNOR U5388 ( .A(p_input[3547]), .B(n5743), .Z(n5746) );
  XNOR U5389 ( .A(n5743), .B(n5568), .Z(n5745) );
  IV U5390 ( .A(p_input[3531]), .Z(n5568) );
  XOR U5391 ( .A(n5747), .B(n5748), .Z(n5743) );
  AND U5392 ( .A(n5749), .B(n5750), .Z(n5748) );
  XNOR U5393 ( .A(p_input[3546]), .B(n5747), .Z(n5750) );
  XNOR U5394 ( .A(n5747), .B(n5577), .Z(n5749) );
  IV U5395 ( .A(p_input[3530]), .Z(n5577) );
  XOR U5396 ( .A(n5751), .B(n5752), .Z(n5747) );
  AND U5397 ( .A(n5753), .B(n5754), .Z(n5752) );
  XNOR U5398 ( .A(p_input[3545]), .B(n5751), .Z(n5754) );
  XNOR U5399 ( .A(n5751), .B(n5586), .Z(n5753) );
  IV U5400 ( .A(p_input[3529]), .Z(n5586) );
  XOR U5401 ( .A(n5755), .B(n5756), .Z(n5751) );
  AND U5402 ( .A(n5757), .B(n5758), .Z(n5756) );
  XNOR U5403 ( .A(p_input[3544]), .B(n5755), .Z(n5758) );
  XNOR U5404 ( .A(n5755), .B(n5595), .Z(n5757) );
  IV U5405 ( .A(p_input[3528]), .Z(n5595) );
  XOR U5406 ( .A(n5759), .B(n5760), .Z(n5755) );
  AND U5407 ( .A(n5761), .B(n5762), .Z(n5760) );
  XNOR U5408 ( .A(p_input[3543]), .B(n5759), .Z(n5762) );
  XNOR U5409 ( .A(n5759), .B(n5604), .Z(n5761) );
  IV U5410 ( .A(p_input[3527]), .Z(n5604) );
  XOR U5411 ( .A(n5763), .B(n5764), .Z(n5759) );
  AND U5412 ( .A(n5765), .B(n5766), .Z(n5764) );
  XNOR U5413 ( .A(p_input[3542]), .B(n5763), .Z(n5766) );
  XNOR U5414 ( .A(n5763), .B(n5613), .Z(n5765) );
  IV U5415 ( .A(p_input[3526]), .Z(n5613) );
  XOR U5416 ( .A(n5767), .B(n5768), .Z(n5763) );
  AND U5417 ( .A(n5769), .B(n5770), .Z(n5768) );
  XNOR U5418 ( .A(p_input[3541]), .B(n5767), .Z(n5770) );
  XNOR U5419 ( .A(n5767), .B(n5622), .Z(n5769) );
  IV U5420 ( .A(p_input[3525]), .Z(n5622) );
  XOR U5421 ( .A(n5771), .B(n5772), .Z(n5767) );
  AND U5422 ( .A(n5773), .B(n5774), .Z(n5772) );
  XNOR U5423 ( .A(p_input[3540]), .B(n5771), .Z(n5774) );
  XNOR U5424 ( .A(n5771), .B(n5631), .Z(n5773) );
  IV U5425 ( .A(p_input[3524]), .Z(n5631) );
  XOR U5426 ( .A(n5775), .B(n5776), .Z(n5771) );
  AND U5427 ( .A(n5777), .B(n5778), .Z(n5776) );
  XNOR U5428 ( .A(p_input[3539]), .B(n5775), .Z(n5778) );
  XNOR U5429 ( .A(n5775), .B(n5640), .Z(n5777) );
  IV U5430 ( .A(p_input[3523]), .Z(n5640) );
  XOR U5431 ( .A(n5779), .B(n5780), .Z(n5775) );
  AND U5432 ( .A(n5781), .B(n5782), .Z(n5780) );
  XNOR U5433 ( .A(p_input[3538]), .B(n5779), .Z(n5782) );
  XNOR U5434 ( .A(n5779), .B(n5649), .Z(n5781) );
  IV U5435 ( .A(p_input[3522]), .Z(n5649) );
  XNOR U5436 ( .A(n5783), .B(n5784), .Z(n5779) );
  AND U5437 ( .A(n5785), .B(n5786), .Z(n5784) );
  XOR U5438 ( .A(p_input[3537]), .B(n5783), .Z(n5786) );
  XNOR U5439 ( .A(p_input[3521]), .B(n5783), .Z(n5785) );
  AND U5440 ( .A(p_input[3536]), .B(n5787), .Z(n5783) );
  IV U5441 ( .A(p_input[3520]), .Z(n5787) );
  XOR U5442 ( .A(n5788), .B(n5789), .Z(n5346) );
  AND U5443 ( .A(n385), .B(n5790), .Z(n5789) );
  XNOR U5444 ( .A(n5791), .B(n5788), .Z(n5790) );
  XOR U5445 ( .A(n5792), .B(n5793), .Z(n385) );
  AND U5446 ( .A(n5794), .B(n5795), .Z(n5793) );
  XNOR U5447 ( .A(n5356), .B(n5792), .Z(n5795) );
  AND U5448 ( .A(p_input[3519]), .B(p_input[3503]), .Z(n5356) );
  XOR U5449 ( .A(n5792), .B(n5357), .Z(n5794) );
  AND U5450 ( .A(p_input[3487]), .B(p_input[3471]), .Z(n5357) );
  XOR U5451 ( .A(n5796), .B(n5797), .Z(n5792) );
  AND U5452 ( .A(n5798), .B(n5799), .Z(n5797) );
  XOR U5453 ( .A(n5796), .B(n5369), .Z(n5799) );
  XNOR U5454 ( .A(p_input[3502]), .B(n5800), .Z(n5369) );
  AND U5455 ( .A(n171), .B(n5801), .Z(n5800) );
  XOR U5456 ( .A(p_input[3518]), .B(p_input[3502]), .Z(n5801) );
  XNOR U5457 ( .A(n5366), .B(n5796), .Z(n5798) );
  XOR U5458 ( .A(n5802), .B(n5803), .Z(n5366) );
  AND U5459 ( .A(n168), .B(n5804), .Z(n5803) );
  XOR U5460 ( .A(p_input[3486]), .B(p_input[3470]), .Z(n5804) );
  XOR U5461 ( .A(n5805), .B(n5806), .Z(n5796) );
  AND U5462 ( .A(n5807), .B(n5808), .Z(n5806) );
  XOR U5463 ( .A(n5805), .B(n5381), .Z(n5808) );
  XNOR U5464 ( .A(p_input[3501]), .B(n5809), .Z(n5381) );
  AND U5465 ( .A(n171), .B(n5810), .Z(n5809) );
  XOR U5466 ( .A(p_input[3517]), .B(p_input[3501]), .Z(n5810) );
  XNOR U5467 ( .A(n5378), .B(n5805), .Z(n5807) );
  XOR U5468 ( .A(n5811), .B(n5812), .Z(n5378) );
  AND U5469 ( .A(n168), .B(n5813), .Z(n5812) );
  XOR U5470 ( .A(p_input[3485]), .B(p_input[3469]), .Z(n5813) );
  XOR U5471 ( .A(n5814), .B(n5815), .Z(n5805) );
  AND U5472 ( .A(n5816), .B(n5817), .Z(n5815) );
  XOR U5473 ( .A(n5814), .B(n5393), .Z(n5817) );
  XNOR U5474 ( .A(p_input[3500]), .B(n5818), .Z(n5393) );
  AND U5475 ( .A(n171), .B(n5819), .Z(n5818) );
  XOR U5476 ( .A(p_input[3516]), .B(p_input[3500]), .Z(n5819) );
  XNOR U5477 ( .A(n5390), .B(n5814), .Z(n5816) );
  XOR U5478 ( .A(n5820), .B(n5821), .Z(n5390) );
  AND U5479 ( .A(n168), .B(n5822), .Z(n5821) );
  XOR U5480 ( .A(p_input[3484]), .B(p_input[3468]), .Z(n5822) );
  XOR U5481 ( .A(n5823), .B(n5824), .Z(n5814) );
  AND U5482 ( .A(n5825), .B(n5826), .Z(n5824) );
  XOR U5483 ( .A(n5823), .B(n5405), .Z(n5826) );
  XNOR U5484 ( .A(p_input[3499]), .B(n5827), .Z(n5405) );
  AND U5485 ( .A(n171), .B(n5828), .Z(n5827) );
  XOR U5486 ( .A(p_input[3515]), .B(p_input[3499]), .Z(n5828) );
  XNOR U5487 ( .A(n5402), .B(n5823), .Z(n5825) );
  XOR U5488 ( .A(n5829), .B(n5830), .Z(n5402) );
  AND U5489 ( .A(n168), .B(n5831), .Z(n5830) );
  XOR U5490 ( .A(p_input[3483]), .B(p_input[3467]), .Z(n5831) );
  XOR U5491 ( .A(n5832), .B(n5833), .Z(n5823) );
  AND U5492 ( .A(n5834), .B(n5835), .Z(n5833) );
  XOR U5493 ( .A(n5832), .B(n5417), .Z(n5835) );
  XNOR U5494 ( .A(p_input[3498]), .B(n5836), .Z(n5417) );
  AND U5495 ( .A(n171), .B(n5837), .Z(n5836) );
  XOR U5496 ( .A(p_input[3514]), .B(p_input[3498]), .Z(n5837) );
  XNOR U5497 ( .A(n5414), .B(n5832), .Z(n5834) );
  XOR U5498 ( .A(n5838), .B(n5839), .Z(n5414) );
  AND U5499 ( .A(n168), .B(n5840), .Z(n5839) );
  XOR U5500 ( .A(p_input[3482]), .B(p_input[3466]), .Z(n5840) );
  XOR U5501 ( .A(n5841), .B(n5842), .Z(n5832) );
  AND U5502 ( .A(n5843), .B(n5844), .Z(n5842) );
  XOR U5503 ( .A(n5841), .B(n5429), .Z(n5844) );
  XNOR U5504 ( .A(p_input[3497]), .B(n5845), .Z(n5429) );
  AND U5505 ( .A(n171), .B(n5846), .Z(n5845) );
  XOR U5506 ( .A(p_input[3513]), .B(p_input[3497]), .Z(n5846) );
  XNOR U5507 ( .A(n5426), .B(n5841), .Z(n5843) );
  XOR U5508 ( .A(n5847), .B(n5848), .Z(n5426) );
  AND U5509 ( .A(n168), .B(n5849), .Z(n5848) );
  XOR U5510 ( .A(p_input[3481]), .B(p_input[3465]), .Z(n5849) );
  XOR U5511 ( .A(n5850), .B(n5851), .Z(n5841) );
  AND U5512 ( .A(n5852), .B(n5853), .Z(n5851) );
  XOR U5513 ( .A(n5850), .B(n5441), .Z(n5853) );
  XNOR U5514 ( .A(p_input[3496]), .B(n5854), .Z(n5441) );
  AND U5515 ( .A(n171), .B(n5855), .Z(n5854) );
  XOR U5516 ( .A(p_input[3512]), .B(p_input[3496]), .Z(n5855) );
  XNOR U5517 ( .A(n5438), .B(n5850), .Z(n5852) );
  XOR U5518 ( .A(n5856), .B(n5857), .Z(n5438) );
  AND U5519 ( .A(n168), .B(n5858), .Z(n5857) );
  XOR U5520 ( .A(p_input[3480]), .B(p_input[3464]), .Z(n5858) );
  XOR U5521 ( .A(n5859), .B(n5860), .Z(n5850) );
  AND U5522 ( .A(n5861), .B(n5862), .Z(n5860) );
  XOR U5523 ( .A(n5859), .B(n5453), .Z(n5862) );
  XNOR U5524 ( .A(p_input[3495]), .B(n5863), .Z(n5453) );
  AND U5525 ( .A(n171), .B(n5864), .Z(n5863) );
  XOR U5526 ( .A(p_input[3511]), .B(p_input[3495]), .Z(n5864) );
  XNOR U5527 ( .A(n5450), .B(n5859), .Z(n5861) );
  XOR U5528 ( .A(n5865), .B(n5866), .Z(n5450) );
  AND U5529 ( .A(n168), .B(n5867), .Z(n5866) );
  XOR U5530 ( .A(p_input[3479]), .B(p_input[3463]), .Z(n5867) );
  XOR U5531 ( .A(n5868), .B(n5869), .Z(n5859) );
  AND U5532 ( .A(n5870), .B(n5871), .Z(n5869) );
  XOR U5533 ( .A(n5868), .B(n5465), .Z(n5871) );
  XNOR U5534 ( .A(p_input[3494]), .B(n5872), .Z(n5465) );
  AND U5535 ( .A(n171), .B(n5873), .Z(n5872) );
  XOR U5536 ( .A(p_input[3510]), .B(p_input[3494]), .Z(n5873) );
  XNOR U5537 ( .A(n5462), .B(n5868), .Z(n5870) );
  XOR U5538 ( .A(n5874), .B(n5875), .Z(n5462) );
  AND U5539 ( .A(n168), .B(n5876), .Z(n5875) );
  XOR U5540 ( .A(p_input[3478]), .B(p_input[3462]), .Z(n5876) );
  XOR U5541 ( .A(n5877), .B(n5878), .Z(n5868) );
  AND U5542 ( .A(n5879), .B(n5880), .Z(n5878) );
  XOR U5543 ( .A(n5877), .B(n5477), .Z(n5880) );
  XNOR U5544 ( .A(p_input[3493]), .B(n5881), .Z(n5477) );
  AND U5545 ( .A(n171), .B(n5882), .Z(n5881) );
  XOR U5546 ( .A(p_input[3509]), .B(p_input[3493]), .Z(n5882) );
  XNOR U5547 ( .A(n5474), .B(n5877), .Z(n5879) );
  XOR U5548 ( .A(n5883), .B(n5884), .Z(n5474) );
  AND U5549 ( .A(n168), .B(n5885), .Z(n5884) );
  XOR U5550 ( .A(p_input[3477]), .B(p_input[3461]), .Z(n5885) );
  XOR U5551 ( .A(n5886), .B(n5887), .Z(n5877) );
  AND U5552 ( .A(n5888), .B(n5889), .Z(n5887) );
  XOR U5553 ( .A(n5886), .B(n5489), .Z(n5889) );
  XNOR U5554 ( .A(p_input[3492]), .B(n5890), .Z(n5489) );
  AND U5555 ( .A(n171), .B(n5891), .Z(n5890) );
  XOR U5556 ( .A(p_input[3508]), .B(p_input[3492]), .Z(n5891) );
  XNOR U5557 ( .A(n5486), .B(n5886), .Z(n5888) );
  XOR U5558 ( .A(n5892), .B(n5893), .Z(n5486) );
  AND U5559 ( .A(n168), .B(n5894), .Z(n5893) );
  XOR U5560 ( .A(p_input[3476]), .B(p_input[3460]), .Z(n5894) );
  XOR U5561 ( .A(n5895), .B(n5896), .Z(n5886) );
  AND U5562 ( .A(n5897), .B(n5898), .Z(n5896) );
  XOR U5563 ( .A(n5895), .B(n5501), .Z(n5898) );
  XNOR U5564 ( .A(p_input[3491]), .B(n5899), .Z(n5501) );
  AND U5565 ( .A(n171), .B(n5900), .Z(n5899) );
  XOR U5566 ( .A(p_input[3507]), .B(p_input[3491]), .Z(n5900) );
  XNOR U5567 ( .A(n5498), .B(n5895), .Z(n5897) );
  XOR U5568 ( .A(n5901), .B(n5902), .Z(n5498) );
  AND U5569 ( .A(n168), .B(n5903), .Z(n5902) );
  XOR U5570 ( .A(p_input[3475]), .B(p_input[3459]), .Z(n5903) );
  XOR U5571 ( .A(n5904), .B(n5905), .Z(n5895) );
  AND U5572 ( .A(n5906), .B(n5907), .Z(n5905) );
  XOR U5573 ( .A(n5904), .B(n5513), .Z(n5907) );
  XNOR U5574 ( .A(p_input[3490]), .B(n5908), .Z(n5513) );
  AND U5575 ( .A(n171), .B(n5909), .Z(n5908) );
  XOR U5576 ( .A(p_input[3506]), .B(p_input[3490]), .Z(n5909) );
  XNOR U5577 ( .A(n5510), .B(n5904), .Z(n5906) );
  XOR U5578 ( .A(n5910), .B(n5911), .Z(n5510) );
  AND U5579 ( .A(n168), .B(n5912), .Z(n5911) );
  XOR U5580 ( .A(p_input[3474]), .B(p_input[3458]), .Z(n5912) );
  XOR U5581 ( .A(n5913), .B(n5914), .Z(n5904) );
  AND U5582 ( .A(n5915), .B(n5916), .Z(n5914) );
  XNOR U5583 ( .A(n5917), .B(n5526), .Z(n5916) );
  XNOR U5584 ( .A(p_input[3489]), .B(n5918), .Z(n5526) );
  AND U5585 ( .A(n171), .B(n5919), .Z(n5918) );
  XNOR U5586 ( .A(p_input[3505]), .B(n5920), .Z(n5919) );
  IV U5587 ( .A(p_input[3489]), .Z(n5920) );
  XNOR U5588 ( .A(n5523), .B(n5913), .Z(n5915) );
  XNOR U5589 ( .A(p_input[3457]), .B(n5921), .Z(n5523) );
  AND U5590 ( .A(n168), .B(n5922), .Z(n5921) );
  XOR U5591 ( .A(p_input[3473]), .B(p_input[3457]), .Z(n5922) );
  IV U5592 ( .A(n5917), .Z(n5913) );
  AND U5593 ( .A(n5788), .B(n5791), .Z(n5917) );
  XOR U5594 ( .A(p_input[3488]), .B(n5923), .Z(n5791) );
  AND U5595 ( .A(n171), .B(n5924), .Z(n5923) );
  XOR U5596 ( .A(p_input[3504]), .B(p_input[3488]), .Z(n5924) );
  XOR U5597 ( .A(n5925), .B(n5926), .Z(n171) );
  AND U5598 ( .A(n5927), .B(n5928), .Z(n5926) );
  XNOR U5599 ( .A(p_input[3519]), .B(n5925), .Z(n5928) );
  XOR U5600 ( .A(n5925), .B(p_input[3503]), .Z(n5927) );
  XOR U5601 ( .A(n5929), .B(n5930), .Z(n5925) );
  AND U5602 ( .A(n5931), .B(n5932), .Z(n5930) );
  XNOR U5603 ( .A(p_input[3518]), .B(n5929), .Z(n5932) );
  XOR U5604 ( .A(n5929), .B(p_input[3502]), .Z(n5931) );
  XOR U5605 ( .A(n5933), .B(n5934), .Z(n5929) );
  AND U5606 ( .A(n5935), .B(n5936), .Z(n5934) );
  XNOR U5607 ( .A(p_input[3517]), .B(n5933), .Z(n5936) );
  XOR U5608 ( .A(n5933), .B(p_input[3501]), .Z(n5935) );
  XOR U5609 ( .A(n5937), .B(n5938), .Z(n5933) );
  AND U5610 ( .A(n5939), .B(n5940), .Z(n5938) );
  XNOR U5611 ( .A(p_input[3516]), .B(n5937), .Z(n5940) );
  XOR U5612 ( .A(n5937), .B(p_input[3500]), .Z(n5939) );
  XOR U5613 ( .A(n5941), .B(n5942), .Z(n5937) );
  AND U5614 ( .A(n5943), .B(n5944), .Z(n5942) );
  XNOR U5615 ( .A(p_input[3515]), .B(n5941), .Z(n5944) );
  XOR U5616 ( .A(n5941), .B(p_input[3499]), .Z(n5943) );
  XOR U5617 ( .A(n5945), .B(n5946), .Z(n5941) );
  AND U5618 ( .A(n5947), .B(n5948), .Z(n5946) );
  XNOR U5619 ( .A(p_input[3514]), .B(n5945), .Z(n5948) );
  XOR U5620 ( .A(n5945), .B(p_input[3498]), .Z(n5947) );
  XOR U5621 ( .A(n5949), .B(n5950), .Z(n5945) );
  AND U5622 ( .A(n5951), .B(n5952), .Z(n5950) );
  XNOR U5623 ( .A(p_input[3513]), .B(n5949), .Z(n5952) );
  XOR U5624 ( .A(n5949), .B(p_input[3497]), .Z(n5951) );
  XOR U5625 ( .A(n5953), .B(n5954), .Z(n5949) );
  AND U5626 ( .A(n5955), .B(n5956), .Z(n5954) );
  XNOR U5627 ( .A(p_input[3512]), .B(n5953), .Z(n5956) );
  XOR U5628 ( .A(n5953), .B(p_input[3496]), .Z(n5955) );
  XOR U5629 ( .A(n5957), .B(n5958), .Z(n5953) );
  AND U5630 ( .A(n5959), .B(n5960), .Z(n5958) );
  XNOR U5631 ( .A(p_input[3511]), .B(n5957), .Z(n5960) );
  XOR U5632 ( .A(n5957), .B(p_input[3495]), .Z(n5959) );
  XOR U5633 ( .A(n5961), .B(n5962), .Z(n5957) );
  AND U5634 ( .A(n5963), .B(n5964), .Z(n5962) );
  XNOR U5635 ( .A(p_input[3510]), .B(n5961), .Z(n5964) );
  XOR U5636 ( .A(n5961), .B(p_input[3494]), .Z(n5963) );
  XOR U5637 ( .A(n5965), .B(n5966), .Z(n5961) );
  AND U5638 ( .A(n5967), .B(n5968), .Z(n5966) );
  XNOR U5639 ( .A(p_input[3509]), .B(n5965), .Z(n5968) );
  XOR U5640 ( .A(n5965), .B(p_input[3493]), .Z(n5967) );
  XOR U5641 ( .A(n5969), .B(n5970), .Z(n5965) );
  AND U5642 ( .A(n5971), .B(n5972), .Z(n5970) );
  XNOR U5643 ( .A(p_input[3508]), .B(n5969), .Z(n5972) );
  XOR U5644 ( .A(n5969), .B(p_input[3492]), .Z(n5971) );
  XOR U5645 ( .A(n5973), .B(n5974), .Z(n5969) );
  AND U5646 ( .A(n5975), .B(n5976), .Z(n5974) );
  XNOR U5647 ( .A(p_input[3507]), .B(n5973), .Z(n5976) );
  XOR U5648 ( .A(n5973), .B(p_input[3491]), .Z(n5975) );
  XOR U5649 ( .A(n5977), .B(n5978), .Z(n5973) );
  AND U5650 ( .A(n5979), .B(n5980), .Z(n5978) );
  XNOR U5651 ( .A(p_input[3506]), .B(n5977), .Z(n5980) );
  XOR U5652 ( .A(n5977), .B(p_input[3490]), .Z(n5979) );
  XNOR U5653 ( .A(n5981), .B(n5982), .Z(n5977) );
  AND U5654 ( .A(n5983), .B(n5984), .Z(n5982) );
  XOR U5655 ( .A(p_input[3505]), .B(n5981), .Z(n5984) );
  XNOR U5656 ( .A(p_input[3489]), .B(n5981), .Z(n5983) );
  AND U5657 ( .A(p_input[3504]), .B(n5985), .Z(n5981) );
  IV U5658 ( .A(p_input[3488]), .Z(n5985) );
  XNOR U5659 ( .A(p_input[3456]), .B(n5986), .Z(n5788) );
  AND U5660 ( .A(n168), .B(n5987), .Z(n5986) );
  XOR U5661 ( .A(p_input[3472]), .B(p_input[3456]), .Z(n5987) );
  XOR U5662 ( .A(n5988), .B(n5989), .Z(n168) );
  AND U5663 ( .A(n5990), .B(n5991), .Z(n5989) );
  XNOR U5664 ( .A(p_input[3487]), .B(n5988), .Z(n5991) );
  XOR U5665 ( .A(n5988), .B(p_input[3471]), .Z(n5990) );
  XOR U5666 ( .A(n5992), .B(n5993), .Z(n5988) );
  AND U5667 ( .A(n5994), .B(n5995), .Z(n5993) );
  XNOR U5668 ( .A(p_input[3486]), .B(n5992), .Z(n5995) );
  XNOR U5669 ( .A(n5992), .B(n5802), .Z(n5994) );
  IV U5670 ( .A(p_input[3470]), .Z(n5802) );
  XOR U5671 ( .A(n5996), .B(n5997), .Z(n5992) );
  AND U5672 ( .A(n5998), .B(n5999), .Z(n5997) );
  XNOR U5673 ( .A(p_input[3485]), .B(n5996), .Z(n5999) );
  XNOR U5674 ( .A(n5996), .B(n5811), .Z(n5998) );
  IV U5675 ( .A(p_input[3469]), .Z(n5811) );
  XOR U5676 ( .A(n6000), .B(n6001), .Z(n5996) );
  AND U5677 ( .A(n6002), .B(n6003), .Z(n6001) );
  XNOR U5678 ( .A(p_input[3484]), .B(n6000), .Z(n6003) );
  XNOR U5679 ( .A(n6000), .B(n5820), .Z(n6002) );
  IV U5680 ( .A(p_input[3468]), .Z(n5820) );
  XOR U5681 ( .A(n6004), .B(n6005), .Z(n6000) );
  AND U5682 ( .A(n6006), .B(n6007), .Z(n6005) );
  XNOR U5683 ( .A(p_input[3483]), .B(n6004), .Z(n6007) );
  XNOR U5684 ( .A(n6004), .B(n5829), .Z(n6006) );
  IV U5685 ( .A(p_input[3467]), .Z(n5829) );
  XOR U5686 ( .A(n6008), .B(n6009), .Z(n6004) );
  AND U5687 ( .A(n6010), .B(n6011), .Z(n6009) );
  XNOR U5688 ( .A(p_input[3482]), .B(n6008), .Z(n6011) );
  XNOR U5689 ( .A(n6008), .B(n5838), .Z(n6010) );
  IV U5690 ( .A(p_input[3466]), .Z(n5838) );
  XOR U5691 ( .A(n6012), .B(n6013), .Z(n6008) );
  AND U5692 ( .A(n6014), .B(n6015), .Z(n6013) );
  XNOR U5693 ( .A(p_input[3481]), .B(n6012), .Z(n6015) );
  XNOR U5694 ( .A(n6012), .B(n5847), .Z(n6014) );
  IV U5695 ( .A(p_input[3465]), .Z(n5847) );
  XOR U5696 ( .A(n6016), .B(n6017), .Z(n6012) );
  AND U5697 ( .A(n6018), .B(n6019), .Z(n6017) );
  XNOR U5698 ( .A(p_input[3480]), .B(n6016), .Z(n6019) );
  XNOR U5699 ( .A(n6016), .B(n5856), .Z(n6018) );
  IV U5700 ( .A(p_input[3464]), .Z(n5856) );
  XOR U5701 ( .A(n6020), .B(n6021), .Z(n6016) );
  AND U5702 ( .A(n6022), .B(n6023), .Z(n6021) );
  XNOR U5703 ( .A(p_input[3479]), .B(n6020), .Z(n6023) );
  XNOR U5704 ( .A(n6020), .B(n5865), .Z(n6022) );
  IV U5705 ( .A(p_input[3463]), .Z(n5865) );
  XOR U5706 ( .A(n6024), .B(n6025), .Z(n6020) );
  AND U5707 ( .A(n6026), .B(n6027), .Z(n6025) );
  XNOR U5708 ( .A(p_input[3478]), .B(n6024), .Z(n6027) );
  XNOR U5709 ( .A(n6024), .B(n5874), .Z(n6026) );
  IV U5710 ( .A(p_input[3462]), .Z(n5874) );
  XOR U5711 ( .A(n6028), .B(n6029), .Z(n6024) );
  AND U5712 ( .A(n6030), .B(n6031), .Z(n6029) );
  XNOR U5713 ( .A(p_input[3477]), .B(n6028), .Z(n6031) );
  XNOR U5714 ( .A(n6028), .B(n5883), .Z(n6030) );
  IV U5715 ( .A(p_input[3461]), .Z(n5883) );
  XOR U5716 ( .A(n6032), .B(n6033), .Z(n6028) );
  AND U5717 ( .A(n6034), .B(n6035), .Z(n6033) );
  XNOR U5718 ( .A(p_input[3476]), .B(n6032), .Z(n6035) );
  XNOR U5719 ( .A(n6032), .B(n5892), .Z(n6034) );
  IV U5720 ( .A(p_input[3460]), .Z(n5892) );
  XOR U5721 ( .A(n6036), .B(n6037), .Z(n6032) );
  AND U5722 ( .A(n6038), .B(n6039), .Z(n6037) );
  XNOR U5723 ( .A(p_input[3475]), .B(n6036), .Z(n6039) );
  XNOR U5724 ( .A(n6036), .B(n5901), .Z(n6038) );
  IV U5725 ( .A(p_input[3459]), .Z(n5901) );
  XOR U5726 ( .A(n6040), .B(n6041), .Z(n6036) );
  AND U5727 ( .A(n6042), .B(n6043), .Z(n6041) );
  XNOR U5728 ( .A(p_input[3474]), .B(n6040), .Z(n6043) );
  XNOR U5729 ( .A(n6040), .B(n5910), .Z(n6042) );
  IV U5730 ( .A(p_input[3458]), .Z(n5910) );
  XNOR U5731 ( .A(n6044), .B(n6045), .Z(n6040) );
  AND U5732 ( .A(n6046), .B(n6047), .Z(n6045) );
  XOR U5733 ( .A(p_input[3473]), .B(n6044), .Z(n6047) );
  XNOR U5734 ( .A(p_input[3457]), .B(n6044), .Z(n6046) );
  AND U5735 ( .A(p_input[3472]), .B(n6048), .Z(n6044) );
  IV U5736 ( .A(p_input[3456]), .Z(n6048) );
  XOR U5737 ( .A(n6049), .B(n6050), .Z(n5164) );
  AND U5738 ( .A(n745), .B(n6051), .Z(n6050) );
  XNOR U5739 ( .A(n6052), .B(n6049), .Z(n6051) );
  XOR U5740 ( .A(n6053), .B(n6054), .Z(n745) );
  AND U5741 ( .A(n6055), .B(n6056), .Z(n6054) );
  XNOR U5742 ( .A(n5176), .B(n6053), .Z(n6056) );
  AND U5743 ( .A(n6057), .B(n6058), .Z(n5176) );
  XOR U5744 ( .A(n6053), .B(n5175), .Z(n6055) );
  AND U5745 ( .A(n6059), .B(n6060), .Z(n5175) );
  XOR U5746 ( .A(n6061), .B(n6062), .Z(n6053) );
  AND U5747 ( .A(n6063), .B(n6064), .Z(n6062) );
  XOR U5748 ( .A(n6061), .B(n5188), .Z(n6064) );
  XOR U5749 ( .A(n6065), .B(n6066), .Z(n5188) );
  AND U5750 ( .A(n391), .B(n6067), .Z(n6066) );
  XOR U5751 ( .A(n6068), .B(n6065), .Z(n6067) );
  XNOR U5752 ( .A(n5185), .B(n6061), .Z(n6063) );
  XOR U5753 ( .A(n6069), .B(n6070), .Z(n5185) );
  AND U5754 ( .A(n388), .B(n6071), .Z(n6070) );
  XOR U5755 ( .A(n6072), .B(n6069), .Z(n6071) );
  XOR U5756 ( .A(n6073), .B(n6074), .Z(n6061) );
  AND U5757 ( .A(n6075), .B(n6076), .Z(n6074) );
  XOR U5758 ( .A(n6073), .B(n5200), .Z(n6076) );
  XOR U5759 ( .A(n6077), .B(n6078), .Z(n5200) );
  AND U5760 ( .A(n391), .B(n6079), .Z(n6078) );
  XOR U5761 ( .A(n6080), .B(n6077), .Z(n6079) );
  XNOR U5762 ( .A(n5197), .B(n6073), .Z(n6075) );
  XOR U5763 ( .A(n6081), .B(n6082), .Z(n5197) );
  AND U5764 ( .A(n388), .B(n6083), .Z(n6082) );
  XOR U5765 ( .A(n6084), .B(n6081), .Z(n6083) );
  XOR U5766 ( .A(n6085), .B(n6086), .Z(n6073) );
  AND U5767 ( .A(n6087), .B(n6088), .Z(n6086) );
  XOR U5768 ( .A(n6085), .B(n5212), .Z(n6088) );
  XOR U5769 ( .A(n6089), .B(n6090), .Z(n5212) );
  AND U5770 ( .A(n391), .B(n6091), .Z(n6090) );
  XOR U5771 ( .A(n6092), .B(n6089), .Z(n6091) );
  XNOR U5772 ( .A(n5209), .B(n6085), .Z(n6087) );
  XOR U5773 ( .A(n6093), .B(n6094), .Z(n5209) );
  AND U5774 ( .A(n388), .B(n6095), .Z(n6094) );
  XOR U5775 ( .A(n6096), .B(n6093), .Z(n6095) );
  XOR U5776 ( .A(n6097), .B(n6098), .Z(n6085) );
  AND U5777 ( .A(n6099), .B(n6100), .Z(n6098) );
  XOR U5778 ( .A(n6097), .B(n5224), .Z(n6100) );
  XOR U5779 ( .A(n6101), .B(n6102), .Z(n5224) );
  AND U5780 ( .A(n391), .B(n6103), .Z(n6102) );
  XOR U5781 ( .A(n6104), .B(n6101), .Z(n6103) );
  XNOR U5782 ( .A(n5221), .B(n6097), .Z(n6099) );
  XOR U5783 ( .A(n6105), .B(n6106), .Z(n5221) );
  AND U5784 ( .A(n388), .B(n6107), .Z(n6106) );
  XOR U5785 ( .A(n6108), .B(n6105), .Z(n6107) );
  XOR U5786 ( .A(n6109), .B(n6110), .Z(n6097) );
  AND U5787 ( .A(n6111), .B(n6112), .Z(n6110) );
  XOR U5788 ( .A(n6109), .B(n5236), .Z(n6112) );
  XOR U5789 ( .A(n6113), .B(n6114), .Z(n5236) );
  AND U5790 ( .A(n391), .B(n6115), .Z(n6114) );
  XOR U5791 ( .A(n6116), .B(n6113), .Z(n6115) );
  XNOR U5792 ( .A(n5233), .B(n6109), .Z(n6111) );
  XOR U5793 ( .A(n6117), .B(n6118), .Z(n5233) );
  AND U5794 ( .A(n388), .B(n6119), .Z(n6118) );
  XOR U5795 ( .A(n6120), .B(n6117), .Z(n6119) );
  XOR U5796 ( .A(n6121), .B(n6122), .Z(n6109) );
  AND U5797 ( .A(n6123), .B(n6124), .Z(n6122) );
  XOR U5798 ( .A(n6121), .B(n5248), .Z(n6124) );
  XOR U5799 ( .A(n6125), .B(n6126), .Z(n5248) );
  AND U5800 ( .A(n391), .B(n6127), .Z(n6126) );
  XOR U5801 ( .A(n6128), .B(n6125), .Z(n6127) );
  XNOR U5802 ( .A(n5245), .B(n6121), .Z(n6123) );
  XOR U5803 ( .A(n6129), .B(n6130), .Z(n5245) );
  AND U5804 ( .A(n388), .B(n6131), .Z(n6130) );
  XOR U5805 ( .A(n6132), .B(n6129), .Z(n6131) );
  XOR U5806 ( .A(n6133), .B(n6134), .Z(n6121) );
  AND U5807 ( .A(n6135), .B(n6136), .Z(n6134) );
  XOR U5808 ( .A(n6133), .B(n5260), .Z(n6136) );
  XOR U5809 ( .A(n6137), .B(n6138), .Z(n5260) );
  AND U5810 ( .A(n391), .B(n6139), .Z(n6138) );
  XOR U5811 ( .A(n6140), .B(n6137), .Z(n6139) );
  XNOR U5812 ( .A(n5257), .B(n6133), .Z(n6135) );
  XOR U5813 ( .A(n6141), .B(n6142), .Z(n5257) );
  AND U5814 ( .A(n388), .B(n6143), .Z(n6142) );
  XOR U5815 ( .A(n6144), .B(n6141), .Z(n6143) );
  XOR U5816 ( .A(n6145), .B(n6146), .Z(n6133) );
  AND U5817 ( .A(n6147), .B(n6148), .Z(n6146) );
  XOR U5818 ( .A(n6145), .B(n5272), .Z(n6148) );
  XOR U5819 ( .A(n6149), .B(n6150), .Z(n5272) );
  AND U5820 ( .A(n391), .B(n6151), .Z(n6150) );
  XOR U5821 ( .A(n6152), .B(n6149), .Z(n6151) );
  XNOR U5822 ( .A(n5269), .B(n6145), .Z(n6147) );
  XOR U5823 ( .A(n6153), .B(n6154), .Z(n5269) );
  AND U5824 ( .A(n388), .B(n6155), .Z(n6154) );
  XOR U5825 ( .A(n6156), .B(n6153), .Z(n6155) );
  XOR U5826 ( .A(n6157), .B(n6158), .Z(n6145) );
  AND U5827 ( .A(n6159), .B(n6160), .Z(n6158) );
  XOR U5828 ( .A(n6157), .B(n5284), .Z(n6160) );
  XOR U5829 ( .A(n6161), .B(n6162), .Z(n5284) );
  AND U5830 ( .A(n391), .B(n6163), .Z(n6162) );
  XOR U5831 ( .A(n6164), .B(n6161), .Z(n6163) );
  XNOR U5832 ( .A(n5281), .B(n6157), .Z(n6159) );
  XOR U5833 ( .A(n6165), .B(n6166), .Z(n5281) );
  AND U5834 ( .A(n388), .B(n6167), .Z(n6166) );
  XOR U5835 ( .A(n6168), .B(n6165), .Z(n6167) );
  XOR U5836 ( .A(n6169), .B(n6170), .Z(n6157) );
  AND U5837 ( .A(n6171), .B(n6172), .Z(n6170) );
  XOR U5838 ( .A(n6169), .B(n5296), .Z(n6172) );
  XOR U5839 ( .A(n6173), .B(n6174), .Z(n5296) );
  AND U5840 ( .A(n391), .B(n6175), .Z(n6174) );
  XOR U5841 ( .A(n6176), .B(n6173), .Z(n6175) );
  XNOR U5842 ( .A(n5293), .B(n6169), .Z(n6171) );
  XOR U5843 ( .A(n6177), .B(n6178), .Z(n5293) );
  AND U5844 ( .A(n388), .B(n6179), .Z(n6178) );
  XOR U5845 ( .A(n6180), .B(n6177), .Z(n6179) );
  XOR U5846 ( .A(n6181), .B(n6182), .Z(n6169) );
  AND U5847 ( .A(n6183), .B(n6184), .Z(n6182) );
  XOR U5848 ( .A(n6181), .B(n5308), .Z(n6184) );
  XOR U5849 ( .A(n6185), .B(n6186), .Z(n5308) );
  AND U5850 ( .A(n391), .B(n6187), .Z(n6186) );
  XOR U5851 ( .A(n6188), .B(n6185), .Z(n6187) );
  XNOR U5852 ( .A(n5305), .B(n6181), .Z(n6183) );
  XOR U5853 ( .A(n6189), .B(n6190), .Z(n5305) );
  AND U5854 ( .A(n388), .B(n6191), .Z(n6190) );
  XOR U5855 ( .A(n6192), .B(n6189), .Z(n6191) );
  XOR U5856 ( .A(n6193), .B(n6194), .Z(n6181) );
  AND U5857 ( .A(n6195), .B(n6196), .Z(n6194) );
  XOR U5858 ( .A(n6193), .B(n5320), .Z(n6196) );
  XOR U5859 ( .A(n6197), .B(n6198), .Z(n5320) );
  AND U5860 ( .A(n391), .B(n6199), .Z(n6198) );
  XOR U5861 ( .A(n6200), .B(n6197), .Z(n6199) );
  XNOR U5862 ( .A(n5317), .B(n6193), .Z(n6195) );
  XOR U5863 ( .A(n6201), .B(n6202), .Z(n5317) );
  AND U5864 ( .A(n388), .B(n6203), .Z(n6202) );
  XOR U5865 ( .A(n6204), .B(n6201), .Z(n6203) );
  XOR U5866 ( .A(n6205), .B(n6206), .Z(n6193) );
  AND U5867 ( .A(n6207), .B(n6208), .Z(n6206) );
  XOR U5868 ( .A(n6205), .B(n5332), .Z(n6208) );
  XOR U5869 ( .A(n6209), .B(n6210), .Z(n5332) );
  AND U5870 ( .A(n391), .B(n6211), .Z(n6210) );
  XOR U5871 ( .A(n6212), .B(n6209), .Z(n6211) );
  XNOR U5872 ( .A(n5329), .B(n6205), .Z(n6207) );
  XOR U5873 ( .A(n6213), .B(n6214), .Z(n5329) );
  AND U5874 ( .A(n388), .B(n6215), .Z(n6214) );
  XOR U5875 ( .A(n6216), .B(n6213), .Z(n6215) );
  XOR U5876 ( .A(n6217), .B(n6218), .Z(n6205) );
  AND U5877 ( .A(n6219), .B(n6220), .Z(n6218) );
  XNOR U5878 ( .A(n6221), .B(n5345), .Z(n6220) );
  XOR U5879 ( .A(n6222), .B(n6223), .Z(n5345) );
  AND U5880 ( .A(n391), .B(n6224), .Z(n6223) );
  XOR U5881 ( .A(n6222), .B(n6225), .Z(n6224) );
  XNOR U5882 ( .A(n5342), .B(n6217), .Z(n6219) );
  XOR U5883 ( .A(n6226), .B(n6227), .Z(n5342) );
  AND U5884 ( .A(n388), .B(n6228), .Z(n6227) );
  XOR U5885 ( .A(n6226), .B(n6229), .Z(n6228) );
  IV U5886 ( .A(n6221), .Z(n6217) );
  AND U5887 ( .A(n6049), .B(n6052), .Z(n6221) );
  XNOR U5888 ( .A(n6230), .B(n6231), .Z(n6052) );
  AND U5889 ( .A(n391), .B(n6232), .Z(n6231) );
  XNOR U5890 ( .A(n6233), .B(n6230), .Z(n6232) );
  XOR U5891 ( .A(n6234), .B(n6235), .Z(n391) );
  AND U5892 ( .A(n6236), .B(n6237), .Z(n6235) );
  XNOR U5893 ( .A(n6057), .B(n6234), .Z(n6237) );
  AND U5894 ( .A(p_input[3455]), .B(p_input[3439]), .Z(n6057) );
  XOR U5895 ( .A(n6234), .B(n6058), .Z(n6236) );
  AND U5896 ( .A(p_input[3423]), .B(p_input[3407]), .Z(n6058) );
  XOR U5897 ( .A(n6238), .B(n6239), .Z(n6234) );
  AND U5898 ( .A(n6240), .B(n6241), .Z(n6239) );
  XOR U5899 ( .A(n6238), .B(n6068), .Z(n6241) );
  XNOR U5900 ( .A(p_input[3438]), .B(n6242), .Z(n6068) );
  AND U5901 ( .A(n179), .B(n6243), .Z(n6242) );
  XOR U5902 ( .A(p_input[3454]), .B(p_input[3438]), .Z(n6243) );
  XNOR U5903 ( .A(n6065), .B(n6238), .Z(n6240) );
  XOR U5904 ( .A(n6244), .B(n6245), .Z(n6065) );
  AND U5905 ( .A(n177), .B(n6246), .Z(n6245) );
  XOR U5906 ( .A(p_input[3422]), .B(p_input[3406]), .Z(n6246) );
  XOR U5907 ( .A(n6247), .B(n6248), .Z(n6238) );
  AND U5908 ( .A(n6249), .B(n6250), .Z(n6248) );
  XOR U5909 ( .A(n6247), .B(n6080), .Z(n6250) );
  XNOR U5910 ( .A(p_input[3437]), .B(n6251), .Z(n6080) );
  AND U5911 ( .A(n179), .B(n6252), .Z(n6251) );
  XOR U5912 ( .A(p_input[3453]), .B(p_input[3437]), .Z(n6252) );
  XNOR U5913 ( .A(n6077), .B(n6247), .Z(n6249) );
  XOR U5914 ( .A(n6253), .B(n6254), .Z(n6077) );
  AND U5915 ( .A(n177), .B(n6255), .Z(n6254) );
  XOR U5916 ( .A(p_input[3421]), .B(p_input[3405]), .Z(n6255) );
  XOR U5917 ( .A(n6256), .B(n6257), .Z(n6247) );
  AND U5918 ( .A(n6258), .B(n6259), .Z(n6257) );
  XOR U5919 ( .A(n6256), .B(n6092), .Z(n6259) );
  XNOR U5920 ( .A(p_input[3436]), .B(n6260), .Z(n6092) );
  AND U5921 ( .A(n179), .B(n6261), .Z(n6260) );
  XOR U5922 ( .A(p_input[3452]), .B(p_input[3436]), .Z(n6261) );
  XNOR U5923 ( .A(n6089), .B(n6256), .Z(n6258) );
  XOR U5924 ( .A(n6262), .B(n6263), .Z(n6089) );
  AND U5925 ( .A(n177), .B(n6264), .Z(n6263) );
  XOR U5926 ( .A(p_input[3420]), .B(p_input[3404]), .Z(n6264) );
  XOR U5927 ( .A(n6265), .B(n6266), .Z(n6256) );
  AND U5928 ( .A(n6267), .B(n6268), .Z(n6266) );
  XOR U5929 ( .A(n6265), .B(n6104), .Z(n6268) );
  XNOR U5930 ( .A(p_input[3435]), .B(n6269), .Z(n6104) );
  AND U5931 ( .A(n179), .B(n6270), .Z(n6269) );
  XOR U5932 ( .A(p_input[3451]), .B(p_input[3435]), .Z(n6270) );
  XNOR U5933 ( .A(n6101), .B(n6265), .Z(n6267) );
  XOR U5934 ( .A(n6271), .B(n6272), .Z(n6101) );
  AND U5935 ( .A(n177), .B(n6273), .Z(n6272) );
  XOR U5936 ( .A(p_input[3419]), .B(p_input[3403]), .Z(n6273) );
  XOR U5937 ( .A(n6274), .B(n6275), .Z(n6265) );
  AND U5938 ( .A(n6276), .B(n6277), .Z(n6275) );
  XOR U5939 ( .A(n6274), .B(n6116), .Z(n6277) );
  XNOR U5940 ( .A(p_input[3434]), .B(n6278), .Z(n6116) );
  AND U5941 ( .A(n179), .B(n6279), .Z(n6278) );
  XOR U5942 ( .A(p_input[3450]), .B(p_input[3434]), .Z(n6279) );
  XNOR U5943 ( .A(n6113), .B(n6274), .Z(n6276) );
  XOR U5944 ( .A(n6280), .B(n6281), .Z(n6113) );
  AND U5945 ( .A(n177), .B(n6282), .Z(n6281) );
  XOR U5946 ( .A(p_input[3418]), .B(p_input[3402]), .Z(n6282) );
  XOR U5947 ( .A(n6283), .B(n6284), .Z(n6274) );
  AND U5948 ( .A(n6285), .B(n6286), .Z(n6284) );
  XOR U5949 ( .A(n6283), .B(n6128), .Z(n6286) );
  XNOR U5950 ( .A(p_input[3433]), .B(n6287), .Z(n6128) );
  AND U5951 ( .A(n179), .B(n6288), .Z(n6287) );
  XOR U5952 ( .A(p_input[3449]), .B(p_input[3433]), .Z(n6288) );
  XNOR U5953 ( .A(n6125), .B(n6283), .Z(n6285) );
  XOR U5954 ( .A(n6289), .B(n6290), .Z(n6125) );
  AND U5955 ( .A(n177), .B(n6291), .Z(n6290) );
  XOR U5956 ( .A(p_input[3417]), .B(p_input[3401]), .Z(n6291) );
  XOR U5957 ( .A(n6292), .B(n6293), .Z(n6283) );
  AND U5958 ( .A(n6294), .B(n6295), .Z(n6293) );
  XOR U5959 ( .A(n6292), .B(n6140), .Z(n6295) );
  XNOR U5960 ( .A(p_input[3432]), .B(n6296), .Z(n6140) );
  AND U5961 ( .A(n179), .B(n6297), .Z(n6296) );
  XOR U5962 ( .A(p_input[3448]), .B(p_input[3432]), .Z(n6297) );
  XNOR U5963 ( .A(n6137), .B(n6292), .Z(n6294) );
  XOR U5964 ( .A(n6298), .B(n6299), .Z(n6137) );
  AND U5965 ( .A(n177), .B(n6300), .Z(n6299) );
  XOR U5966 ( .A(p_input[3416]), .B(p_input[3400]), .Z(n6300) );
  XOR U5967 ( .A(n6301), .B(n6302), .Z(n6292) );
  AND U5968 ( .A(n6303), .B(n6304), .Z(n6302) );
  XOR U5969 ( .A(n6301), .B(n6152), .Z(n6304) );
  XNOR U5970 ( .A(p_input[3431]), .B(n6305), .Z(n6152) );
  AND U5971 ( .A(n179), .B(n6306), .Z(n6305) );
  XOR U5972 ( .A(p_input[3447]), .B(p_input[3431]), .Z(n6306) );
  XNOR U5973 ( .A(n6149), .B(n6301), .Z(n6303) );
  XOR U5974 ( .A(n6307), .B(n6308), .Z(n6149) );
  AND U5975 ( .A(n177), .B(n6309), .Z(n6308) );
  XOR U5976 ( .A(p_input[3415]), .B(p_input[3399]), .Z(n6309) );
  XOR U5977 ( .A(n6310), .B(n6311), .Z(n6301) );
  AND U5978 ( .A(n6312), .B(n6313), .Z(n6311) );
  XOR U5979 ( .A(n6310), .B(n6164), .Z(n6313) );
  XNOR U5980 ( .A(p_input[3430]), .B(n6314), .Z(n6164) );
  AND U5981 ( .A(n179), .B(n6315), .Z(n6314) );
  XOR U5982 ( .A(p_input[3446]), .B(p_input[3430]), .Z(n6315) );
  XNOR U5983 ( .A(n6161), .B(n6310), .Z(n6312) );
  XOR U5984 ( .A(n6316), .B(n6317), .Z(n6161) );
  AND U5985 ( .A(n177), .B(n6318), .Z(n6317) );
  XOR U5986 ( .A(p_input[3414]), .B(p_input[3398]), .Z(n6318) );
  XOR U5987 ( .A(n6319), .B(n6320), .Z(n6310) );
  AND U5988 ( .A(n6321), .B(n6322), .Z(n6320) );
  XOR U5989 ( .A(n6319), .B(n6176), .Z(n6322) );
  XNOR U5990 ( .A(p_input[3429]), .B(n6323), .Z(n6176) );
  AND U5991 ( .A(n179), .B(n6324), .Z(n6323) );
  XOR U5992 ( .A(p_input[3445]), .B(p_input[3429]), .Z(n6324) );
  XNOR U5993 ( .A(n6173), .B(n6319), .Z(n6321) );
  XOR U5994 ( .A(n6325), .B(n6326), .Z(n6173) );
  AND U5995 ( .A(n177), .B(n6327), .Z(n6326) );
  XOR U5996 ( .A(p_input[3413]), .B(p_input[3397]), .Z(n6327) );
  XOR U5997 ( .A(n6328), .B(n6329), .Z(n6319) );
  AND U5998 ( .A(n6330), .B(n6331), .Z(n6329) );
  XOR U5999 ( .A(n6328), .B(n6188), .Z(n6331) );
  XNOR U6000 ( .A(p_input[3428]), .B(n6332), .Z(n6188) );
  AND U6001 ( .A(n179), .B(n6333), .Z(n6332) );
  XOR U6002 ( .A(p_input[3444]), .B(p_input[3428]), .Z(n6333) );
  XNOR U6003 ( .A(n6185), .B(n6328), .Z(n6330) );
  XOR U6004 ( .A(n6334), .B(n6335), .Z(n6185) );
  AND U6005 ( .A(n177), .B(n6336), .Z(n6335) );
  XOR U6006 ( .A(p_input[3412]), .B(p_input[3396]), .Z(n6336) );
  XOR U6007 ( .A(n6337), .B(n6338), .Z(n6328) );
  AND U6008 ( .A(n6339), .B(n6340), .Z(n6338) );
  XOR U6009 ( .A(n6337), .B(n6200), .Z(n6340) );
  XNOR U6010 ( .A(p_input[3427]), .B(n6341), .Z(n6200) );
  AND U6011 ( .A(n179), .B(n6342), .Z(n6341) );
  XOR U6012 ( .A(p_input[3443]), .B(p_input[3427]), .Z(n6342) );
  XNOR U6013 ( .A(n6197), .B(n6337), .Z(n6339) );
  XOR U6014 ( .A(n6343), .B(n6344), .Z(n6197) );
  AND U6015 ( .A(n177), .B(n6345), .Z(n6344) );
  XOR U6016 ( .A(p_input[3411]), .B(p_input[3395]), .Z(n6345) );
  XOR U6017 ( .A(n6346), .B(n6347), .Z(n6337) );
  AND U6018 ( .A(n6348), .B(n6349), .Z(n6347) );
  XOR U6019 ( .A(n6346), .B(n6212), .Z(n6349) );
  XNOR U6020 ( .A(p_input[3426]), .B(n6350), .Z(n6212) );
  AND U6021 ( .A(n179), .B(n6351), .Z(n6350) );
  XOR U6022 ( .A(p_input[3442]), .B(p_input[3426]), .Z(n6351) );
  XNOR U6023 ( .A(n6209), .B(n6346), .Z(n6348) );
  XOR U6024 ( .A(n6352), .B(n6353), .Z(n6209) );
  AND U6025 ( .A(n177), .B(n6354), .Z(n6353) );
  XOR U6026 ( .A(p_input[3410]), .B(p_input[3394]), .Z(n6354) );
  XOR U6027 ( .A(n6355), .B(n6356), .Z(n6346) );
  AND U6028 ( .A(n6357), .B(n6358), .Z(n6356) );
  XNOR U6029 ( .A(n6359), .B(n6225), .Z(n6358) );
  XNOR U6030 ( .A(p_input[3425]), .B(n6360), .Z(n6225) );
  AND U6031 ( .A(n179), .B(n6361), .Z(n6360) );
  XNOR U6032 ( .A(p_input[3441]), .B(n6362), .Z(n6361) );
  IV U6033 ( .A(p_input[3425]), .Z(n6362) );
  XNOR U6034 ( .A(n6222), .B(n6355), .Z(n6357) );
  XNOR U6035 ( .A(p_input[3393]), .B(n6363), .Z(n6222) );
  AND U6036 ( .A(n177), .B(n6364), .Z(n6363) );
  XOR U6037 ( .A(p_input[3409]), .B(p_input[3393]), .Z(n6364) );
  IV U6038 ( .A(n6359), .Z(n6355) );
  AND U6039 ( .A(n6230), .B(n6233), .Z(n6359) );
  XOR U6040 ( .A(p_input[3424]), .B(n6365), .Z(n6233) );
  AND U6041 ( .A(n179), .B(n6366), .Z(n6365) );
  XOR U6042 ( .A(p_input[3440]), .B(p_input[3424]), .Z(n6366) );
  XOR U6043 ( .A(n6367), .B(n6368), .Z(n179) );
  AND U6044 ( .A(n6369), .B(n6370), .Z(n6368) );
  XNOR U6045 ( .A(p_input[3455]), .B(n6367), .Z(n6370) );
  XOR U6046 ( .A(n6367), .B(p_input[3439]), .Z(n6369) );
  XOR U6047 ( .A(n6371), .B(n6372), .Z(n6367) );
  AND U6048 ( .A(n6373), .B(n6374), .Z(n6372) );
  XNOR U6049 ( .A(p_input[3454]), .B(n6371), .Z(n6374) );
  XOR U6050 ( .A(n6371), .B(p_input[3438]), .Z(n6373) );
  XOR U6051 ( .A(n6375), .B(n6376), .Z(n6371) );
  AND U6052 ( .A(n6377), .B(n6378), .Z(n6376) );
  XNOR U6053 ( .A(p_input[3453]), .B(n6375), .Z(n6378) );
  XOR U6054 ( .A(n6375), .B(p_input[3437]), .Z(n6377) );
  XOR U6055 ( .A(n6379), .B(n6380), .Z(n6375) );
  AND U6056 ( .A(n6381), .B(n6382), .Z(n6380) );
  XNOR U6057 ( .A(p_input[3452]), .B(n6379), .Z(n6382) );
  XOR U6058 ( .A(n6379), .B(p_input[3436]), .Z(n6381) );
  XOR U6059 ( .A(n6383), .B(n6384), .Z(n6379) );
  AND U6060 ( .A(n6385), .B(n6386), .Z(n6384) );
  XNOR U6061 ( .A(p_input[3451]), .B(n6383), .Z(n6386) );
  XOR U6062 ( .A(n6383), .B(p_input[3435]), .Z(n6385) );
  XOR U6063 ( .A(n6387), .B(n6388), .Z(n6383) );
  AND U6064 ( .A(n6389), .B(n6390), .Z(n6388) );
  XNOR U6065 ( .A(p_input[3450]), .B(n6387), .Z(n6390) );
  XOR U6066 ( .A(n6387), .B(p_input[3434]), .Z(n6389) );
  XOR U6067 ( .A(n6391), .B(n6392), .Z(n6387) );
  AND U6068 ( .A(n6393), .B(n6394), .Z(n6392) );
  XNOR U6069 ( .A(p_input[3449]), .B(n6391), .Z(n6394) );
  XOR U6070 ( .A(n6391), .B(p_input[3433]), .Z(n6393) );
  XOR U6071 ( .A(n6395), .B(n6396), .Z(n6391) );
  AND U6072 ( .A(n6397), .B(n6398), .Z(n6396) );
  XNOR U6073 ( .A(p_input[3448]), .B(n6395), .Z(n6398) );
  XOR U6074 ( .A(n6395), .B(p_input[3432]), .Z(n6397) );
  XOR U6075 ( .A(n6399), .B(n6400), .Z(n6395) );
  AND U6076 ( .A(n6401), .B(n6402), .Z(n6400) );
  XNOR U6077 ( .A(p_input[3447]), .B(n6399), .Z(n6402) );
  XOR U6078 ( .A(n6399), .B(p_input[3431]), .Z(n6401) );
  XOR U6079 ( .A(n6403), .B(n6404), .Z(n6399) );
  AND U6080 ( .A(n6405), .B(n6406), .Z(n6404) );
  XNOR U6081 ( .A(p_input[3446]), .B(n6403), .Z(n6406) );
  XOR U6082 ( .A(n6403), .B(p_input[3430]), .Z(n6405) );
  XOR U6083 ( .A(n6407), .B(n6408), .Z(n6403) );
  AND U6084 ( .A(n6409), .B(n6410), .Z(n6408) );
  XNOR U6085 ( .A(p_input[3445]), .B(n6407), .Z(n6410) );
  XOR U6086 ( .A(n6407), .B(p_input[3429]), .Z(n6409) );
  XOR U6087 ( .A(n6411), .B(n6412), .Z(n6407) );
  AND U6088 ( .A(n6413), .B(n6414), .Z(n6412) );
  XNOR U6089 ( .A(p_input[3444]), .B(n6411), .Z(n6414) );
  XOR U6090 ( .A(n6411), .B(p_input[3428]), .Z(n6413) );
  XOR U6091 ( .A(n6415), .B(n6416), .Z(n6411) );
  AND U6092 ( .A(n6417), .B(n6418), .Z(n6416) );
  XNOR U6093 ( .A(p_input[3443]), .B(n6415), .Z(n6418) );
  XOR U6094 ( .A(n6415), .B(p_input[3427]), .Z(n6417) );
  XOR U6095 ( .A(n6419), .B(n6420), .Z(n6415) );
  AND U6096 ( .A(n6421), .B(n6422), .Z(n6420) );
  XNOR U6097 ( .A(p_input[3442]), .B(n6419), .Z(n6422) );
  XOR U6098 ( .A(n6419), .B(p_input[3426]), .Z(n6421) );
  XNOR U6099 ( .A(n6423), .B(n6424), .Z(n6419) );
  AND U6100 ( .A(n6425), .B(n6426), .Z(n6424) );
  XOR U6101 ( .A(p_input[3441]), .B(n6423), .Z(n6426) );
  XNOR U6102 ( .A(p_input[3425]), .B(n6423), .Z(n6425) );
  AND U6103 ( .A(p_input[3440]), .B(n6427), .Z(n6423) );
  IV U6104 ( .A(p_input[3424]), .Z(n6427) );
  XNOR U6105 ( .A(p_input[3392]), .B(n6428), .Z(n6230) );
  AND U6106 ( .A(n177), .B(n6429), .Z(n6428) );
  XOR U6107 ( .A(p_input[3408]), .B(p_input[3392]), .Z(n6429) );
  XOR U6108 ( .A(n6430), .B(n6431), .Z(n177) );
  AND U6109 ( .A(n6432), .B(n6433), .Z(n6431) );
  XNOR U6110 ( .A(p_input[3423]), .B(n6430), .Z(n6433) );
  XOR U6111 ( .A(n6430), .B(p_input[3407]), .Z(n6432) );
  XOR U6112 ( .A(n6434), .B(n6435), .Z(n6430) );
  AND U6113 ( .A(n6436), .B(n6437), .Z(n6435) );
  XNOR U6114 ( .A(p_input[3422]), .B(n6434), .Z(n6437) );
  XNOR U6115 ( .A(n6434), .B(n6244), .Z(n6436) );
  IV U6116 ( .A(p_input[3406]), .Z(n6244) );
  XOR U6117 ( .A(n6438), .B(n6439), .Z(n6434) );
  AND U6118 ( .A(n6440), .B(n6441), .Z(n6439) );
  XNOR U6119 ( .A(p_input[3421]), .B(n6438), .Z(n6441) );
  XNOR U6120 ( .A(n6438), .B(n6253), .Z(n6440) );
  IV U6121 ( .A(p_input[3405]), .Z(n6253) );
  XOR U6122 ( .A(n6442), .B(n6443), .Z(n6438) );
  AND U6123 ( .A(n6444), .B(n6445), .Z(n6443) );
  XNOR U6124 ( .A(p_input[3420]), .B(n6442), .Z(n6445) );
  XNOR U6125 ( .A(n6442), .B(n6262), .Z(n6444) );
  IV U6126 ( .A(p_input[3404]), .Z(n6262) );
  XOR U6127 ( .A(n6446), .B(n6447), .Z(n6442) );
  AND U6128 ( .A(n6448), .B(n6449), .Z(n6447) );
  XNOR U6129 ( .A(p_input[3419]), .B(n6446), .Z(n6449) );
  XNOR U6130 ( .A(n6446), .B(n6271), .Z(n6448) );
  IV U6131 ( .A(p_input[3403]), .Z(n6271) );
  XOR U6132 ( .A(n6450), .B(n6451), .Z(n6446) );
  AND U6133 ( .A(n6452), .B(n6453), .Z(n6451) );
  XNOR U6134 ( .A(p_input[3418]), .B(n6450), .Z(n6453) );
  XNOR U6135 ( .A(n6450), .B(n6280), .Z(n6452) );
  IV U6136 ( .A(p_input[3402]), .Z(n6280) );
  XOR U6137 ( .A(n6454), .B(n6455), .Z(n6450) );
  AND U6138 ( .A(n6456), .B(n6457), .Z(n6455) );
  XNOR U6139 ( .A(p_input[3417]), .B(n6454), .Z(n6457) );
  XNOR U6140 ( .A(n6454), .B(n6289), .Z(n6456) );
  IV U6141 ( .A(p_input[3401]), .Z(n6289) );
  XOR U6142 ( .A(n6458), .B(n6459), .Z(n6454) );
  AND U6143 ( .A(n6460), .B(n6461), .Z(n6459) );
  XNOR U6144 ( .A(p_input[3416]), .B(n6458), .Z(n6461) );
  XNOR U6145 ( .A(n6458), .B(n6298), .Z(n6460) );
  IV U6146 ( .A(p_input[3400]), .Z(n6298) );
  XOR U6147 ( .A(n6462), .B(n6463), .Z(n6458) );
  AND U6148 ( .A(n6464), .B(n6465), .Z(n6463) );
  XNOR U6149 ( .A(p_input[3415]), .B(n6462), .Z(n6465) );
  XNOR U6150 ( .A(n6462), .B(n6307), .Z(n6464) );
  IV U6151 ( .A(p_input[3399]), .Z(n6307) );
  XOR U6152 ( .A(n6466), .B(n6467), .Z(n6462) );
  AND U6153 ( .A(n6468), .B(n6469), .Z(n6467) );
  XNOR U6154 ( .A(p_input[3414]), .B(n6466), .Z(n6469) );
  XNOR U6155 ( .A(n6466), .B(n6316), .Z(n6468) );
  IV U6156 ( .A(p_input[3398]), .Z(n6316) );
  XOR U6157 ( .A(n6470), .B(n6471), .Z(n6466) );
  AND U6158 ( .A(n6472), .B(n6473), .Z(n6471) );
  XNOR U6159 ( .A(p_input[3413]), .B(n6470), .Z(n6473) );
  XNOR U6160 ( .A(n6470), .B(n6325), .Z(n6472) );
  IV U6161 ( .A(p_input[3397]), .Z(n6325) );
  XOR U6162 ( .A(n6474), .B(n6475), .Z(n6470) );
  AND U6163 ( .A(n6476), .B(n6477), .Z(n6475) );
  XNOR U6164 ( .A(p_input[3412]), .B(n6474), .Z(n6477) );
  XNOR U6165 ( .A(n6474), .B(n6334), .Z(n6476) );
  IV U6166 ( .A(p_input[3396]), .Z(n6334) );
  XOR U6167 ( .A(n6478), .B(n6479), .Z(n6474) );
  AND U6168 ( .A(n6480), .B(n6481), .Z(n6479) );
  XNOR U6169 ( .A(p_input[3411]), .B(n6478), .Z(n6481) );
  XNOR U6170 ( .A(n6478), .B(n6343), .Z(n6480) );
  IV U6171 ( .A(p_input[3395]), .Z(n6343) );
  XOR U6172 ( .A(n6482), .B(n6483), .Z(n6478) );
  AND U6173 ( .A(n6484), .B(n6485), .Z(n6483) );
  XNOR U6174 ( .A(p_input[3410]), .B(n6482), .Z(n6485) );
  XNOR U6175 ( .A(n6482), .B(n6352), .Z(n6484) );
  IV U6176 ( .A(p_input[3394]), .Z(n6352) );
  XNOR U6177 ( .A(n6486), .B(n6487), .Z(n6482) );
  AND U6178 ( .A(n6488), .B(n6489), .Z(n6487) );
  XOR U6179 ( .A(p_input[3409]), .B(n6486), .Z(n6489) );
  XNOR U6180 ( .A(p_input[3393]), .B(n6486), .Z(n6488) );
  AND U6181 ( .A(p_input[3408]), .B(n6490), .Z(n6486) );
  IV U6182 ( .A(p_input[3392]), .Z(n6490) );
  XOR U6183 ( .A(n6491), .B(n6492), .Z(n6049) );
  AND U6184 ( .A(n388), .B(n6493), .Z(n6492) );
  XNOR U6185 ( .A(n6494), .B(n6491), .Z(n6493) );
  XOR U6186 ( .A(n6495), .B(n6496), .Z(n388) );
  AND U6187 ( .A(n6497), .B(n6498), .Z(n6496) );
  XNOR U6188 ( .A(n6060), .B(n6495), .Z(n6498) );
  AND U6189 ( .A(p_input[3391]), .B(p_input[3375]), .Z(n6060) );
  XOR U6190 ( .A(n6495), .B(n6059), .Z(n6497) );
  AND U6191 ( .A(p_input[3343]), .B(p_input[3359]), .Z(n6059) );
  XOR U6192 ( .A(n6499), .B(n6500), .Z(n6495) );
  AND U6193 ( .A(n6501), .B(n6502), .Z(n6500) );
  XOR U6194 ( .A(n6499), .B(n6072), .Z(n6502) );
  XNOR U6195 ( .A(p_input[3374]), .B(n6503), .Z(n6072) );
  AND U6196 ( .A(n183), .B(n6504), .Z(n6503) );
  XOR U6197 ( .A(p_input[3390]), .B(p_input[3374]), .Z(n6504) );
  XNOR U6198 ( .A(n6069), .B(n6499), .Z(n6501) );
  XOR U6199 ( .A(n6505), .B(n6506), .Z(n6069) );
  AND U6200 ( .A(n180), .B(n6507), .Z(n6506) );
  XOR U6201 ( .A(p_input[3358]), .B(p_input[3342]), .Z(n6507) );
  XOR U6202 ( .A(n6508), .B(n6509), .Z(n6499) );
  AND U6203 ( .A(n6510), .B(n6511), .Z(n6509) );
  XOR U6204 ( .A(n6508), .B(n6084), .Z(n6511) );
  XNOR U6205 ( .A(p_input[3373]), .B(n6512), .Z(n6084) );
  AND U6206 ( .A(n183), .B(n6513), .Z(n6512) );
  XOR U6207 ( .A(p_input[3389]), .B(p_input[3373]), .Z(n6513) );
  XNOR U6208 ( .A(n6081), .B(n6508), .Z(n6510) );
  XOR U6209 ( .A(n6514), .B(n6515), .Z(n6081) );
  AND U6210 ( .A(n180), .B(n6516), .Z(n6515) );
  XOR U6211 ( .A(p_input[3357]), .B(p_input[3341]), .Z(n6516) );
  XOR U6212 ( .A(n6517), .B(n6518), .Z(n6508) );
  AND U6213 ( .A(n6519), .B(n6520), .Z(n6518) );
  XOR U6214 ( .A(n6517), .B(n6096), .Z(n6520) );
  XNOR U6215 ( .A(p_input[3372]), .B(n6521), .Z(n6096) );
  AND U6216 ( .A(n183), .B(n6522), .Z(n6521) );
  XOR U6217 ( .A(p_input[3388]), .B(p_input[3372]), .Z(n6522) );
  XNOR U6218 ( .A(n6093), .B(n6517), .Z(n6519) );
  XOR U6219 ( .A(n6523), .B(n6524), .Z(n6093) );
  AND U6220 ( .A(n180), .B(n6525), .Z(n6524) );
  XOR U6221 ( .A(p_input[3356]), .B(p_input[3340]), .Z(n6525) );
  XOR U6222 ( .A(n6526), .B(n6527), .Z(n6517) );
  AND U6223 ( .A(n6528), .B(n6529), .Z(n6527) );
  XOR U6224 ( .A(n6526), .B(n6108), .Z(n6529) );
  XNOR U6225 ( .A(p_input[3371]), .B(n6530), .Z(n6108) );
  AND U6226 ( .A(n183), .B(n6531), .Z(n6530) );
  XOR U6227 ( .A(p_input[3387]), .B(p_input[3371]), .Z(n6531) );
  XNOR U6228 ( .A(n6105), .B(n6526), .Z(n6528) );
  XOR U6229 ( .A(n6532), .B(n6533), .Z(n6105) );
  AND U6230 ( .A(n180), .B(n6534), .Z(n6533) );
  XOR U6231 ( .A(p_input[3355]), .B(p_input[3339]), .Z(n6534) );
  XOR U6232 ( .A(n6535), .B(n6536), .Z(n6526) );
  AND U6233 ( .A(n6537), .B(n6538), .Z(n6536) );
  XOR U6234 ( .A(n6535), .B(n6120), .Z(n6538) );
  XNOR U6235 ( .A(p_input[3370]), .B(n6539), .Z(n6120) );
  AND U6236 ( .A(n183), .B(n6540), .Z(n6539) );
  XOR U6237 ( .A(p_input[3386]), .B(p_input[3370]), .Z(n6540) );
  XNOR U6238 ( .A(n6117), .B(n6535), .Z(n6537) );
  XOR U6239 ( .A(n6541), .B(n6542), .Z(n6117) );
  AND U6240 ( .A(n180), .B(n6543), .Z(n6542) );
  XOR U6241 ( .A(p_input[3354]), .B(p_input[3338]), .Z(n6543) );
  XOR U6242 ( .A(n6544), .B(n6545), .Z(n6535) );
  AND U6243 ( .A(n6546), .B(n6547), .Z(n6545) );
  XOR U6244 ( .A(n6544), .B(n6132), .Z(n6547) );
  XNOR U6245 ( .A(p_input[3369]), .B(n6548), .Z(n6132) );
  AND U6246 ( .A(n183), .B(n6549), .Z(n6548) );
  XOR U6247 ( .A(p_input[3385]), .B(p_input[3369]), .Z(n6549) );
  XNOR U6248 ( .A(n6129), .B(n6544), .Z(n6546) );
  XOR U6249 ( .A(n6550), .B(n6551), .Z(n6129) );
  AND U6250 ( .A(n180), .B(n6552), .Z(n6551) );
  XOR U6251 ( .A(p_input[3353]), .B(p_input[3337]), .Z(n6552) );
  XOR U6252 ( .A(n6553), .B(n6554), .Z(n6544) );
  AND U6253 ( .A(n6555), .B(n6556), .Z(n6554) );
  XOR U6254 ( .A(n6553), .B(n6144), .Z(n6556) );
  XNOR U6255 ( .A(p_input[3368]), .B(n6557), .Z(n6144) );
  AND U6256 ( .A(n183), .B(n6558), .Z(n6557) );
  XOR U6257 ( .A(p_input[3384]), .B(p_input[3368]), .Z(n6558) );
  XNOR U6258 ( .A(n6141), .B(n6553), .Z(n6555) );
  XOR U6259 ( .A(n6559), .B(n6560), .Z(n6141) );
  AND U6260 ( .A(n180), .B(n6561), .Z(n6560) );
  XOR U6261 ( .A(p_input[3352]), .B(p_input[3336]), .Z(n6561) );
  XOR U6262 ( .A(n6562), .B(n6563), .Z(n6553) );
  AND U6263 ( .A(n6564), .B(n6565), .Z(n6563) );
  XOR U6264 ( .A(n6562), .B(n6156), .Z(n6565) );
  XNOR U6265 ( .A(p_input[3367]), .B(n6566), .Z(n6156) );
  AND U6266 ( .A(n183), .B(n6567), .Z(n6566) );
  XOR U6267 ( .A(p_input[3383]), .B(p_input[3367]), .Z(n6567) );
  XNOR U6268 ( .A(n6153), .B(n6562), .Z(n6564) );
  XOR U6269 ( .A(n6568), .B(n6569), .Z(n6153) );
  AND U6270 ( .A(n180), .B(n6570), .Z(n6569) );
  XOR U6271 ( .A(p_input[3351]), .B(p_input[3335]), .Z(n6570) );
  XOR U6272 ( .A(n6571), .B(n6572), .Z(n6562) );
  AND U6273 ( .A(n6573), .B(n6574), .Z(n6572) );
  XOR U6274 ( .A(n6571), .B(n6168), .Z(n6574) );
  XNOR U6275 ( .A(p_input[3366]), .B(n6575), .Z(n6168) );
  AND U6276 ( .A(n183), .B(n6576), .Z(n6575) );
  XOR U6277 ( .A(p_input[3382]), .B(p_input[3366]), .Z(n6576) );
  XNOR U6278 ( .A(n6165), .B(n6571), .Z(n6573) );
  XOR U6279 ( .A(n6577), .B(n6578), .Z(n6165) );
  AND U6280 ( .A(n180), .B(n6579), .Z(n6578) );
  XOR U6281 ( .A(p_input[3350]), .B(p_input[3334]), .Z(n6579) );
  XOR U6282 ( .A(n6580), .B(n6581), .Z(n6571) );
  AND U6283 ( .A(n6582), .B(n6583), .Z(n6581) );
  XOR U6284 ( .A(n6580), .B(n6180), .Z(n6583) );
  XNOR U6285 ( .A(p_input[3365]), .B(n6584), .Z(n6180) );
  AND U6286 ( .A(n183), .B(n6585), .Z(n6584) );
  XOR U6287 ( .A(p_input[3381]), .B(p_input[3365]), .Z(n6585) );
  XNOR U6288 ( .A(n6177), .B(n6580), .Z(n6582) );
  XOR U6289 ( .A(n6586), .B(n6587), .Z(n6177) );
  AND U6290 ( .A(n180), .B(n6588), .Z(n6587) );
  XOR U6291 ( .A(p_input[3349]), .B(p_input[3333]), .Z(n6588) );
  XOR U6292 ( .A(n6589), .B(n6590), .Z(n6580) );
  AND U6293 ( .A(n6591), .B(n6592), .Z(n6590) );
  XOR U6294 ( .A(n6589), .B(n6192), .Z(n6592) );
  XNOR U6295 ( .A(p_input[3364]), .B(n6593), .Z(n6192) );
  AND U6296 ( .A(n183), .B(n6594), .Z(n6593) );
  XOR U6297 ( .A(p_input[3380]), .B(p_input[3364]), .Z(n6594) );
  XNOR U6298 ( .A(n6189), .B(n6589), .Z(n6591) );
  XOR U6299 ( .A(n6595), .B(n6596), .Z(n6189) );
  AND U6300 ( .A(n180), .B(n6597), .Z(n6596) );
  XOR U6301 ( .A(p_input[3348]), .B(p_input[3332]), .Z(n6597) );
  XOR U6302 ( .A(n6598), .B(n6599), .Z(n6589) );
  AND U6303 ( .A(n6600), .B(n6601), .Z(n6599) );
  XOR U6304 ( .A(n6598), .B(n6204), .Z(n6601) );
  XNOR U6305 ( .A(p_input[3363]), .B(n6602), .Z(n6204) );
  AND U6306 ( .A(n183), .B(n6603), .Z(n6602) );
  XOR U6307 ( .A(p_input[3379]), .B(p_input[3363]), .Z(n6603) );
  XNOR U6308 ( .A(n6201), .B(n6598), .Z(n6600) );
  XOR U6309 ( .A(n6604), .B(n6605), .Z(n6201) );
  AND U6310 ( .A(n180), .B(n6606), .Z(n6605) );
  XOR U6311 ( .A(p_input[3347]), .B(p_input[3331]), .Z(n6606) );
  XOR U6312 ( .A(n6607), .B(n6608), .Z(n6598) );
  AND U6313 ( .A(n6609), .B(n6610), .Z(n6608) );
  XOR U6314 ( .A(n6607), .B(n6216), .Z(n6610) );
  XNOR U6315 ( .A(p_input[3362]), .B(n6611), .Z(n6216) );
  AND U6316 ( .A(n183), .B(n6612), .Z(n6611) );
  XOR U6317 ( .A(p_input[3378]), .B(p_input[3362]), .Z(n6612) );
  XNOR U6318 ( .A(n6213), .B(n6607), .Z(n6609) );
  XOR U6319 ( .A(n6613), .B(n6614), .Z(n6213) );
  AND U6320 ( .A(n180), .B(n6615), .Z(n6614) );
  XOR U6321 ( .A(p_input[3346]), .B(p_input[3330]), .Z(n6615) );
  XOR U6322 ( .A(n6616), .B(n6617), .Z(n6607) );
  AND U6323 ( .A(n6618), .B(n6619), .Z(n6617) );
  XNOR U6324 ( .A(n6620), .B(n6229), .Z(n6619) );
  XNOR U6325 ( .A(p_input[3361]), .B(n6621), .Z(n6229) );
  AND U6326 ( .A(n183), .B(n6622), .Z(n6621) );
  XNOR U6327 ( .A(p_input[3377]), .B(n6623), .Z(n6622) );
  IV U6328 ( .A(p_input[3361]), .Z(n6623) );
  XNOR U6329 ( .A(n6226), .B(n6616), .Z(n6618) );
  XNOR U6330 ( .A(p_input[3329]), .B(n6624), .Z(n6226) );
  AND U6331 ( .A(n180), .B(n6625), .Z(n6624) );
  XOR U6332 ( .A(p_input[3345]), .B(p_input[3329]), .Z(n6625) );
  IV U6333 ( .A(n6620), .Z(n6616) );
  AND U6334 ( .A(n6491), .B(n6494), .Z(n6620) );
  XOR U6335 ( .A(p_input[3360]), .B(n6626), .Z(n6494) );
  AND U6336 ( .A(n183), .B(n6627), .Z(n6626) );
  XOR U6337 ( .A(p_input[3376]), .B(p_input[3360]), .Z(n6627) );
  XOR U6338 ( .A(n6628), .B(n6629), .Z(n183) );
  AND U6339 ( .A(n6630), .B(n6631), .Z(n6629) );
  XNOR U6340 ( .A(p_input[3391]), .B(n6628), .Z(n6631) );
  XOR U6341 ( .A(n6628), .B(p_input[3375]), .Z(n6630) );
  XOR U6342 ( .A(n6632), .B(n6633), .Z(n6628) );
  AND U6343 ( .A(n6634), .B(n6635), .Z(n6633) );
  XNOR U6344 ( .A(p_input[3390]), .B(n6632), .Z(n6635) );
  XOR U6345 ( .A(n6632), .B(p_input[3374]), .Z(n6634) );
  XOR U6346 ( .A(n6636), .B(n6637), .Z(n6632) );
  AND U6347 ( .A(n6638), .B(n6639), .Z(n6637) );
  XNOR U6348 ( .A(p_input[3389]), .B(n6636), .Z(n6639) );
  XOR U6349 ( .A(n6636), .B(p_input[3373]), .Z(n6638) );
  XOR U6350 ( .A(n6640), .B(n6641), .Z(n6636) );
  AND U6351 ( .A(n6642), .B(n6643), .Z(n6641) );
  XNOR U6352 ( .A(p_input[3388]), .B(n6640), .Z(n6643) );
  XOR U6353 ( .A(n6640), .B(p_input[3372]), .Z(n6642) );
  XOR U6354 ( .A(n6644), .B(n6645), .Z(n6640) );
  AND U6355 ( .A(n6646), .B(n6647), .Z(n6645) );
  XNOR U6356 ( .A(p_input[3387]), .B(n6644), .Z(n6647) );
  XOR U6357 ( .A(n6644), .B(p_input[3371]), .Z(n6646) );
  XOR U6358 ( .A(n6648), .B(n6649), .Z(n6644) );
  AND U6359 ( .A(n6650), .B(n6651), .Z(n6649) );
  XNOR U6360 ( .A(p_input[3386]), .B(n6648), .Z(n6651) );
  XOR U6361 ( .A(n6648), .B(p_input[3370]), .Z(n6650) );
  XOR U6362 ( .A(n6652), .B(n6653), .Z(n6648) );
  AND U6363 ( .A(n6654), .B(n6655), .Z(n6653) );
  XNOR U6364 ( .A(p_input[3385]), .B(n6652), .Z(n6655) );
  XOR U6365 ( .A(n6652), .B(p_input[3369]), .Z(n6654) );
  XOR U6366 ( .A(n6656), .B(n6657), .Z(n6652) );
  AND U6367 ( .A(n6658), .B(n6659), .Z(n6657) );
  XNOR U6368 ( .A(p_input[3384]), .B(n6656), .Z(n6659) );
  XOR U6369 ( .A(n6656), .B(p_input[3368]), .Z(n6658) );
  XOR U6370 ( .A(n6660), .B(n6661), .Z(n6656) );
  AND U6371 ( .A(n6662), .B(n6663), .Z(n6661) );
  XNOR U6372 ( .A(p_input[3383]), .B(n6660), .Z(n6663) );
  XOR U6373 ( .A(n6660), .B(p_input[3367]), .Z(n6662) );
  XOR U6374 ( .A(n6664), .B(n6665), .Z(n6660) );
  AND U6375 ( .A(n6666), .B(n6667), .Z(n6665) );
  XNOR U6376 ( .A(p_input[3382]), .B(n6664), .Z(n6667) );
  XOR U6377 ( .A(n6664), .B(p_input[3366]), .Z(n6666) );
  XOR U6378 ( .A(n6668), .B(n6669), .Z(n6664) );
  AND U6379 ( .A(n6670), .B(n6671), .Z(n6669) );
  XNOR U6380 ( .A(p_input[3381]), .B(n6668), .Z(n6671) );
  XOR U6381 ( .A(n6668), .B(p_input[3365]), .Z(n6670) );
  XOR U6382 ( .A(n6672), .B(n6673), .Z(n6668) );
  AND U6383 ( .A(n6674), .B(n6675), .Z(n6673) );
  XNOR U6384 ( .A(p_input[3380]), .B(n6672), .Z(n6675) );
  XOR U6385 ( .A(n6672), .B(p_input[3364]), .Z(n6674) );
  XOR U6386 ( .A(n6676), .B(n6677), .Z(n6672) );
  AND U6387 ( .A(n6678), .B(n6679), .Z(n6677) );
  XNOR U6388 ( .A(p_input[3379]), .B(n6676), .Z(n6679) );
  XOR U6389 ( .A(n6676), .B(p_input[3363]), .Z(n6678) );
  XOR U6390 ( .A(n6680), .B(n6681), .Z(n6676) );
  AND U6391 ( .A(n6682), .B(n6683), .Z(n6681) );
  XNOR U6392 ( .A(p_input[3378]), .B(n6680), .Z(n6683) );
  XOR U6393 ( .A(n6680), .B(p_input[3362]), .Z(n6682) );
  XNOR U6394 ( .A(n6684), .B(n6685), .Z(n6680) );
  AND U6395 ( .A(n6686), .B(n6687), .Z(n6685) );
  XOR U6396 ( .A(p_input[3377]), .B(n6684), .Z(n6687) );
  XNOR U6397 ( .A(p_input[3361]), .B(n6684), .Z(n6686) );
  AND U6398 ( .A(p_input[3376]), .B(n6688), .Z(n6684) );
  IV U6399 ( .A(p_input[3360]), .Z(n6688) );
  XNOR U6400 ( .A(p_input[3328]), .B(n6689), .Z(n6491) );
  AND U6401 ( .A(n180), .B(n6690), .Z(n6689) );
  XOR U6402 ( .A(p_input[3344]), .B(p_input[3328]), .Z(n6690) );
  XOR U6403 ( .A(n6691), .B(n6692), .Z(n180) );
  AND U6404 ( .A(n6693), .B(n6694), .Z(n6692) );
  XNOR U6405 ( .A(p_input[3359]), .B(n6691), .Z(n6694) );
  XOR U6406 ( .A(n6691), .B(p_input[3343]), .Z(n6693) );
  XOR U6407 ( .A(n6695), .B(n6696), .Z(n6691) );
  AND U6408 ( .A(n6697), .B(n6698), .Z(n6696) );
  XNOR U6409 ( .A(p_input[3358]), .B(n6695), .Z(n6698) );
  XNOR U6410 ( .A(n6695), .B(n6505), .Z(n6697) );
  IV U6411 ( .A(p_input[3342]), .Z(n6505) );
  XOR U6412 ( .A(n6699), .B(n6700), .Z(n6695) );
  AND U6413 ( .A(n6701), .B(n6702), .Z(n6700) );
  XNOR U6414 ( .A(p_input[3357]), .B(n6699), .Z(n6702) );
  XNOR U6415 ( .A(n6699), .B(n6514), .Z(n6701) );
  IV U6416 ( .A(p_input[3341]), .Z(n6514) );
  XOR U6417 ( .A(n6703), .B(n6704), .Z(n6699) );
  AND U6418 ( .A(n6705), .B(n6706), .Z(n6704) );
  XNOR U6419 ( .A(p_input[3356]), .B(n6703), .Z(n6706) );
  XNOR U6420 ( .A(n6703), .B(n6523), .Z(n6705) );
  IV U6421 ( .A(p_input[3340]), .Z(n6523) );
  XOR U6422 ( .A(n6707), .B(n6708), .Z(n6703) );
  AND U6423 ( .A(n6709), .B(n6710), .Z(n6708) );
  XNOR U6424 ( .A(p_input[3355]), .B(n6707), .Z(n6710) );
  XNOR U6425 ( .A(n6707), .B(n6532), .Z(n6709) );
  IV U6426 ( .A(p_input[3339]), .Z(n6532) );
  XOR U6427 ( .A(n6711), .B(n6712), .Z(n6707) );
  AND U6428 ( .A(n6713), .B(n6714), .Z(n6712) );
  XNOR U6429 ( .A(p_input[3354]), .B(n6711), .Z(n6714) );
  XNOR U6430 ( .A(n6711), .B(n6541), .Z(n6713) );
  IV U6431 ( .A(p_input[3338]), .Z(n6541) );
  XOR U6432 ( .A(n6715), .B(n6716), .Z(n6711) );
  AND U6433 ( .A(n6717), .B(n6718), .Z(n6716) );
  XNOR U6434 ( .A(p_input[3353]), .B(n6715), .Z(n6718) );
  XNOR U6435 ( .A(n6715), .B(n6550), .Z(n6717) );
  IV U6436 ( .A(p_input[3337]), .Z(n6550) );
  XOR U6437 ( .A(n6719), .B(n6720), .Z(n6715) );
  AND U6438 ( .A(n6721), .B(n6722), .Z(n6720) );
  XNOR U6439 ( .A(p_input[3352]), .B(n6719), .Z(n6722) );
  XNOR U6440 ( .A(n6719), .B(n6559), .Z(n6721) );
  IV U6441 ( .A(p_input[3336]), .Z(n6559) );
  XOR U6442 ( .A(n6723), .B(n6724), .Z(n6719) );
  AND U6443 ( .A(n6725), .B(n6726), .Z(n6724) );
  XNOR U6444 ( .A(p_input[3351]), .B(n6723), .Z(n6726) );
  XNOR U6445 ( .A(n6723), .B(n6568), .Z(n6725) );
  IV U6446 ( .A(p_input[3335]), .Z(n6568) );
  XOR U6447 ( .A(n6727), .B(n6728), .Z(n6723) );
  AND U6448 ( .A(n6729), .B(n6730), .Z(n6728) );
  XNOR U6449 ( .A(p_input[3350]), .B(n6727), .Z(n6730) );
  XNOR U6450 ( .A(n6727), .B(n6577), .Z(n6729) );
  IV U6451 ( .A(p_input[3334]), .Z(n6577) );
  XOR U6452 ( .A(n6731), .B(n6732), .Z(n6727) );
  AND U6453 ( .A(n6733), .B(n6734), .Z(n6732) );
  XNOR U6454 ( .A(p_input[3349]), .B(n6731), .Z(n6734) );
  XNOR U6455 ( .A(n6731), .B(n6586), .Z(n6733) );
  IV U6456 ( .A(p_input[3333]), .Z(n6586) );
  XOR U6457 ( .A(n6735), .B(n6736), .Z(n6731) );
  AND U6458 ( .A(n6737), .B(n6738), .Z(n6736) );
  XNOR U6459 ( .A(p_input[3348]), .B(n6735), .Z(n6738) );
  XNOR U6460 ( .A(n6735), .B(n6595), .Z(n6737) );
  IV U6461 ( .A(p_input[3332]), .Z(n6595) );
  XOR U6462 ( .A(n6739), .B(n6740), .Z(n6735) );
  AND U6463 ( .A(n6741), .B(n6742), .Z(n6740) );
  XNOR U6464 ( .A(p_input[3347]), .B(n6739), .Z(n6742) );
  XNOR U6465 ( .A(n6739), .B(n6604), .Z(n6741) );
  IV U6466 ( .A(p_input[3331]), .Z(n6604) );
  XOR U6467 ( .A(n6743), .B(n6744), .Z(n6739) );
  AND U6468 ( .A(n6745), .B(n6746), .Z(n6744) );
  XNOR U6469 ( .A(p_input[3346]), .B(n6743), .Z(n6746) );
  XNOR U6470 ( .A(n6743), .B(n6613), .Z(n6745) );
  IV U6471 ( .A(p_input[3330]), .Z(n6613) );
  XNOR U6472 ( .A(n6747), .B(n6748), .Z(n6743) );
  AND U6473 ( .A(n6749), .B(n6750), .Z(n6748) );
  XOR U6474 ( .A(p_input[3345]), .B(n6747), .Z(n6750) );
  XNOR U6475 ( .A(p_input[3329]), .B(n6747), .Z(n6749) );
  AND U6476 ( .A(p_input[3344]), .B(n6751), .Z(n6747) );
  IV U6477 ( .A(p_input[3328]), .Z(n6751) );
  XOR U6478 ( .A(n6752), .B(n6753), .Z(n4979) );
  AND U6479 ( .A(n920), .B(n6754), .Z(n6753) );
  XNOR U6480 ( .A(n6755), .B(n6752), .Z(n6754) );
  XOR U6481 ( .A(n6756), .B(n6757), .Z(n920) );
  AND U6482 ( .A(n6758), .B(n6759), .Z(n6757) );
  XNOR U6483 ( .A(n4994), .B(n6756), .Z(n6759) );
  AND U6484 ( .A(n6760), .B(n6761), .Z(n4994) );
  XNOR U6485 ( .A(n6756), .B(n4991), .Z(n6758) );
  IV U6486 ( .A(n6762), .Z(n4991) );
  AND U6487 ( .A(n6763), .B(n6764), .Z(n6762) );
  XOR U6488 ( .A(n6765), .B(n6766), .Z(n6756) );
  AND U6489 ( .A(n6767), .B(n6768), .Z(n6766) );
  XOR U6490 ( .A(n6765), .B(n5006), .Z(n6768) );
  XOR U6491 ( .A(n6769), .B(n6770), .Z(n5006) );
  AND U6492 ( .A(n751), .B(n6771), .Z(n6770) );
  XOR U6493 ( .A(n6772), .B(n6769), .Z(n6771) );
  XNOR U6494 ( .A(n5003), .B(n6765), .Z(n6767) );
  XOR U6495 ( .A(n6773), .B(n6774), .Z(n5003) );
  AND U6496 ( .A(n748), .B(n6775), .Z(n6774) );
  XOR U6497 ( .A(n6776), .B(n6773), .Z(n6775) );
  XOR U6498 ( .A(n6777), .B(n6778), .Z(n6765) );
  AND U6499 ( .A(n6779), .B(n6780), .Z(n6778) );
  XOR U6500 ( .A(n6777), .B(n5018), .Z(n6780) );
  XOR U6501 ( .A(n6781), .B(n6782), .Z(n5018) );
  AND U6502 ( .A(n751), .B(n6783), .Z(n6782) );
  XOR U6503 ( .A(n6784), .B(n6781), .Z(n6783) );
  XNOR U6504 ( .A(n5015), .B(n6777), .Z(n6779) );
  XOR U6505 ( .A(n6785), .B(n6786), .Z(n5015) );
  AND U6506 ( .A(n748), .B(n6787), .Z(n6786) );
  XOR U6507 ( .A(n6788), .B(n6785), .Z(n6787) );
  XOR U6508 ( .A(n6789), .B(n6790), .Z(n6777) );
  AND U6509 ( .A(n6791), .B(n6792), .Z(n6790) );
  XOR U6510 ( .A(n6789), .B(n5030), .Z(n6792) );
  XOR U6511 ( .A(n6793), .B(n6794), .Z(n5030) );
  AND U6512 ( .A(n751), .B(n6795), .Z(n6794) );
  XOR U6513 ( .A(n6796), .B(n6793), .Z(n6795) );
  XNOR U6514 ( .A(n5027), .B(n6789), .Z(n6791) );
  XOR U6515 ( .A(n6797), .B(n6798), .Z(n5027) );
  AND U6516 ( .A(n748), .B(n6799), .Z(n6798) );
  XOR U6517 ( .A(n6800), .B(n6797), .Z(n6799) );
  XOR U6518 ( .A(n6801), .B(n6802), .Z(n6789) );
  AND U6519 ( .A(n6803), .B(n6804), .Z(n6802) );
  XOR U6520 ( .A(n6801), .B(n5042), .Z(n6804) );
  XOR U6521 ( .A(n6805), .B(n6806), .Z(n5042) );
  AND U6522 ( .A(n751), .B(n6807), .Z(n6806) );
  XOR U6523 ( .A(n6808), .B(n6805), .Z(n6807) );
  XNOR U6524 ( .A(n5039), .B(n6801), .Z(n6803) );
  XOR U6525 ( .A(n6809), .B(n6810), .Z(n5039) );
  AND U6526 ( .A(n748), .B(n6811), .Z(n6810) );
  XOR U6527 ( .A(n6812), .B(n6809), .Z(n6811) );
  XOR U6528 ( .A(n6813), .B(n6814), .Z(n6801) );
  AND U6529 ( .A(n6815), .B(n6816), .Z(n6814) );
  XOR U6530 ( .A(n6813), .B(n5054), .Z(n6816) );
  XOR U6531 ( .A(n6817), .B(n6818), .Z(n5054) );
  AND U6532 ( .A(n751), .B(n6819), .Z(n6818) );
  XOR U6533 ( .A(n6820), .B(n6817), .Z(n6819) );
  XNOR U6534 ( .A(n5051), .B(n6813), .Z(n6815) );
  XOR U6535 ( .A(n6821), .B(n6822), .Z(n5051) );
  AND U6536 ( .A(n748), .B(n6823), .Z(n6822) );
  XOR U6537 ( .A(n6824), .B(n6821), .Z(n6823) );
  XOR U6538 ( .A(n6825), .B(n6826), .Z(n6813) );
  AND U6539 ( .A(n6827), .B(n6828), .Z(n6826) );
  XOR U6540 ( .A(n6825), .B(n5066), .Z(n6828) );
  XOR U6541 ( .A(n6829), .B(n6830), .Z(n5066) );
  AND U6542 ( .A(n751), .B(n6831), .Z(n6830) );
  XOR U6543 ( .A(n6832), .B(n6829), .Z(n6831) );
  XNOR U6544 ( .A(n5063), .B(n6825), .Z(n6827) );
  XOR U6545 ( .A(n6833), .B(n6834), .Z(n5063) );
  AND U6546 ( .A(n748), .B(n6835), .Z(n6834) );
  XOR U6547 ( .A(n6836), .B(n6833), .Z(n6835) );
  XOR U6548 ( .A(n6837), .B(n6838), .Z(n6825) );
  AND U6549 ( .A(n6839), .B(n6840), .Z(n6838) );
  XOR U6550 ( .A(n6837), .B(n5078), .Z(n6840) );
  XOR U6551 ( .A(n6841), .B(n6842), .Z(n5078) );
  AND U6552 ( .A(n751), .B(n6843), .Z(n6842) );
  XOR U6553 ( .A(n6844), .B(n6841), .Z(n6843) );
  XNOR U6554 ( .A(n5075), .B(n6837), .Z(n6839) );
  XOR U6555 ( .A(n6845), .B(n6846), .Z(n5075) );
  AND U6556 ( .A(n748), .B(n6847), .Z(n6846) );
  XOR U6557 ( .A(n6848), .B(n6845), .Z(n6847) );
  XOR U6558 ( .A(n6849), .B(n6850), .Z(n6837) );
  AND U6559 ( .A(n6851), .B(n6852), .Z(n6850) );
  XOR U6560 ( .A(n6849), .B(n5090), .Z(n6852) );
  XOR U6561 ( .A(n6853), .B(n6854), .Z(n5090) );
  AND U6562 ( .A(n751), .B(n6855), .Z(n6854) );
  XOR U6563 ( .A(n6856), .B(n6853), .Z(n6855) );
  XNOR U6564 ( .A(n5087), .B(n6849), .Z(n6851) );
  XOR U6565 ( .A(n6857), .B(n6858), .Z(n5087) );
  AND U6566 ( .A(n748), .B(n6859), .Z(n6858) );
  XOR U6567 ( .A(n6860), .B(n6857), .Z(n6859) );
  XOR U6568 ( .A(n6861), .B(n6862), .Z(n6849) );
  AND U6569 ( .A(n6863), .B(n6864), .Z(n6862) );
  XOR U6570 ( .A(n6861), .B(n5102), .Z(n6864) );
  XOR U6571 ( .A(n6865), .B(n6866), .Z(n5102) );
  AND U6572 ( .A(n751), .B(n6867), .Z(n6866) );
  XOR U6573 ( .A(n6868), .B(n6865), .Z(n6867) );
  XNOR U6574 ( .A(n5099), .B(n6861), .Z(n6863) );
  XOR U6575 ( .A(n6869), .B(n6870), .Z(n5099) );
  AND U6576 ( .A(n748), .B(n6871), .Z(n6870) );
  XOR U6577 ( .A(n6872), .B(n6869), .Z(n6871) );
  XOR U6578 ( .A(n6873), .B(n6874), .Z(n6861) );
  AND U6579 ( .A(n6875), .B(n6876), .Z(n6874) );
  XOR U6580 ( .A(n6873), .B(n5114), .Z(n6876) );
  XOR U6581 ( .A(n6877), .B(n6878), .Z(n5114) );
  AND U6582 ( .A(n751), .B(n6879), .Z(n6878) );
  XOR U6583 ( .A(n6880), .B(n6877), .Z(n6879) );
  XNOR U6584 ( .A(n5111), .B(n6873), .Z(n6875) );
  XOR U6585 ( .A(n6881), .B(n6882), .Z(n5111) );
  AND U6586 ( .A(n748), .B(n6883), .Z(n6882) );
  XOR U6587 ( .A(n6884), .B(n6881), .Z(n6883) );
  XOR U6588 ( .A(n6885), .B(n6886), .Z(n6873) );
  AND U6589 ( .A(n6887), .B(n6888), .Z(n6886) );
  XOR U6590 ( .A(n6885), .B(n5126), .Z(n6888) );
  XOR U6591 ( .A(n6889), .B(n6890), .Z(n5126) );
  AND U6592 ( .A(n751), .B(n6891), .Z(n6890) );
  XOR U6593 ( .A(n6892), .B(n6889), .Z(n6891) );
  XNOR U6594 ( .A(n5123), .B(n6885), .Z(n6887) );
  XOR U6595 ( .A(n6893), .B(n6894), .Z(n5123) );
  AND U6596 ( .A(n748), .B(n6895), .Z(n6894) );
  XOR U6597 ( .A(n6896), .B(n6893), .Z(n6895) );
  XOR U6598 ( .A(n6897), .B(n6898), .Z(n6885) );
  AND U6599 ( .A(n6899), .B(n6900), .Z(n6898) );
  XOR U6600 ( .A(n6897), .B(n5138), .Z(n6900) );
  XOR U6601 ( .A(n6901), .B(n6902), .Z(n5138) );
  AND U6602 ( .A(n751), .B(n6903), .Z(n6902) );
  XOR U6603 ( .A(n6904), .B(n6901), .Z(n6903) );
  XNOR U6604 ( .A(n5135), .B(n6897), .Z(n6899) );
  XOR U6605 ( .A(n6905), .B(n6906), .Z(n5135) );
  AND U6606 ( .A(n748), .B(n6907), .Z(n6906) );
  XOR U6607 ( .A(n6908), .B(n6905), .Z(n6907) );
  XOR U6608 ( .A(n6909), .B(n6910), .Z(n6897) );
  AND U6609 ( .A(n6911), .B(n6912), .Z(n6910) );
  XOR U6610 ( .A(n6909), .B(n5150), .Z(n6912) );
  XOR U6611 ( .A(n6913), .B(n6914), .Z(n5150) );
  AND U6612 ( .A(n751), .B(n6915), .Z(n6914) );
  XOR U6613 ( .A(n6916), .B(n6913), .Z(n6915) );
  XNOR U6614 ( .A(n5147), .B(n6909), .Z(n6911) );
  XOR U6615 ( .A(n6917), .B(n6918), .Z(n5147) );
  AND U6616 ( .A(n748), .B(n6919), .Z(n6918) );
  XOR U6617 ( .A(n6920), .B(n6917), .Z(n6919) );
  XOR U6618 ( .A(n6921), .B(n6922), .Z(n6909) );
  AND U6619 ( .A(n6923), .B(n6924), .Z(n6922) );
  XNOR U6620 ( .A(n6925), .B(n5163), .Z(n6924) );
  XOR U6621 ( .A(n6926), .B(n6927), .Z(n5163) );
  AND U6622 ( .A(n751), .B(n6928), .Z(n6927) );
  XOR U6623 ( .A(n6926), .B(n6929), .Z(n6928) );
  XNOR U6624 ( .A(n5160), .B(n6921), .Z(n6923) );
  XOR U6625 ( .A(n6930), .B(n6931), .Z(n5160) );
  AND U6626 ( .A(n748), .B(n6932), .Z(n6931) );
  XOR U6627 ( .A(n6930), .B(n6933), .Z(n6932) );
  IV U6628 ( .A(n6925), .Z(n6921) );
  AND U6629 ( .A(n6752), .B(n6755), .Z(n6925) );
  XNOR U6630 ( .A(n6934), .B(n6935), .Z(n6755) );
  AND U6631 ( .A(n751), .B(n6936), .Z(n6935) );
  XNOR U6632 ( .A(n6937), .B(n6934), .Z(n6936) );
  XOR U6633 ( .A(n6938), .B(n6939), .Z(n751) );
  AND U6634 ( .A(n6940), .B(n6941), .Z(n6939) );
  XNOR U6635 ( .A(n6760), .B(n6938), .Z(n6941) );
  AND U6636 ( .A(n6942), .B(n6943), .Z(n6760) );
  XOR U6637 ( .A(n6938), .B(n6761), .Z(n6940) );
  AND U6638 ( .A(n6944), .B(n6945), .Z(n6761) );
  XOR U6639 ( .A(n6946), .B(n6947), .Z(n6938) );
  AND U6640 ( .A(n6948), .B(n6949), .Z(n6947) );
  XOR U6641 ( .A(n6946), .B(n6772), .Z(n6949) );
  XOR U6642 ( .A(n6950), .B(n6951), .Z(n6772) );
  AND U6643 ( .A(n399), .B(n6952), .Z(n6951) );
  XOR U6644 ( .A(n6953), .B(n6950), .Z(n6952) );
  XNOR U6645 ( .A(n6769), .B(n6946), .Z(n6948) );
  XOR U6646 ( .A(n6954), .B(n6955), .Z(n6769) );
  AND U6647 ( .A(n397), .B(n6956), .Z(n6955) );
  XOR U6648 ( .A(n6957), .B(n6954), .Z(n6956) );
  XOR U6649 ( .A(n6958), .B(n6959), .Z(n6946) );
  AND U6650 ( .A(n6960), .B(n6961), .Z(n6959) );
  XOR U6651 ( .A(n6958), .B(n6784), .Z(n6961) );
  XOR U6652 ( .A(n6962), .B(n6963), .Z(n6784) );
  AND U6653 ( .A(n399), .B(n6964), .Z(n6963) );
  XOR U6654 ( .A(n6965), .B(n6962), .Z(n6964) );
  XNOR U6655 ( .A(n6781), .B(n6958), .Z(n6960) );
  XOR U6656 ( .A(n6966), .B(n6967), .Z(n6781) );
  AND U6657 ( .A(n397), .B(n6968), .Z(n6967) );
  XOR U6658 ( .A(n6969), .B(n6966), .Z(n6968) );
  XOR U6659 ( .A(n6970), .B(n6971), .Z(n6958) );
  AND U6660 ( .A(n6972), .B(n6973), .Z(n6971) );
  XOR U6661 ( .A(n6970), .B(n6796), .Z(n6973) );
  XOR U6662 ( .A(n6974), .B(n6975), .Z(n6796) );
  AND U6663 ( .A(n399), .B(n6976), .Z(n6975) );
  XOR U6664 ( .A(n6977), .B(n6974), .Z(n6976) );
  XNOR U6665 ( .A(n6793), .B(n6970), .Z(n6972) );
  XOR U6666 ( .A(n6978), .B(n6979), .Z(n6793) );
  AND U6667 ( .A(n397), .B(n6980), .Z(n6979) );
  XOR U6668 ( .A(n6981), .B(n6978), .Z(n6980) );
  XOR U6669 ( .A(n6982), .B(n6983), .Z(n6970) );
  AND U6670 ( .A(n6984), .B(n6985), .Z(n6983) );
  XOR U6671 ( .A(n6982), .B(n6808), .Z(n6985) );
  XOR U6672 ( .A(n6986), .B(n6987), .Z(n6808) );
  AND U6673 ( .A(n399), .B(n6988), .Z(n6987) );
  XOR U6674 ( .A(n6989), .B(n6986), .Z(n6988) );
  XNOR U6675 ( .A(n6805), .B(n6982), .Z(n6984) );
  XOR U6676 ( .A(n6990), .B(n6991), .Z(n6805) );
  AND U6677 ( .A(n397), .B(n6992), .Z(n6991) );
  XOR U6678 ( .A(n6993), .B(n6990), .Z(n6992) );
  XOR U6679 ( .A(n6994), .B(n6995), .Z(n6982) );
  AND U6680 ( .A(n6996), .B(n6997), .Z(n6995) );
  XOR U6681 ( .A(n6994), .B(n6820), .Z(n6997) );
  XOR U6682 ( .A(n6998), .B(n6999), .Z(n6820) );
  AND U6683 ( .A(n399), .B(n7000), .Z(n6999) );
  XOR U6684 ( .A(n7001), .B(n6998), .Z(n7000) );
  XNOR U6685 ( .A(n6817), .B(n6994), .Z(n6996) );
  XOR U6686 ( .A(n7002), .B(n7003), .Z(n6817) );
  AND U6687 ( .A(n397), .B(n7004), .Z(n7003) );
  XOR U6688 ( .A(n7005), .B(n7002), .Z(n7004) );
  XOR U6689 ( .A(n7006), .B(n7007), .Z(n6994) );
  AND U6690 ( .A(n7008), .B(n7009), .Z(n7007) );
  XOR U6691 ( .A(n7006), .B(n6832), .Z(n7009) );
  XOR U6692 ( .A(n7010), .B(n7011), .Z(n6832) );
  AND U6693 ( .A(n399), .B(n7012), .Z(n7011) );
  XOR U6694 ( .A(n7013), .B(n7010), .Z(n7012) );
  XNOR U6695 ( .A(n6829), .B(n7006), .Z(n7008) );
  XOR U6696 ( .A(n7014), .B(n7015), .Z(n6829) );
  AND U6697 ( .A(n397), .B(n7016), .Z(n7015) );
  XOR U6698 ( .A(n7017), .B(n7014), .Z(n7016) );
  XOR U6699 ( .A(n7018), .B(n7019), .Z(n7006) );
  AND U6700 ( .A(n7020), .B(n7021), .Z(n7019) );
  XOR U6701 ( .A(n7018), .B(n6844), .Z(n7021) );
  XOR U6702 ( .A(n7022), .B(n7023), .Z(n6844) );
  AND U6703 ( .A(n399), .B(n7024), .Z(n7023) );
  XOR U6704 ( .A(n7025), .B(n7022), .Z(n7024) );
  XNOR U6705 ( .A(n6841), .B(n7018), .Z(n7020) );
  XOR U6706 ( .A(n7026), .B(n7027), .Z(n6841) );
  AND U6707 ( .A(n397), .B(n7028), .Z(n7027) );
  XOR U6708 ( .A(n7029), .B(n7026), .Z(n7028) );
  XOR U6709 ( .A(n7030), .B(n7031), .Z(n7018) );
  AND U6710 ( .A(n7032), .B(n7033), .Z(n7031) );
  XOR U6711 ( .A(n7030), .B(n6856), .Z(n7033) );
  XOR U6712 ( .A(n7034), .B(n7035), .Z(n6856) );
  AND U6713 ( .A(n399), .B(n7036), .Z(n7035) );
  XOR U6714 ( .A(n7037), .B(n7034), .Z(n7036) );
  XNOR U6715 ( .A(n6853), .B(n7030), .Z(n7032) );
  XOR U6716 ( .A(n7038), .B(n7039), .Z(n6853) );
  AND U6717 ( .A(n397), .B(n7040), .Z(n7039) );
  XOR U6718 ( .A(n7041), .B(n7038), .Z(n7040) );
  XOR U6719 ( .A(n7042), .B(n7043), .Z(n7030) );
  AND U6720 ( .A(n7044), .B(n7045), .Z(n7043) );
  XOR U6721 ( .A(n7042), .B(n6868), .Z(n7045) );
  XOR U6722 ( .A(n7046), .B(n7047), .Z(n6868) );
  AND U6723 ( .A(n399), .B(n7048), .Z(n7047) );
  XOR U6724 ( .A(n7049), .B(n7046), .Z(n7048) );
  XNOR U6725 ( .A(n6865), .B(n7042), .Z(n7044) );
  XOR U6726 ( .A(n7050), .B(n7051), .Z(n6865) );
  AND U6727 ( .A(n397), .B(n7052), .Z(n7051) );
  XOR U6728 ( .A(n7053), .B(n7050), .Z(n7052) );
  XOR U6729 ( .A(n7054), .B(n7055), .Z(n7042) );
  AND U6730 ( .A(n7056), .B(n7057), .Z(n7055) );
  XOR U6731 ( .A(n7054), .B(n6880), .Z(n7057) );
  XOR U6732 ( .A(n7058), .B(n7059), .Z(n6880) );
  AND U6733 ( .A(n399), .B(n7060), .Z(n7059) );
  XOR U6734 ( .A(n7061), .B(n7058), .Z(n7060) );
  XNOR U6735 ( .A(n6877), .B(n7054), .Z(n7056) );
  XOR U6736 ( .A(n7062), .B(n7063), .Z(n6877) );
  AND U6737 ( .A(n397), .B(n7064), .Z(n7063) );
  XOR U6738 ( .A(n7065), .B(n7062), .Z(n7064) );
  XOR U6739 ( .A(n7066), .B(n7067), .Z(n7054) );
  AND U6740 ( .A(n7068), .B(n7069), .Z(n7067) );
  XOR U6741 ( .A(n7066), .B(n6892), .Z(n7069) );
  XOR U6742 ( .A(n7070), .B(n7071), .Z(n6892) );
  AND U6743 ( .A(n399), .B(n7072), .Z(n7071) );
  XOR U6744 ( .A(n7073), .B(n7070), .Z(n7072) );
  XNOR U6745 ( .A(n6889), .B(n7066), .Z(n7068) );
  XOR U6746 ( .A(n7074), .B(n7075), .Z(n6889) );
  AND U6747 ( .A(n397), .B(n7076), .Z(n7075) );
  XOR U6748 ( .A(n7077), .B(n7074), .Z(n7076) );
  XOR U6749 ( .A(n7078), .B(n7079), .Z(n7066) );
  AND U6750 ( .A(n7080), .B(n7081), .Z(n7079) );
  XOR U6751 ( .A(n7078), .B(n6904), .Z(n7081) );
  XOR U6752 ( .A(n7082), .B(n7083), .Z(n6904) );
  AND U6753 ( .A(n399), .B(n7084), .Z(n7083) );
  XOR U6754 ( .A(n7085), .B(n7082), .Z(n7084) );
  XNOR U6755 ( .A(n6901), .B(n7078), .Z(n7080) );
  XOR U6756 ( .A(n7086), .B(n7087), .Z(n6901) );
  AND U6757 ( .A(n397), .B(n7088), .Z(n7087) );
  XOR U6758 ( .A(n7089), .B(n7086), .Z(n7088) );
  XOR U6759 ( .A(n7090), .B(n7091), .Z(n7078) );
  AND U6760 ( .A(n7092), .B(n7093), .Z(n7091) );
  XOR U6761 ( .A(n7090), .B(n6916), .Z(n7093) );
  XOR U6762 ( .A(n7094), .B(n7095), .Z(n6916) );
  AND U6763 ( .A(n399), .B(n7096), .Z(n7095) );
  XOR U6764 ( .A(n7097), .B(n7094), .Z(n7096) );
  XNOR U6765 ( .A(n6913), .B(n7090), .Z(n7092) );
  XOR U6766 ( .A(n7098), .B(n7099), .Z(n6913) );
  AND U6767 ( .A(n397), .B(n7100), .Z(n7099) );
  XOR U6768 ( .A(n7101), .B(n7098), .Z(n7100) );
  XOR U6769 ( .A(n7102), .B(n7103), .Z(n7090) );
  AND U6770 ( .A(n7104), .B(n7105), .Z(n7103) );
  XNOR U6771 ( .A(n7106), .B(n6929), .Z(n7105) );
  XOR U6772 ( .A(n7107), .B(n7108), .Z(n6929) );
  AND U6773 ( .A(n399), .B(n7109), .Z(n7108) );
  XOR U6774 ( .A(n7107), .B(n7110), .Z(n7109) );
  XNOR U6775 ( .A(n6926), .B(n7102), .Z(n7104) );
  XOR U6776 ( .A(n7111), .B(n7112), .Z(n6926) );
  AND U6777 ( .A(n397), .B(n7113), .Z(n7112) );
  XOR U6778 ( .A(n7111), .B(n7114), .Z(n7113) );
  IV U6779 ( .A(n7106), .Z(n7102) );
  AND U6780 ( .A(n6934), .B(n6937), .Z(n7106) );
  XNOR U6781 ( .A(n7115), .B(n7116), .Z(n6937) );
  AND U6782 ( .A(n399), .B(n7117), .Z(n7116) );
  XNOR U6783 ( .A(n7118), .B(n7115), .Z(n7117) );
  XOR U6784 ( .A(n7119), .B(n7120), .Z(n399) );
  AND U6785 ( .A(n7121), .B(n7122), .Z(n7120) );
  XNOR U6786 ( .A(n6942), .B(n7119), .Z(n7122) );
  AND U6787 ( .A(p_input[3327]), .B(p_input[3311]), .Z(n6942) );
  XOR U6788 ( .A(n7119), .B(n6943), .Z(n7121) );
  AND U6789 ( .A(p_input[3295]), .B(p_input[3279]), .Z(n6943) );
  XOR U6790 ( .A(n7123), .B(n7124), .Z(n7119) );
  AND U6791 ( .A(n7125), .B(n7126), .Z(n7124) );
  XOR U6792 ( .A(n7123), .B(n6953), .Z(n7126) );
  XNOR U6793 ( .A(p_input[3310]), .B(n7127), .Z(n6953) );
  AND U6794 ( .A(n195), .B(n7128), .Z(n7127) );
  XOR U6795 ( .A(p_input[3326]), .B(p_input[3310]), .Z(n7128) );
  XNOR U6796 ( .A(n6950), .B(n7123), .Z(n7125) );
  XOR U6797 ( .A(n7129), .B(n7130), .Z(n6950) );
  AND U6798 ( .A(n193), .B(n7131), .Z(n7130) );
  XOR U6799 ( .A(p_input[3294]), .B(p_input[3278]), .Z(n7131) );
  XOR U6800 ( .A(n7132), .B(n7133), .Z(n7123) );
  AND U6801 ( .A(n7134), .B(n7135), .Z(n7133) );
  XOR U6802 ( .A(n7132), .B(n6965), .Z(n7135) );
  XNOR U6803 ( .A(p_input[3309]), .B(n7136), .Z(n6965) );
  AND U6804 ( .A(n195), .B(n7137), .Z(n7136) );
  XOR U6805 ( .A(p_input[3325]), .B(p_input[3309]), .Z(n7137) );
  XNOR U6806 ( .A(n6962), .B(n7132), .Z(n7134) );
  XOR U6807 ( .A(n7138), .B(n7139), .Z(n6962) );
  AND U6808 ( .A(n193), .B(n7140), .Z(n7139) );
  XOR U6809 ( .A(p_input[3293]), .B(p_input[3277]), .Z(n7140) );
  XOR U6810 ( .A(n7141), .B(n7142), .Z(n7132) );
  AND U6811 ( .A(n7143), .B(n7144), .Z(n7142) );
  XOR U6812 ( .A(n7141), .B(n6977), .Z(n7144) );
  XNOR U6813 ( .A(p_input[3308]), .B(n7145), .Z(n6977) );
  AND U6814 ( .A(n195), .B(n7146), .Z(n7145) );
  XOR U6815 ( .A(p_input[3324]), .B(p_input[3308]), .Z(n7146) );
  XNOR U6816 ( .A(n6974), .B(n7141), .Z(n7143) );
  XOR U6817 ( .A(n7147), .B(n7148), .Z(n6974) );
  AND U6818 ( .A(n193), .B(n7149), .Z(n7148) );
  XOR U6819 ( .A(p_input[3292]), .B(p_input[3276]), .Z(n7149) );
  XOR U6820 ( .A(n7150), .B(n7151), .Z(n7141) );
  AND U6821 ( .A(n7152), .B(n7153), .Z(n7151) );
  XOR U6822 ( .A(n7150), .B(n6989), .Z(n7153) );
  XNOR U6823 ( .A(p_input[3307]), .B(n7154), .Z(n6989) );
  AND U6824 ( .A(n195), .B(n7155), .Z(n7154) );
  XOR U6825 ( .A(p_input[3323]), .B(p_input[3307]), .Z(n7155) );
  XNOR U6826 ( .A(n6986), .B(n7150), .Z(n7152) );
  XOR U6827 ( .A(n7156), .B(n7157), .Z(n6986) );
  AND U6828 ( .A(n193), .B(n7158), .Z(n7157) );
  XOR U6829 ( .A(p_input[3291]), .B(p_input[3275]), .Z(n7158) );
  XOR U6830 ( .A(n7159), .B(n7160), .Z(n7150) );
  AND U6831 ( .A(n7161), .B(n7162), .Z(n7160) );
  XOR U6832 ( .A(n7159), .B(n7001), .Z(n7162) );
  XNOR U6833 ( .A(p_input[3306]), .B(n7163), .Z(n7001) );
  AND U6834 ( .A(n195), .B(n7164), .Z(n7163) );
  XOR U6835 ( .A(p_input[3322]), .B(p_input[3306]), .Z(n7164) );
  XNOR U6836 ( .A(n6998), .B(n7159), .Z(n7161) );
  XOR U6837 ( .A(n7165), .B(n7166), .Z(n6998) );
  AND U6838 ( .A(n193), .B(n7167), .Z(n7166) );
  XOR U6839 ( .A(p_input[3290]), .B(p_input[3274]), .Z(n7167) );
  XOR U6840 ( .A(n7168), .B(n7169), .Z(n7159) );
  AND U6841 ( .A(n7170), .B(n7171), .Z(n7169) );
  XOR U6842 ( .A(n7168), .B(n7013), .Z(n7171) );
  XNOR U6843 ( .A(p_input[3305]), .B(n7172), .Z(n7013) );
  AND U6844 ( .A(n195), .B(n7173), .Z(n7172) );
  XOR U6845 ( .A(p_input[3321]), .B(p_input[3305]), .Z(n7173) );
  XNOR U6846 ( .A(n7010), .B(n7168), .Z(n7170) );
  XOR U6847 ( .A(n7174), .B(n7175), .Z(n7010) );
  AND U6848 ( .A(n193), .B(n7176), .Z(n7175) );
  XOR U6849 ( .A(p_input[3289]), .B(p_input[3273]), .Z(n7176) );
  XOR U6850 ( .A(n7177), .B(n7178), .Z(n7168) );
  AND U6851 ( .A(n7179), .B(n7180), .Z(n7178) );
  XOR U6852 ( .A(n7177), .B(n7025), .Z(n7180) );
  XNOR U6853 ( .A(p_input[3304]), .B(n7181), .Z(n7025) );
  AND U6854 ( .A(n195), .B(n7182), .Z(n7181) );
  XOR U6855 ( .A(p_input[3320]), .B(p_input[3304]), .Z(n7182) );
  XNOR U6856 ( .A(n7022), .B(n7177), .Z(n7179) );
  XOR U6857 ( .A(n7183), .B(n7184), .Z(n7022) );
  AND U6858 ( .A(n193), .B(n7185), .Z(n7184) );
  XOR U6859 ( .A(p_input[3288]), .B(p_input[3272]), .Z(n7185) );
  XOR U6860 ( .A(n7186), .B(n7187), .Z(n7177) );
  AND U6861 ( .A(n7188), .B(n7189), .Z(n7187) );
  XOR U6862 ( .A(n7186), .B(n7037), .Z(n7189) );
  XNOR U6863 ( .A(p_input[3303]), .B(n7190), .Z(n7037) );
  AND U6864 ( .A(n195), .B(n7191), .Z(n7190) );
  XOR U6865 ( .A(p_input[3319]), .B(p_input[3303]), .Z(n7191) );
  XNOR U6866 ( .A(n7034), .B(n7186), .Z(n7188) );
  XOR U6867 ( .A(n7192), .B(n7193), .Z(n7034) );
  AND U6868 ( .A(n193), .B(n7194), .Z(n7193) );
  XOR U6869 ( .A(p_input[3287]), .B(p_input[3271]), .Z(n7194) );
  XOR U6870 ( .A(n7195), .B(n7196), .Z(n7186) );
  AND U6871 ( .A(n7197), .B(n7198), .Z(n7196) );
  XOR U6872 ( .A(n7195), .B(n7049), .Z(n7198) );
  XNOR U6873 ( .A(p_input[3302]), .B(n7199), .Z(n7049) );
  AND U6874 ( .A(n195), .B(n7200), .Z(n7199) );
  XOR U6875 ( .A(p_input[3318]), .B(p_input[3302]), .Z(n7200) );
  XNOR U6876 ( .A(n7046), .B(n7195), .Z(n7197) );
  XOR U6877 ( .A(n7201), .B(n7202), .Z(n7046) );
  AND U6878 ( .A(n193), .B(n7203), .Z(n7202) );
  XOR U6879 ( .A(p_input[3286]), .B(p_input[3270]), .Z(n7203) );
  XOR U6880 ( .A(n7204), .B(n7205), .Z(n7195) );
  AND U6881 ( .A(n7206), .B(n7207), .Z(n7205) );
  XOR U6882 ( .A(n7204), .B(n7061), .Z(n7207) );
  XNOR U6883 ( .A(p_input[3301]), .B(n7208), .Z(n7061) );
  AND U6884 ( .A(n195), .B(n7209), .Z(n7208) );
  XOR U6885 ( .A(p_input[3317]), .B(p_input[3301]), .Z(n7209) );
  XNOR U6886 ( .A(n7058), .B(n7204), .Z(n7206) );
  XOR U6887 ( .A(n7210), .B(n7211), .Z(n7058) );
  AND U6888 ( .A(n193), .B(n7212), .Z(n7211) );
  XOR U6889 ( .A(p_input[3285]), .B(p_input[3269]), .Z(n7212) );
  XOR U6890 ( .A(n7213), .B(n7214), .Z(n7204) );
  AND U6891 ( .A(n7215), .B(n7216), .Z(n7214) );
  XOR U6892 ( .A(n7213), .B(n7073), .Z(n7216) );
  XNOR U6893 ( .A(p_input[3300]), .B(n7217), .Z(n7073) );
  AND U6894 ( .A(n195), .B(n7218), .Z(n7217) );
  XOR U6895 ( .A(p_input[3316]), .B(p_input[3300]), .Z(n7218) );
  XNOR U6896 ( .A(n7070), .B(n7213), .Z(n7215) );
  XOR U6897 ( .A(n7219), .B(n7220), .Z(n7070) );
  AND U6898 ( .A(n193), .B(n7221), .Z(n7220) );
  XOR U6899 ( .A(p_input[3284]), .B(p_input[3268]), .Z(n7221) );
  XOR U6900 ( .A(n7222), .B(n7223), .Z(n7213) );
  AND U6901 ( .A(n7224), .B(n7225), .Z(n7223) );
  XOR U6902 ( .A(n7222), .B(n7085), .Z(n7225) );
  XNOR U6903 ( .A(p_input[3299]), .B(n7226), .Z(n7085) );
  AND U6904 ( .A(n195), .B(n7227), .Z(n7226) );
  XOR U6905 ( .A(p_input[3315]), .B(p_input[3299]), .Z(n7227) );
  XNOR U6906 ( .A(n7082), .B(n7222), .Z(n7224) );
  XOR U6907 ( .A(n7228), .B(n7229), .Z(n7082) );
  AND U6908 ( .A(n193), .B(n7230), .Z(n7229) );
  XOR U6909 ( .A(p_input[3283]), .B(p_input[3267]), .Z(n7230) );
  XOR U6910 ( .A(n7231), .B(n7232), .Z(n7222) );
  AND U6911 ( .A(n7233), .B(n7234), .Z(n7232) );
  XOR U6912 ( .A(n7231), .B(n7097), .Z(n7234) );
  XNOR U6913 ( .A(p_input[3298]), .B(n7235), .Z(n7097) );
  AND U6914 ( .A(n195), .B(n7236), .Z(n7235) );
  XOR U6915 ( .A(p_input[3314]), .B(p_input[3298]), .Z(n7236) );
  XNOR U6916 ( .A(n7094), .B(n7231), .Z(n7233) );
  XOR U6917 ( .A(n7237), .B(n7238), .Z(n7094) );
  AND U6918 ( .A(n193), .B(n7239), .Z(n7238) );
  XOR U6919 ( .A(p_input[3282]), .B(p_input[3266]), .Z(n7239) );
  XOR U6920 ( .A(n7240), .B(n7241), .Z(n7231) );
  AND U6921 ( .A(n7242), .B(n7243), .Z(n7241) );
  XNOR U6922 ( .A(n7244), .B(n7110), .Z(n7243) );
  XNOR U6923 ( .A(p_input[3297]), .B(n7245), .Z(n7110) );
  AND U6924 ( .A(n195), .B(n7246), .Z(n7245) );
  XNOR U6925 ( .A(p_input[3313]), .B(n7247), .Z(n7246) );
  IV U6926 ( .A(p_input[3297]), .Z(n7247) );
  XNOR U6927 ( .A(n7107), .B(n7240), .Z(n7242) );
  XNOR U6928 ( .A(p_input[3265]), .B(n7248), .Z(n7107) );
  AND U6929 ( .A(n193), .B(n7249), .Z(n7248) );
  XOR U6930 ( .A(p_input[3281]), .B(p_input[3265]), .Z(n7249) );
  IV U6931 ( .A(n7244), .Z(n7240) );
  AND U6932 ( .A(n7115), .B(n7118), .Z(n7244) );
  XOR U6933 ( .A(p_input[3296]), .B(n7250), .Z(n7118) );
  AND U6934 ( .A(n195), .B(n7251), .Z(n7250) );
  XOR U6935 ( .A(p_input[3312]), .B(p_input[3296]), .Z(n7251) );
  XOR U6936 ( .A(n7252), .B(n7253), .Z(n195) );
  AND U6937 ( .A(n7254), .B(n7255), .Z(n7253) );
  XNOR U6938 ( .A(p_input[3327]), .B(n7252), .Z(n7255) );
  XOR U6939 ( .A(n7252), .B(p_input[3311]), .Z(n7254) );
  XOR U6940 ( .A(n7256), .B(n7257), .Z(n7252) );
  AND U6941 ( .A(n7258), .B(n7259), .Z(n7257) );
  XNOR U6942 ( .A(p_input[3326]), .B(n7256), .Z(n7259) );
  XOR U6943 ( .A(n7256), .B(p_input[3310]), .Z(n7258) );
  XOR U6944 ( .A(n7260), .B(n7261), .Z(n7256) );
  AND U6945 ( .A(n7262), .B(n7263), .Z(n7261) );
  XNOR U6946 ( .A(p_input[3325]), .B(n7260), .Z(n7263) );
  XOR U6947 ( .A(n7260), .B(p_input[3309]), .Z(n7262) );
  XOR U6948 ( .A(n7264), .B(n7265), .Z(n7260) );
  AND U6949 ( .A(n7266), .B(n7267), .Z(n7265) );
  XNOR U6950 ( .A(p_input[3324]), .B(n7264), .Z(n7267) );
  XOR U6951 ( .A(n7264), .B(p_input[3308]), .Z(n7266) );
  XOR U6952 ( .A(n7268), .B(n7269), .Z(n7264) );
  AND U6953 ( .A(n7270), .B(n7271), .Z(n7269) );
  XNOR U6954 ( .A(p_input[3323]), .B(n7268), .Z(n7271) );
  XOR U6955 ( .A(n7268), .B(p_input[3307]), .Z(n7270) );
  XOR U6956 ( .A(n7272), .B(n7273), .Z(n7268) );
  AND U6957 ( .A(n7274), .B(n7275), .Z(n7273) );
  XNOR U6958 ( .A(p_input[3322]), .B(n7272), .Z(n7275) );
  XOR U6959 ( .A(n7272), .B(p_input[3306]), .Z(n7274) );
  XOR U6960 ( .A(n7276), .B(n7277), .Z(n7272) );
  AND U6961 ( .A(n7278), .B(n7279), .Z(n7277) );
  XNOR U6962 ( .A(p_input[3321]), .B(n7276), .Z(n7279) );
  XOR U6963 ( .A(n7276), .B(p_input[3305]), .Z(n7278) );
  XOR U6964 ( .A(n7280), .B(n7281), .Z(n7276) );
  AND U6965 ( .A(n7282), .B(n7283), .Z(n7281) );
  XNOR U6966 ( .A(p_input[3320]), .B(n7280), .Z(n7283) );
  XOR U6967 ( .A(n7280), .B(p_input[3304]), .Z(n7282) );
  XOR U6968 ( .A(n7284), .B(n7285), .Z(n7280) );
  AND U6969 ( .A(n7286), .B(n7287), .Z(n7285) );
  XNOR U6970 ( .A(p_input[3319]), .B(n7284), .Z(n7287) );
  XOR U6971 ( .A(n7284), .B(p_input[3303]), .Z(n7286) );
  XOR U6972 ( .A(n7288), .B(n7289), .Z(n7284) );
  AND U6973 ( .A(n7290), .B(n7291), .Z(n7289) );
  XNOR U6974 ( .A(p_input[3318]), .B(n7288), .Z(n7291) );
  XOR U6975 ( .A(n7288), .B(p_input[3302]), .Z(n7290) );
  XOR U6976 ( .A(n7292), .B(n7293), .Z(n7288) );
  AND U6977 ( .A(n7294), .B(n7295), .Z(n7293) );
  XNOR U6978 ( .A(p_input[3317]), .B(n7292), .Z(n7295) );
  XOR U6979 ( .A(n7292), .B(p_input[3301]), .Z(n7294) );
  XOR U6980 ( .A(n7296), .B(n7297), .Z(n7292) );
  AND U6981 ( .A(n7298), .B(n7299), .Z(n7297) );
  XNOR U6982 ( .A(p_input[3316]), .B(n7296), .Z(n7299) );
  XOR U6983 ( .A(n7296), .B(p_input[3300]), .Z(n7298) );
  XOR U6984 ( .A(n7300), .B(n7301), .Z(n7296) );
  AND U6985 ( .A(n7302), .B(n7303), .Z(n7301) );
  XNOR U6986 ( .A(p_input[3315]), .B(n7300), .Z(n7303) );
  XOR U6987 ( .A(n7300), .B(p_input[3299]), .Z(n7302) );
  XOR U6988 ( .A(n7304), .B(n7305), .Z(n7300) );
  AND U6989 ( .A(n7306), .B(n7307), .Z(n7305) );
  XNOR U6990 ( .A(p_input[3314]), .B(n7304), .Z(n7307) );
  XOR U6991 ( .A(n7304), .B(p_input[3298]), .Z(n7306) );
  XNOR U6992 ( .A(n7308), .B(n7309), .Z(n7304) );
  AND U6993 ( .A(n7310), .B(n7311), .Z(n7309) );
  XOR U6994 ( .A(p_input[3313]), .B(n7308), .Z(n7311) );
  XNOR U6995 ( .A(p_input[3297]), .B(n7308), .Z(n7310) );
  AND U6996 ( .A(p_input[3312]), .B(n7312), .Z(n7308) );
  IV U6997 ( .A(p_input[3296]), .Z(n7312) );
  XNOR U6998 ( .A(p_input[3264]), .B(n7313), .Z(n7115) );
  AND U6999 ( .A(n193), .B(n7314), .Z(n7313) );
  XOR U7000 ( .A(p_input[3280]), .B(p_input[3264]), .Z(n7314) );
  XOR U7001 ( .A(n7315), .B(n7316), .Z(n193) );
  AND U7002 ( .A(n7317), .B(n7318), .Z(n7316) );
  XNOR U7003 ( .A(p_input[3295]), .B(n7315), .Z(n7318) );
  XOR U7004 ( .A(n7315), .B(p_input[3279]), .Z(n7317) );
  XOR U7005 ( .A(n7319), .B(n7320), .Z(n7315) );
  AND U7006 ( .A(n7321), .B(n7322), .Z(n7320) );
  XNOR U7007 ( .A(p_input[3294]), .B(n7319), .Z(n7322) );
  XNOR U7008 ( .A(n7319), .B(n7129), .Z(n7321) );
  IV U7009 ( .A(p_input[3278]), .Z(n7129) );
  XOR U7010 ( .A(n7323), .B(n7324), .Z(n7319) );
  AND U7011 ( .A(n7325), .B(n7326), .Z(n7324) );
  XNOR U7012 ( .A(p_input[3293]), .B(n7323), .Z(n7326) );
  XNOR U7013 ( .A(n7323), .B(n7138), .Z(n7325) );
  IV U7014 ( .A(p_input[3277]), .Z(n7138) );
  XOR U7015 ( .A(n7327), .B(n7328), .Z(n7323) );
  AND U7016 ( .A(n7329), .B(n7330), .Z(n7328) );
  XNOR U7017 ( .A(p_input[3292]), .B(n7327), .Z(n7330) );
  XNOR U7018 ( .A(n7327), .B(n7147), .Z(n7329) );
  IV U7019 ( .A(p_input[3276]), .Z(n7147) );
  XOR U7020 ( .A(n7331), .B(n7332), .Z(n7327) );
  AND U7021 ( .A(n7333), .B(n7334), .Z(n7332) );
  XNOR U7022 ( .A(p_input[3291]), .B(n7331), .Z(n7334) );
  XNOR U7023 ( .A(n7331), .B(n7156), .Z(n7333) );
  IV U7024 ( .A(p_input[3275]), .Z(n7156) );
  XOR U7025 ( .A(n7335), .B(n7336), .Z(n7331) );
  AND U7026 ( .A(n7337), .B(n7338), .Z(n7336) );
  XNOR U7027 ( .A(p_input[3290]), .B(n7335), .Z(n7338) );
  XNOR U7028 ( .A(n7335), .B(n7165), .Z(n7337) );
  IV U7029 ( .A(p_input[3274]), .Z(n7165) );
  XOR U7030 ( .A(n7339), .B(n7340), .Z(n7335) );
  AND U7031 ( .A(n7341), .B(n7342), .Z(n7340) );
  XNOR U7032 ( .A(p_input[3289]), .B(n7339), .Z(n7342) );
  XNOR U7033 ( .A(n7339), .B(n7174), .Z(n7341) );
  IV U7034 ( .A(p_input[3273]), .Z(n7174) );
  XOR U7035 ( .A(n7343), .B(n7344), .Z(n7339) );
  AND U7036 ( .A(n7345), .B(n7346), .Z(n7344) );
  XNOR U7037 ( .A(p_input[3288]), .B(n7343), .Z(n7346) );
  XNOR U7038 ( .A(n7343), .B(n7183), .Z(n7345) );
  IV U7039 ( .A(p_input[3272]), .Z(n7183) );
  XOR U7040 ( .A(n7347), .B(n7348), .Z(n7343) );
  AND U7041 ( .A(n7349), .B(n7350), .Z(n7348) );
  XNOR U7042 ( .A(p_input[3287]), .B(n7347), .Z(n7350) );
  XNOR U7043 ( .A(n7347), .B(n7192), .Z(n7349) );
  IV U7044 ( .A(p_input[3271]), .Z(n7192) );
  XOR U7045 ( .A(n7351), .B(n7352), .Z(n7347) );
  AND U7046 ( .A(n7353), .B(n7354), .Z(n7352) );
  XNOR U7047 ( .A(p_input[3286]), .B(n7351), .Z(n7354) );
  XNOR U7048 ( .A(n7351), .B(n7201), .Z(n7353) );
  IV U7049 ( .A(p_input[3270]), .Z(n7201) );
  XOR U7050 ( .A(n7355), .B(n7356), .Z(n7351) );
  AND U7051 ( .A(n7357), .B(n7358), .Z(n7356) );
  XNOR U7052 ( .A(p_input[3285]), .B(n7355), .Z(n7358) );
  XNOR U7053 ( .A(n7355), .B(n7210), .Z(n7357) );
  IV U7054 ( .A(p_input[3269]), .Z(n7210) );
  XOR U7055 ( .A(n7359), .B(n7360), .Z(n7355) );
  AND U7056 ( .A(n7361), .B(n7362), .Z(n7360) );
  XNOR U7057 ( .A(p_input[3284]), .B(n7359), .Z(n7362) );
  XNOR U7058 ( .A(n7359), .B(n7219), .Z(n7361) );
  IV U7059 ( .A(p_input[3268]), .Z(n7219) );
  XOR U7060 ( .A(n7363), .B(n7364), .Z(n7359) );
  AND U7061 ( .A(n7365), .B(n7366), .Z(n7364) );
  XNOR U7062 ( .A(p_input[3283]), .B(n7363), .Z(n7366) );
  XNOR U7063 ( .A(n7363), .B(n7228), .Z(n7365) );
  IV U7064 ( .A(p_input[3267]), .Z(n7228) );
  XOR U7065 ( .A(n7367), .B(n7368), .Z(n7363) );
  AND U7066 ( .A(n7369), .B(n7370), .Z(n7368) );
  XNOR U7067 ( .A(p_input[3282]), .B(n7367), .Z(n7370) );
  XNOR U7068 ( .A(n7367), .B(n7237), .Z(n7369) );
  IV U7069 ( .A(p_input[3266]), .Z(n7237) );
  XNOR U7070 ( .A(n7371), .B(n7372), .Z(n7367) );
  AND U7071 ( .A(n7373), .B(n7374), .Z(n7372) );
  XOR U7072 ( .A(p_input[3281]), .B(n7371), .Z(n7374) );
  XNOR U7073 ( .A(p_input[3265]), .B(n7371), .Z(n7373) );
  AND U7074 ( .A(p_input[3280]), .B(n7375), .Z(n7371) );
  IV U7075 ( .A(p_input[3264]), .Z(n7375) );
  XOR U7076 ( .A(n7376), .B(n7377), .Z(n6934) );
  AND U7077 ( .A(n397), .B(n7378), .Z(n7377) );
  XNOR U7078 ( .A(n7379), .B(n7376), .Z(n7378) );
  XOR U7079 ( .A(n7380), .B(n7381), .Z(n397) );
  AND U7080 ( .A(n7382), .B(n7383), .Z(n7381) );
  XNOR U7081 ( .A(n6944), .B(n7380), .Z(n7383) );
  AND U7082 ( .A(p_input[3263]), .B(p_input[3247]), .Z(n6944) );
  XOR U7083 ( .A(n7380), .B(n6945), .Z(n7382) );
  AND U7084 ( .A(p_input[3231]), .B(p_input[3215]), .Z(n6945) );
  XOR U7085 ( .A(n7384), .B(n7385), .Z(n7380) );
  AND U7086 ( .A(n7386), .B(n7387), .Z(n7385) );
  XOR U7087 ( .A(n7384), .B(n6957), .Z(n7387) );
  XNOR U7088 ( .A(p_input[3246]), .B(n7388), .Z(n6957) );
  AND U7089 ( .A(n199), .B(n7389), .Z(n7388) );
  XOR U7090 ( .A(p_input[3262]), .B(p_input[3246]), .Z(n7389) );
  XNOR U7091 ( .A(n6954), .B(n7384), .Z(n7386) );
  XOR U7092 ( .A(n7390), .B(n7391), .Z(n6954) );
  AND U7093 ( .A(n196), .B(n7392), .Z(n7391) );
  XOR U7094 ( .A(p_input[3230]), .B(p_input[3214]), .Z(n7392) );
  XOR U7095 ( .A(n7393), .B(n7394), .Z(n7384) );
  AND U7096 ( .A(n7395), .B(n7396), .Z(n7394) );
  XOR U7097 ( .A(n7393), .B(n6969), .Z(n7396) );
  XNOR U7098 ( .A(p_input[3245]), .B(n7397), .Z(n6969) );
  AND U7099 ( .A(n199), .B(n7398), .Z(n7397) );
  XOR U7100 ( .A(p_input[3261]), .B(p_input[3245]), .Z(n7398) );
  XNOR U7101 ( .A(n6966), .B(n7393), .Z(n7395) );
  XOR U7102 ( .A(n7399), .B(n7400), .Z(n6966) );
  AND U7103 ( .A(n196), .B(n7401), .Z(n7400) );
  XOR U7104 ( .A(p_input[3229]), .B(p_input[3213]), .Z(n7401) );
  XOR U7105 ( .A(n7402), .B(n7403), .Z(n7393) );
  AND U7106 ( .A(n7404), .B(n7405), .Z(n7403) );
  XOR U7107 ( .A(n7402), .B(n6981), .Z(n7405) );
  XNOR U7108 ( .A(p_input[3244]), .B(n7406), .Z(n6981) );
  AND U7109 ( .A(n199), .B(n7407), .Z(n7406) );
  XOR U7110 ( .A(p_input[3260]), .B(p_input[3244]), .Z(n7407) );
  XNOR U7111 ( .A(n6978), .B(n7402), .Z(n7404) );
  XOR U7112 ( .A(n7408), .B(n7409), .Z(n6978) );
  AND U7113 ( .A(n196), .B(n7410), .Z(n7409) );
  XOR U7114 ( .A(p_input[3228]), .B(p_input[3212]), .Z(n7410) );
  XOR U7115 ( .A(n7411), .B(n7412), .Z(n7402) );
  AND U7116 ( .A(n7413), .B(n7414), .Z(n7412) );
  XOR U7117 ( .A(n7411), .B(n6993), .Z(n7414) );
  XNOR U7118 ( .A(p_input[3243]), .B(n7415), .Z(n6993) );
  AND U7119 ( .A(n199), .B(n7416), .Z(n7415) );
  XOR U7120 ( .A(p_input[3259]), .B(p_input[3243]), .Z(n7416) );
  XNOR U7121 ( .A(n6990), .B(n7411), .Z(n7413) );
  XOR U7122 ( .A(n7417), .B(n7418), .Z(n6990) );
  AND U7123 ( .A(n196), .B(n7419), .Z(n7418) );
  XOR U7124 ( .A(p_input[3227]), .B(p_input[3211]), .Z(n7419) );
  XOR U7125 ( .A(n7420), .B(n7421), .Z(n7411) );
  AND U7126 ( .A(n7422), .B(n7423), .Z(n7421) );
  XOR U7127 ( .A(n7420), .B(n7005), .Z(n7423) );
  XNOR U7128 ( .A(p_input[3242]), .B(n7424), .Z(n7005) );
  AND U7129 ( .A(n199), .B(n7425), .Z(n7424) );
  XOR U7130 ( .A(p_input[3258]), .B(p_input[3242]), .Z(n7425) );
  XNOR U7131 ( .A(n7002), .B(n7420), .Z(n7422) );
  XOR U7132 ( .A(n7426), .B(n7427), .Z(n7002) );
  AND U7133 ( .A(n196), .B(n7428), .Z(n7427) );
  XOR U7134 ( .A(p_input[3226]), .B(p_input[3210]), .Z(n7428) );
  XOR U7135 ( .A(n7429), .B(n7430), .Z(n7420) );
  AND U7136 ( .A(n7431), .B(n7432), .Z(n7430) );
  XOR U7137 ( .A(n7429), .B(n7017), .Z(n7432) );
  XNOR U7138 ( .A(p_input[3241]), .B(n7433), .Z(n7017) );
  AND U7139 ( .A(n199), .B(n7434), .Z(n7433) );
  XOR U7140 ( .A(p_input[3257]), .B(p_input[3241]), .Z(n7434) );
  XNOR U7141 ( .A(n7014), .B(n7429), .Z(n7431) );
  XOR U7142 ( .A(n7435), .B(n7436), .Z(n7014) );
  AND U7143 ( .A(n196), .B(n7437), .Z(n7436) );
  XOR U7144 ( .A(p_input[3225]), .B(p_input[3209]), .Z(n7437) );
  XOR U7145 ( .A(n7438), .B(n7439), .Z(n7429) );
  AND U7146 ( .A(n7440), .B(n7441), .Z(n7439) );
  XOR U7147 ( .A(n7438), .B(n7029), .Z(n7441) );
  XNOR U7148 ( .A(p_input[3240]), .B(n7442), .Z(n7029) );
  AND U7149 ( .A(n199), .B(n7443), .Z(n7442) );
  XOR U7150 ( .A(p_input[3256]), .B(p_input[3240]), .Z(n7443) );
  XNOR U7151 ( .A(n7026), .B(n7438), .Z(n7440) );
  XOR U7152 ( .A(n7444), .B(n7445), .Z(n7026) );
  AND U7153 ( .A(n196), .B(n7446), .Z(n7445) );
  XOR U7154 ( .A(p_input[3224]), .B(p_input[3208]), .Z(n7446) );
  XOR U7155 ( .A(n7447), .B(n7448), .Z(n7438) );
  AND U7156 ( .A(n7449), .B(n7450), .Z(n7448) );
  XOR U7157 ( .A(n7447), .B(n7041), .Z(n7450) );
  XNOR U7158 ( .A(p_input[3239]), .B(n7451), .Z(n7041) );
  AND U7159 ( .A(n199), .B(n7452), .Z(n7451) );
  XOR U7160 ( .A(p_input[3255]), .B(p_input[3239]), .Z(n7452) );
  XNOR U7161 ( .A(n7038), .B(n7447), .Z(n7449) );
  XOR U7162 ( .A(n7453), .B(n7454), .Z(n7038) );
  AND U7163 ( .A(n196), .B(n7455), .Z(n7454) );
  XOR U7164 ( .A(p_input[3223]), .B(p_input[3207]), .Z(n7455) );
  XOR U7165 ( .A(n7456), .B(n7457), .Z(n7447) );
  AND U7166 ( .A(n7458), .B(n7459), .Z(n7457) );
  XOR U7167 ( .A(n7456), .B(n7053), .Z(n7459) );
  XNOR U7168 ( .A(p_input[3238]), .B(n7460), .Z(n7053) );
  AND U7169 ( .A(n199), .B(n7461), .Z(n7460) );
  XOR U7170 ( .A(p_input[3254]), .B(p_input[3238]), .Z(n7461) );
  XNOR U7171 ( .A(n7050), .B(n7456), .Z(n7458) );
  XOR U7172 ( .A(n7462), .B(n7463), .Z(n7050) );
  AND U7173 ( .A(n196), .B(n7464), .Z(n7463) );
  XOR U7174 ( .A(p_input[3222]), .B(p_input[3206]), .Z(n7464) );
  XOR U7175 ( .A(n7465), .B(n7466), .Z(n7456) );
  AND U7176 ( .A(n7467), .B(n7468), .Z(n7466) );
  XOR U7177 ( .A(n7465), .B(n7065), .Z(n7468) );
  XNOR U7178 ( .A(p_input[3237]), .B(n7469), .Z(n7065) );
  AND U7179 ( .A(n199), .B(n7470), .Z(n7469) );
  XOR U7180 ( .A(p_input[3253]), .B(p_input[3237]), .Z(n7470) );
  XNOR U7181 ( .A(n7062), .B(n7465), .Z(n7467) );
  XOR U7182 ( .A(n7471), .B(n7472), .Z(n7062) );
  AND U7183 ( .A(n196), .B(n7473), .Z(n7472) );
  XOR U7184 ( .A(p_input[3221]), .B(p_input[3205]), .Z(n7473) );
  XOR U7185 ( .A(n7474), .B(n7475), .Z(n7465) );
  AND U7186 ( .A(n7476), .B(n7477), .Z(n7475) );
  XOR U7187 ( .A(n7474), .B(n7077), .Z(n7477) );
  XNOR U7188 ( .A(p_input[3236]), .B(n7478), .Z(n7077) );
  AND U7189 ( .A(n199), .B(n7479), .Z(n7478) );
  XOR U7190 ( .A(p_input[3252]), .B(p_input[3236]), .Z(n7479) );
  XNOR U7191 ( .A(n7074), .B(n7474), .Z(n7476) );
  XOR U7192 ( .A(n7480), .B(n7481), .Z(n7074) );
  AND U7193 ( .A(n196), .B(n7482), .Z(n7481) );
  XOR U7194 ( .A(p_input[3220]), .B(p_input[3204]), .Z(n7482) );
  XOR U7195 ( .A(n7483), .B(n7484), .Z(n7474) );
  AND U7196 ( .A(n7485), .B(n7486), .Z(n7484) );
  XOR U7197 ( .A(n7483), .B(n7089), .Z(n7486) );
  XNOR U7198 ( .A(p_input[3235]), .B(n7487), .Z(n7089) );
  AND U7199 ( .A(n199), .B(n7488), .Z(n7487) );
  XOR U7200 ( .A(p_input[3251]), .B(p_input[3235]), .Z(n7488) );
  XNOR U7201 ( .A(n7086), .B(n7483), .Z(n7485) );
  XOR U7202 ( .A(n7489), .B(n7490), .Z(n7086) );
  AND U7203 ( .A(n196), .B(n7491), .Z(n7490) );
  XOR U7204 ( .A(p_input[3219]), .B(p_input[3203]), .Z(n7491) );
  XOR U7205 ( .A(n7492), .B(n7493), .Z(n7483) );
  AND U7206 ( .A(n7494), .B(n7495), .Z(n7493) );
  XOR U7207 ( .A(n7492), .B(n7101), .Z(n7495) );
  XNOR U7208 ( .A(p_input[3234]), .B(n7496), .Z(n7101) );
  AND U7209 ( .A(n199), .B(n7497), .Z(n7496) );
  XOR U7210 ( .A(p_input[3250]), .B(p_input[3234]), .Z(n7497) );
  XNOR U7211 ( .A(n7098), .B(n7492), .Z(n7494) );
  XOR U7212 ( .A(n7498), .B(n7499), .Z(n7098) );
  AND U7213 ( .A(n196), .B(n7500), .Z(n7499) );
  XOR U7214 ( .A(p_input[3218]), .B(p_input[3202]), .Z(n7500) );
  XOR U7215 ( .A(n7501), .B(n7502), .Z(n7492) );
  AND U7216 ( .A(n7503), .B(n7504), .Z(n7502) );
  XNOR U7217 ( .A(n7505), .B(n7114), .Z(n7504) );
  XNOR U7218 ( .A(p_input[3233]), .B(n7506), .Z(n7114) );
  AND U7219 ( .A(n199), .B(n7507), .Z(n7506) );
  XNOR U7220 ( .A(p_input[3249]), .B(n7508), .Z(n7507) );
  IV U7221 ( .A(p_input[3233]), .Z(n7508) );
  XNOR U7222 ( .A(n7111), .B(n7501), .Z(n7503) );
  XNOR U7223 ( .A(p_input[3201]), .B(n7509), .Z(n7111) );
  AND U7224 ( .A(n196), .B(n7510), .Z(n7509) );
  XOR U7225 ( .A(p_input[3217]), .B(p_input[3201]), .Z(n7510) );
  IV U7226 ( .A(n7505), .Z(n7501) );
  AND U7227 ( .A(n7376), .B(n7379), .Z(n7505) );
  XOR U7228 ( .A(p_input[3232]), .B(n7511), .Z(n7379) );
  AND U7229 ( .A(n199), .B(n7512), .Z(n7511) );
  XOR U7230 ( .A(p_input[3248]), .B(p_input[3232]), .Z(n7512) );
  XOR U7231 ( .A(n7513), .B(n7514), .Z(n199) );
  AND U7232 ( .A(n7515), .B(n7516), .Z(n7514) );
  XNOR U7233 ( .A(p_input[3263]), .B(n7513), .Z(n7516) );
  XOR U7234 ( .A(n7513), .B(p_input[3247]), .Z(n7515) );
  XOR U7235 ( .A(n7517), .B(n7518), .Z(n7513) );
  AND U7236 ( .A(n7519), .B(n7520), .Z(n7518) );
  XNOR U7237 ( .A(p_input[3262]), .B(n7517), .Z(n7520) );
  XOR U7238 ( .A(n7517), .B(p_input[3246]), .Z(n7519) );
  XOR U7239 ( .A(n7521), .B(n7522), .Z(n7517) );
  AND U7240 ( .A(n7523), .B(n7524), .Z(n7522) );
  XNOR U7241 ( .A(p_input[3261]), .B(n7521), .Z(n7524) );
  XOR U7242 ( .A(n7521), .B(p_input[3245]), .Z(n7523) );
  XOR U7243 ( .A(n7525), .B(n7526), .Z(n7521) );
  AND U7244 ( .A(n7527), .B(n7528), .Z(n7526) );
  XNOR U7245 ( .A(p_input[3260]), .B(n7525), .Z(n7528) );
  XOR U7246 ( .A(n7525), .B(p_input[3244]), .Z(n7527) );
  XOR U7247 ( .A(n7529), .B(n7530), .Z(n7525) );
  AND U7248 ( .A(n7531), .B(n7532), .Z(n7530) );
  XNOR U7249 ( .A(p_input[3259]), .B(n7529), .Z(n7532) );
  XOR U7250 ( .A(n7529), .B(p_input[3243]), .Z(n7531) );
  XOR U7251 ( .A(n7533), .B(n7534), .Z(n7529) );
  AND U7252 ( .A(n7535), .B(n7536), .Z(n7534) );
  XNOR U7253 ( .A(p_input[3258]), .B(n7533), .Z(n7536) );
  XOR U7254 ( .A(n7533), .B(p_input[3242]), .Z(n7535) );
  XOR U7255 ( .A(n7537), .B(n7538), .Z(n7533) );
  AND U7256 ( .A(n7539), .B(n7540), .Z(n7538) );
  XNOR U7257 ( .A(p_input[3257]), .B(n7537), .Z(n7540) );
  XOR U7258 ( .A(n7537), .B(p_input[3241]), .Z(n7539) );
  XOR U7259 ( .A(n7541), .B(n7542), .Z(n7537) );
  AND U7260 ( .A(n7543), .B(n7544), .Z(n7542) );
  XNOR U7261 ( .A(p_input[3256]), .B(n7541), .Z(n7544) );
  XOR U7262 ( .A(n7541), .B(p_input[3240]), .Z(n7543) );
  XOR U7263 ( .A(n7545), .B(n7546), .Z(n7541) );
  AND U7264 ( .A(n7547), .B(n7548), .Z(n7546) );
  XNOR U7265 ( .A(p_input[3255]), .B(n7545), .Z(n7548) );
  XOR U7266 ( .A(n7545), .B(p_input[3239]), .Z(n7547) );
  XOR U7267 ( .A(n7549), .B(n7550), .Z(n7545) );
  AND U7268 ( .A(n7551), .B(n7552), .Z(n7550) );
  XNOR U7269 ( .A(p_input[3254]), .B(n7549), .Z(n7552) );
  XOR U7270 ( .A(n7549), .B(p_input[3238]), .Z(n7551) );
  XOR U7271 ( .A(n7553), .B(n7554), .Z(n7549) );
  AND U7272 ( .A(n7555), .B(n7556), .Z(n7554) );
  XNOR U7273 ( .A(p_input[3253]), .B(n7553), .Z(n7556) );
  XOR U7274 ( .A(n7553), .B(p_input[3237]), .Z(n7555) );
  XOR U7275 ( .A(n7557), .B(n7558), .Z(n7553) );
  AND U7276 ( .A(n7559), .B(n7560), .Z(n7558) );
  XNOR U7277 ( .A(p_input[3252]), .B(n7557), .Z(n7560) );
  XOR U7278 ( .A(n7557), .B(p_input[3236]), .Z(n7559) );
  XOR U7279 ( .A(n7561), .B(n7562), .Z(n7557) );
  AND U7280 ( .A(n7563), .B(n7564), .Z(n7562) );
  XNOR U7281 ( .A(p_input[3251]), .B(n7561), .Z(n7564) );
  XOR U7282 ( .A(n7561), .B(p_input[3235]), .Z(n7563) );
  XOR U7283 ( .A(n7565), .B(n7566), .Z(n7561) );
  AND U7284 ( .A(n7567), .B(n7568), .Z(n7566) );
  XNOR U7285 ( .A(p_input[3250]), .B(n7565), .Z(n7568) );
  XOR U7286 ( .A(n7565), .B(p_input[3234]), .Z(n7567) );
  XNOR U7287 ( .A(n7569), .B(n7570), .Z(n7565) );
  AND U7288 ( .A(n7571), .B(n7572), .Z(n7570) );
  XOR U7289 ( .A(p_input[3249]), .B(n7569), .Z(n7572) );
  XNOR U7290 ( .A(p_input[3233]), .B(n7569), .Z(n7571) );
  AND U7291 ( .A(p_input[3248]), .B(n7573), .Z(n7569) );
  IV U7292 ( .A(p_input[3232]), .Z(n7573) );
  XNOR U7293 ( .A(p_input[3200]), .B(n7574), .Z(n7376) );
  AND U7294 ( .A(n196), .B(n7575), .Z(n7574) );
  XOR U7295 ( .A(p_input[3216]), .B(p_input[3200]), .Z(n7575) );
  XOR U7296 ( .A(n7576), .B(n7577), .Z(n196) );
  AND U7297 ( .A(n7578), .B(n7579), .Z(n7577) );
  XNOR U7298 ( .A(p_input[3231]), .B(n7576), .Z(n7579) );
  XOR U7299 ( .A(n7576), .B(p_input[3215]), .Z(n7578) );
  XOR U7300 ( .A(n7580), .B(n7581), .Z(n7576) );
  AND U7301 ( .A(n7582), .B(n7583), .Z(n7581) );
  XNOR U7302 ( .A(p_input[3230]), .B(n7580), .Z(n7583) );
  XNOR U7303 ( .A(n7580), .B(n7390), .Z(n7582) );
  IV U7304 ( .A(p_input[3214]), .Z(n7390) );
  XOR U7305 ( .A(n7584), .B(n7585), .Z(n7580) );
  AND U7306 ( .A(n7586), .B(n7587), .Z(n7585) );
  XNOR U7307 ( .A(p_input[3229]), .B(n7584), .Z(n7587) );
  XNOR U7308 ( .A(n7584), .B(n7399), .Z(n7586) );
  IV U7309 ( .A(p_input[3213]), .Z(n7399) );
  XOR U7310 ( .A(n7588), .B(n7589), .Z(n7584) );
  AND U7311 ( .A(n7590), .B(n7591), .Z(n7589) );
  XNOR U7312 ( .A(p_input[3228]), .B(n7588), .Z(n7591) );
  XNOR U7313 ( .A(n7588), .B(n7408), .Z(n7590) );
  IV U7314 ( .A(p_input[3212]), .Z(n7408) );
  XOR U7315 ( .A(n7592), .B(n7593), .Z(n7588) );
  AND U7316 ( .A(n7594), .B(n7595), .Z(n7593) );
  XNOR U7317 ( .A(p_input[3227]), .B(n7592), .Z(n7595) );
  XNOR U7318 ( .A(n7592), .B(n7417), .Z(n7594) );
  IV U7319 ( .A(p_input[3211]), .Z(n7417) );
  XOR U7320 ( .A(n7596), .B(n7597), .Z(n7592) );
  AND U7321 ( .A(n7598), .B(n7599), .Z(n7597) );
  XNOR U7322 ( .A(p_input[3226]), .B(n7596), .Z(n7599) );
  XNOR U7323 ( .A(n7596), .B(n7426), .Z(n7598) );
  IV U7324 ( .A(p_input[3210]), .Z(n7426) );
  XOR U7325 ( .A(n7600), .B(n7601), .Z(n7596) );
  AND U7326 ( .A(n7602), .B(n7603), .Z(n7601) );
  XNOR U7327 ( .A(p_input[3225]), .B(n7600), .Z(n7603) );
  XNOR U7328 ( .A(n7600), .B(n7435), .Z(n7602) );
  IV U7329 ( .A(p_input[3209]), .Z(n7435) );
  XOR U7330 ( .A(n7604), .B(n7605), .Z(n7600) );
  AND U7331 ( .A(n7606), .B(n7607), .Z(n7605) );
  XNOR U7332 ( .A(p_input[3224]), .B(n7604), .Z(n7607) );
  XNOR U7333 ( .A(n7604), .B(n7444), .Z(n7606) );
  IV U7334 ( .A(p_input[3208]), .Z(n7444) );
  XOR U7335 ( .A(n7608), .B(n7609), .Z(n7604) );
  AND U7336 ( .A(n7610), .B(n7611), .Z(n7609) );
  XNOR U7337 ( .A(p_input[3223]), .B(n7608), .Z(n7611) );
  XNOR U7338 ( .A(n7608), .B(n7453), .Z(n7610) );
  IV U7339 ( .A(p_input[3207]), .Z(n7453) );
  XOR U7340 ( .A(n7612), .B(n7613), .Z(n7608) );
  AND U7341 ( .A(n7614), .B(n7615), .Z(n7613) );
  XNOR U7342 ( .A(p_input[3222]), .B(n7612), .Z(n7615) );
  XNOR U7343 ( .A(n7612), .B(n7462), .Z(n7614) );
  IV U7344 ( .A(p_input[3206]), .Z(n7462) );
  XOR U7345 ( .A(n7616), .B(n7617), .Z(n7612) );
  AND U7346 ( .A(n7618), .B(n7619), .Z(n7617) );
  XNOR U7347 ( .A(p_input[3221]), .B(n7616), .Z(n7619) );
  XNOR U7348 ( .A(n7616), .B(n7471), .Z(n7618) );
  IV U7349 ( .A(p_input[3205]), .Z(n7471) );
  XOR U7350 ( .A(n7620), .B(n7621), .Z(n7616) );
  AND U7351 ( .A(n7622), .B(n7623), .Z(n7621) );
  XNOR U7352 ( .A(p_input[3220]), .B(n7620), .Z(n7623) );
  XNOR U7353 ( .A(n7620), .B(n7480), .Z(n7622) );
  IV U7354 ( .A(p_input[3204]), .Z(n7480) );
  XOR U7355 ( .A(n7624), .B(n7625), .Z(n7620) );
  AND U7356 ( .A(n7626), .B(n7627), .Z(n7625) );
  XNOR U7357 ( .A(p_input[3219]), .B(n7624), .Z(n7627) );
  XNOR U7358 ( .A(n7624), .B(n7489), .Z(n7626) );
  IV U7359 ( .A(p_input[3203]), .Z(n7489) );
  XOR U7360 ( .A(n7628), .B(n7629), .Z(n7624) );
  AND U7361 ( .A(n7630), .B(n7631), .Z(n7629) );
  XNOR U7362 ( .A(p_input[3218]), .B(n7628), .Z(n7631) );
  XNOR U7363 ( .A(n7628), .B(n7498), .Z(n7630) );
  IV U7364 ( .A(p_input[3202]), .Z(n7498) );
  XNOR U7365 ( .A(n7632), .B(n7633), .Z(n7628) );
  AND U7366 ( .A(n7634), .B(n7635), .Z(n7633) );
  XOR U7367 ( .A(p_input[3217]), .B(n7632), .Z(n7635) );
  XNOR U7368 ( .A(p_input[3201]), .B(n7632), .Z(n7634) );
  AND U7369 ( .A(p_input[3216]), .B(n7636), .Z(n7632) );
  IV U7370 ( .A(p_input[3200]), .Z(n7636) );
  XOR U7371 ( .A(n7637), .B(n7638), .Z(n6752) );
  AND U7372 ( .A(n748), .B(n7639), .Z(n7638) );
  XNOR U7373 ( .A(n7640), .B(n7637), .Z(n7639) );
  XOR U7374 ( .A(n7641), .B(n7642), .Z(n748) );
  AND U7375 ( .A(n7643), .B(n7644), .Z(n7642) );
  XNOR U7376 ( .A(n6764), .B(n7641), .Z(n7644) );
  AND U7377 ( .A(n7645), .B(n7646), .Z(n6764) );
  XOR U7378 ( .A(n7641), .B(n6763), .Z(n7643) );
  AND U7379 ( .A(n7647), .B(n7648), .Z(n6763) );
  XOR U7380 ( .A(n7649), .B(n7650), .Z(n7641) );
  AND U7381 ( .A(n7651), .B(n7652), .Z(n7650) );
  XOR U7382 ( .A(n7649), .B(n6776), .Z(n7652) );
  XOR U7383 ( .A(n7653), .B(n7654), .Z(n6776) );
  AND U7384 ( .A(n403), .B(n7655), .Z(n7654) );
  XOR U7385 ( .A(n7656), .B(n7653), .Z(n7655) );
  XNOR U7386 ( .A(n6773), .B(n7649), .Z(n7651) );
  XOR U7387 ( .A(n7657), .B(n7658), .Z(n6773) );
  AND U7388 ( .A(n400), .B(n7659), .Z(n7658) );
  XOR U7389 ( .A(n7660), .B(n7657), .Z(n7659) );
  XOR U7390 ( .A(n7661), .B(n7662), .Z(n7649) );
  AND U7391 ( .A(n7663), .B(n7664), .Z(n7662) );
  XOR U7392 ( .A(n7661), .B(n6788), .Z(n7664) );
  XOR U7393 ( .A(n7665), .B(n7666), .Z(n6788) );
  AND U7394 ( .A(n403), .B(n7667), .Z(n7666) );
  XOR U7395 ( .A(n7668), .B(n7665), .Z(n7667) );
  XNOR U7396 ( .A(n6785), .B(n7661), .Z(n7663) );
  XOR U7397 ( .A(n7669), .B(n7670), .Z(n6785) );
  AND U7398 ( .A(n400), .B(n7671), .Z(n7670) );
  XOR U7399 ( .A(n7672), .B(n7669), .Z(n7671) );
  XOR U7400 ( .A(n7673), .B(n7674), .Z(n7661) );
  AND U7401 ( .A(n7675), .B(n7676), .Z(n7674) );
  XOR U7402 ( .A(n7673), .B(n6800), .Z(n7676) );
  XOR U7403 ( .A(n7677), .B(n7678), .Z(n6800) );
  AND U7404 ( .A(n403), .B(n7679), .Z(n7678) );
  XOR U7405 ( .A(n7680), .B(n7677), .Z(n7679) );
  XNOR U7406 ( .A(n6797), .B(n7673), .Z(n7675) );
  XOR U7407 ( .A(n7681), .B(n7682), .Z(n6797) );
  AND U7408 ( .A(n400), .B(n7683), .Z(n7682) );
  XOR U7409 ( .A(n7684), .B(n7681), .Z(n7683) );
  XOR U7410 ( .A(n7685), .B(n7686), .Z(n7673) );
  AND U7411 ( .A(n7687), .B(n7688), .Z(n7686) );
  XOR U7412 ( .A(n7685), .B(n6812), .Z(n7688) );
  XOR U7413 ( .A(n7689), .B(n7690), .Z(n6812) );
  AND U7414 ( .A(n403), .B(n7691), .Z(n7690) );
  XOR U7415 ( .A(n7692), .B(n7689), .Z(n7691) );
  XNOR U7416 ( .A(n6809), .B(n7685), .Z(n7687) );
  XOR U7417 ( .A(n7693), .B(n7694), .Z(n6809) );
  AND U7418 ( .A(n400), .B(n7695), .Z(n7694) );
  XOR U7419 ( .A(n7696), .B(n7693), .Z(n7695) );
  XOR U7420 ( .A(n7697), .B(n7698), .Z(n7685) );
  AND U7421 ( .A(n7699), .B(n7700), .Z(n7698) );
  XOR U7422 ( .A(n7697), .B(n6824), .Z(n7700) );
  XOR U7423 ( .A(n7701), .B(n7702), .Z(n6824) );
  AND U7424 ( .A(n403), .B(n7703), .Z(n7702) );
  XOR U7425 ( .A(n7704), .B(n7701), .Z(n7703) );
  XNOR U7426 ( .A(n6821), .B(n7697), .Z(n7699) );
  XOR U7427 ( .A(n7705), .B(n7706), .Z(n6821) );
  AND U7428 ( .A(n400), .B(n7707), .Z(n7706) );
  XOR U7429 ( .A(n7708), .B(n7705), .Z(n7707) );
  XOR U7430 ( .A(n7709), .B(n7710), .Z(n7697) );
  AND U7431 ( .A(n7711), .B(n7712), .Z(n7710) );
  XOR U7432 ( .A(n7709), .B(n6836), .Z(n7712) );
  XOR U7433 ( .A(n7713), .B(n7714), .Z(n6836) );
  AND U7434 ( .A(n403), .B(n7715), .Z(n7714) );
  XOR U7435 ( .A(n7716), .B(n7713), .Z(n7715) );
  XNOR U7436 ( .A(n6833), .B(n7709), .Z(n7711) );
  XOR U7437 ( .A(n7717), .B(n7718), .Z(n6833) );
  AND U7438 ( .A(n400), .B(n7719), .Z(n7718) );
  XOR U7439 ( .A(n7720), .B(n7717), .Z(n7719) );
  XOR U7440 ( .A(n7721), .B(n7722), .Z(n7709) );
  AND U7441 ( .A(n7723), .B(n7724), .Z(n7722) );
  XOR U7442 ( .A(n7721), .B(n6848), .Z(n7724) );
  XOR U7443 ( .A(n7725), .B(n7726), .Z(n6848) );
  AND U7444 ( .A(n403), .B(n7727), .Z(n7726) );
  XOR U7445 ( .A(n7728), .B(n7725), .Z(n7727) );
  XNOR U7446 ( .A(n6845), .B(n7721), .Z(n7723) );
  XOR U7447 ( .A(n7729), .B(n7730), .Z(n6845) );
  AND U7448 ( .A(n400), .B(n7731), .Z(n7730) );
  XOR U7449 ( .A(n7732), .B(n7729), .Z(n7731) );
  XOR U7450 ( .A(n7733), .B(n7734), .Z(n7721) );
  AND U7451 ( .A(n7735), .B(n7736), .Z(n7734) );
  XOR U7452 ( .A(n7733), .B(n6860), .Z(n7736) );
  XOR U7453 ( .A(n7737), .B(n7738), .Z(n6860) );
  AND U7454 ( .A(n403), .B(n7739), .Z(n7738) );
  XOR U7455 ( .A(n7740), .B(n7737), .Z(n7739) );
  XNOR U7456 ( .A(n6857), .B(n7733), .Z(n7735) );
  XOR U7457 ( .A(n7741), .B(n7742), .Z(n6857) );
  AND U7458 ( .A(n400), .B(n7743), .Z(n7742) );
  XOR U7459 ( .A(n7744), .B(n7741), .Z(n7743) );
  XOR U7460 ( .A(n7745), .B(n7746), .Z(n7733) );
  AND U7461 ( .A(n7747), .B(n7748), .Z(n7746) );
  XOR U7462 ( .A(n7745), .B(n6872), .Z(n7748) );
  XOR U7463 ( .A(n7749), .B(n7750), .Z(n6872) );
  AND U7464 ( .A(n403), .B(n7751), .Z(n7750) );
  XOR U7465 ( .A(n7752), .B(n7749), .Z(n7751) );
  XNOR U7466 ( .A(n6869), .B(n7745), .Z(n7747) );
  XOR U7467 ( .A(n7753), .B(n7754), .Z(n6869) );
  AND U7468 ( .A(n400), .B(n7755), .Z(n7754) );
  XOR U7469 ( .A(n7756), .B(n7753), .Z(n7755) );
  XOR U7470 ( .A(n7757), .B(n7758), .Z(n7745) );
  AND U7471 ( .A(n7759), .B(n7760), .Z(n7758) );
  XOR U7472 ( .A(n7757), .B(n6884), .Z(n7760) );
  XOR U7473 ( .A(n7761), .B(n7762), .Z(n6884) );
  AND U7474 ( .A(n403), .B(n7763), .Z(n7762) );
  XOR U7475 ( .A(n7764), .B(n7761), .Z(n7763) );
  XNOR U7476 ( .A(n6881), .B(n7757), .Z(n7759) );
  XOR U7477 ( .A(n7765), .B(n7766), .Z(n6881) );
  AND U7478 ( .A(n400), .B(n7767), .Z(n7766) );
  XOR U7479 ( .A(n7768), .B(n7765), .Z(n7767) );
  XOR U7480 ( .A(n7769), .B(n7770), .Z(n7757) );
  AND U7481 ( .A(n7771), .B(n7772), .Z(n7770) );
  XOR U7482 ( .A(n7769), .B(n6896), .Z(n7772) );
  XOR U7483 ( .A(n7773), .B(n7774), .Z(n6896) );
  AND U7484 ( .A(n403), .B(n7775), .Z(n7774) );
  XOR U7485 ( .A(n7776), .B(n7773), .Z(n7775) );
  XNOR U7486 ( .A(n6893), .B(n7769), .Z(n7771) );
  XOR U7487 ( .A(n7777), .B(n7778), .Z(n6893) );
  AND U7488 ( .A(n400), .B(n7779), .Z(n7778) );
  XOR U7489 ( .A(n7780), .B(n7777), .Z(n7779) );
  XOR U7490 ( .A(n7781), .B(n7782), .Z(n7769) );
  AND U7491 ( .A(n7783), .B(n7784), .Z(n7782) );
  XOR U7492 ( .A(n7781), .B(n6908), .Z(n7784) );
  XOR U7493 ( .A(n7785), .B(n7786), .Z(n6908) );
  AND U7494 ( .A(n403), .B(n7787), .Z(n7786) );
  XOR U7495 ( .A(n7788), .B(n7785), .Z(n7787) );
  XNOR U7496 ( .A(n6905), .B(n7781), .Z(n7783) );
  XOR U7497 ( .A(n7789), .B(n7790), .Z(n6905) );
  AND U7498 ( .A(n400), .B(n7791), .Z(n7790) );
  XOR U7499 ( .A(n7792), .B(n7789), .Z(n7791) );
  XOR U7500 ( .A(n7793), .B(n7794), .Z(n7781) );
  AND U7501 ( .A(n7795), .B(n7796), .Z(n7794) );
  XOR U7502 ( .A(n7793), .B(n6920), .Z(n7796) );
  XOR U7503 ( .A(n7797), .B(n7798), .Z(n6920) );
  AND U7504 ( .A(n403), .B(n7799), .Z(n7798) );
  XOR U7505 ( .A(n7800), .B(n7797), .Z(n7799) );
  XNOR U7506 ( .A(n6917), .B(n7793), .Z(n7795) );
  XOR U7507 ( .A(n7801), .B(n7802), .Z(n6917) );
  AND U7508 ( .A(n400), .B(n7803), .Z(n7802) );
  XOR U7509 ( .A(n7804), .B(n7801), .Z(n7803) );
  XOR U7510 ( .A(n7805), .B(n7806), .Z(n7793) );
  AND U7511 ( .A(n7807), .B(n7808), .Z(n7806) );
  XNOR U7512 ( .A(n7809), .B(n6933), .Z(n7808) );
  XOR U7513 ( .A(n7810), .B(n7811), .Z(n6933) );
  AND U7514 ( .A(n403), .B(n7812), .Z(n7811) );
  XOR U7515 ( .A(n7810), .B(n7813), .Z(n7812) );
  XNOR U7516 ( .A(n6930), .B(n7805), .Z(n7807) );
  XOR U7517 ( .A(n7814), .B(n7815), .Z(n6930) );
  AND U7518 ( .A(n400), .B(n7816), .Z(n7815) );
  XOR U7519 ( .A(n7814), .B(n7817), .Z(n7816) );
  IV U7520 ( .A(n7809), .Z(n7805) );
  AND U7521 ( .A(n7637), .B(n7640), .Z(n7809) );
  XNOR U7522 ( .A(n7818), .B(n7819), .Z(n7640) );
  AND U7523 ( .A(n403), .B(n7820), .Z(n7819) );
  XNOR U7524 ( .A(n7821), .B(n7818), .Z(n7820) );
  XOR U7525 ( .A(n7822), .B(n7823), .Z(n403) );
  AND U7526 ( .A(n7824), .B(n7825), .Z(n7823) );
  XNOR U7527 ( .A(n7645), .B(n7822), .Z(n7825) );
  AND U7528 ( .A(p_input[3199]), .B(p_input[3183]), .Z(n7645) );
  XOR U7529 ( .A(n7822), .B(n7646), .Z(n7824) );
  AND U7530 ( .A(p_input[3167]), .B(p_input[3151]), .Z(n7646) );
  XOR U7531 ( .A(n7826), .B(n7827), .Z(n7822) );
  AND U7532 ( .A(n7828), .B(n7829), .Z(n7827) );
  XOR U7533 ( .A(n7826), .B(n7656), .Z(n7829) );
  XNOR U7534 ( .A(p_input[3182]), .B(n7830), .Z(n7656) );
  AND U7535 ( .A(n207), .B(n7831), .Z(n7830) );
  XOR U7536 ( .A(p_input[3198]), .B(p_input[3182]), .Z(n7831) );
  XNOR U7537 ( .A(n7653), .B(n7826), .Z(n7828) );
  XOR U7538 ( .A(n7832), .B(n7833), .Z(n7653) );
  AND U7539 ( .A(n205), .B(n7834), .Z(n7833) );
  XOR U7540 ( .A(p_input[3166]), .B(p_input[3150]), .Z(n7834) );
  XOR U7541 ( .A(n7835), .B(n7836), .Z(n7826) );
  AND U7542 ( .A(n7837), .B(n7838), .Z(n7836) );
  XOR U7543 ( .A(n7835), .B(n7668), .Z(n7838) );
  XNOR U7544 ( .A(p_input[3181]), .B(n7839), .Z(n7668) );
  AND U7545 ( .A(n207), .B(n7840), .Z(n7839) );
  XOR U7546 ( .A(p_input[3197]), .B(p_input[3181]), .Z(n7840) );
  XNOR U7547 ( .A(n7665), .B(n7835), .Z(n7837) );
  XOR U7548 ( .A(n7841), .B(n7842), .Z(n7665) );
  AND U7549 ( .A(n205), .B(n7843), .Z(n7842) );
  XOR U7550 ( .A(p_input[3165]), .B(p_input[3149]), .Z(n7843) );
  XOR U7551 ( .A(n7844), .B(n7845), .Z(n7835) );
  AND U7552 ( .A(n7846), .B(n7847), .Z(n7845) );
  XOR U7553 ( .A(n7844), .B(n7680), .Z(n7847) );
  XNOR U7554 ( .A(p_input[3180]), .B(n7848), .Z(n7680) );
  AND U7555 ( .A(n207), .B(n7849), .Z(n7848) );
  XOR U7556 ( .A(p_input[3196]), .B(p_input[3180]), .Z(n7849) );
  XNOR U7557 ( .A(n7677), .B(n7844), .Z(n7846) );
  XOR U7558 ( .A(n7850), .B(n7851), .Z(n7677) );
  AND U7559 ( .A(n205), .B(n7852), .Z(n7851) );
  XOR U7560 ( .A(p_input[3164]), .B(p_input[3148]), .Z(n7852) );
  XOR U7561 ( .A(n7853), .B(n7854), .Z(n7844) );
  AND U7562 ( .A(n7855), .B(n7856), .Z(n7854) );
  XOR U7563 ( .A(n7853), .B(n7692), .Z(n7856) );
  XNOR U7564 ( .A(p_input[3179]), .B(n7857), .Z(n7692) );
  AND U7565 ( .A(n207), .B(n7858), .Z(n7857) );
  XOR U7566 ( .A(p_input[3195]), .B(p_input[3179]), .Z(n7858) );
  XNOR U7567 ( .A(n7689), .B(n7853), .Z(n7855) );
  XOR U7568 ( .A(n7859), .B(n7860), .Z(n7689) );
  AND U7569 ( .A(n205), .B(n7861), .Z(n7860) );
  XOR U7570 ( .A(p_input[3163]), .B(p_input[3147]), .Z(n7861) );
  XOR U7571 ( .A(n7862), .B(n7863), .Z(n7853) );
  AND U7572 ( .A(n7864), .B(n7865), .Z(n7863) );
  XOR U7573 ( .A(n7862), .B(n7704), .Z(n7865) );
  XNOR U7574 ( .A(p_input[3178]), .B(n7866), .Z(n7704) );
  AND U7575 ( .A(n207), .B(n7867), .Z(n7866) );
  XOR U7576 ( .A(p_input[3194]), .B(p_input[3178]), .Z(n7867) );
  XNOR U7577 ( .A(n7701), .B(n7862), .Z(n7864) );
  XOR U7578 ( .A(n7868), .B(n7869), .Z(n7701) );
  AND U7579 ( .A(n205), .B(n7870), .Z(n7869) );
  XOR U7580 ( .A(p_input[3162]), .B(p_input[3146]), .Z(n7870) );
  XOR U7581 ( .A(n7871), .B(n7872), .Z(n7862) );
  AND U7582 ( .A(n7873), .B(n7874), .Z(n7872) );
  XOR U7583 ( .A(n7871), .B(n7716), .Z(n7874) );
  XNOR U7584 ( .A(p_input[3177]), .B(n7875), .Z(n7716) );
  AND U7585 ( .A(n207), .B(n7876), .Z(n7875) );
  XOR U7586 ( .A(p_input[3193]), .B(p_input[3177]), .Z(n7876) );
  XNOR U7587 ( .A(n7713), .B(n7871), .Z(n7873) );
  XOR U7588 ( .A(n7877), .B(n7878), .Z(n7713) );
  AND U7589 ( .A(n205), .B(n7879), .Z(n7878) );
  XOR U7590 ( .A(p_input[3161]), .B(p_input[3145]), .Z(n7879) );
  XOR U7591 ( .A(n7880), .B(n7881), .Z(n7871) );
  AND U7592 ( .A(n7882), .B(n7883), .Z(n7881) );
  XOR U7593 ( .A(n7880), .B(n7728), .Z(n7883) );
  XNOR U7594 ( .A(p_input[3176]), .B(n7884), .Z(n7728) );
  AND U7595 ( .A(n207), .B(n7885), .Z(n7884) );
  XOR U7596 ( .A(p_input[3192]), .B(p_input[3176]), .Z(n7885) );
  XNOR U7597 ( .A(n7725), .B(n7880), .Z(n7882) );
  XOR U7598 ( .A(n7886), .B(n7887), .Z(n7725) );
  AND U7599 ( .A(n205), .B(n7888), .Z(n7887) );
  XOR U7600 ( .A(p_input[3160]), .B(p_input[3144]), .Z(n7888) );
  XOR U7601 ( .A(n7889), .B(n7890), .Z(n7880) );
  AND U7602 ( .A(n7891), .B(n7892), .Z(n7890) );
  XOR U7603 ( .A(n7889), .B(n7740), .Z(n7892) );
  XNOR U7604 ( .A(p_input[3175]), .B(n7893), .Z(n7740) );
  AND U7605 ( .A(n207), .B(n7894), .Z(n7893) );
  XOR U7606 ( .A(p_input[3191]), .B(p_input[3175]), .Z(n7894) );
  XNOR U7607 ( .A(n7737), .B(n7889), .Z(n7891) );
  XOR U7608 ( .A(n7895), .B(n7896), .Z(n7737) );
  AND U7609 ( .A(n205), .B(n7897), .Z(n7896) );
  XOR U7610 ( .A(p_input[3159]), .B(p_input[3143]), .Z(n7897) );
  XOR U7611 ( .A(n7898), .B(n7899), .Z(n7889) );
  AND U7612 ( .A(n7900), .B(n7901), .Z(n7899) );
  XOR U7613 ( .A(n7898), .B(n7752), .Z(n7901) );
  XNOR U7614 ( .A(p_input[3174]), .B(n7902), .Z(n7752) );
  AND U7615 ( .A(n207), .B(n7903), .Z(n7902) );
  XOR U7616 ( .A(p_input[3190]), .B(p_input[3174]), .Z(n7903) );
  XNOR U7617 ( .A(n7749), .B(n7898), .Z(n7900) );
  XOR U7618 ( .A(n7904), .B(n7905), .Z(n7749) );
  AND U7619 ( .A(n205), .B(n7906), .Z(n7905) );
  XOR U7620 ( .A(p_input[3158]), .B(p_input[3142]), .Z(n7906) );
  XOR U7621 ( .A(n7907), .B(n7908), .Z(n7898) );
  AND U7622 ( .A(n7909), .B(n7910), .Z(n7908) );
  XOR U7623 ( .A(n7907), .B(n7764), .Z(n7910) );
  XNOR U7624 ( .A(p_input[3173]), .B(n7911), .Z(n7764) );
  AND U7625 ( .A(n207), .B(n7912), .Z(n7911) );
  XOR U7626 ( .A(p_input[3189]), .B(p_input[3173]), .Z(n7912) );
  XNOR U7627 ( .A(n7761), .B(n7907), .Z(n7909) );
  XOR U7628 ( .A(n7913), .B(n7914), .Z(n7761) );
  AND U7629 ( .A(n205), .B(n7915), .Z(n7914) );
  XOR U7630 ( .A(p_input[3157]), .B(p_input[3141]), .Z(n7915) );
  XOR U7631 ( .A(n7916), .B(n7917), .Z(n7907) );
  AND U7632 ( .A(n7918), .B(n7919), .Z(n7917) );
  XOR U7633 ( .A(n7916), .B(n7776), .Z(n7919) );
  XNOR U7634 ( .A(p_input[3172]), .B(n7920), .Z(n7776) );
  AND U7635 ( .A(n207), .B(n7921), .Z(n7920) );
  XOR U7636 ( .A(p_input[3188]), .B(p_input[3172]), .Z(n7921) );
  XNOR U7637 ( .A(n7773), .B(n7916), .Z(n7918) );
  XOR U7638 ( .A(n7922), .B(n7923), .Z(n7773) );
  AND U7639 ( .A(n205), .B(n7924), .Z(n7923) );
  XOR U7640 ( .A(p_input[3156]), .B(p_input[3140]), .Z(n7924) );
  XOR U7641 ( .A(n7925), .B(n7926), .Z(n7916) );
  AND U7642 ( .A(n7927), .B(n7928), .Z(n7926) );
  XOR U7643 ( .A(n7925), .B(n7788), .Z(n7928) );
  XNOR U7644 ( .A(p_input[3171]), .B(n7929), .Z(n7788) );
  AND U7645 ( .A(n207), .B(n7930), .Z(n7929) );
  XOR U7646 ( .A(p_input[3187]), .B(p_input[3171]), .Z(n7930) );
  XNOR U7647 ( .A(n7785), .B(n7925), .Z(n7927) );
  XOR U7648 ( .A(n7931), .B(n7932), .Z(n7785) );
  AND U7649 ( .A(n205), .B(n7933), .Z(n7932) );
  XOR U7650 ( .A(p_input[3155]), .B(p_input[3139]), .Z(n7933) );
  XOR U7651 ( .A(n7934), .B(n7935), .Z(n7925) );
  AND U7652 ( .A(n7936), .B(n7937), .Z(n7935) );
  XOR U7653 ( .A(n7934), .B(n7800), .Z(n7937) );
  XNOR U7654 ( .A(p_input[3170]), .B(n7938), .Z(n7800) );
  AND U7655 ( .A(n207), .B(n7939), .Z(n7938) );
  XOR U7656 ( .A(p_input[3186]), .B(p_input[3170]), .Z(n7939) );
  XNOR U7657 ( .A(n7797), .B(n7934), .Z(n7936) );
  XOR U7658 ( .A(n7940), .B(n7941), .Z(n7797) );
  AND U7659 ( .A(n205), .B(n7942), .Z(n7941) );
  XOR U7660 ( .A(p_input[3154]), .B(p_input[3138]), .Z(n7942) );
  XOR U7661 ( .A(n7943), .B(n7944), .Z(n7934) );
  AND U7662 ( .A(n7945), .B(n7946), .Z(n7944) );
  XNOR U7663 ( .A(n7947), .B(n7813), .Z(n7946) );
  XNOR U7664 ( .A(p_input[3169]), .B(n7948), .Z(n7813) );
  AND U7665 ( .A(n207), .B(n7949), .Z(n7948) );
  XNOR U7666 ( .A(p_input[3185]), .B(n7950), .Z(n7949) );
  IV U7667 ( .A(p_input[3169]), .Z(n7950) );
  XNOR U7668 ( .A(n7810), .B(n7943), .Z(n7945) );
  XNOR U7669 ( .A(p_input[3137]), .B(n7951), .Z(n7810) );
  AND U7670 ( .A(n205), .B(n7952), .Z(n7951) );
  XOR U7671 ( .A(p_input[3153]), .B(p_input[3137]), .Z(n7952) );
  IV U7672 ( .A(n7947), .Z(n7943) );
  AND U7673 ( .A(n7818), .B(n7821), .Z(n7947) );
  XOR U7674 ( .A(p_input[3168]), .B(n7953), .Z(n7821) );
  AND U7675 ( .A(n207), .B(n7954), .Z(n7953) );
  XOR U7676 ( .A(p_input[3184]), .B(p_input[3168]), .Z(n7954) );
  XOR U7677 ( .A(n7955), .B(n7956), .Z(n207) );
  AND U7678 ( .A(n7957), .B(n7958), .Z(n7956) );
  XNOR U7679 ( .A(p_input[3199]), .B(n7955), .Z(n7958) );
  XOR U7680 ( .A(n7955), .B(p_input[3183]), .Z(n7957) );
  XOR U7681 ( .A(n7959), .B(n7960), .Z(n7955) );
  AND U7682 ( .A(n7961), .B(n7962), .Z(n7960) );
  XNOR U7683 ( .A(p_input[3198]), .B(n7959), .Z(n7962) );
  XOR U7684 ( .A(n7959), .B(p_input[3182]), .Z(n7961) );
  XOR U7685 ( .A(n7963), .B(n7964), .Z(n7959) );
  AND U7686 ( .A(n7965), .B(n7966), .Z(n7964) );
  XNOR U7687 ( .A(p_input[3197]), .B(n7963), .Z(n7966) );
  XOR U7688 ( .A(n7963), .B(p_input[3181]), .Z(n7965) );
  XOR U7689 ( .A(n7967), .B(n7968), .Z(n7963) );
  AND U7690 ( .A(n7969), .B(n7970), .Z(n7968) );
  XNOR U7691 ( .A(p_input[3196]), .B(n7967), .Z(n7970) );
  XOR U7692 ( .A(n7967), .B(p_input[3180]), .Z(n7969) );
  XOR U7693 ( .A(n7971), .B(n7972), .Z(n7967) );
  AND U7694 ( .A(n7973), .B(n7974), .Z(n7972) );
  XNOR U7695 ( .A(p_input[3195]), .B(n7971), .Z(n7974) );
  XOR U7696 ( .A(n7971), .B(p_input[3179]), .Z(n7973) );
  XOR U7697 ( .A(n7975), .B(n7976), .Z(n7971) );
  AND U7698 ( .A(n7977), .B(n7978), .Z(n7976) );
  XNOR U7699 ( .A(p_input[3194]), .B(n7975), .Z(n7978) );
  XOR U7700 ( .A(n7975), .B(p_input[3178]), .Z(n7977) );
  XOR U7701 ( .A(n7979), .B(n7980), .Z(n7975) );
  AND U7702 ( .A(n7981), .B(n7982), .Z(n7980) );
  XNOR U7703 ( .A(p_input[3193]), .B(n7979), .Z(n7982) );
  XOR U7704 ( .A(n7979), .B(p_input[3177]), .Z(n7981) );
  XOR U7705 ( .A(n7983), .B(n7984), .Z(n7979) );
  AND U7706 ( .A(n7985), .B(n7986), .Z(n7984) );
  XNOR U7707 ( .A(p_input[3192]), .B(n7983), .Z(n7986) );
  XOR U7708 ( .A(n7983), .B(p_input[3176]), .Z(n7985) );
  XOR U7709 ( .A(n7987), .B(n7988), .Z(n7983) );
  AND U7710 ( .A(n7989), .B(n7990), .Z(n7988) );
  XNOR U7711 ( .A(p_input[3191]), .B(n7987), .Z(n7990) );
  XOR U7712 ( .A(n7987), .B(p_input[3175]), .Z(n7989) );
  XOR U7713 ( .A(n7991), .B(n7992), .Z(n7987) );
  AND U7714 ( .A(n7993), .B(n7994), .Z(n7992) );
  XNOR U7715 ( .A(p_input[3190]), .B(n7991), .Z(n7994) );
  XOR U7716 ( .A(n7991), .B(p_input[3174]), .Z(n7993) );
  XOR U7717 ( .A(n7995), .B(n7996), .Z(n7991) );
  AND U7718 ( .A(n7997), .B(n7998), .Z(n7996) );
  XNOR U7719 ( .A(p_input[3189]), .B(n7995), .Z(n7998) );
  XOR U7720 ( .A(n7995), .B(p_input[3173]), .Z(n7997) );
  XOR U7721 ( .A(n7999), .B(n8000), .Z(n7995) );
  AND U7722 ( .A(n8001), .B(n8002), .Z(n8000) );
  XNOR U7723 ( .A(p_input[3188]), .B(n7999), .Z(n8002) );
  XOR U7724 ( .A(n7999), .B(p_input[3172]), .Z(n8001) );
  XOR U7725 ( .A(n8003), .B(n8004), .Z(n7999) );
  AND U7726 ( .A(n8005), .B(n8006), .Z(n8004) );
  XNOR U7727 ( .A(p_input[3187]), .B(n8003), .Z(n8006) );
  XOR U7728 ( .A(n8003), .B(p_input[3171]), .Z(n8005) );
  XOR U7729 ( .A(n8007), .B(n8008), .Z(n8003) );
  AND U7730 ( .A(n8009), .B(n8010), .Z(n8008) );
  XNOR U7731 ( .A(p_input[3186]), .B(n8007), .Z(n8010) );
  XOR U7732 ( .A(n8007), .B(p_input[3170]), .Z(n8009) );
  XNOR U7733 ( .A(n8011), .B(n8012), .Z(n8007) );
  AND U7734 ( .A(n8013), .B(n8014), .Z(n8012) );
  XOR U7735 ( .A(p_input[3185]), .B(n8011), .Z(n8014) );
  XNOR U7736 ( .A(p_input[3169]), .B(n8011), .Z(n8013) );
  AND U7737 ( .A(p_input[3184]), .B(n8015), .Z(n8011) );
  IV U7738 ( .A(p_input[3168]), .Z(n8015) );
  XNOR U7739 ( .A(p_input[3136]), .B(n8016), .Z(n7818) );
  AND U7740 ( .A(n205), .B(n8017), .Z(n8016) );
  XOR U7741 ( .A(p_input[3152]), .B(p_input[3136]), .Z(n8017) );
  XOR U7742 ( .A(n8018), .B(n8019), .Z(n205) );
  AND U7743 ( .A(n8020), .B(n8021), .Z(n8019) );
  XNOR U7744 ( .A(p_input[3167]), .B(n8018), .Z(n8021) );
  XOR U7745 ( .A(n8018), .B(p_input[3151]), .Z(n8020) );
  XOR U7746 ( .A(n8022), .B(n8023), .Z(n8018) );
  AND U7747 ( .A(n8024), .B(n8025), .Z(n8023) );
  XNOR U7748 ( .A(p_input[3166]), .B(n8022), .Z(n8025) );
  XNOR U7749 ( .A(n8022), .B(n7832), .Z(n8024) );
  IV U7750 ( .A(p_input[3150]), .Z(n7832) );
  XOR U7751 ( .A(n8026), .B(n8027), .Z(n8022) );
  AND U7752 ( .A(n8028), .B(n8029), .Z(n8027) );
  XNOR U7753 ( .A(p_input[3165]), .B(n8026), .Z(n8029) );
  XNOR U7754 ( .A(n8026), .B(n7841), .Z(n8028) );
  IV U7755 ( .A(p_input[3149]), .Z(n7841) );
  XOR U7756 ( .A(n8030), .B(n8031), .Z(n8026) );
  AND U7757 ( .A(n8032), .B(n8033), .Z(n8031) );
  XNOR U7758 ( .A(p_input[3164]), .B(n8030), .Z(n8033) );
  XNOR U7759 ( .A(n8030), .B(n7850), .Z(n8032) );
  IV U7760 ( .A(p_input[3148]), .Z(n7850) );
  XOR U7761 ( .A(n8034), .B(n8035), .Z(n8030) );
  AND U7762 ( .A(n8036), .B(n8037), .Z(n8035) );
  XNOR U7763 ( .A(p_input[3163]), .B(n8034), .Z(n8037) );
  XNOR U7764 ( .A(n8034), .B(n7859), .Z(n8036) );
  IV U7765 ( .A(p_input[3147]), .Z(n7859) );
  XOR U7766 ( .A(n8038), .B(n8039), .Z(n8034) );
  AND U7767 ( .A(n8040), .B(n8041), .Z(n8039) );
  XNOR U7768 ( .A(p_input[3162]), .B(n8038), .Z(n8041) );
  XNOR U7769 ( .A(n8038), .B(n7868), .Z(n8040) );
  IV U7770 ( .A(p_input[3146]), .Z(n7868) );
  XOR U7771 ( .A(n8042), .B(n8043), .Z(n8038) );
  AND U7772 ( .A(n8044), .B(n8045), .Z(n8043) );
  XNOR U7773 ( .A(p_input[3161]), .B(n8042), .Z(n8045) );
  XNOR U7774 ( .A(n8042), .B(n7877), .Z(n8044) );
  IV U7775 ( .A(p_input[3145]), .Z(n7877) );
  XOR U7776 ( .A(n8046), .B(n8047), .Z(n8042) );
  AND U7777 ( .A(n8048), .B(n8049), .Z(n8047) );
  XNOR U7778 ( .A(p_input[3160]), .B(n8046), .Z(n8049) );
  XNOR U7779 ( .A(n8046), .B(n7886), .Z(n8048) );
  IV U7780 ( .A(p_input[3144]), .Z(n7886) );
  XOR U7781 ( .A(n8050), .B(n8051), .Z(n8046) );
  AND U7782 ( .A(n8052), .B(n8053), .Z(n8051) );
  XNOR U7783 ( .A(p_input[3159]), .B(n8050), .Z(n8053) );
  XNOR U7784 ( .A(n8050), .B(n7895), .Z(n8052) );
  IV U7785 ( .A(p_input[3143]), .Z(n7895) );
  XOR U7786 ( .A(n8054), .B(n8055), .Z(n8050) );
  AND U7787 ( .A(n8056), .B(n8057), .Z(n8055) );
  XNOR U7788 ( .A(p_input[3158]), .B(n8054), .Z(n8057) );
  XNOR U7789 ( .A(n8054), .B(n7904), .Z(n8056) );
  IV U7790 ( .A(p_input[3142]), .Z(n7904) );
  XOR U7791 ( .A(n8058), .B(n8059), .Z(n8054) );
  AND U7792 ( .A(n8060), .B(n8061), .Z(n8059) );
  XNOR U7793 ( .A(p_input[3157]), .B(n8058), .Z(n8061) );
  XNOR U7794 ( .A(n8058), .B(n7913), .Z(n8060) );
  IV U7795 ( .A(p_input[3141]), .Z(n7913) );
  XOR U7796 ( .A(n8062), .B(n8063), .Z(n8058) );
  AND U7797 ( .A(n8064), .B(n8065), .Z(n8063) );
  XNOR U7798 ( .A(p_input[3156]), .B(n8062), .Z(n8065) );
  XNOR U7799 ( .A(n8062), .B(n7922), .Z(n8064) );
  IV U7800 ( .A(p_input[3140]), .Z(n7922) );
  XOR U7801 ( .A(n8066), .B(n8067), .Z(n8062) );
  AND U7802 ( .A(n8068), .B(n8069), .Z(n8067) );
  XNOR U7803 ( .A(p_input[3155]), .B(n8066), .Z(n8069) );
  XNOR U7804 ( .A(n8066), .B(n7931), .Z(n8068) );
  IV U7805 ( .A(p_input[3139]), .Z(n7931) );
  XOR U7806 ( .A(n8070), .B(n8071), .Z(n8066) );
  AND U7807 ( .A(n8072), .B(n8073), .Z(n8071) );
  XNOR U7808 ( .A(p_input[3154]), .B(n8070), .Z(n8073) );
  XNOR U7809 ( .A(n8070), .B(n7940), .Z(n8072) );
  IV U7810 ( .A(p_input[3138]), .Z(n7940) );
  XNOR U7811 ( .A(n8074), .B(n8075), .Z(n8070) );
  AND U7812 ( .A(n8076), .B(n8077), .Z(n8075) );
  XOR U7813 ( .A(p_input[3153]), .B(n8074), .Z(n8077) );
  XNOR U7814 ( .A(p_input[3137]), .B(n8074), .Z(n8076) );
  AND U7815 ( .A(p_input[3152]), .B(n8078), .Z(n8074) );
  IV U7816 ( .A(p_input[3136]), .Z(n8078) );
  XOR U7817 ( .A(n8079), .B(n8080), .Z(n7637) );
  AND U7818 ( .A(n400), .B(n8081), .Z(n8080) );
  XNOR U7819 ( .A(n8082), .B(n8079), .Z(n8081) );
  XOR U7820 ( .A(n8083), .B(n8084), .Z(n400) );
  AND U7821 ( .A(n8085), .B(n8086), .Z(n8084) );
  XNOR U7822 ( .A(n7648), .B(n8083), .Z(n8086) );
  AND U7823 ( .A(p_input[3135]), .B(p_input[3119]), .Z(n7648) );
  XOR U7824 ( .A(n8083), .B(n7647), .Z(n8085) );
  AND U7825 ( .A(p_input[3087]), .B(p_input[3103]), .Z(n7647) );
  XOR U7826 ( .A(n8087), .B(n8088), .Z(n8083) );
  AND U7827 ( .A(n8089), .B(n8090), .Z(n8088) );
  XOR U7828 ( .A(n8087), .B(n7660), .Z(n8090) );
  XNOR U7829 ( .A(p_input[3118]), .B(n8091), .Z(n7660) );
  AND U7830 ( .A(n211), .B(n8092), .Z(n8091) );
  XOR U7831 ( .A(p_input[3134]), .B(p_input[3118]), .Z(n8092) );
  XNOR U7832 ( .A(n7657), .B(n8087), .Z(n8089) );
  XOR U7833 ( .A(n8093), .B(n8094), .Z(n7657) );
  AND U7834 ( .A(n208), .B(n8095), .Z(n8094) );
  XOR U7835 ( .A(p_input[3102]), .B(p_input[3086]), .Z(n8095) );
  XOR U7836 ( .A(n8096), .B(n8097), .Z(n8087) );
  AND U7837 ( .A(n8098), .B(n8099), .Z(n8097) );
  XOR U7838 ( .A(n8096), .B(n7672), .Z(n8099) );
  XNOR U7839 ( .A(p_input[3117]), .B(n8100), .Z(n7672) );
  AND U7840 ( .A(n211), .B(n8101), .Z(n8100) );
  XOR U7841 ( .A(p_input[3133]), .B(p_input[3117]), .Z(n8101) );
  XNOR U7842 ( .A(n7669), .B(n8096), .Z(n8098) );
  XOR U7843 ( .A(n8102), .B(n8103), .Z(n7669) );
  AND U7844 ( .A(n208), .B(n8104), .Z(n8103) );
  XOR U7845 ( .A(p_input[3101]), .B(p_input[3085]), .Z(n8104) );
  XOR U7846 ( .A(n8105), .B(n8106), .Z(n8096) );
  AND U7847 ( .A(n8107), .B(n8108), .Z(n8106) );
  XOR U7848 ( .A(n8105), .B(n7684), .Z(n8108) );
  XNOR U7849 ( .A(p_input[3116]), .B(n8109), .Z(n7684) );
  AND U7850 ( .A(n211), .B(n8110), .Z(n8109) );
  XOR U7851 ( .A(p_input[3132]), .B(p_input[3116]), .Z(n8110) );
  XNOR U7852 ( .A(n7681), .B(n8105), .Z(n8107) );
  XOR U7853 ( .A(n8111), .B(n8112), .Z(n7681) );
  AND U7854 ( .A(n208), .B(n8113), .Z(n8112) );
  XOR U7855 ( .A(p_input[3100]), .B(p_input[3084]), .Z(n8113) );
  XOR U7856 ( .A(n8114), .B(n8115), .Z(n8105) );
  AND U7857 ( .A(n8116), .B(n8117), .Z(n8115) );
  XOR U7858 ( .A(n8114), .B(n7696), .Z(n8117) );
  XNOR U7859 ( .A(p_input[3115]), .B(n8118), .Z(n7696) );
  AND U7860 ( .A(n211), .B(n8119), .Z(n8118) );
  XOR U7861 ( .A(p_input[3131]), .B(p_input[3115]), .Z(n8119) );
  XNOR U7862 ( .A(n7693), .B(n8114), .Z(n8116) );
  XOR U7863 ( .A(n8120), .B(n8121), .Z(n7693) );
  AND U7864 ( .A(n208), .B(n8122), .Z(n8121) );
  XOR U7865 ( .A(p_input[3099]), .B(p_input[3083]), .Z(n8122) );
  XOR U7866 ( .A(n8123), .B(n8124), .Z(n8114) );
  AND U7867 ( .A(n8125), .B(n8126), .Z(n8124) );
  XOR U7868 ( .A(n8123), .B(n7708), .Z(n8126) );
  XNOR U7869 ( .A(p_input[3114]), .B(n8127), .Z(n7708) );
  AND U7870 ( .A(n211), .B(n8128), .Z(n8127) );
  XOR U7871 ( .A(p_input[3130]), .B(p_input[3114]), .Z(n8128) );
  XNOR U7872 ( .A(n7705), .B(n8123), .Z(n8125) );
  XOR U7873 ( .A(n8129), .B(n8130), .Z(n7705) );
  AND U7874 ( .A(n208), .B(n8131), .Z(n8130) );
  XOR U7875 ( .A(p_input[3098]), .B(p_input[3082]), .Z(n8131) );
  XOR U7876 ( .A(n8132), .B(n8133), .Z(n8123) );
  AND U7877 ( .A(n8134), .B(n8135), .Z(n8133) );
  XOR U7878 ( .A(n8132), .B(n7720), .Z(n8135) );
  XNOR U7879 ( .A(p_input[3113]), .B(n8136), .Z(n7720) );
  AND U7880 ( .A(n211), .B(n8137), .Z(n8136) );
  XOR U7881 ( .A(p_input[3129]), .B(p_input[3113]), .Z(n8137) );
  XNOR U7882 ( .A(n7717), .B(n8132), .Z(n8134) );
  XOR U7883 ( .A(n8138), .B(n8139), .Z(n7717) );
  AND U7884 ( .A(n208), .B(n8140), .Z(n8139) );
  XOR U7885 ( .A(p_input[3097]), .B(p_input[3081]), .Z(n8140) );
  XOR U7886 ( .A(n8141), .B(n8142), .Z(n8132) );
  AND U7887 ( .A(n8143), .B(n8144), .Z(n8142) );
  XOR U7888 ( .A(n8141), .B(n7732), .Z(n8144) );
  XNOR U7889 ( .A(p_input[3112]), .B(n8145), .Z(n7732) );
  AND U7890 ( .A(n211), .B(n8146), .Z(n8145) );
  XOR U7891 ( .A(p_input[3128]), .B(p_input[3112]), .Z(n8146) );
  XNOR U7892 ( .A(n7729), .B(n8141), .Z(n8143) );
  XOR U7893 ( .A(n8147), .B(n8148), .Z(n7729) );
  AND U7894 ( .A(n208), .B(n8149), .Z(n8148) );
  XOR U7895 ( .A(p_input[3096]), .B(p_input[3080]), .Z(n8149) );
  XOR U7896 ( .A(n8150), .B(n8151), .Z(n8141) );
  AND U7897 ( .A(n8152), .B(n8153), .Z(n8151) );
  XOR U7898 ( .A(n8150), .B(n7744), .Z(n8153) );
  XNOR U7899 ( .A(p_input[3111]), .B(n8154), .Z(n7744) );
  AND U7900 ( .A(n211), .B(n8155), .Z(n8154) );
  XOR U7901 ( .A(p_input[3127]), .B(p_input[3111]), .Z(n8155) );
  XNOR U7902 ( .A(n7741), .B(n8150), .Z(n8152) );
  XOR U7903 ( .A(n8156), .B(n8157), .Z(n7741) );
  AND U7904 ( .A(n208), .B(n8158), .Z(n8157) );
  XOR U7905 ( .A(p_input[3095]), .B(p_input[3079]), .Z(n8158) );
  XOR U7906 ( .A(n8159), .B(n8160), .Z(n8150) );
  AND U7907 ( .A(n8161), .B(n8162), .Z(n8160) );
  XOR U7908 ( .A(n8159), .B(n7756), .Z(n8162) );
  XNOR U7909 ( .A(p_input[3110]), .B(n8163), .Z(n7756) );
  AND U7910 ( .A(n211), .B(n8164), .Z(n8163) );
  XOR U7911 ( .A(p_input[3126]), .B(p_input[3110]), .Z(n8164) );
  XNOR U7912 ( .A(n7753), .B(n8159), .Z(n8161) );
  XOR U7913 ( .A(n8165), .B(n8166), .Z(n7753) );
  AND U7914 ( .A(n208), .B(n8167), .Z(n8166) );
  XOR U7915 ( .A(p_input[3094]), .B(p_input[3078]), .Z(n8167) );
  XOR U7916 ( .A(n8168), .B(n8169), .Z(n8159) );
  AND U7917 ( .A(n8170), .B(n8171), .Z(n8169) );
  XOR U7918 ( .A(n8168), .B(n7768), .Z(n8171) );
  XNOR U7919 ( .A(p_input[3109]), .B(n8172), .Z(n7768) );
  AND U7920 ( .A(n211), .B(n8173), .Z(n8172) );
  XOR U7921 ( .A(p_input[3125]), .B(p_input[3109]), .Z(n8173) );
  XNOR U7922 ( .A(n7765), .B(n8168), .Z(n8170) );
  XOR U7923 ( .A(n8174), .B(n8175), .Z(n7765) );
  AND U7924 ( .A(n208), .B(n8176), .Z(n8175) );
  XOR U7925 ( .A(p_input[3093]), .B(p_input[3077]), .Z(n8176) );
  XOR U7926 ( .A(n8177), .B(n8178), .Z(n8168) );
  AND U7927 ( .A(n8179), .B(n8180), .Z(n8178) );
  XOR U7928 ( .A(n8177), .B(n7780), .Z(n8180) );
  XNOR U7929 ( .A(p_input[3108]), .B(n8181), .Z(n7780) );
  AND U7930 ( .A(n211), .B(n8182), .Z(n8181) );
  XOR U7931 ( .A(p_input[3124]), .B(p_input[3108]), .Z(n8182) );
  XNOR U7932 ( .A(n7777), .B(n8177), .Z(n8179) );
  XOR U7933 ( .A(n8183), .B(n8184), .Z(n7777) );
  AND U7934 ( .A(n208), .B(n8185), .Z(n8184) );
  XOR U7935 ( .A(p_input[3092]), .B(p_input[3076]), .Z(n8185) );
  XOR U7936 ( .A(n8186), .B(n8187), .Z(n8177) );
  AND U7937 ( .A(n8188), .B(n8189), .Z(n8187) );
  XOR U7938 ( .A(n8186), .B(n7792), .Z(n8189) );
  XNOR U7939 ( .A(p_input[3107]), .B(n8190), .Z(n7792) );
  AND U7940 ( .A(n211), .B(n8191), .Z(n8190) );
  XOR U7941 ( .A(p_input[3123]), .B(p_input[3107]), .Z(n8191) );
  XNOR U7942 ( .A(n7789), .B(n8186), .Z(n8188) );
  XOR U7943 ( .A(n8192), .B(n8193), .Z(n7789) );
  AND U7944 ( .A(n208), .B(n8194), .Z(n8193) );
  XOR U7945 ( .A(p_input[3091]), .B(p_input[3075]), .Z(n8194) );
  XOR U7946 ( .A(n8195), .B(n8196), .Z(n8186) );
  AND U7947 ( .A(n8197), .B(n8198), .Z(n8196) );
  XOR U7948 ( .A(n8195), .B(n7804), .Z(n8198) );
  XNOR U7949 ( .A(p_input[3106]), .B(n8199), .Z(n7804) );
  AND U7950 ( .A(n211), .B(n8200), .Z(n8199) );
  XOR U7951 ( .A(p_input[3122]), .B(p_input[3106]), .Z(n8200) );
  XNOR U7952 ( .A(n7801), .B(n8195), .Z(n8197) );
  XOR U7953 ( .A(n8201), .B(n8202), .Z(n7801) );
  AND U7954 ( .A(n208), .B(n8203), .Z(n8202) );
  XOR U7955 ( .A(p_input[3090]), .B(p_input[3074]), .Z(n8203) );
  XOR U7956 ( .A(n8204), .B(n8205), .Z(n8195) );
  AND U7957 ( .A(n8206), .B(n8207), .Z(n8205) );
  XNOR U7958 ( .A(n8208), .B(n7817), .Z(n8207) );
  XNOR U7959 ( .A(p_input[3105]), .B(n8209), .Z(n7817) );
  AND U7960 ( .A(n211), .B(n8210), .Z(n8209) );
  XNOR U7961 ( .A(p_input[3121]), .B(n8211), .Z(n8210) );
  IV U7962 ( .A(p_input[3105]), .Z(n8211) );
  XNOR U7963 ( .A(n7814), .B(n8204), .Z(n8206) );
  XNOR U7964 ( .A(p_input[3073]), .B(n8212), .Z(n7814) );
  AND U7965 ( .A(n208), .B(n8213), .Z(n8212) );
  XOR U7966 ( .A(p_input[3089]), .B(p_input[3073]), .Z(n8213) );
  IV U7967 ( .A(n8208), .Z(n8204) );
  AND U7968 ( .A(n8079), .B(n8082), .Z(n8208) );
  XOR U7969 ( .A(p_input[3104]), .B(n8214), .Z(n8082) );
  AND U7970 ( .A(n211), .B(n8215), .Z(n8214) );
  XOR U7971 ( .A(p_input[3120]), .B(p_input[3104]), .Z(n8215) );
  XOR U7972 ( .A(n8216), .B(n8217), .Z(n211) );
  AND U7973 ( .A(n8218), .B(n8219), .Z(n8217) );
  XNOR U7974 ( .A(p_input[3135]), .B(n8216), .Z(n8219) );
  XOR U7975 ( .A(n8216), .B(p_input[3119]), .Z(n8218) );
  XOR U7976 ( .A(n8220), .B(n8221), .Z(n8216) );
  AND U7977 ( .A(n8222), .B(n8223), .Z(n8221) );
  XNOR U7978 ( .A(p_input[3134]), .B(n8220), .Z(n8223) );
  XOR U7979 ( .A(n8220), .B(p_input[3118]), .Z(n8222) );
  XOR U7980 ( .A(n8224), .B(n8225), .Z(n8220) );
  AND U7981 ( .A(n8226), .B(n8227), .Z(n8225) );
  XNOR U7982 ( .A(p_input[3133]), .B(n8224), .Z(n8227) );
  XOR U7983 ( .A(n8224), .B(p_input[3117]), .Z(n8226) );
  XOR U7984 ( .A(n8228), .B(n8229), .Z(n8224) );
  AND U7985 ( .A(n8230), .B(n8231), .Z(n8229) );
  XNOR U7986 ( .A(p_input[3132]), .B(n8228), .Z(n8231) );
  XOR U7987 ( .A(n8228), .B(p_input[3116]), .Z(n8230) );
  XOR U7988 ( .A(n8232), .B(n8233), .Z(n8228) );
  AND U7989 ( .A(n8234), .B(n8235), .Z(n8233) );
  XNOR U7990 ( .A(p_input[3131]), .B(n8232), .Z(n8235) );
  XOR U7991 ( .A(n8232), .B(p_input[3115]), .Z(n8234) );
  XOR U7992 ( .A(n8236), .B(n8237), .Z(n8232) );
  AND U7993 ( .A(n8238), .B(n8239), .Z(n8237) );
  XNOR U7994 ( .A(p_input[3130]), .B(n8236), .Z(n8239) );
  XOR U7995 ( .A(n8236), .B(p_input[3114]), .Z(n8238) );
  XOR U7996 ( .A(n8240), .B(n8241), .Z(n8236) );
  AND U7997 ( .A(n8242), .B(n8243), .Z(n8241) );
  XNOR U7998 ( .A(p_input[3129]), .B(n8240), .Z(n8243) );
  XOR U7999 ( .A(n8240), .B(p_input[3113]), .Z(n8242) );
  XOR U8000 ( .A(n8244), .B(n8245), .Z(n8240) );
  AND U8001 ( .A(n8246), .B(n8247), .Z(n8245) );
  XNOR U8002 ( .A(p_input[3128]), .B(n8244), .Z(n8247) );
  XOR U8003 ( .A(n8244), .B(p_input[3112]), .Z(n8246) );
  XOR U8004 ( .A(n8248), .B(n8249), .Z(n8244) );
  AND U8005 ( .A(n8250), .B(n8251), .Z(n8249) );
  XNOR U8006 ( .A(p_input[3127]), .B(n8248), .Z(n8251) );
  XOR U8007 ( .A(n8248), .B(p_input[3111]), .Z(n8250) );
  XOR U8008 ( .A(n8252), .B(n8253), .Z(n8248) );
  AND U8009 ( .A(n8254), .B(n8255), .Z(n8253) );
  XNOR U8010 ( .A(p_input[3126]), .B(n8252), .Z(n8255) );
  XOR U8011 ( .A(n8252), .B(p_input[3110]), .Z(n8254) );
  XOR U8012 ( .A(n8256), .B(n8257), .Z(n8252) );
  AND U8013 ( .A(n8258), .B(n8259), .Z(n8257) );
  XNOR U8014 ( .A(p_input[3125]), .B(n8256), .Z(n8259) );
  XOR U8015 ( .A(n8256), .B(p_input[3109]), .Z(n8258) );
  XOR U8016 ( .A(n8260), .B(n8261), .Z(n8256) );
  AND U8017 ( .A(n8262), .B(n8263), .Z(n8261) );
  XNOR U8018 ( .A(p_input[3124]), .B(n8260), .Z(n8263) );
  XOR U8019 ( .A(n8260), .B(p_input[3108]), .Z(n8262) );
  XOR U8020 ( .A(n8264), .B(n8265), .Z(n8260) );
  AND U8021 ( .A(n8266), .B(n8267), .Z(n8265) );
  XNOR U8022 ( .A(p_input[3123]), .B(n8264), .Z(n8267) );
  XOR U8023 ( .A(n8264), .B(p_input[3107]), .Z(n8266) );
  XOR U8024 ( .A(n8268), .B(n8269), .Z(n8264) );
  AND U8025 ( .A(n8270), .B(n8271), .Z(n8269) );
  XNOR U8026 ( .A(p_input[3122]), .B(n8268), .Z(n8271) );
  XOR U8027 ( .A(n8268), .B(p_input[3106]), .Z(n8270) );
  XNOR U8028 ( .A(n8272), .B(n8273), .Z(n8268) );
  AND U8029 ( .A(n8274), .B(n8275), .Z(n8273) );
  XOR U8030 ( .A(p_input[3121]), .B(n8272), .Z(n8275) );
  XNOR U8031 ( .A(p_input[3105]), .B(n8272), .Z(n8274) );
  AND U8032 ( .A(p_input[3120]), .B(n8276), .Z(n8272) );
  IV U8033 ( .A(p_input[3104]), .Z(n8276) );
  XNOR U8034 ( .A(p_input[3072]), .B(n8277), .Z(n8079) );
  AND U8035 ( .A(n208), .B(n8278), .Z(n8277) );
  XOR U8036 ( .A(p_input[3088]), .B(p_input[3072]), .Z(n8278) );
  XOR U8037 ( .A(n8279), .B(n8280), .Z(n208) );
  AND U8038 ( .A(n8281), .B(n8282), .Z(n8280) );
  XNOR U8039 ( .A(p_input[3103]), .B(n8279), .Z(n8282) );
  XOR U8040 ( .A(n8279), .B(p_input[3087]), .Z(n8281) );
  XOR U8041 ( .A(n8283), .B(n8284), .Z(n8279) );
  AND U8042 ( .A(n8285), .B(n8286), .Z(n8284) );
  XNOR U8043 ( .A(p_input[3102]), .B(n8283), .Z(n8286) );
  XNOR U8044 ( .A(n8283), .B(n8093), .Z(n8285) );
  IV U8045 ( .A(p_input[3086]), .Z(n8093) );
  XOR U8046 ( .A(n8287), .B(n8288), .Z(n8283) );
  AND U8047 ( .A(n8289), .B(n8290), .Z(n8288) );
  XNOR U8048 ( .A(p_input[3101]), .B(n8287), .Z(n8290) );
  XNOR U8049 ( .A(n8287), .B(n8102), .Z(n8289) );
  IV U8050 ( .A(p_input[3085]), .Z(n8102) );
  XOR U8051 ( .A(n8291), .B(n8292), .Z(n8287) );
  AND U8052 ( .A(n8293), .B(n8294), .Z(n8292) );
  XNOR U8053 ( .A(p_input[3100]), .B(n8291), .Z(n8294) );
  XNOR U8054 ( .A(n8291), .B(n8111), .Z(n8293) );
  IV U8055 ( .A(p_input[3084]), .Z(n8111) );
  XOR U8056 ( .A(n8295), .B(n8296), .Z(n8291) );
  AND U8057 ( .A(n8297), .B(n8298), .Z(n8296) );
  XNOR U8058 ( .A(p_input[3099]), .B(n8295), .Z(n8298) );
  XNOR U8059 ( .A(n8295), .B(n8120), .Z(n8297) );
  IV U8060 ( .A(p_input[3083]), .Z(n8120) );
  XOR U8061 ( .A(n8299), .B(n8300), .Z(n8295) );
  AND U8062 ( .A(n8301), .B(n8302), .Z(n8300) );
  XNOR U8063 ( .A(p_input[3098]), .B(n8299), .Z(n8302) );
  XNOR U8064 ( .A(n8299), .B(n8129), .Z(n8301) );
  IV U8065 ( .A(p_input[3082]), .Z(n8129) );
  XOR U8066 ( .A(n8303), .B(n8304), .Z(n8299) );
  AND U8067 ( .A(n8305), .B(n8306), .Z(n8304) );
  XNOR U8068 ( .A(p_input[3097]), .B(n8303), .Z(n8306) );
  XNOR U8069 ( .A(n8303), .B(n8138), .Z(n8305) );
  IV U8070 ( .A(p_input[3081]), .Z(n8138) );
  XOR U8071 ( .A(n8307), .B(n8308), .Z(n8303) );
  AND U8072 ( .A(n8309), .B(n8310), .Z(n8308) );
  XNOR U8073 ( .A(p_input[3096]), .B(n8307), .Z(n8310) );
  XNOR U8074 ( .A(n8307), .B(n8147), .Z(n8309) );
  IV U8075 ( .A(p_input[3080]), .Z(n8147) );
  XOR U8076 ( .A(n8311), .B(n8312), .Z(n8307) );
  AND U8077 ( .A(n8313), .B(n8314), .Z(n8312) );
  XNOR U8078 ( .A(p_input[3095]), .B(n8311), .Z(n8314) );
  XNOR U8079 ( .A(n8311), .B(n8156), .Z(n8313) );
  IV U8080 ( .A(p_input[3079]), .Z(n8156) );
  XOR U8081 ( .A(n8315), .B(n8316), .Z(n8311) );
  AND U8082 ( .A(n8317), .B(n8318), .Z(n8316) );
  XNOR U8083 ( .A(p_input[3094]), .B(n8315), .Z(n8318) );
  XNOR U8084 ( .A(n8315), .B(n8165), .Z(n8317) );
  IV U8085 ( .A(p_input[3078]), .Z(n8165) );
  XOR U8086 ( .A(n8319), .B(n8320), .Z(n8315) );
  AND U8087 ( .A(n8321), .B(n8322), .Z(n8320) );
  XNOR U8088 ( .A(p_input[3093]), .B(n8319), .Z(n8322) );
  XNOR U8089 ( .A(n8319), .B(n8174), .Z(n8321) );
  IV U8090 ( .A(p_input[3077]), .Z(n8174) );
  XOR U8091 ( .A(n8323), .B(n8324), .Z(n8319) );
  AND U8092 ( .A(n8325), .B(n8326), .Z(n8324) );
  XNOR U8093 ( .A(p_input[3092]), .B(n8323), .Z(n8326) );
  XNOR U8094 ( .A(n8323), .B(n8183), .Z(n8325) );
  IV U8095 ( .A(p_input[3076]), .Z(n8183) );
  XOR U8096 ( .A(n8327), .B(n8328), .Z(n8323) );
  AND U8097 ( .A(n8329), .B(n8330), .Z(n8328) );
  XNOR U8098 ( .A(p_input[3091]), .B(n8327), .Z(n8330) );
  XNOR U8099 ( .A(n8327), .B(n8192), .Z(n8329) );
  IV U8100 ( .A(p_input[3075]), .Z(n8192) );
  XOR U8101 ( .A(n8331), .B(n8332), .Z(n8327) );
  AND U8102 ( .A(n8333), .B(n8334), .Z(n8332) );
  XNOR U8103 ( .A(p_input[3090]), .B(n8331), .Z(n8334) );
  XNOR U8104 ( .A(n8331), .B(n8201), .Z(n8333) );
  IV U8105 ( .A(p_input[3074]), .Z(n8201) );
  XNOR U8106 ( .A(n8335), .B(n8336), .Z(n8331) );
  AND U8107 ( .A(n8337), .B(n8338), .Z(n8336) );
  XOR U8108 ( .A(p_input[3089]), .B(n8335), .Z(n8338) );
  XNOR U8109 ( .A(p_input[3073]), .B(n8335), .Z(n8337) );
  AND U8110 ( .A(p_input[3088]), .B(n8339), .Z(n8335) );
  IV U8111 ( .A(p_input[3072]), .Z(n8339) );
  XOR U8112 ( .A(n8340), .B(n8341), .Z(n1248) );
  AND U8113 ( .A(n1045), .B(n8342), .Z(n8341) );
  XNOR U8114 ( .A(n8343), .B(n8340), .Z(n8342) );
  XOR U8115 ( .A(n8344), .B(n8345), .Z(n1045) );
  AND U8116 ( .A(n8346), .B(n8347), .Z(n8345) );
  XOR U8117 ( .A(n8344), .B(n1263), .Z(n8347) );
  XOR U8118 ( .A(n8348), .B(n8349), .Z(n1263) );
  AND U8119 ( .A(n1011), .B(n8350), .Z(n8349) );
  XOR U8120 ( .A(n8351), .B(n8348), .Z(n8350) );
  XNOR U8121 ( .A(n1260), .B(n8344), .Z(n8346) );
  XOR U8122 ( .A(n8352), .B(n8353), .Z(n1260) );
  AND U8123 ( .A(n1008), .B(n8354), .Z(n8353) );
  XOR U8124 ( .A(n8355), .B(n8352), .Z(n8354) );
  XOR U8125 ( .A(n8356), .B(n8357), .Z(n8344) );
  AND U8126 ( .A(n8358), .B(n8359), .Z(n8357) );
  XOR U8127 ( .A(n8356), .B(n1275), .Z(n8359) );
  XOR U8128 ( .A(n8360), .B(n8361), .Z(n1275) );
  AND U8129 ( .A(n1011), .B(n8362), .Z(n8361) );
  XOR U8130 ( .A(n8363), .B(n8360), .Z(n8362) );
  XNOR U8131 ( .A(n1272), .B(n8356), .Z(n8358) );
  XOR U8132 ( .A(n8364), .B(n8365), .Z(n1272) );
  AND U8133 ( .A(n1008), .B(n8366), .Z(n8365) );
  XOR U8134 ( .A(n8367), .B(n8364), .Z(n8366) );
  XOR U8135 ( .A(n8368), .B(n8369), .Z(n8356) );
  AND U8136 ( .A(n8370), .B(n8371), .Z(n8369) );
  XOR U8137 ( .A(n8368), .B(n1287), .Z(n8371) );
  XOR U8138 ( .A(n8372), .B(n8373), .Z(n1287) );
  AND U8139 ( .A(n1011), .B(n8374), .Z(n8373) );
  XOR U8140 ( .A(n8375), .B(n8372), .Z(n8374) );
  XNOR U8141 ( .A(n1284), .B(n8368), .Z(n8370) );
  XOR U8142 ( .A(n8376), .B(n8377), .Z(n1284) );
  AND U8143 ( .A(n1008), .B(n8378), .Z(n8377) );
  XOR U8144 ( .A(n8379), .B(n8376), .Z(n8378) );
  XOR U8145 ( .A(n8380), .B(n8381), .Z(n8368) );
  AND U8146 ( .A(n8382), .B(n8383), .Z(n8381) );
  XOR U8147 ( .A(n8380), .B(n1299), .Z(n8383) );
  XOR U8148 ( .A(n8384), .B(n8385), .Z(n1299) );
  AND U8149 ( .A(n1011), .B(n8386), .Z(n8385) );
  XOR U8150 ( .A(n8387), .B(n8384), .Z(n8386) );
  XNOR U8151 ( .A(n1296), .B(n8380), .Z(n8382) );
  XOR U8152 ( .A(n8388), .B(n8389), .Z(n1296) );
  AND U8153 ( .A(n1008), .B(n8390), .Z(n8389) );
  XOR U8154 ( .A(n8391), .B(n8388), .Z(n8390) );
  XOR U8155 ( .A(n8392), .B(n8393), .Z(n8380) );
  AND U8156 ( .A(n8394), .B(n8395), .Z(n8393) );
  XOR U8157 ( .A(n8392), .B(n1311), .Z(n8395) );
  XOR U8158 ( .A(n8396), .B(n8397), .Z(n1311) );
  AND U8159 ( .A(n1011), .B(n8398), .Z(n8397) );
  XOR U8160 ( .A(n8399), .B(n8396), .Z(n8398) );
  XNOR U8161 ( .A(n1308), .B(n8392), .Z(n8394) );
  XOR U8162 ( .A(n8400), .B(n8401), .Z(n1308) );
  AND U8163 ( .A(n1008), .B(n8402), .Z(n8401) );
  XOR U8164 ( .A(n8403), .B(n8400), .Z(n8402) );
  XOR U8165 ( .A(n8404), .B(n8405), .Z(n8392) );
  AND U8166 ( .A(n8406), .B(n8407), .Z(n8405) );
  XOR U8167 ( .A(n8404), .B(n1323), .Z(n8407) );
  XOR U8168 ( .A(n8408), .B(n8409), .Z(n1323) );
  AND U8169 ( .A(n1011), .B(n8410), .Z(n8409) );
  XOR U8170 ( .A(n8411), .B(n8408), .Z(n8410) );
  XNOR U8171 ( .A(n1320), .B(n8404), .Z(n8406) );
  XOR U8172 ( .A(n8412), .B(n8413), .Z(n1320) );
  AND U8173 ( .A(n1008), .B(n8414), .Z(n8413) );
  XOR U8174 ( .A(n8415), .B(n8412), .Z(n8414) );
  XOR U8175 ( .A(n8416), .B(n8417), .Z(n8404) );
  AND U8176 ( .A(n8418), .B(n8419), .Z(n8417) );
  XOR U8177 ( .A(n8416), .B(n1335), .Z(n8419) );
  XOR U8178 ( .A(n8420), .B(n8421), .Z(n1335) );
  AND U8179 ( .A(n1011), .B(n8422), .Z(n8421) );
  XOR U8180 ( .A(n8423), .B(n8420), .Z(n8422) );
  XNOR U8181 ( .A(n1332), .B(n8416), .Z(n8418) );
  XOR U8182 ( .A(n8424), .B(n8425), .Z(n1332) );
  AND U8183 ( .A(n1008), .B(n8426), .Z(n8425) );
  XOR U8184 ( .A(n8427), .B(n8424), .Z(n8426) );
  XOR U8185 ( .A(n8428), .B(n8429), .Z(n8416) );
  AND U8186 ( .A(n8430), .B(n8431), .Z(n8429) );
  XOR U8187 ( .A(n8428), .B(n1347), .Z(n8431) );
  XOR U8188 ( .A(n8432), .B(n8433), .Z(n1347) );
  AND U8189 ( .A(n1011), .B(n8434), .Z(n8433) );
  XOR U8190 ( .A(n8435), .B(n8432), .Z(n8434) );
  XNOR U8191 ( .A(n1344), .B(n8428), .Z(n8430) );
  XOR U8192 ( .A(n8436), .B(n8437), .Z(n1344) );
  AND U8193 ( .A(n1008), .B(n8438), .Z(n8437) );
  XOR U8194 ( .A(n8439), .B(n8436), .Z(n8438) );
  XOR U8195 ( .A(n8440), .B(n8441), .Z(n8428) );
  AND U8196 ( .A(n8442), .B(n8443), .Z(n8441) );
  XOR U8197 ( .A(n8440), .B(n1359), .Z(n8443) );
  XOR U8198 ( .A(n8444), .B(n8445), .Z(n1359) );
  AND U8199 ( .A(n1011), .B(n8446), .Z(n8445) );
  XOR U8200 ( .A(n8447), .B(n8444), .Z(n8446) );
  XNOR U8201 ( .A(n1356), .B(n8440), .Z(n8442) );
  XOR U8202 ( .A(n8448), .B(n8449), .Z(n1356) );
  AND U8203 ( .A(n1008), .B(n8450), .Z(n8449) );
  XOR U8204 ( .A(n8451), .B(n8448), .Z(n8450) );
  XOR U8205 ( .A(n8452), .B(n8453), .Z(n8440) );
  AND U8206 ( .A(n8454), .B(n8455), .Z(n8453) );
  XOR U8207 ( .A(n8452), .B(n1371), .Z(n8455) );
  XOR U8208 ( .A(n8456), .B(n8457), .Z(n1371) );
  AND U8209 ( .A(n1011), .B(n8458), .Z(n8457) );
  XOR U8210 ( .A(n8459), .B(n8456), .Z(n8458) );
  XNOR U8211 ( .A(n1368), .B(n8452), .Z(n8454) );
  XOR U8212 ( .A(n8460), .B(n8461), .Z(n1368) );
  AND U8213 ( .A(n1008), .B(n8462), .Z(n8461) );
  XOR U8214 ( .A(n8463), .B(n8460), .Z(n8462) );
  XOR U8215 ( .A(n8464), .B(n8465), .Z(n8452) );
  AND U8216 ( .A(n8466), .B(n8467), .Z(n8465) );
  XOR U8217 ( .A(n8464), .B(n1383), .Z(n8467) );
  XOR U8218 ( .A(n8468), .B(n8469), .Z(n1383) );
  AND U8219 ( .A(n1011), .B(n8470), .Z(n8469) );
  XOR U8220 ( .A(n8471), .B(n8468), .Z(n8470) );
  XNOR U8221 ( .A(n1380), .B(n8464), .Z(n8466) );
  XOR U8222 ( .A(n8472), .B(n8473), .Z(n1380) );
  AND U8223 ( .A(n1008), .B(n8474), .Z(n8473) );
  XOR U8224 ( .A(n8475), .B(n8472), .Z(n8474) );
  XOR U8225 ( .A(n8476), .B(n8477), .Z(n8464) );
  AND U8226 ( .A(n8478), .B(n8479), .Z(n8477) );
  XOR U8227 ( .A(n8476), .B(n1395), .Z(n8479) );
  XOR U8228 ( .A(n8480), .B(n8481), .Z(n1395) );
  AND U8229 ( .A(n1011), .B(n8482), .Z(n8481) );
  XOR U8230 ( .A(n8483), .B(n8480), .Z(n8482) );
  XNOR U8231 ( .A(n1392), .B(n8476), .Z(n8478) );
  XOR U8232 ( .A(n8484), .B(n8485), .Z(n1392) );
  AND U8233 ( .A(n1008), .B(n8486), .Z(n8485) );
  XOR U8234 ( .A(n8487), .B(n8484), .Z(n8486) );
  XOR U8235 ( .A(n8488), .B(n8489), .Z(n8476) );
  AND U8236 ( .A(n8490), .B(n8491), .Z(n8489) );
  XOR U8237 ( .A(n8488), .B(n1407), .Z(n8491) );
  XOR U8238 ( .A(n8492), .B(n8493), .Z(n1407) );
  AND U8239 ( .A(n1011), .B(n8494), .Z(n8493) );
  XOR U8240 ( .A(n8495), .B(n8492), .Z(n8494) );
  XNOR U8241 ( .A(n1404), .B(n8488), .Z(n8490) );
  XOR U8242 ( .A(n8496), .B(n8497), .Z(n1404) );
  AND U8243 ( .A(n1008), .B(n8498), .Z(n8497) );
  XOR U8244 ( .A(n8499), .B(n8496), .Z(n8498) );
  XOR U8245 ( .A(n8500), .B(n8501), .Z(n8488) );
  AND U8246 ( .A(n8502), .B(n8503), .Z(n8501) );
  XOR U8247 ( .A(n8500), .B(n1419), .Z(n8503) );
  XOR U8248 ( .A(n8504), .B(n8505), .Z(n1419) );
  AND U8249 ( .A(n1011), .B(n8506), .Z(n8505) );
  XOR U8250 ( .A(n8507), .B(n8504), .Z(n8506) );
  XNOR U8251 ( .A(n1416), .B(n8500), .Z(n8502) );
  XOR U8252 ( .A(n8508), .B(n8509), .Z(n1416) );
  AND U8253 ( .A(n1008), .B(n8510), .Z(n8509) );
  XOR U8254 ( .A(n8511), .B(n8508), .Z(n8510) );
  XOR U8255 ( .A(n8512), .B(n8513), .Z(n8500) );
  AND U8256 ( .A(n8514), .B(n8515), .Z(n8513) );
  XNOR U8257 ( .A(n8516), .B(n1432), .Z(n8515) );
  XOR U8258 ( .A(n8517), .B(n8518), .Z(n1432) );
  AND U8259 ( .A(n1011), .B(n8519), .Z(n8518) );
  XOR U8260 ( .A(n8517), .B(n8520), .Z(n8519) );
  XNOR U8261 ( .A(n1429), .B(n8512), .Z(n8514) );
  XOR U8262 ( .A(n8521), .B(n8522), .Z(n1429) );
  AND U8263 ( .A(n1008), .B(n8523), .Z(n8522) );
  XOR U8264 ( .A(n8521), .B(n8524), .Z(n8523) );
  IV U8265 ( .A(n8516), .Z(n8512) );
  AND U8266 ( .A(n8340), .B(n8343), .Z(n8516) );
  XNOR U8267 ( .A(n8525), .B(n8526), .Z(n8343) );
  AND U8268 ( .A(n1011), .B(n8527), .Z(n8526) );
  XNOR U8269 ( .A(n8528), .B(n8525), .Z(n8527) );
  XOR U8270 ( .A(n8529), .B(n8530), .Z(n1011) );
  AND U8271 ( .A(n8531), .B(n8532), .Z(n8530) );
  XOR U8272 ( .A(n8529), .B(n8351), .Z(n8532) );
  XNOR U8273 ( .A(n8533), .B(n8534), .Z(n8351) );
  AND U8274 ( .A(n8535), .B(n931), .Z(n8534) );
  AND U8275 ( .A(n8533), .B(n8536), .Z(n8535) );
  XNOR U8276 ( .A(n8348), .B(n8529), .Z(n8531) );
  XOR U8277 ( .A(n8537), .B(n8538), .Z(n8348) );
  AND U8278 ( .A(n8539), .B(n929), .Z(n8538) );
  NOR U8279 ( .A(n8537), .B(n8540), .Z(n8539) );
  XOR U8280 ( .A(n8541), .B(n8542), .Z(n8529) );
  AND U8281 ( .A(n8543), .B(n8544), .Z(n8542) );
  XOR U8282 ( .A(n8541), .B(n8363), .Z(n8544) );
  XOR U8283 ( .A(n8545), .B(n8546), .Z(n8363) );
  AND U8284 ( .A(n931), .B(n8547), .Z(n8546) );
  XOR U8285 ( .A(n8548), .B(n8545), .Z(n8547) );
  XNOR U8286 ( .A(n8360), .B(n8541), .Z(n8543) );
  XOR U8287 ( .A(n8549), .B(n8550), .Z(n8360) );
  AND U8288 ( .A(n929), .B(n8551), .Z(n8550) );
  XOR U8289 ( .A(n8552), .B(n8549), .Z(n8551) );
  XOR U8290 ( .A(n8553), .B(n8554), .Z(n8541) );
  AND U8291 ( .A(n8555), .B(n8556), .Z(n8554) );
  XOR U8292 ( .A(n8553), .B(n8375), .Z(n8556) );
  XOR U8293 ( .A(n8557), .B(n8558), .Z(n8375) );
  AND U8294 ( .A(n931), .B(n8559), .Z(n8558) );
  XOR U8295 ( .A(n8560), .B(n8557), .Z(n8559) );
  XNOR U8296 ( .A(n8372), .B(n8553), .Z(n8555) );
  XOR U8297 ( .A(n8561), .B(n8562), .Z(n8372) );
  AND U8298 ( .A(n929), .B(n8563), .Z(n8562) );
  XOR U8299 ( .A(n8564), .B(n8561), .Z(n8563) );
  XOR U8300 ( .A(n8565), .B(n8566), .Z(n8553) );
  AND U8301 ( .A(n8567), .B(n8568), .Z(n8566) );
  XOR U8302 ( .A(n8565), .B(n8387), .Z(n8568) );
  XOR U8303 ( .A(n8569), .B(n8570), .Z(n8387) );
  AND U8304 ( .A(n931), .B(n8571), .Z(n8570) );
  XOR U8305 ( .A(n8572), .B(n8569), .Z(n8571) );
  XNOR U8306 ( .A(n8384), .B(n8565), .Z(n8567) );
  XOR U8307 ( .A(n8573), .B(n8574), .Z(n8384) );
  AND U8308 ( .A(n929), .B(n8575), .Z(n8574) );
  XOR U8309 ( .A(n8576), .B(n8573), .Z(n8575) );
  XOR U8310 ( .A(n8577), .B(n8578), .Z(n8565) );
  AND U8311 ( .A(n8579), .B(n8580), .Z(n8578) );
  XOR U8312 ( .A(n8577), .B(n8399), .Z(n8580) );
  XOR U8313 ( .A(n8581), .B(n8582), .Z(n8399) );
  AND U8314 ( .A(n931), .B(n8583), .Z(n8582) );
  XOR U8315 ( .A(n8584), .B(n8581), .Z(n8583) );
  XNOR U8316 ( .A(n8396), .B(n8577), .Z(n8579) );
  XOR U8317 ( .A(n8585), .B(n8586), .Z(n8396) );
  AND U8318 ( .A(n929), .B(n8587), .Z(n8586) );
  XOR U8319 ( .A(n8588), .B(n8585), .Z(n8587) );
  XOR U8320 ( .A(n8589), .B(n8590), .Z(n8577) );
  AND U8321 ( .A(n8591), .B(n8592), .Z(n8590) );
  XOR U8322 ( .A(n8589), .B(n8411), .Z(n8592) );
  XOR U8323 ( .A(n8593), .B(n8594), .Z(n8411) );
  AND U8324 ( .A(n931), .B(n8595), .Z(n8594) );
  XOR U8325 ( .A(n8596), .B(n8593), .Z(n8595) );
  XNOR U8326 ( .A(n8408), .B(n8589), .Z(n8591) );
  XOR U8327 ( .A(n8597), .B(n8598), .Z(n8408) );
  AND U8328 ( .A(n929), .B(n8599), .Z(n8598) );
  XOR U8329 ( .A(n8600), .B(n8597), .Z(n8599) );
  XOR U8330 ( .A(n8601), .B(n8602), .Z(n8589) );
  AND U8331 ( .A(n8603), .B(n8604), .Z(n8602) );
  XOR U8332 ( .A(n8601), .B(n8423), .Z(n8604) );
  XOR U8333 ( .A(n8605), .B(n8606), .Z(n8423) );
  AND U8334 ( .A(n931), .B(n8607), .Z(n8606) );
  XOR U8335 ( .A(n8608), .B(n8605), .Z(n8607) );
  XNOR U8336 ( .A(n8420), .B(n8601), .Z(n8603) );
  XOR U8337 ( .A(n8609), .B(n8610), .Z(n8420) );
  AND U8338 ( .A(n929), .B(n8611), .Z(n8610) );
  XOR U8339 ( .A(n8612), .B(n8609), .Z(n8611) );
  XOR U8340 ( .A(n8613), .B(n8614), .Z(n8601) );
  AND U8341 ( .A(n8615), .B(n8616), .Z(n8614) );
  XOR U8342 ( .A(n8613), .B(n8435), .Z(n8616) );
  XOR U8343 ( .A(n8617), .B(n8618), .Z(n8435) );
  AND U8344 ( .A(n931), .B(n8619), .Z(n8618) );
  XOR U8345 ( .A(n8620), .B(n8617), .Z(n8619) );
  XNOR U8346 ( .A(n8432), .B(n8613), .Z(n8615) );
  XOR U8347 ( .A(n8621), .B(n8622), .Z(n8432) );
  AND U8348 ( .A(n929), .B(n8623), .Z(n8622) );
  XOR U8349 ( .A(n8624), .B(n8621), .Z(n8623) );
  XOR U8350 ( .A(n8625), .B(n8626), .Z(n8613) );
  AND U8351 ( .A(n8627), .B(n8628), .Z(n8626) );
  XOR U8352 ( .A(n8625), .B(n8447), .Z(n8628) );
  XOR U8353 ( .A(n8629), .B(n8630), .Z(n8447) );
  AND U8354 ( .A(n931), .B(n8631), .Z(n8630) );
  XOR U8355 ( .A(n8632), .B(n8629), .Z(n8631) );
  XNOR U8356 ( .A(n8444), .B(n8625), .Z(n8627) );
  XOR U8357 ( .A(n8633), .B(n8634), .Z(n8444) );
  AND U8358 ( .A(n929), .B(n8635), .Z(n8634) );
  XOR U8359 ( .A(n8636), .B(n8633), .Z(n8635) );
  XOR U8360 ( .A(n8637), .B(n8638), .Z(n8625) );
  AND U8361 ( .A(n8639), .B(n8640), .Z(n8638) );
  XOR U8362 ( .A(n8637), .B(n8459), .Z(n8640) );
  XOR U8363 ( .A(n8641), .B(n8642), .Z(n8459) );
  AND U8364 ( .A(n931), .B(n8643), .Z(n8642) );
  XOR U8365 ( .A(n8644), .B(n8641), .Z(n8643) );
  XNOR U8366 ( .A(n8456), .B(n8637), .Z(n8639) );
  XOR U8367 ( .A(n8645), .B(n8646), .Z(n8456) );
  AND U8368 ( .A(n929), .B(n8647), .Z(n8646) );
  XOR U8369 ( .A(n8648), .B(n8645), .Z(n8647) );
  XOR U8370 ( .A(n8649), .B(n8650), .Z(n8637) );
  AND U8371 ( .A(n8651), .B(n8652), .Z(n8650) );
  XOR U8372 ( .A(n8649), .B(n8471), .Z(n8652) );
  XOR U8373 ( .A(n8653), .B(n8654), .Z(n8471) );
  AND U8374 ( .A(n931), .B(n8655), .Z(n8654) );
  XOR U8375 ( .A(n8656), .B(n8653), .Z(n8655) );
  XNOR U8376 ( .A(n8468), .B(n8649), .Z(n8651) );
  XOR U8377 ( .A(n8657), .B(n8658), .Z(n8468) );
  AND U8378 ( .A(n929), .B(n8659), .Z(n8658) );
  XOR U8379 ( .A(n8660), .B(n8657), .Z(n8659) );
  XOR U8380 ( .A(n8661), .B(n8662), .Z(n8649) );
  AND U8381 ( .A(n8663), .B(n8664), .Z(n8662) );
  XOR U8382 ( .A(n8661), .B(n8483), .Z(n8664) );
  XOR U8383 ( .A(n8665), .B(n8666), .Z(n8483) );
  AND U8384 ( .A(n931), .B(n8667), .Z(n8666) );
  XOR U8385 ( .A(n8668), .B(n8665), .Z(n8667) );
  XNOR U8386 ( .A(n8480), .B(n8661), .Z(n8663) );
  XOR U8387 ( .A(n8669), .B(n8670), .Z(n8480) );
  AND U8388 ( .A(n929), .B(n8671), .Z(n8670) );
  XOR U8389 ( .A(n8672), .B(n8669), .Z(n8671) );
  XOR U8390 ( .A(n8673), .B(n8674), .Z(n8661) );
  AND U8391 ( .A(n8675), .B(n8676), .Z(n8674) );
  XOR U8392 ( .A(n8673), .B(n8495), .Z(n8676) );
  XOR U8393 ( .A(n8677), .B(n8678), .Z(n8495) );
  AND U8394 ( .A(n931), .B(n8679), .Z(n8678) );
  XOR U8395 ( .A(n8680), .B(n8677), .Z(n8679) );
  XNOR U8396 ( .A(n8492), .B(n8673), .Z(n8675) );
  XOR U8397 ( .A(n8681), .B(n8682), .Z(n8492) );
  AND U8398 ( .A(n929), .B(n8683), .Z(n8682) );
  XOR U8399 ( .A(n8684), .B(n8681), .Z(n8683) );
  XOR U8400 ( .A(n8685), .B(n8686), .Z(n8673) );
  AND U8401 ( .A(n8687), .B(n8688), .Z(n8686) );
  XOR U8402 ( .A(n8685), .B(n8507), .Z(n8688) );
  XOR U8403 ( .A(n8689), .B(n8690), .Z(n8507) );
  AND U8404 ( .A(n931), .B(n8691), .Z(n8690) );
  XOR U8405 ( .A(n8692), .B(n8689), .Z(n8691) );
  XNOR U8406 ( .A(n8504), .B(n8685), .Z(n8687) );
  XOR U8407 ( .A(n8693), .B(n8694), .Z(n8504) );
  AND U8408 ( .A(n929), .B(n8695), .Z(n8694) );
  XOR U8409 ( .A(n8696), .B(n8693), .Z(n8695) );
  XOR U8410 ( .A(n8697), .B(n8698), .Z(n8685) );
  AND U8411 ( .A(n8699), .B(n8700), .Z(n8698) );
  XNOR U8412 ( .A(n8701), .B(n8520), .Z(n8700) );
  XOR U8413 ( .A(n8702), .B(n8703), .Z(n8520) );
  AND U8414 ( .A(n931), .B(n8704), .Z(n8703) );
  XOR U8415 ( .A(n8702), .B(n8705), .Z(n8704) );
  XNOR U8416 ( .A(n8517), .B(n8697), .Z(n8699) );
  XOR U8417 ( .A(n8706), .B(n8707), .Z(n8517) );
  AND U8418 ( .A(n929), .B(n8708), .Z(n8707) );
  XOR U8419 ( .A(n8706), .B(n8709), .Z(n8708) );
  IV U8420 ( .A(n8701), .Z(n8697) );
  AND U8421 ( .A(n8525), .B(n8528), .Z(n8701) );
  XNOR U8422 ( .A(n8710), .B(n8711), .Z(n8528) );
  AND U8423 ( .A(n931), .B(n8712), .Z(n8711) );
  XNOR U8424 ( .A(n8713), .B(n8710), .Z(n8712) );
  XOR U8425 ( .A(n8714), .B(n8715), .Z(n931) );
  AND U8426 ( .A(n8716), .B(n8717), .Z(n8715) );
  XOR U8427 ( .A(n8536), .B(n8714), .Z(n8717) );
  IV U8428 ( .A(n8718), .Z(n8536) );
  AND U8429 ( .A(n8719), .B(n8720), .Z(n8718) );
  XOR U8430 ( .A(n8714), .B(n8533), .Z(n8716) );
  AND U8431 ( .A(n8721), .B(n8722), .Z(n8533) );
  XOR U8432 ( .A(n8723), .B(n8724), .Z(n8714) );
  AND U8433 ( .A(n8725), .B(n8726), .Z(n8724) );
  XOR U8434 ( .A(n8723), .B(n8548), .Z(n8726) );
  XOR U8435 ( .A(n8727), .B(n8728), .Z(n8548) );
  AND U8436 ( .A(n763), .B(n8729), .Z(n8728) );
  XOR U8437 ( .A(n8730), .B(n8727), .Z(n8729) );
  XNOR U8438 ( .A(n8545), .B(n8723), .Z(n8725) );
  XOR U8439 ( .A(n8731), .B(n8732), .Z(n8545) );
  AND U8440 ( .A(n761), .B(n8733), .Z(n8732) );
  XOR U8441 ( .A(n8734), .B(n8731), .Z(n8733) );
  XOR U8442 ( .A(n8735), .B(n8736), .Z(n8723) );
  AND U8443 ( .A(n8737), .B(n8738), .Z(n8736) );
  XOR U8444 ( .A(n8735), .B(n8560), .Z(n8738) );
  XOR U8445 ( .A(n8739), .B(n8740), .Z(n8560) );
  AND U8446 ( .A(n763), .B(n8741), .Z(n8740) );
  XOR U8447 ( .A(n8742), .B(n8739), .Z(n8741) );
  XNOR U8448 ( .A(n8557), .B(n8735), .Z(n8737) );
  XOR U8449 ( .A(n8743), .B(n8744), .Z(n8557) );
  AND U8450 ( .A(n761), .B(n8745), .Z(n8744) );
  XOR U8451 ( .A(n8746), .B(n8743), .Z(n8745) );
  XOR U8452 ( .A(n8747), .B(n8748), .Z(n8735) );
  AND U8453 ( .A(n8749), .B(n8750), .Z(n8748) );
  XOR U8454 ( .A(n8747), .B(n8572), .Z(n8750) );
  XOR U8455 ( .A(n8751), .B(n8752), .Z(n8572) );
  AND U8456 ( .A(n763), .B(n8753), .Z(n8752) );
  XOR U8457 ( .A(n8754), .B(n8751), .Z(n8753) );
  XNOR U8458 ( .A(n8569), .B(n8747), .Z(n8749) );
  XOR U8459 ( .A(n8755), .B(n8756), .Z(n8569) );
  AND U8460 ( .A(n761), .B(n8757), .Z(n8756) );
  XOR U8461 ( .A(n8758), .B(n8755), .Z(n8757) );
  XOR U8462 ( .A(n8759), .B(n8760), .Z(n8747) );
  AND U8463 ( .A(n8761), .B(n8762), .Z(n8760) );
  XOR U8464 ( .A(n8759), .B(n8584), .Z(n8762) );
  XOR U8465 ( .A(n8763), .B(n8764), .Z(n8584) );
  AND U8466 ( .A(n763), .B(n8765), .Z(n8764) );
  XOR U8467 ( .A(n8766), .B(n8763), .Z(n8765) );
  XNOR U8468 ( .A(n8581), .B(n8759), .Z(n8761) );
  XOR U8469 ( .A(n8767), .B(n8768), .Z(n8581) );
  AND U8470 ( .A(n761), .B(n8769), .Z(n8768) );
  XOR U8471 ( .A(n8770), .B(n8767), .Z(n8769) );
  XOR U8472 ( .A(n8771), .B(n8772), .Z(n8759) );
  AND U8473 ( .A(n8773), .B(n8774), .Z(n8772) );
  XOR U8474 ( .A(n8771), .B(n8596), .Z(n8774) );
  XOR U8475 ( .A(n8775), .B(n8776), .Z(n8596) );
  AND U8476 ( .A(n763), .B(n8777), .Z(n8776) );
  XOR U8477 ( .A(n8778), .B(n8775), .Z(n8777) );
  XNOR U8478 ( .A(n8593), .B(n8771), .Z(n8773) );
  XOR U8479 ( .A(n8779), .B(n8780), .Z(n8593) );
  AND U8480 ( .A(n761), .B(n8781), .Z(n8780) );
  XOR U8481 ( .A(n8782), .B(n8779), .Z(n8781) );
  XOR U8482 ( .A(n8783), .B(n8784), .Z(n8771) );
  AND U8483 ( .A(n8785), .B(n8786), .Z(n8784) );
  XOR U8484 ( .A(n8783), .B(n8608), .Z(n8786) );
  XOR U8485 ( .A(n8787), .B(n8788), .Z(n8608) );
  AND U8486 ( .A(n763), .B(n8789), .Z(n8788) );
  XOR U8487 ( .A(n8790), .B(n8787), .Z(n8789) );
  XNOR U8488 ( .A(n8605), .B(n8783), .Z(n8785) );
  XOR U8489 ( .A(n8791), .B(n8792), .Z(n8605) );
  AND U8490 ( .A(n761), .B(n8793), .Z(n8792) );
  XOR U8491 ( .A(n8794), .B(n8791), .Z(n8793) );
  XOR U8492 ( .A(n8795), .B(n8796), .Z(n8783) );
  AND U8493 ( .A(n8797), .B(n8798), .Z(n8796) );
  XOR U8494 ( .A(n8795), .B(n8620), .Z(n8798) );
  XOR U8495 ( .A(n8799), .B(n8800), .Z(n8620) );
  AND U8496 ( .A(n763), .B(n8801), .Z(n8800) );
  XOR U8497 ( .A(n8802), .B(n8799), .Z(n8801) );
  XNOR U8498 ( .A(n8617), .B(n8795), .Z(n8797) );
  XOR U8499 ( .A(n8803), .B(n8804), .Z(n8617) );
  AND U8500 ( .A(n761), .B(n8805), .Z(n8804) );
  XOR U8501 ( .A(n8806), .B(n8803), .Z(n8805) );
  XOR U8502 ( .A(n8807), .B(n8808), .Z(n8795) );
  AND U8503 ( .A(n8809), .B(n8810), .Z(n8808) );
  XOR U8504 ( .A(n8807), .B(n8632), .Z(n8810) );
  XOR U8505 ( .A(n8811), .B(n8812), .Z(n8632) );
  AND U8506 ( .A(n763), .B(n8813), .Z(n8812) );
  XOR U8507 ( .A(n8814), .B(n8811), .Z(n8813) );
  XNOR U8508 ( .A(n8629), .B(n8807), .Z(n8809) );
  XOR U8509 ( .A(n8815), .B(n8816), .Z(n8629) );
  AND U8510 ( .A(n761), .B(n8817), .Z(n8816) );
  XOR U8511 ( .A(n8818), .B(n8815), .Z(n8817) );
  XOR U8512 ( .A(n8819), .B(n8820), .Z(n8807) );
  AND U8513 ( .A(n8821), .B(n8822), .Z(n8820) );
  XOR U8514 ( .A(n8819), .B(n8644), .Z(n8822) );
  XOR U8515 ( .A(n8823), .B(n8824), .Z(n8644) );
  AND U8516 ( .A(n763), .B(n8825), .Z(n8824) );
  XOR U8517 ( .A(n8826), .B(n8823), .Z(n8825) );
  XNOR U8518 ( .A(n8641), .B(n8819), .Z(n8821) );
  XOR U8519 ( .A(n8827), .B(n8828), .Z(n8641) );
  AND U8520 ( .A(n761), .B(n8829), .Z(n8828) );
  XOR U8521 ( .A(n8830), .B(n8827), .Z(n8829) );
  XOR U8522 ( .A(n8831), .B(n8832), .Z(n8819) );
  AND U8523 ( .A(n8833), .B(n8834), .Z(n8832) );
  XOR U8524 ( .A(n8831), .B(n8656), .Z(n8834) );
  XOR U8525 ( .A(n8835), .B(n8836), .Z(n8656) );
  AND U8526 ( .A(n763), .B(n8837), .Z(n8836) );
  XOR U8527 ( .A(n8838), .B(n8835), .Z(n8837) );
  XNOR U8528 ( .A(n8653), .B(n8831), .Z(n8833) );
  XOR U8529 ( .A(n8839), .B(n8840), .Z(n8653) );
  AND U8530 ( .A(n761), .B(n8841), .Z(n8840) );
  XOR U8531 ( .A(n8842), .B(n8839), .Z(n8841) );
  XOR U8532 ( .A(n8843), .B(n8844), .Z(n8831) );
  AND U8533 ( .A(n8845), .B(n8846), .Z(n8844) );
  XOR U8534 ( .A(n8843), .B(n8668), .Z(n8846) );
  XOR U8535 ( .A(n8847), .B(n8848), .Z(n8668) );
  AND U8536 ( .A(n763), .B(n8849), .Z(n8848) );
  XOR U8537 ( .A(n8850), .B(n8847), .Z(n8849) );
  XNOR U8538 ( .A(n8665), .B(n8843), .Z(n8845) );
  XOR U8539 ( .A(n8851), .B(n8852), .Z(n8665) );
  AND U8540 ( .A(n761), .B(n8853), .Z(n8852) );
  XOR U8541 ( .A(n8854), .B(n8851), .Z(n8853) );
  XOR U8542 ( .A(n8855), .B(n8856), .Z(n8843) );
  AND U8543 ( .A(n8857), .B(n8858), .Z(n8856) );
  XOR U8544 ( .A(n8855), .B(n8680), .Z(n8858) );
  XOR U8545 ( .A(n8859), .B(n8860), .Z(n8680) );
  AND U8546 ( .A(n763), .B(n8861), .Z(n8860) );
  XOR U8547 ( .A(n8862), .B(n8859), .Z(n8861) );
  XNOR U8548 ( .A(n8677), .B(n8855), .Z(n8857) );
  XOR U8549 ( .A(n8863), .B(n8864), .Z(n8677) );
  AND U8550 ( .A(n761), .B(n8865), .Z(n8864) );
  XOR U8551 ( .A(n8866), .B(n8863), .Z(n8865) );
  XOR U8552 ( .A(n8867), .B(n8868), .Z(n8855) );
  AND U8553 ( .A(n8869), .B(n8870), .Z(n8868) );
  XOR U8554 ( .A(n8867), .B(n8692), .Z(n8870) );
  XOR U8555 ( .A(n8871), .B(n8872), .Z(n8692) );
  AND U8556 ( .A(n763), .B(n8873), .Z(n8872) );
  XOR U8557 ( .A(n8874), .B(n8871), .Z(n8873) );
  XNOR U8558 ( .A(n8689), .B(n8867), .Z(n8869) );
  XOR U8559 ( .A(n8875), .B(n8876), .Z(n8689) );
  AND U8560 ( .A(n761), .B(n8877), .Z(n8876) );
  XOR U8561 ( .A(n8878), .B(n8875), .Z(n8877) );
  XOR U8562 ( .A(n8879), .B(n8880), .Z(n8867) );
  AND U8563 ( .A(n8881), .B(n8882), .Z(n8880) );
  XNOR U8564 ( .A(n8883), .B(n8705), .Z(n8882) );
  XOR U8565 ( .A(n8884), .B(n8885), .Z(n8705) );
  AND U8566 ( .A(n763), .B(n8886), .Z(n8885) );
  XOR U8567 ( .A(n8884), .B(n8887), .Z(n8886) );
  XNOR U8568 ( .A(n8702), .B(n8879), .Z(n8881) );
  XOR U8569 ( .A(n8888), .B(n8889), .Z(n8702) );
  AND U8570 ( .A(n761), .B(n8890), .Z(n8889) );
  XOR U8571 ( .A(n8888), .B(n8891), .Z(n8890) );
  IV U8572 ( .A(n8883), .Z(n8879) );
  AND U8573 ( .A(n8710), .B(n8713), .Z(n8883) );
  XNOR U8574 ( .A(n8892), .B(n8893), .Z(n8713) );
  AND U8575 ( .A(n763), .B(n8894), .Z(n8893) );
  XNOR U8576 ( .A(n8895), .B(n8892), .Z(n8894) );
  XOR U8577 ( .A(n8896), .B(n8897), .Z(n763) );
  AND U8578 ( .A(n8898), .B(n8899), .Z(n8897) );
  XNOR U8579 ( .A(n8719), .B(n8896), .Z(n8899) );
  AND U8580 ( .A(n8900), .B(n8901), .Z(n8719) );
  XOR U8581 ( .A(n8896), .B(n8720), .Z(n8898) );
  AND U8582 ( .A(n8902), .B(n8903), .Z(n8720) );
  XOR U8583 ( .A(n8904), .B(n8905), .Z(n8896) );
  AND U8584 ( .A(n8906), .B(n8907), .Z(n8905) );
  XOR U8585 ( .A(n8904), .B(n8730), .Z(n8907) );
  XOR U8586 ( .A(n8908), .B(n8909), .Z(n8730) );
  AND U8587 ( .A(n419), .B(n8910), .Z(n8909) );
  XOR U8588 ( .A(n8911), .B(n8908), .Z(n8910) );
  XNOR U8589 ( .A(n8727), .B(n8904), .Z(n8906) );
  XOR U8590 ( .A(n8912), .B(n8913), .Z(n8727) );
  AND U8591 ( .A(n417), .B(n8914), .Z(n8913) );
  XOR U8592 ( .A(n8915), .B(n8912), .Z(n8914) );
  XOR U8593 ( .A(n8916), .B(n8917), .Z(n8904) );
  AND U8594 ( .A(n8918), .B(n8919), .Z(n8917) );
  XOR U8595 ( .A(n8916), .B(n8742), .Z(n8919) );
  XOR U8596 ( .A(n8920), .B(n8921), .Z(n8742) );
  AND U8597 ( .A(n419), .B(n8922), .Z(n8921) );
  XOR U8598 ( .A(n8923), .B(n8920), .Z(n8922) );
  XNOR U8599 ( .A(n8739), .B(n8916), .Z(n8918) );
  XOR U8600 ( .A(n8924), .B(n8925), .Z(n8739) );
  AND U8601 ( .A(n417), .B(n8926), .Z(n8925) );
  XOR U8602 ( .A(n8927), .B(n8924), .Z(n8926) );
  XOR U8603 ( .A(n8928), .B(n8929), .Z(n8916) );
  AND U8604 ( .A(n8930), .B(n8931), .Z(n8929) );
  XOR U8605 ( .A(n8928), .B(n8754), .Z(n8931) );
  XOR U8606 ( .A(n8932), .B(n8933), .Z(n8754) );
  AND U8607 ( .A(n419), .B(n8934), .Z(n8933) );
  XOR U8608 ( .A(n8935), .B(n8932), .Z(n8934) );
  XNOR U8609 ( .A(n8751), .B(n8928), .Z(n8930) );
  XOR U8610 ( .A(n8936), .B(n8937), .Z(n8751) );
  AND U8611 ( .A(n417), .B(n8938), .Z(n8937) );
  XOR U8612 ( .A(n8939), .B(n8936), .Z(n8938) );
  XOR U8613 ( .A(n8940), .B(n8941), .Z(n8928) );
  AND U8614 ( .A(n8942), .B(n8943), .Z(n8941) );
  XOR U8615 ( .A(n8940), .B(n8766), .Z(n8943) );
  XOR U8616 ( .A(n8944), .B(n8945), .Z(n8766) );
  AND U8617 ( .A(n419), .B(n8946), .Z(n8945) );
  XOR U8618 ( .A(n8947), .B(n8944), .Z(n8946) );
  XNOR U8619 ( .A(n8763), .B(n8940), .Z(n8942) );
  XOR U8620 ( .A(n8948), .B(n8949), .Z(n8763) );
  AND U8621 ( .A(n417), .B(n8950), .Z(n8949) );
  XOR U8622 ( .A(n8951), .B(n8948), .Z(n8950) );
  XOR U8623 ( .A(n8952), .B(n8953), .Z(n8940) );
  AND U8624 ( .A(n8954), .B(n8955), .Z(n8953) );
  XOR U8625 ( .A(n8952), .B(n8778), .Z(n8955) );
  XOR U8626 ( .A(n8956), .B(n8957), .Z(n8778) );
  AND U8627 ( .A(n419), .B(n8958), .Z(n8957) );
  XOR U8628 ( .A(n8959), .B(n8956), .Z(n8958) );
  XNOR U8629 ( .A(n8775), .B(n8952), .Z(n8954) );
  XOR U8630 ( .A(n8960), .B(n8961), .Z(n8775) );
  AND U8631 ( .A(n417), .B(n8962), .Z(n8961) );
  XOR U8632 ( .A(n8963), .B(n8960), .Z(n8962) );
  XOR U8633 ( .A(n8964), .B(n8965), .Z(n8952) );
  AND U8634 ( .A(n8966), .B(n8967), .Z(n8965) );
  XOR U8635 ( .A(n8964), .B(n8790), .Z(n8967) );
  XOR U8636 ( .A(n8968), .B(n8969), .Z(n8790) );
  AND U8637 ( .A(n419), .B(n8970), .Z(n8969) );
  XOR U8638 ( .A(n8971), .B(n8968), .Z(n8970) );
  XNOR U8639 ( .A(n8787), .B(n8964), .Z(n8966) );
  XOR U8640 ( .A(n8972), .B(n8973), .Z(n8787) );
  AND U8641 ( .A(n417), .B(n8974), .Z(n8973) );
  XOR U8642 ( .A(n8975), .B(n8972), .Z(n8974) );
  XOR U8643 ( .A(n8976), .B(n8977), .Z(n8964) );
  AND U8644 ( .A(n8978), .B(n8979), .Z(n8977) );
  XOR U8645 ( .A(n8976), .B(n8802), .Z(n8979) );
  XOR U8646 ( .A(n8980), .B(n8981), .Z(n8802) );
  AND U8647 ( .A(n419), .B(n8982), .Z(n8981) );
  XOR U8648 ( .A(n8983), .B(n8980), .Z(n8982) );
  XNOR U8649 ( .A(n8799), .B(n8976), .Z(n8978) );
  XOR U8650 ( .A(n8984), .B(n8985), .Z(n8799) );
  AND U8651 ( .A(n417), .B(n8986), .Z(n8985) );
  XOR U8652 ( .A(n8987), .B(n8984), .Z(n8986) );
  XOR U8653 ( .A(n8988), .B(n8989), .Z(n8976) );
  AND U8654 ( .A(n8990), .B(n8991), .Z(n8989) );
  XOR U8655 ( .A(n8988), .B(n8814), .Z(n8991) );
  XOR U8656 ( .A(n8992), .B(n8993), .Z(n8814) );
  AND U8657 ( .A(n419), .B(n8994), .Z(n8993) );
  XOR U8658 ( .A(n8995), .B(n8992), .Z(n8994) );
  XNOR U8659 ( .A(n8811), .B(n8988), .Z(n8990) );
  XOR U8660 ( .A(n8996), .B(n8997), .Z(n8811) );
  AND U8661 ( .A(n417), .B(n8998), .Z(n8997) );
  XOR U8662 ( .A(n8999), .B(n8996), .Z(n8998) );
  XOR U8663 ( .A(n9000), .B(n9001), .Z(n8988) );
  AND U8664 ( .A(n9002), .B(n9003), .Z(n9001) );
  XOR U8665 ( .A(n9000), .B(n8826), .Z(n9003) );
  XOR U8666 ( .A(n9004), .B(n9005), .Z(n8826) );
  AND U8667 ( .A(n419), .B(n9006), .Z(n9005) );
  XOR U8668 ( .A(n9007), .B(n9004), .Z(n9006) );
  XNOR U8669 ( .A(n8823), .B(n9000), .Z(n9002) );
  XOR U8670 ( .A(n9008), .B(n9009), .Z(n8823) );
  AND U8671 ( .A(n417), .B(n9010), .Z(n9009) );
  XOR U8672 ( .A(n9011), .B(n9008), .Z(n9010) );
  XOR U8673 ( .A(n9012), .B(n9013), .Z(n9000) );
  AND U8674 ( .A(n9014), .B(n9015), .Z(n9013) );
  XOR U8675 ( .A(n9012), .B(n8838), .Z(n9015) );
  XOR U8676 ( .A(n9016), .B(n9017), .Z(n8838) );
  AND U8677 ( .A(n419), .B(n9018), .Z(n9017) );
  XOR U8678 ( .A(n9019), .B(n9016), .Z(n9018) );
  XNOR U8679 ( .A(n8835), .B(n9012), .Z(n9014) );
  XOR U8680 ( .A(n9020), .B(n9021), .Z(n8835) );
  AND U8681 ( .A(n417), .B(n9022), .Z(n9021) );
  XOR U8682 ( .A(n9023), .B(n9020), .Z(n9022) );
  XOR U8683 ( .A(n9024), .B(n9025), .Z(n9012) );
  AND U8684 ( .A(n9026), .B(n9027), .Z(n9025) );
  XOR U8685 ( .A(n9024), .B(n8850), .Z(n9027) );
  XOR U8686 ( .A(n9028), .B(n9029), .Z(n8850) );
  AND U8687 ( .A(n419), .B(n9030), .Z(n9029) );
  XOR U8688 ( .A(n9031), .B(n9028), .Z(n9030) );
  XNOR U8689 ( .A(n8847), .B(n9024), .Z(n9026) );
  XOR U8690 ( .A(n9032), .B(n9033), .Z(n8847) );
  AND U8691 ( .A(n417), .B(n9034), .Z(n9033) );
  XOR U8692 ( .A(n9035), .B(n9032), .Z(n9034) );
  XOR U8693 ( .A(n9036), .B(n9037), .Z(n9024) );
  AND U8694 ( .A(n9038), .B(n9039), .Z(n9037) );
  XOR U8695 ( .A(n9036), .B(n8862), .Z(n9039) );
  XOR U8696 ( .A(n9040), .B(n9041), .Z(n8862) );
  AND U8697 ( .A(n419), .B(n9042), .Z(n9041) );
  XOR U8698 ( .A(n9043), .B(n9040), .Z(n9042) );
  XNOR U8699 ( .A(n8859), .B(n9036), .Z(n9038) );
  XOR U8700 ( .A(n9044), .B(n9045), .Z(n8859) );
  AND U8701 ( .A(n417), .B(n9046), .Z(n9045) );
  XOR U8702 ( .A(n9047), .B(n9044), .Z(n9046) );
  XOR U8703 ( .A(n9048), .B(n9049), .Z(n9036) );
  AND U8704 ( .A(n9050), .B(n9051), .Z(n9049) );
  XOR U8705 ( .A(n9048), .B(n8874), .Z(n9051) );
  XOR U8706 ( .A(n9052), .B(n9053), .Z(n8874) );
  AND U8707 ( .A(n419), .B(n9054), .Z(n9053) );
  XOR U8708 ( .A(n9055), .B(n9052), .Z(n9054) );
  XNOR U8709 ( .A(n8871), .B(n9048), .Z(n9050) );
  XOR U8710 ( .A(n9056), .B(n9057), .Z(n8871) );
  AND U8711 ( .A(n417), .B(n9058), .Z(n9057) );
  XOR U8712 ( .A(n9059), .B(n9056), .Z(n9058) );
  XOR U8713 ( .A(n9060), .B(n9061), .Z(n9048) );
  AND U8714 ( .A(n9062), .B(n9063), .Z(n9061) );
  XNOR U8715 ( .A(n9064), .B(n8887), .Z(n9063) );
  XOR U8716 ( .A(n9065), .B(n9066), .Z(n8887) );
  AND U8717 ( .A(n419), .B(n9067), .Z(n9066) );
  XOR U8718 ( .A(n9065), .B(n9068), .Z(n9067) );
  XNOR U8719 ( .A(n8884), .B(n9060), .Z(n9062) );
  XOR U8720 ( .A(n9069), .B(n9070), .Z(n8884) );
  AND U8721 ( .A(n417), .B(n9071), .Z(n9070) );
  XOR U8722 ( .A(n9069), .B(n9072), .Z(n9071) );
  IV U8723 ( .A(n9064), .Z(n9060) );
  AND U8724 ( .A(n8892), .B(n8895), .Z(n9064) );
  XNOR U8725 ( .A(n9073), .B(n9074), .Z(n8895) );
  AND U8726 ( .A(n419), .B(n9075), .Z(n9074) );
  XNOR U8727 ( .A(n9076), .B(n9073), .Z(n9075) );
  XOR U8728 ( .A(n9077), .B(n9078), .Z(n419) );
  AND U8729 ( .A(n9079), .B(n9080), .Z(n9078) );
  XNOR U8730 ( .A(n8900), .B(n9077), .Z(n9080) );
  AND U8731 ( .A(p_input[3071]), .B(p_input[3055]), .Z(n8900) );
  XOR U8732 ( .A(n9077), .B(n8901), .Z(n9079) );
  AND U8733 ( .A(p_input[3039]), .B(p_input[3023]), .Z(n8901) );
  XOR U8734 ( .A(n9081), .B(n9082), .Z(n9077) );
  AND U8735 ( .A(n9083), .B(n9084), .Z(n9082) );
  XOR U8736 ( .A(n9081), .B(n8911), .Z(n9084) );
  XNOR U8737 ( .A(p_input[3054]), .B(n9085), .Z(n8911) );
  AND U8738 ( .A(n231), .B(n9086), .Z(n9085) );
  XOR U8739 ( .A(p_input[3070]), .B(p_input[3054]), .Z(n9086) );
  XNOR U8740 ( .A(n8908), .B(n9081), .Z(n9083) );
  XOR U8741 ( .A(n9087), .B(n9088), .Z(n8908) );
  AND U8742 ( .A(n229), .B(n9089), .Z(n9088) );
  XOR U8743 ( .A(p_input[3038]), .B(p_input[3022]), .Z(n9089) );
  XOR U8744 ( .A(n9090), .B(n9091), .Z(n9081) );
  AND U8745 ( .A(n9092), .B(n9093), .Z(n9091) );
  XOR U8746 ( .A(n9090), .B(n8923), .Z(n9093) );
  XNOR U8747 ( .A(p_input[3053]), .B(n9094), .Z(n8923) );
  AND U8748 ( .A(n231), .B(n9095), .Z(n9094) );
  XOR U8749 ( .A(p_input[3069]), .B(p_input[3053]), .Z(n9095) );
  XNOR U8750 ( .A(n8920), .B(n9090), .Z(n9092) );
  XOR U8751 ( .A(n9096), .B(n9097), .Z(n8920) );
  AND U8752 ( .A(n229), .B(n9098), .Z(n9097) );
  XOR U8753 ( .A(p_input[3037]), .B(p_input[3021]), .Z(n9098) );
  XOR U8754 ( .A(n9099), .B(n9100), .Z(n9090) );
  AND U8755 ( .A(n9101), .B(n9102), .Z(n9100) );
  XOR U8756 ( .A(n9099), .B(n8935), .Z(n9102) );
  XNOR U8757 ( .A(p_input[3052]), .B(n9103), .Z(n8935) );
  AND U8758 ( .A(n231), .B(n9104), .Z(n9103) );
  XOR U8759 ( .A(p_input[3068]), .B(p_input[3052]), .Z(n9104) );
  XNOR U8760 ( .A(n8932), .B(n9099), .Z(n9101) );
  XOR U8761 ( .A(n9105), .B(n9106), .Z(n8932) );
  AND U8762 ( .A(n229), .B(n9107), .Z(n9106) );
  XOR U8763 ( .A(p_input[3036]), .B(p_input[3020]), .Z(n9107) );
  XOR U8764 ( .A(n9108), .B(n9109), .Z(n9099) );
  AND U8765 ( .A(n9110), .B(n9111), .Z(n9109) );
  XOR U8766 ( .A(n9108), .B(n8947), .Z(n9111) );
  XNOR U8767 ( .A(p_input[3051]), .B(n9112), .Z(n8947) );
  AND U8768 ( .A(n231), .B(n9113), .Z(n9112) );
  XOR U8769 ( .A(p_input[3067]), .B(p_input[3051]), .Z(n9113) );
  XNOR U8770 ( .A(n8944), .B(n9108), .Z(n9110) );
  XOR U8771 ( .A(n9114), .B(n9115), .Z(n8944) );
  AND U8772 ( .A(n229), .B(n9116), .Z(n9115) );
  XOR U8773 ( .A(p_input[3035]), .B(p_input[3019]), .Z(n9116) );
  XOR U8774 ( .A(n9117), .B(n9118), .Z(n9108) );
  AND U8775 ( .A(n9119), .B(n9120), .Z(n9118) );
  XOR U8776 ( .A(n9117), .B(n8959), .Z(n9120) );
  XNOR U8777 ( .A(p_input[3050]), .B(n9121), .Z(n8959) );
  AND U8778 ( .A(n231), .B(n9122), .Z(n9121) );
  XOR U8779 ( .A(p_input[3066]), .B(p_input[3050]), .Z(n9122) );
  XNOR U8780 ( .A(n8956), .B(n9117), .Z(n9119) );
  XOR U8781 ( .A(n9123), .B(n9124), .Z(n8956) );
  AND U8782 ( .A(n229), .B(n9125), .Z(n9124) );
  XOR U8783 ( .A(p_input[3034]), .B(p_input[3018]), .Z(n9125) );
  XOR U8784 ( .A(n9126), .B(n9127), .Z(n9117) );
  AND U8785 ( .A(n9128), .B(n9129), .Z(n9127) );
  XOR U8786 ( .A(n9126), .B(n8971), .Z(n9129) );
  XNOR U8787 ( .A(p_input[3049]), .B(n9130), .Z(n8971) );
  AND U8788 ( .A(n231), .B(n9131), .Z(n9130) );
  XOR U8789 ( .A(p_input[3065]), .B(p_input[3049]), .Z(n9131) );
  XNOR U8790 ( .A(n8968), .B(n9126), .Z(n9128) );
  XOR U8791 ( .A(n9132), .B(n9133), .Z(n8968) );
  AND U8792 ( .A(n229), .B(n9134), .Z(n9133) );
  XOR U8793 ( .A(p_input[3033]), .B(p_input[3017]), .Z(n9134) );
  XOR U8794 ( .A(n9135), .B(n9136), .Z(n9126) );
  AND U8795 ( .A(n9137), .B(n9138), .Z(n9136) );
  XOR U8796 ( .A(n9135), .B(n8983), .Z(n9138) );
  XNOR U8797 ( .A(p_input[3048]), .B(n9139), .Z(n8983) );
  AND U8798 ( .A(n231), .B(n9140), .Z(n9139) );
  XOR U8799 ( .A(p_input[3064]), .B(p_input[3048]), .Z(n9140) );
  XNOR U8800 ( .A(n8980), .B(n9135), .Z(n9137) );
  XOR U8801 ( .A(n9141), .B(n9142), .Z(n8980) );
  AND U8802 ( .A(n229), .B(n9143), .Z(n9142) );
  XOR U8803 ( .A(p_input[3032]), .B(p_input[3016]), .Z(n9143) );
  XOR U8804 ( .A(n9144), .B(n9145), .Z(n9135) );
  AND U8805 ( .A(n9146), .B(n9147), .Z(n9145) );
  XOR U8806 ( .A(n9144), .B(n8995), .Z(n9147) );
  XNOR U8807 ( .A(p_input[3047]), .B(n9148), .Z(n8995) );
  AND U8808 ( .A(n231), .B(n9149), .Z(n9148) );
  XOR U8809 ( .A(p_input[3063]), .B(p_input[3047]), .Z(n9149) );
  XNOR U8810 ( .A(n8992), .B(n9144), .Z(n9146) );
  XOR U8811 ( .A(n9150), .B(n9151), .Z(n8992) );
  AND U8812 ( .A(n229), .B(n9152), .Z(n9151) );
  XOR U8813 ( .A(p_input[3031]), .B(p_input[3015]), .Z(n9152) );
  XOR U8814 ( .A(n9153), .B(n9154), .Z(n9144) );
  AND U8815 ( .A(n9155), .B(n9156), .Z(n9154) );
  XOR U8816 ( .A(n9153), .B(n9007), .Z(n9156) );
  XNOR U8817 ( .A(p_input[3046]), .B(n9157), .Z(n9007) );
  AND U8818 ( .A(n231), .B(n9158), .Z(n9157) );
  XOR U8819 ( .A(p_input[3062]), .B(p_input[3046]), .Z(n9158) );
  XNOR U8820 ( .A(n9004), .B(n9153), .Z(n9155) );
  XOR U8821 ( .A(n9159), .B(n9160), .Z(n9004) );
  AND U8822 ( .A(n229), .B(n9161), .Z(n9160) );
  XOR U8823 ( .A(p_input[3030]), .B(p_input[3014]), .Z(n9161) );
  XOR U8824 ( .A(n9162), .B(n9163), .Z(n9153) );
  AND U8825 ( .A(n9164), .B(n9165), .Z(n9163) );
  XOR U8826 ( .A(n9162), .B(n9019), .Z(n9165) );
  XNOR U8827 ( .A(p_input[3045]), .B(n9166), .Z(n9019) );
  AND U8828 ( .A(n231), .B(n9167), .Z(n9166) );
  XOR U8829 ( .A(p_input[3061]), .B(p_input[3045]), .Z(n9167) );
  XNOR U8830 ( .A(n9016), .B(n9162), .Z(n9164) );
  XOR U8831 ( .A(n9168), .B(n9169), .Z(n9016) );
  AND U8832 ( .A(n229), .B(n9170), .Z(n9169) );
  XOR U8833 ( .A(p_input[3029]), .B(p_input[3013]), .Z(n9170) );
  XOR U8834 ( .A(n9171), .B(n9172), .Z(n9162) );
  AND U8835 ( .A(n9173), .B(n9174), .Z(n9172) );
  XOR U8836 ( .A(n9171), .B(n9031), .Z(n9174) );
  XNOR U8837 ( .A(p_input[3044]), .B(n9175), .Z(n9031) );
  AND U8838 ( .A(n231), .B(n9176), .Z(n9175) );
  XOR U8839 ( .A(p_input[3060]), .B(p_input[3044]), .Z(n9176) );
  XNOR U8840 ( .A(n9028), .B(n9171), .Z(n9173) );
  XOR U8841 ( .A(n9177), .B(n9178), .Z(n9028) );
  AND U8842 ( .A(n229), .B(n9179), .Z(n9178) );
  XOR U8843 ( .A(p_input[3028]), .B(p_input[3012]), .Z(n9179) );
  XOR U8844 ( .A(n9180), .B(n9181), .Z(n9171) );
  AND U8845 ( .A(n9182), .B(n9183), .Z(n9181) );
  XOR U8846 ( .A(n9180), .B(n9043), .Z(n9183) );
  XNOR U8847 ( .A(p_input[3043]), .B(n9184), .Z(n9043) );
  AND U8848 ( .A(n231), .B(n9185), .Z(n9184) );
  XOR U8849 ( .A(p_input[3059]), .B(p_input[3043]), .Z(n9185) );
  XNOR U8850 ( .A(n9040), .B(n9180), .Z(n9182) );
  XOR U8851 ( .A(n9186), .B(n9187), .Z(n9040) );
  AND U8852 ( .A(n229), .B(n9188), .Z(n9187) );
  XOR U8853 ( .A(p_input[3027]), .B(p_input[3011]), .Z(n9188) );
  XOR U8854 ( .A(n9189), .B(n9190), .Z(n9180) );
  AND U8855 ( .A(n9191), .B(n9192), .Z(n9190) );
  XOR U8856 ( .A(n9189), .B(n9055), .Z(n9192) );
  XNOR U8857 ( .A(p_input[3042]), .B(n9193), .Z(n9055) );
  AND U8858 ( .A(n231), .B(n9194), .Z(n9193) );
  XOR U8859 ( .A(p_input[3058]), .B(p_input[3042]), .Z(n9194) );
  XNOR U8860 ( .A(n9052), .B(n9189), .Z(n9191) );
  XOR U8861 ( .A(n9195), .B(n9196), .Z(n9052) );
  AND U8862 ( .A(n229), .B(n9197), .Z(n9196) );
  XOR U8863 ( .A(p_input[3026]), .B(p_input[3010]), .Z(n9197) );
  XOR U8864 ( .A(n9198), .B(n9199), .Z(n9189) );
  AND U8865 ( .A(n9200), .B(n9201), .Z(n9199) );
  XNOR U8866 ( .A(n9202), .B(n9068), .Z(n9201) );
  XNOR U8867 ( .A(p_input[3041]), .B(n9203), .Z(n9068) );
  AND U8868 ( .A(n231), .B(n9204), .Z(n9203) );
  XNOR U8869 ( .A(p_input[3057]), .B(n9205), .Z(n9204) );
  IV U8870 ( .A(p_input[3041]), .Z(n9205) );
  XNOR U8871 ( .A(n9065), .B(n9198), .Z(n9200) );
  XNOR U8872 ( .A(p_input[3009]), .B(n9206), .Z(n9065) );
  AND U8873 ( .A(n229), .B(n9207), .Z(n9206) );
  XOR U8874 ( .A(p_input[3025]), .B(p_input[3009]), .Z(n9207) );
  IV U8875 ( .A(n9202), .Z(n9198) );
  AND U8876 ( .A(n9073), .B(n9076), .Z(n9202) );
  XOR U8877 ( .A(p_input[3040]), .B(n9208), .Z(n9076) );
  AND U8878 ( .A(n231), .B(n9209), .Z(n9208) );
  XOR U8879 ( .A(p_input[3056]), .B(p_input[3040]), .Z(n9209) );
  XOR U8880 ( .A(n9210), .B(n9211), .Z(n231) );
  AND U8881 ( .A(n9212), .B(n9213), .Z(n9211) );
  XNOR U8882 ( .A(p_input[3071]), .B(n9210), .Z(n9213) );
  XOR U8883 ( .A(n9210), .B(p_input[3055]), .Z(n9212) );
  XOR U8884 ( .A(n9214), .B(n9215), .Z(n9210) );
  AND U8885 ( .A(n9216), .B(n9217), .Z(n9215) );
  XNOR U8886 ( .A(p_input[3070]), .B(n9214), .Z(n9217) );
  XOR U8887 ( .A(n9214), .B(p_input[3054]), .Z(n9216) );
  XOR U8888 ( .A(n9218), .B(n9219), .Z(n9214) );
  AND U8889 ( .A(n9220), .B(n9221), .Z(n9219) );
  XNOR U8890 ( .A(p_input[3069]), .B(n9218), .Z(n9221) );
  XOR U8891 ( .A(n9218), .B(p_input[3053]), .Z(n9220) );
  XOR U8892 ( .A(n9222), .B(n9223), .Z(n9218) );
  AND U8893 ( .A(n9224), .B(n9225), .Z(n9223) );
  XNOR U8894 ( .A(p_input[3068]), .B(n9222), .Z(n9225) );
  XOR U8895 ( .A(n9222), .B(p_input[3052]), .Z(n9224) );
  XOR U8896 ( .A(n9226), .B(n9227), .Z(n9222) );
  AND U8897 ( .A(n9228), .B(n9229), .Z(n9227) );
  XNOR U8898 ( .A(p_input[3067]), .B(n9226), .Z(n9229) );
  XOR U8899 ( .A(n9226), .B(p_input[3051]), .Z(n9228) );
  XOR U8900 ( .A(n9230), .B(n9231), .Z(n9226) );
  AND U8901 ( .A(n9232), .B(n9233), .Z(n9231) );
  XNOR U8902 ( .A(p_input[3066]), .B(n9230), .Z(n9233) );
  XOR U8903 ( .A(n9230), .B(p_input[3050]), .Z(n9232) );
  XOR U8904 ( .A(n9234), .B(n9235), .Z(n9230) );
  AND U8905 ( .A(n9236), .B(n9237), .Z(n9235) );
  XNOR U8906 ( .A(p_input[3065]), .B(n9234), .Z(n9237) );
  XOR U8907 ( .A(n9234), .B(p_input[3049]), .Z(n9236) );
  XOR U8908 ( .A(n9238), .B(n9239), .Z(n9234) );
  AND U8909 ( .A(n9240), .B(n9241), .Z(n9239) );
  XNOR U8910 ( .A(p_input[3064]), .B(n9238), .Z(n9241) );
  XOR U8911 ( .A(n9238), .B(p_input[3048]), .Z(n9240) );
  XOR U8912 ( .A(n9242), .B(n9243), .Z(n9238) );
  AND U8913 ( .A(n9244), .B(n9245), .Z(n9243) );
  XNOR U8914 ( .A(p_input[3063]), .B(n9242), .Z(n9245) );
  XOR U8915 ( .A(n9242), .B(p_input[3047]), .Z(n9244) );
  XOR U8916 ( .A(n9246), .B(n9247), .Z(n9242) );
  AND U8917 ( .A(n9248), .B(n9249), .Z(n9247) );
  XNOR U8918 ( .A(p_input[3062]), .B(n9246), .Z(n9249) );
  XOR U8919 ( .A(n9246), .B(p_input[3046]), .Z(n9248) );
  XOR U8920 ( .A(n9250), .B(n9251), .Z(n9246) );
  AND U8921 ( .A(n9252), .B(n9253), .Z(n9251) );
  XNOR U8922 ( .A(p_input[3061]), .B(n9250), .Z(n9253) );
  XOR U8923 ( .A(n9250), .B(p_input[3045]), .Z(n9252) );
  XOR U8924 ( .A(n9254), .B(n9255), .Z(n9250) );
  AND U8925 ( .A(n9256), .B(n9257), .Z(n9255) );
  XNOR U8926 ( .A(p_input[3060]), .B(n9254), .Z(n9257) );
  XOR U8927 ( .A(n9254), .B(p_input[3044]), .Z(n9256) );
  XOR U8928 ( .A(n9258), .B(n9259), .Z(n9254) );
  AND U8929 ( .A(n9260), .B(n9261), .Z(n9259) );
  XNOR U8930 ( .A(p_input[3059]), .B(n9258), .Z(n9261) );
  XOR U8931 ( .A(n9258), .B(p_input[3043]), .Z(n9260) );
  XOR U8932 ( .A(n9262), .B(n9263), .Z(n9258) );
  AND U8933 ( .A(n9264), .B(n9265), .Z(n9263) );
  XNOR U8934 ( .A(p_input[3058]), .B(n9262), .Z(n9265) );
  XOR U8935 ( .A(n9262), .B(p_input[3042]), .Z(n9264) );
  XNOR U8936 ( .A(n9266), .B(n9267), .Z(n9262) );
  AND U8937 ( .A(n9268), .B(n9269), .Z(n9267) );
  XOR U8938 ( .A(p_input[3057]), .B(n9266), .Z(n9269) );
  XNOR U8939 ( .A(p_input[3041]), .B(n9266), .Z(n9268) );
  AND U8940 ( .A(p_input[3056]), .B(n9270), .Z(n9266) );
  IV U8941 ( .A(p_input[3040]), .Z(n9270) );
  XNOR U8942 ( .A(p_input[3008]), .B(n9271), .Z(n9073) );
  AND U8943 ( .A(n229), .B(n9272), .Z(n9271) );
  XOR U8944 ( .A(p_input[3024]), .B(p_input[3008]), .Z(n9272) );
  XOR U8945 ( .A(n9273), .B(n9274), .Z(n229) );
  AND U8946 ( .A(n9275), .B(n9276), .Z(n9274) );
  XNOR U8947 ( .A(p_input[3039]), .B(n9273), .Z(n9276) );
  XOR U8948 ( .A(n9273), .B(p_input[3023]), .Z(n9275) );
  XOR U8949 ( .A(n9277), .B(n9278), .Z(n9273) );
  AND U8950 ( .A(n9279), .B(n9280), .Z(n9278) );
  XNOR U8951 ( .A(p_input[3038]), .B(n9277), .Z(n9280) );
  XNOR U8952 ( .A(n9277), .B(n9087), .Z(n9279) );
  IV U8953 ( .A(p_input[3022]), .Z(n9087) );
  XOR U8954 ( .A(n9281), .B(n9282), .Z(n9277) );
  AND U8955 ( .A(n9283), .B(n9284), .Z(n9282) );
  XNOR U8956 ( .A(p_input[3037]), .B(n9281), .Z(n9284) );
  XNOR U8957 ( .A(n9281), .B(n9096), .Z(n9283) );
  IV U8958 ( .A(p_input[3021]), .Z(n9096) );
  XOR U8959 ( .A(n9285), .B(n9286), .Z(n9281) );
  AND U8960 ( .A(n9287), .B(n9288), .Z(n9286) );
  XNOR U8961 ( .A(p_input[3036]), .B(n9285), .Z(n9288) );
  XNOR U8962 ( .A(n9285), .B(n9105), .Z(n9287) );
  IV U8963 ( .A(p_input[3020]), .Z(n9105) );
  XOR U8964 ( .A(n9289), .B(n9290), .Z(n9285) );
  AND U8965 ( .A(n9291), .B(n9292), .Z(n9290) );
  XNOR U8966 ( .A(p_input[3035]), .B(n9289), .Z(n9292) );
  XNOR U8967 ( .A(n9289), .B(n9114), .Z(n9291) );
  IV U8968 ( .A(p_input[3019]), .Z(n9114) );
  XOR U8969 ( .A(n9293), .B(n9294), .Z(n9289) );
  AND U8970 ( .A(n9295), .B(n9296), .Z(n9294) );
  XNOR U8971 ( .A(p_input[3034]), .B(n9293), .Z(n9296) );
  XNOR U8972 ( .A(n9293), .B(n9123), .Z(n9295) );
  IV U8973 ( .A(p_input[3018]), .Z(n9123) );
  XOR U8974 ( .A(n9297), .B(n9298), .Z(n9293) );
  AND U8975 ( .A(n9299), .B(n9300), .Z(n9298) );
  XNOR U8976 ( .A(p_input[3033]), .B(n9297), .Z(n9300) );
  XNOR U8977 ( .A(n9297), .B(n9132), .Z(n9299) );
  IV U8978 ( .A(p_input[3017]), .Z(n9132) );
  XOR U8979 ( .A(n9301), .B(n9302), .Z(n9297) );
  AND U8980 ( .A(n9303), .B(n9304), .Z(n9302) );
  XNOR U8981 ( .A(p_input[3032]), .B(n9301), .Z(n9304) );
  XNOR U8982 ( .A(n9301), .B(n9141), .Z(n9303) );
  IV U8983 ( .A(p_input[3016]), .Z(n9141) );
  XOR U8984 ( .A(n9305), .B(n9306), .Z(n9301) );
  AND U8985 ( .A(n9307), .B(n9308), .Z(n9306) );
  XNOR U8986 ( .A(p_input[3031]), .B(n9305), .Z(n9308) );
  XNOR U8987 ( .A(n9305), .B(n9150), .Z(n9307) );
  IV U8988 ( .A(p_input[3015]), .Z(n9150) );
  XOR U8989 ( .A(n9309), .B(n9310), .Z(n9305) );
  AND U8990 ( .A(n9311), .B(n9312), .Z(n9310) );
  XNOR U8991 ( .A(p_input[3030]), .B(n9309), .Z(n9312) );
  XNOR U8992 ( .A(n9309), .B(n9159), .Z(n9311) );
  IV U8993 ( .A(p_input[3014]), .Z(n9159) );
  XOR U8994 ( .A(n9313), .B(n9314), .Z(n9309) );
  AND U8995 ( .A(n9315), .B(n9316), .Z(n9314) );
  XNOR U8996 ( .A(p_input[3029]), .B(n9313), .Z(n9316) );
  XNOR U8997 ( .A(n9313), .B(n9168), .Z(n9315) );
  IV U8998 ( .A(p_input[3013]), .Z(n9168) );
  XOR U8999 ( .A(n9317), .B(n9318), .Z(n9313) );
  AND U9000 ( .A(n9319), .B(n9320), .Z(n9318) );
  XNOR U9001 ( .A(p_input[3028]), .B(n9317), .Z(n9320) );
  XNOR U9002 ( .A(n9317), .B(n9177), .Z(n9319) );
  IV U9003 ( .A(p_input[3012]), .Z(n9177) );
  XOR U9004 ( .A(n9321), .B(n9322), .Z(n9317) );
  AND U9005 ( .A(n9323), .B(n9324), .Z(n9322) );
  XNOR U9006 ( .A(p_input[3027]), .B(n9321), .Z(n9324) );
  XNOR U9007 ( .A(n9321), .B(n9186), .Z(n9323) );
  IV U9008 ( .A(p_input[3011]), .Z(n9186) );
  XOR U9009 ( .A(n9325), .B(n9326), .Z(n9321) );
  AND U9010 ( .A(n9327), .B(n9328), .Z(n9326) );
  XNOR U9011 ( .A(p_input[3026]), .B(n9325), .Z(n9328) );
  XNOR U9012 ( .A(n9325), .B(n9195), .Z(n9327) );
  IV U9013 ( .A(p_input[3010]), .Z(n9195) );
  XNOR U9014 ( .A(n9329), .B(n9330), .Z(n9325) );
  AND U9015 ( .A(n9331), .B(n9332), .Z(n9330) );
  XOR U9016 ( .A(p_input[3025]), .B(n9329), .Z(n9332) );
  XNOR U9017 ( .A(p_input[3009]), .B(n9329), .Z(n9331) );
  AND U9018 ( .A(p_input[3024]), .B(n9333), .Z(n9329) );
  IV U9019 ( .A(p_input[3008]), .Z(n9333) );
  XOR U9020 ( .A(n9334), .B(n9335), .Z(n8892) );
  AND U9021 ( .A(n417), .B(n9336), .Z(n9335) );
  XNOR U9022 ( .A(n9337), .B(n9334), .Z(n9336) );
  XOR U9023 ( .A(n9338), .B(n9339), .Z(n417) );
  AND U9024 ( .A(n9340), .B(n9341), .Z(n9339) );
  XNOR U9025 ( .A(n8902), .B(n9338), .Z(n9341) );
  AND U9026 ( .A(p_input[3007]), .B(p_input[2991]), .Z(n8902) );
  XOR U9027 ( .A(n9338), .B(n8903), .Z(n9340) );
  AND U9028 ( .A(p_input[2975]), .B(p_input[2959]), .Z(n8903) );
  XOR U9029 ( .A(n9342), .B(n9343), .Z(n9338) );
  AND U9030 ( .A(n9344), .B(n9345), .Z(n9343) );
  XOR U9031 ( .A(n9342), .B(n8915), .Z(n9345) );
  XNOR U9032 ( .A(p_input[2990]), .B(n9346), .Z(n8915) );
  AND U9033 ( .A(n235), .B(n9347), .Z(n9346) );
  XOR U9034 ( .A(p_input[3006]), .B(p_input[2990]), .Z(n9347) );
  XNOR U9035 ( .A(n8912), .B(n9342), .Z(n9344) );
  XOR U9036 ( .A(n9348), .B(n9349), .Z(n8912) );
  AND U9037 ( .A(n232), .B(n9350), .Z(n9349) );
  XOR U9038 ( .A(p_input[2974]), .B(p_input[2958]), .Z(n9350) );
  XOR U9039 ( .A(n9351), .B(n9352), .Z(n9342) );
  AND U9040 ( .A(n9353), .B(n9354), .Z(n9352) );
  XOR U9041 ( .A(n9351), .B(n8927), .Z(n9354) );
  XNOR U9042 ( .A(p_input[2989]), .B(n9355), .Z(n8927) );
  AND U9043 ( .A(n235), .B(n9356), .Z(n9355) );
  XOR U9044 ( .A(p_input[3005]), .B(p_input[2989]), .Z(n9356) );
  XNOR U9045 ( .A(n8924), .B(n9351), .Z(n9353) );
  XOR U9046 ( .A(n9357), .B(n9358), .Z(n8924) );
  AND U9047 ( .A(n232), .B(n9359), .Z(n9358) );
  XOR U9048 ( .A(p_input[2973]), .B(p_input[2957]), .Z(n9359) );
  XOR U9049 ( .A(n9360), .B(n9361), .Z(n9351) );
  AND U9050 ( .A(n9362), .B(n9363), .Z(n9361) );
  XOR U9051 ( .A(n9360), .B(n8939), .Z(n9363) );
  XNOR U9052 ( .A(p_input[2988]), .B(n9364), .Z(n8939) );
  AND U9053 ( .A(n235), .B(n9365), .Z(n9364) );
  XOR U9054 ( .A(p_input[3004]), .B(p_input[2988]), .Z(n9365) );
  XNOR U9055 ( .A(n8936), .B(n9360), .Z(n9362) );
  XOR U9056 ( .A(n9366), .B(n9367), .Z(n8936) );
  AND U9057 ( .A(n232), .B(n9368), .Z(n9367) );
  XOR U9058 ( .A(p_input[2972]), .B(p_input[2956]), .Z(n9368) );
  XOR U9059 ( .A(n9369), .B(n9370), .Z(n9360) );
  AND U9060 ( .A(n9371), .B(n9372), .Z(n9370) );
  XOR U9061 ( .A(n9369), .B(n8951), .Z(n9372) );
  XNOR U9062 ( .A(p_input[2987]), .B(n9373), .Z(n8951) );
  AND U9063 ( .A(n235), .B(n9374), .Z(n9373) );
  XOR U9064 ( .A(p_input[3003]), .B(p_input[2987]), .Z(n9374) );
  XNOR U9065 ( .A(n8948), .B(n9369), .Z(n9371) );
  XOR U9066 ( .A(n9375), .B(n9376), .Z(n8948) );
  AND U9067 ( .A(n232), .B(n9377), .Z(n9376) );
  XOR U9068 ( .A(p_input[2971]), .B(p_input[2955]), .Z(n9377) );
  XOR U9069 ( .A(n9378), .B(n9379), .Z(n9369) );
  AND U9070 ( .A(n9380), .B(n9381), .Z(n9379) );
  XOR U9071 ( .A(n9378), .B(n8963), .Z(n9381) );
  XNOR U9072 ( .A(p_input[2986]), .B(n9382), .Z(n8963) );
  AND U9073 ( .A(n235), .B(n9383), .Z(n9382) );
  XOR U9074 ( .A(p_input[3002]), .B(p_input[2986]), .Z(n9383) );
  XNOR U9075 ( .A(n8960), .B(n9378), .Z(n9380) );
  XOR U9076 ( .A(n9384), .B(n9385), .Z(n8960) );
  AND U9077 ( .A(n232), .B(n9386), .Z(n9385) );
  XOR U9078 ( .A(p_input[2970]), .B(p_input[2954]), .Z(n9386) );
  XOR U9079 ( .A(n9387), .B(n9388), .Z(n9378) );
  AND U9080 ( .A(n9389), .B(n9390), .Z(n9388) );
  XOR U9081 ( .A(n9387), .B(n8975), .Z(n9390) );
  XNOR U9082 ( .A(p_input[2985]), .B(n9391), .Z(n8975) );
  AND U9083 ( .A(n235), .B(n9392), .Z(n9391) );
  XOR U9084 ( .A(p_input[3001]), .B(p_input[2985]), .Z(n9392) );
  XNOR U9085 ( .A(n8972), .B(n9387), .Z(n9389) );
  XOR U9086 ( .A(n9393), .B(n9394), .Z(n8972) );
  AND U9087 ( .A(n232), .B(n9395), .Z(n9394) );
  XOR U9088 ( .A(p_input[2969]), .B(p_input[2953]), .Z(n9395) );
  XOR U9089 ( .A(n9396), .B(n9397), .Z(n9387) );
  AND U9090 ( .A(n9398), .B(n9399), .Z(n9397) );
  XOR U9091 ( .A(n9396), .B(n8987), .Z(n9399) );
  XNOR U9092 ( .A(p_input[2984]), .B(n9400), .Z(n8987) );
  AND U9093 ( .A(n235), .B(n9401), .Z(n9400) );
  XOR U9094 ( .A(p_input[3000]), .B(p_input[2984]), .Z(n9401) );
  XNOR U9095 ( .A(n8984), .B(n9396), .Z(n9398) );
  XOR U9096 ( .A(n9402), .B(n9403), .Z(n8984) );
  AND U9097 ( .A(n232), .B(n9404), .Z(n9403) );
  XOR U9098 ( .A(p_input[2968]), .B(p_input[2952]), .Z(n9404) );
  XOR U9099 ( .A(n9405), .B(n9406), .Z(n9396) );
  AND U9100 ( .A(n9407), .B(n9408), .Z(n9406) );
  XOR U9101 ( .A(n9405), .B(n8999), .Z(n9408) );
  XNOR U9102 ( .A(p_input[2983]), .B(n9409), .Z(n8999) );
  AND U9103 ( .A(n235), .B(n9410), .Z(n9409) );
  XOR U9104 ( .A(p_input[2999]), .B(p_input[2983]), .Z(n9410) );
  XNOR U9105 ( .A(n8996), .B(n9405), .Z(n9407) );
  XOR U9106 ( .A(n9411), .B(n9412), .Z(n8996) );
  AND U9107 ( .A(n232), .B(n9413), .Z(n9412) );
  XOR U9108 ( .A(p_input[2967]), .B(p_input[2951]), .Z(n9413) );
  XOR U9109 ( .A(n9414), .B(n9415), .Z(n9405) );
  AND U9110 ( .A(n9416), .B(n9417), .Z(n9415) );
  XOR U9111 ( .A(n9414), .B(n9011), .Z(n9417) );
  XNOR U9112 ( .A(p_input[2982]), .B(n9418), .Z(n9011) );
  AND U9113 ( .A(n235), .B(n9419), .Z(n9418) );
  XOR U9114 ( .A(p_input[2998]), .B(p_input[2982]), .Z(n9419) );
  XNOR U9115 ( .A(n9008), .B(n9414), .Z(n9416) );
  XOR U9116 ( .A(n9420), .B(n9421), .Z(n9008) );
  AND U9117 ( .A(n232), .B(n9422), .Z(n9421) );
  XOR U9118 ( .A(p_input[2966]), .B(p_input[2950]), .Z(n9422) );
  XOR U9119 ( .A(n9423), .B(n9424), .Z(n9414) );
  AND U9120 ( .A(n9425), .B(n9426), .Z(n9424) );
  XOR U9121 ( .A(n9423), .B(n9023), .Z(n9426) );
  XNOR U9122 ( .A(p_input[2981]), .B(n9427), .Z(n9023) );
  AND U9123 ( .A(n235), .B(n9428), .Z(n9427) );
  XOR U9124 ( .A(p_input[2997]), .B(p_input[2981]), .Z(n9428) );
  XNOR U9125 ( .A(n9020), .B(n9423), .Z(n9425) );
  XOR U9126 ( .A(n9429), .B(n9430), .Z(n9020) );
  AND U9127 ( .A(n232), .B(n9431), .Z(n9430) );
  XOR U9128 ( .A(p_input[2965]), .B(p_input[2949]), .Z(n9431) );
  XOR U9129 ( .A(n9432), .B(n9433), .Z(n9423) );
  AND U9130 ( .A(n9434), .B(n9435), .Z(n9433) );
  XOR U9131 ( .A(n9432), .B(n9035), .Z(n9435) );
  XNOR U9132 ( .A(p_input[2980]), .B(n9436), .Z(n9035) );
  AND U9133 ( .A(n235), .B(n9437), .Z(n9436) );
  XOR U9134 ( .A(p_input[2996]), .B(p_input[2980]), .Z(n9437) );
  XNOR U9135 ( .A(n9032), .B(n9432), .Z(n9434) );
  XOR U9136 ( .A(n9438), .B(n9439), .Z(n9032) );
  AND U9137 ( .A(n232), .B(n9440), .Z(n9439) );
  XOR U9138 ( .A(p_input[2964]), .B(p_input[2948]), .Z(n9440) );
  XOR U9139 ( .A(n9441), .B(n9442), .Z(n9432) );
  AND U9140 ( .A(n9443), .B(n9444), .Z(n9442) );
  XOR U9141 ( .A(n9441), .B(n9047), .Z(n9444) );
  XNOR U9142 ( .A(p_input[2979]), .B(n9445), .Z(n9047) );
  AND U9143 ( .A(n235), .B(n9446), .Z(n9445) );
  XOR U9144 ( .A(p_input[2995]), .B(p_input[2979]), .Z(n9446) );
  XNOR U9145 ( .A(n9044), .B(n9441), .Z(n9443) );
  XOR U9146 ( .A(n9447), .B(n9448), .Z(n9044) );
  AND U9147 ( .A(n232), .B(n9449), .Z(n9448) );
  XOR U9148 ( .A(p_input[2963]), .B(p_input[2947]), .Z(n9449) );
  XOR U9149 ( .A(n9450), .B(n9451), .Z(n9441) );
  AND U9150 ( .A(n9452), .B(n9453), .Z(n9451) );
  XOR U9151 ( .A(n9450), .B(n9059), .Z(n9453) );
  XNOR U9152 ( .A(p_input[2978]), .B(n9454), .Z(n9059) );
  AND U9153 ( .A(n235), .B(n9455), .Z(n9454) );
  XOR U9154 ( .A(p_input[2994]), .B(p_input[2978]), .Z(n9455) );
  XNOR U9155 ( .A(n9056), .B(n9450), .Z(n9452) );
  XOR U9156 ( .A(n9456), .B(n9457), .Z(n9056) );
  AND U9157 ( .A(n232), .B(n9458), .Z(n9457) );
  XOR U9158 ( .A(p_input[2962]), .B(p_input[2946]), .Z(n9458) );
  XOR U9159 ( .A(n9459), .B(n9460), .Z(n9450) );
  AND U9160 ( .A(n9461), .B(n9462), .Z(n9460) );
  XNOR U9161 ( .A(n9463), .B(n9072), .Z(n9462) );
  XNOR U9162 ( .A(p_input[2977]), .B(n9464), .Z(n9072) );
  AND U9163 ( .A(n235), .B(n9465), .Z(n9464) );
  XNOR U9164 ( .A(p_input[2993]), .B(n9466), .Z(n9465) );
  IV U9165 ( .A(p_input[2977]), .Z(n9466) );
  XNOR U9166 ( .A(n9069), .B(n9459), .Z(n9461) );
  XNOR U9167 ( .A(p_input[2945]), .B(n9467), .Z(n9069) );
  AND U9168 ( .A(n232), .B(n9468), .Z(n9467) );
  XOR U9169 ( .A(p_input[2961]), .B(p_input[2945]), .Z(n9468) );
  IV U9170 ( .A(n9463), .Z(n9459) );
  AND U9171 ( .A(n9334), .B(n9337), .Z(n9463) );
  XOR U9172 ( .A(p_input[2976]), .B(n9469), .Z(n9337) );
  AND U9173 ( .A(n235), .B(n9470), .Z(n9469) );
  XOR U9174 ( .A(p_input[2992]), .B(p_input[2976]), .Z(n9470) );
  XOR U9175 ( .A(n9471), .B(n9472), .Z(n235) );
  AND U9176 ( .A(n9473), .B(n9474), .Z(n9472) );
  XNOR U9177 ( .A(p_input[3007]), .B(n9471), .Z(n9474) );
  XOR U9178 ( .A(n9471), .B(p_input[2991]), .Z(n9473) );
  XOR U9179 ( .A(n9475), .B(n9476), .Z(n9471) );
  AND U9180 ( .A(n9477), .B(n9478), .Z(n9476) );
  XNOR U9181 ( .A(p_input[3006]), .B(n9475), .Z(n9478) );
  XOR U9182 ( .A(n9475), .B(p_input[2990]), .Z(n9477) );
  XOR U9183 ( .A(n9479), .B(n9480), .Z(n9475) );
  AND U9184 ( .A(n9481), .B(n9482), .Z(n9480) );
  XNOR U9185 ( .A(p_input[3005]), .B(n9479), .Z(n9482) );
  XOR U9186 ( .A(n9479), .B(p_input[2989]), .Z(n9481) );
  XOR U9187 ( .A(n9483), .B(n9484), .Z(n9479) );
  AND U9188 ( .A(n9485), .B(n9486), .Z(n9484) );
  XNOR U9189 ( .A(p_input[3004]), .B(n9483), .Z(n9486) );
  XOR U9190 ( .A(n9483), .B(p_input[2988]), .Z(n9485) );
  XOR U9191 ( .A(n9487), .B(n9488), .Z(n9483) );
  AND U9192 ( .A(n9489), .B(n9490), .Z(n9488) );
  XNOR U9193 ( .A(p_input[3003]), .B(n9487), .Z(n9490) );
  XOR U9194 ( .A(n9487), .B(p_input[2987]), .Z(n9489) );
  XOR U9195 ( .A(n9491), .B(n9492), .Z(n9487) );
  AND U9196 ( .A(n9493), .B(n9494), .Z(n9492) );
  XNOR U9197 ( .A(p_input[3002]), .B(n9491), .Z(n9494) );
  XOR U9198 ( .A(n9491), .B(p_input[2986]), .Z(n9493) );
  XOR U9199 ( .A(n9495), .B(n9496), .Z(n9491) );
  AND U9200 ( .A(n9497), .B(n9498), .Z(n9496) );
  XNOR U9201 ( .A(p_input[3001]), .B(n9495), .Z(n9498) );
  XOR U9202 ( .A(n9495), .B(p_input[2985]), .Z(n9497) );
  XOR U9203 ( .A(n9499), .B(n9500), .Z(n9495) );
  AND U9204 ( .A(n9501), .B(n9502), .Z(n9500) );
  XNOR U9205 ( .A(p_input[3000]), .B(n9499), .Z(n9502) );
  XOR U9206 ( .A(n9499), .B(p_input[2984]), .Z(n9501) );
  XOR U9207 ( .A(n9503), .B(n9504), .Z(n9499) );
  AND U9208 ( .A(n9505), .B(n9506), .Z(n9504) );
  XNOR U9209 ( .A(p_input[2999]), .B(n9503), .Z(n9506) );
  XOR U9210 ( .A(n9503), .B(p_input[2983]), .Z(n9505) );
  XOR U9211 ( .A(n9507), .B(n9508), .Z(n9503) );
  AND U9212 ( .A(n9509), .B(n9510), .Z(n9508) );
  XNOR U9213 ( .A(p_input[2998]), .B(n9507), .Z(n9510) );
  XOR U9214 ( .A(n9507), .B(p_input[2982]), .Z(n9509) );
  XOR U9215 ( .A(n9511), .B(n9512), .Z(n9507) );
  AND U9216 ( .A(n9513), .B(n9514), .Z(n9512) );
  XNOR U9217 ( .A(p_input[2997]), .B(n9511), .Z(n9514) );
  XOR U9218 ( .A(n9511), .B(p_input[2981]), .Z(n9513) );
  XOR U9219 ( .A(n9515), .B(n9516), .Z(n9511) );
  AND U9220 ( .A(n9517), .B(n9518), .Z(n9516) );
  XNOR U9221 ( .A(p_input[2996]), .B(n9515), .Z(n9518) );
  XOR U9222 ( .A(n9515), .B(p_input[2980]), .Z(n9517) );
  XOR U9223 ( .A(n9519), .B(n9520), .Z(n9515) );
  AND U9224 ( .A(n9521), .B(n9522), .Z(n9520) );
  XNOR U9225 ( .A(p_input[2995]), .B(n9519), .Z(n9522) );
  XOR U9226 ( .A(n9519), .B(p_input[2979]), .Z(n9521) );
  XOR U9227 ( .A(n9523), .B(n9524), .Z(n9519) );
  AND U9228 ( .A(n9525), .B(n9526), .Z(n9524) );
  XNOR U9229 ( .A(p_input[2994]), .B(n9523), .Z(n9526) );
  XOR U9230 ( .A(n9523), .B(p_input[2978]), .Z(n9525) );
  XNOR U9231 ( .A(n9527), .B(n9528), .Z(n9523) );
  AND U9232 ( .A(n9529), .B(n9530), .Z(n9528) );
  XOR U9233 ( .A(p_input[2993]), .B(n9527), .Z(n9530) );
  XNOR U9234 ( .A(p_input[2977]), .B(n9527), .Z(n9529) );
  AND U9235 ( .A(p_input[2992]), .B(n9531), .Z(n9527) );
  IV U9236 ( .A(p_input[2976]), .Z(n9531) );
  XNOR U9237 ( .A(p_input[2944]), .B(n9532), .Z(n9334) );
  AND U9238 ( .A(n232), .B(n9533), .Z(n9532) );
  XOR U9239 ( .A(p_input[2960]), .B(p_input[2944]), .Z(n9533) );
  XOR U9240 ( .A(n9534), .B(n9535), .Z(n232) );
  AND U9241 ( .A(n9536), .B(n9537), .Z(n9535) );
  XNOR U9242 ( .A(p_input[2975]), .B(n9534), .Z(n9537) );
  XOR U9243 ( .A(n9534), .B(p_input[2959]), .Z(n9536) );
  XOR U9244 ( .A(n9538), .B(n9539), .Z(n9534) );
  AND U9245 ( .A(n9540), .B(n9541), .Z(n9539) );
  XNOR U9246 ( .A(p_input[2974]), .B(n9538), .Z(n9541) );
  XNOR U9247 ( .A(n9538), .B(n9348), .Z(n9540) );
  IV U9248 ( .A(p_input[2958]), .Z(n9348) );
  XOR U9249 ( .A(n9542), .B(n9543), .Z(n9538) );
  AND U9250 ( .A(n9544), .B(n9545), .Z(n9543) );
  XNOR U9251 ( .A(p_input[2973]), .B(n9542), .Z(n9545) );
  XNOR U9252 ( .A(n9542), .B(n9357), .Z(n9544) );
  IV U9253 ( .A(p_input[2957]), .Z(n9357) );
  XOR U9254 ( .A(n9546), .B(n9547), .Z(n9542) );
  AND U9255 ( .A(n9548), .B(n9549), .Z(n9547) );
  XNOR U9256 ( .A(p_input[2972]), .B(n9546), .Z(n9549) );
  XNOR U9257 ( .A(n9546), .B(n9366), .Z(n9548) );
  IV U9258 ( .A(p_input[2956]), .Z(n9366) );
  XOR U9259 ( .A(n9550), .B(n9551), .Z(n9546) );
  AND U9260 ( .A(n9552), .B(n9553), .Z(n9551) );
  XNOR U9261 ( .A(p_input[2971]), .B(n9550), .Z(n9553) );
  XNOR U9262 ( .A(n9550), .B(n9375), .Z(n9552) );
  IV U9263 ( .A(p_input[2955]), .Z(n9375) );
  XOR U9264 ( .A(n9554), .B(n9555), .Z(n9550) );
  AND U9265 ( .A(n9556), .B(n9557), .Z(n9555) );
  XNOR U9266 ( .A(p_input[2970]), .B(n9554), .Z(n9557) );
  XNOR U9267 ( .A(n9554), .B(n9384), .Z(n9556) );
  IV U9268 ( .A(p_input[2954]), .Z(n9384) );
  XOR U9269 ( .A(n9558), .B(n9559), .Z(n9554) );
  AND U9270 ( .A(n9560), .B(n9561), .Z(n9559) );
  XNOR U9271 ( .A(p_input[2969]), .B(n9558), .Z(n9561) );
  XNOR U9272 ( .A(n9558), .B(n9393), .Z(n9560) );
  IV U9273 ( .A(p_input[2953]), .Z(n9393) );
  XOR U9274 ( .A(n9562), .B(n9563), .Z(n9558) );
  AND U9275 ( .A(n9564), .B(n9565), .Z(n9563) );
  XNOR U9276 ( .A(p_input[2968]), .B(n9562), .Z(n9565) );
  XNOR U9277 ( .A(n9562), .B(n9402), .Z(n9564) );
  IV U9278 ( .A(p_input[2952]), .Z(n9402) );
  XOR U9279 ( .A(n9566), .B(n9567), .Z(n9562) );
  AND U9280 ( .A(n9568), .B(n9569), .Z(n9567) );
  XNOR U9281 ( .A(p_input[2967]), .B(n9566), .Z(n9569) );
  XNOR U9282 ( .A(n9566), .B(n9411), .Z(n9568) );
  IV U9283 ( .A(p_input[2951]), .Z(n9411) );
  XOR U9284 ( .A(n9570), .B(n9571), .Z(n9566) );
  AND U9285 ( .A(n9572), .B(n9573), .Z(n9571) );
  XNOR U9286 ( .A(p_input[2966]), .B(n9570), .Z(n9573) );
  XNOR U9287 ( .A(n9570), .B(n9420), .Z(n9572) );
  IV U9288 ( .A(p_input[2950]), .Z(n9420) );
  XOR U9289 ( .A(n9574), .B(n9575), .Z(n9570) );
  AND U9290 ( .A(n9576), .B(n9577), .Z(n9575) );
  XNOR U9291 ( .A(p_input[2965]), .B(n9574), .Z(n9577) );
  XNOR U9292 ( .A(n9574), .B(n9429), .Z(n9576) );
  IV U9293 ( .A(p_input[2949]), .Z(n9429) );
  XOR U9294 ( .A(n9578), .B(n9579), .Z(n9574) );
  AND U9295 ( .A(n9580), .B(n9581), .Z(n9579) );
  XNOR U9296 ( .A(p_input[2964]), .B(n9578), .Z(n9581) );
  XNOR U9297 ( .A(n9578), .B(n9438), .Z(n9580) );
  IV U9298 ( .A(p_input[2948]), .Z(n9438) );
  XOR U9299 ( .A(n9582), .B(n9583), .Z(n9578) );
  AND U9300 ( .A(n9584), .B(n9585), .Z(n9583) );
  XNOR U9301 ( .A(p_input[2963]), .B(n9582), .Z(n9585) );
  XNOR U9302 ( .A(n9582), .B(n9447), .Z(n9584) );
  IV U9303 ( .A(p_input[2947]), .Z(n9447) );
  XOR U9304 ( .A(n9586), .B(n9587), .Z(n9582) );
  AND U9305 ( .A(n9588), .B(n9589), .Z(n9587) );
  XNOR U9306 ( .A(p_input[2962]), .B(n9586), .Z(n9589) );
  XNOR U9307 ( .A(n9586), .B(n9456), .Z(n9588) );
  IV U9308 ( .A(p_input[2946]), .Z(n9456) );
  XNOR U9309 ( .A(n9590), .B(n9591), .Z(n9586) );
  AND U9310 ( .A(n9592), .B(n9593), .Z(n9591) );
  XOR U9311 ( .A(p_input[2961]), .B(n9590), .Z(n9593) );
  XNOR U9312 ( .A(p_input[2945]), .B(n9590), .Z(n9592) );
  AND U9313 ( .A(p_input[2960]), .B(n9594), .Z(n9590) );
  IV U9314 ( .A(p_input[2944]), .Z(n9594) );
  XOR U9315 ( .A(n9595), .B(n9596), .Z(n8710) );
  AND U9316 ( .A(n761), .B(n9597), .Z(n9596) );
  XNOR U9317 ( .A(n9598), .B(n9595), .Z(n9597) );
  XOR U9318 ( .A(n9599), .B(n9600), .Z(n761) );
  AND U9319 ( .A(n9601), .B(n9602), .Z(n9600) );
  XNOR U9320 ( .A(n8722), .B(n9599), .Z(n9602) );
  AND U9321 ( .A(n9603), .B(n9604), .Z(n8722) );
  XOR U9322 ( .A(n9599), .B(n8721), .Z(n9601) );
  AND U9323 ( .A(n9605), .B(n9606), .Z(n8721) );
  XOR U9324 ( .A(n9607), .B(n9608), .Z(n9599) );
  AND U9325 ( .A(n9609), .B(n9610), .Z(n9608) );
  XOR U9326 ( .A(n9607), .B(n8734), .Z(n9610) );
  XOR U9327 ( .A(n9611), .B(n9612), .Z(n8734) );
  AND U9328 ( .A(n423), .B(n9613), .Z(n9612) );
  XOR U9329 ( .A(n9614), .B(n9611), .Z(n9613) );
  XNOR U9330 ( .A(n8731), .B(n9607), .Z(n9609) );
  XOR U9331 ( .A(n9615), .B(n9616), .Z(n8731) );
  AND U9332 ( .A(n420), .B(n9617), .Z(n9616) );
  XOR U9333 ( .A(n9618), .B(n9615), .Z(n9617) );
  XOR U9334 ( .A(n9619), .B(n9620), .Z(n9607) );
  AND U9335 ( .A(n9621), .B(n9622), .Z(n9620) );
  XOR U9336 ( .A(n9619), .B(n8746), .Z(n9622) );
  XOR U9337 ( .A(n9623), .B(n9624), .Z(n8746) );
  AND U9338 ( .A(n423), .B(n9625), .Z(n9624) );
  XOR U9339 ( .A(n9626), .B(n9623), .Z(n9625) );
  XNOR U9340 ( .A(n8743), .B(n9619), .Z(n9621) );
  XOR U9341 ( .A(n9627), .B(n9628), .Z(n8743) );
  AND U9342 ( .A(n420), .B(n9629), .Z(n9628) );
  XOR U9343 ( .A(n9630), .B(n9627), .Z(n9629) );
  XOR U9344 ( .A(n9631), .B(n9632), .Z(n9619) );
  AND U9345 ( .A(n9633), .B(n9634), .Z(n9632) );
  XOR U9346 ( .A(n9631), .B(n8758), .Z(n9634) );
  XOR U9347 ( .A(n9635), .B(n9636), .Z(n8758) );
  AND U9348 ( .A(n423), .B(n9637), .Z(n9636) );
  XOR U9349 ( .A(n9638), .B(n9635), .Z(n9637) );
  XNOR U9350 ( .A(n8755), .B(n9631), .Z(n9633) );
  XOR U9351 ( .A(n9639), .B(n9640), .Z(n8755) );
  AND U9352 ( .A(n420), .B(n9641), .Z(n9640) );
  XOR U9353 ( .A(n9642), .B(n9639), .Z(n9641) );
  XOR U9354 ( .A(n9643), .B(n9644), .Z(n9631) );
  AND U9355 ( .A(n9645), .B(n9646), .Z(n9644) );
  XOR U9356 ( .A(n9643), .B(n8770), .Z(n9646) );
  XOR U9357 ( .A(n9647), .B(n9648), .Z(n8770) );
  AND U9358 ( .A(n423), .B(n9649), .Z(n9648) );
  XOR U9359 ( .A(n9650), .B(n9647), .Z(n9649) );
  XNOR U9360 ( .A(n8767), .B(n9643), .Z(n9645) );
  XOR U9361 ( .A(n9651), .B(n9652), .Z(n8767) );
  AND U9362 ( .A(n420), .B(n9653), .Z(n9652) );
  XOR U9363 ( .A(n9654), .B(n9651), .Z(n9653) );
  XOR U9364 ( .A(n9655), .B(n9656), .Z(n9643) );
  AND U9365 ( .A(n9657), .B(n9658), .Z(n9656) );
  XOR U9366 ( .A(n9655), .B(n8782), .Z(n9658) );
  XOR U9367 ( .A(n9659), .B(n9660), .Z(n8782) );
  AND U9368 ( .A(n423), .B(n9661), .Z(n9660) );
  XOR U9369 ( .A(n9662), .B(n9659), .Z(n9661) );
  XNOR U9370 ( .A(n8779), .B(n9655), .Z(n9657) );
  XOR U9371 ( .A(n9663), .B(n9664), .Z(n8779) );
  AND U9372 ( .A(n420), .B(n9665), .Z(n9664) );
  XOR U9373 ( .A(n9666), .B(n9663), .Z(n9665) );
  XOR U9374 ( .A(n9667), .B(n9668), .Z(n9655) );
  AND U9375 ( .A(n9669), .B(n9670), .Z(n9668) );
  XOR U9376 ( .A(n9667), .B(n8794), .Z(n9670) );
  XOR U9377 ( .A(n9671), .B(n9672), .Z(n8794) );
  AND U9378 ( .A(n423), .B(n9673), .Z(n9672) );
  XOR U9379 ( .A(n9674), .B(n9671), .Z(n9673) );
  XNOR U9380 ( .A(n8791), .B(n9667), .Z(n9669) );
  XOR U9381 ( .A(n9675), .B(n9676), .Z(n8791) );
  AND U9382 ( .A(n420), .B(n9677), .Z(n9676) );
  XOR U9383 ( .A(n9678), .B(n9675), .Z(n9677) );
  XOR U9384 ( .A(n9679), .B(n9680), .Z(n9667) );
  AND U9385 ( .A(n9681), .B(n9682), .Z(n9680) );
  XOR U9386 ( .A(n9679), .B(n8806), .Z(n9682) );
  XOR U9387 ( .A(n9683), .B(n9684), .Z(n8806) );
  AND U9388 ( .A(n423), .B(n9685), .Z(n9684) );
  XOR U9389 ( .A(n9686), .B(n9683), .Z(n9685) );
  XNOR U9390 ( .A(n8803), .B(n9679), .Z(n9681) );
  XOR U9391 ( .A(n9687), .B(n9688), .Z(n8803) );
  AND U9392 ( .A(n420), .B(n9689), .Z(n9688) );
  XOR U9393 ( .A(n9690), .B(n9687), .Z(n9689) );
  XOR U9394 ( .A(n9691), .B(n9692), .Z(n9679) );
  AND U9395 ( .A(n9693), .B(n9694), .Z(n9692) );
  XOR U9396 ( .A(n9691), .B(n8818), .Z(n9694) );
  XOR U9397 ( .A(n9695), .B(n9696), .Z(n8818) );
  AND U9398 ( .A(n423), .B(n9697), .Z(n9696) );
  XOR U9399 ( .A(n9698), .B(n9695), .Z(n9697) );
  XNOR U9400 ( .A(n8815), .B(n9691), .Z(n9693) );
  XOR U9401 ( .A(n9699), .B(n9700), .Z(n8815) );
  AND U9402 ( .A(n420), .B(n9701), .Z(n9700) );
  XOR U9403 ( .A(n9702), .B(n9699), .Z(n9701) );
  XOR U9404 ( .A(n9703), .B(n9704), .Z(n9691) );
  AND U9405 ( .A(n9705), .B(n9706), .Z(n9704) );
  XOR U9406 ( .A(n9703), .B(n8830), .Z(n9706) );
  XOR U9407 ( .A(n9707), .B(n9708), .Z(n8830) );
  AND U9408 ( .A(n423), .B(n9709), .Z(n9708) );
  XOR U9409 ( .A(n9710), .B(n9707), .Z(n9709) );
  XNOR U9410 ( .A(n8827), .B(n9703), .Z(n9705) );
  XOR U9411 ( .A(n9711), .B(n9712), .Z(n8827) );
  AND U9412 ( .A(n420), .B(n9713), .Z(n9712) );
  XOR U9413 ( .A(n9714), .B(n9711), .Z(n9713) );
  XOR U9414 ( .A(n9715), .B(n9716), .Z(n9703) );
  AND U9415 ( .A(n9717), .B(n9718), .Z(n9716) );
  XOR U9416 ( .A(n9715), .B(n8842), .Z(n9718) );
  XOR U9417 ( .A(n9719), .B(n9720), .Z(n8842) );
  AND U9418 ( .A(n423), .B(n9721), .Z(n9720) );
  XOR U9419 ( .A(n9722), .B(n9719), .Z(n9721) );
  XNOR U9420 ( .A(n8839), .B(n9715), .Z(n9717) );
  XOR U9421 ( .A(n9723), .B(n9724), .Z(n8839) );
  AND U9422 ( .A(n420), .B(n9725), .Z(n9724) );
  XOR U9423 ( .A(n9726), .B(n9723), .Z(n9725) );
  XOR U9424 ( .A(n9727), .B(n9728), .Z(n9715) );
  AND U9425 ( .A(n9729), .B(n9730), .Z(n9728) );
  XOR U9426 ( .A(n9727), .B(n8854), .Z(n9730) );
  XOR U9427 ( .A(n9731), .B(n9732), .Z(n8854) );
  AND U9428 ( .A(n423), .B(n9733), .Z(n9732) );
  XOR U9429 ( .A(n9734), .B(n9731), .Z(n9733) );
  XNOR U9430 ( .A(n8851), .B(n9727), .Z(n9729) );
  XOR U9431 ( .A(n9735), .B(n9736), .Z(n8851) );
  AND U9432 ( .A(n420), .B(n9737), .Z(n9736) );
  XOR U9433 ( .A(n9738), .B(n9735), .Z(n9737) );
  XOR U9434 ( .A(n9739), .B(n9740), .Z(n9727) );
  AND U9435 ( .A(n9741), .B(n9742), .Z(n9740) );
  XOR U9436 ( .A(n9739), .B(n8866), .Z(n9742) );
  XOR U9437 ( .A(n9743), .B(n9744), .Z(n8866) );
  AND U9438 ( .A(n423), .B(n9745), .Z(n9744) );
  XOR U9439 ( .A(n9746), .B(n9743), .Z(n9745) );
  XNOR U9440 ( .A(n8863), .B(n9739), .Z(n9741) );
  XOR U9441 ( .A(n9747), .B(n9748), .Z(n8863) );
  AND U9442 ( .A(n420), .B(n9749), .Z(n9748) );
  XOR U9443 ( .A(n9750), .B(n9747), .Z(n9749) );
  XOR U9444 ( .A(n9751), .B(n9752), .Z(n9739) );
  AND U9445 ( .A(n9753), .B(n9754), .Z(n9752) );
  XOR U9446 ( .A(n9751), .B(n8878), .Z(n9754) );
  XOR U9447 ( .A(n9755), .B(n9756), .Z(n8878) );
  AND U9448 ( .A(n423), .B(n9757), .Z(n9756) );
  XOR U9449 ( .A(n9758), .B(n9755), .Z(n9757) );
  XNOR U9450 ( .A(n8875), .B(n9751), .Z(n9753) );
  XOR U9451 ( .A(n9759), .B(n9760), .Z(n8875) );
  AND U9452 ( .A(n420), .B(n9761), .Z(n9760) );
  XOR U9453 ( .A(n9762), .B(n9759), .Z(n9761) );
  XOR U9454 ( .A(n9763), .B(n9764), .Z(n9751) );
  AND U9455 ( .A(n9765), .B(n9766), .Z(n9764) );
  XNOR U9456 ( .A(n9767), .B(n8891), .Z(n9766) );
  XOR U9457 ( .A(n9768), .B(n9769), .Z(n8891) );
  AND U9458 ( .A(n423), .B(n9770), .Z(n9769) );
  XOR U9459 ( .A(n9768), .B(n9771), .Z(n9770) );
  XNOR U9460 ( .A(n8888), .B(n9763), .Z(n9765) );
  XOR U9461 ( .A(n9772), .B(n9773), .Z(n8888) );
  AND U9462 ( .A(n420), .B(n9774), .Z(n9773) );
  XOR U9463 ( .A(n9772), .B(n9775), .Z(n9774) );
  IV U9464 ( .A(n9767), .Z(n9763) );
  AND U9465 ( .A(n9595), .B(n9598), .Z(n9767) );
  XNOR U9466 ( .A(n9776), .B(n9777), .Z(n9598) );
  AND U9467 ( .A(n423), .B(n9778), .Z(n9777) );
  XNOR U9468 ( .A(n9779), .B(n9776), .Z(n9778) );
  XOR U9469 ( .A(n9780), .B(n9781), .Z(n423) );
  AND U9470 ( .A(n9782), .B(n9783), .Z(n9781) );
  XNOR U9471 ( .A(n9603), .B(n9780), .Z(n9783) );
  AND U9472 ( .A(p_input[2943]), .B(p_input[2927]), .Z(n9603) );
  XOR U9473 ( .A(n9780), .B(n9604), .Z(n9782) );
  AND U9474 ( .A(p_input[2911]), .B(p_input[2895]), .Z(n9604) );
  XOR U9475 ( .A(n9784), .B(n9785), .Z(n9780) );
  AND U9476 ( .A(n9786), .B(n9787), .Z(n9785) );
  XOR U9477 ( .A(n9784), .B(n9614), .Z(n9787) );
  XNOR U9478 ( .A(p_input[2926]), .B(n9788), .Z(n9614) );
  AND U9479 ( .A(n243), .B(n9789), .Z(n9788) );
  XOR U9480 ( .A(p_input[2942]), .B(p_input[2926]), .Z(n9789) );
  XNOR U9481 ( .A(n9611), .B(n9784), .Z(n9786) );
  XOR U9482 ( .A(n9790), .B(n9791), .Z(n9611) );
  AND U9483 ( .A(n241), .B(n9792), .Z(n9791) );
  XOR U9484 ( .A(p_input[2910]), .B(p_input[2894]), .Z(n9792) );
  XOR U9485 ( .A(n9793), .B(n9794), .Z(n9784) );
  AND U9486 ( .A(n9795), .B(n9796), .Z(n9794) );
  XOR U9487 ( .A(n9793), .B(n9626), .Z(n9796) );
  XNOR U9488 ( .A(p_input[2925]), .B(n9797), .Z(n9626) );
  AND U9489 ( .A(n243), .B(n9798), .Z(n9797) );
  XOR U9490 ( .A(p_input[2941]), .B(p_input[2925]), .Z(n9798) );
  XNOR U9491 ( .A(n9623), .B(n9793), .Z(n9795) );
  XOR U9492 ( .A(n9799), .B(n9800), .Z(n9623) );
  AND U9493 ( .A(n241), .B(n9801), .Z(n9800) );
  XOR U9494 ( .A(p_input[2909]), .B(p_input[2893]), .Z(n9801) );
  XOR U9495 ( .A(n9802), .B(n9803), .Z(n9793) );
  AND U9496 ( .A(n9804), .B(n9805), .Z(n9803) );
  XOR U9497 ( .A(n9802), .B(n9638), .Z(n9805) );
  XNOR U9498 ( .A(p_input[2924]), .B(n9806), .Z(n9638) );
  AND U9499 ( .A(n243), .B(n9807), .Z(n9806) );
  XOR U9500 ( .A(p_input[2940]), .B(p_input[2924]), .Z(n9807) );
  XNOR U9501 ( .A(n9635), .B(n9802), .Z(n9804) );
  XOR U9502 ( .A(n9808), .B(n9809), .Z(n9635) );
  AND U9503 ( .A(n241), .B(n9810), .Z(n9809) );
  XOR U9504 ( .A(p_input[2908]), .B(p_input[2892]), .Z(n9810) );
  XOR U9505 ( .A(n9811), .B(n9812), .Z(n9802) );
  AND U9506 ( .A(n9813), .B(n9814), .Z(n9812) );
  XOR U9507 ( .A(n9811), .B(n9650), .Z(n9814) );
  XNOR U9508 ( .A(p_input[2923]), .B(n9815), .Z(n9650) );
  AND U9509 ( .A(n243), .B(n9816), .Z(n9815) );
  XOR U9510 ( .A(p_input[2939]), .B(p_input[2923]), .Z(n9816) );
  XNOR U9511 ( .A(n9647), .B(n9811), .Z(n9813) );
  XOR U9512 ( .A(n9817), .B(n9818), .Z(n9647) );
  AND U9513 ( .A(n241), .B(n9819), .Z(n9818) );
  XOR U9514 ( .A(p_input[2907]), .B(p_input[2891]), .Z(n9819) );
  XOR U9515 ( .A(n9820), .B(n9821), .Z(n9811) );
  AND U9516 ( .A(n9822), .B(n9823), .Z(n9821) );
  XOR U9517 ( .A(n9820), .B(n9662), .Z(n9823) );
  XNOR U9518 ( .A(p_input[2922]), .B(n9824), .Z(n9662) );
  AND U9519 ( .A(n243), .B(n9825), .Z(n9824) );
  XOR U9520 ( .A(p_input[2938]), .B(p_input[2922]), .Z(n9825) );
  XNOR U9521 ( .A(n9659), .B(n9820), .Z(n9822) );
  XOR U9522 ( .A(n9826), .B(n9827), .Z(n9659) );
  AND U9523 ( .A(n241), .B(n9828), .Z(n9827) );
  XOR U9524 ( .A(p_input[2906]), .B(p_input[2890]), .Z(n9828) );
  XOR U9525 ( .A(n9829), .B(n9830), .Z(n9820) );
  AND U9526 ( .A(n9831), .B(n9832), .Z(n9830) );
  XOR U9527 ( .A(n9829), .B(n9674), .Z(n9832) );
  XNOR U9528 ( .A(p_input[2921]), .B(n9833), .Z(n9674) );
  AND U9529 ( .A(n243), .B(n9834), .Z(n9833) );
  XOR U9530 ( .A(p_input[2937]), .B(p_input[2921]), .Z(n9834) );
  XNOR U9531 ( .A(n9671), .B(n9829), .Z(n9831) );
  XOR U9532 ( .A(n9835), .B(n9836), .Z(n9671) );
  AND U9533 ( .A(n241), .B(n9837), .Z(n9836) );
  XOR U9534 ( .A(p_input[2905]), .B(p_input[2889]), .Z(n9837) );
  XOR U9535 ( .A(n9838), .B(n9839), .Z(n9829) );
  AND U9536 ( .A(n9840), .B(n9841), .Z(n9839) );
  XOR U9537 ( .A(n9838), .B(n9686), .Z(n9841) );
  XNOR U9538 ( .A(p_input[2920]), .B(n9842), .Z(n9686) );
  AND U9539 ( .A(n243), .B(n9843), .Z(n9842) );
  XOR U9540 ( .A(p_input[2936]), .B(p_input[2920]), .Z(n9843) );
  XNOR U9541 ( .A(n9683), .B(n9838), .Z(n9840) );
  XOR U9542 ( .A(n9844), .B(n9845), .Z(n9683) );
  AND U9543 ( .A(n241), .B(n9846), .Z(n9845) );
  XOR U9544 ( .A(p_input[2904]), .B(p_input[2888]), .Z(n9846) );
  XOR U9545 ( .A(n9847), .B(n9848), .Z(n9838) );
  AND U9546 ( .A(n9849), .B(n9850), .Z(n9848) );
  XOR U9547 ( .A(n9847), .B(n9698), .Z(n9850) );
  XNOR U9548 ( .A(p_input[2919]), .B(n9851), .Z(n9698) );
  AND U9549 ( .A(n243), .B(n9852), .Z(n9851) );
  XOR U9550 ( .A(p_input[2935]), .B(p_input[2919]), .Z(n9852) );
  XNOR U9551 ( .A(n9695), .B(n9847), .Z(n9849) );
  XOR U9552 ( .A(n9853), .B(n9854), .Z(n9695) );
  AND U9553 ( .A(n241), .B(n9855), .Z(n9854) );
  XOR U9554 ( .A(p_input[2903]), .B(p_input[2887]), .Z(n9855) );
  XOR U9555 ( .A(n9856), .B(n9857), .Z(n9847) );
  AND U9556 ( .A(n9858), .B(n9859), .Z(n9857) );
  XOR U9557 ( .A(n9856), .B(n9710), .Z(n9859) );
  XNOR U9558 ( .A(p_input[2918]), .B(n9860), .Z(n9710) );
  AND U9559 ( .A(n243), .B(n9861), .Z(n9860) );
  XOR U9560 ( .A(p_input[2934]), .B(p_input[2918]), .Z(n9861) );
  XNOR U9561 ( .A(n9707), .B(n9856), .Z(n9858) );
  XOR U9562 ( .A(n9862), .B(n9863), .Z(n9707) );
  AND U9563 ( .A(n241), .B(n9864), .Z(n9863) );
  XOR U9564 ( .A(p_input[2902]), .B(p_input[2886]), .Z(n9864) );
  XOR U9565 ( .A(n9865), .B(n9866), .Z(n9856) );
  AND U9566 ( .A(n9867), .B(n9868), .Z(n9866) );
  XOR U9567 ( .A(n9865), .B(n9722), .Z(n9868) );
  XNOR U9568 ( .A(p_input[2917]), .B(n9869), .Z(n9722) );
  AND U9569 ( .A(n243), .B(n9870), .Z(n9869) );
  XOR U9570 ( .A(p_input[2933]), .B(p_input[2917]), .Z(n9870) );
  XNOR U9571 ( .A(n9719), .B(n9865), .Z(n9867) );
  XOR U9572 ( .A(n9871), .B(n9872), .Z(n9719) );
  AND U9573 ( .A(n241), .B(n9873), .Z(n9872) );
  XOR U9574 ( .A(p_input[2901]), .B(p_input[2885]), .Z(n9873) );
  XOR U9575 ( .A(n9874), .B(n9875), .Z(n9865) );
  AND U9576 ( .A(n9876), .B(n9877), .Z(n9875) );
  XOR U9577 ( .A(n9874), .B(n9734), .Z(n9877) );
  XNOR U9578 ( .A(p_input[2916]), .B(n9878), .Z(n9734) );
  AND U9579 ( .A(n243), .B(n9879), .Z(n9878) );
  XOR U9580 ( .A(p_input[2932]), .B(p_input[2916]), .Z(n9879) );
  XNOR U9581 ( .A(n9731), .B(n9874), .Z(n9876) );
  XOR U9582 ( .A(n9880), .B(n9881), .Z(n9731) );
  AND U9583 ( .A(n241), .B(n9882), .Z(n9881) );
  XOR U9584 ( .A(p_input[2900]), .B(p_input[2884]), .Z(n9882) );
  XOR U9585 ( .A(n9883), .B(n9884), .Z(n9874) );
  AND U9586 ( .A(n9885), .B(n9886), .Z(n9884) );
  XOR U9587 ( .A(n9883), .B(n9746), .Z(n9886) );
  XNOR U9588 ( .A(p_input[2915]), .B(n9887), .Z(n9746) );
  AND U9589 ( .A(n243), .B(n9888), .Z(n9887) );
  XOR U9590 ( .A(p_input[2931]), .B(p_input[2915]), .Z(n9888) );
  XNOR U9591 ( .A(n9743), .B(n9883), .Z(n9885) );
  XOR U9592 ( .A(n9889), .B(n9890), .Z(n9743) );
  AND U9593 ( .A(n241), .B(n9891), .Z(n9890) );
  XOR U9594 ( .A(p_input[2899]), .B(p_input[2883]), .Z(n9891) );
  XOR U9595 ( .A(n9892), .B(n9893), .Z(n9883) );
  AND U9596 ( .A(n9894), .B(n9895), .Z(n9893) );
  XOR U9597 ( .A(n9892), .B(n9758), .Z(n9895) );
  XNOR U9598 ( .A(p_input[2914]), .B(n9896), .Z(n9758) );
  AND U9599 ( .A(n243), .B(n9897), .Z(n9896) );
  XOR U9600 ( .A(p_input[2930]), .B(p_input[2914]), .Z(n9897) );
  XNOR U9601 ( .A(n9755), .B(n9892), .Z(n9894) );
  XOR U9602 ( .A(n9898), .B(n9899), .Z(n9755) );
  AND U9603 ( .A(n241), .B(n9900), .Z(n9899) );
  XOR U9604 ( .A(p_input[2898]), .B(p_input[2882]), .Z(n9900) );
  XOR U9605 ( .A(n9901), .B(n9902), .Z(n9892) );
  AND U9606 ( .A(n9903), .B(n9904), .Z(n9902) );
  XNOR U9607 ( .A(n9905), .B(n9771), .Z(n9904) );
  XNOR U9608 ( .A(p_input[2913]), .B(n9906), .Z(n9771) );
  AND U9609 ( .A(n243), .B(n9907), .Z(n9906) );
  XNOR U9610 ( .A(p_input[2929]), .B(n9908), .Z(n9907) );
  IV U9611 ( .A(p_input[2913]), .Z(n9908) );
  XNOR U9612 ( .A(n9768), .B(n9901), .Z(n9903) );
  XNOR U9613 ( .A(p_input[2881]), .B(n9909), .Z(n9768) );
  AND U9614 ( .A(n241), .B(n9910), .Z(n9909) );
  XOR U9615 ( .A(p_input[2897]), .B(p_input[2881]), .Z(n9910) );
  IV U9616 ( .A(n9905), .Z(n9901) );
  AND U9617 ( .A(n9776), .B(n9779), .Z(n9905) );
  XOR U9618 ( .A(p_input[2912]), .B(n9911), .Z(n9779) );
  AND U9619 ( .A(n243), .B(n9912), .Z(n9911) );
  XOR U9620 ( .A(p_input[2928]), .B(p_input[2912]), .Z(n9912) );
  XOR U9621 ( .A(n9913), .B(n9914), .Z(n243) );
  AND U9622 ( .A(n9915), .B(n9916), .Z(n9914) );
  XNOR U9623 ( .A(p_input[2943]), .B(n9913), .Z(n9916) );
  XOR U9624 ( .A(n9913), .B(p_input[2927]), .Z(n9915) );
  XOR U9625 ( .A(n9917), .B(n9918), .Z(n9913) );
  AND U9626 ( .A(n9919), .B(n9920), .Z(n9918) );
  XNOR U9627 ( .A(p_input[2942]), .B(n9917), .Z(n9920) );
  XOR U9628 ( .A(n9917), .B(p_input[2926]), .Z(n9919) );
  XOR U9629 ( .A(n9921), .B(n9922), .Z(n9917) );
  AND U9630 ( .A(n9923), .B(n9924), .Z(n9922) );
  XNOR U9631 ( .A(p_input[2941]), .B(n9921), .Z(n9924) );
  XOR U9632 ( .A(n9921), .B(p_input[2925]), .Z(n9923) );
  XOR U9633 ( .A(n9925), .B(n9926), .Z(n9921) );
  AND U9634 ( .A(n9927), .B(n9928), .Z(n9926) );
  XNOR U9635 ( .A(p_input[2940]), .B(n9925), .Z(n9928) );
  XOR U9636 ( .A(n9925), .B(p_input[2924]), .Z(n9927) );
  XOR U9637 ( .A(n9929), .B(n9930), .Z(n9925) );
  AND U9638 ( .A(n9931), .B(n9932), .Z(n9930) );
  XNOR U9639 ( .A(p_input[2939]), .B(n9929), .Z(n9932) );
  XOR U9640 ( .A(n9929), .B(p_input[2923]), .Z(n9931) );
  XOR U9641 ( .A(n9933), .B(n9934), .Z(n9929) );
  AND U9642 ( .A(n9935), .B(n9936), .Z(n9934) );
  XNOR U9643 ( .A(p_input[2938]), .B(n9933), .Z(n9936) );
  XOR U9644 ( .A(n9933), .B(p_input[2922]), .Z(n9935) );
  XOR U9645 ( .A(n9937), .B(n9938), .Z(n9933) );
  AND U9646 ( .A(n9939), .B(n9940), .Z(n9938) );
  XNOR U9647 ( .A(p_input[2937]), .B(n9937), .Z(n9940) );
  XOR U9648 ( .A(n9937), .B(p_input[2921]), .Z(n9939) );
  XOR U9649 ( .A(n9941), .B(n9942), .Z(n9937) );
  AND U9650 ( .A(n9943), .B(n9944), .Z(n9942) );
  XNOR U9651 ( .A(p_input[2936]), .B(n9941), .Z(n9944) );
  XOR U9652 ( .A(n9941), .B(p_input[2920]), .Z(n9943) );
  XOR U9653 ( .A(n9945), .B(n9946), .Z(n9941) );
  AND U9654 ( .A(n9947), .B(n9948), .Z(n9946) );
  XNOR U9655 ( .A(p_input[2935]), .B(n9945), .Z(n9948) );
  XOR U9656 ( .A(n9945), .B(p_input[2919]), .Z(n9947) );
  XOR U9657 ( .A(n9949), .B(n9950), .Z(n9945) );
  AND U9658 ( .A(n9951), .B(n9952), .Z(n9950) );
  XNOR U9659 ( .A(p_input[2934]), .B(n9949), .Z(n9952) );
  XOR U9660 ( .A(n9949), .B(p_input[2918]), .Z(n9951) );
  XOR U9661 ( .A(n9953), .B(n9954), .Z(n9949) );
  AND U9662 ( .A(n9955), .B(n9956), .Z(n9954) );
  XNOR U9663 ( .A(p_input[2933]), .B(n9953), .Z(n9956) );
  XOR U9664 ( .A(n9953), .B(p_input[2917]), .Z(n9955) );
  XOR U9665 ( .A(n9957), .B(n9958), .Z(n9953) );
  AND U9666 ( .A(n9959), .B(n9960), .Z(n9958) );
  XNOR U9667 ( .A(p_input[2932]), .B(n9957), .Z(n9960) );
  XOR U9668 ( .A(n9957), .B(p_input[2916]), .Z(n9959) );
  XOR U9669 ( .A(n9961), .B(n9962), .Z(n9957) );
  AND U9670 ( .A(n9963), .B(n9964), .Z(n9962) );
  XNOR U9671 ( .A(p_input[2931]), .B(n9961), .Z(n9964) );
  XOR U9672 ( .A(n9961), .B(p_input[2915]), .Z(n9963) );
  XOR U9673 ( .A(n9965), .B(n9966), .Z(n9961) );
  AND U9674 ( .A(n9967), .B(n9968), .Z(n9966) );
  XNOR U9675 ( .A(p_input[2930]), .B(n9965), .Z(n9968) );
  XOR U9676 ( .A(n9965), .B(p_input[2914]), .Z(n9967) );
  XNOR U9677 ( .A(n9969), .B(n9970), .Z(n9965) );
  AND U9678 ( .A(n9971), .B(n9972), .Z(n9970) );
  XOR U9679 ( .A(p_input[2929]), .B(n9969), .Z(n9972) );
  XNOR U9680 ( .A(p_input[2913]), .B(n9969), .Z(n9971) );
  AND U9681 ( .A(p_input[2928]), .B(n9973), .Z(n9969) );
  IV U9682 ( .A(p_input[2912]), .Z(n9973) );
  XNOR U9683 ( .A(p_input[2880]), .B(n9974), .Z(n9776) );
  AND U9684 ( .A(n241), .B(n9975), .Z(n9974) );
  XOR U9685 ( .A(p_input[2896]), .B(p_input[2880]), .Z(n9975) );
  XOR U9686 ( .A(n9976), .B(n9977), .Z(n241) );
  AND U9687 ( .A(n9978), .B(n9979), .Z(n9977) );
  XNOR U9688 ( .A(p_input[2911]), .B(n9976), .Z(n9979) );
  XOR U9689 ( .A(n9976), .B(p_input[2895]), .Z(n9978) );
  XOR U9690 ( .A(n9980), .B(n9981), .Z(n9976) );
  AND U9691 ( .A(n9982), .B(n9983), .Z(n9981) );
  XNOR U9692 ( .A(p_input[2910]), .B(n9980), .Z(n9983) );
  XNOR U9693 ( .A(n9980), .B(n9790), .Z(n9982) );
  IV U9694 ( .A(p_input[2894]), .Z(n9790) );
  XOR U9695 ( .A(n9984), .B(n9985), .Z(n9980) );
  AND U9696 ( .A(n9986), .B(n9987), .Z(n9985) );
  XNOR U9697 ( .A(p_input[2909]), .B(n9984), .Z(n9987) );
  XNOR U9698 ( .A(n9984), .B(n9799), .Z(n9986) );
  IV U9699 ( .A(p_input[2893]), .Z(n9799) );
  XOR U9700 ( .A(n9988), .B(n9989), .Z(n9984) );
  AND U9701 ( .A(n9990), .B(n9991), .Z(n9989) );
  XNOR U9702 ( .A(p_input[2908]), .B(n9988), .Z(n9991) );
  XNOR U9703 ( .A(n9988), .B(n9808), .Z(n9990) );
  IV U9704 ( .A(p_input[2892]), .Z(n9808) );
  XOR U9705 ( .A(n9992), .B(n9993), .Z(n9988) );
  AND U9706 ( .A(n9994), .B(n9995), .Z(n9993) );
  XNOR U9707 ( .A(p_input[2907]), .B(n9992), .Z(n9995) );
  XNOR U9708 ( .A(n9992), .B(n9817), .Z(n9994) );
  IV U9709 ( .A(p_input[2891]), .Z(n9817) );
  XOR U9710 ( .A(n9996), .B(n9997), .Z(n9992) );
  AND U9711 ( .A(n9998), .B(n9999), .Z(n9997) );
  XNOR U9712 ( .A(p_input[2906]), .B(n9996), .Z(n9999) );
  XNOR U9713 ( .A(n9996), .B(n9826), .Z(n9998) );
  IV U9714 ( .A(p_input[2890]), .Z(n9826) );
  XOR U9715 ( .A(n10000), .B(n10001), .Z(n9996) );
  AND U9716 ( .A(n10002), .B(n10003), .Z(n10001) );
  XNOR U9717 ( .A(p_input[2905]), .B(n10000), .Z(n10003) );
  XNOR U9718 ( .A(n10000), .B(n9835), .Z(n10002) );
  IV U9719 ( .A(p_input[2889]), .Z(n9835) );
  XOR U9720 ( .A(n10004), .B(n10005), .Z(n10000) );
  AND U9721 ( .A(n10006), .B(n10007), .Z(n10005) );
  XNOR U9722 ( .A(p_input[2904]), .B(n10004), .Z(n10007) );
  XNOR U9723 ( .A(n10004), .B(n9844), .Z(n10006) );
  IV U9724 ( .A(p_input[2888]), .Z(n9844) );
  XOR U9725 ( .A(n10008), .B(n10009), .Z(n10004) );
  AND U9726 ( .A(n10010), .B(n10011), .Z(n10009) );
  XNOR U9727 ( .A(p_input[2903]), .B(n10008), .Z(n10011) );
  XNOR U9728 ( .A(n10008), .B(n9853), .Z(n10010) );
  IV U9729 ( .A(p_input[2887]), .Z(n9853) );
  XOR U9730 ( .A(n10012), .B(n10013), .Z(n10008) );
  AND U9731 ( .A(n10014), .B(n10015), .Z(n10013) );
  XNOR U9732 ( .A(p_input[2902]), .B(n10012), .Z(n10015) );
  XNOR U9733 ( .A(n10012), .B(n9862), .Z(n10014) );
  IV U9734 ( .A(p_input[2886]), .Z(n9862) );
  XOR U9735 ( .A(n10016), .B(n10017), .Z(n10012) );
  AND U9736 ( .A(n10018), .B(n10019), .Z(n10017) );
  XNOR U9737 ( .A(p_input[2901]), .B(n10016), .Z(n10019) );
  XNOR U9738 ( .A(n10016), .B(n9871), .Z(n10018) );
  IV U9739 ( .A(p_input[2885]), .Z(n9871) );
  XOR U9740 ( .A(n10020), .B(n10021), .Z(n10016) );
  AND U9741 ( .A(n10022), .B(n10023), .Z(n10021) );
  XNOR U9742 ( .A(p_input[2900]), .B(n10020), .Z(n10023) );
  XNOR U9743 ( .A(n10020), .B(n9880), .Z(n10022) );
  IV U9744 ( .A(p_input[2884]), .Z(n9880) );
  XOR U9745 ( .A(n10024), .B(n10025), .Z(n10020) );
  AND U9746 ( .A(n10026), .B(n10027), .Z(n10025) );
  XNOR U9747 ( .A(p_input[2899]), .B(n10024), .Z(n10027) );
  XNOR U9748 ( .A(n10024), .B(n9889), .Z(n10026) );
  IV U9749 ( .A(p_input[2883]), .Z(n9889) );
  XOR U9750 ( .A(n10028), .B(n10029), .Z(n10024) );
  AND U9751 ( .A(n10030), .B(n10031), .Z(n10029) );
  XNOR U9752 ( .A(p_input[2898]), .B(n10028), .Z(n10031) );
  XNOR U9753 ( .A(n10028), .B(n9898), .Z(n10030) );
  IV U9754 ( .A(p_input[2882]), .Z(n9898) );
  XNOR U9755 ( .A(n10032), .B(n10033), .Z(n10028) );
  AND U9756 ( .A(n10034), .B(n10035), .Z(n10033) );
  XOR U9757 ( .A(p_input[2897]), .B(n10032), .Z(n10035) );
  XNOR U9758 ( .A(p_input[2881]), .B(n10032), .Z(n10034) );
  AND U9759 ( .A(p_input[2896]), .B(n10036), .Z(n10032) );
  IV U9760 ( .A(p_input[2880]), .Z(n10036) );
  XOR U9761 ( .A(n10037), .B(n10038), .Z(n9595) );
  AND U9762 ( .A(n420), .B(n10039), .Z(n10038) );
  XNOR U9763 ( .A(n10040), .B(n10037), .Z(n10039) );
  XOR U9764 ( .A(n10041), .B(n10042), .Z(n420) );
  AND U9765 ( .A(n10043), .B(n10044), .Z(n10042) );
  XNOR U9766 ( .A(n9606), .B(n10041), .Z(n10044) );
  AND U9767 ( .A(p_input[2879]), .B(p_input[2863]), .Z(n9606) );
  XOR U9768 ( .A(n10041), .B(n9605), .Z(n10043) );
  AND U9769 ( .A(p_input[2831]), .B(p_input[2847]), .Z(n9605) );
  XOR U9770 ( .A(n10045), .B(n10046), .Z(n10041) );
  AND U9771 ( .A(n10047), .B(n10048), .Z(n10046) );
  XOR U9772 ( .A(n10045), .B(n9618), .Z(n10048) );
  XNOR U9773 ( .A(p_input[2862]), .B(n10049), .Z(n9618) );
  AND U9774 ( .A(n247), .B(n10050), .Z(n10049) );
  XOR U9775 ( .A(p_input[2878]), .B(p_input[2862]), .Z(n10050) );
  XNOR U9776 ( .A(n9615), .B(n10045), .Z(n10047) );
  XOR U9777 ( .A(n10051), .B(n10052), .Z(n9615) );
  AND U9778 ( .A(n244), .B(n10053), .Z(n10052) );
  XOR U9779 ( .A(p_input[2846]), .B(p_input[2830]), .Z(n10053) );
  XOR U9780 ( .A(n10054), .B(n10055), .Z(n10045) );
  AND U9781 ( .A(n10056), .B(n10057), .Z(n10055) );
  XOR U9782 ( .A(n10054), .B(n9630), .Z(n10057) );
  XNOR U9783 ( .A(p_input[2861]), .B(n10058), .Z(n9630) );
  AND U9784 ( .A(n247), .B(n10059), .Z(n10058) );
  XOR U9785 ( .A(p_input[2877]), .B(p_input[2861]), .Z(n10059) );
  XNOR U9786 ( .A(n9627), .B(n10054), .Z(n10056) );
  XOR U9787 ( .A(n10060), .B(n10061), .Z(n9627) );
  AND U9788 ( .A(n244), .B(n10062), .Z(n10061) );
  XOR U9789 ( .A(p_input[2845]), .B(p_input[2829]), .Z(n10062) );
  XOR U9790 ( .A(n10063), .B(n10064), .Z(n10054) );
  AND U9791 ( .A(n10065), .B(n10066), .Z(n10064) );
  XOR U9792 ( .A(n10063), .B(n9642), .Z(n10066) );
  XNOR U9793 ( .A(p_input[2860]), .B(n10067), .Z(n9642) );
  AND U9794 ( .A(n247), .B(n10068), .Z(n10067) );
  XOR U9795 ( .A(p_input[2876]), .B(p_input[2860]), .Z(n10068) );
  XNOR U9796 ( .A(n9639), .B(n10063), .Z(n10065) );
  XOR U9797 ( .A(n10069), .B(n10070), .Z(n9639) );
  AND U9798 ( .A(n244), .B(n10071), .Z(n10070) );
  XOR U9799 ( .A(p_input[2844]), .B(p_input[2828]), .Z(n10071) );
  XOR U9800 ( .A(n10072), .B(n10073), .Z(n10063) );
  AND U9801 ( .A(n10074), .B(n10075), .Z(n10073) );
  XOR U9802 ( .A(n10072), .B(n9654), .Z(n10075) );
  XNOR U9803 ( .A(p_input[2859]), .B(n10076), .Z(n9654) );
  AND U9804 ( .A(n247), .B(n10077), .Z(n10076) );
  XOR U9805 ( .A(p_input[2875]), .B(p_input[2859]), .Z(n10077) );
  XNOR U9806 ( .A(n9651), .B(n10072), .Z(n10074) );
  XOR U9807 ( .A(n10078), .B(n10079), .Z(n9651) );
  AND U9808 ( .A(n244), .B(n10080), .Z(n10079) );
  XOR U9809 ( .A(p_input[2843]), .B(p_input[2827]), .Z(n10080) );
  XOR U9810 ( .A(n10081), .B(n10082), .Z(n10072) );
  AND U9811 ( .A(n10083), .B(n10084), .Z(n10082) );
  XOR U9812 ( .A(n10081), .B(n9666), .Z(n10084) );
  XNOR U9813 ( .A(p_input[2858]), .B(n10085), .Z(n9666) );
  AND U9814 ( .A(n247), .B(n10086), .Z(n10085) );
  XOR U9815 ( .A(p_input[2874]), .B(p_input[2858]), .Z(n10086) );
  XNOR U9816 ( .A(n9663), .B(n10081), .Z(n10083) );
  XOR U9817 ( .A(n10087), .B(n10088), .Z(n9663) );
  AND U9818 ( .A(n244), .B(n10089), .Z(n10088) );
  XOR U9819 ( .A(p_input[2842]), .B(p_input[2826]), .Z(n10089) );
  XOR U9820 ( .A(n10090), .B(n10091), .Z(n10081) );
  AND U9821 ( .A(n10092), .B(n10093), .Z(n10091) );
  XOR U9822 ( .A(n10090), .B(n9678), .Z(n10093) );
  XNOR U9823 ( .A(p_input[2857]), .B(n10094), .Z(n9678) );
  AND U9824 ( .A(n247), .B(n10095), .Z(n10094) );
  XOR U9825 ( .A(p_input[2873]), .B(p_input[2857]), .Z(n10095) );
  XNOR U9826 ( .A(n9675), .B(n10090), .Z(n10092) );
  XOR U9827 ( .A(n10096), .B(n10097), .Z(n9675) );
  AND U9828 ( .A(n244), .B(n10098), .Z(n10097) );
  XOR U9829 ( .A(p_input[2841]), .B(p_input[2825]), .Z(n10098) );
  XOR U9830 ( .A(n10099), .B(n10100), .Z(n10090) );
  AND U9831 ( .A(n10101), .B(n10102), .Z(n10100) );
  XOR U9832 ( .A(n10099), .B(n9690), .Z(n10102) );
  XNOR U9833 ( .A(p_input[2856]), .B(n10103), .Z(n9690) );
  AND U9834 ( .A(n247), .B(n10104), .Z(n10103) );
  XOR U9835 ( .A(p_input[2872]), .B(p_input[2856]), .Z(n10104) );
  XNOR U9836 ( .A(n9687), .B(n10099), .Z(n10101) );
  XOR U9837 ( .A(n10105), .B(n10106), .Z(n9687) );
  AND U9838 ( .A(n244), .B(n10107), .Z(n10106) );
  XOR U9839 ( .A(p_input[2840]), .B(p_input[2824]), .Z(n10107) );
  XOR U9840 ( .A(n10108), .B(n10109), .Z(n10099) );
  AND U9841 ( .A(n10110), .B(n10111), .Z(n10109) );
  XOR U9842 ( .A(n10108), .B(n9702), .Z(n10111) );
  XNOR U9843 ( .A(p_input[2855]), .B(n10112), .Z(n9702) );
  AND U9844 ( .A(n247), .B(n10113), .Z(n10112) );
  XOR U9845 ( .A(p_input[2871]), .B(p_input[2855]), .Z(n10113) );
  XNOR U9846 ( .A(n9699), .B(n10108), .Z(n10110) );
  XOR U9847 ( .A(n10114), .B(n10115), .Z(n9699) );
  AND U9848 ( .A(n244), .B(n10116), .Z(n10115) );
  XOR U9849 ( .A(p_input[2839]), .B(p_input[2823]), .Z(n10116) );
  XOR U9850 ( .A(n10117), .B(n10118), .Z(n10108) );
  AND U9851 ( .A(n10119), .B(n10120), .Z(n10118) );
  XOR U9852 ( .A(n10117), .B(n9714), .Z(n10120) );
  XNOR U9853 ( .A(p_input[2854]), .B(n10121), .Z(n9714) );
  AND U9854 ( .A(n247), .B(n10122), .Z(n10121) );
  XOR U9855 ( .A(p_input[2870]), .B(p_input[2854]), .Z(n10122) );
  XNOR U9856 ( .A(n9711), .B(n10117), .Z(n10119) );
  XOR U9857 ( .A(n10123), .B(n10124), .Z(n9711) );
  AND U9858 ( .A(n244), .B(n10125), .Z(n10124) );
  XOR U9859 ( .A(p_input[2838]), .B(p_input[2822]), .Z(n10125) );
  XOR U9860 ( .A(n10126), .B(n10127), .Z(n10117) );
  AND U9861 ( .A(n10128), .B(n10129), .Z(n10127) );
  XOR U9862 ( .A(n10126), .B(n9726), .Z(n10129) );
  XNOR U9863 ( .A(p_input[2853]), .B(n10130), .Z(n9726) );
  AND U9864 ( .A(n247), .B(n10131), .Z(n10130) );
  XOR U9865 ( .A(p_input[2869]), .B(p_input[2853]), .Z(n10131) );
  XNOR U9866 ( .A(n9723), .B(n10126), .Z(n10128) );
  XOR U9867 ( .A(n10132), .B(n10133), .Z(n9723) );
  AND U9868 ( .A(n244), .B(n10134), .Z(n10133) );
  XOR U9869 ( .A(p_input[2837]), .B(p_input[2821]), .Z(n10134) );
  XOR U9870 ( .A(n10135), .B(n10136), .Z(n10126) );
  AND U9871 ( .A(n10137), .B(n10138), .Z(n10136) );
  XOR U9872 ( .A(n10135), .B(n9738), .Z(n10138) );
  XNOR U9873 ( .A(p_input[2852]), .B(n10139), .Z(n9738) );
  AND U9874 ( .A(n247), .B(n10140), .Z(n10139) );
  XOR U9875 ( .A(p_input[2868]), .B(p_input[2852]), .Z(n10140) );
  XNOR U9876 ( .A(n9735), .B(n10135), .Z(n10137) );
  XOR U9877 ( .A(n10141), .B(n10142), .Z(n9735) );
  AND U9878 ( .A(n244), .B(n10143), .Z(n10142) );
  XOR U9879 ( .A(p_input[2836]), .B(p_input[2820]), .Z(n10143) );
  XOR U9880 ( .A(n10144), .B(n10145), .Z(n10135) );
  AND U9881 ( .A(n10146), .B(n10147), .Z(n10145) );
  XOR U9882 ( .A(n10144), .B(n9750), .Z(n10147) );
  XNOR U9883 ( .A(p_input[2851]), .B(n10148), .Z(n9750) );
  AND U9884 ( .A(n247), .B(n10149), .Z(n10148) );
  XOR U9885 ( .A(p_input[2867]), .B(p_input[2851]), .Z(n10149) );
  XNOR U9886 ( .A(n9747), .B(n10144), .Z(n10146) );
  XOR U9887 ( .A(n10150), .B(n10151), .Z(n9747) );
  AND U9888 ( .A(n244), .B(n10152), .Z(n10151) );
  XOR U9889 ( .A(p_input[2835]), .B(p_input[2819]), .Z(n10152) );
  XOR U9890 ( .A(n10153), .B(n10154), .Z(n10144) );
  AND U9891 ( .A(n10155), .B(n10156), .Z(n10154) );
  XOR U9892 ( .A(n10153), .B(n9762), .Z(n10156) );
  XNOR U9893 ( .A(p_input[2850]), .B(n10157), .Z(n9762) );
  AND U9894 ( .A(n247), .B(n10158), .Z(n10157) );
  XOR U9895 ( .A(p_input[2866]), .B(p_input[2850]), .Z(n10158) );
  XNOR U9896 ( .A(n9759), .B(n10153), .Z(n10155) );
  XOR U9897 ( .A(n10159), .B(n10160), .Z(n9759) );
  AND U9898 ( .A(n244), .B(n10161), .Z(n10160) );
  XOR U9899 ( .A(p_input[2834]), .B(p_input[2818]), .Z(n10161) );
  XOR U9900 ( .A(n10162), .B(n10163), .Z(n10153) );
  AND U9901 ( .A(n10164), .B(n10165), .Z(n10163) );
  XNOR U9902 ( .A(n10166), .B(n9775), .Z(n10165) );
  XNOR U9903 ( .A(p_input[2849]), .B(n10167), .Z(n9775) );
  AND U9904 ( .A(n247), .B(n10168), .Z(n10167) );
  XNOR U9905 ( .A(p_input[2865]), .B(n10169), .Z(n10168) );
  IV U9906 ( .A(p_input[2849]), .Z(n10169) );
  XNOR U9907 ( .A(n9772), .B(n10162), .Z(n10164) );
  XNOR U9908 ( .A(p_input[2817]), .B(n10170), .Z(n9772) );
  AND U9909 ( .A(n244), .B(n10171), .Z(n10170) );
  XOR U9910 ( .A(p_input[2833]), .B(p_input[2817]), .Z(n10171) );
  IV U9911 ( .A(n10166), .Z(n10162) );
  AND U9912 ( .A(n10037), .B(n10040), .Z(n10166) );
  XOR U9913 ( .A(p_input[2848]), .B(n10172), .Z(n10040) );
  AND U9914 ( .A(n247), .B(n10173), .Z(n10172) );
  XOR U9915 ( .A(p_input[2864]), .B(p_input[2848]), .Z(n10173) );
  XOR U9916 ( .A(n10174), .B(n10175), .Z(n247) );
  AND U9917 ( .A(n10176), .B(n10177), .Z(n10175) );
  XNOR U9918 ( .A(p_input[2879]), .B(n10174), .Z(n10177) );
  XOR U9919 ( .A(n10174), .B(p_input[2863]), .Z(n10176) );
  XOR U9920 ( .A(n10178), .B(n10179), .Z(n10174) );
  AND U9921 ( .A(n10180), .B(n10181), .Z(n10179) );
  XNOR U9922 ( .A(p_input[2878]), .B(n10178), .Z(n10181) );
  XOR U9923 ( .A(n10178), .B(p_input[2862]), .Z(n10180) );
  XOR U9924 ( .A(n10182), .B(n10183), .Z(n10178) );
  AND U9925 ( .A(n10184), .B(n10185), .Z(n10183) );
  XNOR U9926 ( .A(p_input[2877]), .B(n10182), .Z(n10185) );
  XOR U9927 ( .A(n10182), .B(p_input[2861]), .Z(n10184) );
  XOR U9928 ( .A(n10186), .B(n10187), .Z(n10182) );
  AND U9929 ( .A(n10188), .B(n10189), .Z(n10187) );
  XNOR U9930 ( .A(p_input[2876]), .B(n10186), .Z(n10189) );
  XOR U9931 ( .A(n10186), .B(p_input[2860]), .Z(n10188) );
  XOR U9932 ( .A(n10190), .B(n10191), .Z(n10186) );
  AND U9933 ( .A(n10192), .B(n10193), .Z(n10191) );
  XNOR U9934 ( .A(p_input[2875]), .B(n10190), .Z(n10193) );
  XOR U9935 ( .A(n10190), .B(p_input[2859]), .Z(n10192) );
  XOR U9936 ( .A(n10194), .B(n10195), .Z(n10190) );
  AND U9937 ( .A(n10196), .B(n10197), .Z(n10195) );
  XNOR U9938 ( .A(p_input[2874]), .B(n10194), .Z(n10197) );
  XOR U9939 ( .A(n10194), .B(p_input[2858]), .Z(n10196) );
  XOR U9940 ( .A(n10198), .B(n10199), .Z(n10194) );
  AND U9941 ( .A(n10200), .B(n10201), .Z(n10199) );
  XNOR U9942 ( .A(p_input[2873]), .B(n10198), .Z(n10201) );
  XOR U9943 ( .A(n10198), .B(p_input[2857]), .Z(n10200) );
  XOR U9944 ( .A(n10202), .B(n10203), .Z(n10198) );
  AND U9945 ( .A(n10204), .B(n10205), .Z(n10203) );
  XNOR U9946 ( .A(p_input[2872]), .B(n10202), .Z(n10205) );
  XOR U9947 ( .A(n10202), .B(p_input[2856]), .Z(n10204) );
  XOR U9948 ( .A(n10206), .B(n10207), .Z(n10202) );
  AND U9949 ( .A(n10208), .B(n10209), .Z(n10207) );
  XNOR U9950 ( .A(p_input[2871]), .B(n10206), .Z(n10209) );
  XOR U9951 ( .A(n10206), .B(p_input[2855]), .Z(n10208) );
  XOR U9952 ( .A(n10210), .B(n10211), .Z(n10206) );
  AND U9953 ( .A(n10212), .B(n10213), .Z(n10211) );
  XNOR U9954 ( .A(p_input[2870]), .B(n10210), .Z(n10213) );
  XOR U9955 ( .A(n10210), .B(p_input[2854]), .Z(n10212) );
  XOR U9956 ( .A(n10214), .B(n10215), .Z(n10210) );
  AND U9957 ( .A(n10216), .B(n10217), .Z(n10215) );
  XNOR U9958 ( .A(p_input[2869]), .B(n10214), .Z(n10217) );
  XOR U9959 ( .A(n10214), .B(p_input[2853]), .Z(n10216) );
  XOR U9960 ( .A(n10218), .B(n10219), .Z(n10214) );
  AND U9961 ( .A(n10220), .B(n10221), .Z(n10219) );
  XNOR U9962 ( .A(p_input[2868]), .B(n10218), .Z(n10221) );
  XOR U9963 ( .A(n10218), .B(p_input[2852]), .Z(n10220) );
  XOR U9964 ( .A(n10222), .B(n10223), .Z(n10218) );
  AND U9965 ( .A(n10224), .B(n10225), .Z(n10223) );
  XNOR U9966 ( .A(p_input[2867]), .B(n10222), .Z(n10225) );
  XOR U9967 ( .A(n10222), .B(p_input[2851]), .Z(n10224) );
  XOR U9968 ( .A(n10226), .B(n10227), .Z(n10222) );
  AND U9969 ( .A(n10228), .B(n10229), .Z(n10227) );
  XNOR U9970 ( .A(p_input[2866]), .B(n10226), .Z(n10229) );
  XOR U9971 ( .A(n10226), .B(p_input[2850]), .Z(n10228) );
  XNOR U9972 ( .A(n10230), .B(n10231), .Z(n10226) );
  AND U9973 ( .A(n10232), .B(n10233), .Z(n10231) );
  XOR U9974 ( .A(p_input[2865]), .B(n10230), .Z(n10233) );
  XNOR U9975 ( .A(p_input[2849]), .B(n10230), .Z(n10232) );
  AND U9976 ( .A(p_input[2864]), .B(n10234), .Z(n10230) );
  IV U9977 ( .A(p_input[2848]), .Z(n10234) );
  XNOR U9978 ( .A(p_input[2816]), .B(n10235), .Z(n10037) );
  AND U9979 ( .A(n244), .B(n10236), .Z(n10235) );
  XOR U9980 ( .A(p_input[2832]), .B(p_input[2816]), .Z(n10236) );
  XOR U9981 ( .A(n10237), .B(n10238), .Z(n244) );
  AND U9982 ( .A(n10239), .B(n10240), .Z(n10238) );
  XNOR U9983 ( .A(p_input[2847]), .B(n10237), .Z(n10240) );
  XOR U9984 ( .A(n10237), .B(p_input[2831]), .Z(n10239) );
  XOR U9985 ( .A(n10241), .B(n10242), .Z(n10237) );
  AND U9986 ( .A(n10243), .B(n10244), .Z(n10242) );
  XNOR U9987 ( .A(p_input[2846]), .B(n10241), .Z(n10244) );
  XNOR U9988 ( .A(n10241), .B(n10051), .Z(n10243) );
  IV U9989 ( .A(p_input[2830]), .Z(n10051) );
  XOR U9990 ( .A(n10245), .B(n10246), .Z(n10241) );
  AND U9991 ( .A(n10247), .B(n10248), .Z(n10246) );
  XNOR U9992 ( .A(p_input[2845]), .B(n10245), .Z(n10248) );
  XNOR U9993 ( .A(n10245), .B(n10060), .Z(n10247) );
  IV U9994 ( .A(p_input[2829]), .Z(n10060) );
  XOR U9995 ( .A(n10249), .B(n10250), .Z(n10245) );
  AND U9996 ( .A(n10251), .B(n10252), .Z(n10250) );
  XNOR U9997 ( .A(p_input[2844]), .B(n10249), .Z(n10252) );
  XNOR U9998 ( .A(n10249), .B(n10069), .Z(n10251) );
  IV U9999 ( .A(p_input[2828]), .Z(n10069) );
  XOR U10000 ( .A(n10253), .B(n10254), .Z(n10249) );
  AND U10001 ( .A(n10255), .B(n10256), .Z(n10254) );
  XNOR U10002 ( .A(p_input[2843]), .B(n10253), .Z(n10256) );
  XNOR U10003 ( .A(n10253), .B(n10078), .Z(n10255) );
  IV U10004 ( .A(p_input[2827]), .Z(n10078) );
  XOR U10005 ( .A(n10257), .B(n10258), .Z(n10253) );
  AND U10006 ( .A(n10259), .B(n10260), .Z(n10258) );
  XNOR U10007 ( .A(p_input[2842]), .B(n10257), .Z(n10260) );
  XNOR U10008 ( .A(n10257), .B(n10087), .Z(n10259) );
  IV U10009 ( .A(p_input[2826]), .Z(n10087) );
  XOR U10010 ( .A(n10261), .B(n10262), .Z(n10257) );
  AND U10011 ( .A(n10263), .B(n10264), .Z(n10262) );
  XNOR U10012 ( .A(p_input[2841]), .B(n10261), .Z(n10264) );
  XNOR U10013 ( .A(n10261), .B(n10096), .Z(n10263) );
  IV U10014 ( .A(p_input[2825]), .Z(n10096) );
  XOR U10015 ( .A(n10265), .B(n10266), .Z(n10261) );
  AND U10016 ( .A(n10267), .B(n10268), .Z(n10266) );
  XNOR U10017 ( .A(p_input[2840]), .B(n10265), .Z(n10268) );
  XNOR U10018 ( .A(n10265), .B(n10105), .Z(n10267) );
  IV U10019 ( .A(p_input[2824]), .Z(n10105) );
  XOR U10020 ( .A(n10269), .B(n10270), .Z(n10265) );
  AND U10021 ( .A(n10271), .B(n10272), .Z(n10270) );
  XNOR U10022 ( .A(p_input[2839]), .B(n10269), .Z(n10272) );
  XNOR U10023 ( .A(n10269), .B(n10114), .Z(n10271) );
  IV U10024 ( .A(p_input[2823]), .Z(n10114) );
  XOR U10025 ( .A(n10273), .B(n10274), .Z(n10269) );
  AND U10026 ( .A(n10275), .B(n10276), .Z(n10274) );
  XNOR U10027 ( .A(p_input[2838]), .B(n10273), .Z(n10276) );
  XNOR U10028 ( .A(n10273), .B(n10123), .Z(n10275) );
  IV U10029 ( .A(p_input[2822]), .Z(n10123) );
  XOR U10030 ( .A(n10277), .B(n10278), .Z(n10273) );
  AND U10031 ( .A(n10279), .B(n10280), .Z(n10278) );
  XNOR U10032 ( .A(p_input[2837]), .B(n10277), .Z(n10280) );
  XNOR U10033 ( .A(n10277), .B(n10132), .Z(n10279) );
  IV U10034 ( .A(p_input[2821]), .Z(n10132) );
  XOR U10035 ( .A(n10281), .B(n10282), .Z(n10277) );
  AND U10036 ( .A(n10283), .B(n10284), .Z(n10282) );
  XNOR U10037 ( .A(p_input[2836]), .B(n10281), .Z(n10284) );
  XNOR U10038 ( .A(n10281), .B(n10141), .Z(n10283) );
  IV U10039 ( .A(p_input[2820]), .Z(n10141) );
  XOR U10040 ( .A(n10285), .B(n10286), .Z(n10281) );
  AND U10041 ( .A(n10287), .B(n10288), .Z(n10286) );
  XNOR U10042 ( .A(p_input[2835]), .B(n10285), .Z(n10288) );
  XNOR U10043 ( .A(n10285), .B(n10150), .Z(n10287) );
  IV U10044 ( .A(p_input[2819]), .Z(n10150) );
  XOR U10045 ( .A(n10289), .B(n10290), .Z(n10285) );
  AND U10046 ( .A(n10291), .B(n10292), .Z(n10290) );
  XNOR U10047 ( .A(p_input[2834]), .B(n10289), .Z(n10292) );
  XNOR U10048 ( .A(n10289), .B(n10159), .Z(n10291) );
  IV U10049 ( .A(p_input[2818]), .Z(n10159) );
  XNOR U10050 ( .A(n10293), .B(n10294), .Z(n10289) );
  AND U10051 ( .A(n10295), .B(n10296), .Z(n10294) );
  XOR U10052 ( .A(p_input[2833]), .B(n10293), .Z(n10296) );
  XNOR U10053 ( .A(p_input[2817]), .B(n10293), .Z(n10295) );
  AND U10054 ( .A(p_input[2832]), .B(n10297), .Z(n10293) );
  IV U10055 ( .A(p_input[2816]), .Z(n10297) );
  XOR U10056 ( .A(n10298), .B(n10299), .Z(n8525) );
  AND U10057 ( .A(n929), .B(n10300), .Z(n10299) );
  XNOR U10058 ( .A(n10301), .B(n10298), .Z(n10300) );
  XOR U10059 ( .A(n10302), .B(n10303), .Z(n929) );
  AND U10060 ( .A(n10304), .B(n10305), .Z(n10303) );
  XNOR U10061 ( .A(n8540), .B(n10302), .Z(n10305) );
  AND U10062 ( .A(n10306), .B(n10307), .Z(n8540) );
  XNOR U10063 ( .A(n10302), .B(n8537), .Z(n10304) );
  IV U10064 ( .A(n10308), .Z(n8537) );
  AND U10065 ( .A(n10309), .B(n10310), .Z(n10308) );
  XOR U10066 ( .A(n10311), .B(n10312), .Z(n10302) );
  AND U10067 ( .A(n10313), .B(n10314), .Z(n10312) );
  XOR U10068 ( .A(n10311), .B(n8552), .Z(n10314) );
  XOR U10069 ( .A(n10315), .B(n10316), .Z(n8552) );
  AND U10070 ( .A(n767), .B(n10317), .Z(n10316) );
  XOR U10071 ( .A(n10318), .B(n10315), .Z(n10317) );
  XNOR U10072 ( .A(n8549), .B(n10311), .Z(n10313) );
  XOR U10073 ( .A(n10319), .B(n10320), .Z(n8549) );
  AND U10074 ( .A(n764), .B(n10321), .Z(n10320) );
  XOR U10075 ( .A(n10322), .B(n10319), .Z(n10321) );
  XOR U10076 ( .A(n10323), .B(n10324), .Z(n10311) );
  AND U10077 ( .A(n10325), .B(n10326), .Z(n10324) );
  XOR U10078 ( .A(n10323), .B(n8564), .Z(n10326) );
  XOR U10079 ( .A(n10327), .B(n10328), .Z(n8564) );
  AND U10080 ( .A(n767), .B(n10329), .Z(n10328) );
  XOR U10081 ( .A(n10330), .B(n10327), .Z(n10329) );
  XNOR U10082 ( .A(n8561), .B(n10323), .Z(n10325) );
  XOR U10083 ( .A(n10331), .B(n10332), .Z(n8561) );
  AND U10084 ( .A(n764), .B(n10333), .Z(n10332) );
  XOR U10085 ( .A(n10334), .B(n10331), .Z(n10333) );
  XOR U10086 ( .A(n10335), .B(n10336), .Z(n10323) );
  AND U10087 ( .A(n10337), .B(n10338), .Z(n10336) );
  XOR U10088 ( .A(n10335), .B(n8576), .Z(n10338) );
  XOR U10089 ( .A(n10339), .B(n10340), .Z(n8576) );
  AND U10090 ( .A(n767), .B(n10341), .Z(n10340) );
  XOR U10091 ( .A(n10342), .B(n10339), .Z(n10341) );
  XNOR U10092 ( .A(n8573), .B(n10335), .Z(n10337) );
  XOR U10093 ( .A(n10343), .B(n10344), .Z(n8573) );
  AND U10094 ( .A(n764), .B(n10345), .Z(n10344) );
  XOR U10095 ( .A(n10346), .B(n10343), .Z(n10345) );
  XOR U10096 ( .A(n10347), .B(n10348), .Z(n10335) );
  AND U10097 ( .A(n10349), .B(n10350), .Z(n10348) );
  XOR U10098 ( .A(n10347), .B(n8588), .Z(n10350) );
  XOR U10099 ( .A(n10351), .B(n10352), .Z(n8588) );
  AND U10100 ( .A(n767), .B(n10353), .Z(n10352) );
  XOR U10101 ( .A(n10354), .B(n10351), .Z(n10353) );
  XNOR U10102 ( .A(n8585), .B(n10347), .Z(n10349) );
  XOR U10103 ( .A(n10355), .B(n10356), .Z(n8585) );
  AND U10104 ( .A(n764), .B(n10357), .Z(n10356) );
  XOR U10105 ( .A(n10358), .B(n10355), .Z(n10357) );
  XOR U10106 ( .A(n10359), .B(n10360), .Z(n10347) );
  AND U10107 ( .A(n10361), .B(n10362), .Z(n10360) );
  XOR U10108 ( .A(n10359), .B(n8600), .Z(n10362) );
  XOR U10109 ( .A(n10363), .B(n10364), .Z(n8600) );
  AND U10110 ( .A(n767), .B(n10365), .Z(n10364) );
  XOR U10111 ( .A(n10366), .B(n10363), .Z(n10365) );
  XNOR U10112 ( .A(n8597), .B(n10359), .Z(n10361) );
  XOR U10113 ( .A(n10367), .B(n10368), .Z(n8597) );
  AND U10114 ( .A(n764), .B(n10369), .Z(n10368) );
  XOR U10115 ( .A(n10370), .B(n10367), .Z(n10369) );
  XOR U10116 ( .A(n10371), .B(n10372), .Z(n10359) );
  AND U10117 ( .A(n10373), .B(n10374), .Z(n10372) );
  XOR U10118 ( .A(n10371), .B(n8612), .Z(n10374) );
  XOR U10119 ( .A(n10375), .B(n10376), .Z(n8612) );
  AND U10120 ( .A(n767), .B(n10377), .Z(n10376) );
  XOR U10121 ( .A(n10378), .B(n10375), .Z(n10377) );
  XNOR U10122 ( .A(n8609), .B(n10371), .Z(n10373) );
  XOR U10123 ( .A(n10379), .B(n10380), .Z(n8609) );
  AND U10124 ( .A(n764), .B(n10381), .Z(n10380) );
  XOR U10125 ( .A(n10382), .B(n10379), .Z(n10381) );
  XOR U10126 ( .A(n10383), .B(n10384), .Z(n10371) );
  AND U10127 ( .A(n10385), .B(n10386), .Z(n10384) );
  XOR U10128 ( .A(n10383), .B(n8624), .Z(n10386) );
  XOR U10129 ( .A(n10387), .B(n10388), .Z(n8624) );
  AND U10130 ( .A(n767), .B(n10389), .Z(n10388) );
  XOR U10131 ( .A(n10390), .B(n10387), .Z(n10389) );
  XNOR U10132 ( .A(n8621), .B(n10383), .Z(n10385) );
  XOR U10133 ( .A(n10391), .B(n10392), .Z(n8621) );
  AND U10134 ( .A(n764), .B(n10393), .Z(n10392) );
  XOR U10135 ( .A(n10394), .B(n10391), .Z(n10393) );
  XOR U10136 ( .A(n10395), .B(n10396), .Z(n10383) );
  AND U10137 ( .A(n10397), .B(n10398), .Z(n10396) );
  XOR U10138 ( .A(n10395), .B(n8636), .Z(n10398) );
  XOR U10139 ( .A(n10399), .B(n10400), .Z(n8636) );
  AND U10140 ( .A(n767), .B(n10401), .Z(n10400) );
  XOR U10141 ( .A(n10402), .B(n10399), .Z(n10401) );
  XNOR U10142 ( .A(n8633), .B(n10395), .Z(n10397) );
  XOR U10143 ( .A(n10403), .B(n10404), .Z(n8633) );
  AND U10144 ( .A(n764), .B(n10405), .Z(n10404) );
  XOR U10145 ( .A(n10406), .B(n10403), .Z(n10405) );
  XOR U10146 ( .A(n10407), .B(n10408), .Z(n10395) );
  AND U10147 ( .A(n10409), .B(n10410), .Z(n10408) );
  XOR U10148 ( .A(n10407), .B(n8648), .Z(n10410) );
  XOR U10149 ( .A(n10411), .B(n10412), .Z(n8648) );
  AND U10150 ( .A(n767), .B(n10413), .Z(n10412) );
  XOR U10151 ( .A(n10414), .B(n10411), .Z(n10413) );
  XNOR U10152 ( .A(n8645), .B(n10407), .Z(n10409) );
  XOR U10153 ( .A(n10415), .B(n10416), .Z(n8645) );
  AND U10154 ( .A(n764), .B(n10417), .Z(n10416) );
  XOR U10155 ( .A(n10418), .B(n10415), .Z(n10417) );
  XOR U10156 ( .A(n10419), .B(n10420), .Z(n10407) );
  AND U10157 ( .A(n10421), .B(n10422), .Z(n10420) );
  XOR U10158 ( .A(n10419), .B(n8660), .Z(n10422) );
  XOR U10159 ( .A(n10423), .B(n10424), .Z(n8660) );
  AND U10160 ( .A(n767), .B(n10425), .Z(n10424) );
  XOR U10161 ( .A(n10426), .B(n10423), .Z(n10425) );
  XNOR U10162 ( .A(n8657), .B(n10419), .Z(n10421) );
  XOR U10163 ( .A(n10427), .B(n10428), .Z(n8657) );
  AND U10164 ( .A(n764), .B(n10429), .Z(n10428) );
  XOR U10165 ( .A(n10430), .B(n10427), .Z(n10429) );
  XOR U10166 ( .A(n10431), .B(n10432), .Z(n10419) );
  AND U10167 ( .A(n10433), .B(n10434), .Z(n10432) );
  XOR U10168 ( .A(n10431), .B(n8672), .Z(n10434) );
  XOR U10169 ( .A(n10435), .B(n10436), .Z(n8672) );
  AND U10170 ( .A(n767), .B(n10437), .Z(n10436) );
  XOR U10171 ( .A(n10438), .B(n10435), .Z(n10437) );
  XNOR U10172 ( .A(n8669), .B(n10431), .Z(n10433) );
  XOR U10173 ( .A(n10439), .B(n10440), .Z(n8669) );
  AND U10174 ( .A(n764), .B(n10441), .Z(n10440) );
  XOR U10175 ( .A(n10442), .B(n10439), .Z(n10441) );
  XOR U10176 ( .A(n10443), .B(n10444), .Z(n10431) );
  AND U10177 ( .A(n10445), .B(n10446), .Z(n10444) );
  XOR U10178 ( .A(n10443), .B(n8684), .Z(n10446) );
  XOR U10179 ( .A(n10447), .B(n10448), .Z(n8684) );
  AND U10180 ( .A(n767), .B(n10449), .Z(n10448) );
  XOR U10181 ( .A(n10450), .B(n10447), .Z(n10449) );
  XNOR U10182 ( .A(n8681), .B(n10443), .Z(n10445) );
  XOR U10183 ( .A(n10451), .B(n10452), .Z(n8681) );
  AND U10184 ( .A(n764), .B(n10453), .Z(n10452) );
  XOR U10185 ( .A(n10454), .B(n10451), .Z(n10453) );
  XOR U10186 ( .A(n10455), .B(n10456), .Z(n10443) );
  AND U10187 ( .A(n10457), .B(n10458), .Z(n10456) );
  XOR U10188 ( .A(n10455), .B(n8696), .Z(n10458) );
  XOR U10189 ( .A(n10459), .B(n10460), .Z(n8696) );
  AND U10190 ( .A(n767), .B(n10461), .Z(n10460) );
  XOR U10191 ( .A(n10462), .B(n10459), .Z(n10461) );
  XNOR U10192 ( .A(n8693), .B(n10455), .Z(n10457) );
  XOR U10193 ( .A(n10463), .B(n10464), .Z(n8693) );
  AND U10194 ( .A(n764), .B(n10465), .Z(n10464) );
  XOR U10195 ( .A(n10466), .B(n10463), .Z(n10465) );
  XOR U10196 ( .A(n10467), .B(n10468), .Z(n10455) );
  AND U10197 ( .A(n10469), .B(n10470), .Z(n10468) );
  XNOR U10198 ( .A(n10471), .B(n8709), .Z(n10470) );
  XOR U10199 ( .A(n10472), .B(n10473), .Z(n8709) );
  AND U10200 ( .A(n767), .B(n10474), .Z(n10473) );
  XOR U10201 ( .A(n10472), .B(n10475), .Z(n10474) );
  XNOR U10202 ( .A(n8706), .B(n10467), .Z(n10469) );
  XOR U10203 ( .A(n10476), .B(n10477), .Z(n8706) );
  AND U10204 ( .A(n764), .B(n10478), .Z(n10477) );
  XOR U10205 ( .A(n10476), .B(n10479), .Z(n10478) );
  IV U10206 ( .A(n10471), .Z(n10467) );
  AND U10207 ( .A(n10298), .B(n10301), .Z(n10471) );
  XNOR U10208 ( .A(n10480), .B(n10481), .Z(n10301) );
  AND U10209 ( .A(n767), .B(n10482), .Z(n10481) );
  XNOR U10210 ( .A(n10483), .B(n10480), .Z(n10482) );
  XOR U10211 ( .A(n10484), .B(n10485), .Z(n767) );
  AND U10212 ( .A(n10486), .B(n10487), .Z(n10485) );
  XNOR U10213 ( .A(n10306), .B(n10484), .Z(n10487) );
  AND U10214 ( .A(n10488), .B(n10489), .Z(n10306) );
  XOR U10215 ( .A(n10484), .B(n10307), .Z(n10486) );
  AND U10216 ( .A(n10490), .B(n10491), .Z(n10307) );
  XOR U10217 ( .A(n10492), .B(n10493), .Z(n10484) );
  AND U10218 ( .A(n10494), .B(n10495), .Z(n10493) );
  XOR U10219 ( .A(n10492), .B(n10318), .Z(n10495) );
  XOR U10220 ( .A(n10496), .B(n10497), .Z(n10318) );
  AND U10221 ( .A(n431), .B(n10498), .Z(n10497) );
  XOR U10222 ( .A(n10499), .B(n10496), .Z(n10498) );
  XNOR U10223 ( .A(n10315), .B(n10492), .Z(n10494) );
  XOR U10224 ( .A(n10500), .B(n10501), .Z(n10315) );
  AND U10225 ( .A(n429), .B(n10502), .Z(n10501) );
  XOR U10226 ( .A(n10503), .B(n10500), .Z(n10502) );
  XOR U10227 ( .A(n10504), .B(n10505), .Z(n10492) );
  AND U10228 ( .A(n10506), .B(n10507), .Z(n10505) );
  XOR U10229 ( .A(n10504), .B(n10330), .Z(n10507) );
  XOR U10230 ( .A(n10508), .B(n10509), .Z(n10330) );
  AND U10231 ( .A(n431), .B(n10510), .Z(n10509) );
  XOR U10232 ( .A(n10511), .B(n10508), .Z(n10510) );
  XNOR U10233 ( .A(n10327), .B(n10504), .Z(n10506) );
  XOR U10234 ( .A(n10512), .B(n10513), .Z(n10327) );
  AND U10235 ( .A(n429), .B(n10514), .Z(n10513) );
  XOR U10236 ( .A(n10515), .B(n10512), .Z(n10514) );
  XOR U10237 ( .A(n10516), .B(n10517), .Z(n10504) );
  AND U10238 ( .A(n10518), .B(n10519), .Z(n10517) );
  XOR U10239 ( .A(n10516), .B(n10342), .Z(n10519) );
  XOR U10240 ( .A(n10520), .B(n10521), .Z(n10342) );
  AND U10241 ( .A(n431), .B(n10522), .Z(n10521) );
  XOR U10242 ( .A(n10523), .B(n10520), .Z(n10522) );
  XNOR U10243 ( .A(n10339), .B(n10516), .Z(n10518) );
  XOR U10244 ( .A(n10524), .B(n10525), .Z(n10339) );
  AND U10245 ( .A(n429), .B(n10526), .Z(n10525) );
  XOR U10246 ( .A(n10527), .B(n10524), .Z(n10526) );
  XOR U10247 ( .A(n10528), .B(n10529), .Z(n10516) );
  AND U10248 ( .A(n10530), .B(n10531), .Z(n10529) );
  XOR U10249 ( .A(n10528), .B(n10354), .Z(n10531) );
  XOR U10250 ( .A(n10532), .B(n10533), .Z(n10354) );
  AND U10251 ( .A(n431), .B(n10534), .Z(n10533) );
  XOR U10252 ( .A(n10535), .B(n10532), .Z(n10534) );
  XNOR U10253 ( .A(n10351), .B(n10528), .Z(n10530) );
  XOR U10254 ( .A(n10536), .B(n10537), .Z(n10351) );
  AND U10255 ( .A(n429), .B(n10538), .Z(n10537) );
  XOR U10256 ( .A(n10539), .B(n10536), .Z(n10538) );
  XOR U10257 ( .A(n10540), .B(n10541), .Z(n10528) );
  AND U10258 ( .A(n10542), .B(n10543), .Z(n10541) );
  XOR U10259 ( .A(n10540), .B(n10366), .Z(n10543) );
  XOR U10260 ( .A(n10544), .B(n10545), .Z(n10366) );
  AND U10261 ( .A(n431), .B(n10546), .Z(n10545) );
  XOR U10262 ( .A(n10547), .B(n10544), .Z(n10546) );
  XNOR U10263 ( .A(n10363), .B(n10540), .Z(n10542) );
  XOR U10264 ( .A(n10548), .B(n10549), .Z(n10363) );
  AND U10265 ( .A(n429), .B(n10550), .Z(n10549) );
  XOR U10266 ( .A(n10551), .B(n10548), .Z(n10550) );
  XOR U10267 ( .A(n10552), .B(n10553), .Z(n10540) );
  AND U10268 ( .A(n10554), .B(n10555), .Z(n10553) );
  XOR U10269 ( .A(n10552), .B(n10378), .Z(n10555) );
  XOR U10270 ( .A(n10556), .B(n10557), .Z(n10378) );
  AND U10271 ( .A(n431), .B(n10558), .Z(n10557) );
  XOR U10272 ( .A(n10559), .B(n10556), .Z(n10558) );
  XNOR U10273 ( .A(n10375), .B(n10552), .Z(n10554) );
  XOR U10274 ( .A(n10560), .B(n10561), .Z(n10375) );
  AND U10275 ( .A(n429), .B(n10562), .Z(n10561) );
  XOR U10276 ( .A(n10563), .B(n10560), .Z(n10562) );
  XOR U10277 ( .A(n10564), .B(n10565), .Z(n10552) );
  AND U10278 ( .A(n10566), .B(n10567), .Z(n10565) );
  XOR U10279 ( .A(n10564), .B(n10390), .Z(n10567) );
  XOR U10280 ( .A(n10568), .B(n10569), .Z(n10390) );
  AND U10281 ( .A(n431), .B(n10570), .Z(n10569) );
  XOR U10282 ( .A(n10571), .B(n10568), .Z(n10570) );
  XNOR U10283 ( .A(n10387), .B(n10564), .Z(n10566) );
  XOR U10284 ( .A(n10572), .B(n10573), .Z(n10387) );
  AND U10285 ( .A(n429), .B(n10574), .Z(n10573) );
  XOR U10286 ( .A(n10575), .B(n10572), .Z(n10574) );
  XOR U10287 ( .A(n10576), .B(n10577), .Z(n10564) );
  AND U10288 ( .A(n10578), .B(n10579), .Z(n10577) );
  XOR U10289 ( .A(n10576), .B(n10402), .Z(n10579) );
  XOR U10290 ( .A(n10580), .B(n10581), .Z(n10402) );
  AND U10291 ( .A(n431), .B(n10582), .Z(n10581) );
  XOR U10292 ( .A(n10583), .B(n10580), .Z(n10582) );
  XNOR U10293 ( .A(n10399), .B(n10576), .Z(n10578) );
  XOR U10294 ( .A(n10584), .B(n10585), .Z(n10399) );
  AND U10295 ( .A(n429), .B(n10586), .Z(n10585) );
  XOR U10296 ( .A(n10587), .B(n10584), .Z(n10586) );
  XOR U10297 ( .A(n10588), .B(n10589), .Z(n10576) );
  AND U10298 ( .A(n10590), .B(n10591), .Z(n10589) );
  XOR U10299 ( .A(n10588), .B(n10414), .Z(n10591) );
  XOR U10300 ( .A(n10592), .B(n10593), .Z(n10414) );
  AND U10301 ( .A(n431), .B(n10594), .Z(n10593) );
  XOR U10302 ( .A(n10595), .B(n10592), .Z(n10594) );
  XNOR U10303 ( .A(n10411), .B(n10588), .Z(n10590) );
  XOR U10304 ( .A(n10596), .B(n10597), .Z(n10411) );
  AND U10305 ( .A(n429), .B(n10598), .Z(n10597) );
  XOR U10306 ( .A(n10599), .B(n10596), .Z(n10598) );
  XOR U10307 ( .A(n10600), .B(n10601), .Z(n10588) );
  AND U10308 ( .A(n10602), .B(n10603), .Z(n10601) );
  XOR U10309 ( .A(n10600), .B(n10426), .Z(n10603) );
  XOR U10310 ( .A(n10604), .B(n10605), .Z(n10426) );
  AND U10311 ( .A(n431), .B(n10606), .Z(n10605) );
  XOR U10312 ( .A(n10607), .B(n10604), .Z(n10606) );
  XNOR U10313 ( .A(n10423), .B(n10600), .Z(n10602) );
  XOR U10314 ( .A(n10608), .B(n10609), .Z(n10423) );
  AND U10315 ( .A(n429), .B(n10610), .Z(n10609) );
  XOR U10316 ( .A(n10611), .B(n10608), .Z(n10610) );
  XOR U10317 ( .A(n10612), .B(n10613), .Z(n10600) );
  AND U10318 ( .A(n10614), .B(n10615), .Z(n10613) );
  XOR U10319 ( .A(n10612), .B(n10438), .Z(n10615) );
  XOR U10320 ( .A(n10616), .B(n10617), .Z(n10438) );
  AND U10321 ( .A(n431), .B(n10618), .Z(n10617) );
  XOR U10322 ( .A(n10619), .B(n10616), .Z(n10618) );
  XNOR U10323 ( .A(n10435), .B(n10612), .Z(n10614) );
  XOR U10324 ( .A(n10620), .B(n10621), .Z(n10435) );
  AND U10325 ( .A(n429), .B(n10622), .Z(n10621) );
  XOR U10326 ( .A(n10623), .B(n10620), .Z(n10622) );
  XOR U10327 ( .A(n10624), .B(n10625), .Z(n10612) );
  AND U10328 ( .A(n10626), .B(n10627), .Z(n10625) );
  XOR U10329 ( .A(n10624), .B(n10450), .Z(n10627) );
  XOR U10330 ( .A(n10628), .B(n10629), .Z(n10450) );
  AND U10331 ( .A(n431), .B(n10630), .Z(n10629) );
  XOR U10332 ( .A(n10631), .B(n10628), .Z(n10630) );
  XNOR U10333 ( .A(n10447), .B(n10624), .Z(n10626) );
  XOR U10334 ( .A(n10632), .B(n10633), .Z(n10447) );
  AND U10335 ( .A(n429), .B(n10634), .Z(n10633) );
  XOR U10336 ( .A(n10635), .B(n10632), .Z(n10634) );
  XOR U10337 ( .A(n10636), .B(n10637), .Z(n10624) );
  AND U10338 ( .A(n10638), .B(n10639), .Z(n10637) );
  XOR U10339 ( .A(n10636), .B(n10462), .Z(n10639) );
  XOR U10340 ( .A(n10640), .B(n10641), .Z(n10462) );
  AND U10341 ( .A(n431), .B(n10642), .Z(n10641) );
  XOR U10342 ( .A(n10643), .B(n10640), .Z(n10642) );
  XNOR U10343 ( .A(n10459), .B(n10636), .Z(n10638) );
  XOR U10344 ( .A(n10644), .B(n10645), .Z(n10459) );
  AND U10345 ( .A(n429), .B(n10646), .Z(n10645) );
  XOR U10346 ( .A(n10647), .B(n10644), .Z(n10646) );
  XOR U10347 ( .A(n10648), .B(n10649), .Z(n10636) );
  AND U10348 ( .A(n10650), .B(n10651), .Z(n10649) );
  XNOR U10349 ( .A(n10652), .B(n10475), .Z(n10651) );
  XOR U10350 ( .A(n10653), .B(n10654), .Z(n10475) );
  AND U10351 ( .A(n431), .B(n10655), .Z(n10654) );
  XOR U10352 ( .A(n10653), .B(n10656), .Z(n10655) );
  XNOR U10353 ( .A(n10472), .B(n10648), .Z(n10650) );
  XOR U10354 ( .A(n10657), .B(n10658), .Z(n10472) );
  AND U10355 ( .A(n429), .B(n10659), .Z(n10658) );
  XOR U10356 ( .A(n10657), .B(n10660), .Z(n10659) );
  IV U10357 ( .A(n10652), .Z(n10648) );
  AND U10358 ( .A(n10480), .B(n10483), .Z(n10652) );
  XNOR U10359 ( .A(n10661), .B(n10662), .Z(n10483) );
  AND U10360 ( .A(n431), .B(n10663), .Z(n10662) );
  XNOR U10361 ( .A(n10664), .B(n10661), .Z(n10663) );
  XOR U10362 ( .A(n10665), .B(n10666), .Z(n431) );
  AND U10363 ( .A(n10667), .B(n10668), .Z(n10666) );
  XNOR U10364 ( .A(n10488), .B(n10665), .Z(n10668) );
  AND U10365 ( .A(p_input[2815]), .B(p_input[2799]), .Z(n10488) );
  XOR U10366 ( .A(n10665), .B(n10489), .Z(n10667) );
  AND U10367 ( .A(p_input[2783]), .B(p_input[2767]), .Z(n10489) );
  XOR U10368 ( .A(n10669), .B(n10670), .Z(n10665) );
  AND U10369 ( .A(n10671), .B(n10672), .Z(n10670) );
  XOR U10370 ( .A(n10669), .B(n10499), .Z(n10672) );
  XNOR U10371 ( .A(p_input[2798]), .B(n10673), .Z(n10499) );
  AND U10372 ( .A(n259), .B(n10674), .Z(n10673) );
  XOR U10373 ( .A(p_input[2814]), .B(p_input[2798]), .Z(n10674) );
  XNOR U10374 ( .A(n10496), .B(n10669), .Z(n10671) );
  XOR U10375 ( .A(n10675), .B(n10676), .Z(n10496) );
  AND U10376 ( .A(n257), .B(n10677), .Z(n10676) );
  XOR U10377 ( .A(p_input[2782]), .B(p_input[2766]), .Z(n10677) );
  XOR U10378 ( .A(n10678), .B(n10679), .Z(n10669) );
  AND U10379 ( .A(n10680), .B(n10681), .Z(n10679) );
  XOR U10380 ( .A(n10678), .B(n10511), .Z(n10681) );
  XNOR U10381 ( .A(p_input[2797]), .B(n10682), .Z(n10511) );
  AND U10382 ( .A(n259), .B(n10683), .Z(n10682) );
  XOR U10383 ( .A(p_input[2813]), .B(p_input[2797]), .Z(n10683) );
  XNOR U10384 ( .A(n10508), .B(n10678), .Z(n10680) );
  XOR U10385 ( .A(n10684), .B(n10685), .Z(n10508) );
  AND U10386 ( .A(n257), .B(n10686), .Z(n10685) );
  XOR U10387 ( .A(p_input[2781]), .B(p_input[2765]), .Z(n10686) );
  XOR U10388 ( .A(n10687), .B(n10688), .Z(n10678) );
  AND U10389 ( .A(n10689), .B(n10690), .Z(n10688) );
  XOR U10390 ( .A(n10687), .B(n10523), .Z(n10690) );
  XNOR U10391 ( .A(p_input[2796]), .B(n10691), .Z(n10523) );
  AND U10392 ( .A(n259), .B(n10692), .Z(n10691) );
  XOR U10393 ( .A(p_input[2812]), .B(p_input[2796]), .Z(n10692) );
  XNOR U10394 ( .A(n10520), .B(n10687), .Z(n10689) );
  XOR U10395 ( .A(n10693), .B(n10694), .Z(n10520) );
  AND U10396 ( .A(n257), .B(n10695), .Z(n10694) );
  XOR U10397 ( .A(p_input[2780]), .B(p_input[2764]), .Z(n10695) );
  XOR U10398 ( .A(n10696), .B(n10697), .Z(n10687) );
  AND U10399 ( .A(n10698), .B(n10699), .Z(n10697) );
  XOR U10400 ( .A(n10696), .B(n10535), .Z(n10699) );
  XNOR U10401 ( .A(p_input[2795]), .B(n10700), .Z(n10535) );
  AND U10402 ( .A(n259), .B(n10701), .Z(n10700) );
  XOR U10403 ( .A(p_input[2811]), .B(p_input[2795]), .Z(n10701) );
  XNOR U10404 ( .A(n10532), .B(n10696), .Z(n10698) );
  XOR U10405 ( .A(n10702), .B(n10703), .Z(n10532) );
  AND U10406 ( .A(n257), .B(n10704), .Z(n10703) );
  XOR U10407 ( .A(p_input[2779]), .B(p_input[2763]), .Z(n10704) );
  XOR U10408 ( .A(n10705), .B(n10706), .Z(n10696) );
  AND U10409 ( .A(n10707), .B(n10708), .Z(n10706) );
  XOR U10410 ( .A(n10705), .B(n10547), .Z(n10708) );
  XNOR U10411 ( .A(p_input[2794]), .B(n10709), .Z(n10547) );
  AND U10412 ( .A(n259), .B(n10710), .Z(n10709) );
  XOR U10413 ( .A(p_input[2810]), .B(p_input[2794]), .Z(n10710) );
  XNOR U10414 ( .A(n10544), .B(n10705), .Z(n10707) );
  XOR U10415 ( .A(n10711), .B(n10712), .Z(n10544) );
  AND U10416 ( .A(n257), .B(n10713), .Z(n10712) );
  XOR U10417 ( .A(p_input[2778]), .B(p_input[2762]), .Z(n10713) );
  XOR U10418 ( .A(n10714), .B(n10715), .Z(n10705) );
  AND U10419 ( .A(n10716), .B(n10717), .Z(n10715) );
  XOR U10420 ( .A(n10714), .B(n10559), .Z(n10717) );
  XNOR U10421 ( .A(p_input[2793]), .B(n10718), .Z(n10559) );
  AND U10422 ( .A(n259), .B(n10719), .Z(n10718) );
  XOR U10423 ( .A(p_input[2809]), .B(p_input[2793]), .Z(n10719) );
  XNOR U10424 ( .A(n10556), .B(n10714), .Z(n10716) );
  XOR U10425 ( .A(n10720), .B(n10721), .Z(n10556) );
  AND U10426 ( .A(n257), .B(n10722), .Z(n10721) );
  XOR U10427 ( .A(p_input[2777]), .B(p_input[2761]), .Z(n10722) );
  XOR U10428 ( .A(n10723), .B(n10724), .Z(n10714) );
  AND U10429 ( .A(n10725), .B(n10726), .Z(n10724) );
  XOR U10430 ( .A(n10723), .B(n10571), .Z(n10726) );
  XNOR U10431 ( .A(p_input[2792]), .B(n10727), .Z(n10571) );
  AND U10432 ( .A(n259), .B(n10728), .Z(n10727) );
  XOR U10433 ( .A(p_input[2808]), .B(p_input[2792]), .Z(n10728) );
  XNOR U10434 ( .A(n10568), .B(n10723), .Z(n10725) );
  XOR U10435 ( .A(n10729), .B(n10730), .Z(n10568) );
  AND U10436 ( .A(n257), .B(n10731), .Z(n10730) );
  XOR U10437 ( .A(p_input[2776]), .B(p_input[2760]), .Z(n10731) );
  XOR U10438 ( .A(n10732), .B(n10733), .Z(n10723) );
  AND U10439 ( .A(n10734), .B(n10735), .Z(n10733) );
  XOR U10440 ( .A(n10732), .B(n10583), .Z(n10735) );
  XNOR U10441 ( .A(p_input[2791]), .B(n10736), .Z(n10583) );
  AND U10442 ( .A(n259), .B(n10737), .Z(n10736) );
  XOR U10443 ( .A(p_input[2807]), .B(p_input[2791]), .Z(n10737) );
  XNOR U10444 ( .A(n10580), .B(n10732), .Z(n10734) );
  XOR U10445 ( .A(n10738), .B(n10739), .Z(n10580) );
  AND U10446 ( .A(n257), .B(n10740), .Z(n10739) );
  XOR U10447 ( .A(p_input[2775]), .B(p_input[2759]), .Z(n10740) );
  XOR U10448 ( .A(n10741), .B(n10742), .Z(n10732) );
  AND U10449 ( .A(n10743), .B(n10744), .Z(n10742) );
  XOR U10450 ( .A(n10741), .B(n10595), .Z(n10744) );
  XNOR U10451 ( .A(p_input[2790]), .B(n10745), .Z(n10595) );
  AND U10452 ( .A(n259), .B(n10746), .Z(n10745) );
  XOR U10453 ( .A(p_input[2806]), .B(p_input[2790]), .Z(n10746) );
  XNOR U10454 ( .A(n10592), .B(n10741), .Z(n10743) );
  XOR U10455 ( .A(n10747), .B(n10748), .Z(n10592) );
  AND U10456 ( .A(n257), .B(n10749), .Z(n10748) );
  XOR U10457 ( .A(p_input[2774]), .B(p_input[2758]), .Z(n10749) );
  XOR U10458 ( .A(n10750), .B(n10751), .Z(n10741) );
  AND U10459 ( .A(n10752), .B(n10753), .Z(n10751) );
  XOR U10460 ( .A(n10750), .B(n10607), .Z(n10753) );
  XNOR U10461 ( .A(p_input[2789]), .B(n10754), .Z(n10607) );
  AND U10462 ( .A(n259), .B(n10755), .Z(n10754) );
  XOR U10463 ( .A(p_input[2805]), .B(p_input[2789]), .Z(n10755) );
  XNOR U10464 ( .A(n10604), .B(n10750), .Z(n10752) );
  XOR U10465 ( .A(n10756), .B(n10757), .Z(n10604) );
  AND U10466 ( .A(n257), .B(n10758), .Z(n10757) );
  XOR U10467 ( .A(p_input[2773]), .B(p_input[2757]), .Z(n10758) );
  XOR U10468 ( .A(n10759), .B(n10760), .Z(n10750) );
  AND U10469 ( .A(n10761), .B(n10762), .Z(n10760) );
  XOR U10470 ( .A(n10759), .B(n10619), .Z(n10762) );
  XNOR U10471 ( .A(p_input[2788]), .B(n10763), .Z(n10619) );
  AND U10472 ( .A(n259), .B(n10764), .Z(n10763) );
  XOR U10473 ( .A(p_input[2804]), .B(p_input[2788]), .Z(n10764) );
  XNOR U10474 ( .A(n10616), .B(n10759), .Z(n10761) );
  XOR U10475 ( .A(n10765), .B(n10766), .Z(n10616) );
  AND U10476 ( .A(n257), .B(n10767), .Z(n10766) );
  XOR U10477 ( .A(p_input[2772]), .B(p_input[2756]), .Z(n10767) );
  XOR U10478 ( .A(n10768), .B(n10769), .Z(n10759) );
  AND U10479 ( .A(n10770), .B(n10771), .Z(n10769) );
  XOR U10480 ( .A(n10768), .B(n10631), .Z(n10771) );
  XNOR U10481 ( .A(p_input[2787]), .B(n10772), .Z(n10631) );
  AND U10482 ( .A(n259), .B(n10773), .Z(n10772) );
  XOR U10483 ( .A(p_input[2803]), .B(p_input[2787]), .Z(n10773) );
  XNOR U10484 ( .A(n10628), .B(n10768), .Z(n10770) );
  XOR U10485 ( .A(n10774), .B(n10775), .Z(n10628) );
  AND U10486 ( .A(n257), .B(n10776), .Z(n10775) );
  XOR U10487 ( .A(p_input[2771]), .B(p_input[2755]), .Z(n10776) );
  XOR U10488 ( .A(n10777), .B(n10778), .Z(n10768) );
  AND U10489 ( .A(n10779), .B(n10780), .Z(n10778) );
  XOR U10490 ( .A(n10777), .B(n10643), .Z(n10780) );
  XNOR U10491 ( .A(p_input[2786]), .B(n10781), .Z(n10643) );
  AND U10492 ( .A(n259), .B(n10782), .Z(n10781) );
  XOR U10493 ( .A(p_input[2802]), .B(p_input[2786]), .Z(n10782) );
  XNOR U10494 ( .A(n10640), .B(n10777), .Z(n10779) );
  XOR U10495 ( .A(n10783), .B(n10784), .Z(n10640) );
  AND U10496 ( .A(n257), .B(n10785), .Z(n10784) );
  XOR U10497 ( .A(p_input[2770]), .B(p_input[2754]), .Z(n10785) );
  XOR U10498 ( .A(n10786), .B(n10787), .Z(n10777) );
  AND U10499 ( .A(n10788), .B(n10789), .Z(n10787) );
  XNOR U10500 ( .A(n10790), .B(n10656), .Z(n10789) );
  XNOR U10501 ( .A(p_input[2785]), .B(n10791), .Z(n10656) );
  AND U10502 ( .A(n259), .B(n10792), .Z(n10791) );
  XNOR U10503 ( .A(p_input[2801]), .B(n10793), .Z(n10792) );
  IV U10504 ( .A(p_input[2785]), .Z(n10793) );
  XNOR U10505 ( .A(n10653), .B(n10786), .Z(n10788) );
  XNOR U10506 ( .A(p_input[2753]), .B(n10794), .Z(n10653) );
  AND U10507 ( .A(n257), .B(n10795), .Z(n10794) );
  XOR U10508 ( .A(p_input[2769]), .B(p_input[2753]), .Z(n10795) );
  IV U10509 ( .A(n10790), .Z(n10786) );
  AND U10510 ( .A(n10661), .B(n10664), .Z(n10790) );
  XOR U10511 ( .A(p_input[2784]), .B(n10796), .Z(n10664) );
  AND U10512 ( .A(n259), .B(n10797), .Z(n10796) );
  XOR U10513 ( .A(p_input[2800]), .B(p_input[2784]), .Z(n10797) );
  XOR U10514 ( .A(n10798), .B(n10799), .Z(n259) );
  AND U10515 ( .A(n10800), .B(n10801), .Z(n10799) );
  XNOR U10516 ( .A(p_input[2815]), .B(n10798), .Z(n10801) );
  XOR U10517 ( .A(n10798), .B(p_input[2799]), .Z(n10800) );
  XOR U10518 ( .A(n10802), .B(n10803), .Z(n10798) );
  AND U10519 ( .A(n10804), .B(n10805), .Z(n10803) );
  XNOR U10520 ( .A(p_input[2814]), .B(n10802), .Z(n10805) );
  XOR U10521 ( .A(n10802), .B(p_input[2798]), .Z(n10804) );
  XOR U10522 ( .A(n10806), .B(n10807), .Z(n10802) );
  AND U10523 ( .A(n10808), .B(n10809), .Z(n10807) );
  XNOR U10524 ( .A(p_input[2813]), .B(n10806), .Z(n10809) );
  XOR U10525 ( .A(n10806), .B(p_input[2797]), .Z(n10808) );
  XOR U10526 ( .A(n10810), .B(n10811), .Z(n10806) );
  AND U10527 ( .A(n10812), .B(n10813), .Z(n10811) );
  XNOR U10528 ( .A(p_input[2812]), .B(n10810), .Z(n10813) );
  XOR U10529 ( .A(n10810), .B(p_input[2796]), .Z(n10812) );
  XOR U10530 ( .A(n10814), .B(n10815), .Z(n10810) );
  AND U10531 ( .A(n10816), .B(n10817), .Z(n10815) );
  XNOR U10532 ( .A(p_input[2811]), .B(n10814), .Z(n10817) );
  XOR U10533 ( .A(n10814), .B(p_input[2795]), .Z(n10816) );
  XOR U10534 ( .A(n10818), .B(n10819), .Z(n10814) );
  AND U10535 ( .A(n10820), .B(n10821), .Z(n10819) );
  XNOR U10536 ( .A(p_input[2810]), .B(n10818), .Z(n10821) );
  XOR U10537 ( .A(n10818), .B(p_input[2794]), .Z(n10820) );
  XOR U10538 ( .A(n10822), .B(n10823), .Z(n10818) );
  AND U10539 ( .A(n10824), .B(n10825), .Z(n10823) );
  XNOR U10540 ( .A(p_input[2809]), .B(n10822), .Z(n10825) );
  XOR U10541 ( .A(n10822), .B(p_input[2793]), .Z(n10824) );
  XOR U10542 ( .A(n10826), .B(n10827), .Z(n10822) );
  AND U10543 ( .A(n10828), .B(n10829), .Z(n10827) );
  XNOR U10544 ( .A(p_input[2808]), .B(n10826), .Z(n10829) );
  XOR U10545 ( .A(n10826), .B(p_input[2792]), .Z(n10828) );
  XOR U10546 ( .A(n10830), .B(n10831), .Z(n10826) );
  AND U10547 ( .A(n10832), .B(n10833), .Z(n10831) );
  XNOR U10548 ( .A(p_input[2807]), .B(n10830), .Z(n10833) );
  XOR U10549 ( .A(n10830), .B(p_input[2791]), .Z(n10832) );
  XOR U10550 ( .A(n10834), .B(n10835), .Z(n10830) );
  AND U10551 ( .A(n10836), .B(n10837), .Z(n10835) );
  XNOR U10552 ( .A(p_input[2806]), .B(n10834), .Z(n10837) );
  XOR U10553 ( .A(n10834), .B(p_input[2790]), .Z(n10836) );
  XOR U10554 ( .A(n10838), .B(n10839), .Z(n10834) );
  AND U10555 ( .A(n10840), .B(n10841), .Z(n10839) );
  XNOR U10556 ( .A(p_input[2805]), .B(n10838), .Z(n10841) );
  XOR U10557 ( .A(n10838), .B(p_input[2789]), .Z(n10840) );
  XOR U10558 ( .A(n10842), .B(n10843), .Z(n10838) );
  AND U10559 ( .A(n10844), .B(n10845), .Z(n10843) );
  XNOR U10560 ( .A(p_input[2804]), .B(n10842), .Z(n10845) );
  XOR U10561 ( .A(n10842), .B(p_input[2788]), .Z(n10844) );
  XOR U10562 ( .A(n10846), .B(n10847), .Z(n10842) );
  AND U10563 ( .A(n10848), .B(n10849), .Z(n10847) );
  XNOR U10564 ( .A(p_input[2803]), .B(n10846), .Z(n10849) );
  XOR U10565 ( .A(n10846), .B(p_input[2787]), .Z(n10848) );
  XOR U10566 ( .A(n10850), .B(n10851), .Z(n10846) );
  AND U10567 ( .A(n10852), .B(n10853), .Z(n10851) );
  XNOR U10568 ( .A(p_input[2802]), .B(n10850), .Z(n10853) );
  XOR U10569 ( .A(n10850), .B(p_input[2786]), .Z(n10852) );
  XNOR U10570 ( .A(n10854), .B(n10855), .Z(n10850) );
  AND U10571 ( .A(n10856), .B(n10857), .Z(n10855) );
  XOR U10572 ( .A(p_input[2801]), .B(n10854), .Z(n10857) );
  XNOR U10573 ( .A(p_input[2785]), .B(n10854), .Z(n10856) );
  AND U10574 ( .A(p_input[2800]), .B(n10858), .Z(n10854) );
  IV U10575 ( .A(p_input[2784]), .Z(n10858) );
  XNOR U10576 ( .A(p_input[2752]), .B(n10859), .Z(n10661) );
  AND U10577 ( .A(n257), .B(n10860), .Z(n10859) );
  XOR U10578 ( .A(p_input[2768]), .B(p_input[2752]), .Z(n10860) );
  XOR U10579 ( .A(n10861), .B(n10862), .Z(n257) );
  AND U10580 ( .A(n10863), .B(n10864), .Z(n10862) );
  XNOR U10581 ( .A(p_input[2783]), .B(n10861), .Z(n10864) );
  XOR U10582 ( .A(n10861), .B(p_input[2767]), .Z(n10863) );
  XOR U10583 ( .A(n10865), .B(n10866), .Z(n10861) );
  AND U10584 ( .A(n10867), .B(n10868), .Z(n10866) );
  XNOR U10585 ( .A(p_input[2782]), .B(n10865), .Z(n10868) );
  XNOR U10586 ( .A(n10865), .B(n10675), .Z(n10867) );
  IV U10587 ( .A(p_input[2766]), .Z(n10675) );
  XOR U10588 ( .A(n10869), .B(n10870), .Z(n10865) );
  AND U10589 ( .A(n10871), .B(n10872), .Z(n10870) );
  XNOR U10590 ( .A(p_input[2781]), .B(n10869), .Z(n10872) );
  XNOR U10591 ( .A(n10869), .B(n10684), .Z(n10871) );
  IV U10592 ( .A(p_input[2765]), .Z(n10684) );
  XOR U10593 ( .A(n10873), .B(n10874), .Z(n10869) );
  AND U10594 ( .A(n10875), .B(n10876), .Z(n10874) );
  XNOR U10595 ( .A(p_input[2780]), .B(n10873), .Z(n10876) );
  XNOR U10596 ( .A(n10873), .B(n10693), .Z(n10875) );
  IV U10597 ( .A(p_input[2764]), .Z(n10693) );
  XOR U10598 ( .A(n10877), .B(n10878), .Z(n10873) );
  AND U10599 ( .A(n10879), .B(n10880), .Z(n10878) );
  XNOR U10600 ( .A(p_input[2779]), .B(n10877), .Z(n10880) );
  XNOR U10601 ( .A(n10877), .B(n10702), .Z(n10879) );
  IV U10602 ( .A(p_input[2763]), .Z(n10702) );
  XOR U10603 ( .A(n10881), .B(n10882), .Z(n10877) );
  AND U10604 ( .A(n10883), .B(n10884), .Z(n10882) );
  XNOR U10605 ( .A(p_input[2778]), .B(n10881), .Z(n10884) );
  XNOR U10606 ( .A(n10881), .B(n10711), .Z(n10883) );
  IV U10607 ( .A(p_input[2762]), .Z(n10711) );
  XOR U10608 ( .A(n10885), .B(n10886), .Z(n10881) );
  AND U10609 ( .A(n10887), .B(n10888), .Z(n10886) );
  XNOR U10610 ( .A(p_input[2777]), .B(n10885), .Z(n10888) );
  XNOR U10611 ( .A(n10885), .B(n10720), .Z(n10887) );
  IV U10612 ( .A(p_input[2761]), .Z(n10720) );
  XOR U10613 ( .A(n10889), .B(n10890), .Z(n10885) );
  AND U10614 ( .A(n10891), .B(n10892), .Z(n10890) );
  XNOR U10615 ( .A(p_input[2776]), .B(n10889), .Z(n10892) );
  XNOR U10616 ( .A(n10889), .B(n10729), .Z(n10891) );
  IV U10617 ( .A(p_input[2760]), .Z(n10729) );
  XOR U10618 ( .A(n10893), .B(n10894), .Z(n10889) );
  AND U10619 ( .A(n10895), .B(n10896), .Z(n10894) );
  XNOR U10620 ( .A(p_input[2775]), .B(n10893), .Z(n10896) );
  XNOR U10621 ( .A(n10893), .B(n10738), .Z(n10895) );
  IV U10622 ( .A(p_input[2759]), .Z(n10738) );
  XOR U10623 ( .A(n10897), .B(n10898), .Z(n10893) );
  AND U10624 ( .A(n10899), .B(n10900), .Z(n10898) );
  XNOR U10625 ( .A(p_input[2774]), .B(n10897), .Z(n10900) );
  XNOR U10626 ( .A(n10897), .B(n10747), .Z(n10899) );
  IV U10627 ( .A(p_input[2758]), .Z(n10747) );
  XOR U10628 ( .A(n10901), .B(n10902), .Z(n10897) );
  AND U10629 ( .A(n10903), .B(n10904), .Z(n10902) );
  XNOR U10630 ( .A(p_input[2773]), .B(n10901), .Z(n10904) );
  XNOR U10631 ( .A(n10901), .B(n10756), .Z(n10903) );
  IV U10632 ( .A(p_input[2757]), .Z(n10756) );
  XOR U10633 ( .A(n10905), .B(n10906), .Z(n10901) );
  AND U10634 ( .A(n10907), .B(n10908), .Z(n10906) );
  XNOR U10635 ( .A(p_input[2772]), .B(n10905), .Z(n10908) );
  XNOR U10636 ( .A(n10905), .B(n10765), .Z(n10907) );
  IV U10637 ( .A(p_input[2756]), .Z(n10765) );
  XOR U10638 ( .A(n10909), .B(n10910), .Z(n10905) );
  AND U10639 ( .A(n10911), .B(n10912), .Z(n10910) );
  XNOR U10640 ( .A(p_input[2771]), .B(n10909), .Z(n10912) );
  XNOR U10641 ( .A(n10909), .B(n10774), .Z(n10911) );
  IV U10642 ( .A(p_input[2755]), .Z(n10774) );
  XOR U10643 ( .A(n10913), .B(n10914), .Z(n10909) );
  AND U10644 ( .A(n10915), .B(n10916), .Z(n10914) );
  XNOR U10645 ( .A(p_input[2770]), .B(n10913), .Z(n10916) );
  XNOR U10646 ( .A(n10913), .B(n10783), .Z(n10915) );
  IV U10647 ( .A(p_input[2754]), .Z(n10783) );
  XNOR U10648 ( .A(n10917), .B(n10918), .Z(n10913) );
  AND U10649 ( .A(n10919), .B(n10920), .Z(n10918) );
  XOR U10650 ( .A(p_input[2769]), .B(n10917), .Z(n10920) );
  XNOR U10651 ( .A(p_input[2753]), .B(n10917), .Z(n10919) );
  AND U10652 ( .A(p_input[2768]), .B(n10921), .Z(n10917) );
  IV U10653 ( .A(p_input[2752]), .Z(n10921) );
  XOR U10654 ( .A(n10922), .B(n10923), .Z(n10480) );
  AND U10655 ( .A(n429), .B(n10924), .Z(n10923) );
  XNOR U10656 ( .A(n10925), .B(n10922), .Z(n10924) );
  XOR U10657 ( .A(n10926), .B(n10927), .Z(n429) );
  AND U10658 ( .A(n10928), .B(n10929), .Z(n10927) );
  XNOR U10659 ( .A(n10490), .B(n10926), .Z(n10929) );
  AND U10660 ( .A(p_input[2751]), .B(p_input[2735]), .Z(n10490) );
  XOR U10661 ( .A(n10926), .B(n10491), .Z(n10928) );
  AND U10662 ( .A(p_input[2719]), .B(p_input[2703]), .Z(n10491) );
  XOR U10663 ( .A(n10930), .B(n10931), .Z(n10926) );
  AND U10664 ( .A(n10932), .B(n10933), .Z(n10931) );
  XOR U10665 ( .A(n10930), .B(n10503), .Z(n10933) );
  XNOR U10666 ( .A(p_input[2734]), .B(n10934), .Z(n10503) );
  AND U10667 ( .A(n263), .B(n10935), .Z(n10934) );
  XOR U10668 ( .A(p_input[2750]), .B(p_input[2734]), .Z(n10935) );
  XNOR U10669 ( .A(n10500), .B(n10930), .Z(n10932) );
  XOR U10670 ( .A(n10936), .B(n10937), .Z(n10500) );
  AND U10671 ( .A(n260), .B(n10938), .Z(n10937) );
  XOR U10672 ( .A(p_input[2718]), .B(p_input[2702]), .Z(n10938) );
  XOR U10673 ( .A(n10939), .B(n10940), .Z(n10930) );
  AND U10674 ( .A(n10941), .B(n10942), .Z(n10940) );
  XOR U10675 ( .A(n10939), .B(n10515), .Z(n10942) );
  XNOR U10676 ( .A(p_input[2733]), .B(n10943), .Z(n10515) );
  AND U10677 ( .A(n263), .B(n10944), .Z(n10943) );
  XOR U10678 ( .A(p_input[2749]), .B(p_input[2733]), .Z(n10944) );
  XNOR U10679 ( .A(n10512), .B(n10939), .Z(n10941) );
  XOR U10680 ( .A(n10945), .B(n10946), .Z(n10512) );
  AND U10681 ( .A(n260), .B(n10947), .Z(n10946) );
  XOR U10682 ( .A(p_input[2717]), .B(p_input[2701]), .Z(n10947) );
  XOR U10683 ( .A(n10948), .B(n10949), .Z(n10939) );
  AND U10684 ( .A(n10950), .B(n10951), .Z(n10949) );
  XOR U10685 ( .A(n10948), .B(n10527), .Z(n10951) );
  XNOR U10686 ( .A(p_input[2732]), .B(n10952), .Z(n10527) );
  AND U10687 ( .A(n263), .B(n10953), .Z(n10952) );
  XOR U10688 ( .A(p_input[2748]), .B(p_input[2732]), .Z(n10953) );
  XNOR U10689 ( .A(n10524), .B(n10948), .Z(n10950) );
  XOR U10690 ( .A(n10954), .B(n10955), .Z(n10524) );
  AND U10691 ( .A(n260), .B(n10956), .Z(n10955) );
  XOR U10692 ( .A(p_input[2716]), .B(p_input[2700]), .Z(n10956) );
  XOR U10693 ( .A(n10957), .B(n10958), .Z(n10948) );
  AND U10694 ( .A(n10959), .B(n10960), .Z(n10958) );
  XOR U10695 ( .A(n10957), .B(n10539), .Z(n10960) );
  XNOR U10696 ( .A(p_input[2731]), .B(n10961), .Z(n10539) );
  AND U10697 ( .A(n263), .B(n10962), .Z(n10961) );
  XOR U10698 ( .A(p_input[2747]), .B(p_input[2731]), .Z(n10962) );
  XNOR U10699 ( .A(n10536), .B(n10957), .Z(n10959) );
  XOR U10700 ( .A(n10963), .B(n10964), .Z(n10536) );
  AND U10701 ( .A(n260), .B(n10965), .Z(n10964) );
  XOR U10702 ( .A(p_input[2715]), .B(p_input[2699]), .Z(n10965) );
  XOR U10703 ( .A(n10966), .B(n10967), .Z(n10957) );
  AND U10704 ( .A(n10968), .B(n10969), .Z(n10967) );
  XOR U10705 ( .A(n10966), .B(n10551), .Z(n10969) );
  XNOR U10706 ( .A(p_input[2730]), .B(n10970), .Z(n10551) );
  AND U10707 ( .A(n263), .B(n10971), .Z(n10970) );
  XOR U10708 ( .A(p_input[2746]), .B(p_input[2730]), .Z(n10971) );
  XNOR U10709 ( .A(n10548), .B(n10966), .Z(n10968) );
  XOR U10710 ( .A(n10972), .B(n10973), .Z(n10548) );
  AND U10711 ( .A(n260), .B(n10974), .Z(n10973) );
  XOR U10712 ( .A(p_input[2714]), .B(p_input[2698]), .Z(n10974) );
  XOR U10713 ( .A(n10975), .B(n10976), .Z(n10966) );
  AND U10714 ( .A(n10977), .B(n10978), .Z(n10976) );
  XOR U10715 ( .A(n10975), .B(n10563), .Z(n10978) );
  XNOR U10716 ( .A(p_input[2729]), .B(n10979), .Z(n10563) );
  AND U10717 ( .A(n263), .B(n10980), .Z(n10979) );
  XOR U10718 ( .A(p_input[2745]), .B(p_input[2729]), .Z(n10980) );
  XNOR U10719 ( .A(n10560), .B(n10975), .Z(n10977) );
  XOR U10720 ( .A(n10981), .B(n10982), .Z(n10560) );
  AND U10721 ( .A(n260), .B(n10983), .Z(n10982) );
  XOR U10722 ( .A(p_input[2713]), .B(p_input[2697]), .Z(n10983) );
  XOR U10723 ( .A(n10984), .B(n10985), .Z(n10975) );
  AND U10724 ( .A(n10986), .B(n10987), .Z(n10985) );
  XOR U10725 ( .A(n10984), .B(n10575), .Z(n10987) );
  XNOR U10726 ( .A(p_input[2728]), .B(n10988), .Z(n10575) );
  AND U10727 ( .A(n263), .B(n10989), .Z(n10988) );
  XOR U10728 ( .A(p_input[2744]), .B(p_input[2728]), .Z(n10989) );
  XNOR U10729 ( .A(n10572), .B(n10984), .Z(n10986) );
  XOR U10730 ( .A(n10990), .B(n10991), .Z(n10572) );
  AND U10731 ( .A(n260), .B(n10992), .Z(n10991) );
  XOR U10732 ( .A(p_input[2712]), .B(p_input[2696]), .Z(n10992) );
  XOR U10733 ( .A(n10993), .B(n10994), .Z(n10984) );
  AND U10734 ( .A(n10995), .B(n10996), .Z(n10994) );
  XOR U10735 ( .A(n10993), .B(n10587), .Z(n10996) );
  XNOR U10736 ( .A(p_input[2727]), .B(n10997), .Z(n10587) );
  AND U10737 ( .A(n263), .B(n10998), .Z(n10997) );
  XOR U10738 ( .A(p_input[2743]), .B(p_input[2727]), .Z(n10998) );
  XNOR U10739 ( .A(n10584), .B(n10993), .Z(n10995) );
  XOR U10740 ( .A(n10999), .B(n11000), .Z(n10584) );
  AND U10741 ( .A(n260), .B(n11001), .Z(n11000) );
  XOR U10742 ( .A(p_input[2711]), .B(p_input[2695]), .Z(n11001) );
  XOR U10743 ( .A(n11002), .B(n11003), .Z(n10993) );
  AND U10744 ( .A(n11004), .B(n11005), .Z(n11003) );
  XOR U10745 ( .A(n11002), .B(n10599), .Z(n11005) );
  XNOR U10746 ( .A(p_input[2726]), .B(n11006), .Z(n10599) );
  AND U10747 ( .A(n263), .B(n11007), .Z(n11006) );
  XOR U10748 ( .A(p_input[2742]), .B(p_input[2726]), .Z(n11007) );
  XNOR U10749 ( .A(n10596), .B(n11002), .Z(n11004) );
  XOR U10750 ( .A(n11008), .B(n11009), .Z(n10596) );
  AND U10751 ( .A(n260), .B(n11010), .Z(n11009) );
  XOR U10752 ( .A(p_input[2710]), .B(p_input[2694]), .Z(n11010) );
  XOR U10753 ( .A(n11011), .B(n11012), .Z(n11002) );
  AND U10754 ( .A(n11013), .B(n11014), .Z(n11012) );
  XOR U10755 ( .A(n11011), .B(n10611), .Z(n11014) );
  XNOR U10756 ( .A(p_input[2725]), .B(n11015), .Z(n10611) );
  AND U10757 ( .A(n263), .B(n11016), .Z(n11015) );
  XOR U10758 ( .A(p_input[2741]), .B(p_input[2725]), .Z(n11016) );
  XNOR U10759 ( .A(n10608), .B(n11011), .Z(n11013) );
  XOR U10760 ( .A(n11017), .B(n11018), .Z(n10608) );
  AND U10761 ( .A(n260), .B(n11019), .Z(n11018) );
  XOR U10762 ( .A(p_input[2709]), .B(p_input[2693]), .Z(n11019) );
  XOR U10763 ( .A(n11020), .B(n11021), .Z(n11011) );
  AND U10764 ( .A(n11022), .B(n11023), .Z(n11021) );
  XOR U10765 ( .A(n11020), .B(n10623), .Z(n11023) );
  XNOR U10766 ( .A(p_input[2724]), .B(n11024), .Z(n10623) );
  AND U10767 ( .A(n263), .B(n11025), .Z(n11024) );
  XOR U10768 ( .A(p_input[2740]), .B(p_input[2724]), .Z(n11025) );
  XNOR U10769 ( .A(n10620), .B(n11020), .Z(n11022) );
  XOR U10770 ( .A(n11026), .B(n11027), .Z(n10620) );
  AND U10771 ( .A(n260), .B(n11028), .Z(n11027) );
  XOR U10772 ( .A(p_input[2708]), .B(p_input[2692]), .Z(n11028) );
  XOR U10773 ( .A(n11029), .B(n11030), .Z(n11020) );
  AND U10774 ( .A(n11031), .B(n11032), .Z(n11030) );
  XOR U10775 ( .A(n11029), .B(n10635), .Z(n11032) );
  XNOR U10776 ( .A(p_input[2723]), .B(n11033), .Z(n10635) );
  AND U10777 ( .A(n263), .B(n11034), .Z(n11033) );
  XOR U10778 ( .A(p_input[2739]), .B(p_input[2723]), .Z(n11034) );
  XNOR U10779 ( .A(n10632), .B(n11029), .Z(n11031) );
  XOR U10780 ( .A(n11035), .B(n11036), .Z(n10632) );
  AND U10781 ( .A(n260), .B(n11037), .Z(n11036) );
  XOR U10782 ( .A(p_input[2707]), .B(p_input[2691]), .Z(n11037) );
  XOR U10783 ( .A(n11038), .B(n11039), .Z(n11029) );
  AND U10784 ( .A(n11040), .B(n11041), .Z(n11039) );
  XOR U10785 ( .A(n11038), .B(n10647), .Z(n11041) );
  XNOR U10786 ( .A(p_input[2722]), .B(n11042), .Z(n10647) );
  AND U10787 ( .A(n263), .B(n11043), .Z(n11042) );
  XOR U10788 ( .A(p_input[2738]), .B(p_input[2722]), .Z(n11043) );
  XNOR U10789 ( .A(n10644), .B(n11038), .Z(n11040) );
  XOR U10790 ( .A(n11044), .B(n11045), .Z(n10644) );
  AND U10791 ( .A(n260), .B(n11046), .Z(n11045) );
  XOR U10792 ( .A(p_input[2706]), .B(p_input[2690]), .Z(n11046) );
  XOR U10793 ( .A(n11047), .B(n11048), .Z(n11038) );
  AND U10794 ( .A(n11049), .B(n11050), .Z(n11048) );
  XNOR U10795 ( .A(n11051), .B(n10660), .Z(n11050) );
  XNOR U10796 ( .A(p_input[2721]), .B(n11052), .Z(n10660) );
  AND U10797 ( .A(n263), .B(n11053), .Z(n11052) );
  XNOR U10798 ( .A(p_input[2737]), .B(n11054), .Z(n11053) );
  IV U10799 ( .A(p_input[2721]), .Z(n11054) );
  XNOR U10800 ( .A(n10657), .B(n11047), .Z(n11049) );
  XNOR U10801 ( .A(p_input[2689]), .B(n11055), .Z(n10657) );
  AND U10802 ( .A(n260), .B(n11056), .Z(n11055) );
  XOR U10803 ( .A(p_input[2705]), .B(p_input[2689]), .Z(n11056) );
  IV U10804 ( .A(n11051), .Z(n11047) );
  AND U10805 ( .A(n10922), .B(n10925), .Z(n11051) );
  XOR U10806 ( .A(p_input[2720]), .B(n11057), .Z(n10925) );
  AND U10807 ( .A(n263), .B(n11058), .Z(n11057) );
  XOR U10808 ( .A(p_input[2736]), .B(p_input[2720]), .Z(n11058) );
  XOR U10809 ( .A(n11059), .B(n11060), .Z(n263) );
  AND U10810 ( .A(n11061), .B(n11062), .Z(n11060) );
  XNOR U10811 ( .A(p_input[2751]), .B(n11059), .Z(n11062) );
  XOR U10812 ( .A(n11059), .B(p_input[2735]), .Z(n11061) );
  XOR U10813 ( .A(n11063), .B(n11064), .Z(n11059) );
  AND U10814 ( .A(n11065), .B(n11066), .Z(n11064) );
  XNOR U10815 ( .A(p_input[2750]), .B(n11063), .Z(n11066) );
  XOR U10816 ( .A(n11063), .B(p_input[2734]), .Z(n11065) );
  XOR U10817 ( .A(n11067), .B(n11068), .Z(n11063) );
  AND U10818 ( .A(n11069), .B(n11070), .Z(n11068) );
  XNOR U10819 ( .A(p_input[2749]), .B(n11067), .Z(n11070) );
  XOR U10820 ( .A(n11067), .B(p_input[2733]), .Z(n11069) );
  XOR U10821 ( .A(n11071), .B(n11072), .Z(n11067) );
  AND U10822 ( .A(n11073), .B(n11074), .Z(n11072) );
  XNOR U10823 ( .A(p_input[2748]), .B(n11071), .Z(n11074) );
  XOR U10824 ( .A(n11071), .B(p_input[2732]), .Z(n11073) );
  XOR U10825 ( .A(n11075), .B(n11076), .Z(n11071) );
  AND U10826 ( .A(n11077), .B(n11078), .Z(n11076) );
  XNOR U10827 ( .A(p_input[2747]), .B(n11075), .Z(n11078) );
  XOR U10828 ( .A(n11075), .B(p_input[2731]), .Z(n11077) );
  XOR U10829 ( .A(n11079), .B(n11080), .Z(n11075) );
  AND U10830 ( .A(n11081), .B(n11082), .Z(n11080) );
  XNOR U10831 ( .A(p_input[2746]), .B(n11079), .Z(n11082) );
  XOR U10832 ( .A(n11079), .B(p_input[2730]), .Z(n11081) );
  XOR U10833 ( .A(n11083), .B(n11084), .Z(n11079) );
  AND U10834 ( .A(n11085), .B(n11086), .Z(n11084) );
  XNOR U10835 ( .A(p_input[2745]), .B(n11083), .Z(n11086) );
  XOR U10836 ( .A(n11083), .B(p_input[2729]), .Z(n11085) );
  XOR U10837 ( .A(n11087), .B(n11088), .Z(n11083) );
  AND U10838 ( .A(n11089), .B(n11090), .Z(n11088) );
  XNOR U10839 ( .A(p_input[2744]), .B(n11087), .Z(n11090) );
  XOR U10840 ( .A(n11087), .B(p_input[2728]), .Z(n11089) );
  XOR U10841 ( .A(n11091), .B(n11092), .Z(n11087) );
  AND U10842 ( .A(n11093), .B(n11094), .Z(n11092) );
  XNOR U10843 ( .A(p_input[2743]), .B(n11091), .Z(n11094) );
  XOR U10844 ( .A(n11091), .B(p_input[2727]), .Z(n11093) );
  XOR U10845 ( .A(n11095), .B(n11096), .Z(n11091) );
  AND U10846 ( .A(n11097), .B(n11098), .Z(n11096) );
  XNOR U10847 ( .A(p_input[2742]), .B(n11095), .Z(n11098) );
  XOR U10848 ( .A(n11095), .B(p_input[2726]), .Z(n11097) );
  XOR U10849 ( .A(n11099), .B(n11100), .Z(n11095) );
  AND U10850 ( .A(n11101), .B(n11102), .Z(n11100) );
  XNOR U10851 ( .A(p_input[2741]), .B(n11099), .Z(n11102) );
  XOR U10852 ( .A(n11099), .B(p_input[2725]), .Z(n11101) );
  XOR U10853 ( .A(n11103), .B(n11104), .Z(n11099) );
  AND U10854 ( .A(n11105), .B(n11106), .Z(n11104) );
  XNOR U10855 ( .A(p_input[2740]), .B(n11103), .Z(n11106) );
  XOR U10856 ( .A(n11103), .B(p_input[2724]), .Z(n11105) );
  XOR U10857 ( .A(n11107), .B(n11108), .Z(n11103) );
  AND U10858 ( .A(n11109), .B(n11110), .Z(n11108) );
  XNOR U10859 ( .A(p_input[2739]), .B(n11107), .Z(n11110) );
  XOR U10860 ( .A(n11107), .B(p_input[2723]), .Z(n11109) );
  XOR U10861 ( .A(n11111), .B(n11112), .Z(n11107) );
  AND U10862 ( .A(n11113), .B(n11114), .Z(n11112) );
  XNOR U10863 ( .A(p_input[2738]), .B(n11111), .Z(n11114) );
  XOR U10864 ( .A(n11111), .B(p_input[2722]), .Z(n11113) );
  XNOR U10865 ( .A(n11115), .B(n11116), .Z(n11111) );
  AND U10866 ( .A(n11117), .B(n11118), .Z(n11116) );
  XOR U10867 ( .A(p_input[2737]), .B(n11115), .Z(n11118) );
  XNOR U10868 ( .A(p_input[2721]), .B(n11115), .Z(n11117) );
  AND U10869 ( .A(p_input[2736]), .B(n11119), .Z(n11115) );
  IV U10870 ( .A(p_input[2720]), .Z(n11119) );
  XNOR U10871 ( .A(p_input[2688]), .B(n11120), .Z(n10922) );
  AND U10872 ( .A(n260), .B(n11121), .Z(n11120) );
  XOR U10873 ( .A(p_input[2704]), .B(p_input[2688]), .Z(n11121) );
  XOR U10874 ( .A(n11122), .B(n11123), .Z(n260) );
  AND U10875 ( .A(n11124), .B(n11125), .Z(n11123) );
  XNOR U10876 ( .A(p_input[2719]), .B(n11122), .Z(n11125) );
  XOR U10877 ( .A(n11122), .B(p_input[2703]), .Z(n11124) );
  XOR U10878 ( .A(n11126), .B(n11127), .Z(n11122) );
  AND U10879 ( .A(n11128), .B(n11129), .Z(n11127) );
  XNOR U10880 ( .A(p_input[2718]), .B(n11126), .Z(n11129) );
  XNOR U10881 ( .A(n11126), .B(n10936), .Z(n11128) );
  IV U10882 ( .A(p_input[2702]), .Z(n10936) );
  XOR U10883 ( .A(n11130), .B(n11131), .Z(n11126) );
  AND U10884 ( .A(n11132), .B(n11133), .Z(n11131) );
  XNOR U10885 ( .A(p_input[2717]), .B(n11130), .Z(n11133) );
  XNOR U10886 ( .A(n11130), .B(n10945), .Z(n11132) );
  IV U10887 ( .A(p_input[2701]), .Z(n10945) );
  XOR U10888 ( .A(n11134), .B(n11135), .Z(n11130) );
  AND U10889 ( .A(n11136), .B(n11137), .Z(n11135) );
  XNOR U10890 ( .A(p_input[2716]), .B(n11134), .Z(n11137) );
  XNOR U10891 ( .A(n11134), .B(n10954), .Z(n11136) );
  IV U10892 ( .A(p_input[2700]), .Z(n10954) );
  XOR U10893 ( .A(n11138), .B(n11139), .Z(n11134) );
  AND U10894 ( .A(n11140), .B(n11141), .Z(n11139) );
  XNOR U10895 ( .A(p_input[2715]), .B(n11138), .Z(n11141) );
  XNOR U10896 ( .A(n11138), .B(n10963), .Z(n11140) );
  IV U10897 ( .A(p_input[2699]), .Z(n10963) );
  XOR U10898 ( .A(n11142), .B(n11143), .Z(n11138) );
  AND U10899 ( .A(n11144), .B(n11145), .Z(n11143) );
  XNOR U10900 ( .A(p_input[2714]), .B(n11142), .Z(n11145) );
  XNOR U10901 ( .A(n11142), .B(n10972), .Z(n11144) );
  IV U10902 ( .A(p_input[2698]), .Z(n10972) );
  XOR U10903 ( .A(n11146), .B(n11147), .Z(n11142) );
  AND U10904 ( .A(n11148), .B(n11149), .Z(n11147) );
  XNOR U10905 ( .A(p_input[2713]), .B(n11146), .Z(n11149) );
  XNOR U10906 ( .A(n11146), .B(n10981), .Z(n11148) );
  IV U10907 ( .A(p_input[2697]), .Z(n10981) );
  XOR U10908 ( .A(n11150), .B(n11151), .Z(n11146) );
  AND U10909 ( .A(n11152), .B(n11153), .Z(n11151) );
  XNOR U10910 ( .A(p_input[2712]), .B(n11150), .Z(n11153) );
  XNOR U10911 ( .A(n11150), .B(n10990), .Z(n11152) );
  IV U10912 ( .A(p_input[2696]), .Z(n10990) );
  XOR U10913 ( .A(n11154), .B(n11155), .Z(n11150) );
  AND U10914 ( .A(n11156), .B(n11157), .Z(n11155) );
  XNOR U10915 ( .A(p_input[2711]), .B(n11154), .Z(n11157) );
  XNOR U10916 ( .A(n11154), .B(n10999), .Z(n11156) );
  IV U10917 ( .A(p_input[2695]), .Z(n10999) );
  XOR U10918 ( .A(n11158), .B(n11159), .Z(n11154) );
  AND U10919 ( .A(n11160), .B(n11161), .Z(n11159) );
  XNOR U10920 ( .A(p_input[2710]), .B(n11158), .Z(n11161) );
  XNOR U10921 ( .A(n11158), .B(n11008), .Z(n11160) );
  IV U10922 ( .A(p_input[2694]), .Z(n11008) );
  XOR U10923 ( .A(n11162), .B(n11163), .Z(n11158) );
  AND U10924 ( .A(n11164), .B(n11165), .Z(n11163) );
  XNOR U10925 ( .A(p_input[2709]), .B(n11162), .Z(n11165) );
  XNOR U10926 ( .A(n11162), .B(n11017), .Z(n11164) );
  IV U10927 ( .A(p_input[2693]), .Z(n11017) );
  XOR U10928 ( .A(n11166), .B(n11167), .Z(n11162) );
  AND U10929 ( .A(n11168), .B(n11169), .Z(n11167) );
  XNOR U10930 ( .A(p_input[2708]), .B(n11166), .Z(n11169) );
  XNOR U10931 ( .A(n11166), .B(n11026), .Z(n11168) );
  IV U10932 ( .A(p_input[2692]), .Z(n11026) );
  XOR U10933 ( .A(n11170), .B(n11171), .Z(n11166) );
  AND U10934 ( .A(n11172), .B(n11173), .Z(n11171) );
  XNOR U10935 ( .A(p_input[2707]), .B(n11170), .Z(n11173) );
  XNOR U10936 ( .A(n11170), .B(n11035), .Z(n11172) );
  IV U10937 ( .A(p_input[2691]), .Z(n11035) );
  XOR U10938 ( .A(n11174), .B(n11175), .Z(n11170) );
  AND U10939 ( .A(n11176), .B(n11177), .Z(n11175) );
  XNOR U10940 ( .A(p_input[2706]), .B(n11174), .Z(n11177) );
  XNOR U10941 ( .A(n11174), .B(n11044), .Z(n11176) );
  IV U10942 ( .A(p_input[2690]), .Z(n11044) );
  XNOR U10943 ( .A(n11178), .B(n11179), .Z(n11174) );
  AND U10944 ( .A(n11180), .B(n11181), .Z(n11179) );
  XOR U10945 ( .A(p_input[2705]), .B(n11178), .Z(n11181) );
  XNOR U10946 ( .A(p_input[2689]), .B(n11178), .Z(n11180) );
  AND U10947 ( .A(p_input[2704]), .B(n11182), .Z(n11178) );
  IV U10948 ( .A(p_input[2688]), .Z(n11182) );
  XOR U10949 ( .A(n11183), .B(n11184), .Z(n10298) );
  AND U10950 ( .A(n764), .B(n11185), .Z(n11184) );
  XNOR U10951 ( .A(n11186), .B(n11183), .Z(n11185) );
  XOR U10952 ( .A(n11187), .B(n11188), .Z(n764) );
  AND U10953 ( .A(n11189), .B(n11190), .Z(n11188) );
  XNOR U10954 ( .A(n10310), .B(n11187), .Z(n11190) );
  AND U10955 ( .A(n11191), .B(n11192), .Z(n10310) );
  XOR U10956 ( .A(n11187), .B(n10309), .Z(n11189) );
  AND U10957 ( .A(n11193), .B(n11194), .Z(n10309) );
  XOR U10958 ( .A(n11195), .B(n11196), .Z(n11187) );
  AND U10959 ( .A(n11197), .B(n11198), .Z(n11196) );
  XOR U10960 ( .A(n11195), .B(n10322), .Z(n11198) );
  XOR U10961 ( .A(n11199), .B(n11200), .Z(n10322) );
  AND U10962 ( .A(n435), .B(n11201), .Z(n11200) );
  XOR U10963 ( .A(n11202), .B(n11199), .Z(n11201) );
  XNOR U10964 ( .A(n10319), .B(n11195), .Z(n11197) );
  XOR U10965 ( .A(n11203), .B(n11204), .Z(n10319) );
  AND U10966 ( .A(n432), .B(n11205), .Z(n11204) );
  XOR U10967 ( .A(n11206), .B(n11203), .Z(n11205) );
  XOR U10968 ( .A(n11207), .B(n11208), .Z(n11195) );
  AND U10969 ( .A(n11209), .B(n11210), .Z(n11208) );
  XOR U10970 ( .A(n11207), .B(n10334), .Z(n11210) );
  XOR U10971 ( .A(n11211), .B(n11212), .Z(n10334) );
  AND U10972 ( .A(n435), .B(n11213), .Z(n11212) );
  XOR U10973 ( .A(n11214), .B(n11211), .Z(n11213) );
  XNOR U10974 ( .A(n10331), .B(n11207), .Z(n11209) );
  XOR U10975 ( .A(n11215), .B(n11216), .Z(n10331) );
  AND U10976 ( .A(n432), .B(n11217), .Z(n11216) );
  XOR U10977 ( .A(n11218), .B(n11215), .Z(n11217) );
  XOR U10978 ( .A(n11219), .B(n11220), .Z(n11207) );
  AND U10979 ( .A(n11221), .B(n11222), .Z(n11220) );
  XOR U10980 ( .A(n11219), .B(n10346), .Z(n11222) );
  XOR U10981 ( .A(n11223), .B(n11224), .Z(n10346) );
  AND U10982 ( .A(n435), .B(n11225), .Z(n11224) );
  XOR U10983 ( .A(n11226), .B(n11223), .Z(n11225) );
  XNOR U10984 ( .A(n10343), .B(n11219), .Z(n11221) );
  XOR U10985 ( .A(n11227), .B(n11228), .Z(n10343) );
  AND U10986 ( .A(n432), .B(n11229), .Z(n11228) );
  XOR U10987 ( .A(n11230), .B(n11227), .Z(n11229) );
  XOR U10988 ( .A(n11231), .B(n11232), .Z(n11219) );
  AND U10989 ( .A(n11233), .B(n11234), .Z(n11232) );
  XOR U10990 ( .A(n11231), .B(n10358), .Z(n11234) );
  XOR U10991 ( .A(n11235), .B(n11236), .Z(n10358) );
  AND U10992 ( .A(n435), .B(n11237), .Z(n11236) );
  XOR U10993 ( .A(n11238), .B(n11235), .Z(n11237) );
  XNOR U10994 ( .A(n10355), .B(n11231), .Z(n11233) );
  XOR U10995 ( .A(n11239), .B(n11240), .Z(n10355) );
  AND U10996 ( .A(n432), .B(n11241), .Z(n11240) );
  XOR U10997 ( .A(n11242), .B(n11239), .Z(n11241) );
  XOR U10998 ( .A(n11243), .B(n11244), .Z(n11231) );
  AND U10999 ( .A(n11245), .B(n11246), .Z(n11244) );
  XOR U11000 ( .A(n11243), .B(n10370), .Z(n11246) );
  XOR U11001 ( .A(n11247), .B(n11248), .Z(n10370) );
  AND U11002 ( .A(n435), .B(n11249), .Z(n11248) );
  XOR U11003 ( .A(n11250), .B(n11247), .Z(n11249) );
  XNOR U11004 ( .A(n10367), .B(n11243), .Z(n11245) );
  XOR U11005 ( .A(n11251), .B(n11252), .Z(n10367) );
  AND U11006 ( .A(n432), .B(n11253), .Z(n11252) );
  XOR U11007 ( .A(n11254), .B(n11251), .Z(n11253) );
  XOR U11008 ( .A(n11255), .B(n11256), .Z(n11243) );
  AND U11009 ( .A(n11257), .B(n11258), .Z(n11256) );
  XOR U11010 ( .A(n11255), .B(n10382), .Z(n11258) );
  XOR U11011 ( .A(n11259), .B(n11260), .Z(n10382) );
  AND U11012 ( .A(n435), .B(n11261), .Z(n11260) );
  XOR U11013 ( .A(n11262), .B(n11259), .Z(n11261) );
  XNOR U11014 ( .A(n10379), .B(n11255), .Z(n11257) );
  XOR U11015 ( .A(n11263), .B(n11264), .Z(n10379) );
  AND U11016 ( .A(n432), .B(n11265), .Z(n11264) );
  XOR U11017 ( .A(n11266), .B(n11263), .Z(n11265) );
  XOR U11018 ( .A(n11267), .B(n11268), .Z(n11255) );
  AND U11019 ( .A(n11269), .B(n11270), .Z(n11268) );
  XOR U11020 ( .A(n11267), .B(n10394), .Z(n11270) );
  XOR U11021 ( .A(n11271), .B(n11272), .Z(n10394) );
  AND U11022 ( .A(n435), .B(n11273), .Z(n11272) );
  XOR U11023 ( .A(n11274), .B(n11271), .Z(n11273) );
  XNOR U11024 ( .A(n10391), .B(n11267), .Z(n11269) );
  XOR U11025 ( .A(n11275), .B(n11276), .Z(n10391) );
  AND U11026 ( .A(n432), .B(n11277), .Z(n11276) );
  XOR U11027 ( .A(n11278), .B(n11275), .Z(n11277) );
  XOR U11028 ( .A(n11279), .B(n11280), .Z(n11267) );
  AND U11029 ( .A(n11281), .B(n11282), .Z(n11280) );
  XOR U11030 ( .A(n11279), .B(n10406), .Z(n11282) );
  XOR U11031 ( .A(n11283), .B(n11284), .Z(n10406) );
  AND U11032 ( .A(n435), .B(n11285), .Z(n11284) );
  XOR U11033 ( .A(n11286), .B(n11283), .Z(n11285) );
  XNOR U11034 ( .A(n10403), .B(n11279), .Z(n11281) );
  XOR U11035 ( .A(n11287), .B(n11288), .Z(n10403) );
  AND U11036 ( .A(n432), .B(n11289), .Z(n11288) );
  XOR U11037 ( .A(n11290), .B(n11287), .Z(n11289) );
  XOR U11038 ( .A(n11291), .B(n11292), .Z(n11279) );
  AND U11039 ( .A(n11293), .B(n11294), .Z(n11292) );
  XOR U11040 ( .A(n11291), .B(n10418), .Z(n11294) );
  XOR U11041 ( .A(n11295), .B(n11296), .Z(n10418) );
  AND U11042 ( .A(n435), .B(n11297), .Z(n11296) );
  XOR U11043 ( .A(n11298), .B(n11295), .Z(n11297) );
  XNOR U11044 ( .A(n10415), .B(n11291), .Z(n11293) );
  XOR U11045 ( .A(n11299), .B(n11300), .Z(n10415) );
  AND U11046 ( .A(n432), .B(n11301), .Z(n11300) );
  XOR U11047 ( .A(n11302), .B(n11299), .Z(n11301) );
  XOR U11048 ( .A(n11303), .B(n11304), .Z(n11291) );
  AND U11049 ( .A(n11305), .B(n11306), .Z(n11304) );
  XOR U11050 ( .A(n11303), .B(n10430), .Z(n11306) );
  XOR U11051 ( .A(n11307), .B(n11308), .Z(n10430) );
  AND U11052 ( .A(n435), .B(n11309), .Z(n11308) );
  XOR U11053 ( .A(n11310), .B(n11307), .Z(n11309) );
  XNOR U11054 ( .A(n10427), .B(n11303), .Z(n11305) );
  XOR U11055 ( .A(n11311), .B(n11312), .Z(n10427) );
  AND U11056 ( .A(n432), .B(n11313), .Z(n11312) );
  XOR U11057 ( .A(n11314), .B(n11311), .Z(n11313) );
  XOR U11058 ( .A(n11315), .B(n11316), .Z(n11303) );
  AND U11059 ( .A(n11317), .B(n11318), .Z(n11316) );
  XOR U11060 ( .A(n11315), .B(n10442), .Z(n11318) );
  XOR U11061 ( .A(n11319), .B(n11320), .Z(n10442) );
  AND U11062 ( .A(n435), .B(n11321), .Z(n11320) );
  XOR U11063 ( .A(n11322), .B(n11319), .Z(n11321) );
  XNOR U11064 ( .A(n10439), .B(n11315), .Z(n11317) );
  XOR U11065 ( .A(n11323), .B(n11324), .Z(n10439) );
  AND U11066 ( .A(n432), .B(n11325), .Z(n11324) );
  XOR U11067 ( .A(n11326), .B(n11323), .Z(n11325) );
  XOR U11068 ( .A(n11327), .B(n11328), .Z(n11315) );
  AND U11069 ( .A(n11329), .B(n11330), .Z(n11328) );
  XOR U11070 ( .A(n11327), .B(n10454), .Z(n11330) );
  XOR U11071 ( .A(n11331), .B(n11332), .Z(n10454) );
  AND U11072 ( .A(n435), .B(n11333), .Z(n11332) );
  XOR U11073 ( .A(n11334), .B(n11331), .Z(n11333) );
  XNOR U11074 ( .A(n10451), .B(n11327), .Z(n11329) );
  XOR U11075 ( .A(n11335), .B(n11336), .Z(n10451) );
  AND U11076 ( .A(n432), .B(n11337), .Z(n11336) );
  XOR U11077 ( .A(n11338), .B(n11335), .Z(n11337) );
  XOR U11078 ( .A(n11339), .B(n11340), .Z(n11327) );
  AND U11079 ( .A(n11341), .B(n11342), .Z(n11340) );
  XOR U11080 ( .A(n11339), .B(n10466), .Z(n11342) );
  XOR U11081 ( .A(n11343), .B(n11344), .Z(n10466) );
  AND U11082 ( .A(n435), .B(n11345), .Z(n11344) );
  XOR U11083 ( .A(n11346), .B(n11343), .Z(n11345) );
  XNOR U11084 ( .A(n10463), .B(n11339), .Z(n11341) );
  XOR U11085 ( .A(n11347), .B(n11348), .Z(n10463) );
  AND U11086 ( .A(n432), .B(n11349), .Z(n11348) );
  XOR U11087 ( .A(n11350), .B(n11347), .Z(n11349) );
  XOR U11088 ( .A(n11351), .B(n11352), .Z(n11339) );
  AND U11089 ( .A(n11353), .B(n11354), .Z(n11352) );
  XNOR U11090 ( .A(n11355), .B(n10479), .Z(n11354) );
  XOR U11091 ( .A(n11356), .B(n11357), .Z(n10479) );
  AND U11092 ( .A(n435), .B(n11358), .Z(n11357) );
  XOR U11093 ( .A(n11356), .B(n11359), .Z(n11358) );
  XNOR U11094 ( .A(n10476), .B(n11351), .Z(n11353) );
  XOR U11095 ( .A(n11360), .B(n11361), .Z(n10476) );
  AND U11096 ( .A(n432), .B(n11362), .Z(n11361) );
  XOR U11097 ( .A(n11360), .B(n11363), .Z(n11362) );
  IV U11098 ( .A(n11355), .Z(n11351) );
  AND U11099 ( .A(n11183), .B(n11186), .Z(n11355) );
  XNOR U11100 ( .A(n11364), .B(n11365), .Z(n11186) );
  AND U11101 ( .A(n435), .B(n11366), .Z(n11365) );
  XNOR U11102 ( .A(n11367), .B(n11364), .Z(n11366) );
  XOR U11103 ( .A(n11368), .B(n11369), .Z(n435) );
  AND U11104 ( .A(n11370), .B(n11371), .Z(n11369) );
  XNOR U11105 ( .A(n11191), .B(n11368), .Z(n11371) );
  AND U11106 ( .A(p_input[2687]), .B(p_input[2671]), .Z(n11191) );
  XOR U11107 ( .A(n11368), .B(n11192), .Z(n11370) );
  AND U11108 ( .A(p_input[2655]), .B(p_input[2639]), .Z(n11192) );
  XOR U11109 ( .A(n11372), .B(n11373), .Z(n11368) );
  AND U11110 ( .A(n11374), .B(n11375), .Z(n11373) );
  XOR U11111 ( .A(n11372), .B(n11202), .Z(n11375) );
  XNOR U11112 ( .A(p_input[2670]), .B(n11376), .Z(n11202) );
  AND U11113 ( .A(n271), .B(n11377), .Z(n11376) );
  XOR U11114 ( .A(p_input[2686]), .B(p_input[2670]), .Z(n11377) );
  XNOR U11115 ( .A(n11199), .B(n11372), .Z(n11374) );
  XOR U11116 ( .A(n11378), .B(n11379), .Z(n11199) );
  AND U11117 ( .A(n269), .B(n11380), .Z(n11379) );
  XOR U11118 ( .A(p_input[2654]), .B(p_input[2638]), .Z(n11380) );
  XOR U11119 ( .A(n11381), .B(n11382), .Z(n11372) );
  AND U11120 ( .A(n11383), .B(n11384), .Z(n11382) );
  XOR U11121 ( .A(n11381), .B(n11214), .Z(n11384) );
  XNOR U11122 ( .A(p_input[2669]), .B(n11385), .Z(n11214) );
  AND U11123 ( .A(n271), .B(n11386), .Z(n11385) );
  XOR U11124 ( .A(p_input[2685]), .B(p_input[2669]), .Z(n11386) );
  XNOR U11125 ( .A(n11211), .B(n11381), .Z(n11383) );
  XOR U11126 ( .A(n11387), .B(n11388), .Z(n11211) );
  AND U11127 ( .A(n269), .B(n11389), .Z(n11388) );
  XOR U11128 ( .A(p_input[2653]), .B(p_input[2637]), .Z(n11389) );
  XOR U11129 ( .A(n11390), .B(n11391), .Z(n11381) );
  AND U11130 ( .A(n11392), .B(n11393), .Z(n11391) );
  XOR U11131 ( .A(n11390), .B(n11226), .Z(n11393) );
  XNOR U11132 ( .A(p_input[2668]), .B(n11394), .Z(n11226) );
  AND U11133 ( .A(n271), .B(n11395), .Z(n11394) );
  XOR U11134 ( .A(p_input[2684]), .B(p_input[2668]), .Z(n11395) );
  XNOR U11135 ( .A(n11223), .B(n11390), .Z(n11392) );
  XOR U11136 ( .A(n11396), .B(n11397), .Z(n11223) );
  AND U11137 ( .A(n269), .B(n11398), .Z(n11397) );
  XOR U11138 ( .A(p_input[2652]), .B(p_input[2636]), .Z(n11398) );
  XOR U11139 ( .A(n11399), .B(n11400), .Z(n11390) );
  AND U11140 ( .A(n11401), .B(n11402), .Z(n11400) );
  XOR U11141 ( .A(n11399), .B(n11238), .Z(n11402) );
  XNOR U11142 ( .A(p_input[2667]), .B(n11403), .Z(n11238) );
  AND U11143 ( .A(n271), .B(n11404), .Z(n11403) );
  XOR U11144 ( .A(p_input[2683]), .B(p_input[2667]), .Z(n11404) );
  XNOR U11145 ( .A(n11235), .B(n11399), .Z(n11401) );
  XOR U11146 ( .A(n11405), .B(n11406), .Z(n11235) );
  AND U11147 ( .A(n269), .B(n11407), .Z(n11406) );
  XOR U11148 ( .A(p_input[2651]), .B(p_input[2635]), .Z(n11407) );
  XOR U11149 ( .A(n11408), .B(n11409), .Z(n11399) );
  AND U11150 ( .A(n11410), .B(n11411), .Z(n11409) );
  XOR U11151 ( .A(n11408), .B(n11250), .Z(n11411) );
  XNOR U11152 ( .A(p_input[2666]), .B(n11412), .Z(n11250) );
  AND U11153 ( .A(n271), .B(n11413), .Z(n11412) );
  XOR U11154 ( .A(p_input[2682]), .B(p_input[2666]), .Z(n11413) );
  XNOR U11155 ( .A(n11247), .B(n11408), .Z(n11410) );
  XOR U11156 ( .A(n11414), .B(n11415), .Z(n11247) );
  AND U11157 ( .A(n269), .B(n11416), .Z(n11415) );
  XOR U11158 ( .A(p_input[2650]), .B(p_input[2634]), .Z(n11416) );
  XOR U11159 ( .A(n11417), .B(n11418), .Z(n11408) );
  AND U11160 ( .A(n11419), .B(n11420), .Z(n11418) );
  XOR U11161 ( .A(n11417), .B(n11262), .Z(n11420) );
  XNOR U11162 ( .A(p_input[2665]), .B(n11421), .Z(n11262) );
  AND U11163 ( .A(n271), .B(n11422), .Z(n11421) );
  XOR U11164 ( .A(p_input[2681]), .B(p_input[2665]), .Z(n11422) );
  XNOR U11165 ( .A(n11259), .B(n11417), .Z(n11419) );
  XOR U11166 ( .A(n11423), .B(n11424), .Z(n11259) );
  AND U11167 ( .A(n269), .B(n11425), .Z(n11424) );
  XOR U11168 ( .A(p_input[2649]), .B(p_input[2633]), .Z(n11425) );
  XOR U11169 ( .A(n11426), .B(n11427), .Z(n11417) );
  AND U11170 ( .A(n11428), .B(n11429), .Z(n11427) );
  XOR U11171 ( .A(n11426), .B(n11274), .Z(n11429) );
  XNOR U11172 ( .A(p_input[2664]), .B(n11430), .Z(n11274) );
  AND U11173 ( .A(n271), .B(n11431), .Z(n11430) );
  XOR U11174 ( .A(p_input[2680]), .B(p_input[2664]), .Z(n11431) );
  XNOR U11175 ( .A(n11271), .B(n11426), .Z(n11428) );
  XOR U11176 ( .A(n11432), .B(n11433), .Z(n11271) );
  AND U11177 ( .A(n269), .B(n11434), .Z(n11433) );
  XOR U11178 ( .A(p_input[2648]), .B(p_input[2632]), .Z(n11434) );
  XOR U11179 ( .A(n11435), .B(n11436), .Z(n11426) );
  AND U11180 ( .A(n11437), .B(n11438), .Z(n11436) );
  XOR U11181 ( .A(n11435), .B(n11286), .Z(n11438) );
  XNOR U11182 ( .A(p_input[2663]), .B(n11439), .Z(n11286) );
  AND U11183 ( .A(n271), .B(n11440), .Z(n11439) );
  XOR U11184 ( .A(p_input[2679]), .B(p_input[2663]), .Z(n11440) );
  XNOR U11185 ( .A(n11283), .B(n11435), .Z(n11437) );
  XOR U11186 ( .A(n11441), .B(n11442), .Z(n11283) );
  AND U11187 ( .A(n269), .B(n11443), .Z(n11442) );
  XOR U11188 ( .A(p_input[2647]), .B(p_input[2631]), .Z(n11443) );
  XOR U11189 ( .A(n11444), .B(n11445), .Z(n11435) );
  AND U11190 ( .A(n11446), .B(n11447), .Z(n11445) );
  XOR U11191 ( .A(n11444), .B(n11298), .Z(n11447) );
  XNOR U11192 ( .A(p_input[2662]), .B(n11448), .Z(n11298) );
  AND U11193 ( .A(n271), .B(n11449), .Z(n11448) );
  XOR U11194 ( .A(p_input[2678]), .B(p_input[2662]), .Z(n11449) );
  XNOR U11195 ( .A(n11295), .B(n11444), .Z(n11446) );
  XOR U11196 ( .A(n11450), .B(n11451), .Z(n11295) );
  AND U11197 ( .A(n269), .B(n11452), .Z(n11451) );
  XOR U11198 ( .A(p_input[2646]), .B(p_input[2630]), .Z(n11452) );
  XOR U11199 ( .A(n11453), .B(n11454), .Z(n11444) );
  AND U11200 ( .A(n11455), .B(n11456), .Z(n11454) );
  XOR U11201 ( .A(n11453), .B(n11310), .Z(n11456) );
  XNOR U11202 ( .A(p_input[2661]), .B(n11457), .Z(n11310) );
  AND U11203 ( .A(n271), .B(n11458), .Z(n11457) );
  XOR U11204 ( .A(p_input[2677]), .B(p_input[2661]), .Z(n11458) );
  XNOR U11205 ( .A(n11307), .B(n11453), .Z(n11455) );
  XOR U11206 ( .A(n11459), .B(n11460), .Z(n11307) );
  AND U11207 ( .A(n269), .B(n11461), .Z(n11460) );
  XOR U11208 ( .A(p_input[2645]), .B(p_input[2629]), .Z(n11461) );
  XOR U11209 ( .A(n11462), .B(n11463), .Z(n11453) );
  AND U11210 ( .A(n11464), .B(n11465), .Z(n11463) );
  XOR U11211 ( .A(n11462), .B(n11322), .Z(n11465) );
  XNOR U11212 ( .A(p_input[2660]), .B(n11466), .Z(n11322) );
  AND U11213 ( .A(n271), .B(n11467), .Z(n11466) );
  XOR U11214 ( .A(p_input[2676]), .B(p_input[2660]), .Z(n11467) );
  XNOR U11215 ( .A(n11319), .B(n11462), .Z(n11464) );
  XOR U11216 ( .A(n11468), .B(n11469), .Z(n11319) );
  AND U11217 ( .A(n269), .B(n11470), .Z(n11469) );
  XOR U11218 ( .A(p_input[2644]), .B(p_input[2628]), .Z(n11470) );
  XOR U11219 ( .A(n11471), .B(n11472), .Z(n11462) );
  AND U11220 ( .A(n11473), .B(n11474), .Z(n11472) );
  XOR U11221 ( .A(n11471), .B(n11334), .Z(n11474) );
  XNOR U11222 ( .A(p_input[2659]), .B(n11475), .Z(n11334) );
  AND U11223 ( .A(n271), .B(n11476), .Z(n11475) );
  XOR U11224 ( .A(p_input[2675]), .B(p_input[2659]), .Z(n11476) );
  XNOR U11225 ( .A(n11331), .B(n11471), .Z(n11473) );
  XOR U11226 ( .A(n11477), .B(n11478), .Z(n11331) );
  AND U11227 ( .A(n269), .B(n11479), .Z(n11478) );
  XOR U11228 ( .A(p_input[2643]), .B(p_input[2627]), .Z(n11479) );
  XOR U11229 ( .A(n11480), .B(n11481), .Z(n11471) );
  AND U11230 ( .A(n11482), .B(n11483), .Z(n11481) );
  XOR U11231 ( .A(n11480), .B(n11346), .Z(n11483) );
  XNOR U11232 ( .A(p_input[2658]), .B(n11484), .Z(n11346) );
  AND U11233 ( .A(n271), .B(n11485), .Z(n11484) );
  XOR U11234 ( .A(p_input[2674]), .B(p_input[2658]), .Z(n11485) );
  XNOR U11235 ( .A(n11343), .B(n11480), .Z(n11482) );
  XOR U11236 ( .A(n11486), .B(n11487), .Z(n11343) );
  AND U11237 ( .A(n269), .B(n11488), .Z(n11487) );
  XOR U11238 ( .A(p_input[2642]), .B(p_input[2626]), .Z(n11488) );
  XOR U11239 ( .A(n11489), .B(n11490), .Z(n11480) );
  AND U11240 ( .A(n11491), .B(n11492), .Z(n11490) );
  XNOR U11241 ( .A(n11493), .B(n11359), .Z(n11492) );
  XNOR U11242 ( .A(p_input[2657]), .B(n11494), .Z(n11359) );
  AND U11243 ( .A(n271), .B(n11495), .Z(n11494) );
  XNOR U11244 ( .A(p_input[2673]), .B(n11496), .Z(n11495) );
  IV U11245 ( .A(p_input[2657]), .Z(n11496) );
  XNOR U11246 ( .A(n11356), .B(n11489), .Z(n11491) );
  XNOR U11247 ( .A(p_input[2625]), .B(n11497), .Z(n11356) );
  AND U11248 ( .A(n269), .B(n11498), .Z(n11497) );
  XOR U11249 ( .A(p_input[2641]), .B(p_input[2625]), .Z(n11498) );
  IV U11250 ( .A(n11493), .Z(n11489) );
  AND U11251 ( .A(n11364), .B(n11367), .Z(n11493) );
  XOR U11252 ( .A(p_input[2656]), .B(n11499), .Z(n11367) );
  AND U11253 ( .A(n271), .B(n11500), .Z(n11499) );
  XOR U11254 ( .A(p_input[2672]), .B(p_input[2656]), .Z(n11500) );
  XOR U11255 ( .A(n11501), .B(n11502), .Z(n271) );
  AND U11256 ( .A(n11503), .B(n11504), .Z(n11502) );
  XNOR U11257 ( .A(p_input[2687]), .B(n11501), .Z(n11504) );
  XOR U11258 ( .A(n11501), .B(p_input[2671]), .Z(n11503) );
  XOR U11259 ( .A(n11505), .B(n11506), .Z(n11501) );
  AND U11260 ( .A(n11507), .B(n11508), .Z(n11506) );
  XNOR U11261 ( .A(p_input[2686]), .B(n11505), .Z(n11508) );
  XOR U11262 ( .A(n11505), .B(p_input[2670]), .Z(n11507) );
  XOR U11263 ( .A(n11509), .B(n11510), .Z(n11505) );
  AND U11264 ( .A(n11511), .B(n11512), .Z(n11510) );
  XNOR U11265 ( .A(p_input[2685]), .B(n11509), .Z(n11512) );
  XOR U11266 ( .A(n11509), .B(p_input[2669]), .Z(n11511) );
  XOR U11267 ( .A(n11513), .B(n11514), .Z(n11509) );
  AND U11268 ( .A(n11515), .B(n11516), .Z(n11514) );
  XNOR U11269 ( .A(p_input[2684]), .B(n11513), .Z(n11516) );
  XOR U11270 ( .A(n11513), .B(p_input[2668]), .Z(n11515) );
  XOR U11271 ( .A(n11517), .B(n11518), .Z(n11513) );
  AND U11272 ( .A(n11519), .B(n11520), .Z(n11518) );
  XNOR U11273 ( .A(p_input[2683]), .B(n11517), .Z(n11520) );
  XOR U11274 ( .A(n11517), .B(p_input[2667]), .Z(n11519) );
  XOR U11275 ( .A(n11521), .B(n11522), .Z(n11517) );
  AND U11276 ( .A(n11523), .B(n11524), .Z(n11522) );
  XNOR U11277 ( .A(p_input[2682]), .B(n11521), .Z(n11524) );
  XOR U11278 ( .A(n11521), .B(p_input[2666]), .Z(n11523) );
  XOR U11279 ( .A(n11525), .B(n11526), .Z(n11521) );
  AND U11280 ( .A(n11527), .B(n11528), .Z(n11526) );
  XNOR U11281 ( .A(p_input[2681]), .B(n11525), .Z(n11528) );
  XOR U11282 ( .A(n11525), .B(p_input[2665]), .Z(n11527) );
  XOR U11283 ( .A(n11529), .B(n11530), .Z(n11525) );
  AND U11284 ( .A(n11531), .B(n11532), .Z(n11530) );
  XNOR U11285 ( .A(p_input[2680]), .B(n11529), .Z(n11532) );
  XOR U11286 ( .A(n11529), .B(p_input[2664]), .Z(n11531) );
  XOR U11287 ( .A(n11533), .B(n11534), .Z(n11529) );
  AND U11288 ( .A(n11535), .B(n11536), .Z(n11534) );
  XNOR U11289 ( .A(p_input[2679]), .B(n11533), .Z(n11536) );
  XOR U11290 ( .A(n11533), .B(p_input[2663]), .Z(n11535) );
  XOR U11291 ( .A(n11537), .B(n11538), .Z(n11533) );
  AND U11292 ( .A(n11539), .B(n11540), .Z(n11538) );
  XNOR U11293 ( .A(p_input[2678]), .B(n11537), .Z(n11540) );
  XOR U11294 ( .A(n11537), .B(p_input[2662]), .Z(n11539) );
  XOR U11295 ( .A(n11541), .B(n11542), .Z(n11537) );
  AND U11296 ( .A(n11543), .B(n11544), .Z(n11542) );
  XNOR U11297 ( .A(p_input[2677]), .B(n11541), .Z(n11544) );
  XOR U11298 ( .A(n11541), .B(p_input[2661]), .Z(n11543) );
  XOR U11299 ( .A(n11545), .B(n11546), .Z(n11541) );
  AND U11300 ( .A(n11547), .B(n11548), .Z(n11546) );
  XNOR U11301 ( .A(p_input[2676]), .B(n11545), .Z(n11548) );
  XOR U11302 ( .A(n11545), .B(p_input[2660]), .Z(n11547) );
  XOR U11303 ( .A(n11549), .B(n11550), .Z(n11545) );
  AND U11304 ( .A(n11551), .B(n11552), .Z(n11550) );
  XNOR U11305 ( .A(p_input[2675]), .B(n11549), .Z(n11552) );
  XOR U11306 ( .A(n11549), .B(p_input[2659]), .Z(n11551) );
  XOR U11307 ( .A(n11553), .B(n11554), .Z(n11549) );
  AND U11308 ( .A(n11555), .B(n11556), .Z(n11554) );
  XNOR U11309 ( .A(p_input[2674]), .B(n11553), .Z(n11556) );
  XOR U11310 ( .A(n11553), .B(p_input[2658]), .Z(n11555) );
  XNOR U11311 ( .A(n11557), .B(n11558), .Z(n11553) );
  AND U11312 ( .A(n11559), .B(n11560), .Z(n11558) );
  XOR U11313 ( .A(p_input[2673]), .B(n11557), .Z(n11560) );
  XNOR U11314 ( .A(p_input[2657]), .B(n11557), .Z(n11559) );
  AND U11315 ( .A(p_input[2672]), .B(n11561), .Z(n11557) );
  IV U11316 ( .A(p_input[2656]), .Z(n11561) );
  XNOR U11317 ( .A(p_input[2624]), .B(n11562), .Z(n11364) );
  AND U11318 ( .A(n269), .B(n11563), .Z(n11562) );
  XOR U11319 ( .A(p_input[2640]), .B(p_input[2624]), .Z(n11563) );
  XOR U11320 ( .A(n11564), .B(n11565), .Z(n269) );
  AND U11321 ( .A(n11566), .B(n11567), .Z(n11565) );
  XNOR U11322 ( .A(p_input[2655]), .B(n11564), .Z(n11567) );
  XOR U11323 ( .A(n11564), .B(p_input[2639]), .Z(n11566) );
  XOR U11324 ( .A(n11568), .B(n11569), .Z(n11564) );
  AND U11325 ( .A(n11570), .B(n11571), .Z(n11569) );
  XNOR U11326 ( .A(p_input[2654]), .B(n11568), .Z(n11571) );
  XNOR U11327 ( .A(n11568), .B(n11378), .Z(n11570) );
  IV U11328 ( .A(p_input[2638]), .Z(n11378) );
  XOR U11329 ( .A(n11572), .B(n11573), .Z(n11568) );
  AND U11330 ( .A(n11574), .B(n11575), .Z(n11573) );
  XNOR U11331 ( .A(p_input[2653]), .B(n11572), .Z(n11575) );
  XNOR U11332 ( .A(n11572), .B(n11387), .Z(n11574) );
  IV U11333 ( .A(p_input[2637]), .Z(n11387) );
  XOR U11334 ( .A(n11576), .B(n11577), .Z(n11572) );
  AND U11335 ( .A(n11578), .B(n11579), .Z(n11577) );
  XNOR U11336 ( .A(p_input[2652]), .B(n11576), .Z(n11579) );
  XNOR U11337 ( .A(n11576), .B(n11396), .Z(n11578) );
  IV U11338 ( .A(p_input[2636]), .Z(n11396) );
  XOR U11339 ( .A(n11580), .B(n11581), .Z(n11576) );
  AND U11340 ( .A(n11582), .B(n11583), .Z(n11581) );
  XNOR U11341 ( .A(p_input[2651]), .B(n11580), .Z(n11583) );
  XNOR U11342 ( .A(n11580), .B(n11405), .Z(n11582) );
  IV U11343 ( .A(p_input[2635]), .Z(n11405) );
  XOR U11344 ( .A(n11584), .B(n11585), .Z(n11580) );
  AND U11345 ( .A(n11586), .B(n11587), .Z(n11585) );
  XNOR U11346 ( .A(p_input[2650]), .B(n11584), .Z(n11587) );
  XNOR U11347 ( .A(n11584), .B(n11414), .Z(n11586) );
  IV U11348 ( .A(p_input[2634]), .Z(n11414) );
  XOR U11349 ( .A(n11588), .B(n11589), .Z(n11584) );
  AND U11350 ( .A(n11590), .B(n11591), .Z(n11589) );
  XNOR U11351 ( .A(p_input[2649]), .B(n11588), .Z(n11591) );
  XNOR U11352 ( .A(n11588), .B(n11423), .Z(n11590) );
  IV U11353 ( .A(p_input[2633]), .Z(n11423) );
  XOR U11354 ( .A(n11592), .B(n11593), .Z(n11588) );
  AND U11355 ( .A(n11594), .B(n11595), .Z(n11593) );
  XNOR U11356 ( .A(p_input[2648]), .B(n11592), .Z(n11595) );
  XNOR U11357 ( .A(n11592), .B(n11432), .Z(n11594) );
  IV U11358 ( .A(p_input[2632]), .Z(n11432) );
  XOR U11359 ( .A(n11596), .B(n11597), .Z(n11592) );
  AND U11360 ( .A(n11598), .B(n11599), .Z(n11597) );
  XNOR U11361 ( .A(p_input[2647]), .B(n11596), .Z(n11599) );
  XNOR U11362 ( .A(n11596), .B(n11441), .Z(n11598) );
  IV U11363 ( .A(p_input[2631]), .Z(n11441) );
  XOR U11364 ( .A(n11600), .B(n11601), .Z(n11596) );
  AND U11365 ( .A(n11602), .B(n11603), .Z(n11601) );
  XNOR U11366 ( .A(p_input[2646]), .B(n11600), .Z(n11603) );
  XNOR U11367 ( .A(n11600), .B(n11450), .Z(n11602) );
  IV U11368 ( .A(p_input[2630]), .Z(n11450) );
  XOR U11369 ( .A(n11604), .B(n11605), .Z(n11600) );
  AND U11370 ( .A(n11606), .B(n11607), .Z(n11605) );
  XNOR U11371 ( .A(p_input[2645]), .B(n11604), .Z(n11607) );
  XNOR U11372 ( .A(n11604), .B(n11459), .Z(n11606) );
  IV U11373 ( .A(p_input[2629]), .Z(n11459) );
  XOR U11374 ( .A(n11608), .B(n11609), .Z(n11604) );
  AND U11375 ( .A(n11610), .B(n11611), .Z(n11609) );
  XNOR U11376 ( .A(p_input[2644]), .B(n11608), .Z(n11611) );
  XNOR U11377 ( .A(n11608), .B(n11468), .Z(n11610) );
  IV U11378 ( .A(p_input[2628]), .Z(n11468) );
  XOR U11379 ( .A(n11612), .B(n11613), .Z(n11608) );
  AND U11380 ( .A(n11614), .B(n11615), .Z(n11613) );
  XNOR U11381 ( .A(p_input[2643]), .B(n11612), .Z(n11615) );
  XNOR U11382 ( .A(n11612), .B(n11477), .Z(n11614) );
  IV U11383 ( .A(p_input[2627]), .Z(n11477) );
  XOR U11384 ( .A(n11616), .B(n11617), .Z(n11612) );
  AND U11385 ( .A(n11618), .B(n11619), .Z(n11617) );
  XNOR U11386 ( .A(p_input[2642]), .B(n11616), .Z(n11619) );
  XNOR U11387 ( .A(n11616), .B(n11486), .Z(n11618) );
  IV U11388 ( .A(p_input[2626]), .Z(n11486) );
  XNOR U11389 ( .A(n11620), .B(n11621), .Z(n11616) );
  AND U11390 ( .A(n11622), .B(n11623), .Z(n11621) );
  XOR U11391 ( .A(p_input[2641]), .B(n11620), .Z(n11623) );
  XNOR U11392 ( .A(p_input[2625]), .B(n11620), .Z(n11622) );
  AND U11393 ( .A(p_input[2640]), .B(n11624), .Z(n11620) );
  IV U11394 ( .A(p_input[2624]), .Z(n11624) );
  XOR U11395 ( .A(n11625), .B(n11626), .Z(n11183) );
  AND U11396 ( .A(n432), .B(n11627), .Z(n11626) );
  XNOR U11397 ( .A(n11628), .B(n11625), .Z(n11627) );
  XOR U11398 ( .A(n11629), .B(n11630), .Z(n432) );
  AND U11399 ( .A(n11631), .B(n11632), .Z(n11630) );
  XNOR U11400 ( .A(n11194), .B(n11629), .Z(n11632) );
  AND U11401 ( .A(p_input[2623]), .B(p_input[2607]), .Z(n11194) );
  XOR U11402 ( .A(n11629), .B(n11193), .Z(n11631) );
  AND U11403 ( .A(p_input[2575]), .B(p_input[2591]), .Z(n11193) );
  XOR U11404 ( .A(n11633), .B(n11634), .Z(n11629) );
  AND U11405 ( .A(n11635), .B(n11636), .Z(n11634) );
  XOR U11406 ( .A(n11633), .B(n11206), .Z(n11636) );
  XNOR U11407 ( .A(p_input[2606]), .B(n11637), .Z(n11206) );
  AND U11408 ( .A(n275), .B(n11638), .Z(n11637) );
  XOR U11409 ( .A(p_input[2622]), .B(p_input[2606]), .Z(n11638) );
  XNOR U11410 ( .A(n11203), .B(n11633), .Z(n11635) );
  XOR U11411 ( .A(n11639), .B(n11640), .Z(n11203) );
  AND U11412 ( .A(n272), .B(n11641), .Z(n11640) );
  XOR U11413 ( .A(p_input[2590]), .B(p_input[2574]), .Z(n11641) );
  XOR U11414 ( .A(n11642), .B(n11643), .Z(n11633) );
  AND U11415 ( .A(n11644), .B(n11645), .Z(n11643) );
  XOR U11416 ( .A(n11642), .B(n11218), .Z(n11645) );
  XNOR U11417 ( .A(p_input[2605]), .B(n11646), .Z(n11218) );
  AND U11418 ( .A(n275), .B(n11647), .Z(n11646) );
  XOR U11419 ( .A(p_input[2621]), .B(p_input[2605]), .Z(n11647) );
  XNOR U11420 ( .A(n11215), .B(n11642), .Z(n11644) );
  XOR U11421 ( .A(n11648), .B(n11649), .Z(n11215) );
  AND U11422 ( .A(n272), .B(n11650), .Z(n11649) );
  XOR U11423 ( .A(p_input[2589]), .B(p_input[2573]), .Z(n11650) );
  XOR U11424 ( .A(n11651), .B(n11652), .Z(n11642) );
  AND U11425 ( .A(n11653), .B(n11654), .Z(n11652) );
  XOR U11426 ( .A(n11651), .B(n11230), .Z(n11654) );
  XNOR U11427 ( .A(p_input[2604]), .B(n11655), .Z(n11230) );
  AND U11428 ( .A(n275), .B(n11656), .Z(n11655) );
  XOR U11429 ( .A(p_input[2620]), .B(p_input[2604]), .Z(n11656) );
  XNOR U11430 ( .A(n11227), .B(n11651), .Z(n11653) );
  XOR U11431 ( .A(n11657), .B(n11658), .Z(n11227) );
  AND U11432 ( .A(n272), .B(n11659), .Z(n11658) );
  XOR U11433 ( .A(p_input[2588]), .B(p_input[2572]), .Z(n11659) );
  XOR U11434 ( .A(n11660), .B(n11661), .Z(n11651) );
  AND U11435 ( .A(n11662), .B(n11663), .Z(n11661) );
  XOR U11436 ( .A(n11660), .B(n11242), .Z(n11663) );
  XNOR U11437 ( .A(p_input[2603]), .B(n11664), .Z(n11242) );
  AND U11438 ( .A(n275), .B(n11665), .Z(n11664) );
  XOR U11439 ( .A(p_input[2619]), .B(p_input[2603]), .Z(n11665) );
  XNOR U11440 ( .A(n11239), .B(n11660), .Z(n11662) );
  XOR U11441 ( .A(n11666), .B(n11667), .Z(n11239) );
  AND U11442 ( .A(n272), .B(n11668), .Z(n11667) );
  XOR U11443 ( .A(p_input[2587]), .B(p_input[2571]), .Z(n11668) );
  XOR U11444 ( .A(n11669), .B(n11670), .Z(n11660) );
  AND U11445 ( .A(n11671), .B(n11672), .Z(n11670) );
  XOR U11446 ( .A(n11669), .B(n11254), .Z(n11672) );
  XNOR U11447 ( .A(p_input[2602]), .B(n11673), .Z(n11254) );
  AND U11448 ( .A(n275), .B(n11674), .Z(n11673) );
  XOR U11449 ( .A(p_input[2618]), .B(p_input[2602]), .Z(n11674) );
  XNOR U11450 ( .A(n11251), .B(n11669), .Z(n11671) );
  XOR U11451 ( .A(n11675), .B(n11676), .Z(n11251) );
  AND U11452 ( .A(n272), .B(n11677), .Z(n11676) );
  XOR U11453 ( .A(p_input[2586]), .B(p_input[2570]), .Z(n11677) );
  XOR U11454 ( .A(n11678), .B(n11679), .Z(n11669) );
  AND U11455 ( .A(n11680), .B(n11681), .Z(n11679) );
  XOR U11456 ( .A(n11678), .B(n11266), .Z(n11681) );
  XNOR U11457 ( .A(p_input[2601]), .B(n11682), .Z(n11266) );
  AND U11458 ( .A(n275), .B(n11683), .Z(n11682) );
  XOR U11459 ( .A(p_input[2617]), .B(p_input[2601]), .Z(n11683) );
  XNOR U11460 ( .A(n11263), .B(n11678), .Z(n11680) );
  XOR U11461 ( .A(n11684), .B(n11685), .Z(n11263) );
  AND U11462 ( .A(n272), .B(n11686), .Z(n11685) );
  XOR U11463 ( .A(p_input[2585]), .B(p_input[2569]), .Z(n11686) );
  XOR U11464 ( .A(n11687), .B(n11688), .Z(n11678) );
  AND U11465 ( .A(n11689), .B(n11690), .Z(n11688) );
  XOR U11466 ( .A(n11687), .B(n11278), .Z(n11690) );
  XNOR U11467 ( .A(p_input[2600]), .B(n11691), .Z(n11278) );
  AND U11468 ( .A(n275), .B(n11692), .Z(n11691) );
  XOR U11469 ( .A(p_input[2616]), .B(p_input[2600]), .Z(n11692) );
  XNOR U11470 ( .A(n11275), .B(n11687), .Z(n11689) );
  XOR U11471 ( .A(n11693), .B(n11694), .Z(n11275) );
  AND U11472 ( .A(n272), .B(n11695), .Z(n11694) );
  XOR U11473 ( .A(p_input[2584]), .B(p_input[2568]), .Z(n11695) );
  XOR U11474 ( .A(n11696), .B(n11697), .Z(n11687) );
  AND U11475 ( .A(n11698), .B(n11699), .Z(n11697) );
  XOR U11476 ( .A(n11696), .B(n11290), .Z(n11699) );
  XNOR U11477 ( .A(p_input[2599]), .B(n11700), .Z(n11290) );
  AND U11478 ( .A(n275), .B(n11701), .Z(n11700) );
  XOR U11479 ( .A(p_input[2615]), .B(p_input[2599]), .Z(n11701) );
  XNOR U11480 ( .A(n11287), .B(n11696), .Z(n11698) );
  XOR U11481 ( .A(n11702), .B(n11703), .Z(n11287) );
  AND U11482 ( .A(n272), .B(n11704), .Z(n11703) );
  XOR U11483 ( .A(p_input[2583]), .B(p_input[2567]), .Z(n11704) );
  XOR U11484 ( .A(n11705), .B(n11706), .Z(n11696) );
  AND U11485 ( .A(n11707), .B(n11708), .Z(n11706) );
  XOR U11486 ( .A(n11705), .B(n11302), .Z(n11708) );
  XNOR U11487 ( .A(p_input[2598]), .B(n11709), .Z(n11302) );
  AND U11488 ( .A(n275), .B(n11710), .Z(n11709) );
  XOR U11489 ( .A(p_input[2614]), .B(p_input[2598]), .Z(n11710) );
  XNOR U11490 ( .A(n11299), .B(n11705), .Z(n11707) );
  XOR U11491 ( .A(n11711), .B(n11712), .Z(n11299) );
  AND U11492 ( .A(n272), .B(n11713), .Z(n11712) );
  XOR U11493 ( .A(p_input[2582]), .B(p_input[2566]), .Z(n11713) );
  XOR U11494 ( .A(n11714), .B(n11715), .Z(n11705) );
  AND U11495 ( .A(n11716), .B(n11717), .Z(n11715) );
  XOR U11496 ( .A(n11714), .B(n11314), .Z(n11717) );
  XNOR U11497 ( .A(p_input[2597]), .B(n11718), .Z(n11314) );
  AND U11498 ( .A(n275), .B(n11719), .Z(n11718) );
  XOR U11499 ( .A(p_input[2613]), .B(p_input[2597]), .Z(n11719) );
  XNOR U11500 ( .A(n11311), .B(n11714), .Z(n11716) );
  XOR U11501 ( .A(n11720), .B(n11721), .Z(n11311) );
  AND U11502 ( .A(n272), .B(n11722), .Z(n11721) );
  XOR U11503 ( .A(p_input[2581]), .B(p_input[2565]), .Z(n11722) );
  XOR U11504 ( .A(n11723), .B(n11724), .Z(n11714) );
  AND U11505 ( .A(n11725), .B(n11726), .Z(n11724) );
  XOR U11506 ( .A(n11723), .B(n11326), .Z(n11726) );
  XNOR U11507 ( .A(p_input[2596]), .B(n11727), .Z(n11326) );
  AND U11508 ( .A(n275), .B(n11728), .Z(n11727) );
  XOR U11509 ( .A(p_input[2612]), .B(p_input[2596]), .Z(n11728) );
  XNOR U11510 ( .A(n11323), .B(n11723), .Z(n11725) );
  XOR U11511 ( .A(n11729), .B(n11730), .Z(n11323) );
  AND U11512 ( .A(n272), .B(n11731), .Z(n11730) );
  XOR U11513 ( .A(p_input[2580]), .B(p_input[2564]), .Z(n11731) );
  XOR U11514 ( .A(n11732), .B(n11733), .Z(n11723) );
  AND U11515 ( .A(n11734), .B(n11735), .Z(n11733) );
  XOR U11516 ( .A(n11732), .B(n11338), .Z(n11735) );
  XNOR U11517 ( .A(p_input[2595]), .B(n11736), .Z(n11338) );
  AND U11518 ( .A(n275), .B(n11737), .Z(n11736) );
  XOR U11519 ( .A(p_input[2611]), .B(p_input[2595]), .Z(n11737) );
  XNOR U11520 ( .A(n11335), .B(n11732), .Z(n11734) );
  XOR U11521 ( .A(n11738), .B(n11739), .Z(n11335) );
  AND U11522 ( .A(n272), .B(n11740), .Z(n11739) );
  XOR U11523 ( .A(p_input[2579]), .B(p_input[2563]), .Z(n11740) );
  XOR U11524 ( .A(n11741), .B(n11742), .Z(n11732) );
  AND U11525 ( .A(n11743), .B(n11744), .Z(n11742) );
  XOR U11526 ( .A(n11741), .B(n11350), .Z(n11744) );
  XNOR U11527 ( .A(p_input[2594]), .B(n11745), .Z(n11350) );
  AND U11528 ( .A(n275), .B(n11746), .Z(n11745) );
  XOR U11529 ( .A(p_input[2610]), .B(p_input[2594]), .Z(n11746) );
  XNOR U11530 ( .A(n11347), .B(n11741), .Z(n11743) );
  XOR U11531 ( .A(n11747), .B(n11748), .Z(n11347) );
  AND U11532 ( .A(n272), .B(n11749), .Z(n11748) );
  XOR U11533 ( .A(p_input[2578]), .B(p_input[2562]), .Z(n11749) );
  XOR U11534 ( .A(n11750), .B(n11751), .Z(n11741) );
  AND U11535 ( .A(n11752), .B(n11753), .Z(n11751) );
  XNOR U11536 ( .A(n11754), .B(n11363), .Z(n11753) );
  XNOR U11537 ( .A(p_input[2593]), .B(n11755), .Z(n11363) );
  AND U11538 ( .A(n275), .B(n11756), .Z(n11755) );
  XNOR U11539 ( .A(p_input[2609]), .B(n11757), .Z(n11756) );
  IV U11540 ( .A(p_input[2593]), .Z(n11757) );
  XNOR U11541 ( .A(n11360), .B(n11750), .Z(n11752) );
  XNOR U11542 ( .A(p_input[2561]), .B(n11758), .Z(n11360) );
  AND U11543 ( .A(n272), .B(n11759), .Z(n11758) );
  XOR U11544 ( .A(p_input[2577]), .B(p_input[2561]), .Z(n11759) );
  IV U11545 ( .A(n11754), .Z(n11750) );
  AND U11546 ( .A(n11625), .B(n11628), .Z(n11754) );
  XOR U11547 ( .A(p_input[2592]), .B(n11760), .Z(n11628) );
  AND U11548 ( .A(n275), .B(n11761), .Z(n11760) );
  XOR U11549 ( .A(p_input[2608]), .B(p_input[2592]), .Z(n11761) );
  XOR U11550 ( .A(n11762), .B(n11763), .Z(n275) );
  AND U11551 ( .A(n11764), .B(n11765), .Z(n11763) );
  XNOR U11552 ( .A(p_input[2623]), .B(n11762), .Z(n11765) );
  XOR U11553 ( .A(n11762), .B(p_input[2607]), .Z(n11764) );
  XOR U11554 ( .A(n11766), .B(n11767), .Z(n11762) );
  AND U11555 ( .A(n11768), .B(n11769), .Z(n11767) );
  XNOR U11556 ( .A(p_input[2622]), .B(n11766), .Z(n11769) );
  XOR U11557 ( .A(n11766), .B(p_input[2606]), .Z(n11768) );
  XOR U11558 ( .A(n11770), .B(n11771), .Z(n11766) );
  AND U11559 ( .A(n11772), .B(n11773), .Z(n11771) );
  XNOR U11560 ( .A(p_input[2621]), .B(n11770), .Z(n11773) );
  XOR U11561 ( .A(n11770), .B(p_input[2605]), .Z(n11772) );
  XOR U11562 ( .A(n11774), .B(n11775), .Z(n11770) );
  AND U11563 ( .A(n11776), .B(n11777), .Z(n11775) );
  XNOR U11564 ( .A(p_input[2620]), .B(n11774), .Z(n11777) );
  XOR U11565 ( .A(n11774), .B(p_input[2604]), .Z(n11776) );
  XOR U11566 ( .A(n11778), .B(n11779), .Z(n11774) );
  AND U11567 ( .A(n11780), .B(n11781), .Z(n11779) );
  XNOR U11568 ( .A(p_input[2619]), .B(n11778), .Z(n11781) );
  XOR U11569 ( .A(n11778), .B(p_input[2603]), .Z(n11780) );
  XOR U11570 ( .A(n11782), .B(n11783), .Z(n11778) );
  AND U11571 ( .A(n11784), .B(n11785), .Z(n11783) );
  XNOR U11572 ( .A(p_input[2618]), .B(n11782), .Z(n11785) );
  XOR U11573 ( .A(n11782), .B(p_input[2602]), .Z(n11784) );
  XOR U11574 ( .A(n11786), .B(n11787), .Z(n11782) );
  AND U11575 ( .A(n11788), .B(n11789), .Z(n11787) );
  XNOR U11576 ( .A(p_input[2617]), .B(n11786), .Z(n11789) );
  XOR U11577 ( .A(n11786), .B(p_input[2601]), .Z(n11788) );
  XOR U11578 ( .A(n11790), .B(n11791), .Z(n11786) );
  AND U11579 ( .A(n11792), .B(n11793), .Z(n11791) );
  XNOR U11580 ( .A(p_input[2616]), .B(n11790), .Z(n11793) );
  XOR U11581 ( .A(n11790), .B(p_input[2600]), .Z(n11792) );
  XOR U11582 ( .A(n11794), .B(n11795), .Z(n11790) );
  AND U11583 ( .A(n11796), .B(n11797), .Z(n11795) );
  XNOR U11584 ( .A(p_input[2615]), .B(n11794), .Z(n11797) );
  XOR U11585 ( .A(n11794), .B(p_input[2599]), .Z(n11796) );
  XOR U11586 ( .A(n11798), .B(n11799), .Z(n11794) );
  AND U11587 ( .A(n11800), .B(n11801), .Z(n11799) );
  XNOR U11588 ( .A(p_input[2614]), .B(n11798), .Z(n11801) );
  XOR U11589 ( .A(n11798), .B(p_input[2598]), .Z(n11800) );
  XOR U11590 ( .A(n11802), .B(n11803), .Z(n11798) );
  AND U11591 ( .A(n11804), .B(n11805), .Z(n11803) );
  XNOR U11592 ( .A(p_input[2613]), .B(n11802), .Z(n11805) );
  XOR U11593 ( .A(n11802), .B(p_input[2597]), .Z(n11804) );
  XOR U11594 ( .A(n11806), .B(n11807), .Z(n11802) );
  AND U11595 ( .A(n11808), .B(n11809), .Z(n11807) );
  XNOR U11596 ( .A(p_input[2612]), .B(n11806), .Z(n11809) );
  XOR U11597 ( .A(n11806), .B(p_input[2596]), .Z(n11808) );
  XOR U11598 ( .A(n11810), .B(n11811), .Z(n11806) );
  AND U11599 ( .A(n11812), .B(n11813), .Z(n11811) );
  XNOR U11600 ( .A(p_input[2611]), .B(n11810), .Z(n11813) );
  XOR U11601 ( .A(n11810), .B(p_input[2595]), .Z(n11812) );
  XOR U11602 ( .A(n11814), .B(n11815), .Z(n11810) );
  AND U11603 ( .A(n11816), .B(n11817), .Z(n11815) );
  XNOR U11604 ( .A(p_input[2610]), .B(n11814), .Z(n11817) );
  XOR U11605 ( .A(n11814), .B(p_input[2594]), .Z(n11816) );
  XNOR U11606 ( .A(n11818), .B(n11819), .Z(n11814) );
  AND U11607 ( .A(n11820), .B(n11821), .Z(n11819) );
  XOR U11608 ( .A(p_input[2609]), .B(n11818), .Z(n11821) );
  XNOR U11609 ( .A(p_input[2593]), .B(n11818), .Z(n11820) );
  AND U11610 ( .A(p_input[2608]), .B(n11822), .Z(n11818) );
  IV U11611 ( .A(p_input[2592]), .Z(n11822) );
  XNOR U11612 ( .A(p_input[2560]), .B(n11823), .Z(n11625) );
  AND U11613 ( .A(n272), .B(n11824), .Z(n11823) );
  XOR U11614 ( .A(p_input[2576]), .B(p_input[2560]), .Z(n11824) );
  XOR U11615 ( .A(n11825), .B(n11826), .Z(n272) );
  AND U11616 ( .A(n11827), .B(n11828), .Z(n11826) );
  XNOR U11617 ( .A(p_input[2591]), .B(n11825), .Z(n11828) );
  XOR U11618 ( .A(n11825), .B(p_input[2575]), .Z(n11827) );
  XOR U11619 ( .A(n11829), .B(n11830), .Z(n11825) );
  AND U11620 ( .A(n11831), .B(n11832), .Z(n11830) );
  XNOR U11621 ( .A(p_input[2590]), .B(n11829), .Z(n11832) );
  XNOR U11622 ( .A(n11829), .B(n11639), .Z(n11831) );
  IV U11623 ( .A(p_input[2574]), .Z(n11639) );
  XOR U11624 ( .A(n11833), .B(n11834), .Z(n11829) );
  AND U11625 ( .A(n11835), .B(n11836), .Z(n11834) );
  XNOR U11626 ( .A(p_input[2589]), .B(n11833), .Z(n11836) );
  XNOR U11627 ( .A(n11833), .B(n11648), .Z(n11835) );
  IV U11628 ( .A(p_input[2573]), .Z(n11648) );
  XOR U11629 ( .A(n11837), .B(n11838), .Z(n11833) );
  AND U11630 ( .A(n11839), .B(n11840), .Z(n11838) );
  XNOR U11631 ( .A(p_input[2588]), .B(n11837), .Z(n11840) );
  XNOR U11632 ( .A(n11837), .B(n11657), .Z(n11839) );
  IV U11633 ( .A(p_input[2572]), .Z(n11657) );
  XOR U11634 ( .A(n11841), .B(n11842), .Z(n11837) );
  AND U11635 ( .A(n11843), .B(n11844), .Z(n11842) );
  XNOR U11636 ( .A(p_input[2587]), .B(n11841), .Z(n11844) );
  XNOR U11637 ( .A(n11841), .B(n11666), .Z(n11843) );
  IV U11638 ( .A(p_input[2571]), .Z(n11666) );
  XOR U11639 ( .A(n11845), .B(n11846), .Z(n11841) );
  AND U11640 ( .A(n11847), .B(n11848), .Z(n11846) );
  XNOR U11641 ( .A(p_input[2586]), .B(n11845), .Z(n11848) );
  XNOR U11642 ( .A(n11845), .B(n11675), .Z(n11847) );
  IV U11643 ( .A(p_input[2570]), .Z(n11675) );
  XOR U11644 ( .A(n11849), .B(n11850), .Z(n11845) );
  AND U11645 ( .A(n11851), .B(n11852), .Z(n11850) );
  XNOR U11646 ( .A(p_input[2585]), .B(n11849), .Z(n11852) );
  XNOR U11647 ( .A(n11849), .B(n11684), .Z(n11851) );
  IV U11648 ( .A(p_input[2569]), .Z(n11684) );
  XOR U11649 ( .A(n11853), .B(n11854), .Z(n11849) );
  AND U11650 ( .A(n11855), .B(n11856), .Z(n11854) );
  XNOR U11651 ( .A(p_input[2584]), .B(n11853), .Z(n11856) );
  XNOR U11652 ( .A(n11853), .B(n11693), .Z(n11855) );
  IV U11653 ( .A(p_input[2568]), .Z(n11693) );
  XOR U11654 ( .A(n11857), .B(n11858), .Z(n11853) );
  AND U11655 ( .A(n11859), .B(n11860), .Z(n11858) );
  XNOR U11656 ( .A(p_input[2583]), .B(n11857), .Z(n11860) );
  XNOR U11657 ( .A(n11857), .B(n11702), .Z(n11859) );
  IV U11658 ( .A(p_input[2567]), .Z(n11702) );
  XOR U11659 ( .A(n11861), .B(n11862), .Z(n11857) );
  AND U11660 ( .A(n11863), .B(n11864), .Z(n11862) );
  XNOR U11661 ( .A(p_input[2582]), .B(n11861), .Z(n11864) );
  XNOR U11662 ( .A(n11861), .B(n11711), .Z(n11863) );
  IV U11663 ( .A(p_input[2566]), .Z(n11711) );
  XOR U11664 ( .A(n11865), .B(n11866), .Z(n11861) );
  AND U11665 ( .A(n11867), .B(n11868), .Z(n11866) );
  XNOR U11666 ( .A(p_input[2581]), .B(n11865), .Z(n11868) );
  XNOR U11667 ( .A(n11865), .B(n11720), .Z(n11867) );
  IV U11668 ( .A(p_input[2565]), .Z(n11720) );
  XOR U11669 ( .A(n11869), .B(n11870), .Z(n11865) );
  AND U11670 ( .A(n11871), .B(n11872), .Z(n11870) );
  XNOR U11671 ( .A(p_input[2580]), .B(n11869), .Z(n11872) );
  XNOR U11672 ( .A(n11869), .B(n11729), .Z(n11871) );
  IV U11673 ( .A(p_input[2564]), .Z(n11729) );
  XOR U11674 ( .A(n11873), .B(n11874), .Z(n11869) );
  AND U11675 ( .A(n11875), .B(n11876), .Z(n11874) );
  XNOR U11676 ( .A(p_input[2579]), .B(n11873), .Z(n11876) );
  XNOR U11677 ( .A(n11873), .B(n11738), .Z(n11875) );
  IV U11678 ( .A(p_input[2563]), .Z(n11738) );
  XOR U11679 ( .A(n11877), .B(n11878), .Z(n11873) );
  AND U11680 ( .A(n11879), .B(n11880), .Z(n11878) );
  XNOR U11681 ( .A(p_input[2578]), .B(n11877), .Z(n11880) );
  XNOR U11682 ( .A(n11877), .B(n11747), .Z(n11879) );
  IV U11683 ( .A(p_input[2562]), .Z(n11747) );
  XNOR U11684 ( .A(n11881), .B(n11882), .Z(n11877) );
  AND U11685 ( .A(n11883), .B(n11884), .Z(n11882) );
  XOR U11686 ( .A(p_input[2577]), .B(n11881), .Z(n11884) );
  XNOR U11687 ( .A(p_input[2561]), .B(n11881), .Z(n11883) );
  AND U11688 ( .A(p_input[2576]), .B(n11885), .Z(n11881) );
  IV U11689 ( .A(p_input[2560]), .Z(n11885) );
  XOR U11690 ( .A(n11886), .B(n11887), .Z(n8340) );
  AND U11691 ( .A(n1008), .B(n11888), .Z(n11887) );
  XNOR U11692 ( .A(n11889), .B(n11886), .Z(n11888) );
  XOR U11693 ( .A(n11890), .B(n11891), .Z(n1008) );
  AND U11694 ( .A(n11892), .B(n11893), .Z(n11891) );
  XOR U11695 ( .A(n11890), .B(n8355), .Z(n11893) );
  XNOR U11696 ( .A(n11894), .B(n11895), .Z(n8355) );
  AND U11697 ( .A(n11896), .B(n935), .Z(n11895) );
  AND U11698 ( .A(n11894), .B(n11897), .Z(n11896) );
  XNOR U11699 ( .A(n8352), .B(n11890), .Z(n11892) );
  XOR U11700 ( .A(n11898), .B(n11899), .Z(n8352) );
  AND U11701 ( .A(n11900), .B(n932), .Z(n11899) );
  NOR U11702 ( .A(n11898), .B(n11901), .Z(n11900) );
  XOR U11703 ( .A(n11902), .B(n11903), .Z(n11890) );
  AND U11704 ( .A(n11904), .B(n11905), .Z(n11903) );
  XOR U11705 ( .A(n11902), .B(n8367), .Z(n11905) );
  XOR U11706 ( .A(n11906), .B(n11907), .Z(n8367) );
  AND U11707 ( .A(n935), .B(n11908), .Z(n11907) );
  XOR U11708 ( .A(n11909), .B(n11906), .Z(n11908) );
  XNOR U11709 ( .A(n8364), .B(n11902), .Z(n11904) );
  XOR U11710 ( .A(n11910), .B(n11911), .Z(n8364) );
  AND U11711 ( .A(n932), .B(n11912), .Z(n11911) );
  XOR U11712 ( .A(n11913), .B(n11910), .Z(n11912) );
  XOR U11713 ( .A(n11914), .B(n11915), .Z(n11902) );
  AND U11714 ( .A(n11916), .B(n11917), .Z(n11915) );
  XOR U11715 ( .A(n11914), .B(n8379), .Z(n11917) );
  XOR U11716 ( .A(n11918), .B(n11919), .Z(n8379) );
  AND U11717 ( .A(n935), .B(n11920), .Z(n11919) );
  XOR U11718 ( .A(n11921), .B(n11918), .Z(n11920) );
  XNOR U11719 ( .A(n8376), .B(n11914), .Z(n11916) );
  XOR U11720 ( .A(n11922), .B(n11923), .Z(n8376) );
  AND U11721 ( .A(n932), .B(n11924), .Z(n11923) );
  XOR U11722 ( .A(n11925), .B(n11922), .Z(n11924) );
  XOR U11723 ( .A(n11926), .B(n11927), .Z(n11914) );
  AND U11724 ( .A(n11928), .B(n11929), .Z(n11927) );
  XOR U11725 ( .A(n11926), .B(n8391), .Z(n11929) );
  XOR U11726 ( .A(n11930), .B(n11931), .Z(n8391) );
  AND U11727 ( .A(n935), .B(n11932), .Z(n11931) );
  XOR U11728 ( .A(n11933), .B(n11930), .Z(n11932) );
  XNOR U11729 ( .A(n8388), .B(n11926), .Z(n11928) );
  XOR U11730 ( .A(n11934), .B(n11935), .Z(n8388) );
  AND U11731 ( .A(n932), .B(n11936), .Z(n11935) );
  XOR U11732 ( .A(n11937), .B(n11934), .Z(n11936) );
  XOR U11733 ( .A(n11938), .B(n11939), .Z(n11926) );
  AND U11734 ( .A(n11940), .B(n11941), .Z(n11939) );
  XOR U11735 ( .A(n11938), .B(n8403), .Z(n11941) );
  XOR U11736 ( .A(n11942), .B(n11943), .Z(n8403) );
  AND U11737 ( .A(n935), .B(n11944), .Z(n11943) );
  XOR U11738 ( .A(n11945), .B(n11942), .Z(n11944) );
  XNOR U11739 ( .A(n8400), .B(n11938), .Z(n11940) );
  XOR U11740 ( .A(n11946), .B(n11947), .Z(n8400) );
  AND U11741 ( .A(n932), .B(n11948), .Z(n11947) );
  XOR U11742 ( .A(n11949), .B(n11946), .Z(n11948) );
  XOR U11743 ( .A(n11950), .B(n11951), .Z(n11938) );
  AND U11744 ( .A(n11952), .B(n11953), .Z(n11951) );
  XOR U11745 ( .A(n11950), .B(n8415), .Z(n11953) );
  XOR U11746 ( .A(n11954), .B(n11955), .Z(n8415) );
  AND U11747 ( .A(n935), .B(n11956), .Z(n11955) );
  XOR U11748 ( .A(n11957), .B(n11954), .Z(n11956) );
  XNOR U11749 ( .A(n8412), .B(n11950), .Z(n11952) );
  XOR U11750 ( .A(n11958), .B(n11959), .Z(n8412) );
  AND U11751 ( .A(n932), .B(n11960), .Z(n11959) );
  XOR U11752 ( .A(n11961), .B(n11958), .Z(n11960) );
  XOR U11753 ( .A(n11962), .B(n11963), .Z(n11950) );
  AND U11754 ( .A(n11964), .B(n11965), .Z(n11963) );
  XOR U11755 ( .A(n11962), .B(n8427), .Z(n11965) );
  XOR U11756 ( .A(n11966), .B(n11967), .Z(n8427) );
  AND U11757 ( .A(n935), .B(n11968), .Z(n11967) );
  XOR U11758 ( .A(n11969), .B(n11966), .Z(n11968) );
  XNOR U11759 ( .A(n8424), .B(n11962), .Z(n11964) );
  XOR U11760 ( .A(n11970), .B(n11971), .Z(n8424) );
  AND U11761 ( .A(n932), .B(n11972), .Z(n11971) );
  XOR U11762 ( .A(n11973), .B(n11970), .Z(n11972) );
  XOR U11763 ( .A(n11974), .B(n11975), .Z(n11962) );
  AND U11764 ( .A(n11976), .B(n11977), .Z(n11975) );
  XOR U11765 ( .A(n11974), .B(n8439), .Z(n11977) );
  XOR U11766 ( .A(n11978), .B(n11979), .Z(n8439) );
  AND U11767 ( .A(n935), .B(n11980), .Z(n11979) );
  XOR U11768 ( .A(n11981), .B(n11978), .Z(n11980) );
  XNOR U11769 ( .A(n8436), .B(n11974), .Z(n11976) );
  XOR U11770 ( .A(n11982), .B(n11983), .Z(n8436) );
  AND U11771 ( .A(n932), .B(n11984), .Z(n11983) );
  XOR U11772 ( .A(n11985), .B(n11982), .Z(n11984) );
  XOR U11773 ( .A(n11986), .B(n11987), .Z(n11974) );
  AND U11774 ( .A(n11988), .B(n11989), .Z(n11987) );
  XOR U11775 ( .A(n11986), .B(n8451), .Z(n11989) );
  XOR U11776 ( .A(n11990), .B(n11991), .Z(n8451) );
  AND U11777 ( .A(n935), .B(n11992), .Z(n11991) );
  XOR U11778 ( .A(n11993), .B(n11990), .Z(n11992) );
  XNOR U11779 ( .A(n8448), .B(n11986), .Z(n11988) );
  XOR U11780 ( .A(n11994), .B(n11995), .Z(n8448) );
  AND U11781 ( .A(n932), .B(n11996), .Z(n11995) );
  XOR U11782 ( .A(n11997), .B(n11994), .Z(n11996) );
  XOR U11783 ( .A(n11998), .B(n11999), .Z(n11986) );
  AND U11784 ( .A(n12000), .B(n12001), .Z(n11999) );
  XOR U11785 ( .A(n11998), .B(n8463), .Z(n12001) );
  XOR U11786 ( .A(n12002), .B(n12003), .Z(n8463) );
  AND U11787 ( .A(n935), .B(n12004), .Z(n12003) );
  XOR U11788 ( .A(n12005), .B(n12002), .Z(n12004) );
  XNOR U11789 ( .A(n8460), .B(n11998), .Z(n12000) );
  XOR U11790 ( .A(n12006), .B(n12007), .Z(n8460) );
  AND U11791 ( .A(n932), .B(n12008), .Z(n12007) );
  XOR U11792 ( .A(n12009), .B(n12006), .Z(n12008) );
  XOR U11793 ( .A(n12010), .B(n12011), .Z(n11998) );
  AND U11794 ( .A(n12012), .B(n12013), .Z(n12011) );
  XOR U11795 ( .A(n12010), .B(n8475), .Z(n12013) );
  XOR U11796 ( .A(n12014), .B(n12015), .Z(n8475) );
  AND U11797 ( .A(n935), .B(n12016), .Z(n12015) );
  XOR U11798 ( .A(n12017), .B(n12014), .Z(n12016) );
  XNOR U11799 ( .A(n8472), .B(n12010), .Z(n12012) );
  XOR U11800 ( .A(n12018), .B(n12019), .Z(n8472) );
  AND U11801 ( .A(n932), .B(n12020), .Z(n12019) );
  XOR U11802 ( .A(n12021), .B(n12018), .Z(n12020) );
  XOR U11803 ( .A(n12022), .B(n12023), .Z(n12010) );
  AND U11804 ( .A(n12024), .B(n12025), .Z(n12023) );
  XOR U11805 ( .A(n12022), .B(n8487), .Z(n12025) );
  XOR U11806 ( .A(n12026), .B(n12027), .Z(n8487) );
  AND U11807 ( .A(n935), .B(n12028), .Z(n12027) );
  XOR U11808 ( .A(n12029), .B(n12026), .Z(n12028) );
  XNOR U11809 ( .A(n8484), .B(n12022), .Z(n12024) );
  XOR U11810 ( .A(n12030), .B(n12031), .Z(n8484) );
  AND U11811 ( .A(n932), .B(n12032), .Z(n12031) );
  XOR U11812 ( .A(n12033), .B(n12030), .Z(n12032) );
  XOR U11813 ( .A(n12034), .B(n12035), .Z(n12022) );
  AND U11814 ( .A(n12036), .B(n12037), .Z(n12035) );
  XOR U11815 ( .A(n12034), .B(n8499), .Z(n12037) );
  XOR U11816 ( .A(n12038), .B(n12039), .Z(n8499) );
  AND U11817 ( .A(n935), .B(n12040), .Z(n12039) );
  XOR U11818 ( .A(n12041), .B(n12038), .Z(n12040) );
  XNOR U11819 ( .A(n8496), .B(n12034), .Z(n12036) );
  XOR U11820 ( .A(n12042), .B(n12043), .Z(n8496) );
  AND U11821 ( .A(n932), .B(n12044), .Z(n12043) );
  XOR U11822 ( .A(n12045), .B(n12042), .Z(n12044) );
  XOR U11823 ( .A(n12046), .B(n12047), .Z(n12034) );
  AND U11824 ( .A(n12048), .B(n12049), .Z(n12047) );
  XOR U11825 ( .A(n12046), .B(n8511), .Z(n12049) );
  XOR U11826 ( .A(n12050), .B(n12051), .Z(n8511) );
  AND U11827 ( .A(n935), .B(n12052), .Z(n12051) );
  XOR U11828 ( .A(n12053), .B(n12050), .Z(n12052) );
  XNOR U11829 ( .A(n8508), .B(n12046), .Z(n12048) );
  XOR U11830 ( .A(n12054), .B(n12055), .Z(n8508) );
  AND U11831 ( .A(n932), .B(n12056), .Z(n12055) );
  XOR U11832 ( .A(n12057), .B(n12054), .Z(n12056) );
  XOR U11833 ( .A(n12058), .B(n12059), .Z(n12046) );
  AND U11834 ( .A(n12060), .B(n12061), .Z(n12059) );
  XNOR U11835 ( .A(n12062), .B(n8524), .Z(n12061) );
  XOR U11836 ( .A(n12063), .B(n12064), .Z(n8524) );
  AND U11837 ( .A(n935), .B(n12065), .Z(n12064) );
  XOR U11838 ( .A(n12063), .B(n12066), .Z(n12065) );
  XNOR U11839 ( .A(n8521), .B(n12058), .Z(n12060) );
  XOR U11840 ( .A(n12067), .B(n12068), .Z(n8521) );
  AND U11841 ( .A(n932), .B(n12069), .Z(n12068) );
  XOR U11842 ( .A(n12067), .B(n12070), .Z(n12069) );
  IV U11843 ( .A(n12062), .Z(n12058) );
  AND U11844 ( .A(n11886), .B(n11889), .Z(n12062) );
  XNOR U11845 ( .A(n12071), .B(n12072), .Z(n11889) );
  AND U11846 ( .A(n935), .B(n12073), .Z(n12072) );
  XNOR U11847 ( .A(n12074), .B(n12071), .Z(n12073) );
  XOR U11848 ( .A(n12075), .B(n12076), .Z(n935) );
  AND U11849 ( .A(n12077), .B(n12078), .Z(n12076) );
  XOR U11850 ( .A(n11897), .B(n12075), .Z(n12078) );
  IV U11851 ( .A(n12079), .Z(n11897) );
  AND U11852 ( .A(n12080), .B(n12081), .Z(n12079) );
  XOR U11853 ( .A(n12075), .B(n11894), .Z(n12077) );
  AND U11854 ( .A(n12082), .B(n12083), .Z(n11894) );
  XOR U11855 ( .A(n12084), .B(n12085), .Z(n12075) );
  AND U11856 ( .A(n12086), .B(n12087), .Z(n12085) );
  XOR U11857 ( .A(n12084), .B(n11909), .Z(n12087) );
  XOR U11858 ( .A(n12088), .B(n12089), .Z(n11909) );
  AND U11859 ( .A(n775), .B(n12090), .Z(n12089) );
  XOR U11860 ( .A(n12091), .B(n12088), .Z(n12090) );
  XNOR U11861 ( .A(n11906), .B(n12084), .Z(n12086) );
  XOR U11862 ( .A(n12092), .B(n12093), .Z(n11906) );
  AND U11863 ( .A(n773), .B(n12094), .Z(n12093) );
  XOR U11864 ( .A(n12095), .B(n12092), .Z(n12094) );
  XOR U11865 ( .A(n12096), .B(n12097), .Z(n12084) );
  AND U11866 ( .A(n12098), .B(n12099), .Z(n12097) );
  XOR U11867 ( .A(n12096), .B(n11921), .Z(n12099) );
  XOR U11868 ( .A(n12100), .B(n12101), .Z(n11921) );
  AND U11869 ( .A(n775), .B(n12102), .Z(n12101) );
  XOR U11870 ( .A(n12103), .B(n12100), .Z(n12102) );
  XNOR U11871 ( .A(n11918), .B(n12096), .Z(n12098) );
  XOR U11872 ( .A(n12104), .B(n12105), .Z(n11918) );
  AND U11873 ( .A(n773), .B(n12106), .Z(n12105) );
  XOR U11874 ( .A(n12107), .B(n12104), .Z(n12106) );
  XOR U11875 ( .A(n12108), .B(n12109), .Z(n12096) );
  AND U11876 ( .A(n12110), .B(n12111), .Z(n12109) );
  XOR U11877 ( .A(n12108), .B(n11933), .Z(n12111) );
  XOR U11878 ( .A(n12112), .B(n12113), .Z(n11933) );
  AND U11879 ( .A(n775), .B(n12114), .Z(n12113) );
  XOR U11880 ( .A(n12115), .B(n12112), .Z(n12114) );
  XNOR U11881 ( .A(n11930), .B(n12108), .Z(n12110) );
  XOR U11882 ( .A(n12116), .B(n12117), .Z(n11930) );
  AND U11883 ( .A(n773), .B(n12118), .Z(n12117) );
  XOR U11884 ( .A(n12119), .B(n12116), .Z(n12118) );
  XOR U11885 ( .A(n12120), .B(n12121), .Z(n12108) );
  AND U11886 ( .A(n12122), .B(n12123), .Z(n12121) );
  XOR U11887 ( .A(n12120), .B(n11945), .Z(n12123) );
  XOR U11888 ( .A(n12124), .B(n12125), .Z(n11945) );
  AND U11889 ( .A(n775), .B(n12126), .Z(n12125) );
  XOR U11890 ( .A(n12127), .B(n12124), .Z(n12126) );
  XNOR U11891 ( .A(n11942), .B(n12120), .Z(n12122) );
  XOR U11892 ( .A(n12128), .B(n12129), .Z(n11942) );
  AND U11893 ( .A(n773), .B(n12130), .Z(n12129) );
  XOR U11894 ( .A(n12131), .B(n12128), .Z(n12130) );
  XOR U11895 ( .A(n12132), .B(n12133), .Z(n12120) );
  AND U11896 ( .A(n12134), .B(n12135), .Z(n12133) );
  XOR U11897 ( .A(n12132), .B(n11957), .Z(n12135) );
  XOR U11898 ( .A(n12136), .B(n12137), .Z(n11957) );
  AND U11899 ( .A(n775), .B(n12138), .Z(n12137) );
  XOR U11900 ( .A(n12139), .B(n12136), .Z(n12138) );
  XNOR U11901 ( .A(n11954), .B(n12132), .Z(n12134) );
  XOR U11902 ( .A(n12140), .B(n12141), .Z(n11954) );
  AND U11903 ( .A(n773), .B(n12142), .Z(n12141) );
  XOR U11904 ( .A(n12143), .B(n12140), .Z(n12142) );
  XOR U11905 ( .A(n12144), .B(n12145), .Z(n12132) );
  AND U11906 ( .A(n12146), .B(n12147), .Z(n12145) );
  XOR U11907 ( .A(n12144), .B(n11969), .Z(n12147) );
  XOR U11908 ( .A(n12148), .B(n12149), .Z(n11969) );
  AND U11909 ( .A(n775), .B(n12150), .Z(n12149) );
  XOR U11910 ( .A(n12151), .B(n12148), .Z(n12150) );
  XNOR U11911 ( .A(n11966), .B(n12144), .Z(n12146) );
  XOR U11912 ( .A(n12152), .B(n12153), .Z(n11966) );
  AND U11913 ( .A(n773), .B(n12154), .Z(n12153) );
  XOR U11914 ( .A(n12155), .B(n12152), .Z(n12154) );
  XOR U11915 ( .A(n12156), .B(n12157), .Z(n12144) );
  AND U11916 ( .A(n12158), .B(n12159), .Z(n12157) );
  XOR U11917 ( .A(n12156), .B(n11981), .Z(n12159) );
  XOR U11918 ( .A(n12160), .B(n12161), .Z(n11981) );
  AND U11919 ( .A(n775), .B(n12162), .Z(n12161) );
  XOR U11920 ( .A(n12163), .B(n12160), .Z(n12162) );
  XNOR U11921 ( .A(n11978), .B(n12156), .Z(n12158) );
  XOR U11922 ( .A(n12164), .B(n12165), .Z(n11978) );
  AND U11923 ( .A(n773), .B(n12166), .Z(n12165) );
  XOR U11924 ( .A(n12167), .B(n12164), .Z(n12166) );
  XOR U11925 ( .A(n12168), .B(n12169), .Z(n12156) );
  AND U11926 ( .A(n12170), .B(n12171), .Z(n12169) );
  XOR U11927 ( .A(n12168), .B(n11993), .Z(n12171) );
  XOR U11928 ( .A(n12172), .B(n12173), .Z(n11993) );
  AND U11929 ( .A(n775), .B(n12174), .Z(n12173) );
  XOR U11930 ( .A(n12175), .B(n12172), .Z(n12174) );
  XNOR U11931 ( .A(n11990), .B(n12168), .Z(n12170) );
  XOR U11932 ( .A(n12176), .B(n12177), .Z(n11990) );
  AND U11933 ( .A(n773), .B(n12178), .Z(n12177) );
  XOR U11934 ( .A(n12179), .B(n12176), .Z(n12178) );
  XOR U11935 ( .A(n12180), .B(n12181), .Z(n12168) );
  AND U11936 ( .A(n12182), .B(n12183), .Z(n12181) );
  XOR U11937 ( .A(n12180), .B(n12005), .Z(n12183) );
  XOR U11938 ( .A(n12184), .B(n12185), .Z(n12005) );
  AND U11939 ( .A(n775), .B(n12186), .Z(n12185) );
  XOR U11940 ( .A(n12187), .B(n12184), .Z(n12186) );
  XNOR U11941 ( .A(n12002), .B(n12180), .Z(n12182) );
  XOR U11942 ( .A(n12188), .B(n12189), .Z(n12002) );
  AND U11943 ( .A(n773), .B(n12190), .Z(n12189) );
  XOR U11944 ( .A(n12191), .B(n12188), .Z(n12190) );
  XOR U11945 ( .A(n12192), .B(n12193), .Z(n12180) );
  AND U11946 ( .A(n12194), .B(n12195), .Z(n12193) );
  XOR U11947 ( .A(n12192), .B(n12017), .Z(n12195) );
  XOR U11948 ( .A(n12196), .B(n12197), .Z(n12017) );
  AND U11949 ( .A(n775), .B(n12198), .Z(n12197) );
  XOR U11950 ( .A(n12199), .B(n12196), .Z(n12198) );
  XNOR U11951 ( .A(n12014), .B(n12192), .Z(n12194) );
  XOR U11952 ( .A(n12200), .B(n12201), .Z(n12014) );
  AND U11953 ( .A(n773), .B(n12202), .Z(n12201) );
  XOR U11954 ( .A(n12203), .B(n12200), .Z(n12202) );
  XOR U11955 ( .A(n12204), .B(n12205), .Z(n12192) );
  AND U11956 ( .A(n12206), .B(n12207), .Z(n12205) );
  XOR U11957 ( .A(n12204), .B(n12029), .Z(n12207) );
  XOR U11958 ( .A(n12208), .B(n12209), .Z(n12029) );
  AND U11959 ( .A(n775), .B(n12210), .Z(n12209) );
  XOR U11960 ( .A(n12211), .B(n12208), .Z(n12210) );
  XNOR U11961 ( .A(n12026), .B(n12204), .Z(n12206) );
  XOR U11962 ( .A(n12212), .B(n12213), .Z(n12026) );
  AND U11963 ( .A(n773), .B(n12214), .Z(n12213) );
  XOR U11964 ( .A(n12215), .B(n12212), .Z(n12214) );
  XOR U11965 ( .A(n12216), .B(n12217), .Z(n12204) );
  AND U11966 ( .A(n12218), .B(n12219), .Z(n12217) );
  XOR U11967 ( .A(n12216), .B(n12041), .Z(n12219) );
  XOR U11968 ( .A(n12220), .B(n12221), .Z(n12041) );
  AND U11969 ( .A(n775), .B(n12222), .Z(n12221) );
  XOR U11970 ( .A(n12223), .B(n12220), .Z(n12222) );
  XNOR U11971 ( .A(n12038), .B(n12216), .Z(n12218) );
  XOR U11972 ( .A(n12224), .B(n12225), .Z(n12038) );
  AND U11973 ( .A(n773), .B(n12226), .Z(n12225) );
  XOR U11974 ( .A(n12227), .B(n12224), .Z(n12226) );
  XOR U11975 ( .A(n12228), .B(n12229), .Z(n12216) );
  AND U11976 ( .A(n12230), .B(n12231), .Z(n12229) );
  XOR U11977 ( .A(n12228), .B(n12053), .Z(n12231) );
  XOR U11978 ( .A(n12232), .B(n12233), .Z(n12053) );
  AND U11979 ( .A(n775), .B(n12234), .Z(n12233) );
  XOR U11980 ( .A(n12235), .B(n12232), .Z(n12234) );
  XNOR U11981 ( .A(n12050), .B(n12228), .Z(n12230) );
  XOR U11982 ( .A(n12236), .B(n12237), .Z(n12050) );
  AND U11983 ( .A(n773), .B(n12238), .Z(n12237) );
  XOR U11984 ( .A(n12239), .B(n12236), .Z(n12238) );
  XOR U11985 ( .A(n12240), .B(n12241), .Z(n12228) );
  AND U11986 ( .A(n12242), .B(n12243), .Z(n12241) );
  XNOR U11987 ( .A(n12244), .B(n12066), .Z(n12243) );
  XOR U11988 ( .A(n12245), .B(n12246), .Z(n12066) );
  AND U11989 ( .A(n775), .B(n12247), .Z(n12246) );
  XOR U11990 ( .A(n12245), .B(n12248), .Z(n12247) );
  XNOR U11991 ( .A(n12063), .B(n12240), .Z(n12242) );
  XOR U11992 ( .A(n12249), .B(n12250), .Z(n12063) );
  AND U11993 ( .A(n773), .B(n12251), .Z(n12250) );
  XOR U11994 ( .A(n12249), .B(n12252), .Z(n12251) );
  IV U11995 ( .A(n12244), .Z(n12240) );
  AND U11996 ( .A(n12071), .B(n12074), .Z(n12244) );
  XNOR U11997 ( .A(n12253), .B(n12254), .Z(n12074) );
  AND U11998 ( .A(n775), .B(n12255), .Z(n12254) );
  XNOR U11999 ( .A(n12256), .B(n12253), .Z(n12255) );
  XOR U12000 ( .A(n12257), .B(n12258), .Z(n775) );
  AND U12001 ( .A(n12259), .B(n12260), .Z(n12258) );
  XNOR U12002 ( .A(n12080), .B(n12257), .Z(n12260) );
  AND U12003 ( .A(n12261), .B(n12262), .Z(n12080) );
  XOR U12004 ( .A(n12257), .B(n12081), .Z(n12259) );
  AND U12005 ( .A(n12263), .B(n12264), .Z(n12081) );
  XOR U12006 ( .A(n12265), .B(n12266), .Z(n12257) );
  AND U12007 ( .A(n12267), .B(n12268), .Z(n12266) );
  XOR U12008 ( .A(n12265), .B(n12091), .Z(n12268) );
  XOR U12009 ( .A(n12269), .B(n12270), .Z(n12091) );
  AND U12010 ( .A(n447), .B(n12271), .Z(n12270) );
  XOR U12011 ( .A(n12272), .B(n12269), .Z(n12271) );
  XNOR U12012 ( .A(n12088), .B(n12265), .Z(n12267) );
  XOR U12013 ( .A(n12273), .B(n12274), .Z(n12088) );
  AND U12014 ( .A(n445), .B(n12275), .Z(n12274) );
  XOR U12015 ( .A(n12276), .B(n12273), .Z(n12275) );
  XOR U12016 ( .A(n12277), .B(n12278), .Z(n12265) );
  AND U12017 ( .A(n12279), .B(n12280), .Z(n12278) );
  XOR U12018 ( .A(n12277), .B(n12103), .Z(n12280) );
  XOR U12019 ( .A(n12281), .B(n12282), .Z(n12103) );
  AND U12020 ( .A(n447), .B(n12283), .Z(n12282) );
  XOR U12021 ( .A(n12284), .B(n12281), .Z(n12283) );
  XNOR U12022 ( .A(n12100), .B(n12277), .Z(n12279) );
  XOR U12023 ( .A(n12285), .B(n12286), .Z(n12100) );
  AND U12024 ( .A(n445), .B(n12287), .Z(n12286) );
  XOR U12025 ( .A(n12288), .B(n12285), .Z(n12287) );
  XOR U12026 ( .A(n12289), .B(n12290), .Z(n12277) );
  AND U12027 ( .A(n12291), .B(n12292), .Z(n12290) );
  XOR U12028 ( .A(n12289), .B(n12115), .Z(n12292) );
  XOR U12029 ( .A(n12293), .B(n12294), .Z(n12115) );
  AND U12030 ( .A(n447), .B(n12295), .Z(n12294) );
  XOR U12031 ( .A(n12296), .B(n12293), .Z(n12295) );
  XNOR U12032 ( .A(n12112), .B(n12289), .Z(n12291) );
  XOR U12033 ( .A(n12297), .B(n12298), .Z(n12112) );
  AND U12034 ( .A(n445), .B(n12299), .Z(n12298) );
  XOR U12035 ( .A(n12300), .B(n12297), .Z(n12299) );
  XOR U12036 ( .A(n12301), .B(n12302), .Z(n12289) );
  AND U12037 ( .A(n12303), .B(n12304), .Z(n12302) );
  XOR U12038 ( .A(n12301), .B(n12127), .Z(n12304) );
  XOR U12039 ( .A(n12305), .B(n12306), .Z(n12127) );
  AND U12040 ( .A(n447), .B(n12307), .Z(n12306) );
  XOR U12041 ( .A(n12308), .B(n12305), .Z(n12307) );
  XNOR U12042 ( .A(n12124), .B(n12301), .Z(n12303) );
  XOR U12043 ( .A(n12309), .B(n12310), .Z(n12124) );
  AND U12044 ( .A(n445), .B(n12311), .Z(n12310) );
  XOR U12045 ( .A(n12312), .B(n12309), .Z(n12311) );
  XOR U12046 ( .A(n12313), .B(n12314), .Z(n12301) );
  AND U12047 ( .A(n12315), .B(n12316), .Z(n12314) );
  XOR U12048 ( .A(n12313), .B(n12139), .Z(n12316) );
  XOR U12049 ( .A(n12317), .B(n12318), .Z(n12139) );
  AND U12050 ( .A(n447), .B(n12319), .Z(n12318) );
  XOR U12051 ( .A(n12320), .B(n12317), .Z(n12319) );
  XNOR U12052 ( .A(n12136), .B(n12313), .Z(n12315) );
  XOR U12053 ( .A(n12321), .B(n12322), .Z(n12136) );
  AND U12054 ( .A(n445), .B(n12323), .Z(n12322) );
  XOR U12055 ( .A(n12324), .B(n12321), .Z(n12323) );
  XOR U12056 ( .A(n12325), .B(n12326), .Z(n12313) );
  AND U12057 ( .A(n12327), .B(n12328), .Z(n12326) );
  XOR U12058 ( .A(n12325), .B(n12151), .Z(n12328) );
  XOR U12059 ( .A(n12329), .B(n12330), .Z(n12151) );
  AND U12060 ( .A(n447), .B(n12331), .Z(n12330) );
  XOR U12061 ( .A(n12332), .B(n12329), .Z(n12331) );
  XNOR U12062 ( .A(n12148), .B(n12325), .Z(n12327) );
  XOR U12063 ( .A(n12333), .B(n12334), .Z(n12148) );
  AND U12064 ( .A(n445), .B(n12335), .Z(n12334) );
  XOR U12065 ( .A(n12336), .B(n12333), .Z(n12335) );
  XOR U12066 ( .A(n12337), .B(n12338), .Z(n12325) );
  AND U12067 ( .A(n12339), .B(n12340), .Z(n12338) );
  XOR U12068 ( .A(n12337), .B(n12163), .Z(n12340) );
  XOR U12069 ( .A(n12341), .B(n12342), .Z(n12163) );
  AND U12070 ( .A(n447), .B(n12343), .Z(n12342) );
  XOR U12071 ( .A(n12344), .B(n12341), .Z(n12343) );
  XNOR U12072 ( .A(n12160), .B(n12337), .Z(n12339) );
  XOR U12073 ( .A(n12345), .B(n12346), .Z(n12160) );
  AND U12074 ( .A(n445), .B(n12347), .Z(n12346) );
  XOR U12075 ( .A(n12348), .B(n12345), .Z(n12347) );
  XOR U12076 ( .A(n12349), .B(n12350), .Z(n12337) );
  AND U12077 ( .A(n12351), .B(n12352), .Z(n12350) );
  XOR U12078 ( .A(n12349), .B(n12175), .Z(n12352) );
  XOR U12079 ( .A(n12353), .B(n12354), .Z(n12175) );
  AND U12080 ( .A(n447), .B(n12355), .Z(n12354) );
  XOR U12081 ( .A(n12356), .B(n12353), .Z(n12355) );
  XNOR U12082 ( .A(n12172), .B(n12349), .Z(n12351) );
  XOR U12083 ( .A(n12357), .B(n12358), .Z(n12172) );
  AND U12084 ( .A(n445), .B(n12359), .Z(n12358) );
  XOR U12085 ( .A(n12360), .B(n12357), .Z(n12359) );
  XOR U12086 ( .A(n12361), .B(n12362), .Z(n12349) );
  AND U12087 ( .A(n12363), .B(n12364), .Z(n12362) );
  XOR U12088 ( .A(n12361), .B(n12187), .Z(n12364) );
  XOR U12089 ( .A(n12365), .B(n12366), .Z(n12187) );
  AND U12090 ( .A(n447), .B(n12367), .Z(n12366) );
  XOR U12091 ( .A(n12368), .B(n12365), .Z(n12367) );
  XNOR U12092 ( .A(n12184), .B(n12361), .Z(n12363) );
  XOR U12093 ( .A(n12369), .B(n12370), .Z(n12184) );
  AND U12094 ( .A(n445), .B(n12371), .Z(n12370) );
  XOR U12095 ( .A(n12372), .B(n12369), .Z(n12371) );
  XOR U12096 ( .A(n12373), .B(n12374), .Z(n12361) );
  AND U12097 ( .A(n12375), .B(n12376), .Z(n12374) );
  XOR U12098 ( .A(n12373), .B(n12199), .Z(n12376) );
  XOR U12099 ( .A(n12377), .B(n12378), .Z(n12199) );
  AND U12100 ( .A(n447), .B(n12379), .Z(n12378) );
  XOR U12101 ( .A(n12380), .B(n12377), .Z(n12379) );
  XNOR U12102 ( .A(n12196), .B(n12373), .Z(n12375) );
  XOR U12103 ( .A(n12381), .B(n12382), .Z(n12196) );
  AND U12104 ( .A(n445), .B(n12383), .Z(n12382) );
  XOR U12105 ( .A(n12384), .B(n12381), .Z(n12383) );
  XOR U12106 ( .A(n12385), .B(n12386), .Z(n12373) );
  AND U12107 ( .A(n12387), .B(n12388), .Z(n12386) );
  XOR U12108 ( .A(n12385), .B(n12211), .Z(n12388) );
  XOR U12109 ( .A(n12389), .B(n12390), .Z(n12211) );
  AND U12110 ( .A(n447), .B(n12391), .Z(n12390) );
  XOR U12111 ( .A(n12392), .B(n12389), .Z(n12391) );
  XNOR U12112 ( .A(n12208), .B(n12385), .Z(n12387) );
  XOR U12113 ( .A(n12393), .B(n12394), .Z(n12208) );
  AND U12114 ( .A(n445), .B(n12395), .Z(n12394) );
  XOR U12115 ( .A(n12396), .B(n12393), .Z(n12395) );
  XOR U12116 ( .A(n12397), .B(n12398), .Z(n12385) );
  AND U12117 ( .A(n12399), .B(n12400), .Z(n12398) );
  XOR U12118 ( .A(n12397), .B(n12223), .Z(n12400) );
  XOR U12119 ( .A(n12401), .B(n12402), .Z(n12223) );
  AND U12120 ( .A(n447), .B(n12403), .Z(n12402) );
  XOR U12121 ( .A(n12404), .B(n12401), .Z(n12403) );
  XNOR U12122 ( .A(n12220), .B(n12397), .Z(n12399) );
  XOR U12123 ( .A(n12405), .B(n12406), .Z(n12220) );
  AND U12124 ( .A(n445), .B(n12407), .Z(n12406) );
  XOR U12125 ( .A(n12408), .B(n12405), .Z(n12407) );
  XOR U12126 ( .A(n12409), .B(n12410), .Z(n12397) );
  AND U12127 ( .A(n12411), .B(n12412), .Z(n12410) );
  XOR U12128 ( .A(n12409), .B(n12235), .Z(n12412) );
  XOR U12129 ( .A(n12413), .B(n12414), .Z(n12235) );
  AND U12130 ( .A(n447), .B(n12415), .Z(n12414) );
  XOR U12131 ( .A(n12416), .B(n12413), .Z(n12415) );
  XNOR U12132 ( .A(n12232), .B(n12409), .Z(n12411) );
  XOR U12133 ( .A(n12417), .B(n12418), .Z(n12232) );
  AND U12134 ( .A(n445), .B(n12419), .Z(n12418) );
  XOR U12135 ( .A(n12420), .B(n12417), .Z(n12419) );
  XOR U12136 ( .A(n12421), .B(n12422), .Z(n12409) );
  AND U12137 ( .A(n12423), .B(n12424), .Z(n12422) );
  XNOR U12138 ( .A(n12425), .B(n12248), .Z(n12424) );
  XOR U12139 ( .A(n12426), .B(n12427), .Z(n12248) );
  AND U12140 ( .A(n447), .B(n12428), .Z(n12427) );
  XOR U12141 ( .A(n12426), .B(n12429), .Z(n12428) );
  XNOR U12142 ( .A(n12245), .B(n12421), .Z(n12423) );
  XOR U12143 ( .A(n12430), .B(n12431), .Z(n12245) );
  AND U12144 ( .A(n445), .B(n12432), .Z(n12431) );
  XOR U12145 ( .A(n12430), .B(n12433), .Z(n12432) );
  IV U12146 ( .A(n12425), .Z(n12421) );
  AND U12147 ( .A(n12253), .B(n12256), .Z(n12425) );
  XNOR U12148 ( .A(n12434), .B(n12435), .Z(n12256) );
  AND U12149 ( .A(n447), .B(n12436), .Z(n12435) );
  XNOR U12150 ( .A(n12437), .B(n12434), .Z(n12436) );
  XOR U12151 ( .A(n12438), .B(n12439), .Z(n447) );
  AND U12152 ( .A(n12440), .B(n12441), .Z(n12439) );
  XNOR U12153 ( .A(n12261), .B(n12438), .Z(n12441) );
  AND U12154 ( .A(p_input[2559]), .B(p_input[2543]), .Z(n12261) );
  XOR U12155 ( .A(n12438), .B(n12262), .Z(n12440) );
  AND U12156 ( .A(p_input[2527]), .B(p_input[2511]), .Z(n12262) );
  XOR U12157 ( .A(n12442), .B(n12443), .Z(n12438) );
  AND U12158 ( .A(n12444), .B(n12445), .Z(n12443) );
  XOR U12159 ( .A(n12442), .B(n12272), .Z(n12445) );
  XNOR U12160 ( .A(p_input[2542]), .B(n12446), .Z(n12272) );
  AND U12161 ( .A(n291), .B(n12447), .Z(n12446) );
  XOR U12162 ( .A(p_input[2558]), .B(p_input[2542]), .Z(n12447) );
  XNOR U12163 ( .A(n12269), .B(n12442), .Z(n12444) );
  XOR U12164 ( .A(n12448), .B(n12449), .Z(n12269) );
  AND U12165 ( .A(n289), .B(n12450), .Z(n12449) );
  XOR U12166 ( .A(p_input[2526]), .B(p_input[2510]), .Z(n12450) );
  XOR U12167 ( .A(n12451), .B(n12452), .Z(n12442) );
  AND U12168 ( .A(n12453), .B(n12454), .Z(n12452) );
  XOR U12169 ( .A(n12451), .B(n12284), .Z(n12454) );
  XNOR U12170 ( .A(p_input[2541]), .B(n12455), .Z(n12284) );
  AND U12171 ( .A(n291), .B(n12456), .Z(n12455) );
  XOR U12172 ( .A(p_input[2557]), .B(p_input[2541]), .Z(n12456) );
  XNOR U12173 ( .A(n12281), .B(n12451), .Z(n12453) );
  XOR U12174 ( .A(n12457), .B(n12458), .Z(n12281) );
  AND U12175 ( .A(n289), .B(n12459), .Z(n12458) );
  XOR U12176 ( .A(p_input[2525]), .B(p_input[2509]), .Z(n12459) );
  XOR U12177 ( .A(n12460), .B(n12461), .Z(n12451) );
  AND U12178 ( .A(n12462), .B(n12463), .Z(n12461) );
  XOR U12179 ( .A(n12460), .B(n12296), .Z(n12463) );
  XNOR U12180 ( .A(p_input[2540]), .B(n12464), .Z(n12296) );
  AND U12181 ( .A(n291), .B(n12465), .Z(n12464) );
  XOR U12182 ( .A(p_input[2556]), .B(p_input[2540]), .Z(n12465) );
  XNOR U12183 ( .A(n12293), .B(n12460), .Z(n12462) );
  XOR U12184 ( .A(n12466), .B(n12467), .Z(n12293) );
  AND U12185 ( .A(n289), .B(n12468), .Z(n12467) );
  XOR U12186 ( .A(p_input[2524]), .B(p_input[2508]), .Z(n12468) );
  XOR U12187 ( .A(n12469), .B(n12470), .Z(n12460) );
  AND U12188 ( .A(n12471), .B(n12472), .Z(n12470) );
  XOR U12189 ( .A(n12469), .B(n12308), .Z(n12472) );
  XNOR U12190 ( .A(p_input[2539]), .B(n12473), .Z(n12308) );
  AND U12191 ( .A(n291), .B(n12474), .Z(n12473) );
  XOR U12192 ( .A(p_input[2555]), .B(p_input[2539]), .Z(n12474) );
  XNOR U12193 ( .A(n12305), .B(n12469), .Z(n12471) );
  XOR U12194 ( .A(n12475), .B(n12476), .Z(n12305) );
  AND U12195 ( .A(n289), .B(n12477), .Z(n12476) );
  XOR U12196 ( .A(p_input[2523]), .B(p_input[2507]), .Z(n12477) );
  XOR U12197 ( .A(n12478), .B(n12479), .Z(n12469) );
  AND U12198 ( .A(n12480), .B(n12481), .Z(n12479) );
  XOR U12199 ( .A(n12478), .B(n12320), .Z(n12481) );
  XNOR U12200 ( .A(p_input[2538]), .B(n12482), .Z(n12320) );
  AND U12201 ( .A(n291), .B(n12483), .Z(n12482) );
  XOR U12202 ( .A(p_input[2554]), .B(p_input[2538]), .Z(n12483) );
  XNOR U12203 ( .A(n12317), .B(n12478), .Z(n12480) );
  XOR U12204 ( .A(n12484), .B(n12485), .Z(n12317) );
  AND U12205 ( .A(n289), .B(n12486), .Z(n12485) );
  XOR U12206 ( .A(p_input[2522]), .B(p_input[2506]), .Z(n12486) );
  XOR U12207 ( .A(n12487), .B(n12488), .Z(n12478) );
  AND U12208 ( .A(n12489), .B(n12490), .Z(n12488) );
  XOR U12209 ( .A(n12487), .B(n12332), .Z(n12490) );
  XNOR U12210 ( .A(p_input[2537]), .B(n12491), .Z(n12332) );
  AND U12211 ( .A(n291), .B(n12492), .Z(n12491) );
  XOR U12212 ( .A(p_input[2553]), .B(p_input[2537]), .Z(n12492) );
  XNOR U12213 ( .A(n12329), .B(n12487), .Z(n12489) );
  XOR U12214 ( .A(n12493), .B(n12494), .Z(n12329) );
  AND U12215 ( .A(n289), .B(n12495), .Z(n12494) );
  XOR U12216 ( .A(p_input[2521]), .B(p_input[2505]), .Z(n12495) );
  XOR U12217 ( .A(n12496), .B(n12497), .Z(n12487) );
  AND U12218 ( .A(n12498), .B(n12499), .Z(n12497) );
  XOR U12219 ( .A(n12496), .B(n12344), .Z(n12499) );
  XNOR U12220 ( .A(p_input[2536]), .B(n12500), .Z(n12344) );
  AND U12221 ( .A(n291), .B(n12501), .Z(n12500) );
  XOR U12222 ( .A(p_input[2552]), .B(p_input[2536]), .Z(n12501) );
  XNOR U12223 ( .A(n12341), .B(n12496), .Z(n12498) );
  XOR U12224 ( .A(n12502), .B(n12503), .Z(n12341) );
  AND U12225 ( .A(n289), .B(n12504), .Z(n12503) );
  XOR U12226 ( .A(p_input[2520]), .B(p_input[2504]), .Z(n12504) );
  XOR U12227 ( .A(n12505), .B(n12506), .Z(n12496) );
  AND U12228 ( .A(n12507), .B(n12508), .Z(n12506) );
  XOR U12229 ( .A(n12505), .B(n12356), .Z(n12508) );
  XNOR U12230 ( .A(p_input[2535]), .B(n12509), .Z(n12356) );
  AND U12231 ( .A(n291), .B(n12510), .Z(n12509) );
  XOR U12232 ( .A(p_input[2551]), .B(p_input[2535]), .Z(n12510) );
  XNOR U12233 ( .A(n12353), .B(n12505), .Z(n12507) );
  XOR U12234 ( .A(n12511), .B(n12512), .Z(n12353) );
  AND U12235 ( .A(n289), .B(n12513), .Z(n12512) );
  XOR U12236 ( .A(p_input[2519]), .B(p_input[2503]), .Z(n12513) );
  XOR U12237 ( .A(n12514), .B(n12515), .Z(n12505) );
  AND U12238 ( .A(n12516), .B(n12517), .Z(n12515) );
  XOR U12239 ( .A(n12514), .B(n12368), .Z(n12517) );
  XNOR U12240 ( .A(p_input[2534]), .B(n12518), .Z(n12368) );
  AND U12241 ( .A(n291), .B(n12519), .Z(n12518) );
  XOR U12242 ( .A(p_input[2550]), .B(p_input[2534]), .Z(n12519) );
  XNOR U12243 ( .A(n12365), .B(n12514), .Z(n12516) );
  XOR U12244 ( .A(n12520), .B(n12521), .Z(n12365) );
  AND U12245 ( .A(n289), .B(n12522), .Z(n12521) );
  XOR U12246 ( .A(p_input[2518]), .B(p_input[2502]), .Z(n12522) );
  XOR U12247 ( .A(n12523), .B(n12524), .Z(n12514) );
  AND U12248 ( .A(n12525), .B(n12526), .Z(n12524) );
  XOR U12249 ( .A(n12523), .B(n12380), .Z(n12526) );
  XNOR U12250 ( .A(p_input[2533]), .B(n12527), .Z(n12380) );
  AND U12251 ( .A(n291), .B(n12528), .Z(n12527) );
  XOR U12252 ( .A(p_input[2549]), .B(p_input[2533]), .Z(n12528) );
  XNOR U12253 ( .A(n12377), .B(n12523), .Z(n12525) );
  XOR U12254 ( .A(n12529), .B(n12530), .Z(n12377) );
  AND U12255 ( .A(n289), .B(n12531), .Z(n12530) );
  XOR U12256 ( .A(p_input[2517]), .B(p_input[2501]), .Z(n12531) );
  XOR U12257 ( .A(n12532), .B(n12533), .Z(n12523) );
  AND U12258 ( .A(n12534), .B(n12535), .Z(n12533) );
  XOR U12259 ( .A(n12532), .B(n12392), .Z(n12535) );
  XNOR U12260 ( .A(p_input[2532]), .B(n12536), .Z(n12392) );
  AND U12261 ( .A(n291), .B(n12537), .Z(n12536) );
  XOR U12262 ( .A(p_input[2548]), .B(p_input[2532]), .Z(n12537) );
  XNOR U12263 ( .A(n12389), .B(n12532), .Z(n12534) );
  XOR U12264 ( .A(n12538), .B(n12539), .Z(n12389) );
  AND U12265 ( .A(n289), .B(n12540), .Z(n12539) );
  XOR U12266 ( .A(p_input[2516]), .B(p_input[2500]), .Z(n12540) );
  XOR U12267 ( .A(n12541), .B(n12542), .Z(n12532) );
  AND U12268 ( .A(n12543), .B(n12544), .Z(n12542) );
  XOR U12269 ( .A(n12541), .B(n12404), .Z(n12544) );
  XNOR U12270 ( .A(p_input[2531]), .B(n12545), .Z(n12404) );
  AND U12271 ( .A(n291), .B(n12546), .Z(n12545) );
  XOR U12272 ( .A(p_input[2547]), .B(p_input[2531]), .Z(n12546) );
  XNOR U12273 ( .A(n12401), .B(n12541), .Z(n12543) );
  XOR U12274 ( .A(n12547), .B(n12548), .Z(n12401) );
  AND U12275 ( .A(n289), .B(n12549), .Z(n12548) );
  XOR U12276 ( .A(p_input[2515]), .B(p_input[2499]), .Z(n12549) );
  XOR U12277 ( .A(n12550), .B(n12551), .Z(n12541) );
  AND U12278 ( .A(n12552), .B(n12553), .Z(n12551) );
  XOR U12279 ( .A(n12550), .B(n12416), .Z(n12553) );
  XNOR U12280 ( .A(p_input[2530]), .B(n12554), .Z(n12416) );
  AND U12281 ( .A(n291), .B(n12555), .Z(n12554) );
  XOR U12282 ( .A(p_input[2546]), .B(p_input[2530]), .Z(n12555) );
  XNOR U12283 ( .A(n12413), .B(n12550), .Z(n12552) );
  XOR U12284 ( .A(n12556), .B(n12557), .Z(n12413) );
  AND U12285 ( .A(n289), .B(n12558), .Z(n12557) );
  XOR U12286 ( .A(p_input[2514]), .B(p_input[2498]), .Z(n12558) );
  XOR U12287 ( .A(n12559), .B(n12560), .Z(n12550) );
  AND U12288 ( .A(n12561), .B(n12562), .Z(n12560) );
  XNOR U12289 ( .A(n12563), .B(n12429), .Z(n12562) );
  XNOR U12290 ( .A(p_input[2529]), .B(n12564), .Z(n12429) );
  AND U12291 ( .A(n291), .B(n12565), .Z(n12564) );
  XNOR U12292 ( .A(p_input[2545]), .B(n12566), .Z(n12565) );
  IV U12293 ( .A(p_input[2529]), .Z(n12566) );
  XNOR U12294 ( .A(n12426), .B(n12559), .Z(n12561) );
  XNOR U12295 ( .A(p_input[2497]), .B(n12567), .Z(n12426) );
  AND U12296 ( .A(n289), .B(n12568), .Z(n12567) );
  XOR U12297 ( .A(p_input[2513]), .B(p_input[2497]), .Z(n12568) );
  IV U12298 ( .A(n12563), .Z(n12559) );
  AND U12299 ( .A(n12434), .B(n12437), .Z(n12563) );
  XOR U12300 ( .A(p_input[2528]), .B(n12569), .Z(n12437) );
  AND U12301 ( .A(n291), .B(n12570), .Z(n12569) );
  XOR U12302 ( .A(p_input[2544]), .B(p_input[2528]), .Z(n12570) );
  XOR U12303 ( .A(n12571), .B(n12572), .Z(n291) );
  AND U12304 ( .A(n12573), .B(n12574), .Z(n12572) );
  XNOR U12305 ( .A(p_input[2559]), .B(n12571), .Z(n12574) );
  XOR U12306 ( .A(n12571), .B(p_input[2543]), .Z(n12573) );
  XOR U12307 ( .A(n12575), .B(n12576), .Z(n12571) );
  AND U12308 ( .A(n12577), .B(n12578), .Z(n12576) );
  XNOR U12309 ( .A(p_input[2558]), .B(n12575), .Z(n12578) );
  XOR U12310 ( .A(n12575), .B(p_input[2542]), .Z(n12577) );
  XOR U12311 ( .A(n12579), .B(n12580), .Z(n12575) );
  AND U12312 ( .A(n12581), .B(n12582), .Z(n12580) );
  XNOR U12313 ( .A(p_input[2557]), .B(n12579), .Z(n12582) );
  XOR U12314 ( .A(n12579), .B(p_input[2541]), .Z(n12581) );
  XOR U12315 ( .A(n12583), .B(n12584), .Z(n12579) );
  AND U12316 ( .A(n12585), .B(n12586), .Z(n12584) );
  XNOR U12317 ( .A(p_input[2556]), .B(n12583), .Z(n12586) );
  XOR U12318 ( .A(n12583), .B(p_input[2540]), .Z(n12585) );
  XOR U12319 ( .A(n12587), .B(n12588), .Z(n12583) );
  AND U12320 ( .A(n12589), .B(n12590), .Z(n12588) );
  XNOR U12321 ( .A(p_input[2555]), .B(n12587), .Z(n12590) );
  XOR U12322 ( .A(n12587), .B(p_input[2539]), .Z(n12589) );
  XOR U12323 ( .A(n12591), .B(n12592), .Z(n12587) );
  AND U12324 ( .A(n12593), .B(n12594), .Z(n12592) );
  XNOR U12325 ( .A(p_input[2554]), .B(n12591), .Z(n12594) );
  XOR U12326 ( .A(n12591), .B(p_input[2538]), .Z(n12593) );
  XOR U12327 ( .A(n12595), .B(n12596), .Z(n12591) );
  AND U12328 ( .A(n12597), .B(n12598), .Z(n12596) );
  XNOR U12329 ( .A(p_input[2553]), .B(n12595), .Z(n12598) );
  XOR U12330 ( .A(n12595), .B(p_input[2537]), .Z(n12597) );
  XOR U12331 ( .A(n12599), .B(n12600), .Z(n12595) );
  AND U12332 ( .A(n12601), .B(n12602), .Z(n12600) );
  XNOR U12333 ( .A(p_input[2552]), .B(n12599), .Z(n12602) );
  XOR U12334 ( .A(n12599), .B(p_input[2536]), .Z(n12601) );
  XOR U12335 ( .A(n12603), .B(n12604), .Z(n12599) );
  AND U12336 ( .A(n12605), .B(n12606), .Z(n12604) );
  XNOR U12337 ( .A(p_input[2551]), .B(n12603), .Z(n12606) );
  XOR U12338 ( .A(n12603), .B(p_input[2535]), .Z(n12605) );
  XOR U12339 ( .A(n12607), .B(n12608), .Z(n12603) );
  AND U12340 ( .A(n12609), .B(n12610), .Z(n12608) );
  XNOR U12341 ( .A(p_input[2550]), .B(n12607), .Z(n12610) );
  XOR U12342 ( .A(n12607), .B(p_input[2534]), .Z(n12609) );
  XOR U12343 ( .A(n12611), .B(n12612), .Z(n12607) );
  AND U12344 ( .A(n12613), .B(n12614), .Z(n12612) );
  XNOR U12345 ( .A(p_input[2549]), .B(n12611), .Z(n12614) );
  XOR U12346 ( .A(n12611), .B(p_input[2533]), .Z(n12613) );
  XOR U12347 ( .A(n12615), .B(n12616), .Z(n12611) );
  AND U12348 ( .A(n12617), .B(n12618), .Z(n12616) );
  XNOR U12349 ( .A(p_input[2548]), .B(n12615), .Z(n12618) );
  XOR U12350 ( .A(n12615), .B(p_input[2532]), .Z(n12617) );
  XOR U12351 ( .A(n12619), .B(n12620), .Z(n12615) );
  AND U12352 ( .A(n12621), .B(n12622), .Z(n12620) );
  XNOR U12353 ( .A(p_input[2547]), .B(n12619), .Z(n12622) );
  XOR U12354 ( .A(n12619), .B(p_input[2531]), .Z(n12621) );
  XOR U12355 ( .A(n12623), .B(n12624), .Z(n12619) );
  AND U12356 ( .A(n12625), .B(n12626), .Z(n12624) );
  XNOR U12357 ( .A(p_input[2546]), .B(n12623), .Z(n12626) );
  XOR U12358 ( .A(n12623), .B(p_input[2530]), .Z(n12625) );
  XNOR U12359 ( .A(n12627), .B(n12628), .Z(n12623) );
  AND U12360 ( .A(n12629), .B(n12630), .Z(n12628) );
  XOR U12361 ( .A(p_input[2545]), .B(n12627), .Z(n12630) );
  XNOR U12362 ( .A(p_input[2529]), .B(n12627), .Z(n12629) );
  AND U12363 ( .A(p_input[2544]), .B(n12631), .Z(n12627) );
  IV U12364 ( .A(p_input[2528]), .Z(n12631) );
  XNOR U12365 ( .A(p_input[2496]), .B(n12632), .Z(n12434) );
  AND U12366 ( .A(n289), .B(n12633), .Z(n12632) );
  XOR U12367 ( .A(p_input[2512]), .B(p_input[2496]), .Z(n12633) );
  XOR U12368 ( .A(n12634), .B(n12635), .Z(n289) );
  AND U12369 ( .A(n12636), .B(n12637), .Z(n12635) );
  XNOR U12370 ( .A(p_input[2527]), .B(n12634), .Z(n12637) );
  XOR U12371 ( .A(n12634), .B(p_input[2511]), .Z(n12636) );
  XOR U12372 ( .A(n12638), .B(n12639), .Z(n12634) );
  AND U12373 ( .A(n12640), .B(n12641), .Z(n12639) );
  XNOR U12374 ( .A(p_input[2526]), .B(n12638), .Z(n12641) );
  XNOR U12375 ( .A(n12638), .B(n12448), .Z(n12640) );
  IV U12376 ( .A(p_input[2510]), .Z(n12448) );
  XOR U12377 ( .A(n12642), .B(n12643), .Z(n12638) );
  AND U12378 ( .A(n12644), .B(n12645), .Z(n12643) );
  XNOR U12379 ( .A(p_input[2525]), .B(n12642), .Z(n12645) );
  XNOR U12380 ( .A(n12642), .B(n12457), .Z(n12644) );
  IV U12381 ( .A(p_input[2509]), .Z(n12457) );
  XOR U12382 ( .A(n12646), .B(n12647), .Z(n12642) );
  AND U12383 ( .A(n12648), .B(n12649), .Z(n12647) );
  XNOR U12384 ( .A(p_input[2524]), .B(n12646), .Z(n12649) );
  XNOR U12385 ( .A(n12646), .B(n12466), .Z(n12648) );
  IV U12386 ( .A(p_input[2508]), .Z(n12466) );
  XOR U12387 ( .A(n12650), .B(n12651), .Z(n12646) );
  AND U12388 ( .A(n12652), .B(n12653), .Z(n12651) );
  XNOR U12389 ( .A(p_input[2523]), .B(n12650), .Z(n12653) );
  XNOR U12390 ( .A(n12650), .B(n12475), .Z(n12652) );
  IV U12391 ( .A(p_input[2507]), .Z(n12475) );
  XOR U12392 ( .A(n12654), .B(n12655), .Z(n12650) );
  AND U12393 ( .A(n12656), .B(n12657), .Z(n12655) );
  XNOR U12394 ( .A(p_input[2522]), .B(n12654), .Z(n12657) );
  XNOR U12395 ( .A(n12654), .B(n12484), .Z(n12656) );
  IV U12396 ( .A(p_input[2506]), .Z(n12484) );
  XOR U12397 ( .A(n12658), .B(n12659), .Z(n12654) );
  AND U12398 ( .A(n12660), .B(n12661), .Z(n12659) );
  XNOR U12399 ( .A(p_input[2521]), .B(n12658), .Z(n12661) );
  XNOR U12400 ( .A(n12658), .B(n12493), .Z(n12660) );
  IV U12401 ( .A(p_input[2505]), .Z(n12493) );
  XOR U12402 ( .A(n12662), .B(n12663), .Z(n12658) );
  AND U12403 ( .A(n12664), .B(n12665), .Z(n12663) );
  XNOR U12404 ( .A(p_input[2520]), .B(n12662), .Z(n12665) );
  XNOR U12405 ( .A(n12662), .B(n12502), .Z(n12664) );
  IV U12406 ( .A(p_input[2504]), .Z(n12502) );
  XOR U12407 ( .A(n12666), .B(n12667), .Z(n12662) );
  AND U12408 ( .A(n12668), .B(n12669), .Z(n12667) );
  XNOR U12409 ( .A(p_input[2519]), .B(n12666), .Z(n12669) );
  XNOR U12410 ( .A(n12666), .B(n12511), .Z(n12668) );
  IV U12411 ( .A(p_input[2503]), .Z(n12511) );
  XOR U12412 ( .A(n12670), .B(n12671), .Z(n12666) );
  AND U12413 ( .A(n12672), .B(n12673), .Z(n12671) );
  XNOR U12414 ( .A(p_input[2518]), .B(n12670), .Z(n12673) );
  XNOR U12415 ( .A(n12670), .B(n12520), .Z(n12672) );
  IV U12416 ( .A(p_input[2502]), .Z(n12520) );
  XOR U12417 ( .A(n12674), .B(n12675), .Z(n12670) );
  AND U12418 ( .A(n12676), .B(n12677), .Z(n12675) );
  XNOR U12419 ( .A(p_input[2517]), .B(n12674), .Z(n12677) );
  XNOR U12420 ( .A(n12674), .B(n12529), .Z(n12676) );
  IV U12421 ( .A(p_input[2501]), .Z(n12529) );
  XOR U12422 ( .A(n12678), .B(n12679), .Z(n12674) );
  AND U12423 ( .A(n12680), .B(n12681), .Z(n12679) );
  XNOR U12424 ( .A(p_input[2516]), .B(n12678), .Z(n12681) );
  XNOR U12425 ( .A(n12678), .B(n12538), .Z(n12680) );
  IV U12426 ( .A(p_input[2500]), .Z(n12538) );
  XOR U12427 ( .A(n12682), .B(n12683), .Z(n12678) );
  AND U12428 ( .A(n12684), .B(n12685), .Z(n12683) );
  XNOR U12429 ( .A(p_input[2515]), .B(n12682), .Z(n12685) );
  XNOR U12430 ( .A(n12682), .B(n12547), .Z(n12684) );
  IV U12431 ( .A(p_input[2499]), .Z(n12547) );
  XOR U12432 ( .A(n12686), .B(n12687), .Z(n12682) );
  AND U12433 ( .A(n12688), .B(n12689), .Z(n12687) );
  XNOR U12434 ( .A(p_input[2514]), .B(n12686), .Z(n12689) );
  XNOR U12435 ( .A(n12686), .B(n12556), .Z(n12688) );
  IV U12436 ( .A(p_input[2498]), .Z(n12556) );
  XNOR U12437 ( .A(n12690), .B(n12691), .Z(n12686) );
  AND U12438 ( .A(n12692), .B(n12693), .Z(n12691) );
  XOR U12439 ( .A(p_input[2513]), .B(n12690), .Z(n12693) );
  XNOR U12440 ( .A(p_input[2497]), .B(n12690), .Z(n12692) );
  AND U12441 ( .A(p_input[2512]), .B(n12694), .Z(n12690) );
  IV U12442 ( .A(p_input[2496]), .Z(n12694) );
  XOR U12443 ( .A(n12695), .B(n12696), .Z(n12253) );
  AND U12444 ( .A(n445), .B(n12697), .Z(n12696) );
  XNOR U12445 ( .A(n12698), .B(n12695), .Z(n12697) );
  XOR U12446 ( .A(n12699), .B(n12700), .Z(n445) );
  AND U12447 ( .A(n12701), .B(n12702), .Z(n12700) );
  XNOR U12448 ( .A(n12263), .B(n12699), .Z(n12702) );
  AND U12449 ( .A(p_input[2495]), .B(p_input[2479]), .Z(n12263) );
  XOR U12450 ( .A(n12699), .B(n12264), .Z(n12701) );
  AND U12451 ( .A(p_input[2463]), .B(p_input[2447]), .Z(n12264) );
  XOR U12452 ( .A(n12703), .B(n12704), .Z(n12699) );
  AND U12453 ( .A(n12705), .B(n12706), .Z(n12704) );
  XOR U12454 ( .A(n12703), .B(n12276), .Z(n12706) );
  XNOR U12455 ( .A(p_input[2478]), .B(n12707), .Z(n12276) );
  AND U12456 ( .A(n295), .B(n12708), .Z(n12707) );
  XOR U12457 ( .A(p_input[2494]), .B(p_input[2478]), .Z(n12708) );
  XNOR U12458 ( .A(n12273), .B(n12703), .Z(n12705) );
  XOR U12459 ( .A(n12709), .B(n12710), .Z(n12273) );
  AND U12460 ( .A(n292), .B(n12711), .Z(n12710) );
  XOR U12461 ( .A(p_input[2462]), .B(p_input[2446]), .Z(n12711) );
  XOR U12462 ( .A(n12712), .B(n12713), .Z(n12703) );
  AND U12463 ( .A(n12714), .B(n12715), .Z(n12713) );
  XOR U12464 ( .A(n12712), .B(n12288), .Z(n12715) );
  XNOR U12465 ( .A(p_input[2477]), .B(n12716), .Z(n12288) );
  AND U12466 ( .A(n295), .B(n12717), .Z(n12716) );
  XOR U12467 ( .A(p_input[2493]), .B(p_input[2477]), .Z(n12717) );
  XNOR U12468 ( .A(n12285), .B(n12712), .Z(n12714) );
  XOR U12469 ( .A(n12718), .B(n12719), .Z(n12285) );
  AND U12470 ( .A(n292), .B(n12720), .Z(n12719) );
  XOR U12471 ( .A(p_input[2461]), .B(p_input[2445]), .Z(n12720) );
  XOR U12472 ( .A(n12721), .B(n12722), .Z(n12712) );
  AND U12473 ( .A(n12723), .B(n12724), .Z(n12722) );
  XOR U12474 ( .A(n12721), .B(n12300), .Z(n12724) );
  XNOR U12475 ( .A(p_input[2476]), .B(n12725), .Z(n12300) );
  AND U12476 ( .A(n295), .B(n12726), .Z(n12725) );
  XOR U12477 ( .A(p_input[2492]), .B(p_input[2476]), .Z(n12726) );
  XNOR U12478 ( .A(n12297), .B(n12721), .Z(n12723) );
  XOR U12479 ( .A(n12727), .B(n12728), .Z(n12297) );
  AND U12480 ( .A(n292), .B(n12729), .Z(n12728) );
  XOR U12481 ( .A(p_input[2460]), .B(p_input[2444]), .Z(n12729) );
  XOR U12482 ( .A(n12730), .B(n12731), .Z(n12721) );
  AND U12483 ( .A(n12732), .B(n12733), .Z(n12731) );
  XOR U12484 ( .A(n12730), .B(n12312), .Z(n12733) );
  XNOR U12485 ( .A(p_input[2475]), .B(n12734), .Z(n12312) );
  AND U12486 ( .A(n295), .B(n12735), .Z(n12734) );
  XOR U12487 ( .A(p_input[2491]), .B(p_input[2475]), .Z(n12735) );
  XNOR U12488 ( .A(n12309), .B(n12730), .Z(n12732) );
  XOR U12489 ( .A(n12736), .B(n12737), .Z(n12309) );
  AND U12490 ( .A(n292), .B(n12738), .Z(n12737) );
  XOR U12491 ( .A(p_input[2459]), .B(p_input[2443]), .Z(n12738) );
  XOR U12492 ( .A(n12739), .B(n12740), .Z(n12730) );
  AND U12493 ( .A(n12741), .B(n12742), .Z(n12740) );
  XOR U12494 ( .A(n12739), .B(n12324), .Z(n12742) );
  XNOR U12495 ( .A(p_input[2474]), .B(n12743), .Z(n12324) );
  AND U12496 ( .A(n295), .B(n12744), .Z(n12743) );
  XOR U12497 ( .A(p_input[2490]), .B(p_input[2474]), .Z(n12744) );
  XNOR U12498 ( .A(n12321), .B(n12739), .Z(n12741) );
  XOR U12499 ( .A(n12745), .B(n12746), .Z(n12321) );
  AND U12500 ( .A(n292), .B(n12747), .Z(n12746) );
  XOR U12501 ( .A(p_input[2458]), .B(p_input[2442]), .Z(n12747) );
  XOR U12502 ( .A(n12748), .B(n12749), .Z(n12739) );
  AND U12503 ( .A(n12750), .B(n12751), .Z(n12749) );
  XOR U12504 ( .A(n12748), .B(n12336), .Z(n12751) );
  XNOR U12505 ( .A(p_input[2473]), .B(n12752), .Z(n12336) );
  AND U12506 ( .A(n295), .B(n12753), .Z(n12752) );
  XOR U12507 ( .A(p_input[2489]), .B(p_input[2473]), .Z(n12753) );
  XNOR U12508 ( .A(n12333), .B(n12748), .Z(n12750) );
  XOR U12509 ( .A(n12754), .B(n12755), .Z(n12333) );
  AND U12510 ( .A(n292), .B(n12756), .Z(n12755) );
  XOR U12511 ( .A(p_input[2457]), .B(p_input[2441]), .Z(n12756) );
  XOR U12512 ( .A(n12757), .B(n12758), .Z(n12748) );
  AND U12513 ( .A(n12759), .B(n12760), .Z(n12758) );
  XOR U12514 ( .A(n12757), .B(n12348), .Z(n12760) );
  XNOR U12515 ( .A(p_input[2472]), .B(n12761), .Z(n12348) );
  AND U12516 ( .A(n295), .B(n12762), .Z(n12761) );
  XOR U12517 ( .A(p_input[2488]), .B(p_input[2472]), .Z(n12762) );
  XNOR U12518 ( .A(n12345), .B(n12757), .Z(n12759) );
  XOR U12519 ( .A(n12763), .B(n12764), .Z(n12345) );
  AND U12520 ( .A(n292), .B(n12765), .Z(n12764) );
  XOR U12521 ( .A(p_input[2456]), .B(p_input[2440]), .Z(n12765) );
  XOR U12522 ( .A(n12766), .B(n12767), .Z(n12757) );
  AND U12523 ( .A(n12768), .B(n12769), .Z(n12767) );
  XOR U12524 ( .A(n12766), .B(n12360), .Z(n12769) );
  XNOR U12525 ( .A(p_input[2471]), .B(n12770), .Z(n12360) );
  AND U12526 ( .A(n295), .B(n12771), .Z(n12770) );
  XOR U12527 ( .A(p_input[2487]), .B(p_input[2471]), .Z(n12771) );
  XNOR U12528 ( .A(n12357), .B(n12766), .Z(n12768) );
  XOR U12529 ( .A(n12772), .B(n12773), .Z(n12357) );
  AND U12530 ( .A(n292), .B(n12774), .Z(n12773) );
  XOR U12531 ( .A(p_input[2455]), .B(p_input[2439]), .Z(n12774) );
  XOR U12532 ( .A(n12775), .B(n12776), .Z(n12766) );
  AND U12533 ( .A(n12777), .B(n12778), .Z(n12776) );
  XOR U12534 ( .A(n12775), .B(n12372), .Z(n12778) );
  XNOR U12535 ( .A(p_input[2470]), .B(n12779), .Z(n12372) );
  AND U12536 ( .A(n295), .B(n12780), .Z(n12779) );
  XOR U12537 ( .A(p_input[2486]), .B(p_input[2470]), .Z(n12780) );
  XNOR U12538 ( .A(n12369), .B(n12775), .Z(n12777) );
  XOR U12539 ( .A(n12781), .B(n12782), .Z(n12369) );
  AND U12540 ( .A(n292), .B(n12783), .Z(n12782) );
  XOR U12541 ( .A(p_input[2454]), .B(p_input[2438]), .Z(n12783) );
  XOR U12542 ( .A(n12784), .B(n12785), .Z(n12775) );
  AND U12543 ( .A(n12786), .B(n12787), .Z(n12785) );
  XOR U12544 ( .A(n12784), .B(n12384), .Z(n12787) );
  XNOR U12545 ( .A(p_input[2469]), .B(n12788), .Z(n12384) );
  AND U12546 ( .A(n295), .B(n12789), .Z(n12788) );
  XOR U12547 ( .A(p_input[2485]), .B(p_input[2469]), .Z(n12789) );
  XNOR U12548 ( .A(n12381), .B(n12784), .Z(n12786) );
  XOR U12549 ( .A(n12790), .B(n12791), .Z(n12381) );
  AND U12550 ( .A(n292), .B(n12792), .Z(n12791) );
  XOR U12551 ( .A(p_input[2453]), .B(p_input[2437]), .Z(n12792) );
  XOR U12552 ( .A(n12793), .B(n12794), .Z(n12784) );
  AND U12553 ( .A(n12795), .B(n12796), .Z(n12794) );
  XOR U12554 ( .A(n12793), .B(n12396), .Z(n12796) );
  XNOR U12555 ( .A(p_input[2468]), .B(n12797), .Z(n12396) );
  AND U12556 ( .A(n295), .B(n12798), .Z(n12797) );
  XOR U12557 ( .A(p_input[2484]), .B(p_input[2468]), .Z(n12798) );
  XNOR U12558 ( .A(n12393), .B(n12793), .Z(n12795) );
  XOR U12559 ( .A(n12799), .B(n12800), .Z(n12393) );
  AND U12560 ( .A(n292), .B(n12801), .Z(n12800) );
  XOR U12561 ( .A(p_input[2452]), .B(p_input[2436]), .Z(n12801) );
  XOR U12562 ( .A(n12802), .B(n12803), .Z(n12793) );
  AND U12563 ( .A(n12804), .B(n12805), .Z(n12803) );
  XOR U12564 ( .A(n12802), .B(n12408), .Z(n12805) );
  XNOR U12565 ( .A(p_input[2467]), .B(n12806), .Z(n12408) );
  AND U12566 ( .A(n295), .B(n12807), .Z(n12806) );
  XOR U12567 ( .A(p_input[2483]), .B(p_input[2467]), .Z(n12807) );
  XNOR U12568 ( .A(n12405), .B(n12802), .Z(n12804) );
  XOR U12569 ( .A(n12808), .B(n12809), .Z(n12405) );
  AND U12570 ( .A(n292), .B(n12810), .Z(n12809) );
  XOR U12571 ( .A(p_input[2451]), .B(p_input[2435]), .Z(n12810) );
  XOR U12572 ( .A(n12811), .B(n12812), .Z(n12802) );
  AND U12573 ( .A(n12813), .B(n12814), .Z(n12812) );
  XOR U12574 ( .A(n12811), .B(n12420), .Z(n12814) );
  XNOR U12575 ( .A(p_input[2466]), .B(n12815), .Z(n12420) );
  AND U12576 ( .A(n295), .B(n12816), .Z(n12815) );
  XOR U12577 ( .A(p_input[2482]), .B(p_input[2466]), .Z(n12816) );
  XNOR U12578 ( .A(n12417), .B(n12811), .Z(n12813) );
  XOR U12579 ( .A(n12817), .B(n12818), .Z(n12417) );
  AND U12580 ( .A(n292), .B(n12819), .Z(n12818) );
  XOR U12581 ( .A(p_input[2450]), .B(p_input[2434]), .Z(n12819) );
  XOR U12582 ( .A(n12820), .B(n12821), .Z(n12811) );
  AND U12583 ( .A(n12822), .B(n12823), .Z(n12821) );
  XNOR U12584 ( .A(n12824), .B(n12433), .Z(n12823) );
  XNOR U12585 ( .A(p_input[2465]), .B(n12825), .Z(n12433) );
  AND U12586 ( .A(n295), .B(n12826), .Z(n12825) );
  XNOR U12587 ( .A(p_input[2481]), .B(n12827), .Z(n12826) );
  IV U12588 ( .A(p_input[2465]), .Z(n12827) );
  XNOR U12589 ( .A(n12430), .B(n12820), .Z(n12822) );
  XNOR U12590 ( .A(p_input[2433]), .B(n12828), .Z(n12430) );
  AND U12591 ( .A(n292), .B(n12829), .Z(n12828) );
  XOR U12592 ( .A(p_input[2449]), .B(p_input[2433]), .Z(n12829) );
  IV U12593 ( .A(n12824), .Z(n12820) );
  AND U12594 ( .A(n12695), .B(n12698), .Z(n12824) );
  XOR U12595 ( .A(p_input[2464]), .B(n12830), .Z(n12698) );
  AND U12596 ( .A(n295), .B(n12831), .Z(n12830) );
  XOR U12597 ( .A(p_input[2480]), .B(p_input[2464]), .Z(n12831) );
  XOR U12598 ( .A(n12832), .B(n12833), .Z(n295) );
  AND U12599 ( .A(n12834), .B(n12835), .Z(n12833) );
  XNOR U12600 ( .A(p_input[2495]), .B(n12832), .Z(n12835) );
  XOR U12601 ( .A(n12832), .B(p_input[2479]), .Z(n12834) );
  XOR U12602 ( .A(n12836), .B(n12837), .Z(n12832) );
  AND U12603 ( .A(n12838), .B(n12839), .Z(n12837) );
  XNOR U12604 ( .A(p_input[2494]), .B(n12836), .Z(n12839) );
  XOR U12605 ( .A(n12836), .B(p_input[2478]), .Z(n12838) );
  XOR U12606 ( .A(n12840), .B(n12841), .Z(n12836) );
  AND U12607 ( .A(n12842), .B(n12843), .Z(n12841) );
  XNOR U12608 ( .A(p_input[2493]), .B(n12840), .Z(n12843) );
  XOR U12609 ( .A(n12840), .B(p_input[2477]), .Z(n12842) );
  XOR U12610 ( .A(n12844), .B(n12845), .Z(n12840) );
  AND U12611 ( .A(n12846), .B(n12847), .Z(n12845) );
  XNOR U12612 ( .A(p_input[2492]), .B(n12844), .Z(n12847) );
  XOR U12613 ( .A(n12844), .B(p_input[2476]), .Z(n12846) );
  XOR U12614 ( .A(n12848), .B(n12849), .Z(n12844) );
  AND U12615 ( .A(n12850), .B(n12851), .Z(n12849) );
  XNOR U12616 ( .A(p_input[2491]), .B(n12848), .Z(n12851) );
  XOR U12617 ( .A(n12848), .B(p_input[2475]), .Z(n12850) );
  XOR U12618 ( .A(n12852), .B(n12853), .Z(n12848) );
  AND U12619 ( .A(n12854), .B(n12855), .Z(n12853) );
  XNOR U12620 ( .A(p_input[2490]), .B(n12852), .Z(n12855) );
  XOR U12621 ( .A(n12852), .B(p_input[2474]), .Z(n12854) );
  XOR U12622 ( .A(n12856), .B(n12857), .Z(n12852) );
  AND U12623 ( .A(n12858), .B(n12859), .Z(n12857) );
  XNOR U12624 ( .A(p_input[2489]), .B(n12856), .Z(n12859) );
  XOR U12625 ( .A(n12856), .B(p_input[2473]), .Z(n12858) );
  XOR U12626 ( .A(n12860), .B(n12861), .Z(n12856) );
  AND U12627 ( .A(n12862), .B(n12863), .Z(n12861) );
  XNOR U12628 ( .A(p_input[2488]), .B(n12860), .Z(n12863) );
  XOR U12629 ( .A(n12860), .B(p_input[2472]), .Z(n12862) );
  XOR U12630 ( .A(n12864), .B(n12865), .Z(n12860) );
  AND U12631 ( .A(n12866), .B(n12867), .Z(n12865) );
  XNOR U12632 ( .A(p_input[2487]), .B(n12864), .Z(n12867) );
  XOR U12633 ( .A(n12864), .B(p_input[2471]), .Z(n12866) );
  XOR U12634 ( .A(n12868), .B(n12869), .Z(n12864) );
  AND U12635 ( .A(n12870), .B(n12871), .Z(n12869) );
  XNOR U12636 ( .A(p_input[2486]), .B(n12868), .Z(n12871) );
  XOR U12637 ( .A(n12868), .B(p_input[2470]), .Z(n12870) );
  XOR U12638 ( .A(n12872), .B(n12873), .Z(n12868) );
  AND U12639 ( .A(n12874), .B(n12875), .Z(n12873) );
  XNOR U12640 ( .A(p_input[2485]), .B(n12872), .Z(n12875) );
  XOR U12641 ( .A(n12872), .B(p_input[2469]), .Z(n12874) );
  XOR U12642 ( .A(n12876), .B(n12877), .Z(n12872) );
  AND U12643 ( .A(n12878), .B(n12879), .Z(n12877) );
  XNOR U12644 ( .A(p_input[2484]), .B(n12876), .Z(n12879) );
  XOR U12645 ( .A(n12876), .B(p_input[2468]), .Z(n12878) );
  XOR U12646 ( .A(n12880), .B(n12881), .Z(n12876) );
  AND U12647 ( .A(n12882), .B(n12883), .Z(n12881) );
  XNOR U12648 ( .A(p_input[2483]), .B(n12880), .Z(n12883) );
  XOR U12649 ( .A(n12880), .B(p_input[2467]), .Z(n12882) );
  XOR U12650 ( .A(n12884), .B(n12885), .Z(n12880) );
  AND U12651 ( .A(n12886), .B(n12887), .Z(n12885) );
  XNOR U12652 ( .A(p_input[2482]), .B(n12884), .Z(n12887) );
  XOR U12653 ( .A(n12884), .B(p_input[2466]), .Z(n12886) );
  XNOR U12654 ( .A(n12888), .B(n12889), .Z(n12884) );
  AND U12655 ( .A(n12890), .B(n12891), .Z(n12889) );
  XOR U12656 ( .A(p_input[2481]), .B(n12888), .Z(n12891) );
  XNOR U12657 ( .A(p_input[2465]), .B(n12888), .Z(n12890) );
  AND U12658 ( .A(p_input[2480]), .B(n12892), .Z(n12888) );
  IV U12659 ( .A(p_input[2464]), .Z(n12892) );
  XNOR U12660 ( .A(p_input[2432]), .B(n12893), .Z(n12695) );
  AND U12661 ( .A(n292), .B(n12894), .Z(n12893) );
  XOR U12662 ( .A(p_input[2448]), .B(p_input[2432]), .Z(n12894) );
  XOR U12663 ( .A(n12895), .B(n12896), .Z(n292) );
  AND U12664 ( .A(n12897), .B(n12898), .Z(n12896) );
  XNOR U12665 ( .A(p_input[2463]), .B(n12895), .Z(n12898) );
  XOR U12666 ( .A(n12895), .B(p_input[2447]), .Z(n12897) );
  XOR U12667 ( .A(n12899), .B(n12900), .Z(n12895) );
  AND U12668 ( .A(n12901), .B(n12902), .Z(n12900) );
  XNOR U12669 ( .A(p_input[2462]), .B(n12899), .Z(n12902) );
  XNOR U12670 ( .A(n12899), .B(n12709), .Z(n12901) );
  IV U12671 ( .A(p_input[2446]), .Z(n12709) );
  XOR U12672 ( .A(n12903), .B(n12904), .Z(n12899) );
  AND U12673 ( .A(n12905), .B(n12906), .Z(n12904) );
  XNOR U12674 ( .A(p_input[2461]), .B(n12903), .Z(n12906) );
  XNOR U12675 ( .A(n12903), .B(n12718), .Z(n12905) );
  IV U12676 ( .A(p_input[2445]), .Z(n12718) );
  XOR U12677 ( .A(n12907), .B(n12908), .Z(n12903) );
  AND U12678 ( .A(n12909), .B(n12910), .Z(n12908) );
  XNOR U12679 ( .A(p_input[2460]), .B(n12907), .Z(n12910) );
  XNOR U12680 ( .A(n12907), .B(n12727), .Z(n12909) );
  IV U12681 ( .A(p_input[2444]), .Z(n12727) );
  XOR U12682 ( .A(n12911), .B(n12912), .Z(n12907) );
  AND U12683 ( .A(n12913), .B(n12914), .Z(n12912) );
  XNOR U12684 ( .A(p_input[2459]), .B(n12911), .Z(n12914) );
  XNOR U12685 ( .A(n12911), .B(n12736), .Z(n12913) );
  IV U12686 ( .A(p_input[2443]), .Z(n12736) );
  XOR U12687 ( .A(n12915), .B(n12916), .Z(n12911) );
  AND U12688 ( .A(n12917), .B(n12918), .Z(n12916) );
  XNOR U12689 ( .A(p_input[2458]), .B(n12915), .Z(n12918) );
  XNOR U12690 ( .A(n12915), .B(n12745), .Z(n12917) );
  IV U12691 ( .A(p_input[2442]), .Z(n12745) );
  XOR U12692 ( .A(n12919), .B(n12920), .Z(n12915) );
  AND U12693 ( .A(n12921), .B(n12922), .Z(n12920) );
  XNOR U12694 ( .A(p_input[2457]), .B(n12919), .Z(n12922) );
  XNOR U12695 ( .A(n12919), .B(n12754), .Z(n12921) );
  IV U12696 ( .A(p_input[2441]), .Z(n12754) );
  XOR U12697 ( .A(n12923), .B(n12924), .Z(n12919) );
  AND U12698 ( .A(n12925), .B(n12926), .Z(n12924) );
  XNOR U12699 ( .A(p_input[2456]), .B(n12923), .Z(n12926) );
  XNOR U12700 ( .A(n12923), .B(n12763), .Z(n12925) );
  IV U12701 ( .A(p_input[2440]), .Z(n12763) );
  XOR U12702 ( .A(n12927), .B(n12928), .Z(n12923) );
  AND U12703 ( .A(n12929), .B(n12930), .Z(n12928) );
  XNOR U12704 ( .A(p_input[2455]), .B(n12927), .Z(n12930) );
  XNOR U12705 ( .A(n12927), .B(n12772), .Z(n12929) );
  IV U12706 ( .A(p_input[2439]), .Z(n12772) );
  XOR U12707 ( .A(n12931), .B(n12932), .Z(n12927) );
  AND U12708 ( .A(n12933), .B(n12934), .Z(n12932) );
  XNOR U12709 ( .A(p_input[2454]), .B(n12931), .Z(n12934) );
  XNOR U12710 ( .A(n12931), .B(n12781), .Z(n12933) );
  IV U12711 ( .A(p_input[2438]), .Z(n12781) );
  XOR U12712 ( .A(n12935), .B(n12936), .Z(n12931) );
  AND U12713 ( .A(n12937), .B(n12938), .Z(n12936) );
  XNOR U12714 ( .A(p_input[2453]), .B(n12935), .Z(n12938) );
  XNOR U12715 ( .A(n12935), .B(n12790), .Z(n12937) );
  IV U12716 ( .A(p_input[2437]), .Z(n12790) );
  XOR U12717 ( .A(n12939), .B(n12940), .Z(n12935) );
  AND U12718 ( .A(n12941), .B(n12942), .Z(n12940) );
  XNOR U12719 ( .A(p_input[2452]), .B(n12939), .Z(n12942) );
  XNOR U12720 ( .A(n12939), .B(n12799), .Z(n12941) );
  IV U12721 ( .A(p_input[2436]), .Z(n12799) );
  XOR U12722 ( .A(n12943), .B(n12944), .Z(n12939) );
  AND U12723 ( .A(n12945), .B(n12946), .Z(n12944) );
  XNOR U12724 ( .A(p_input[2451]), .B(n12943), .Z(n12946) );
  XNOR U12725 ( .A(n12943), .B(n12808), .Z(n12945) );
  IV U12726 ( .A(p_input[2435]), .Z(n12808) );
  XOR U12727 ( .A(n12947), .B(n12948), .Z(n12943) );
  AND U12728 ( .A(n12949), .B(n12950), .Z(n12948) );
  XNOR U12729 ( .A(p_input[2450]), .B(n12947), .Z(n12950) );
  XNOR U12730 ( .A(n12947), .B(n12817), .Z(n12949) );
  IV U12731 ( .A(p_input[2434]), .Z(n12817) );
  XNOR U12732 ( .A(n12951), .B(n12952), .Z(n12947) );
  AND U12733 ( .A(n12953), .B(n12954), .Z(n12952) );
  XOR U12734 ( .A(p_input[2449]), .B(n12951), .Z(n12954) );
  XNOR U12735 ( .A(p_input[2433]), .B(n12951), .Z(n12953) );
  AND U12736 ( .A(p_input[2448]), .B(n12955), .Z(n12951) );
  IV U12737 ( .A(p_input[2432]), .Z(n12955) );
  XOR U12738 ( .A(n12956), .B(n12957), .Z(n12071) );
  AND U12739 ( .A(n773), .B(n12958), .Z(n12957) );
  XNOR U12740 ( .A(n12959), .B(n12956), .Z(n12958) );
  XOR U12741 ( .A(n12960), .B(n12961), .Z(n773) );
  AND U12742 ( .A(n12962), .B(n12963), .Z(n12961) );
  XNOR U12743 ( .A(n12083), .B(n12960), .Z(n12963) );
  AND U12744 ( .A(n12964), .B(n12965), .Z(n12083) );
  XOR U12745 ( .A(n12960), .B(n12082), .Z(n12962) );
  AND U12746 ( .A(n12966), .B(n12967), .Z(n12082) );
  XOR U12747 ( .A(n12968), .B(n12969), .Z(n12960) );
  AND U12748 ( .A(n12970), .B(n12971), .Z(n12969) );
  XOR U12749 ( .A(n12968), .B(n12095), .Z(n12971) );
  XOR U12750 ( .A(n12972), .B(n12973), .Z(n12095) );
  AND U12751 ( .A(n451), .B(n12974), .Z(n12973) );
  XOR U12752 ( .A(n12975), .B(n12972), .Z(n12974) );
  XNOR U12753 ( .A(n12092), .B(n12968), .Z(n12970) );
  XOR U12754 ( .A(n12976), .B(n12977), .Z(n12092) );
  AND U12755 ( .A(n448), .B(n12978), .Z(n12977) );
  XOR U12756 ( .A(n12979), .B(n12976), .Z(n12978) );
  XOR U12757 ( .A(n12980), .B(n12981), .Z(n12968) );
  AND U12758 ( .A(n12982), .B(n12983), .Z(n12981) );
  XOR U12759 ( .A(n12980), .B(n12107), .Z(n12983) );
  XOR U12760 ( .A(n12984), .B(n12985), .Z(n12107) );
  AND U12761 ( .A(n451), .B(n12986), .Z(n12985) );
  XOR U12762 ( .A(n12987), .B(n12984), .Z(n12986) );
  XNOR U12763 ( .A(n12104), .B(n12980), .Z(n12982) );
  XOR U12764 ( .A(n12988), .B(n12989), .Z(n12104) );
  AND U12765 ( .A(n448), .B(n12990), .Z(n12989) );
  XOR U12766 ( .A(n12991), .B(n12988), .Z(n12990) );
  XOR U12767 ( .A(n12992), .B(n12993), .Z(n12980) );
  AND U12768 ( .A(n12994), .B(n12995), .Z(n12993) );
  XOR U12769 ( .A(n12992), .B(n12119), .Z(n12995) );
  XOR U12770 ( .A(n12996), .B(n12997), .Z(n12119) );
  AND U12771 ( .A(n451), .B(n12998), .Z(n12997) );
  XOR U12772 ( .A(n12999), .B(n12996), .Z(n12998) );
  XNOR U12773 ( .A(n12116), .B(n12992), .Z(n12994) );
  XOR U12774 ( .A(n13000), .B(n13001), .Z(n12116) );
  AND U12775 ( .A(n448), .B(n13002), .Z(n13001) );
  XOR U12776 ( .A(n13003), .B(n13000), .Z(n13002) );
  XOR U12777 ( .A(n13004), .B(n13005), .Z(n12992) );
  AND U12778 ( .A(n13006), .B(n13007), .Z(n13005) );
  XOR U12779 ( .A(n13004), .B(n12131), .Z(n13007) );
  XOR U12780 ( .A(n13008), .B(n13009), .Z(n12131) );
  AND U12781 ( .A(n451), .B(n13010), .Z(n13009) );
  XOR U12782 ( .A(n13011), .B(n13008), .Z(n13010) );
  XNOR U12783 ( .A(n12128), .B(n13004), .Z(n13006) );
  XOR U12784 ( .A(n13012), .B(n13013), .Z(n12128) );
  AND U12785 ( .A(n448), .B(n13014), .Z(n13013) );
  XOR U12786 ( .A(n13015), .B(n13012), .Z(n13014) );
  XOR U12787 ( .A(n13016), .B(n13017), .Z(n13004) );
  AND U12788 ( .A(n13018), .B(n13019), .Z(n13017) );
  XOR U12789 ( .A(n13016), .B(n12143), .Z(n13019) );
  XOR U12790 ( .A(n13020), .B(n13021), .Z(n12143) );
  AND U12791 ( .A(n451), .B(n13022), .Z(n13021) );
  XOR U12792 ( .A(n13023), .B(n13020), .Z(n13022) );
  XNOR U12793 ( .A(n12140), .B(n13016), .Z(n13018) );
  XOR U12794 ( .A(n13024), .B(n13025), .Z(n12140) );
  AND U12795 ( .A(n448), .B(n13026), .Z(n13025) );
  XOR U12796 ( .A(n13027), .B(n13024), .Z(n13026) );
  XOR U12797 ( .A(n13028), .B(n13029), .Z(n13016) );
  AND U12798 ( .A(n13030), .B(n13031), .Z(n13029) );
  XOR U12799 ( .A(n13028), .B(n12155), .Z(n13031) );
  XOR U12800 ( .A(n13032), .B(n13033), .Z(n12155) );
  AND U12801 ( .A(n451), .B(n13034), .Z(n13033) );
  XOR U12802 ( .A(n13035), .B(n13032), .Z(n13034) );
  XNOR U12803 ( .A(n12152), .B(n13028), .Z(n13030) );
  XOR U12804 ( .A(n13036), .B(n13037), .Z(n12152) );
  AND U12805 ( .A(n448), .B(n13038), .Z(n13037) );
  XOR U12806 ( .A(n13039), .B(n13036), .Z(n13038) );
  XOR U12807 ( .A(n13040), .B(n13041), .Z(n13028) );
  AND U12808 ( .A(n13042), .B(n13043), .Z(n13041) );
  XOR U12809 ( .A(n13040), .B(n12167), .Z(n13043) );
  XOR U12810 ( .A(n13044), .B(n13045), .Z(n12167) );
  AND U12811 ( .A(n451), .B(n13046), .Z(n13045) );
  XOR U12812 ( .A(n13047), .B(n13044), .Z(n13046) );
  XNOR U12813 ( .A(n12164), .B(n13040), .Z(n13042) );
  XOR U12814 ( .A(n13048), .B(n13049), .Z(n12164) );
  AND U12815 ( .A(n448), .B(n13050), .Z(n13049) );
  XOR U12816 ( .A(n13051), .B(n13048), .Z(n13050) );
  XOR U12817 ( .A(n13052), .B(n13053), .Z(n13040) );
  AND U12818 ( .A(n13054), .B(n13055), .Z(n13053) );
  XOR U12819 ( .A(n13052), .B(n12179), .Z(n13055) );
  XOR U12820 ( .A(n13056), .B(n13057), .Z(n12179) );
  AND U12821 ( .A(n451), .B(n13058), .Z(n13057) );
  XOR U12822 ( .A(n13059), .B(n13056), .Z(n13058) );
  XNOR U12823 ( .A(n12176), .B(n13052), .Z(n13054) );
  XOR U12824 ( .A(n13060), .B(n13061), .Z(n12176) );
  AND U12825 ( .A(n448), .B(n13062), .Z(n13061) );
  XOR U12826 ( .A(n13063), .B(n13060), .Z(n13062) );
  XOR U12827 ( .A(n13064), .B(n13065), .Z(n13052) );
  AND U12828 ( .A(n13066), .B(n13067), .Z(n13065) );
  XOR U12829 ( .A(n13064), .B(n12191), .Z(n13067) );
  XOR U12830 ( .A(n13068), .B(n13069), .Z(n12191) );
  AND U12831 ( .A(n451), .B(n13070), .Z(n13069) );
  XOR U12832 ( .A(n13071), .B(n13068), .Z(n13070) );
  XNOR U12833 ( .A(n12188), .B(n13064), .Z(n13066) );
  XOR U12834 ( .A(n13072), .B(n13073), .Z(n12188) );
  AND U12835 ( .A(n448), .B(n13074), .Z(n13073) );
  XOR U12836 ( .A(n13075), .B(n13072), .Z(n13074) );
  XOR U12837 ( .A(n13076), .B(n13077), .Z(n13064) );
  AND U12838 ( .A(n13078), .B(n13079), .Z(n13077) );
  XOR U12839 ( .A(n13076), .B(n12203), .Z(n13079) );
  XOR U12840 ( .A(n13080), .B(n13081), .Z(n12203) );
  AND U12841 ( .A(n451), .B(n13082), .Z(n13081) );
  XOR U12842 ( .A(n13083), .B(n13080), .Z(n13082) );
  XNOR U12843 ( .A(n12200), .B(n13076), .Z(n13078) );
  XOR U12844 ( .A(n13084), .B(n13085), .Z(n12200) );
  AND U12845 ( .A(n448), .B(n13086), .Z(n13085) );
  XOR U12846 ( .A(n13087), .B(n13084), .Z(n13086) );
  XOR U12847 ( .A(n13088), .B(n13089), .Z(n13076) );
  AND U12848 ( .A(n13090), .B(n13091), .Z(n13089) );
  XOR U12849 ( .A(n13088), .B(n12215), .Z(n13091) );
  XOR U12850 ( .A(n13092), .B(n13093), .Z(n12215) );
  AND U12851 ( .A(n451), .B(n13094), .Z(n13093) );
  XOR U12852 ( .A(n13095), .B(n13092), .Z(n13094) );
  XNOR U12853 ( .A(n12212), .B(n13088), .Z(n13090) );
  XOR U12854 ( .A(n13096), .B(n13097), .Z(n12212) );
  AND U12855 ( .A(n448), .B(n13098), .Z(n13097) );
  XOR U12856 ( .A(n13099), .B(n13096), .Z(n13098) );
  XOR U12857 ( .A(n13100), .B(n13101), .Z(n13088) );
  AND U12858 ( .A(n13102), .B(n13103), .Z(n13101) );
  XOR U12859 ( .A(n13100), .B(n12227), .Z(n13103) );
  XOR U12860 ( .A(n13104), .B(n13105), .Z(n12227) );
  AND U12861 ( .A(n451), .B(n13106), .Z(n13105) );
  XOR U12862 ( .A(n13107), .B(n13104), .Z(n13106) );
  XNOR U12863 ( .A(n12224), .B(n13100), .Z(n13102) );
  XOR U12864 ( .A(n13108), .B(n13109), .Z(n12224) );
  AND U12865 ( .A(n448), .B(n13110), .Z(n13109) );
  XOR U12866 ( .A(n13111), .B(n13108), .Z(n13110) );
  XOR U12867 ( .A(n13112), .B(n13113), .Z(n13100) );
  AND U12868 ( .A(n13114), .B(n13115), .Z(n13113) );
  XOR U12869 ( .A(n13112), .B(n12239), .Z(n13115) );
  XOR U12870 ( .A(n13116), .B(n13117), .Z(n12239) );
  AND U12871 ( .A(n451), .B(n13118), .Z(n13117) );
  XOR U12872 ( .A(n13119), .B(n13116), .Z(n13118) );
  XNOR U12873 ( .A(n12236), .B(n13112), .Z(n13114) );
  XOR U12874 ( .A(n13120), .B(n13121), .Z(n12236) );
  AND U12875 ( .A(n448), .B(n13122), .Z(n13121) );
  XOR U12876 ( .A(n13123), .B(n13120), .Z(n13122) );
  XOR U12877 ( .A(n13124), .B(n13125), .Z(n13112) );
  AND U12878 ( .A(n13126), .B(n13127), .Z(n13125) );
  XNOR U12879 ( .A(n13128), .B(n12252), .Z(n13127) );
  XOR U12880 ( .A(n13129), .B(n13130), .Z(n12252) );
  AND U12881 ( .A(n451), .B(n13131), .Z(n13130) );
  XOR U12882 ( .A(n13129), .B(n13132), .Z(n13131) );
  XNOR U12883 ( .A(n12249), .B(n13124), .Z(n13126) );
  XOR U12884 ( .A(n13133), .B(n13134), .Z(n12249) );
  AND U12885 ( .A(n448), .B(n13135), .Z(n13134) );
  XOR U12886 ( .A(n13133), .B(n13136), .Z(n13135) );
  IV U12887 ( .A(n13128), .Z(n13124) );
  AND U12888 ( .A(n12956), .B(n12959), .Z(n13128) );
  XNOR U12889 ( .A(n13137), .B(n13138), .Z(n12959) );
  AND U12890 ( .A(n451), .B(n13139), .Z(n13138) );
  XNOR U12891 ( .A(n13140), .B(n13137), .Z(n13139) );
  XOR U12892 ( .A(n13141), .B(n13142), .Z(n451) );
  AND U12893 ( .A(n13143), .B(n13144), .Z(n13142) );
  XNOR U12894 ( .A(n12964), .B(n13141), .Z(n13144) );
  AND U12895 ( .A(p_input[2431]), .B(p_input[2415]), .Z(n12964) );
  XOR U12896 ( .A(n13141), .B(n12965), .Z(n13143) );
  AND U12897 ( .A(p_input[2399]), .B(p_input[2383]), .Z(n12965) );
  XOR U12898 ( .A(n13145), .B(n13146), .Z(n13141) );
  AND U12899 ( .A(n13147), .B(n13148), .Z(n13146) );
  XOR U12900 ( .A(n13145), .B(n12975), .Z(n13148) );
  XNOR U12901 ( .A(p_input[2414]), .B(n13149), .Z(n12975) );
  AND U12902 ( .A(n303), .B(n13150), .Z(n13149) );
  XOR U12903 ( .A(p_input[2430]), .B(p_input[2414]), .Z(n13150) );
  XNOR U12904 ( .A(n12972), .B(n13145), .Z(n13147) );
  XOR U12905 ( .A(n13151), .B(n13152), .Z(n12972) );
  AND U12906 ( .A(n301), .B(n13153), .Z(n13152) );
  XOR U12907 ( .A(p_input[2398]), .B(p_input[2382]), .Z(n13153) );
  XOR U12908 ( .A(n13154), .B(n13155), .Z(n13145) );
  AND U12909 ( .A(n13156), .B(n13157), .Z(n13155) );
  XOR U12910 ( .A(n13154), .B(n12987), .Z(n13157) );
  XNOR U12911 ( .A(p_input[2413]), .B(n13158), .Z(n12987) );
  AND U12912 ( .A(n303), .B(n13159), .Z(n13158) );
  XOR U12913 ( .A(p_input[2429]), .B(p_input[2413]), .Z(n13159) );
  XNOR U12914 ( .A(n12984), .B(n13154), .Z(n13156) );
  XOR U12915 ( .A(n13160), .B(n13161), .Z(n12984) );
  AND U12916 ( .A(n301), .B(n13162), .Z(n13161) );
  XOR U12917 ( .A(p_input[2397]), .B(p_input[2381]), .Z(n13162) );
  XOR U12918 ( .A(n13163), .B(n13164), .Z(n13154) );
  AND U12919 ( .A(n13165), .B(n13166), .Z(n13164) );
  XOR U12920 ( .A(n13163), .B(n12999), .Z(n13166) );
  XNOR U12921 ( .A(p_input[2412]), .B(n13167), .Z(n12999) );
  AND U12922 ( .A(n303), .B(n13168), .Z(n13167) );
  XOR U12923 ( .A(p_input[2428]), .B(p_input[2412]), .Z(n13168) );
  XNOR U12924 ( .A(n12996), .B(n13163), .Z(n13165) );
  XOR U12925 ( .A(n13169), .B(n13170), .Z(n12996) );
  AND U12926 ( .A(n301), .B(n13171), .Z(n13170) );
  XOR U12927 ( .A(p_input[2396]), .B(p_input[2380]), .Z(n13171) );
  XOR U12928 ( .A(n13172), .B(n13173), .Z(n13163) );
  AND U12929 ( .A(n13174), .B(n13175), .Z(n13173) );
  XOR U12930 ( .A(n13172), .B(n13011), .Z(n13175) );
  XNOR U12931 ( .A(p_input[2411]), .B(n13176), .Z(n13011) );
  AND U12932 ( .A(n303), .B(n13177), .Z(n13176) );
  XOR U12933 ( .A(p_input[2427]), .B(p_input[2411]), .Z(n13177) );
  XNOR U12934 ( .A(n13008), .B(n13172), .Z(n13174) );
  XOR U12935 ( .A(n13178), .B(n13179), .Z(n13008) );
  AND U12936 ( .A(n301), .B(n13180), .Z(n13179) );
  XOR U12937 ( .A(p_input[2395]), .B(p_input[2379]), .Z(n13180) );
  XOR U12938 ( .A(n13181), .B(n13182), .Z(n13172) );
  AND U12939 ( .A(n13183), .B(n13184), .Z(n13182) );
  XOR U12940 ( .A(n13181), .B(n13023), .Z(n13184) );
  XNOR U12941 ( .A(p_input[2410]), .B(n13185), .Z(n13023) );
  AND U12942 ( .A(n303), .B(n13186), .Z(n13185) );
  XOR U12943 ( .A(p_input[2426]), .B(p_input[2410]), .Z(n13186) );
  XNOR U12944 ( .A(n13020), .B(n13181), .Z(n13183) );
  XOR U12945 ( .A(n13187), .B(n13188), .Z(n13020) );
  AND U12946 ( .A(n301), .B(n13189), .Z(n13188) );
  XOR U12947 ( .A(p_input[2394]), .B(p_input[2378]), .Z(n13189) );
  XOR U12948 ( .A(n13190), .B(n13191), .Z(n13181) );
  AND U12949 ( .A(n13192), .B(n13193), .Z(n13191) );
  XOR U12950 ( .A(n13190), .B(n13035), .Z(n13193) );
  XNOR U12951 ( .A(p_input[2409]), .B(n13194), .Z(n13035) );
  AND U12952 ( .A(n303), .B(n13195), .Z(n13194) );
  XOR U12953 ( .A(p_input[2425]), .B(p_input[2409]), .Z(n13195) );
  XNOR U12954 ( .A(n13032), .B(n13190), .Z(n13192) );
  XOR U12955 ( .A(n13196), .B(n13197), .Z(n13032) );
  AND U12956 ( .A(n301), .B(n13198), .Z(n13197) );
  XOR U12957 ( .A(p_input[2393]), .B(p_input[2377]), .Z(n13198) );
  XOR U12958 ( .A(n13199), .B(n13200), .Z(n13190) );
  AND U12959 ( .A(n13201), .B(n13202), .Z(n13200) );
  XOR U12960 ( .A(n13199), .B(n13047), .Z(n13202) );
  XNOR U12961 ( .A(p_input[2408]), .B(n13203), .Z(n13047) );
  AND U12962 ( .A(n303), .B(n13204), .Z(n13203) );
  XOR U12963 ( .A(p_input[2424]), .B(p_input[2408]), .Z(n13204) );
  XNOR U12964 ( .A(n13044), .B(n13199), .Z(n13201) );
  XOR U12965 ( .A(n13205), .B(n13206), .Z(n13044) );
  AND U12966 ( .A(n301), .B(n13207), .Z(n13206) );
  XOR U12967 ( .A(p_input[2392]), .B(p_input[2376]), .Z(n13207) );
  XOR U12968 ( .A(n13208), .B(n13209), .Z(n13199) );
  AND U12969 ( .A(n13210), .B(n13211), .Z(n13209) );
  XOR U12970 ( .A(n13208), .B(n13059), .Z(n13211) );
  XNOR U12971 ( .A(p_input[2407]), .B(n13212), .Z(n13059) );
  AND U12972 ( .A(n303), .B(n13213), .Z(n13212) );
  XOR U12973 ( .A(p_input[2423]), .B(p_input[2407]), .Z(n13213) );
  XNOR U12974 ( .A(n13056), .B(n13208), .Z(n13210) );
  XOR U12975 ( .A(n13214), .B(n13215), .Z(n13056) );
  AND U12976 ( .A(n301), .B(n13216), .Z(n13215) );
  XOR U12977 ( .A(p_input[2391]), .B(p_input[2375]), .Z(n13216) );
  XOR U12978 ( .A(n13217), .B(n13218), .Z(n13208) );
  AND U12979 ( .A(n13219), .B(n13220), .Z(n13218) );
  XOR U12980 ( .A(n13217), .B(n13071), .Z(n13220) );
  XNOR U12981 ( .A(p_input[2406]), .B(n13221), .Z(n13071) );
  AND U12982 ( .A(n303), .B(n13222), .Z(n13221) );
  XOR U12983 ( .A(p_input[2422]), .B(p_input[2406]), .Z(n13222) );
  XNOR U12984 ( .A(n13068), .B(n13217), .Z(n13219) );
  XOR U12985 ( .A(n13223), .B(n13224), .Z(n13068) );
  AND U12986 ( .A(n301), .B(n13225), .Z(n13224) );
  XOR U12987 ( .A(p_input[2390]), .B(p_input[2374]), .Z(n13225) );
  XOR U12988 ( .A(n13226), .B(n13227), .Z(n13217) );
  AND U12989 ( .A(n13228), .B(n13229), .Z(n13227) );
  XOR U12990 ( .A(n13226), .B(n13083), .Z(n13229) );
  XNOR U12991 ( .A(p_input[2405]), .B(n13230), .Z(n13083) );
  AND U12992 ( .A(n303), .B(n13231), .Z(n13230) );
  XOR U12993 ( .A(p_input[2421]), .B(p_input[2405]), .Z(n13231) );
  XNOR U12994 ( .A(n13080), .B(n13226), .Z(n13228) );
  XOR U12995 ( .A(n13232), .B(n13233), .Z(n13080) );
  AND U12996 ( .A(n301), .B(n13234), .Z(n13233) );
  XOR U12997 ( .A(p_input[2389]), .B(p_input[2373]), .Z(n13234) );
  XOR U12998 ( .A(n13235), .B(n13236), .Z(n13226) );
  AND U12999 ( .A(n13237), .B(n13238), .Z(n13236) );
  XOR U13000 ( .A(n13235), .B(n13095), .Z(n13238) );
  XNOR U13001 ( .A(p_input[2404]), .B(n13239), .Z(n13095) );
  AND U13002 ( .A(n303), .B(n13240), .Z(n13239) );
  XOR U13003 ( .A(p_input[2420]), .B(p_input[2404]), .Z(n13240) );
  XNOR U13004 ( .A(n13092), .B(n13235), .Z(n13237) );
  XOR U13005 ( .A(n13241), .B(n13242), .Z(n13092) );
  AND U13006 ( .A(n301), .B(n13243), .Z(n13242) );
  XOR U13007 ( .A(p_input[2388]), .B(p_input[2372]), .Z(n13243) );
  XOR U13008 ( .A(n13244), .B(n13245), .Z(n13235) );
  AND U13009 ( .A(n13246), .B(n13247), .Z(n13245) );
  XOR U13010 ( .A(n13244), .B(n13107), .Z(n13247) );
  XNOR U13011 ( .A(p_input[2403]), .B(n13248), .Z(n13107) );
  AND U13012 ( .A(n303), .B(n13249), .Z(n13248) );
  XOR U13013 ( .A(p_input[2419]), .B(p_input[2403]), .Z(n13249) );
  XNOR U13014 ( .A(n13104), .B(n13244), .Z(n13246) );
  XOR U13015 ( .A(n13250), .B(n13251), .Z(n13104) );
  AND U13016 ( .A(n301), .B(n13252), .Z(n13251) );
  XOR U13017 ( .A(p_input[2387]), .B(p_input[2371]), .Z(n13252) );
  XOR U13018 ( .A(n13253), .B(n13254), .Z(n13244) );
  AND U13019 ( .A(n13255), .B(n13256), .Z(n13254) );
  XOR U13020 ( .A(n13253), .B(n13119), .Z(n13256) );
  XNOR U13021 ( .A(p_input[2402]), .B(n13257), .Z(n13119) );
  AND U13022 ( .A(n303), .B(n13258), .Z(n13257) );
  XOR U13023 ( .A(p_input[2418]), .B(p_input[2402]), .Z(n13258) );
  XNOR U13024 ( .A(n13116), .B(n13253), .Z(n13255) );
  XOR U13025 ( .A(n13259), .B(n13260), .Z(n13116) );
  AND U13026 ( .A(n301), .B(n13261), .Z(n13260) );
  XOR U13027 ( .A(p_input[2386]), .B(p_input[2370]), .Z(n13261) );
  XOR U13028 ( .A(n13262), .B(n13263), .Z(n13253) );
  AND U13029 ( .A(n13264), .B(n13265), .Z(n13263) );
  XNOR U13030 ( .A(n13266), .B(n13132), .Z(n13265) );
  XNOR U13031 ( .A(p_input[2401]), .B(n13267), .Z(n13132) );
  AND U13032 ( .A(n303), .B(n13268), .Z(n13267) );
  XNOR U13033 ( .A(p_input[2417]), .B(n13269), .Z(n13268) );
  IV U13034 ( .A(p_input[2401]), .Z(n13269) );
  XNOR U13035 ( .A(n13129), .B(n13262), .Z(n13264) );
  XNOR U13036 ( .A(p_input[2369]), .B(n13270), .Z(n13129) );
  AND U13037 ( .A(n301), .B(n13271), .Z(n13270) );
  XOR U13038 ( .A(p_input[2385]), .B(p_input[2369]), .Z(n13271) );
  IV U13039 ( .A(n13266), .Z(n13262) );
  AND U13040 ( .A(n13137), .B(n13140), .Z(n13266) );
  XOR U13041 ( .A(p_input[2400]), .B(n13272), .Z(n13140) );
  AND U13042 ( .A(n303), .B(n13273), .Z(n13272) );
  XOR U13043 ( .A(p_input[2416]), .B(p_input[2400]), .Z(n13273) );
  XOR U13044 ( .A(n13274), .B(n13275), .Z(n303) );
  AND U13045 ( .A(n13276), .B(n13277), .Z(n13275) );
  XNOR U13046 ( .A(p_input[2431]), .B(n13274), .Z(n13277) );
  XOR U13047 ( .A(n13274), .B(p_input[2415]), .Z(n13276) );
  XOR U13048 ( .A(n13278), .B(n13279), .Z(n13274) );
  AND U13049 ( .A(n13280), .B(n13281), .Z(n13279) );
  XNOR U13050 ( .A(p_input[2430]), .B(n13278), .Z(n13281) );
  XOR U13051 ( .A(n13278), .B(p_input[2414]), .Z(n13280) );
  XOR U13052 ( .A(n13282), .B(n13283), .Z(n13278) );
  AND U13053 ( .A(n13284), .B(n13285), .Z(n13283) );
  XNOR U13054 ( .A(p_input[2429]), .B(n13282), .Z(n13285) );
  XOR U13055 ( .A(n13282), .B(p_input[2413]), .Z(n13284) );
  XOR U13056 ( .A(n13286), .B(n13287), .Z(n13282) );
  AND U13057 ( .A(n13288), .B(n13289), .Z(n13287) );
  XNOR U13058 ( .A(p_input[2428]), .B(n13286), .Z(n13289) );
  XOR U13059 ( .A(n13286), .B(p_input[2412]), .Z(n13288) );
  XOR U13060 ( .A(n13290), .B(n13291), .Z(n13286) );
  AND U13061 ( .A(n13292), .B(n13293), .Z(n13291) );
  XNOR U13062 ( .A(p_input[2427]), .B(n13290), .Z(n13293) );
  XOR U13063 ( .A(n13290), .B(p_input[2411]), .Z(n13292) );
  XOR U13064 ( .A(n13294), .B(n13295), .Z(n13290) );
  AND U13065 ( .A(n13296), .B(n13297), .Z(n13295) );
  XNOR U13066 ( .A(p_input[2426]), .B(n13294), .Z(n13297) );
  XOR U13067 ( .A(n13294), .B(p_input[2410]), .Z(n13296) );
  XOR U13068 ( .A(n13298), .B(n13299), .Z(n13294) );
  AND U13069 ( .A(n13300), .B(n13301), .Z(n13299) );
  XNOR U13070 ( .A(p_input[2425]), .B(n13298), .Z(n13301) );
  XOR U13071 ( .A(n13298), .B(p_input[2409]), .Z(n13300) );
  XOR U13072 ( .A(n13302), .B(n13303), .Z(n13298) );
  AND U13073 ( .A(n13304), .B(n13305), .Z(n13303) );
  XNOR U13074 ( .A(p_input[2424]), .B(n13302), .Z(n13305) );
  XOR U13075 ( .A(n13302), .B(p_input[2408]), .Z(n13304) );
  XOR U13076 ( .A(n13306), .B(n13307), .Z(n13302) );
  AND U13077 ( .A(n13308), .B(n13309), .Z(n13307) );
  XNOR U13078 ( .A(p_input[2423]), .B(n13306), .Z(n13309) );
  XOR U13079 ( .A(n13306), .B(p_input[2407]), .Z(n13308) );
  XOR U13080 ( .A(n13310), .B(n13311), .Z(n13306) );
  AND U13081 ( .A(n13312), .B(n13313), .Z(n13311) );
  XNOR U13082 ( .A(p_input[2422]), .B(n13310), .Z(n13313) );
  XOR U13083 ( .A(n13310), .B(p_input[2406]), .Z(n13312) );
  XOR U13084 ( .A(n13314), .B(n13315), .Z(n13310) );
  AND U13085 ( .A(n13316), .B(n13317), .Z(n13315) );
  XNOR U13086 ( .A(p_input[2421]), .B(n13314), .Z(n13317) );
  XOR U13087 ( .A(n13314), .B(p_input[2405]), .Z(n13316) );
  XOR U13088 ( .A(n13318), .B(n13319), .Z(n13314) );
  AND U13089 ( .A(n13320), .B(n13321), .Z(n13319) );
  XNOR U13090 ( .A(p_input[2420]), .B(n13318), .Z(n13321) );
  XOR U13091 ( .A(n13318), .B(p_input[2404]), .Z(n13320) );
  XOR U13092 ( .A(n13322), .B(n13323), .Z(n13318) );
  AND U13093 ( .A(n13324), .B(n13325), .Z(n13323) );
  XNOR U13094 ( .A(p_input[2419]), .B(n13322), .Z(n13325) );
  XOR U13095 ( .A(n13322), .B(p_input[2403]), .Z(n13324) );
  XOR U13096 ( .A(n13326), .B(n13327), .Z(n13322) );
  AND U13097 ( .A(n13328), .B(n13329), .Z(n13327) );
  XNOR U13098 ( .A(p_input[2418]), .B(n13326), .Z(n13329) );
  XOR U13099 ( .A(n13326), .B(p_input[2402]), .Z(n13328) );
  XNOR U13100 ( .A(n13330), .B(n13331), .Z(n13326) );
  AND U13101 ( .A(n13332), .B(n13333), .Z(n13331) );
  XOR U13102 ( .A(p_input[2417]), .B(n13330), .Z(n13333) );
  XNOR U13103 ( .A(p_input[2401]), .B(n13330), .Z(n13332) );
  AND U13104 ( .A(p_input[2416]), .B(n13334), .Z(n13330) );
  IV U13105 ( .A(p_input[2400]), .Z(n13334) );
  XNOR U13106 ( .A(p_input[2368]), .B(n13335), .Z(n13137) );
  AND U13107 ( .A(n301), .B(n13336), .Z(n13335) );
  XOR U13108 ( .A(p_input[2384]), .B(p_input[2368]), .Z(n13336) );
  XOR U13109 ( .A(n13337), .B(n13338), .Z(n301) );
  AND U13110 ( .A(n13339), .B(n13340), .Z(n13338) );
  XNOR U13111 ( .A(p_input[2399]), .B(n13337), .Z(n13340) );
  XOR U13112 ( .A(n13337), .B(p_input[2383]), .Z(n13339) );
  XOR U13113 ( .A(n13341), .B(n13342), .Z(n13337) );
  AND U13114 ( .A(n13343), .B(n13344), .Z(n13342) );
  XNOR U13115 ( .A(p_input[2398]), .B(n13341), .Z(n13344) );
  XNOR U13116 ( .A(n13341), .B(n13151), .Z(n13343) );
  IV U13117 ( .A(p_input[2382]), .Z(n13151) );
  XOR U13118 ( .A(n13345), .B(n13346), .Z(n13341) );
  AND U13119 ( .A(n13347), .B(n13348), .Z(n13346) );
  XNOR U13120 ( .A(p_input[2397]), .B(n13345), .Z(n13348) );
  XNOR U13121 ( .A(n13345), .B(n13160), .Z(n13347) );
  IV U13122 ( .A(p_input[2381]), .Z(n13160) );
  XOR U13123 ( .A(n13349), .B(n13350), .Z(n13345) );
  AND U13124 ( .A(n13351), .B(n13352), .Z(n13350) );
  XNOR U13125 ( .A(p_input[2396]), .B(n13349), .Z(n13352) );
  XNOR U13126 ( .A(n13349), .B(n13169), .Z(n13351) );
  IV U13127 ( .A(p_input[2380]), .Z(n13169) );
  XOR U13128 ( .A(n13353), .B(n13354), .Z(n13349) );
  AND U13129 ( .A(n13355), .B(n13356), .Z(n13354) );
  XNOR U13130 ( .A(p_input[2395]), .B(n13353), .Z(n13356) );
  XNOR U13131 ( .A(n13353), .B(n13178), .Z(n13355) );
  IV U13132 ( .A(p_input[2379]), .Z(n13178) );
  XOR U13133 ( .A(n13357), .B(n13358), .Z(n13353) );
  AND U13134 ( .A(n13359), .B(n13360), .Z(n13358) );
  XNOR U13135 ( .A(p_input[2394]), .B(n13357), .Z(n13360) );
  XNOR U13136 ( .A(n13357), .B(n13187), .Z(n13359) );
  IV U13137 ( .A(p_input[2378]), .Z(n13187) );
  XOR U13138 ( .A(n13361), .B(n13362), .Z(n13357) );
  AND U13139 ( .A(n13363), .B(n13364), .Z(n13362) );
  XNOR U13140 ( .A(p_input[2393]), .B(n13361), .Z(n13364) );
  XNOR U13141 ( .A(n13361), .B(n13196), .Z(n13363) );
  IV U13142 ( .A(p_input[2377]), .Z(n13196) );
  XOR U13143 ( .A(n13365), .B(n13366), .Z(n13361) );
  AND U13144 ( .A(n13367), .B(n13368), .Z(n13366) );
  XNOR U13145 ( .A(p_input[2392]), .B(n13365), .Z(n13368) );
  XNOR U13146 ( .A(n13365), .B(n13205), .Z(n13367) );
  IV U13147 ( .A(p_input[2376]), .Z(n13205) );
  XOR U13148 ( .A(n13369), .B(n13370), .Z(n13365) );
  AND U13149 ( .A(n13371), .B(n13372), .Z(n13370) );
  XNOR U13150 ( .A(p_input[2391]), .B(n13369), .Z(n13372) );
  XNOR U13151 ( .A(n13369), .B(n13214), .Z(n13371) );
  IV U13152 ( .A(p_input[2375]), .Z(n13214) );
  XOR U13153 ( .A(n13373), .B(n13374), .Z(n13369) );
  AND U13154 ( .A(n13375), .B(n13376), .Z(n13374) );
  XNOR U13155 ( .A(p_input[2390]), .B(n13373), .Z(n13376) );
  XNOR U13156 ( .A(n13373), .B(n13223), .Z(n13375) );
  IV U13157 ( .A(p_input[2374]), .Z(n13223) );
  XOR U13158 ( .A(n13377), .B(n13378), .Z(n13373) );
  AND U13159 ( .A(n13379), .B(n13380), .Z(n13378) );
  XNOR U13160 ( .A(p_input[2389]), .B(n13377), .Z(n13380) );
  XNOR U13161 ( .A(n13377), .B(n13232), .Z(n13379) );
  IV U13162 ( .A(p_input[2373]), .Z(n13232) );
  XOR U13163 ( .A(n13381), .B(n13382), .Z(n13377) );
  AND U13164 ( .A(n13383), .B(n13384), .Z(n13382) );
  XNOR U13165 ( .A(p_input[2388]), .B(n13381), .Z(n13384) );
  XNOR U13166 ( .A(n13381), .B(n13241), .Z(n13383) );
  IV U13167 ( .A(p_input[2372]), .Z(n13241) );
  XOR U13168 ( .A(n13385), .B(n13386), .Z(n13381) );
  AND U13169 ( .A(n13387), .B(n13388), .Z(n13386) );
  XNOR U13170 ( .A(p_input[2387]), .B(n13385), .Z(n13388) );
  XNOR U13171 ( .A(n13385), .B(n13250), .Z(n13387) );
  IV U13172 ( .A(p_input[2371]), .Z(n13250) );
  XOR U13173 ( .A(n13389), .B(n13390), .Z(n13385) );
  AND U13174 ( .A(n13391), .B(n13392), .Z(n13390) );
  XNOR U13175 ( .A(p_input[2386]), .B(n13389), .Z(n13392) );
  XNOR U13176 ( .A(n13389), .B(n13259), .Z(n13391) );
  IV U13177 ( .A(p_input[2370]), .Z(n13259) );
  XNOR U13178 ( .A(n13393), .B(n13394), .Z(n13389) );
  AND U13179 ( .A(n13395), .B(n13396), .Z(n13394) );
  XOR U13180 ( .A(p_input[2385]), .B(n13393), .Z(n13396) );
  XNOR U13181 ( .A(p_input[2369]), .B(n13393), .Z(n13395) );
  AND U13182 ( .A(p_input[2384]), .B(n13397), .Z(n13393) );
  IV U13183 ( .A(p_input[2368]), .Z(n13397) );
  XOR U13184 ( .A(n13398), .B(n13399), .Z(n12956) );
  AND U13185 ( .A(n448), .B(n13400), .Z(n13399) );
  XNOR U13186 ( .A(n13401), .B(n13398), .Z(n13400) );
  XOR U13187 ( .A(n13402), .B(n13403), .Z(n448) );
  AND U13188 ( .A(n13404), .B(n13405), .Z(n13403) );
  XNOR U13189 ( .A(n12967), .B(n13402), .Z(n13405) );
  AND U13190 ( .A(p_input[2367]), .B(p_input[2351]), .Z(n12967) );
  XOR U13191 ( .A(n13402), .B(n12966), .Z(n13404) );
  AND U13192 ( .A(p_input[2319]), .B(p_input[2335]), .Z(n12966) );
  XOR U13193 ( .A(n13406), .B(n13407), .Z(n13402) );
  AND U13194 ( .A(n13408), .B(n13409), .Z(n13407) );
  XOR U13195 ( .A(n13406), .B(n12979), .Z(n13409) );
  XNOR U13196 ( .A(p_input[2350]), .B(n13410), .Z(n12979) );
  AND U13197 ( .A(n307), .B(n13411), .Z(n13410) );
  XOR U13198 ( .A(p_input[2366]), .B(p_input[2350]), .Z(n13411) );
  XNOR U13199 ( .A(n12976), .B(n13406), .Z(n13408) );
  XOR U13200 ( .A(n13412), .B(n13413), .Z(n12976) );
  AND U13201 ( .A(n304), .B(n13414), .Z(n13413) );
  XOR U13202 ( .A(p_input[2334]), .B(p_input[2318]), .Z(n13414) );
  XOR U13203 ( .A(n13415), .B(n13416), .Z(n13406) );
  AND U13204 ( .A(n13417), .B(n13418), .Z(n13416) );
  XOR U13205 ( .A(n13415), .B(n12991), .Z(n13418) );
  XNOR U13206 ( .A(p_input[2349]), .B(n13419), .Z(n12991) );
  AND U13207 ( .A(n307), .B(n13420), .Z(n13419) );
  XOR U13208 ( .A(p_input[2365]), .B(p_input[2349]), .Z(n13420) );
  XNOR U13209 ( .A(n12988), .B(n13415), .Z(n13417) );
  XOR U13210 ( .A(n13421), .B(n13422), .Z(n12988) );
  AND U13211 ( .A(n304), .B(n13423), .Z(n13422) );
  XOR U13212 ( .A(p_input[2333]), .B(p_input[2317]), .Z(n13423) );
  XOR U13213 ( .A(n13424), .B(n13425), .Z(n13415) );
  AND U13214 ( .A(n13426), .B(n13427), .Z(n13425) );
  XOR U13215 ( .A(n13424), .B(n13003), .Z(n13427) );
  XNOR U13216 ( .A(p_input[2348]), .B(n13428), .Z(n13003) );
  AND U13217 ( .A(n307), .B(n13429), .Z(n13428) );
  XOR U13218 ( .A(p_input[2364]), .B(p_input[2348]), .Z(n13429) );
  XNOR U13219 ( .A(n13000), .B(n13424), .Z(n13426) );
  XOR U13220 ( .A(n13430), .B(n13431), .Z(n13000) );
  AND U13221 ( .A(n304), .B(n13432), .Z(n13431) );
  XOR U13222 ( .A(p_input[2332]), .B(p_input[2316]), .Z(n13432) );
  XOR U13223 ( .A(n13433), .B(n13434), .Z(n13424) );
  AND U13224 ( .A(n13435), .B(n13436), .Z(n13434) );
  XOR U13225 ( .A(n13433), .B(n13015), .Z(n13436) );
  XNOR U13226 ( .A(p_input[2347]), .B(n13437), .Z(n13015) );
  AND U13227 ( .A(n307), .B(n13438), .Z(n13437) );
  XOR U13228 ( .A(p_input[2363]), .B(p_input[2347]), .Z(n13438) );
  XNOR U13229 ( .A(n13012), .B(n13433), .Z(n13435) );
  XOR U13230 ( .A(n13439), .B(n13440), .Z(n13012) );
  AND U13231 ( .A(n304), .B(n13441), .Z(n13440) );
  XOR U13232 ( .A(p_input[2331]), .B(p_input[2315]), .Z(n13441) );
  XOR U13233 ( .A(n13442), .B(n13443), .Z(n13433) );
  AND U13234 ( .A(n13444), .B(n13445), .Z(n13443) );
  XOR U13235 ( .A(n13442), .B(n13027), .Z(n13445) );
  XNOR U13236 ( .A(p_input[2346]), .B(n13446), .Z(n13027) );
  AND U13237 ( .A(n307), .B(n13447), .Z(n13446) );
  XOR U13238 ( .A(p_input[2362]), .B(p_input[2346]), .Z(n13447) );
  XNOR U13239 ( .A(n13024), .B(n13442), .Z(n13444) );
  XOR U13240 ( .A(n13448), .B(n13449), .Z(n13024) );
  AND U13241 ( .A(n304), .B(n13450), .Z(n13449) );
  XOR U13242 ( .A(p_input[2330]), .B(p_input[2314]), .Z(n13450) );
  XOR U13243 ( .A(n13451), .B(n13452), .Z(n13442) );
  AND U13244 ( .A(n13453), .B(n13454), .Z(n13452) );
  XOR U13245 ( .A(n13451), .B(n13039), .Z(n13454) );
  XNOR U13246 ( .A(p_input[2345]), .B(n13455), .Z(n13039) );
  AND U13247 ( .A(n307), .B(n13456), .Z(n13455) );
  XOR U13248 ( .A(p_input[2361]), .B(p_input[2345]), .Z(n13456) );
  XNOR U13249 ( .A(n13036), .B(n13451), .Z(n13453) );
  XOR U13250 ( .A(n13457), .B(n13458), .Z(n13036) );
  AND U13251 ( .A(n304), .B(n13459), .Z(n13458) );
  XOR U13252 ( .A(p_input[2329]), .B(p_input[2313]), .Z(n13459) );
  XOR U13253 ( .A(n13460), .B(n13461), .Z(n13451) );
  AND U13254 ( .A(n13462), .B(n13463), .Z(n13461) );
  XOR U13255 ( .A(n13460), .B(n13051), .Z(n13463) );
  XNOR U13256 ( .A(p_input[2344]), .B(n13464), .Z(n13051) );
  AND U13257 ( .A(n307), .B(n13465), .Z(n13464) );
  XOR U13258 ( .A(p_input[2360]), .B(p_input[2344]), .Z(n13465) );
  XNOR U13259 ( .A(n13048), .B(n13460), .Z(n13462) );
  XOR U13260 ( .A(n13466), .B(n13467), .Z(n13048) );
  AND U13261 ( .A(n304), .B(n13468), .Z(n13467) );
  XOR U13262 ( .A(p_input[2328]), .B(p_input[2312]), .Z(n13468) );
  XOR U13263 ( .A(n13469), .B(n13470), .Z(n13460) );
  AND U13264 ( .A(n13471), .B(n13472), .Z(n13470) );
  XOR U13265 ( .A(n13469), .B(n13063), .Z(n13472) );
  XNOR U13266 ( .A(p_input[2343]), .B(n13473), .Z(n13063) );
  AND U13267 ( .A(n307), .B(n13474), .Z(n13473) );
  XOR U13268 ( .A(p_input[2359]), .B(p_input[2343]), .Z(n13474) );
  XNOR U13269 ( .A(n13060), .B(n13469), .Z(n13471) );
  XOR U13270 ( .A(n13475), .B(n13476), .Z(n13060) );
  AND U13271 ( .A(n304), .B(n13477), .Z(n13476) );
  XOR U13272 ( .A(p_input[2327]), .B(p_input[2311]), .Z(n13477) );
  XOR U13273 ( .A(n13478), .B(n13479), .Z(n13469) );
  AND U13274 ( .A(n13480), .B(n13481), .Z(n13479) );
  XOR U13275 ( .A(n13478), .B(n13075), .Z(n13481) );
  XNOR U13276 ( .A(p_input[2342]), .B(n13482), .Z(n13075) );
  AND U13277 ( .A(n307), .B(n13483), .Z(n13482) );
  XOR U13278 ( .A(p_input[2358]), .B(p_input[2342]), .Z(n13483) );
  XNOR U13279 ( .A(n13072), .B(n13478), .Z(n13480) );
  XOR U13280 ( .A(n13484), .B(n13485), .Z(n13072) );
  AND U13281 ( .A(n304), .B(n13486), .Z(n13485) );
  XOR U13282 ( .A(p_input[2326]), .B(p_input[2310]), .Z(n13486) );
  XOR U13283 ( .A(n13487), .B(n13488), .Z(n13478) );
  AND U13284 ( .A(n13489), .B(n13490), .Z(n13488) );
  XOR U13285 ( .A(n13487), .B(n13087), .Z(n13490) );
  XNOR U13286 ( .A(p_input[2341]), .B(n13491), .Z(n13087) );
  AND U13287 ( .A(n307), .B(n13492), .Z(n13491) );
  XOR U13288 ( .A(p_input[2357]), .B(p_input[2341]), .Z(n13492) );
  XNOR U13289 ( .A(n13084), .B(n13487), .Z(n13489) );
  XOR U13290 ( .A(n13493), .B(n13494), .Z(n13084) );
  AND U13291 ( .A(n304), .B(n13495), .Z(n13494) );
  XOR U13292 ( .A(p_input[2325]), .B(p_input[2309]), .Z(n13495) );
  XOR U13293 ( .A(n13496), .B(n13497), .Z(n13487) );
  AND U13294 ( .A(n13498), .B(n13499), .Z(n13497) );
  XOR U13295 ( .A(n13496), .B(n13099), .Z(n13499) );
  XNOR U13296 ( .A(p_input[2340]), .B(n13500), .Z(n13099) );
  AND U13297 ( .A(n307), .B(n13501), .Z(n13500) );
  XOR U13298 ( .A(p_input[2356]), .B(p_input[2340]), .Z(n13501) );
  XNOR U13299 ( .A(n13096), .B(n13496), .Z(n13498) );
  XOR U13300 ( .A(n13502), .B(n13503), .Z(n13096) );
  AND U13301 ( .A(n304), .B(n13504), .Z(n13503) );
  XOR U13302 ( .A(p_input[2324]), .B(p_input[2308]), .Z(n13504) );
  XOR U13303 ( .A(n13505), .B(n13506), .Z(n13496) );
  AND U13304 ( .A(n13507), .B(n13508), .Z(n13506) );
  XOR U13305 ( .A(n13505), .B(n13111), .Z(n13508) );
  XNOR U13306 ( .A(p_input[2339]), .B(n13509), .Z(n13111) );
  AND U13307 ( .A(n307), .B(n13510), .Z(n13509) );
  XOR U13308 ( .A(p_input[2355]), .B(p_input[2339]), .Z(n13510) );
  XNOR U13309 ( .A(n13108), .B(n13505), .Z(n13507) );
  XOR U13310 ( .A(n13511), .B(n13512), .Z(n13108) );
  AND U13311 ( .A(n304), .B(n13513), .Z(n13512) );
  XOR U13312 ( .A(p_input[2323]), .B(p_input[2307]), .Z(n13513) );
  XOR U13313 ( .A(n13514), .B(n13515), .Z(n13505) );
  AND U13314 ( .A(n13516), .B(n13517), .Z(n13515) );
  XOR U13315 ( .A(n13514), .B(n13123), .Z(n13517) );
  XNOR U13316 ( .A(p_input[2338]), .B(n13518), .Z(n13123) );
  AND U13317 ( .A(n307), .B(n13519), .Z(n13518) );
  XOR U13318 ( .A(p_input[2354]), .B(p_input[2338]), .Z(n13519) );
  XNOR U13319 ( .A(n13120), .B(n13514), .Z(n13516) );
  XOR U13320 ( .A(n13520), .B(n13521), .Z(n13120) );
  AND U13321 ( .A(n304), .B(n13522), .Z(n13521) );
  XOR U13322 ( .A(p_input[2322]), .B(p_input[2306]), .Z(n13522) );
  XOR U13323 ( .A(n13523), .B(n13524), .Z(n13514) );
  AND U13324 ( .A(n13525), .B(n13526), .Z(n13524) );
  XNOR U13325 ( .A(n13527), .B(n13136), .Z(n13526) );
  XNOR U13326 ( .A(p_input[2337]), .B(n13528), .Z(n13136) );
  AND U13327 ( .A(n307), .B(n13529), .Z(n13528) );
  XNOR U13328 ( .A(p_input[2353]), .B(n13530), .Z(n13529) );
  IV U13329 ( .A(p_input[2337]), .Z(n13530) );
  XNOR U13330 ( .A(n13133), .B(n13523), .Z(n13525) );
  XNOR U13331 ( .A(p_input[2305]), .B(n13531), .Z(n13133) );
  AND U13332 ( .A(n304), .B(n13532), .Z(n13531) );
  XOR U13333 ( .A(p_input[2321]), .B(p_input[2305]), .Z(n13532) );
  IV U13334 ( .A(n13527), .Z(n13523) );
  AND U13335 ( .A(n13398), .B(n13401), .Z(n13527) );
  XOR U13336 ( .A(p_input[2336]), .B(n13533), .Z(n13401) );
  AND U13337 ( .A(n307), .B(n13534), .Z(n13533) );
  XOR U13338 ( .A(p_input[2352]), .B(p_input[2336]), .Z(n13534) );
  XOR U13339 ( .A(n13535), .B(n13536), .Z(n307) );
  AND U13340 ( .A(n13537), .B(n13538), .Z(n13536) );
  XNOR U13341 ( .A(p_input[2367]), .B(n13535), .Z(n13538) );
  XOR U13342 ( .A(n13535), .B(p_input[2351]), .Z(n13537) );
  XOR U13343 ( .A(n13539), .B(n13540), .Z(n13535) );
  AND U13344 ( .A(n13541), .B(n13542), .Z(n13540) );
  XNOR U13345 ( .A(p_input[2366]), .B(n13539), .Z(n13542) );
  XOR U13346 ( .A(n13539), .B(p_input[2350]), .Z(n13541) );
  XOR U13347 ( .A(n13543), .B(n13544), .Z(n13539) );
  AND U13348 ( .A(n13545), .B(n13546), .Z(n13544) );
  XNOR U13349 ( .A(p_input[2365]), .B(n13543), .Z(n13546) );
  XOR U13350 ( .A(n13543), .B(p_input[2349]), .Z(n13545) );
  XOR U13351 ( .A(n13547), .B(n13548), .Z(n13543) );
  AND U13352 ( .A(n13549), .B(n13550), .Z(n13548) );
  XNOR U13353 ( .A(p_input[2364]), .B(n13547), .Z(n13550) );
  XOR U13354 ( .A(n13547), .B(p_input[2348]), .Z(n13549) );
  XOR U13355 ( .A(n13551), .B(n13552), .Z(n13547) );
  AND U13356 ( .A(n13553), .B(n13554), .Z(n13552) );
  XNOR U13357 ( .A(p_input[2363]), .B(n13551), .Z(n13554) );
  XOR U13358 ( .A(n13551), .B(p_input[2347]), .Z(n13553) );
  XOR U13359 ( .A(n13555), .B(n13556), .Z(n13551) );
  AND U13360 ( .A(n13557), .B(n13558), .Z(n13556) );
  XNOR U13361 ( .A(p_input[2362]), .B(n13555), .Z(n13558) );
  XOR U13362 ( .A(n13555), .B(p_input[2346]), .Z(n13557) );
  XOR U13363 ( .A(n13559), .B(n13560), .Z(n13555) );
  AND U13364 ( .A(n13561), .B(n13562), .Z(n13560) );
  XNOR U13365 ( .A(p_input[2361]), .B(n13559), .Z(n13562) );
  XOR U13366 ( .A(n13559), .B(p_input[2345]), .Z(n13561) );
  XOR U13367 ( .A(n13563), .B(n13564), .Z(n13559) );
  AND U13368 ( .A(n13565), .B(n13566), .Z(n13564) );
  XNOR U13369 ( .A(p_input[2360]), .B(n13563), .Z(n13566) );
  XOR U13370 ( .A(n13563), .B(p_input[2344]), .Z(n13565) );
  XOR U13371 ( .A(n13567), .B(n13568), .Z(n13563) );
  AND U13372 ( .A(n13569), .B(n13570), .Z(n13568) );
  XNOR U13373 ( .A(p_input[2359]), .B(n13567), .Z(n13570) );
  XOR U13374 ( .A(n13567), .B(p_input[2343]), .Z(n13569) );
  XOR U13375 ( .A(n13571), .B(n13572), .Z(n13567) );
  AND U13376 ( .A(n13573), .B(n13574), .Z(n13572) );
  XNOR U13377 ( .A(p_input[2358]), .B(n13571), .Z(n13574) );
  XOR U13378 ( .A(n13571), .B(p_input[2342]), .Z(n13573) );
  XOR U13379 ( .A(n13575), .B(n13576), .Z(n13571) );
  AND U13380 ( .A(n13577), .B(n13578), .Z(n13576) );
  XNOR U13381 ( .A(p_input[2357]), .B(n13575), .Z(n13578) );
  XOR U13382 ( .A(n13575), .B(p_input[2341]), .Z(n13577) );
  XOR U13383 ( .A(n13579), .B(n13580), .Z(n13575) );
  AND U13384 ( .A(n13581), .B(n13582), .Z(n13580) );
  XNOR U13385 ( .A(p_input[2356]), .B(n13579), .Z(n13582) );
  XOR U13386 ( .A(n13579), .B(p_input[2340]), .Z(n13581) );
  XOR U13387 ( .A(n13583), .B(n13584), .Z(n13579) );
  AND U13388 ( .A(n13585), .B(n13586), .Z(n13584) );
  XNOR U13389 ( .A(p_input[2355]), .B(n13583), .Z(n13586) );
  XOR U13390 ( .A(n13583), .B(p_input[2339]), .Z(n13585) );
  XOR U13391 ( .A(n13587), .B(n13588), .Z(n13583) );
  AND U13392 ( .A(n13589), .B(n13590), .Z(n13588) );
  XNOR U13393 ( .A(p_input[2354]), .B(n13587), .Z(n13590) );
  XOR U13394 ( .A(n13587), .B(p_input[2338]), .Z(n13589) );
  XNOR U13395 ( .A(n13591), .B(n13592), .Z(n13587) );
  AND U13396 ( .A(n13593), .B(n13594), .Z(n13592) );
  XOR U13397 ( .A(p_input[2353]), .B(n13591), .Z(n13594) );
  XNOR U13398 ( .A(p_input[2337]), .B(n13591), .Z(n13593) );
  AND U13399 ( .A(p_input[2352]), .B(n13595), .Z(n13591) );
  IV U13400 ( .A(p_input[2336]), .Z(n13595) );
  XNOR U13401 ( .A(p_input[2304]), .B(n13596), .Z(n13398) );
  AND U13402 ( .A(n304), .B(n13597), .Z(n13596) );
  XOR U13403 ( .A(p_input[2320]), .B(p_input[2304]), .Z(n13597) );
  XOR U13404 ( .A(n13598), .B(n13599), .Z(n304) );
  AND U13405 ( .A(n13600), .B(n13601), .Z(n13599) );
  XNOR U13406 ( .A(p_input[2335]), .B(n13598), .Z(n13601) );
  XOR U13407 ( .A(n13598), .B(p_input[2319]), .Z(n13600) );
  XOR U13408 ( .A(n13602), .B(n13603), .Z(n13598) );
  AND U13409 ( .A(n13604), .B(n13605), .Z(n13603) );
  XNOR U13410 ( .A(p_input[2334]), .B(n13602), .Z(n13605) );
  XNOR U13411 ( .A(n13602), .B(n13412), .Z(n13604) );
  IV U13412 ( .A(p_input[2318]), .Z(n13412) );
  XOR U13413 ( .A(n13606), .B(n13607), .Z(n13602) );
  AND U13414 ( .A(n13608), .B(n13609), .Z(n13607) );
  XNOR U13415 ( .A(p_input[2333]), .B(n13606), .Z(n13609) );
  XNOR U13416 ( .A(n13606), .B(n13421), .Z(n13608) );
  IV U13417 ( .A(p_input[2317]), .Z(n13421) );
  XOR U13418 ( .A(n13610), .B(n13611), .Z(n13606) );
  AND U13419 ( .A(n13612), .B(n13613), .Z(n13611) );
  XNOR U13420 ( .A(p_input[2332]), .B(n13610), .Z(n13613) );
  XNOR U13421 ( .A(n13610), .B(n13430), .Z(n13612) );
  IV U13422 ( .A(p_input[2316]), .Z(n13430) );
  XOR U13423 ( .A(n13614), .B(n13615), .Z(n13610) );
  AND U13424 ( .A(n13616), .B(n13617), .Z(n13615) );
  XNOR U13425 ( .A(p_input[2331]), .B(n13614), .Z(n13617) );
  XNOR U13426 ( .A(n13614), .B(n13439), .Z(n13616) );
  IV U13427 ( .A(p_input[2315]), .Z(n13439) );
  XOR U13428 ( .A(n13618), .B(n13619), .Z(n13614) );
  AND U13429 ( .A(n13620), .B(n13621), .Z(n13619) );
  XNOR U13430 ( .A(p_input[2330]), .B(n13618), .Z(n13621) );
  XNOR U13431 ( .A(n13618), .B(n13448), .Z(n13620) );
  IV U13432 ( .A(p_input[2314]), .Z(n13448) );
  XOR U13433 ( .A(n13622), .B(n13623), .Z(n13618) );
  AND U13434 ( .A(n13624), .B(n13625), .Z(n13623) );
  XNOR U13435 ( .A(p_input[2329]), .B(n13622), .Z(n13625) );
  XNOR U13436 ( .A(n13622), .B(n13457), .Z(n13624) );
  IV U13437 ( .A(p_input[2313]), .Z(n13457) );
  XOR U13438 ( .A(n13626), .B(n13627), .Z(n13622) );
  AND U13439 ( .A(n13628), .B(n13629), .Z(n13627) );
  XNOR U13440 ( .A(p_input[2328]), .B(n13626), .Z(n13629) );
  XNOR U13441 ( .A(n13626), .B(n13466), .Z(n13628) );
  IV U13442 ( .A(p_input[2312]), .Z(n13466) );
  XOR U13443 ( .A(n13630), .B(n13631), .Z(n13626) );
  AND U13444 ( .A(n13632), .B(n13633), .Z(n13631) );
  XNOR U13445 ( .A(p_input[2327]), .B(n13630), .Z(n13633) );
  XNOR U13446 ( .A(n13630), .B(n13475), .Z(n13632) );
  IV U13447 ( .A(p_input[2311]), .Z(n13475) );
  XOR U13448 ( .A(n13634), .B(n13635), .Z(n13630) );
  AND U13449 ( .A(n13636), .B(n13637), .Z(n13635) );
  XNOR U13450 ( .A(p_input[2326]), .B(n13634), .Z(n13637) );
  XNOR U13451 ( .A(n13634), .B(n13484), .Z(n13636) );
  IV U13452 ( .A(p_input[2310]), .Z(n13484) );
  XOR U13453 ( .A(n13638), .B(n13639), .Z(n13634) );
  AND U13454 ( .A(n13640), .B(n13641), .Z(n13639) );
  XNOR U13455 ( .A(p_input[2325]), .B(n13638), .Z(n13641) );
  XNOR U13456 ( .A(n13638), .B(n13493), .Z(n13640) );
  IV U13457 ( .A(p_input[2309]), .Z(n13493) );
  XOR U13458 ( .A(n13642), .B(n13643), .Z(n13638) );
  AND U13459 ( .A(n13644), .B(n13645), .Z(n13643) );
  XNOR U13460 ( .A(p_input[2324]), .B(n13642), .Z(n13645) );
  XNOR U13461 ( .A(n13642), .B(n13502), .Z(n13644) );
  IV U13462 ( .A(p_input[2308]), .Z(n13502) );
  XOR U13463 ( .A(n13646), .B(n13647), .Z(n13642) );
  AND U13464 ( .A(n13648), .B(n13649), .Z(n13647) );
  XNOR U13465 ( .A(p_input[2323]), .B(n13646), .Z(n13649) );
  XNOR U13466 ( .A(n13646), .B(n13511), .Z(n13648) );
  IV U13467 ( .A(p_input[2307]), .Z(n13511) );
  XOR U13468 ( .A(n13650), .B(n13651), .Z(n13646) );
  AND U13469 ( .A(n13652), .B(n13653), .Z(n13651) );
  XNOR U13470 ( .A(p_input[2322]), .B(n13650), .Z(n13653) );
  XNOR U13471 ( .A(n13650), .B(n13520), .Z(n13652) );
  IV U13472 ( .A(p_input[2306]), .Z(n13520) );
  XNOR U13473 ( .A(n13654), .B(n13655), .Z(n13650) );
  AND U13474 ( .A(n13656), .B(n13657), .Z(n13655) );
  XOR U13475 ( .A(p_input[2321]), .B(n13654), .Z(n13657) );
  XNOR U13476 ( .A(p_input[2305]), .B(n13654), .Z(n13656) );
  AND U13477 ( .A(p_input[2320]), .B(n13658), .Z(n13654) );
  IV U13478 ( .A(p_input[2304]), .Z(n13658) );
  XOR U13479 ( .A(n13659), .B(n13660), .Z(n11886) );
  AND U13480 ( .A(n932), .B(n13661), .Z(n13660) );
  XNOR U13481 ( .A(n13662), .B(n13659), .Z(n13661) );
  XOR U13482 ( .A(n13663), .B(n13664), .Z(n932) );
  AND U13483 ( .A(n13665), .B(n13666), .Z(n13664) );
  XNOR U13484 ( .A(n11901), .B(n13663), .Z(n13666) );
  AND U13485 ( .A(n13667), .B(n13668), .Z(n11901) );
  XNOR U13486 ( .A(n13663), .B(n11898), .Z(n13665) );
  IV U13487 ( .A(n13669), .Z(n11898) );
  AND U13488 ( .A(n13670), .B(n13671), .Z(n13669) );
  XOR U13489 ( .A(n13672), .B(n13673), .Z(n13663) );
  AND U13490 ( .A(n13674), .B(n13675), .Z(n13673) );
  XOR U13491 ( .A(n13672), .B(n11913), .Z(n13675) );
  XOR U13492 ( .A(n13676), .B(n13677), .Z(n11913) );
  AND U13493 ( .A(n779), .B(n13678), .Z(n13677) );
  XOR U13494 ( .A(n13679), .B(n13676), .Z(n13678) );
  XNOR U13495 ( .A(n11910), .B(n13672), .Z(n13674) );
  XOR U13496 ( .A(n13680), .B(n13681), .Z(n11910) );
  AND U13497 ( .A(n776), .B(n13682), .Z(n13681) );
  XOR U13498 ( .A(n13683), .B(n13680), .Z(n13682) );
  XOR U13499 ( .A(n13684), .B(n13685), .Z(n13672) );
  AND U13500 ( .A(n13686), .B(n13687), .Z(n13685) );
  XOR U13501 ( .A(n13684), .B(n11925), .Z(n13687) );
  XOR U13502 ( .A(n13688), .B(n13689), .Z(n11925) );
  AND U13503 ( .A(n779), .B(n13690), .Z(n13689) );
  XOR U13504 ( .A(n13691), .B(n13688), .Z(n13690) );
  XNOR U13505 ( .A(n11922), .B(n13684), .Z(n13686) );
  XOR U13506 ( .A(n13692), .B(n13693), .Z(n11922) );
  AND U13507 ( .A(n776), .B(n13694), .Z(n13693) );
  XOR U13508 ( .A(n13695), .B(n13692), .Z(n13694) );
  XOR U13509 ( .A(n13696), .B(n13697), .Z(n13684) );
  AND U13510 ( .A(n13698), .B(n13699), .Z(n13697) );
  XOR U13511 ( .A(n13696), .B(n11937), .Z(n13699) );
  XOR U13512 ( .A(n13700), .B(n13701), .Z(n11937) );
  AND U13513 ( .A(n779), .B(n13702), .Z(n13701) );
  XOR U13514 ( .A(n13703), .B(n13700), .Z(n13702) );
  XNOR U13515 ( .A(n11934), .B(n13696), .Z(n13698) );
  XOR U13516 ( .A(n13704), .B(n13705), .Z(n11934) );
  AND U13517 ( .A(n776), .B(n13706), .Z(n13705) );
  XOR U13518 ( .A(n13707), .B(n13704), .Z(n13706) );
  XOR U13519 ( .A(n13708), .B(n13709), .Z(n13696) );
  AND U13520 ( .A(n13710), .B(n13711), .Z(n13709) );
  XOR U13521 ( .A(n13708), .B(n11949), .Z(n13711) );
  XOR U13522 ( .A(n13712), .B(n13713), .Z(n11949) );
  AND U13523 ( .A(n779), .B(n13714), .Z(n13713) );
  XOR U13524 ( .A(n13715), .B(n13712), .Z(n13714) );
  XNOR U13525 ( .A(n11946), .B(n13708), .Z(n13710) );
  XOR U13526 ( .A(n13716), .B(n13717), .Z(n11946) );
  AND U13527 ( .A(n776), .B(n13718), .Z(n13717) );
  XOR U13528 ( .A(n13719), .B(n13716), .Z(n13718) );
  XOR U13529 ( .A(n13720), .B(n13721), .Z(n13708) );
  AND U13530 ( .A(n13722), .B(n13723), .Z(n13721) );
  XOR U13531 ( .A(n13720), .B(n11961), .Z(n13723) );
  XOR U13532 ( .A(n13724), .B(n13725), .Z(n11961) );
  AND U13533 ( .A(n779), .B(n13726), .Z(n13725) );
  XOR U13534 ( .A(n13727), .B(n13724), .Z(n13726) );
  XNOR U13535 ( .A(n11958), .B(n13720), .Z(n13722) );
  XOR U13536 ( .A(n13728), .B(n13729), .Z(n11958) );
  AND U13537 ( .A(n776), .B(n13730), .Z(n13729) );
  XOR U13538 ( .A(n13731), .B(n13728), .Z(n13730) );
  XOR U13539 ( .A(n13732), .B(n13733), .Z(n13720) );
  AND U13540 ( .A(n13734), .B(n13735), .Z(n13733) );
  XOR U13541 ( .A(n13732), .B(n11973), .Z(n13735) );
  XOR U13542 ( .A(n13736), .B(n13737), .Z(n11973) );
  AND U13543 ( .A(n779), .B(n13738), .Z(n13737) );
  XOR U13544 ( .A(n13739), .B(n13736), .Z(n13738) );
  XNOR U13545 ( .A(n11970), .B(n13732), .Z(n13734) );
  XOR U13546 ( .A(n13740), .B(n13741), .Z(n11970) );
  AND U13547 ( .A(n776), .B(n13742), .Z(n13741) );
  XOR U13548 ( .A(n13743), .B(n13740), .Z(n13742) );
  XOR U13549 ( .A(n13744), .B(n13745), .Z(n13732) );
  AND U13550 ( .A(n13746), .B(n13747), .Z(n13745) );
  XOR U13551 ( .A(n13744), .B(n11985), .Z(n13747) );
  XOR U13552 ( .A(n13748), .B(n13749), .Z(n11985) );
  AND U13553 ( .A(n779), .B(n13750), .Z(n13749) );
  XOR U13554 ( .A(n13751), .B(n13748), .Z(n13750) );
  XNOR U13555 ( .A(n11982), .B(n13744), .Z(n13746) );
  XOR U13556 ( .A(n13752), .B(n13753), .Z(n11982) );
  AND U13557 ( .A(n776), .B(n13754), .Z(n13753) );
  XOR U13558 ( .A(n13755), .B(n13752), .Z(n13754) );
  XOR U13559 ( .A(n13756), .B(n13757), .Z(n13744) );
  AND U13560 ( .A(n13758), .B(n13759), .Z(n13757) );
  XOR U13561 ( .A(n13756), .B(n11997), .Z(n13759) );
  XOR U13562 ( .A(n13760), .B(n13761), .Z(n11997) );
  AND U13563 ( .A(n779), .B(n13762), .Z(n13761) );
  XOR U13564 ( .A(n13763), .B(n13760), .Z(n13762) );
  XNOR U13565 ( .A(n11994), .B(n13756), .Z(n13758) );
  XOR U13566 ( .A(n13764), .B(n13765), .Z(n11994) );
  AND U13567 ( .A(n776), .B(n13766), .Z(n13765) );
  XOR U13568 ( .A(n13767), .B(n13764), .Z(n13766) );
  XOR U13569 ( .A(n13768), .B(n13769), .Z(n13756) );
  AND U13570 ( .A(n13770), .B(n13771), .Z(n13769) );
  XOR U13571 ( .A(n13768), .B(n12009), .Z(n13771) );
  XOR U13572 ( .A(n13772), .B(n13773), .Z(n12009) );
  AND U13573 ( .A(n779), .B(n13774), .Z(n13773) );
  XOR U13574 ( .A(n13775), .B(n13772), .Z(n13774) );
  XNOR U13575 ( .A(n12006), .B(n13768), .Z(n13770) );
  XOR U13576 ( .A(n13776), .B(n13777), .Z(n12006) );
  AND U13577 ( .A(n776), .B(n13778), .Z(n13777) );
  XOR U13578 ( .A(n13779), .B(n13776), .Z(n13778) );
  XOR U13579 ( .A(n13780), .B(n13781), .Z(n13768) );
  AND U13580 ( .A(n13782), .B(n13783), .Z(n13781) );
  XOR U13581 ( .A(n13780), .B(n12021), .Z(n13783) );
  XOR U13582 ( .A(n13784), .B(n13785), .Z(n12021) );
  AND U13583 ( .A(n779), .B(n13786), .Z(n13785) );
  XOR U13584 ( .A(n13787), .B(n13784), .Z(n13786) );
  XNOR U13585 ( .A(n12018), .B(n13780), .Z(n13782) );
  XOR U13586 ( .A(n13788), .B(n13789), .Z(n12018) );
  AND U13587 ( .A(n776), .B(n13790), .Z(n13789) );
  XOR U13588 ( .A(n13791), .B(n13788), .Z(n13790) );
  XOR U13589 ( .A(n13792), .B(n13793), .Z(n13780) );
  AND U13590 ( .A(n13794), .B(n13795), .Z(n13793) );
  XOR U13591 ( .A(n13792), .B(n12033), .Z(n13795) );
  XOR U13592 ( .A(n13796), .B(n13797), .Z(n12033) );
  AND U13593 ( .A(n779), .B(n13798), .Z(n13797) );
  XOR U13594 ( .A(n13799), .B(n13796), .Z(n13798) );
  XNOR U13595 ( .A(n12030), .B(n13792), .Z(n13794) );
  XOR U13596 ( .A(n13800), .B(n13801), .Z(n12030) );
  AND U13597 ( .A(n776), .B(n13802), .Z(n13801) );
  XOR U13598 ( .A(n13803), .B(n13800), .Z(n13802) );
  XOR U13599 ( .A(n13804), .B(n13805), .Z(n13792) );
  AND U13600 ( .A(n13806), .B(n13807), .Z(n13805) );
  XOR U13601 ( .A(n13804), .B(n12045), .Z(n13807) );
  XOR U13602 ( .A(n13808), .B(n13809), .Z(n12045) );
  AND U13603 ( .A(n779), .B(n13810), .Z(n13809) );
  XOR U13604 ( .A(n13811), .B(n13808), .Z(n13810) );
  XNOR U13605 ( .A(n12042), .B(n13804), .Z(n13806) );
  XOR U13606 ( .A(n13812), .B(n13813), .Z(n12042) );
  AND U13607 ( .A(n776), .B(n13814), .Z(n13813) );
  XOR U13608 ( .A(n13815), .B(n13812), .Z(n13814) );
  XOR U13609 ( .A(n13816), .B(n13817), .Z(n13804) );
  AND U13610 ( .A(n13818), .B(n13819), .Z(n13817) );
  XOR U13611 ( .A(n13816), .B(n12057), .Z(n13819) );
  XOR U13612 ( .A(n13820), .B(n13821), .Z(n12057) );
  AND U13613 ( .A(n779), .B(n13822), .Z(n13821) );
  XOR U13614 ( .A(n13823), .B(n13820), .Z(n13822) );
  XNOR U13615 ( .A(n12054), .B(n13816), .Z(n13818) );
  XOR U13616 ( .A(n13824), .B(n13825), .Z(n12054) );
  AND U13617 ( .A(n776), .B(n13826), .Z(n13825) );
  XOR U13618 ( .A(n13827), .B(n13824), .Z(n13826) );
  XOR U13619 ( .A(n13828), .B(n13829), .Z(n13816) );
  AND U13620 ( .A(n13830), .B(n13831), .Z(n13829) );
  XNOR U13621 ( .A(n13832), .B(n12070), .Z(n13831) );
  XOR U13622 ( .A(n13833), .B(n13834), .Z(n12070) );
  AND U13623 ( .A(n779), .B(n13835), .Z(n13834) );
  XOR U13624 ( .A(n13833), .B(n13836), .Z(n13835) );
  XNOR U13625 ( .A(n12067), .B(n13828), .Z(n13830) );
  XOR U13626 ( .A(n13837), .B(n13838), .Z(n12067) );
  AND U13627 ( .A(n776), .B(n13839), .Z(n13838) );
  XOR U13628 ( .A(n13837), .B(n13840), .Z(n13839) );
  IV U13629 ( .A(n13832), .Z(n13828) );
  AND U13630 ( .A(n13659), .B(n13662), .Z(n13832) );
  XNOR U13631 ( .A(n13841), .B(n13842), .Z(n13662) );
  AND U13632 ( .A(n779), .B(n13843), .Z(n13842) );
  XNOR U13633 ( .A(n13844), .B(n13841), .Z(n13843) );
  XOR U13634 ( .A(n13845), .B(n13846), .Z(n779) );
  AND U13635 ( .A(n13847), .B(n13848), .Z(n13846) );
  XNOR U13636 ( .A(n13667), .B(n13845), .Z(n13848) );
  AND U13637 ( .A(n13849), .B(n13850), .Z(n13667) );
  XOR U13638 ( .A(n13845), .B(n13668), .Z(n13847) );
  AND U13639 ( .A(n13851), .B(n13852), .Z(n13668) );
  XOR U13640 ( .A(n13853), .B(n13854), .Z(n13845) );
  AND U13641 ( .A(n13855), .B(n13856), .Z(n13854) );
  XOR U13642 ( .A(n13853), .B(n13679), .Z(n13856) );
  XOR U13643 ( .A(n13857), .B(n13858), .Z(n13679) );
  AND U13644 ( .A(n459), .B(n13859), .Z(n13858) );
  XOR U13645 ( .A(n13860), .B(n13857), .Z(n13859) );
  XNOR U13646 ( .A(n13676), .B(n13853), .Z(n13855) );
  XOR U13647 ( .A(n13861), .B(n13862), .Z(n13676) );
  AND U13648 ( .A(n457), .B(n13863), .Z(n13862) );
  XOR U13649 ( .A(n13864), .B(n13861), .Z(n13863) );
  XOR U13650 ( .A(n13865), .B(n13866), .Z(n13853) );
  AND U13651 ( .A(n13867), .B(n13868), .Z(n13866) );
  XOR U13652 ( .A(n13865), .B(n13691), .Z(n13868) );
  XOR U13653 ( .A(n13869), .B(n13870), .Z(n13691) );
  AND U13654 ( .A(n459), .B(n13871), .Z(n13870) );
  XOR U13655 ( .A(n13872), .B(n13869), .Z(n13871) );
  XNOR U13656 ( .A(n13688), .B(n13865), .Z(n13867) );
  XOR U13657 ( .A(n13873), .B(n13874), .Z(n13688) );
  AND U13658 ( .A(n457), .B(n13875), .Z(n13874) );
  XOR U13659 ( .A(n13876), .B(n13873), .Z(n13875) );
  XOR U13660 ( .A(n13877), .B(n13878), .Z(n13865) );
  AND U13661 ( .A(n13879), .B(n13880), .Z(n13878) );
  XOR U13662 ( .A(n13877), .B(n13703), .Z(n13880) );
  XOR U13663 ( .A(n13881), .B(n13882), .Z(n13703) );
  AND U13664 ( .A(n459), .B(n13883), .Z(n13882) );
  XOR U13665 ( .A(n13884), .B(n13881), .Z(n13883) );
  XNOR U13666 ( .A(n13700), .B(n13877), .Z(n13879) );
  XOR U13667 ( .A(n13885), .B(n13886), .Z(n13700) );
  AND U13668 ( .A(n457), .B(n13887), .Z(n13886) );
  XOR U13669 ( .A(n13888), .B(n13885), .Z(n13887) );
  XOR U13670 ( .A(n13889), .B(n13890), .Z(n13877) );
  AND U13671 ( .A(n13891), .B(n13892), .Z(n13890) );
  XOR U13672 ( .A(n13889), .B(n13715), .Z(n13892) );
  XOR U13673 ( .A(n13893), .B(n13894), .Z(n13715) );
  AND U13674 ( .A(n459), .B(n13895), .Z(n13894) );
  XOR U13675 ( .A(n13896), .B(n13893), .Z(n13895) );
  XNOR U13676 ( .A(n13712), .B(n13889), .Z(n13891) );
  XOR U13677 ( .A(n13897), .B(n13898), .Z(n13712) );
  AND U13678 ( .A(n457), .B(n13899), .Z(n13898) );
  XOR U13679 ( .A(n13900), .B(n13897), .Z(n13899) );
  XOR U13680 ( .A(n13901), .B(n13902), .Z(n13889) );
  AND U13681 ( .A(n13903), .B(n13904), .Z(n13902) );
  XOR U13682 ( .A(n13901), .B(n13727), .Z(n13904) );
  XOR U13683 ( .A(n13905), .B(n13906), .Z(n13727) );
  AND U13684 ( .A(n459), .B(n13907), .Z(n13906) );
  XOR U13685 ( .A(n13908), .B(n13905), .Z(n13907) );
  XNOR U13686 ( .A(n13724), .B(n13901), .Z(n13903) );
  XOR U13687 ( .A(n13909), .B(n13910), .Z(n13724) );
  AND U13688 ( .A(n457), .B(n13911), .Z(n13910) );
  XOR U13689 ( .A(n13912), .B(n13909), .Z(n13911) );
  XOR U13690 ( .A(n13913), .B(n13914), .Z(n13901) );
  AND U13691 ( .A(n13915), .B(n13916), .Z(n13914) );
  XOR U13692 ( .A(n13913), .B(n13739), .Z(n13916) );
  XOR U13693 ( .A(n13917), .B(n13918), .Z(n13739) );
  AND U13694 ( .A(n459), .B(n13919), .Z(n13918) );
  XOR U13695 ( .A(n13920), .B(n13917), .Z(n13919) );
  XNOR U13696 ( .A(n13736), .B(n13913), .Z(n13915) );
  XOR U13697 ( .A(n13921), .B(n13922), .Z(n13736) );
  AND U13698 ( .A(n457), .B(n13923), .Z(n13922) );
  XOR U13699 ( .A(n13924), .B(n13921), .Z(n13923) );
  XOR U13700 ( .A(n13925), .B(n13926), .Z(n13913) );
  AND U13701 ( .A(n13927), .B(n13928), .Z(n13926) );
  XOR U13702 ( .A(n13925), .B(n13751), .Z(n13928) );
  XOR U13703 ( .A(n13929), .B(n13930), .Z(n13751) );
  AND U13704 ( .A(n459), .B(n13931), .Z(n13930) );
  XOR U13705 ( .A(n13932), .B(n13929), .Z(n13931) );
  XNOR U13706 ( .A(n13748), .B(n13925), .Z(n13927) );
  XOR U13707 ( .A(n13933), .B(n13934), .Z(n13748) );
  AND U13708 ( .A(n457), .B(n13935), .Z(n13934) );
  XOR U13709 ( .A(n13936), .B(n13933), .Z(n13935) );
  XOR U13710 ( .A(n13937), .B(n13938), .Z(n13925) );
  AND U13711 ( .A(n13939), .B(n13940), .Z(n13938) );
  XOR U13712 ( .A(n13937), .B(n13763), .Z(n13940) );
  XOR U13713 ( .A(n13941), .B(n13942), .Z(n13763) );
  AND U13714 ( .A(n459), .B(n13943), .Z(n13942) );
  XOR U13715 ( .A(n13944), .B(n13941), .Z(n13943) );
  XNOR U13716 ( .A(n13760), .B(n13937), .Z(n13939) );
  XOR U13717 ( .A(n13945), .B(n13946), .Z(n13760) );
  AND U13718 ( .A(n457), .B(n13947), .Z(n13946) );
  XOR U13719 ( .A(n13948), .B(n13945), .Z(n13947) );
  XOR U13720 ( .A(n13949), .B(n13950), .Z(n13937) );
  AND U13721 ( .A(n13951), .B(n13952), .Z(n13950) );
  XOR U13722 ( .A(n13949), .B(n13775), .Z(n13952) );
  XOR U13723 ( .A(n13953), .B(n13954), .Z(n13775) );
  AND U13724 ( .A(n459), .B(n13955), .Z(n13954) );
  XOR U13725 ( .A(n13956), .B(n13953), .Z(n13955) );
  XNOR U13726 ( .A(n13772), .B(n13949), .Z(n13951) );
  XOR U13727 ( .A(n13957), .B(n13958), .Z(n13772) );
  AND U13728 ( .A(n457), .B(n13959), .Z(n13958) );
  XOR U13729 ( .A(n13960), .B(n13957), .Z(n13959) );
  XOR U13730 ( .A(n13961), .B(n13962), .Z(n13949) );
  AND U13731 ( .A(n13963), .B(n13964), .Z(n13962) );
  XOR U13732 ( .A(n13961), .B(n13787), .Z(n13964) );
  XOR U13733 ( .A(n13965), .B(n13966), .Z(n13787) );
  AND U13734 ( .A(n459), .B(n13967), .Z(n13966) );
  XOR U13735 ( .A(n13968), .B(n13965), .Z(n13967) );
  XNOR U13736 ( .A(n13784), .B(n13961), .Z(n13963) );
  XOR U13737 ( .A(n13969), .B(n13970), .Z(n13784) );
  AND U13738 ( .A(n457), .B(n13971), .Z(n13970) );
  XOR U13739 ( .A(n13972), .B(n13969), .Z(n13971) );
  XOR U13740 ( .A(n13973), .B(n13974), .Z(n13961) );
  AND U13741 ( .A(n13975), .B(n13976), .Z(n13974) );
  XOR U13742 ( .A(n13973), .B(n13799), .Z(n13976) );
  XOR U13743 ( .A(n13977), .B(n13978), .Z(n13799) );
  AND U13744 ( .A(n459), .B(n13979), .Z(n13978) );
  XOR U13745 ( .A(n13980), .B(n13977), .Z(n13979) );
  XNOR U13746 ( .A(n13796), .B(n13973), .Z(n13975) );
  XOR U13747 ( .A(n13981), .B(n13982), .Z(n13796) );
  AND U13748 ( .A(n457), .B(n13983), .Z(n13982) );
  XOR U13749 ( .A(n13984), .B(n13981), .Z(n13983) );
  XOR U13750 ( .A(n13985), .B(n13986), .Z(n13973) );
  AND U13751 ( .A(n13987), .B(n13988), .Z(n13986) );
  XOR U13752 ( .A(n13985), .B(n13811), .Z(n13988) );
  XOR U13753 ( .A(n13989), .B(n13990), .Z(n13811) );
  AND U13754 ( .A(n459), .B(n13991), .Z(n13990) );
  XOR U13755 ( .A(n13992), .B(n13989), .Z(n13991) );
  XNOR U13756 ( .A(n13808), .B(n13985), .Z(n13987) );
  XOR U13757 ( .A(n13993), .B(n13994), .Z(n13808) );
  AND U13758 ( .A(n457), .B(n13995), .Z(n13994) );
  XOR U13759 ( .A(n13996), .B(n13993), .Z(n13995) );
  XOR U13760 ( .A(n13997), .B(n13998), .Z(n13985) );
  AND U13761 ( .A(n13999), .B(n14000), .Z(n13998) );
  XOR U13762 ( .A(n13997), .B(n13823), .Z(n14000) );
  XOR U13763 ( .A(n14001), .B(n14002), .Z(n13823) );
  AND U13764 ( .A(n459), .B(n14003), .Z(n14002) );
  XOR U13765 ( .A(n14004), .B(n14001), .Z(n14003) );
  XNOR U13766 ( .A(n13820), .B(n13997), .Z(n13999) );
  XOR U13767 ( .A(n14005), .B(n14006), .Z(n13820) );
  AND U13768 ( .A(n457), .B(n14007), .Z(n14006) );
  XOR U13769 ( .A(n14008), .B(n14005), .Z(n14007) );
  XOR U13770 ( .A(n14009), .B(n14010), .Z(n13997) );
  AND U13771 ( .A(n14011), .B(n14012), .Z(n14010) );
  XNOR U13772 ( .A(n14013), .B(n13836), .Z(n14012) );
  XOR U13773 ( .A(n14014), .B(n14015), .Z(n13836) );
  AND U13774 ( .A(n459), .B(n14016), .Z(n14015) );
  XOR U13775 ( .A(n14014), .B(n14017), .Z(n14016) );
  XNOR U13776 ( .A(n13833), .B(n14009), .Z(n14011) );
  XOR U13777 ( .A(n14018), .B(n14019), .Z(n13833) );
  AND U13778 ( .A(n457), .B(n14020), .Z(n14019) );
  XOR U13779 ( .A(n14018), .B(n14021), .Z(n14020) );
  IV U13780 ( .A(n14013), .Z(n14009) );
  AND U13781 ( .A(n13841), .B(n13844), .Z(n14013) );
  XNOR U13782 ( .A(n14022), .B(n14023), .Z(n13844) );
  AND U13783 ( .A(n459), .B(n14024), .Z(n14023) );
  XNOR U13784 ( .A(n14025), .B(n14022), .Z(n14024) );
  XOR U13785 ( .A(n14026), .B(n14027), .Z(n459) );
  AND U13786 ( .A(n14028), .B(n14029), .Z(n14027) );
  XNOR U13787 ( .A(n13849), .B(n14026), .Z(n14029) );
  AND U13788 ( .A(p_input[2303]), .B(p_input[2287]), .Z(n13849) );
  XOR U13789 ( .A(n14026), .B(n13850), .Z(n14028) );
  AND U13790 ( .A(p_input[2271]), .B(p_input[2255]), .Z(n13850) );
  XOR U13791 ( .A(n14030), .B(n14031), .Z(n14026) );
  AND U13792 ( .A(n14032), .B(n14033), .Z(n14031) );
  XOR U13793 ( .A(n14030), .B(n13860), .Z(n14033) );
  XNOR U13794 ( .A(p_input[2286]), .B(n14034), .Z(n13860) );
  AND U13795 ( .A(n319), .B(n14035), .Z(n14034) );
  XOR U13796 ( .A(p_input[2302]), .B(p_input[2286]), .Z(n14035) );
  XNOR U13797 ( .A(n13857), .B(n14030), .Z(n14032) );
  XOR U13798 ( .A(n14036), .B(n14037), .Z(n13857) );
  AND U13799 ( .A(n317), .B(n14038), .Z(n14037) );
  XOR U13800 ( .A(p_input[2270]), .B(p_input[2254]), .Z(n14038) );
  XOR U13801 ( .A(n14039), .B(n14040), .Z(n14030) );
  AND U13802 ( .A(n14041), .B(n14042), .Z(n14040) );
  XOR U13803 ( .A(n14039), .B(n13872), .Z(n14042) );
  XNOR U13804 ( .A(p_input[2285]), .B(n14043), .Z(n13872) );
  AND U13805 ( .A(n319), .B(n14044), .Z(n14043) );
  XOR U13806 ( .A(p_input[2301]), .B(p_input[2285]), .Z(n14044) );
  XNOR U13807 ( .A(n13869), .B(n14039), .Z(n14041) );
  XOR U13808 ( .A(n14045), .B(n14046), .Z(n13869) );
  AND U13809 ( .A(n317), .B(n14047), .Z(n14046) );
  XOR U13810 ( .A(p_input[2269]), .B(p_input[2253]), .Z(n14047) );
  XOR U13811 ( .A(n14048), .B(n14049), .Z(n14039) );
  AND U13812 ( .A(n14050), .B(n14051), .Z(n14049) );
  XOR U13813 ( .A(n14048), .B(n13884), .Z(n14051) );
  XNOR U13814 ( .A(p_input[2284]), .B(n14052), .Z(n13884) );
  AND U13815 ( .A(n319), .B(n14053), .Z(n14052) );
  XOR U13816 ( .A(p_input[2300]), .B(p_input[2284]), .Z(n14053) );
  XNOR U13817 ( .A(n13881), .B(n14048), .Z(n14050) );
  XOR U13818 ( .A(n14054), .B(n14055), .Z(n13881) );
  AND U13819 ( .A(n317), .B(n14056), .Z(n14055) );
  XOR U13820 ( .A(p_input[2268]), .B(p_input[2252]), .Z(n14056) );
  XOR U13821 ( .A(n14057), .B(n14058), .Z(n14048) );
  AND U13822 ( .A(n14059), .B(n14060), .Z(n14058) );
  XOR U13823 ( .A(n14057), .B(n13896), .Z(n14060) );
  XNOR U13824 ( .A(p_input[2283]), .B(n14061), .Z(n13896) );
  AND U13825 ( .A(n319), .B(n14062), .Z(n14061) );
  XOR U13826 ( .A(p_input[2299]), .B(p_input[2283]), .Z(n14062) );
  XNOR U13827 ( .A(n13893), .B(n14057), .Z(n14059) );
  XOR U13828 ( .A(n14063), .B(n14064), .Z(n13893) );
  AND U13829 ( .A(n317), .B(n14065), .Z(n14064) );
  XOR U13830 ( .A(p_input[2267]), .B(p_input[2251]), .Z(n14065) );
  XOR U13831 ( .A(n14066), .B(n14067), .Z(n14057) );
  AND U13832 ( .A(n14068), .B(n14069), .Z(n14067) );
  XOR U13833 ( .A(n14066), .B(n13908), .Z(n14069) );
  XNOR U13834 ( .A(p_input[2282]), .B(n14070), .Z(n13908) );
  AND U13835 ( .A(n319), .B(n14071), .Z(n14070) );
  XOR U13836 ( .A(p_input[2298]), .B(p_input[2282]), .Z(n14071) );
  XNOR U13837 ( .A(n13905), .B(n14066), .Z(n14068) );
  XOR U13838 ( .A(n14072), .B(n14073), .Z(n13905) );
  AND U13839 ( .A(n317), .B(n14074), .Z(n14073) );
  XOR U13840 ( .A(p_input[2266]), .B(p_input[2250]), .Z(n14074) );
  XOR U13841 ( .A(n14075), .B(n14076), .Z(n14066) );
  AND U13842 ( .A(n14077), .B(n14078), .Z(n14076) );
  XOR U13843 ( .A(n14075), .B(n13920), .Z(n14078) );
  XNOR U13844 ( .A(p_input[2281]), .B(n14079), .Z(n13920) );
  AND U13845 ( .A(n319), .B(n14080), .Z(n14079) );
  XOR U13846 ( .A(p_input[2297]), .B(p_input[2281]), .Z(n14080) );
  XNOR U13847 ( .A(n13917), .B(n14075), .Z(n14077) );
  XOR U13848 ( .A(n14081), .B(n14082), .Z(n13917) );
  AND U13849 ( .A(n317), .B(n14083), .Z(n14082) );
  XOR U13850 ( .A(p_input[2265]), .B(p_input[2249]), .Z(n14083) );
  XOR U13851 ( .A(n14084), .B(n14085), .Z(n14075) );
  AND U13852 ( .A(n14086), .B(n14087), .Z(n14085) );
  XOR U13853 ( .A(n14084), .B(n13932), .Z(n14087) );
  XNOR U13854 ( .A(p_input[2280]), .B(n14088), .Z(n13932) );
  AND U13855 ( .A(n319), .B(n14089), .Z(n14088) );
  XOR U13856 ( .A(p_input[2296]), .B(p_input[2280]), .Z(n14089) );
  XNOR U13857 ( .A(n13929), .B(n14084), .Z(n14086) );
  XOR U13858 ( .A(n14090), .B(n14091), .Z(n13929) );
  AND U13859 ( .A(n317), .B(n14092), .Z(n14091) );
  XOR U13860 ( .A(p_input[2264]), .B(p_input[2248]), .Z(n14092) );
  XOR U13861 ( .A(n14093), .B(n14094), .Z(n14084) );
  AND U13862 ( .A(n14095), .B(n14096), .Z(n14094) );
  XOR U13863 ( .A(n14093), .B(n13944), .Z(n14096) );
  XNOR U13864 ( .A(p_input[2279]), .B(n14097), .Z(n13944) );
  AND U13865 ( .A(n319), .B(n14098), .Z(n14097) );
  XOR U13866 ( .A(p_input[2295]), .B(p_input[2279]), .Z(n14098) );
  XNOR U13867 ( .A(n13941), .B(n14093), .Z(n14095) );
  XOR U13868 ( .A(n14099), .B(n14100), .Z(n13941) );
  AND U13869 ( .A(n317), .B(n14101), .Z(n14100) );
  XOR U13870 ( .A(p_input[2263]), .B(p_input[2247]), .Z(n14101) );
  XOR U13871 ( .A(n14102), .B(n14103), .Z(n14093) );
  AND U13872 ( .A(n14104), .B(n14105), .Z(n14103) );
  XOR U13873 ( .A(n14102), .B(n13956), .Z(n14105) );
  XNOR U13874 ( .A(p_input[2278]), .B(n14106), .Z(n13956) );
  AND U13875 ( .A(n319), .B(n14107), .Z(n14106) );
  XOR U13876 ( .A(p_input[2294]), .B(p_input[2278]), .Z(n14107) );
  XNOR U13877 ( .A(n13953), .B(n14102), .Z(n14104) );
  XOR U13878 ( .A(n14108), .B(n14109), .Z(n13953) );
  AND U13879 ( .A(n317), .B(n14110), .Z(n14109) );
  XOR U13880 ( .A(p_input[2262]), .B(p_input[2246]), .Z(n14110) );
  XOR U13881 ( .A(n14111), .B(n14112), .Z(n14102) );
  AND U13882 ( .A(n14113), .B(n14114), .Z(n14112) );
  XOR U13883 ( .A(n14111), .B(n13968), .Z(n14114) );
  XNOR U13884 ( .A(p_input[2277]), .B(n14115), .Z(n13968) );
  AND U13885 ( .A(n319), .B(n14116), .Z(n14115) );
  XOR U13886 ( .A(p_input[2293]), .B(p_input[2277]), .Z(n14116) );
  XNOR U13887 ( .A(n13965), .B(n14111), .Z(n14113) );
  XOR U13888 ( .A(n14117), .B(n14118), .Z(n13965) );
  AND U13889 ( .A(n317), .B(n14119), .Z(n14118) );
  XOR U13890 ( .A(p_input[2261]), .B(p_input[2245]), .Z(n14119) );
  XOR U13891 ( .A(n14120), .B(n14121), .Z(n14111) );
  AND U13892 ( .A(n14122), .B(n14123), .Z(n14121) );
  XOR U13893 ( .A(n14120), .B(n13980), .Z(n14123) );
  XNOR U13894 ( .A(p_input[2276]), .B(n14124), .Z(n13980) );
  AND U13895 ( .A(n319), .B(n14125), .Z(n14124) );
  XOR U13896 ( .A(p_input[2292]), .B(p_input[2276]), .Z(n14125) );
  XNOR U13897 ( .A(n13977), .B(n14120), .Z(n14122) );
  XOR U13898 ( .A(n14126), .B(n14127), .Z(n13977) );
  AND U13899 ( .A(n317), .B(n14128), .Z(n14127) );
  XOR U13900 ( .A(p_input[2260]), .B(p_input[2244]), .Z(n14128) );
  XOR U13901 ( .A(n14129), .B(n14130), .Z(n14120) );
  AND U13902 ( .A(n14131), .B(n14132), .Z(n14130) );
  XOR U13903 ( .A(n14129), .B(n13992), .Z(n14132) );
  XNOR U13904 ( .A(p_input[2275]), .B(n14133), .Z(n13992) );
  AND U13905 ( .A(n319), .B(n14134), .Z(n14133) );
  XOR U13906 ( .A(p_input[2291]), .B(p_input[2275]), .Z(n14134) );
  XNOR U13907 ( .A(n13989), .B(n14129), .Z(n14131) );
  XOR U13908 ( .A(n14135), .B(n14136), .Z(n13989) );
  AND U13909 ( .A(n317), .B(n14137), .Z(n14136) );
  XOR U13910 ( .A(p_input[2259]), .B(p_input[2243]), .Z(n14137) );
  XOR U13911 ( .A(n14138), .B(n14139), .Z(n14129) );
  AND U13912 ( .A(n14140), .B(n14141), .Z(n14139) );
  XOR U13913 ( .A(n14138), .B(n14004), .Z(n14141) );
  XNOR U13914 ( .A(p_input[2274]), .B(n14142), .Z(n14004) );
  AND U13915 ( .A(n319), .B(n14143), .Z(n14142) );
  XOR U13916 ( .A(p_input[2290]), .B(p_input[2274]), .Z(n14143) );
  XNOR U13917 ( .A(n14001), .B(n14138), .Z(n14140) );
  XOR U13918 ( .A(n14144), .B(n14145), .Z(n14001) );
  AND U13919 ( .A(n317), .B(n14146), .Z(n14145) );
  XOR U13920 ( .A(p_input[2258]), .B(p_input[2242]), .Z(n14146) );
  XOR U13921 ( .A(n14147), .B(n14148), .Z(n14138) );
  AND U13922 ( .A(n14149), .B(n14150), .Z(n14148) );
  XNOR U13923 ( .A(n14151), .B(n14017), .Z(n14150) );
  XNOR U13924 ( .A(p_input[2273]), .B(n14152), .Z(n14017) );
  AND U13925 ( .A(n319), .B(n14153), .Z(n14152) );
  XNOR U13926 ( .A(p_input[2289]), .B(n14154), .Z(n14153) );
  IV U13927 ( .A(p_input[2273]), .Z(n14154) );
  XNOR U13928 ( .A(n14014), .B(n14147), .Z(n14149) );
  XNOR U13929 ( .A(p_input[2241]), .B(n14155), .Z(n14014) );
  AND U13930 ( .A(n317), .B(n14156), .Z(n14155) );
  XOR U13931 ( .A(p_input[2257]), .B(p_input[2241]), .Z(n14156) );
  IV U13932 ( .A(n14151), .Z(n14147) );
  AND U13933 ( .A(n14022), .B(n14025), .Z(n14151) );
  XOR U13934 ( .A(p_input[2272]), .B(n14157), .Z(n14025) );
  AND U13935 ( .A(n319), .B(n14158), .Z(n14157) );
  XOR U13936 ( .A(p_input[2288]), .B(p_input[2272]), .Z(n14158) );
  XOR U13937 ( .A(n14159), .B(n14160), .Z(n319) );
  AND U13938 ( .A(n14161), .B(n14162), .Z(n14160) );
  XNOR U13939 ( .A(p_input[2303]), .B(n14159), .Z(n14162) );
  XOR U13940 ( .A(n14159), .B(p_input[2287]), .Z(n14161) );
  XOR U13941 ( .A(n14163), .B(n14164), .Z(n14159) );
  AND U13942 ( .A(n14165), .B(n14166), .Z(n14164) );
  XNOR U13943 ( .A(p_input[2302]), .B(n14163), .Z(n14166) );
  XOR U13944 ( .A(n14163), .B(p_input[2286]), .Z(n14165) );
  XOR U13945 ( .A(n14167), .B(n14168), .Z(n14163) );
  AND U13946 ( .A(n14169), .B(n14170), .Z(n14168) );
  XNOR U13947 ( .A(p_input[2301]), .B(n14167), .Z(n14170) );
  XOR U13948 ( .A(n14167), .B(p_input[2285]), .Z(n14169) );
  XOR U13949 ( .A(n14171), .B(n14172), .Z(n14167) );
  AND U13950 ( .A(n14173), .B(n14174), .Z(n14172) );
  XNOR U13951 ( .A(p_input[2300]), .B(n14171), .Z(n14174) );
  XOR U13952 ( .A(n14171), .B(p_input[2284]), .Z(n14173) );
  XOR U13953 ( .A(n14175), .B(n14176), .Z(n14171) );
  AND U13954 ( .A(n14177), .B(n14178), .Z(n14176) );
  XNOR U13955 ( .A(p_input[2299]), .B(n14175), .Z(n14178) );
  XOR U13956 ( .A(n14175), .B(p_input[2283]), .Z(n14177) );
  XOR U13957 ( .A(n14179), .B(n14180), .Z(n14175) );
  AND U13958 ( .A(n14181), .B(n14182), .Z(n14180) );
  XNOR U13959 ( .A(p_input[2298]), .B(n14179), .Z(n14182) );
  XOR U13960 ( .A(n14179), .B(p_input[2282]), .Z(n14181) );
  XOR U13961 ( .A(n14183), .B(n14184), .Z(n14179) );
  AND U13962 ( .A(n14185), .B(n14186), .Z(n14184) );
  XNOR U13963 ( .A(p_input[2297]), .B(n14183), .Z(n14186) );
  XOR U13964 ( .A(n14183), .B(p_input[2281]), .Z(n14185) );
  XOR U13965 ( .A(n14187), .B(n14188), .Z(n14183) );
  AND U13966 ( .A(n14189), .B(n14190), .Z(n14188) );
  XNOR U13967 ( .A(p_input[2296]), .B(n14187), .Z(n14190) );
  XOR U13968 ( .A(n14187), .B(p_input[2280]), .Z(n14189) );
  XOR U13969 ( .A(n14191), .B(n14192), .Z(n14187) );
  AND U13970 ( .A(n14193), .B(n14194), .Z(n14192) );
  XNOR U13971 ( .A(p_input[2295]), .B(n14191), .Z(n14194) );
  XOR U13972 ( .A(n14191), .B(p_input[2279]), .Z(n14193) );
  XOR U13973 ( .A(n14195), .B(n14196), .Z(n14191) );
  AND U13974 ( .A(n14197), .B(n14198), .Z(n14196) );
  XNOR U13975 ( .A(p_input[2294]), .B(n14195), .Z(n14198) );
  XOR U13976 ( .A(n14195), .B(p_input[2278]), .Z(n14197) );
  XOR U13977 ( .A(n14199), .B(n14200), .Z(n14195) );
  AND U13978 ( .A(n14201), .B(n14202), .Z(n14200) );
  XNOR U13979 ( .A(p_input[2293]), .B(n14199), .Z(n14202) );
  XOR U13980 ( .A(n14199), .B(p_input[2277]), .Z(n14201) );
  XOR U13981 ( .A(n14203), .B(n14204), .Z(n14199) );
  AND U13982 ( .A(n14205), .B(n14206), .Z(n14204) );
  XNOR U13983 ( .A(p_input[2292]), .B(n14203), .Z(n14206) );
  XOR U13984 ( .A(n14203), .B(p_input[2276]), .Z(n14205) );
  XOR U13985 ( .A(n14207), .B(n14208), .Z(n14203) );
  AND U13986 ( .A(n14209), .B(n14210), .Z(n14208) );
  XNOR U13987 ( .A(p_input[2291]), .B(n14207), .Z(n14210) );
  XOR U13988 ( .A(n14207), .B(p_input[2275]), .Z(n14209) );
  XOR U13989 ( .A(n14211), .B(n14212), .Z(n14207) );
  AND U13990 ( .A(n14213), .B(n14214), .Z(n14212) );
  XNOR U13991 ( .A(p_input[2290]), .B(n14211), .Z(n14214) );
  XOR U13992 ( .A(n14211), .B(p_input[2274]), .Z(n14213) );
  XNOR U13993 ( .A(n14215), .B(n14216), .Z(n14211) );
  AND U13994 ( .A(n14217), .B(n14218), .Z(n14216) );
  XOR U13995 ( .A(p_input[2289]), .B(n14215), .Z(n14218) );
  XNOR U13996 ( .A(p_input[2273]), .B(n14215), .Z(n14217) );
  AND U13997 ( .A(p_input[2288]), .B(n14219), .Z(n14215) );
  IV U13998 ( .A(p_input[2272]), .Z(n14219) );
  XNOR U13999 ( .A(p_input[2240]), .B(n14220), .Z(n14022) );
  AND U14000 ( .A(n317), .B(n14221), .Z(n14220) );
  XOR U14001 ( .A(p_input[2256]), .B(p_input[2240]), .Z(n14221) );
  XOR U14002 ( .A(n14222), .B(n14223), .Z(n317) );
  AND U14003 ( .A(n14224), .B(n14225), .Z(n14223) );
  XNOR U14004 ( .A(p_input[2271]), .B(n14222), .Z(n14225) );
  XOR U14005 ( .A(n14222), .B(p_input[2255]), .Z(n14224) );
  XOR U14006 ( .A(n14226), .B(n14227), .Z(n14222) );
  AND U14007 ( .A(n14228), .B(n14229), .Z(n14227) );
  XNOR U14008 ( .A(p_input[2270]), .B(n14226), .Z(n14229) );
  XNOR U14009 ( .A(n14226), .B(n14036), .Z(n14228) );
  IV U14010 ( .A(p_input[2254]), .Z(n14036) );
  XOR U14011 ( .A(n14230), .B(n14231), .Z(n14226) );
  AND U14012 ( .A(n14232), .B(n14233), .Z(n14231) );
  XNOR U14013 ( .A(p_input[2269]), .B(n14230), .Z(n14233) );
  XNOR U14014 ( .A(n14230), .B(n14045), .Z(n14232) );
  IV U14015 ( .A(p_input[2253]), .Z(n14045) );
  XOR U14016 ( .A(n14234), .B(n14235), .Z(n14230) );
  AND U14017 ( .A(n14236), .B(n14237), .Z(n14235) );
  XNOR U14018 ( .A(p_input[2268]), .B(n14234), .Z(n14237) );
  XNOR U14019 ( .A(n14234), .B(n14054), .Z(n14236) );
  IV U14020 ( .A(p_input[2252]), .Z(n14054) );
  XOR U14021 ( .A(n14238), .B(n14239), .Z(n14234) );
  AND U14022 ( .A(n14240), .B(n14241), .Z(n14239) );
  XNOR U14023 ( .A(p_input[2267]), .B(n14238), .Z(n14241) );
  XNOR U14024 ( .A(n14238), .B(n14063), .Z(n14240) );
  IV U14025 ( .A(p_input[2251]), .Z(n14063) );
  XOR U14026 ( .A(n14242), .B(n14243), .Z(n14238) );
  AND U14027 ( .A(n14244), .B(n14245), .Z(n14243) );
  XNOR U14028 ( .A(p_input[2266]), .B(n14242), .Z(n14245) );
  XNOR U14029 ( .A(n14242), .B(n14072), .Z(n14244) );
  IV U14030 ( .A(p_input[2250]), .Z(n14072) );
  XOR U14031 ( .A(n14246), .B(n14247), .Z(n14242) );
  AND U14032 ( .A(n14248), .B(n14249), .Z(n14247) );
  XNOR U14033 ( .A(p_input[2265]), .B(n14246), .Z(n14249) );
  XNOR U14034 ( .A(n14246), .B(n14081), .Z(n14248) );
  IV U14035 ( .A(p_input[2249]), .Z(n14081) );
  XOR U14036 ( .A(n14250), .B(n14251), .Z(n14246) );
  AND U14037 ( .A(n14252), .B(n14253), .Z(n14251) );
  XNOR U14038 ( .A(p_input[2264]), .B(n14250), .Z(n14253) );
  XNOR U14039 ( .A(n14250), .B(n14090), .Z(n14252) );
  IV U14040 ( .A(p_input[2248]), .Z(n14090) );
  XOR U14041 ( .A(n14254), .B(n14255), .Z(n14250) );
  AND U14042 ( .A(n14256), .B(n14257), .Z(n14255) );
  XNOR U14043 ( .A(p_input[2263]), .B(n14254), .Z(n14257) );
  XNOR U14044 ( .A(n14254), .B(n14099), .Z(n14256) );
  IV U14045 ( .A(p_input[2247]), .Z(n14099) );
  XOR U14046 ( .A(n14258), .B(n14259), .Z(n14254) );
  AND U14047 ( .A(n14260), .B(n14261), .Z(n14259) );
  XNOR U14048 ( .A(p_input[2262]), .B(n14258), .Z(n14261) );
  XNOR U14049 ( .A(n14258), .B(n14108), .Z(n14260) );
  IV U14050 ( .A(p_input[2246]), .Z(n14108) );
  XOR U14051 ( .A(n14262), .B(n14263), .Z(n14258) );
  AND U14052 ( .A(n14264), .B(n14265), .Z(n14263) );
  XNOR U14053 ( .A(p_input[2261]), .B(n14262), .Z(n14265) );
  XNOR U14054 ( .A(n14262), .B(n14117), .Z(n14264) );
  IV U14055 ( .A(p_input[2245]), .Z(n14117) );
  XOR U14056 ( .A(n14266), .B(n14267), .Z(n14262) );
  AND U14057 ( .A(n14268), .B(n14269), .Z(n14267) );
  XNOR U14058 ( .A(p_input[2260]), .B(n14266), .Z(n14269) );
  XNOR U14059 ( .A(n14266), .B(n14126), .Z(n14268) );
  IV U14060 ( .A(p_input[2244]), .Z(n14126) );
  XOR U14061 ( .A(n14270), .B(n14271), .Z(n14266) );
  AND U14062 ( .A(n14272), .B(n14273), .Z(n14271) );
  XNOR U14063 ( .A(p_input[2259]), .B(n14270), .Z(n14273) );
  XNOR U14064 ( .A(n14270), .B(n14135), .Z(n14272) );
  IV U14065 ( .A(p_input[2243]), .Z(n14135) );
  XOR U14066 ( .A(n14274), .B(n14275), .Z(n14270) );
  AND U14067 ( .A(n14276), .B(n14277), .Z(n14275) );
  XNOR U14068 ( .A(p_input[2258]), .B(n14274), .Z(n14277) );
  XNOR U14069 ( .A(n14274), .B(n14144), .Z(n14276) );
  IV U14070 ( .A(p_input[2242]), .Z(n14144) );
  XNOR U14071 ( .A(n14278), .B(n14279), .Z(n14274) );
  AND U14072 ( .A(n14280), .B(n14281), .Z(n14279) );
  XOR U14073 ( .A(p_input[2257]), .B(n14278), .Z(n14281) );
  XNOR U14074 ( .A(p_input[2241]), .B(n14278), .Z(n14280) );
  AND U14075 ( .A(p_input[2256]), .B(n14282), .Z(n14278) );
  IV U14076 ( .A(p_input[2240]), .Z(n14282) );
  XOR U14077 ( .A(n14283), .B(n14284), .Z(n13841) );
  AND U14078 ( .A(n457), .B(n14285), .Z(n14284) );
  XNOR U14079 ( .A(n14286), .B(n14283), .Z(n14285) );
  XOR U14080 ( .A(n14287), .B(n14288), .Z(n457) );
  AND U14081 ( .A(n14289), .B(n14290), .Z(n14288) );
  XNOR U14082 ( .A(n13851), .B(n14287), .Z(n14290) );
  AND U14083 ( .A(p_input[2239]), .B(p_input[2223]), .Z(n13851) );
  XOR U14084 ( .A(n14287), .B(n13852), .Z(n14289) );
  AND U14085 ( .A(p_input[2207]), .B(p_input[2191]), .Z(n13852) );
  XOR U14086 ( .A(n14291), .B(n14292), .Z(n14287) );
  AND U14087 ( .A(n14293), .B(n14294), .Z(n14292) );
  XOR U14088 ( .A(n14291), .B(n13864), .Z(n14294) );
  XNOR U14089 ( .A(p_input[2222]), .B(n14295), .Z(n13864) );
  AND U14090 ( .A(n323), .B(n14296), .Z(n14295) );
  XOR U14091 ( .A(p_input[2238]), .B(p_input[2222]), .Z(n14296) );
  XNOR U14092 ( .A(n13861), .B(n14291), .Z(n14293) );
  XOR U14093 ( .A(n14297), .B(n14298), .Z(n13861) );
  AND U14094 ( .A(n320), .B(n14299), .Z(n14298) );
  XOR U14095 ( .A(p_input[2206]), .B(p_input[2190]), .Z(n14299) );
  XOR U14096 ( .A(n14300), .B(n14301), .Z(n14291) );
  AND U14097 ( .A(n14302), .B(n14303), .Z(n14301) );
  XOR U14098 ( .A(n14300), .B(n13876), .Z(n14303) );
  XNOR U14099 ( .A(p_input[2221]), .B(n14304), .Z(n13876) );
  AND U14100 ( .A(n323), .B(n14305), .Z(n14304) );
  XOR U14101 ( .A(p_input[2237]), .B(p_input[2221]), .Z(n14305) );
  XNOR U14102 ( .A(n13873), .B(n14300), .Z(n14302) );
  XOR U14103 ( .A(n14306), .B(n14307), .Z(n13873) );
  AND U14104 ( .A(n320), .B(n14308), .Z(n14307) );
  XOR U14105 ( .A(p_input[2205]), .B(p_input[2189]), .Z(n14308) );
  XOR U14106 ( .A(n14309), .B(n14310), .Z(n14300) );
  AND U14107 ( .A(n14311), .B(n14312), .Z(n14310) );
  XOR U14108 ( .A(n14309), .B(n13888), .Z(n14312) );
  XNOR U14109 ( .A(p_input[2220]), .B(n14313), .Z(n13888) );
  AND U14110 ( .A(n323), .B(n14314), .Z(n14313) );
  XOR U14111 ( .A(p_input[2236]), .B(p_input[2220]), .Z(n14314) );
  XNOR U14112 ( .A(n13885), .B(n14309), .Z(n14311) );
  XOR U14113 ( .A(n14315), .B(n14316), .Z(n13885) );
  AND U14114 ( .A(n320), .B(n14317), .Z(n14316) );
  XOR U14115 ( .A(p_input[2204]), .B(p_input[2188]), .Z(n14317) );
  XOR U14116 ( .A(n14318), .B(n14319), .Z(n14309) );
  AND U14117 ( .A(n14320), .B(n14321), .Z(n14319) );
  XOR U14118 ( .A(n14318), .B(n13900), .Z(n14321) );
  XNOR U14119 ( .A(p_input[2219]), .B(n14322), .Z(n13900) );
  AND U14120 ( .A(n323), .B(n14323), .Z(n14322) );
  XOR U14121 ( .A(p_input[2235]), .B(p_input[2219]), .Z(n14323) );
  XNOR U14122 ( .A(n13897), .B(n14318), .Z(n14320) );
  XOR U14123 ( .A(n14324), .B(n14325), .Z(n13897) );
  AND U14124 ( .A(n320), .B(n14326), .Z(n14325) );
  XOR U14125 ( .A(p_input[2203]), .B(p_input[2187]), .Z(n14326) );
  XOR U14126 ( .A(n14327), .B(n14328), .Z(n14318) );
  AND U14127 ( .A(n14329), .B(n14330), .Z(n14328) );
  XOR U14128 ( .A(n14327), .B(n13912), .Z(n14330) );
  XNOR U14129 ( .A(p_input[2218]), .B(n14331), .Z(n13912) );
  AND U14130 ( .A(n323), .B(n14332), .Z(n14331) );
  XOR U14131 ( .A(p_input[2234]), .B(p_input[2218]), .Z(n14332) );
  XNOR U14132 ( .A(n13909), .B(n14327), .Z(n14329) );
  XOR U14133 ( .A(n14333), .B(n14334), .Z(n13909) );
  AND U14134 ( .A(n320), .B(n14335), .Z(n14334) );
  XOR U14135 ( .A(p_input[2202]), .B(p_input[2186]), .Z(n14335) );
  XOR U14136 ( .A(n14336), .B(n14337), .Z(n14327) );
  AND U14137 ( .A(n14338), .B(n14339), .Z(n14337) );
  XOR U14138 ( .A(n14336), .B(n13924), .Z(n14339) );
  XNOR U14139 ( .A(p_input[2217]), .B(n14340), .Z(n13924) );
  AND U14140 ( .A(n323), .B(n14341), .Z(n14340) );
  XOR U14141 ( .A(p_input[2233]), .B(p_input[2217]), .Z(n14341) );
  XNOR U14142 ( .A(n13921), .B(n14336), .Z(n14338) );
  XOR U14143 ( .A(n14342), .B(n14343), .Z(n13921) );
  AND U14144 ( .A(n320), .B(n14344), .Z(n14343) );
  XOR U14145 ( .A(p_input[2201]), .B(p_input[2185]), .Z(n14344) );
  XOR U14146 ( .A(n14345), .B(n14346), .Z(n14336) );
  AND U14147 ( .A(n14347), .B(n14348), .Z(n14346) );
  XOR U14148 ( .A(n14345), .B(n13936), .Z(n14348) );
  XNOR U14149 ( .A(p_input[2216]), .B(n14349), .Z(n13936) );
  AND U14150 ( .A(n323), .B(n14350), .Z(n14349) );
  XOR U14151 ( .A(p_input[2232]), .B(p_input[2216]), .Z(n14350) );
  XNOR U14152 ( .A(n13933), .B(n14345), .Z(n14347) );
  XOR U14153 ( .A(n14351), .B(n14352), .Z(n13933) );
  AND U14154 ( .A(n320), .B(n14353), .Z(n14352) );
  XOR U14155 ( .A(p_input[2200]), .B(p_input[2184]), .Z(n14353) );
  XOR U14156 ( .A(n14354), .B(n14355), .Z(n14345) );
  AND U14157 ( .A(n14356), .B(n14357), .Z(n14355) );
  XOR U14158 ( .A(n14354), .B(n13948), .Z(n14357) );
  XNOR U14159 ( .A(p_input[2215]), .B(n14358), .Z(n13948) );
  AND U14160 ( .A(n323), .B(n14359), .Z(n14358) );
  XOR U14161 ( .A(p_input[2231]), .B(p_input[2215]), .Z(n14359) );
  XNOR U14162 ( .A(n13945), .B(n14354), .Z(n14356) );
  XOR U14163 ( .A(n14360), .B(n14361), .Z(n13945) );
  AND U14164 ( .A(n320), .B(n14362), .Z(n14361) );
  XOR U14165 ( .A(p_input[2199]), .B(p_input[2183]), .Z(n14362) );
  XOR U14166 ( .A(n14363), .B(n14364), .Z(n14354) );
  AND U14167 ( .A(n14365), .B(n14366), .Z(n14364) );
  XOR U14168 ( .A(n14363), .B(n13960), .Z(n14366) );
  XNOR U14169 ( .A(p_input[2214]), .B(n14367), .Z(n13960) );
  AND U14170 ( .A(n323), .B(n14368), .Z(n14367) );
  XOR U14171 ( .A(p_input[2230]), .B(p_input[2214]), .Z(n14368) );
  XNOR U14172 ( .A(n13957), .B(n14363), .Z(n14365) );
  XOR U14173 ( .A(n14369), .B(n14370), .Z(n13957) );
  AND U14174 ( .A(n320), .B(n14371), .Z(n14370) );
  XOR U14175 ( .A(p_input[2198]), .B(p_input[2182]), .Z(n14371) );
  XOR U14176 ( .A(n14372), .B(n14373), .Z(n14363) );
  AND U14177 ( .A(n14374), .B(n14375), .Z(n14373) );
  XOR U14178 ( .A(n14372), .B(n13972), .Z(n14375) );
  XNOR U14179 ( .A(p_input[2213]), .B(n14376), .Z(n13972) );
  AND U14180 ( .A(n323), .B(n14377), .Z(n14376) );
  XOR U14181 ( .A(p_input[2229]), .B(p_input[2213]), .Z(n14377) );
  XNOR U14182 ( .A(n13969), .B(n14372), .Z(n14374) );
  XOR U14183 ( .A(n14378), .B(n14379), .Z(n13969) );
  AND U14184 ( .A(n320), .B(n14380), .Z(n14379) );
  XOR U14185 ( .A(p_input[2197]), .B(p_input[2181]), .Z(n14380) );
  XOR U14186 ( .A(n14381), .B(n14382), .Z(n14372) );
  AND U14187 ( .A(n14383), .B(n14384), .Z(n14382) );
  XOR U14188 ( .A(n14381), .B(n13984), .Z(n14384) );
  XNOR U14189 ( .A(p_input[2212]), .B(n14385), .Z(n13984) );
  AND U14190 ( .A(n323), .B(n14386), .Z(n14385) );
  XOR U14191 ( .A(p_input[2228]), .B(p_input[2212]), .Z(n14386) );
  XNOR U14192 ( .A(n13981), .B(n14381), .Z(n14383) );
  XOR U14193 ( .A(n14387), .B(n14388), .Z(n13981) );
  AND U14194 ( .A(n320), .B(n14389), .Z(n14388) );
  XOR U14195 ( .A(p_input[2196]), .B(p_input[2180]), .Z(n14389) );
  XOR U14196 ( .A(n14390), .B(n14391), .Z(n14381) );
  AND U14197 ( .A(n14392), .B(n14393), .Z(n14391) );
  XOR U14198 ( .A(n14390), .B(n13996), .Z(n14393) );
  XNOR U14199 ( .A(p_input[2211]), .B(n14394), .Z(n13996) );
  AND U14200 ( .A(n323), .B(n14395), .Z(n14394) );
  XOR U14201 ( .A(p_input[2227]), .B(p_input[2211]), .Z(n14395) );
  XNOR U14202 ( .A(n13993), .B(n14390), .Z(n14392) );
  XOR U14203 ( .A(n14396), .B(n14397), .Z(n13993) );
  AND U14204 ( .A(n320), .B(n14398), .Z(n14397) );
  XOR U14205 ( .A(p_input[2195]), .B(p_input[2179]), .Z(n14398) );
  XOR U14206 ( .A(n14399), .B(n14400), .Z(n14390) );
  AND U14207 ( .A(n14401), .B(n14402), .Z(n14400) );
  XOR U14208 ( .A(n14399), .B(n14008), .Z(n14402) );
  XNOR U14209 ( .A(p_input[2210]), .B(n14403), .Z(n14008) );
  AND U14210 ( .A(n323), .B(n14404), .Z(n14403) );
  XOR U14211 ( .A(p_input[2226]), .B(p_input[2210]), .Z(n14404) );
  XNOR U14212 ( .A(n14005), .B(n14399), .Z(n14401) );
  XOR U14213 ( .A(n14405), .B(n14406), .Z(n14005) );
  AND U14214 ( .A(n320), .B(n14407), .Z(n14406) );
  XOR U14215 ( .A(p_input[2194]), .B(p_input[2178]), .Z(n14407) );
  XOR U14216 ( .A(n14408), .B(n14409), .Z(n14399) );
  AND U14217 ( .A(n14410), .B(n14411), .Z(n14409) );
  XNOR U14218 ( .A(n14412), .B(n14021), .Z(n14411) );
  XNOR U14219 ( .A(p_input[2209]), .B(n14413), .Z(n14021) );
  AND U14220 ( .A(n323), .B(n14414), .Z(n14413) );
  XNOR U14221 ( .A(p_input[2225]), .B(n14415), .Z(n14414) );
  IV U14222 ( .A(p_input[2209]), .Z(n14415) );
  XNOR U14223 ( .A(n14018), .B(n14408), .Z(n14410) );
  XNOR U14224 ( .A(p_input[2177]), .B(n14416), .Z(n14018) );
  AND U14225 ( .A(n320), .B(n14417), .Z(n14416) );
  XOR U14226 ( .A(p_input[2193]), .B(p_input[2177]), .Z(n14417) );
  IV U14227 ( .A(n14412), .Z(n14408) );
  AND U14228 ( .A(n14283), .B(n14286), .Z(n14412) );
  XOR U14229 ( .A(p_input[2208]), .B(n14418), .Z(n14286) );
  AND U14230 ( .A(n323), .B(n14419), .Z(n14418) );
  XOR U14231 ( .A(p_input[2224]), .B(p_input[2208]), .Z(n14419) );
  XOR U14232 ( .A(n14420), .B(n14421), .Z(n323) );
  AND U14233 ( .A(n14422), .B(n14423), .Z(n14421) );
  XNOR U14234 ( .A(p_input[2239]), .B(n14420), .Z(n14423) );
  XOR U14235 ( .A(n14420), .B(p_input[2223]), .Z(n14422) );
  XOR U14236 ( .A(n14424), .B(n14425), .Z(n14420) );
  AND U14237 ( .A(n14426), .B(n14427), .Z(n14425) );
  XNOR U14238 ( .A(p_input[2238]), .B(n14424), .Z(n14427) );
  XOR U14239 ( .A(n14424), .B(p_input[2222]), .Z(n14426) );
  XOR U14240 ( .A(n14428), .B(n14429), .Z(n14424) );
  AND U14241 ( .A(n14430), .B(n14431), .Z(n14429) );
  XNOR U14242 ( .A(p_input[2237]), .B(n14428), .Z(n14431) );
  XOR U14243 ( .A(n14428), .B(p_input[2221]), .Z(n14430) );
  XOR U14244 ( .A(n14432), .B(n14433), .Z(n14428) );
  AND U14245 ( .A(n14434), .B(n14435), .Z(n14433) );
  XNOR U14246 ( .A(p_input[2236]), .B(n14432), .Z(n14435) );
  XOR U14247 ( .A(n14432), .B(p_input[2220]), .Z(n14434) );
  XOR U14248 ( .A(n14436), .B(n14437), .Z(n14432) );
  AND U14249 ( .A(n14438), .B(n14439), .Z(n14437) );
  XNOR U14250 ( .A(p_input[2235]), .B(n14436), .Z(n14439) );
  XOR U14251 ( .A(n14436), .B(p_input[2219]), .Z(n14438) );
  XOR U14252 ( .A(n14440), .B(n14441), .Z(n14436) );
  AND U14253 ( .A(n14442), .B(n14443), .Z(n14441) );
  XNOR U14254 ( .A(p_input[2234]), .B(n14440), .Z(n14443) );
  XOR U14255 ( .A(n14440), .B(p_input[2218]), .Z(n14442) );
  XOR U14256 ( .A(n14444), .B(n14445), .Z(n14440) );
  AND U14257 ( .A(n14446), .B(n14447), .Z(n14445) );
  XNOR U14258 ( .A(p_input[2233]), .B(n14444), .Z(n14447) );
  XOR U14259 ( .A(n14444), .B(p_input[2217]), .Z(n14446) );
  XOR U14260 ( .A(n14448), .B(n14449), .Z(n14444) );
  AND U14261 ( .A(n14450), .B(n14451), .Z(n14449) );
  XNOR U14262 ( .A(p_input[2232]), .B(n14448), .Z(n14451) );
  XOR U14263 ( .A(n14448), .B(p_input[2216]), .Z(n14450) );
  XOR U14264 ( .A(n14452), .B(n14453), .Z(n14448) );
  AND U14265 ( .A(n14454), .B(n14455), .Z(n14453) );
  XNOR U14266 ( .A(p_input[2231]), .B(n14452), .Z(n14455) );
  XOR U14267 ( .A(n14452), .B(p_input[2215]), .Z(n14454) );
  XOR U14268 ( .A(n14456), .B(n14457), .Z(n14452) );
  AND U14269 ( .A(n14458), .B(n14459), .Z(n14457) );
  XNOR U14270 ( .A(p_input[2230]), .B(n14456), .Z(n14459) );
  XOR U14271 ( .A(n14456), .B(p_input[2214]), .Z(n14458) );
  XOR U14272 ( .A(n14460), .B(n14461), .Z(n14456) );
  AND U14273 ( .A(n14462), .B(n14463), .Z(n14461) );
  XNOR U14274 ( .A(p_input[2229]), .B(n14460), .Z(n14463) );
  XOR U14275 ( .A(n14460), .B(p_input[2213]), .Z(n14462) );
  XOR U14276 ( .A(n14464), .B(n14465), .Z(n14460) );
  AND U14277 ( .A(n14466), .B(n14467), .Z(n14465) );
  XNOR U14278 ( .A(p_input[2228]), .B(n14464), .Z(n14467) );
  XOR U14279 ( .A(n14464), .B(p_input[2212]), .Z(n14466) );
  XOR U14280 ( .A(n14468), .B(n14469), .Z(n14464) );
  AND U14281 ( .A(n14470), .B(n14471), .Z(n14469) );
  XNOR U14282 ( .A(p_input[2227]), .B(n14468), .Z(n14471) );
  XOR U14283 ( .A(n14468), .B(p_input[2211]), .Z(n14470) );
  XOR U14284 ( .A(n14472), .B(n14473), .Z(n14468) );
  AND U14285 ( .A(n14474), .B(n14475), .Z(n14473) );
  XNOR U14286 ( .A(p_input[2226]), .B(n14472), .Z(n14475) );
  XOR U14287 ( .A(n14472), .B(p_input[2210]), .Z(n14474) );
  XNOR U14288 ( .A(n14476), .B(n14477), .Z(n14472) );
  AND U14289 ( .A(n14478), .B(n14479), .Z(n14477) );
  XOR U14290 ( .A(p_input[2225]), .B(n14476), .Z(n14479) );
  XNOR U14291 ( .A(p_input[2209]), .B(n14476), .Z(n14478) );
  AND U14292 ( .A(p_input[2224]), .B(n14480), .Z(n14476) );
  IV U14293 ( .A(p_input[2208]), .Z(n14480) );
  XNOR U14294 ( .A(p_input[2176]), .B(n14481), .Z(n14283) );
  AND U14295 ( .A(n320), .B(n14482), .Z(n14481) );
  XOR U14296 ( .A(p_input[2192]), .B(p_input[2176]), .Z(n14482) );
  XOR U14297 ( .A(n14483), .B(n14484), .Z(n320) );
  AND U14298 ( .A(n14485), .B(n14486), .Z(n14484) );
  XNOR U14299 ( .A(p_input[2207]), .B(n14483), .Z(n14486) );
  XOR U14300 ( .A(n14483), .B(p_input[2191]), .Z(n14485) );
  XOR U14301 ( .A(n14487), .B(n14488), .Z(n14483) );
  AND U14302 ( .A(n14489), .B(n14490), .Z(n14488) );
  XNOR U14303 ( .A(p_input[2206]), .B(n14487), .Z(n14490) );
  XNOR U14304 ( .A(n14487), .B(n14297), .Z(n14489) );
  IV U14305 ( .A(p_input[2190]), .Z(n14297) );
  XOR U14306 ( .A(n14491), .B(n14492), .Z(n14487) );
  AND U14307 ( .A(n14493), .B(n14494), .Z(n14492) );
  XNOR U14308 ( .A(p_input[2205]), .B(n14491), .Z(n14494) );
  XNOR U14309 ( .A(n14491), .B(n14306), .Z(n14493) );
  IV U14310 ( .A(p_input[2189]), .Z(n14306) );
  XOR U14311 ( .A(n14495), .B(n14496), .Z(n14491) );
  AND U14312 ( .A(n14497), .B(n14498), .Z(n14496) );
  XNOR U14313 ( .A(p_input[2204]), .B(n14495), .Z(n14498) );
  XNOR U14314 ( .A(n14495), .B(n14315), .Z(n14497) );
  IV U14315 ( .A(p_input[2188]), .Z(n14315) );
  XOR U14316 ( .A(n14499), .B(n14500), .Z(n14495) );
  AND U14317 ( .A(n14501), .B(n14502), .Z(n14500) );
  XNOR U14318 ( .A(p_input[2203]), .B(n14499), .Z(n14502) );
  XNOR U14319 ( .A(n14499), .B(n14324), .Z(n14501) );
  IV U14320 ( .A(p_input[2187]), .Z(n14324) );
  XOR U14321 ( .A(n14503), .B(n14504), .Z(n14499) );
  AND U14322 ( .A(n14505), .B(n14506), .Z(n14504) );
  XNOR U14323 ( .A(p_input[2202]), .B(n14503), .Z(n14506) );
  XNOR U14324 ( .A(n14503), .B(n14333), .Z(n14505) );
  IV U14325 ( .A(p_input[2186]), .Z(n14333) );
  XOR U14326 ( .A(n14507), .B(n14508), .Z(n14503) );
  AND U14327 ( .A(n14509), .B(n14510), .Z(n14508) );
  XNOR U14328 ( .A(p_input[2201]), .B(n14507), .Z(n14510) );
  XNOR U14329 ( .A(n14507), .B(n14342), .Z(n14509) );
  IV U14330 ( .A(p_input[2185]), .Z(n14342) );
  XOR U14331 ( .A(n14511), .B(n14512), .Z(n14507) );
  AND U14332 ( .A(n14513), .B(n14514), .Z(n14512) );
  XNOR U14333 ( .A(p_input[2200]), .B(n14511), .Z(n14514) );
  XNOR U14334 ( .A(n14511), .B(n14351), .Z(n14513) );
  IV U14335 ( .A(p_input[2184]), .Z(n14351) );
  XOR U14336 ( .A(n14515), .B(n14516), .Z(n14511) );
  AND U14337 ( .A(n14517), .B(n14518), .Z(n14516) );
  XNOR U14338 ( .A(p_input[2199]), .B(n14515), .Z(n14518) );
  XNOR U14339 ( .A(n14515), .B(n14360), .Z(n14517) );
  IV U14340 ( .A(p_input[2183]), .Z(n14360) );
  XOR U14341 ( .A(n14519), .B(n14520), .Z(n14515) );
  AND U14342 ( .A(n14521), .B(n14522), .Z(n14520) );
  XNOR U14343 ( .A(p_input[2198]), .B(n14519), .Z(n14522) );
  XNOR U14344 ( .A(n14519), .B(n14369), .Z(n14521) );
  IV U14345 ( .A(p_input[2182]), .Z(n14369) );
  XOR U14346 ( .A(n14523), .B(n14524), .Z(n14519) );
  AND U14347 ( .A(n14525), .B(n14526), .Z(n14524) );
  XNOR U14348 ( .A(p_input[2197]), .B(n14523), .Z(n14526) );
  XNOR U14349 ( .A(n14523), .B(n14378), .Z(n14525) );
  IV U14350 ( .A(p_input[2181]), .Z(n14378) );
  XOR U14351 ( .A(n14527), .B(n14528), .Z(n14523) );
  AND U14352 ( .A(n14529), .B(n14530), .Z(n14528) );
  XNOR U14353 ( .A(p_input[2196]), .B(n14527), .Z(n14530) );
  XNOR U14354 ( .A(n14527), .B(n14387), .Z(n14529) );
  IV U14355 ( .A(p_input[2180]), .Z(n14387) );
  XOR U14356 ( .A(n14531), .B(n14532), .Z(n14527) );
  AND U14357 ( .A(n14533), .B(n14534), .Z(n14532) );
  XNOR U14358 ( .A(p_input[2195]), .B(n14531), .Z(n14534) );
  XNOR U14359 ( .A(n14531), .B(n14396), .Z(n14533) );
  IV U14360 ( .A(p_input[2179]), .Z(n14396) );
  XOR U14361 ( .A(n14535), .B(n14536), .Z(n14531) );
  AND U14362 ( .A(n14537), .B(n14538), .Z(n14536) );
  XNOR U14363 ( .A(p_input[2194]), .B(n14535), .Z(n14538) );
  XNOR U14364 ( .A(n14535), .B(n14405), .Z(n14537) );
  IV U14365 ( .A(p_input[2178]), .Z(n14405) );
  XNOR U14366 ( .A(n14539), .B(n14540), .Z(n14535) );
  AND U14367 ( .A(n14541), .B(n14542), .Z(n14540) );
  XOR U14368 ( .A(p_input[2193]), .B(n14539), .Z(n14542) );
  XNOR U14369 ( .A(p_input[2177]), .B(n14539), .Z(n14541) );
  AND U14370 ( .A(p_input[2192]), .B(n14543), .Z(n14539) );
  IV U14371 ( .A(p_input[2176]), .Z(n14543) );
  XOR U14372 ( .A(n14544), .B(n14545), .Z(n13659) );
  AND U14373 ( .A(n776), .B(n14546), .Z(n14545) );
  XNOR U14374 ( .A(n14547), .B(n14544), .Z(n14546) );
  XOR U14375 ( .A(n14548), .B(n14549), .Z(n776) );
  AND U14376 ( .A(n14550), .B(n14551), .Z(n14549) );
  XNOR U14377 ( .A(n13671), .B(n14548), .Z(n14551) );
  AND U14378 ( .A(n14552), .B(n14553), .Z(n13671) );
  XOR U14379 ( .A(n14548), .B(n13670), .Z(n14550) );
  AND U14380 ( .A(n14554), .B(n14555), .Z(n13670) );
  XOR U14381 ( .A(n14556), .B(n14557), .Z(n14548) );
  AND U14382 ( .A(n14558), .B(n14559), .Z(n14557) );
  XOR U14383 ( .A(n14556), .B(n13683), .Z(n14559) );
  XOR U14384 ( .A(n14560), .B(n14561), .Z(n13683) );
  AND U14385 ( .A(n463), .B(n14562), .Z(n14561) );
  XOR U14386 ( .A(n14563), .B(n14560), .Z(n14562) );
  XNOR U14387 ( .A(n13680), .B(n14556), .Z(n14558) );
  XOR U14388 ( .A(n14564), .B(n14565), .Z(n13680) );
  AND U14389 ( .A(n460), .B(n14566), .Z(n14565) );
  XOR U14390 ( .A(n14567), .B(n14564), .Z(n14566) );
  XOR U14391 ( .A(n14568), .B(n14569), .Z(n14556) );
  AND U14392 ( .A(n14570), .B(n14571), .Z(n14569) );
  XOR U14393 ( .A(n14568), .B(n13695), .Z(n14571) );
  XOR U14394 ( .A(n14572), .B(n14573), .Z(n13695) );
  AND U14395 ( .A(n463), .B(n14574), .Z(n14573) );
  XOR U14396 ( .A(n14575), .B(n14572), .Z(n14574) );
  XNOR U14397 ( .A(n13692), .B(n14568), .Z(n14570) );
  XOR U14398 ( .A(n14576), .B(n14577), .Z(n13692) );
  AND U14399 ( .A(n460), .B(n14578), .Z(n14577) );
  XOR U14400 ( .A(n14579), .B(n14576), .Z(n14578) );
  XOR U14401 ( .A(n14580), .B(n14581), .Z(n14568) );
  AND U14402 ( .A(n14582), .B(n14583), .Z(n14581) );
  XOR U14403 ( .A(n14580), .B(n13707), .Z(n14583) );
  XOR U14404 ( .A(n14584), .B(n14585), .Z(n13707) );
  AND U14405 ( .A(n463), .B(n14586), .Z(n14585) );
  XOR U14406 ( .A(n14587), .B(n14584), .Z(n14586) );
  XNOR U14407 ( .A(n13704), .B(n14580), .Z(n14582) );
  XOR U14408 ( .A(n14588), .B(n14589), .Z(n13704) );
  AND U14409 ( .A(n460), .B(n14590), .Z(n14589) );
  XOR U14410 ( .A(n14591), .B(n14588), .Z(n14590) );
  XOR U14411 ( .A(n14592), .B(n14593), .Z(n14580) );
  AND U14412 ( .A(n14594), .B(n14595), .Z(n14593) );
  XOR U14413 ( .A(n14592), .B(n13719), .Z(n14595) );
  XOR U14414 ( .A(n14596), .B(n14597), .Z(n13719) );
  AND U14415 ( .A(n463), .B(n14598), .Z(n14597) );
  XOR U14416 ( .A(n14599), .B(n14596), .Z(n14598) );
  XNOR U14417 ( .A(n13716), .B(n14592), .Z(n14594) );
  XOR U14418 ( .A(n14600), .B(n14601), .Z(n13716) );
  AND U14419 ( .A(n460), .B(n14602), .Z(n14601) );
  XOR U14420 ( .A(n14603), .B(n14600), .Z(n14602) );
  XOR U14421 ( .A(n14604), .B(n14605), .Z(n14592) );
  AND U14422 ( .A(n14606), .B(n14607), .Z(n14605) );
  XOR U14423 ( .A(n14604), .B(n13731), .Z(n14607) );
  XOR U14424 ( .A(n14608), .B(n14609), .Z(n13731) );
  AND U14425 ( .A(n463), .B(n14610), .Z(n14609) );
  XOR U14426 ( .A(n14611), .B(n14608), .Z(n14610) );
  XNOR U14427 ( .A(n13728), .B(n14604), .Z(n14606) );
  XOR U14428 ( .A(n14612), .B(n14613), .Z(n13728) );
  AND U14429 ( .A(n460), .B(n14614), .Z(n14613) );
  XOR U14430 ( .A(n14615), .B(n14612), .Z(n14614) );
  XOR U14431 ( .A(n14616), .B(n14617), .Z(n14604) );
  AND U14432 ( .A(n14618), .B(n14619), .Z(n14617) );
  XOR U14433 ( .A(n14616), .B(n13743), .Z(n14619) );
  XOR U14434 ( .A(n14620), .B(n14621), .Z(n13743) );
  AND U14435 ( .A(n463), .B(n14622), .Z(n14621) );
  XOR U14436 ( .A(n14623), .B(n14620), .Z(n14622) );
  XNOR U14437 ( .A(n13740), .B(n14616), .Z(n14618) );
  XOR U14438 ( .A(n14624), .B(n14625), .Z(n13740) );
  AND U14439 ( .A(n460), .B(n14626), .Z(n14625) );
  XOR U14440 ( .A(n14627), .B(n14624), .Z(n14626) );
  XOR U14441 ( .A(n14628), .B(n14629), .Z(n14616) );
  AND U14442 ( .A(n14630), .B(n14631), .Z(n14629) );
  XOR U14443 ( .A(n14628), .B(n13755), .Z(n14631) );
  XOR U14444 ( .A(n14632), .B(n14633), .Z(n13755) );
  AND U14445 ( .A(n463), .B(n14634), .Z(n14633) );
  XOR U14446 ( .A(n14635), .B(n14632), .Z(n14634) );
  XNOR U14447 ( .A(n13752), .B(n14628), .Z(n14630) );
  XOR U14448 ( .A(n14636), .B(n14637), .Z(n13752) );
  AND U14449 ( .A(n460), .B(n14638), .Z(n14637) );
  XOR U14450 ( .A(n14639), .B(n14636), .Z(n14638) );
  XOR U14451 ( .A(n14640), .B(n14641), .Z(n14628) );
  AND U14452 ( .A(n14642), .B(n14643), .Z(n14641) );
  XOR U14453 ( .A(n14640), .B(n13767), .Z(n14643) );
  XOR U14454 ( .A(n14644), .B(n14645), .Z(n13767) );
  AND U14455 ( .A(n463), .B(n14646), .Z(n14645) );
  XOR U14456 ( .A(n14647), .B(n14644), .Z(n14646) );
  XNOR U14457 ( .A(n13764), .B(n14640), .Z(n14642) );
  XOR U14458 ( .A(n14648), .B(n14649), .Z(n13764) );
  AND U14459 ( .A(n460), .B(n14650), .Z(n14649) );
  XOR U14460 ( .A(n14651), .B(n14648), .Z(n14650) );
  XOR U14461 ( .A(n14652), .B(n14653), .Z(n14640) );
  AND U14462 ( .A(n14654), .B(n14655), .Z(n14653) );
  XOR U14463 ( .A(n14652), .B(n13779), .Z(n14655) );
  XOR U14464 ( .A(n14656), .B(n14657), .Z(n13779) );
  AND U14465 ( .A(n463), .B(n14658), .Z(n14657) );
  XOR U14466 ( .A(n14659), .B(n14656), .Z(n14658) );
  XNOR U14467 ( .A(n13776), .B(n14652), .Z(n14654) );
  XOR U14468 ( .A(n14660), .B(n14661), .Z(n13776) );
  AND U14469 ( .A(n460), .B(n14662), .Z(n14661) );
  XOR U14470 ( .A(n14663), .B(n14660), .Z(n14662) );
  XOR U14471 ( .A(n14664), .B(n14665), .Z(n14652) );
  AND U14472 ( .A(n14666), .B(n14667), .Z(n14665) );
  XOR U14473 ( .A(n14664), .B(n13791), .Z(n14667) );
  XOR U14474 ( .A(n14668), .B(n14669), .Z(n13791) );
  AND U14475 ( .A(n463), .B(n14670), .Z(n14669) );
  XOR U14476 ( .A(n14671), .B(n14668), .Z(n14670) );
  XNOR U14477 ( .A(n13788), .B(n14664), .Z(n14666) );
  XOR U14478 ( .A(n14672), .B(n14673), .Z(n13788) );
  AND U14479 ( .A(n460), .B(n14674), .Z(n14673) );
  XOR U14480 ( .A(n14675), .B(n14672), .Z(n14674) );
  XOR U14481 ( .A(n14676), .B(n14677), .Z(n14664) );
  AND U14482 ( .A(n14678), .B(n14679), .Z(n14677) );
  XOR U14483 ( .A(n14676), .B(n13803), .Z(n14679) );
  XOR U14484 ( .A(n14680), .B(n14681), .Z(n13803) );
  AND U14485 ( .A(n463), .B(n14682), .Z(n14681) );
  XOR U14486 ( .A(n14683), .B(n14680), .Z(n14682) );
  XNOR U14487 ( .A(n13800), .B(n14676), .Z(n14678) );
  XOR U14488 ( .A(n14684), .B(n14685), .Z(n13800) );
  AND U14489 ( .A(n460), .B(n14686), .Z(n14685) );
  XOR U14490 ( .A(n14687), .B(n14684), .Z(n14686) );
  XOR U14491 ( .A(n14688), .B(n14689), .Z(n14676) );
  AND U14492 ( .A(n14690), .B(n14691), .Z(n14689) );
  XOR U14493 ( .A(n14688), .B(n13815), .Z(n14691) );
  XOR U14494 ( .A(n14692), .B(n14693), .Z(n13815) );
  AND U14495 ( .A(n463), .B(n14694), .Z(n14693) );
  XOR U14496 ( .A(n14695), .B(n14692), .Z(n14694) );
  XNOR U14497 ( .A(n13812), .B(n14688), .Z(n14690) );
  XOR U14498 ( .A(n14696), .B(n14697), .Z(n13812) );
  AND U14499 ( .A(n460), .B(n14698), .Z(n14697) );
  XOR U14500 ( .A(n14699), .B(n14696), .Z(n14698) );
  XOR U14501 ( .A(n14700), .B(n14701), .Z(n14688) );
  AND U14502 ( .A(n14702), .B(n14703), .Z(n14701) );
  XOR U14503 ( .A(n14700), .B(n13827), .Z(n14703) );
  XOR U14504 ( .A(n14704), .B(n14705), .Z(n13827) );
  AND U14505 ( .A(n463), .B(n14706), .Z(n14705) );
  XOR U14506 ( .A(n14707), .B(n14704), .Z(n14706) );
  XNOR U14507 ( .A(n13824), .B(n14700), .Z(n14702) );
  XOR U14508 ( .A(n14708), .B(n14709), .Z(n13824) );
  AND U14509 ( .A(n460), .B(n14710), .Z(n14709) );
  XOR U14510 ( .A(n14711), .B(n14708), .Z(n14710) );
  XOR U14511 ( .A(n14712), .B(n14713), .Z(n14700) );
  AND U14512 ( .A(n14714), .B(n14715), .Z(n14713) );
  XNOR U14513 ( .A(n14716), .B(n13840), .Z(n14715) );
  XOR U14514 ( .A(n14717), .B(n14718), .Z(n13840) );
  AND U14515 ( .A(n463), .B(n14719), .Z(n14718) );
  XOR U14516 ( .A(n14717), .B(n14720), .Z(n14719) );
  XNOR U14517 ( .A(n13837), .B(n14712), .Z(n14714) );
  XOR U14518 ( .A(n14721), .B(n14722), .Z(n13837) );
  AND U14519 ( .A(n460), .B(n14723), .Z(n14722) );
  XOR U14520 ( .A(n14721), .B(n14724), .Z(n14723) );
  IV U14521 ( .A(n14716), .Z(n14712) );
  AND U14522 ( .A(n14544), .B(n14547), .Z(n14716) );
  XNOR U14523 ( .A(n14725), .B(n14726), .Z(n14547) );
  AND U14524 ( .A(n463), .B(n14727), .Z(n14726) );
  XNOR U14525 ( .A(n14728), .B(n14725), .Z(n14727) );
  XOR U14526 ( .A(n14729), .B(n14730), .Z(n463) );
  AND U14527 ( .A(n14731), .B(n14732), .Z(n14730) );
  XNOR U14528 ( .A(n14552), .B(n14729), .Z(n14732) );
  AND U14529 ( .A(p_input[2175]), .B(p_input[2159]), .Z(n14552) );
  XOR U14530 ( .A(n14729), .B(n14553), .Z(n14731) );
  AND U14531 ( .A(p_input[2143]), .B(p_input[2127]), .Z(n14553) );
  XOR U14532 ( .A(n14733), .B(n14734), .Z(n14729) );
  AND U14533 ( .A(n14735), .B(n14736), .Z(n14734) );
  XOR U14534 ( .A(n14733), .B(n14563), .Z(n14736) );
  XNOR U14535 ( .A(p_input[2158]), .B(n14737), .Z(n14563) );
  AND U14536 ( .A(n331), .B(n14738), .Z(n14737) );
  XOR U14537 ( .A(p_input[2174]), .B(p_input[2158]), .Z(n14738) );
  XNOR U14538 ( .A(n14560), .B(n14733), .Z(n14735) );
  XOR U14539 ( .A(n14739), .B(n14740), .Z(n14560) );
  AND U14540 ( .A(n329), .B(n14741), .Z(n14740) );
  XOR U14541 ( .A(p_input[2142]), .B(p_input[2126]), .Z(n14741) );
  XOR U14542 ( .A(n14742), .B(n14743), .Z(n14733) );
  AND U14543 ( .A(n14744), .B(n14745), .Z(n14743) );
  XOR U14544 ( .A(n14742), .B(n14575), .Z(n14745) );
  XNOR U14545 ( .A(p_input[2157]), .B(n14746), .Z(n14575) );
  AND U14546 ( .A(n331), .B(n14747), .Z(n14746) );
  XOR U14547 ( .A(p_input[2173]), .B(p_input[2157]), .Z(n14747) );
  XNOR U14548 ( .A(n14572), .B(n14742), .Z(n14744) );
  XOR U14549 ( .A(n14748), .B(n14749), .Z(n14572) );
  AND U14550 ( .A(n329), .B(n14750), .Z(n14749) );
  XOR U14551 ( .A(p_input[2141]), .B(p_input[2125]), .Z(n14750) );
  XOR U14552 ( .A(n14751), .B(n14752), .Z(n14742) );
  AND U14553 ( .A(n14753), .B(n14754), .Z(n14752) );
  XOR U14554 ( .A(n14751), .B(n14587), .Z(n14754) );
  XNOR U14555 ( .A(p_input[2156]), .B(n14755), .Z(n14587) );
  AND U14556 ( .A(n331), .B(n14756), .Z(n14755) );
  XOR U14557 ( .A(p_input[2172]), .B(p_input[2156]), .Z(n14756) );
  XNOR U14558 ( .A(n14584), .B(n14751), .Z(n14753) );
  XOR U14559 ( .A(n14757), .B(n14758), .Z(n14584) );
  AND U14560 ( .A(n329), .B(n14759), .Z(n14758) );
  XOR U14561 ( .A(p_input[2140]), .B(p_input[2124]), .Z(n14759) );
  XOR U14562 ( .A(n14760), .B(n14761), .Z(n14751) );
  AND U14563 ( .A(n14762), .B(n14763), .Z(n14761) );
  XOR U14564 ( .A(n14760), .B(n14599), .Z(n14763) );
  XNOR U14565 ( .A(p_input[2155]), .B(n14764), .Z(n14599) );
  AND U14566 ( .A(n331), .B(n14765), .Z(n14764) );
  XOR U14567 ( .A(p_input[2171]), .B(p_input[2155]), .Z(n14765) );
  XNOR U14568 ( .A(n14596), .B(n14760), .Z(n14762) );
  XOR U14569 ( .A(n14766), .B(n14767), .Z(n14596) );
  AND U14570 ( .A(n329), .B(n14768), .Z(n14767) );
  XOR U14571 ( .A(p_input[2139]), .B(p_input[2123]), .Z(n14768) );
  XOR U14572 ( .A(n14769), .B(n14770), .Z(n14760) );
  AND U14573 ( .A(n14771), .B(n14772), .Z(n14770) );
  XOR U14574 ( .A(n14769), .B(n14611), .Z(n14772) );
  XNOR U14575 ( .A(p_input[2154]), .B(n14773), .Z(n14611) );
  AND U14576 ( .A(n331), .B(n14774), .Z(n14773) );
  XOR U14577 ( .A(p_input[2170]), .B(p_input[2154]), .Z(n14774) );
  XNOR U14578 ( .A(n14608), .B(n14769), .Z(n14771) );
  XOR U14579 ( .A(n14775), .B(n14776), .Z(n14608) );
  AND U14580 ( .A(n329), .B(n14777), .Z(n14776) );
  XOR U14581 ( .A(p_input[2138]), .B(p_input[2122]), .Z(n14777) );
  XOR U14582 ( .A(n14778), .B(n14779), .Z(n14769) );
  AND U14583 ( .A(n14780), .B(n14781), .Z(n14779) );
  XOR U14584 ( .A(n14778), .B(n14623), .Z(n14781) );
  XNOR U14585 ( .A(p_input[2153]), .B(n14782), .Z(n14623) );
  AND U14586 ( .A(n331), .B(n14783), .Z(n14782) );
  XOR U14587 ( .A(p_input[2169]), .B(p_input[2153]), .Z(n14783) );
  XNOR U14588 ( .A(n14620), .B(n14778), .Z(n14780) );
  XOR U14589 ( .A(n14784), .B(n14785), .Z(n14620) );
  AND U14590 ( .A(n329), .B(n14786), .Z(n14785) );
  XOR U14591 ( .A(p_input[2137]), .B(p_input[2121]), .Z(n14786) );
  XOR U14592 ( .A(n14787), .B(n14788), .Z(n14778) );
  AND U14593 ( .A(n14789), .B(n14790), .Z(n14788) );
  XOR U14594 ( .A(n14787), .B(n14635), .Z(n14790) );
  XNOR U14595 ( .A(p_input[2152]), .B(n14791), .Z(n14635) );
  AND U14596 ( .A(n331), .B(n14792), .Z(n14791) );
  XOR U14597 ( .A(p_input[2168]), .B(p_input[2152]), .Z(n14792) );
  XNOR U14598 ( .A(n14632), .B(n14787), .Z(n14789) );
  XOR U14599 ( .A(n14793), .B(n14794), .Z(n14632) );
  AND U14600 ( .A(n329), .B(n14795), .Z(n14794) );
  XOR U14601 ( .A(p_input[2136]), .B(p_input[2120]), .Z(n14795) );
  XOR U14602 ( .A(n14796), .B(n14797), .Z(n14787) );
  AND U14603 ( .A(n14798), .B(n14799), .Z(n14797) );
  XOR U14604 ( .A(n14796), .B(n14647), .Z(n14799) );
  XNOR U14605 ( .A(p_input[2151]), .B(n14800), .Z(n14647) );
  AND U14606 ( .A(n331), .B(n14801), .Z(n14800) );
  XOR U14607 ( .A(p_input[2167]), .B(p_input[2151]), .Z(n14801) );
  XNOR U14608 ( .A(n14644), .B(n14796), .Z(n14798) );
  XOR U14609 ( .A(n14802), .B(n14803), .Z(n14644) );
  AND U14610 ( .A(n329), .B(n14804), .Z(n14803) );
  XOR U14611 ( .A(p_input[2135]), .B(p_input[2119]), .Z(n14804) );
  XOR U14612 ( .A(n14805), .B(n14806), .Z(n14796) );
  AND U14613 ( .A(n14807), .B(n14808), .Z(n14806) );
  XOR U14614 ( .A(n14805), .B(n14659), .Z(n14808) );
  XNOR U14615 ( .A(p_input[2150]), .B(n14809), .Z(n14659) );
  AND U14616 ( .A(n331), .B(n14810), .Z(n14809) );
  XOR U14617 ( .A(p_input[2166]), .B(p_input[2150]), .Z(n14810) );
  XNOR U14618 ( .A(n14656), .B(n14805), .Z(n14807) );
  XOR U14619 ( .A(n14811), .B(n14812), .Z(n14656) );
  AND U14620 ( .A(n329), .B(n14813), .Z(n14812) );
  XOR U14621 ( .A(p_input[2134]), .B(p_input[2118]), .Z(n14813) );
  XOR U14622 ( .A(n14814), .B(n14815), .Z(n14805) );
  AND U14623 ( .A(n14816), .B(n14817), .Z(n14815) );
  XOR U14624 ( .A(n14814), .B(n14671), .Z(n14817) );
  XNOR U14625 ( .A(p_input[2149]), .B(n14818), .Z(n14671) );
  AND U14626 ( .A(n331), .B(n14819), .Z(n14818) );
  XOR U14627 ( .A(p_input[2165]), .B(p_input[2149]), .Z(n14819) );
  XNOR U14628 ( .A(n14668), .B(n14814), .Z(n14816) );
  XOR U14629 ( .A(n14820), .B(n14821), .Z(n14668) );
  AND U14630 ( .A(n329), .B(n14822), .Z(n14821) );
  XOR U14631 ( .A(p_input[2133]), .B(p_input[2117]), .Z(n14822) );
  XOR U14632 ( .A(n14823), .B(n14824), .Z(n14814) );
  AND U14633 ( .A(n14825), .B(n14826), .Z(n14824) );
  XOR U14634 ( .A(n14823), .B(n14683), .Z(n14826) );
  XNOR U14635 ( .A(p_input[2148]), .B(n14827), .Z(n14683) );
  AND U14636 ( .A(n331), .B(n14828), .Z(n14827) );
  XOR U14637 ( .A(p_input[2164]), .B(p_input[2148]), .Z(n14828) );
  XNOR U14638 ( .A(n14680), .B(n14823), .Z(n14825) );
  XOR U14639 ( .A(n14829), .B(n14830), .Z(n14680) );
  AND U14640 ( .A(n329), .B(n14831), .Z(n14830) );
  XOR U14641 ( .A(p_input[2132]), .B(p_input[2116]), .Z(n14831) );
  XOR U14642 ( .A(n14832), .B(n14833), .Z(n14823) );
  AND U14643 ( .A(n14834), .B(n14835), .Z(n14833) );
  XOR U14644 ( .A(n14832), .B(n14695), .Z(n14835) );
  XNOR U14645 ( .A(p_input[2147]), .B(n14836), .Z(n14695) );
  AND U14646 ( .A(n331), .B(n14837), .Z(n14836) );
  XOR U14647 ( .A(p_input[2163]), .B(p_input[2147]), .Z(n14837) );
  XNOR U14648 ( .A(n14692), .B(n14832), .Z(n14834) );
  XOR U14649 ( .A(n14838), .B(n14839), .Z(n14692) );
  AND U14650 ( .A(n329), .B(n14840), .Z(n14839) );
  XOR U14651 ( .A(p_input[2131]), .B(p_input[2115]), .Z(n14840) );
  XOR U14652 ( .A(n14841), .B(n14842), .Z(n14832) );
  AND U14653 ( .A(n14843), .B(n14844), .Z(n14842) );
  XOR U14654 ( .A(n14841), .B(n14707), .Z(n14844) );
  XNOR U14655 ( .A(p_input[2146]), .B(n14845), .Z(n14707) );
  AND U14656 ( .A(n331), .B(n14846), .Z(n14845) );
  XOR U14657 ( .A(p_input[2162]), .B(p_input[2146]), .Z(n14846) );
  XNOR U14658 ( .A(n14704), .B(n14841), .Z(n14843) );
  XOR U14659 ( .A(n14847), .B(n14848), .Z(n14704) );
  AND U14660 ( .A(n329), .B(n14849), .Z(n14848) );
  XOR U14661 ( .A(p_input[2130]), .B(p_input[2114]), .Z(n14849) );
  XOR U14662 ( .A(n14850), .B(n14851), .Z(n14841) );
  AND U14663 ( .A(n14852), .B(n14853), .Z(n14851) );
  XNOR U14664 ( .A(n14854), .B(n14720), .Z(n14853) );
  XNOR U14665 ( .A(p_input[2145]), .B(n14855), .Z(n14720) );
  AND U14666 ( .A(n331), .B(n14856), .Z(n14855) );
  XNOR U14667 ( .A(p_input[2161]), .B(n14857), .Z(n14856) );
  IV U14668 ( .A(p_input[2145]), .Z(n14857) );
  XNOR U14669 ( .A(n14717), .B(n14850), .Z(n14852) );
  XNOR U14670 ( .A(p_input[2113]), .B(n14858), .Z(n14717) );
  AND U14671 ( .A(n329), .B(n14859), .Z(n14858) );
  XOR U14672 ( .A(p_input[2129]), .B(p_input[2113]), .Z(n14859) );
  IV U14673 ( .A(n14854), .Z(n14850) );
  AND U14674 ( .A(n14725), .B(n14728), .Z(n14854) );
  XOR U14675 ( .A(p_input[2144]), .B(n14860), .Z(n14728) );
  AND U14676 ( .A(n331), .B(n14861), .Z(n14860) );
  XOR U14677 ( .A(p_input[2160]), .B(p_input[2144]), .Z(n14861) );
  XOR U14678 ( .A(n14862), .B(n14863), .Z(n331) );
  AND U14679 ( .A(n14864), .B(n14865), .Z(n14863) );
  XNOR U14680 ( .A(p_input[2175]), .B(n14862), .Z(n14865) );
  XOR U14681 ( .A(n14862), .B(p_input[2159]), .Z(n14864) );
  XOR U14682 ( .A(n14866), .B(n14867), .Z(n14862) );
  AND U14683 ( .A(n14868), .B(n14869), .Z(n14867) );
  XNOR U14684 ( .A(p_input[2174]), .B(n14866), .Z(n14869) );
  XOR U14685 ( .A(n14866), .B(p_input[2158]), .Z(n14868) );
  XOR U14686 ( .A(n14870), .B(n14871), .Z(n14866) );
  AND U14687 ( .A(n14872), .B(n14873), .Z(n14871) );
  XNOR U14688 ( .A(p_input[2173]), .B(n14870), .Z(n14873) );
  XOR U14689 ( .A(n14870), .B(p_input[2157]), .Z(n14872) );
  XOR U14690 ( .A(n14874), .B(n14875), .Z(n14870) );
  AND U14691 ( .A(n14876), .B(n14877), .Z(n14875) );
  XNOR U14692 ( .A(p_input[2172]), .B(n14874), .Z(n14877) );
  XOR U14693 ( .A(n14874), .B(p_input[2156]), .Z(n14876) );
  XOR U14694 ( .A(n14878), .B(n14879), .Z(n14874) );
  AND U14695 ( .A(n14880), .B(n14881), .Z(n14879) );
  XNOR U14696 ( .A(p_input[2171]), .B(n14878), .Z(n14881) );
  XOR U14697 ( .A(n14878), .B(p_input[2155]), .Z(n14880) );
  XOR U14698 ( .A(n14882), .B(n14883), .Z(n14878) );
  AND U14699 ( .A(n14884), .B(n14885), .Z(n14883) );
  XNOR U14700 ( .A(p_input[2170]), .B(n14882), .Z(n14885) );
  XOR U14701 ( .A(n14882), .B(p_input[2154]), .Z(n14884) );
  XOR U14702 ( .A(n14886), .B(n14887), .Z(n14882) );
  AND U14703 ( .A(n14888), .B(n14889), .Z(n14887) );
  XNOR U14704 ( .A(p_input[2169]), .B(n14886), .Z(n14889) );
  XOR U14705 ( .A(n14886), .B(p_input[2153]), .Z(n14888) );
  XOR U14706 ( .A(n14890), .B(n14891), .Z(n14886) );
  AND U14707 ( .A(n14892), .B(n14893), .Z(n14891) );
  XNOR U14708 ( .A(p_input[2168]), .B(n14890), .Z(n14893) );
  XOR U14709 ( .A(n14890), .B(p_input[2152]), .Z(n14892) );
  XOR U14710 ( .A(n14894), .B(n14895), .Z(n14890) );
  AND U14711 ( .A(n14896), .B(n14897), .Z(n14895) );
  XNOR U14712 ( .A(p_input[2167]), .B(n14894), .Z(n14897) );
  XOR U14713 ( .A(n14894), .B(p_input[2151]), .Z(n14896) );
  XOR U14714 ( .A(n14898), .B(n14899), .Z(n14894) );
  AND U14715 ( .A(n14900), .B(n14901), .Z(n14899) );
  XNOR U14716 ( .A(p_input[2166]), .B(n14898), .Z(n14901) );
  XOR U14717 ( .A(n14898), .B(p_input[2150]), .Z(n14900) );
  XOR U14718 ( .A(n14902), .B(n14903), .Z(n14898) );
  AND U14719 ( .A(n14904), .B(n14905), .Z(n14903) );
  XNOR U14720 ( .A(p_input[2165]), .B(n14902), .Z(n14905) );
  XOR U14721 ( .A(n14902), .B(p_input[2149]), .Z(n14904) );
  XOR U14722 ( .A(n14906), .B(n14907), .Z(n14902) );
  AND U14723 ( .A(n14908), .B(n14909), .Z(n14907) );
  XNOR U14724 ( .A(p_input[2164]), .B(n14906), .Z(n14909) );
  XOR U14725 ( .A(n14906), .B(p_input[2148]), .Z(n14908) );
  XOR U14726 ( .A(n14910), .B(n14911), .Z(n14906) );
  AND U14727 ( .A(n14912), .B(n14913), .Z(n14911) );
  XNOR U14728 ( .A(p_input[2163]), .B(n14910), .Z(n14913) );
  XOR U14729 ( .A(n14910), .B(p_input[2147]), .Z(n14912) );
  XOR U14730 ( .A(n14914), .B(n14915), .Z(n14910) );
  AND U14731 ( .A(n14916), .B(n14917), .Z(n14915) );
  XNOR U14732 ( .A(p_input[2162]), .B(n14914), .Z(n14917) );
  XOR U14733 ( .A(n14914), .B(p_input[2146]), .Z(n14916) );
  XNOR U14734 ( .A(n14918), .B(n14919), .Z(n14914) );
  AND U14735 ( .A(n14920), .B(n14921), .Z(n14919) );
  XOR U14736 ( .A(p_input[2161]), .B(n14918), .Z(n14921) );
  XNOR U14737 ( .A(p_input[2145]), .B(n14918), .Z(n14920) );
  AND U14738 ( .A(p_input[2160]), .B(n14922), .Z(n14918) );
  IV U14739 ( .A(p_input[2144]), .Z(n14922) );
  XNOR U14740 ( .A(p_input[2112]), .B(n14923), .Z(n14725) );
  AND U14741 ( .A(n329), .B(n14924), .Z(n14923) );
  XOR U14742 ( .A(p_input[2128]), .B(p_input[2112]), .Z(n14924) );
  XOR U14743 ( .A(n14925), .B(n14926), .Z(n329) );
  AND U14744 ( .A(n14927), .B(n14928), .Z(n14926) );
  XNOR U14745 ( .A(p_input[2143]), .B(n14925), .Z(n14928) );
  XOR U14746 ( .A(n14925), .B(p_input[2127]), .Z(n14927) );
  XOR U14747 ( .A(n14929), .B(n14930), .Z(n14925) );
  AND U14748 ( .A(n14931), .B(n14932), .Z(n14930) );
  XNOR U14749 ( .A(p_input[2142]), .B(n14929), .Z(n14932) );
  XNOR U14750 ( .A(n14929), .B(n14739), .Z(n14931) );
  IV U14751 ( .A(p_input[2126]), .Z(n14739) );
  XOR U14752 ( .A(n14933), .B(n14934), .Z(n14929) );
  AND U14753 ( .A(n14935), .B(n14936), .Z(n14934) );
  XNOR U14754 ( .A(p_input[2141]), .B(n14933), .Z(n14936) );
  XNOR U14755 ( .A(n14933), .B(n14748), .Z(n14935) );
  IV U14756 ( .A(p_input[2125]), .Z(n14748) );
  XOR U14757 ( .A(n14937), .B(n14938), .Z(n14933) );
  AND U14758 ( .A(n14939), .B(n14940), .Z(n14938) );
  XNOR U14759 ( .A(p_input[2140]), .B(n14937), .Z(n14940) );
  XNOR U14760 ( .A(n14937), .B(n14757), .Z(n14939) );
  IV U14761 ( .A(p_input[2124]), .Z(n14757) );
  XOR U14762 ( .A(n14941), .B(n14942), .Z(n14937) );
  AND U14763 ( .A(n14943), .B(n14944), .Z(n14942) );
  XNOR U14764 ( .A(p_input[2139]), .B(n14941), .Z(n14944) );
  XNOR U14765 ( .A(n14941), .B(n14766), .Z(n14943) );
  IV U14766 ( .A(p_input[2123]), .Z(n14766) );
  XOR U14767 ( .A(n14945), .B(n14946), .Z(n14941) );
  AND U14768 ( .A(n14947), .B(n14948), .Z(n14946) );
  XNOR U14769 ( .A(p_input[2138]), .B(n14945), .Z(n14948) );
  XNOR U14770 ( .A(n14945), .B(n14775), .Z(n14947) );
  IV U14771 ( .A(p_input[2122]), .Z(n14775) );
  XOR U14772 ( .A(n14949), .B(n14950), .Z(n14945) );
  AND U14773 ( .A(n14951), .B(n14952), .Z(n14950) );
  XNOR U14774 ( .A(p_input[2137]), .B(n14949), .Z(n14952) );
  XNOR U14775 ( .A(n14949), .B(n14784), .Z(n14951) );
  IV U14776 ( .A(p_input[2121]), .Z(n14784) );
  XOR U14777 ( .A(n14953), .B(n14954), .Z(n14949) );
  AND U14778 ( .A(n14955), .B(n14956), .Z(n14954) );
  XNOR U14779 ( .A(p_input[2136]), .B(n14953), .Z(n14956) );
  XNOR U14780 ( .A(n14953), .B(n14793), .Z(n14955) );
  IV U14781 ( .A(p_input[2120]), .Z(n14793) );
  XOR U14782 ( .A(n14957), .B(n14958), .Z(n14953) );
  AND U14783 ( .A(n14959), .B(n14960), .Z(n14958) );
  XNOR U14784 ( .A(p_input[2135]), .B(n14957), .Z(n14960) );
  XNOR U14785 ( .A(n14957), .B(n14802), .Z(n14959) );
  IV U14786 ( .A(p_input[2119]), .Z(n14802) );
  XOR U14787 ( .A(n14961), .B(n14962), .Z(n14957) );
  AND U14788 ( .A(n14963), .B(n14964), .Z(n14962) );
  XNOR U14789 ( .A(p_input[2134]), .B(n14961), .Z(n14964) );
  XNOR U14790 ( .A(n14961), .B(n14811), .Z(n14963) );
  IV U14791 ( .A(p_input[2118]), .Z(n14811) );
  XOR U14792 ( .A(n14965), .B(n14966), .Z(n14961) );
  AND U14793 ( .A(n14967), .B(n14968), .Z(n14966) );
  XNOR U14794 ( .A(p_input[2133]), .B(n14965), .Z(n14968) );
  XNOR U14795 ( .A(n14965), .B(n14820), .Z(n14967) );
  IV U14796 ( .A(p_input[2117]), .Z(n14820) );
  XOR U14797 ( .A(n14969), .B(n14970), .Z(n14965) );
  AND U14798 ( .A(n14971), .B(n14972), .Z(n14970) );
  XNOR U14799 ( .A(p_input[2132]), .B(n14969), .Z(n14972) );
  XNOR U14800 ( .A(n14969), .B(n14829), .Z(n14971) );
  IV U14801 ( .A(p_input[2116]), .Z(n14829) );
  XOR U14802 ( .A(n14973), .B(n14974), .Z(n14969) );
  AND U14803 ( .A(n14975), .B(n14976), .Z(n14974) );
  XNOR U14804 ( .A(p_input[2131]), .B(n14973), .Z(n14976) );
  XNOR U14805 ( .A(n14973), .B(n14838), .Z(n14975) );
  IV U14806 ( .A(p_input[2115]), .Z(n14838) );
  XOR U14807 ( .A(n14977), .B(n14978), .Z(n14973) );
  AND U14808 ( .A(n14979), .B(n14980), .Z(n14978) );
  XNOR U14809 ( .A(p_input[2130]), .B(n14977), .Z(n14980) );
  XNOR U14810 ( .A(n14977), .B(n14847), .Z(n14979) );
  IV U14811 ( .A(p_input[2114]), .Z(n14847) );
  XNOR U14812 ( .A(n14981), .B(n14982), .Z(n14977) );
  AND U14813 ( .A(n14983), .B(n14984), .Z(n14982) );
  XOR U14814 ( .A(p_input[2129]), .B(n14981), .Z(n14984) );
  XNOR U14815 ( .A(p_input[2113]), .B(n14981), .Z(n14983) );
  AND U14816 ( .A(p_input[2128]), .B(n14985), .Z(n14981) );
  IV U14817 ( .A(p_input[2112]), .Z(n14985) );
  XOR U14818 ( .A(n14986), .B(n14987), .Z(n14544) );
  AND U14819 ( .A(n460), .B(n14988), .Z(n14987) );
  XNOR U14820 ( .A(n14989), .B(n14986), .Z(n14988) );
  XOR U14821 ( .A(n14990), .B(n14991), .Z(n460) );
  AND U14822 ( .A(n14992), .B(n14993), .Z(n14991) );
  XNOR U14823 ( .A(n14555), .B(n14990), .Z(n14993) );
  AND U14824 ( .A(p_input[2111]), .B(p_input[2095]), .Z(n14555) );
  XOR U14825 ( .A(n14990), .B(n14554), .Z(n14992) );
  AND U14826 ( .A(p_input[2063]), .B(p_input[2079]), .Z(n14554) );
  XOR U14827 ( .A(n14994), .B(n14995), .Z(n14990) );
  AND U14828 ( .A(n14996), .B(n14997), .Z(n14995) );
  XOR U14829 ( .A(n14994), .B(n14567), .Z(n14997) );
  XNOR U14830 ( .A(p_input[2094]), .B(n14998), .Z(n14567) );
  AND U14831 ( .A(n335), .B(n14999), .Z(n14998) );
  XOR U14832 ( .A(p_input[2110]), .B(p_input[2094]), .Z(n14999) );
  XNOR U14833 ( .A(n14564), .B(n14994), .Z(n14996) );
  XOR U14834 ( .A(n15000), .B(n15001), .Z(n14564) );
  AND U14835 ( .A(n332), .B(n15002), .Z(n15001) );
  XOR U14836 ( .A(p_input[2078]), .B(p_input[2062]), .Z(n15002) );
  XOR U14837 ( .A(n15003), .B(n15004), .Z(n14994) );
  AND U14838 ( .A(n15005), .B(n15006), .Z(n15004) );
  XOR U14839 ( .A(n15003), .B(n14579), .Z(n15006) );
  XNOR U14840 ( .A(p_input[2093]), .B(n15007), .Z(n14579) );
  AND U14841 ( .A(n335), .B(n15008), .Z(n15007) );
  XOR U14842 ( .A(p_input[2109]), .B(p_input[2093]), .Z(n15008) );
  XNOR U14843 ( .A(n14576), .B(n15003), .Z(n15005) );
  XOR U14844 ( .A(n15009), .B(n15010), .Z(n14576) );
  AND U14845 ( .A(n332), .B(n15011), .Z(n15010) );
  XOR U14846 ( .A(p_input[2077]), .B(p_input[2061]), .Z(n15011) );
  XOR U14847 ( .A(n15012), .B(n15013), .Z(n15003) );
  AND U14848 ( .A(n15014), .B(n15015), .Z(n15013) );
  XOR U14849 ( .A(n15012), .B(n14591), .Z(n15015) );
  XNOR U14850 ( .A(p_input[2092]), .B(n15016), .Z(n14591) );
  AND U14851 ( .A(n335), .B(n15017), .Z(n15016) );
  XOR U14852 ( .A(p_input[2108]), .B(p_input[2092]), .Z(n15017) );
  XNOR U14853 ( .A(n14588), .B(n15012), .Z(n15014) );
  XOR U14854 ( .A(n15018), .B(n15019), .Z(n14588) );
  AND U14855 ( .A(n332), .B(n15020), .Z(n15019) );
  XOR U14856 ( .A(p_input[2076]), .B(p_input[2060]), .Z(n15020) );
  XOR U14857 ( .A(n15021), .B(n15022), .Z(n15012) );
  AND U14858 ( .A(n15023), .B(n15024), .Z(n15022) );
  XOR U14859 ( .A(n15021), .B(n14603), .Z(n15024) );
  XNOR U14860 ( .A(p_input[2091]), .B(n15025), .Z(n14603) );
  AND U14861 ( .A(n335), .B(n15026), .Z(n15025) );
  XOR U14862 ( .A(p_input[2107]), .B(p_input[2091]), .Z(n15026) );
  XNOR U14863 ( .A(n14600), .B(n15021), .Z(n15023) );
  XOR U14864 ( .A(n15027), .B(n15028), .Z(n14600) );
  AND U14865 ( .A(n332), .B(n15029), .Z(n15028) );
  XOR U14866 ( .A(p_input[2075]), .B(p_input[2059]), .Z(n15029) );
  XOR U14867 ( .A(n15030), .B(n15031), .Z(n15021) );
  AND U14868 ( .A(n15032), .B(n15033), .Z(n15031) );
  XOR U14869 ( .A(n15030), .B(n14615), .Z(n15033) );
  XNOR U14870 ( .A(p_input[2090]), .B(n15034), .Z(n14615) );
  AND U14871 ( .A(n335), .B(n15035), .Z(n15034) );
  XOR U14872 ( .A(p_input[2106]), .B(p_input[2090]), .Z(n15035) );
  XNOR U14873 ( .A(n14612), .B(n15030), .Z(n15032) );
  XOR U14874 ( .A(n15036), .B(n15037), .Z(n14612) );
  AND U14875 ( .A(n332), .B(n15038), .Z(n15037) );
  XOR U14876 ( .A(p_input[2074]), .B(p_input[2058]), .Z(n15038) );
  XOR U14877 ( .A(n15039), .B(n15040), .Z(n15030) );
  AND U14878 ( .A(n15041), .B(n15042), .Z(n15040) );
  XOR U14879 ( .A(n15039), .B(n14627), .Z(n15042) );
  XNOR U14880 ( .A(p_input[2089]), .B(n15043), .Z(n14627) );
  AND U14881 ( .A(n335), .B(n15044), .Z(n15043) );
  XOR U14882 ( .A(p_input[2105]), .B(p_input[2089]), .Z(n15044) );
  XNOR U14883 ( .A(n14624), .B(n15039), .Z(n15041) );
  XOR U14884 ( .A(n15045), .B(n15046), .Z(n14624) );
  AND U14885 ( .A(n332), .B(n15047), .Z(n15046) );
  XOR U14886 ( .A(p_input[2073]), .B(p_input[2057]), .Z(n15047) );
  XOR U14887 ( .A(n15048), .B(n15049), .Z(n15039) );
  AND U14888 ( .A(n15050), .B(n15051), .Z(n15049) );
  XOR U14889 ( .A(n15048), .B(n14639), .Z(n15051) );
  XNOR U14890 ( .A(p_input[2088]), .B(n15052), .Z(n14639) );
  AND U14891 ( .A(n335), .B(n15053), .Z(n15052) );
  XOR U14892 ( .A(p_input[2104]), .B(p_input[2088]), .Z(n15053) );
  XNOR U14893 ( .A(n14636), .B(n15048), .Z(n15050) );
  XOR U14894 ( .A(n15054), .B(n15055), .Z(n14636) );
  AND U14895 ( .A(n332), .B(n15056), .Z(n15055) );
  XOR U14896 ( .A(p_input[2072]), .B(p_input[2056]), .Z(n15056) );
  XOR U14897 ( .A(n15057), .B(n15058), .Z(n15048) );
  AND U14898 ( .A(n15059), .B(n15060), .Z(n15058) );
  XOR U14899 ( .A(n15057), .B(n14651), .Z(n15060) );
  XNOR U14900 ( .A(p_input[2087]), .B(n15061), .Z(n14651) );
  AND U14901 ( .A(n335), .B(n15062), .Z(n15061) );
  XOR U14902 ( .A(p_input[2103]), .B(p_input[2087]), .Z(n15062) );
  XNOR U14903 ( .A(n14648), .B(n15057), .Z(n15059) );
  XOR U14904 ( .A(n15063), .B(n15064), .Z(n14648) );
  AND U14905 ( .A(n332), .B(n15065), .Z(n15064) );
  XOR U14906 ( .A(p_input[2071]), .B(p_input[2055]), .Z(n15065) );
  XOR U14907 ( .A(n15066), .B(n15067), .Z(n15057) );
  AND U14908 ( .A(n15068), .B(n15069), .Z(n15067) );
  XOR U14909 ( .A(n15066), .B(n14663), .Z(n15069) );
  XNOR U14910 ( .A(p_input[2086]), .B(n15070), .Z(n14663) );
  AND U14911 ( .A(n335), .B(n15071), .Z(n15070) );
  XOR U14912 ( .A(p_input[2102]), .B(p_input[2086]), .Z(n15071) );
  XNOR U14913 ( .A(n14660), .B(n15066), .Z(n15068) );
  XOR U14914 ( .A(n15072), .B(n15073), .Z(n14660) );
  AND U14915 ( .A(n332), .B(n15074), .Z(n15073) );
  XOR U14916 ( .A(p_input[2070]), .B(p_input[2054]), .Z(n15074) );
  XOR U14917 ( .A(n15075), .B(n15076), .Z(n15066) );
  AND U14918 ( .A(n15077), .B(n15078), .Z(n15076) );
  XOR U14919 ( .A(n15075), .B(n14675), .Z(n15078) );
  XNOR U14920 ( .A(p_input[2085]), .B(n15079), .Z(n14675) );
  AND U14921 ( .A(n335), .B(n15080), .Z(n15079) );
  XOR U14922 ( .A(p_input[2101]), .B(p_input[2085]), .Z(n15080) );
  XNOR U14923 ( .A(n14672), .B(n15075), .Z(n15077) );
  XOR U14924 ( .A(n15081), .B(n15082), .Z(n14672) );
  AND U14925 ( .A(n332), .B(n15083), .Z(n15082) );
  XOR U14926 ( .A(p_input[2069]), .B(p_input[2053]), .Z(n15083) );
  XOR U14927 ( .A(n15084), .B(n15085), .Z(n15075) );
  AND U14928 ( .A(n15086), .B(n15087), .Z(n15085) );
  XOR U14929 ( .A(n15084), .B(n14687), .Z(n15087) );
  XNOR U14930 ( .A(p_input[2084]), .B(n15088), .Z(n14687) );
  AND U14931 ( .A(n335), .B(n15089), .Z(n15088) );
  XOR U14932 ( .A(p_input[2100]), .B(p_input[2084]), .Z(n15089) );
  XNOR U14933 ( .A(n14684), .B(n15084), .Z(n15086) );
  XOR U14934 ( .A(n15090), .B(n15091), .Z(n14684) );
  AND U14935 ( .A(n332), .B(n15092), .Z(n15091) );
  XOR U14936 ( .A(p_input[2068]), .B(p_input[2052]), .Z(n15092) );
  XOR U14937 ( .A(n15093), .B(n15094), .Z(n15084) );
  AND U14938 ( .A(n15095), .B(n15096), .Z(n15094) );
  XOR U14939 ( .A(n15093), .B(n14699), .Z(n15096) );
  XNOR U14940 ( .A(p_input[2083]), .B(n15097), .Z(n14699) );
  AND U14941 ( .A(n335), .B(n15098), .Z(n15097) );
  XOR U14942 ( .A(p_input[2099]), .B(p_input[2083]), .Z(n15098) );
  XNOR U14943 ( .A(n14696), .B(n15093), .Z(n15095) );
  XOR U14944 ( .A(n15099), .B(n15100), .Z(n14696) );
  AND U14945 ( .A(n332), .B(n15101), .Z(n15100) );
  XOR U14946 ( .A(p_input[2067]), .B(p_input[2051]), .Z(n15101) );
  XOR U14947 ( .A(n15102), .B(n15103), .Z(n15093) );
  AND U14948 ( .A(n15104), .B(n15105), .Z(n15103) );
  XOR U14949 ( .A(n15102), .B(n14711), .Z(n15105) );
  XNOR U14950 ( .A(p_input[2082]), .B(n15106), .Z(n14711) );
  AND U14951 ( .A(n335), .B(n15107), .Z(n15106) );
  XOR U14952 ( .A(p_input[2098]), .B(p_input[2082]), .Z(n15107) );
  XNOR U14953 ( .A(n14708), .B(n15102), .Z(n15104) );
  XOR U14954 ( .A(n15108), .B(n15109), .Z(n14708) );
  AND U14955 ( .A(n332), .B(n15110), .Z(n15109) );
  XOR U14956 ( .A(p_input[2066]), .B(p_input[2050]), .Z(n15110) );
  XOR U14957 ( .A(n15111), .B(n15112), .Z(n15102) );
  AND U14958 ( .A(n15113), .B(n15114), .Z(n15112) );
  XNOR U14959 ( .A(n15115), .B(n14724), .Z(n15114) );
  XNOR U14960 ( .A(p_input[2081]), .B(n15116), .Z(n14724) );
  AND U14961 ( .A(n335), .B(n15117), .Z(n15116) );
  XNOR U14962 ( .A(p_input[2097]), .B(n15118), .Z(n15117) );
  IV U14963 ( .A(p_input[2081]), .Z(n15118) );
  XNOR U14964 ( .A(n14721), .B(n15111), .Z(n15113) );
  XNOR U14965 ( .A(p_input[2049]), .B(n15119), .Z(n14721) );
  AND U14966 ( .A(n332), .B(n15120), .Z(n15119) );
  XOR U14967 ( .A(p_input[2065]), .B(p_input[2049]), .Z(n15120) );
  IV U14968 ( .A(n15115), .Z(n15111) );
  AND U14969 ( .A(n14986), .B(n14989), .Z(n15115) );
  XOR U14970 ( .A(p_input[2080]), .B(n15121), .Z(n14989) );
  AND U14971 ( .A(n335), .B(n15122), .Z(n15121) );
  XOR U14972 ( .A(p_input[2096]), .B(p_input[2080]), .Z(n15122) );
  XOR U14973 ( .A(n15123), .B(n15124), .Z(n335) );
  AND U14974 ( .A(n15125), .B(n15126), .Z(n15124) );
  XNOR U14975 ( .A(p_input[2111]), .B(n15123), .Z(n15126) );
  XOR U14976 ( .A(n15123), .B(p_input[2095]), .Z(n15125) );
  XOR U14977 ( .A(n15127), .B(n15128), .Z(n15123) );
  AND U14978 ( .A(n15129), .B(n15130), .Z(n15128) );
  XNOR U14979 ( .A(p_input[2110]), .B(n15127), .Z(n15130) );
  XOR U14980 ( .A(n15127), .B(p_input[2094]), .Z(n15129) );
  XOR U14981 ( .A(n15131), .B(n15132), .Z(n15127) );
  AND U14982 ( .A(n15133), .B(n15134), .Z(n15132) );
  XNOR U14983 ( .A(p_input[2109]), .B(n15131), .Z(n15134) );
  XOR U14984 ( .A(n15131), .B(p_input[2093]), .Z(n15133) );
  XOR U14985 ( .A(n15135), .B(n15136), .Z(n15131) );
  AND U14986 ( .A(n15137), .B(n15138), .Z(n15136) );
  XNOR U14987 ( .A(p_input[2108]), .B(n15135), .Z(n15138) );
  XOR U14988 ( .A(n15135), .B(p_input[2092]), .Z(n15137) );
  XOR U14989 ( .A(n15139), .B(n15140), .Z(n15135) );
  AND U14990 ( .A(n15141), .B(n15142), .Z(n15140) );
  XNOR U14991 ( .A(p_input[2107]), .B(n15139), .Z(n15142) );
  XOR U14992 ( .A(n15139), .B(p_input[2091]), .Z(n15141) );
  XOR U14993 ( .A(n15143), .B(n15144), .Z(n15139) );
  AND U14994 ( .A(n15145), .B(n15146), .Z(n15144) );
  XNOR U14995 ( .A(p_input[2106]), .B(n15143), .Z(n15146) );
  XOR U14996 ( .A(n15143), .B(p_input[2090]), .Z(n15145) );
  XOR U14997 ( .A(n15147), .B(n15148), .Z(n15143) );
  AND U14998 ( .A(n15149), .B(n15150), .Z(n15148) );
  XNOR U14999 ( .A(p_input[2105]), .B(n15147), .Z(n15150) );
  XOR U15000 ( .A(n15147), .B(p_input[2089]), .Z(n15149) );
  XOR U15001 ( .A(n15151), .B(n15152), .Z(n15147) );
  AND U15002 ( .A(n15153), .B(n15154), .Z(n15152) );
  XNOR U15003 ( .A(p_input[2104]), .B(n15151), .Z(n15154) );
  XOR U15004 ( .A(n15151), .B(p_input[2088]), .Z(n15153) );
  XOR U15005 ( .A(n15155), .B(n15156), .Z(n15151) );
  AND U15006 ( .A(n15157), .B(n15158), .Z(n15156) );
  XNOR U15007 ( .A(p_input[2103]), .B(n15155), .Z(n15158) );
  XOR U15008 ( .A(n15155), .B(p_input[2087]), .Z(n15157) );
  XOR U15009 ( .A(n15159), .B(n15160), .Z(n15155) );
  AND U15010 ( .A(n15161), .B(n15162), .Z(n15160) );
  XNOR U15011 ( .A(p_input[2102]), .B(n15159), .Z(n15162) );
  XOR U15012 ( .A(n15159), .B(p_input[2086]), .Z(n15161) );
  XOR U15013 ( .A(n15163), .B(n15164), .Z(n15159) );
  AND U15014 ( .A(n15165), .B(n15166), .Z(n15164) );
  XNOR U15015 ( .A(p_input[2101]), .B(n15163), .Z(n15166) );
  XOR U15016 ( .A(n15163), .B(p_input[2085]), .Z(n15165) );
  XOR U15017 ( .A(n15167), .B(n15168), .Z(n15163) );
  AND U15018 ( .A(n15169), .B(n15170), .Z(n15168) );
  XNOR U15019 ( .A(p_input[2100]), .B(n15167), .Z(n15170) );
  XOR U15020 ( .A(n15167), .B(p_input[2084]), .Z(n15169) );
  XOR U15021 ( .A(n15171), .B(n15172), .Z(n15167) );
  AND U15022 ( .A(n15173), .B(n15174), .Z(n15172) );
  XNOR U15023 ( .A(p_input[2099]), .B(n15171), .Z(n15174) );
  XOR U15024 ( .A(n15171), .B(p_input[2083]), .Z(n15173) );
  XOR U15025 ( .A(n15175), .B(n15176), .Z(n15171) );
  AND U15026 ( .A(n15177), .B(n15178), .Z(n15176) );
  XNOR U15027 ( .A(p_input[2098]), .B(n15175), .Z(n15178) );
  XOR U15028 ( .A(n15175), .B(p_input[2082]), .Z(n15177) );
  XNOR U15029 ( .A(n15179), .B(n15180), .Z(n15175) );
  AND U15030 ( .A(n15181), .B(n15182), .Z(n15180) );
  XOR U15031 ( .A(p_input[2097]), .B(n15179), .Z(n15182) );
  XNOR U15032 ( .A(p_input[2081]), .B(n15179), .Z(n15181) );
  AND U15033 ( .A(p_input[2096]), .B(n15183), .Z(n15179) );
  IV U15034 ( .A(p_input[2080]), .Z(n15183) );
  XNOR U15035 ( .A(p_input[2048]), .B(n15184), .Z(n14986) );
  AND U15036 ( .A(n332), .B(n15185), .Z(n15184) );
  XOR U15037 ( .A(p_input[2064]), .B(p_input[2048]), .Z(n15185) );
  XOR U15038 ( .A(n15186), .B(n15187), .Z(n332) );
  AND U15039 ( .A(n15188), .B(n15189), .Z(n15187) );
  XNOR U15040 ( .A(p_input[2079]), .B(n15186), .Z(n15189) );
  XOR U15041 ( .A(n15186), .B(p_input[2063]), .Z(n15188) );
  XOR U15042 ( .A(n15190), .B(n15191), .Z(n15186) );
  AND U15043 ( .A(n15192), .B(n15193), .Z(n15191) );
  XNOR U15044 ( .A(p_input[2078]), .B(n15190), .Z(n15193) );
  XNOR U15045 ( .A(n15190), .B(n15000), .Z(n15192) );
  IV U15046 ( .A(p_input[2062]), .Z(n15000) );
  XOR U15047 ( .A(n15194), .B(n15195), .Z(n15190) );
  AND U15048 ( .A(n15196), .B(n15197), .Z(n15195) );
  XNOR U15049 ( .A(p_input[2077]), .B(n15194), .Z(n15197) );
  XNOR U15050 ( .A(n15194), .B(n15009), .Z(n15196) );
  IV U15051 ( .A(p_input[2061]), .Z(n15009) );
  XOR U15052 ( .A(n15198), .B(n15199), .Z(n15194) );
  AND U15053 ( .A(n15200), .B(n15201), .Z(n15199) );
  XNOR U15054 ( .A(p_input[2076]), .B(n15198), .Z(n15201) );
  XNOR U15055 ( .A(n15198), .B(n15018), .Z(n15200) );
  IV U15056 ( .A(p_input[2060]), .Z(n15018) );
  XOR U15057 ( .A(n15202), .B(n15203), .Z(n15198) );
  AND U15058 ( .A(n15204), .B(n15205), .Z(n15203) );
  XNOR U15059 ( .A(p_input[2075]), .B(n15202), .Z(n15205) );
  XNOR U15060 ( .A(n15202), .B(n15027), .Z(n15204) );
  IV U15061 ( .A(p_input[2059]), .Z(n15027) );
  XOR U15062 ( .A(n15206), .B(n15207), .Z(n15202) );
  AND U15063 ( .A(n15208), .B(n15209), .Z(n15207) );
  XNOR U15064 ( .A(p_input[2074]), .B(n15206), .Z(n15209) );
  XNOR U15065 ( .A(n15206), .B(n15036), .Z(n15208) );
  IV U15066 ( .A(p_input[2058]), .Z(n15036) );
  XOR U15067 ( .A(n15210), .B(n15211), .Z(n15206) );
  AND U15068 ( .A(n15212), .B(n15213), .Z(n15211) );
  XNOR U15069 ( .A(p_input[2073]), .B(n15210), .Z(n15213) );
  XNOR U15070 ( .A(n15210), .B(n15045), .Z(n15212) );
  IV U15071 ( .A(p_input[2057]), .Z(n15045) );
  XOR U15072 ( .A(n15214), .B(n15215), .Z(n15210) );
  AND U15073 ( .A(n15216), .B(n15217), .Z(n15215) );
  XNOR U15074 ( .A(p_input[2072]), .B(n15214), .Z(n15217) );
  XNOR U15075 ( .A(n15214), .B(n15054), .Z(n15216) );
  IV U15076 ( .A(p_input[2056]), .Z(n15054) );
  XOR U15077 ( .A(n15218), .B(n15219), .Z(n15214) );
  AND U15078 ( .A(n15220), .B(n15221), .Z(n15219) );
  XNOR U15079 ( .A(p_input[2071]), .B(n15218), .Z(n15221) );
  XNOR U15080 ( .A(n15218), .B(n15063), .Z(n15220) );
  IV U15081 ( .A(p_input[2055]), .Z(n15063) );
  XOR U15082 ( .A(n15222), .B(n15223), .Z(n15218) );
  AND U15083 ( .A(n15224), .B(n15225), .Z(n15223) );
  XNOR U15084 ( .A(p_input[2070]), .B(n15222), .Z(n15225) );
  XNOR U15085 ( .A(n15222), .B(n15072), .Z(n15224) );
  IV U15086 ( .A(p_input[2054]), .Z(n15072) );
  XOR U15087 ( .A(n15226), .B(n15227), .Z(n15222) );
  AND U15088 ( .A(n15228), .B(n15229), .Z(n15227) );
  XNOR U15089 ( .A(p_input[2069]), .B(n15226), .Z(n15229) );
  XNOR U15090 ( .A(n15226), .B(n15081), .Z(n15228) );
  IV U15091 ( .A(p_input[2053]), .Z(n15081) );
  XOR U15092 ( .A(n15230), .B(n15231), .Z(n15226) );
  AND U15093 ( .A(n15232), .B(n15233), .Z(n15231) );
  XNOR U15094 ( .A(p_input[2068]), .B(n15230), .Z(n15233) );
  XNOR U15095 ( .A(n15230), .B(n15090), .Z(n15232) );
  IV U15096 ( .A(p_input[2052]), .Z(n15090) );
  XOR U15097 ( .A(n15234), .B(n15235), .Z(n15230) );
  AND U15098 ( .A(n15236), .B(n15237), .Z(n15235) );
  XNOR U15099 ( .A(p_input[2067]), .B(n15234), .Z(n15237) );
  XNOR U15100 ( .A(n15234), .B(n15099), .Z(n15236) );
  IV U15101 ( .A(p_input[2051]), .Z(n15099) );
  XOR U15102 ( .A(n15238), .B(n15239), .Z(n15234) );
  AND U15103 ( .A(n15240), .B(n15241), .Z(n15239) );
  XNOR U15104 ( .A(p_input[2066]), .B(n15238), .Z(n15241) );
  XNOR U15105 ( .A(n15238), .B(n15108), .Z(n15240) );
  IV U15106 ( .A(p_input[2050]), .Z(n15108) );
  XNOR U15107 ( .A(n15242), .B(n15243), .Z(n15238) );
  AND U15108 ( .A(n15244), .B(n15245), .Z(n15243) );
  XOR U15109 ( .A(p_input[2065]), .B(n15242), .Z(n15245) );
  XNOR U15110 ( .A(p_input[2049]), .B(n15242), .Z(n15244) );
  AND U15111 ( .A(p_input[2064]), .B(n15246), .Z(n15242) );
  IV U15112 ( .A(p_input[2048]), .Z(n15246) );
  XOR U15113 ( .A(n15247), .B(n15248), .Z(n7) );
  AND U15114 ( .A(n1060), .B(n15249), .Z(n15248) );
  XNOR U15115 ( .A(n15250), .B(n15247), .Z(n15249) );
  XOR U15116 ( .A(n15251), .B(n15252), .Z(n1060) );
  AND U15117 ( .A(n15253), .B(n15254), .Z(n15252) );
  XOR U15118 ( .A(n15251), .B(n1079), .Z(n15254) );
  XOR U15119 ( .A(n15255), .B(n15256), .Z(n1079) );
  AND U15120 ( .A(n1051), .B(n15257), .Z(n15256) );
  XOR U15121 ( .A(n15258), .B(n15255), .Z(n15257) );
  XNOR U15122 ( .A(n1076), .B(n15251), .Z(n15253) );
  XOR U15123 ( .A(n15259), .B(n15260), .Z(n1076) );
  AND U15124 ( .A(n1048), .B(n15261), .Z(n15260) );
  XOR U15125 ( .A(n15262), .B(n15259), .Z(n15261) );
  XOR U15126 ( .A(n15263), .B(n15264), .Z(n15251) );
  AND U15127 ( .A(n15265), .B(n15266), .Z(n15264) );
  XOR U15128 ( .A(n15263), .B(n1091), .Z(n15266) );
  XOR U15129 ( .A(n15267), .B(n15268), .Z(n1091) );
  AND U15130 ( .A(n1051), .B(n15269), .Z(n15268) );
  XOR U15131 ( .A(n15270), .B(n15267), .Z(n15269) );
  XNOR U15132 ( .A(n1088), .B(n15263), .Z(n15265) );
  XOR U15133 ( .A(n15271), .B(n15272), .Z(n1088) );
  AND U15134 ( .A(n1048), .B(n15273), .Z(n15272) );
  XOR U15135 ( .A(n15274), .B(n15271), .Z(n15273) );
  XOR U15136 ( .A(n15275), .B(n15276), .Z(n15263) );
  AND U15137 ( .A(n15277), .B(n15278), .Z(n15276) );
  XOR U15138 ( .A(n15275), .B(n1103), .Z(n15278) );
  XOR U15139 ( .A(n15279), .B(n15280), .Z(n1103) );
  AND U15140 ( .A(n1051), .B(n15281), .Z(n15280) );
  XOR U15141 ( .A(n15282), .B(n15279), .Z(n15281) );
  XNOR U15142 ( .A(n1100), .B(n15275), .Z(n15277) );
  XOR U15143 ( .A(n15283), .B(n15284), .Z(n1100) );
  AND U15144 ( .A(n1048), .B(n15285), .Z(n15284) );
  XOR U15145 ( .A(n15286), .B(n15283), .Z(n15285) );
  XOR U15146 ( .A(n15287), .B(n15288), .Z(n15275) );
  AND U15147 ( .A(n15289), .B(n15290), .Z(n15288) );
  XOR U15148 ( .A(n15287), .B(n1115), .Z(n15290) );
  XOR U15149 ( .A(n15291), .B(n15292), .Z(n1115) );
  AND U15150 ( .A(n1051), .B(n15293), .Z(n15292) );
  XOR U15151 ( .A(n15294), .B(n15291), .Z(n15293) );
  XNOR U15152 ( .A(n1112), .B(n15287), .Z(n15289) );
  XOR U15153 ( .A(n15295), .B(n15296), .Z(n1112) );
  AND U15154 ( .A(n1048), .B(n15297), .Z(n15296) );
  XOR U15155 ( .A(n15298), .B(n15295), .Z(n15297) );
  XOR U15156 ( .A(n15299), .B(n15300), .Z(n15287) );
  AND U15157 ( .A(n15301), .B(n15302), .Z(n15300) );
  XOR U15158 ( .A(n15299), .B(n1127), .Z(n15302) );
  XOR U15159 ( .A(n15303), .B(n15304), .Z(n1127) );
  AND U15160 ( .A(n1051), .B(n15305), .Z(n15304) );
  XOR U15161 ( .A(n15306), .B(n15303), .Z(n15305) );
  XNOR U15162 ( .A(n1124), .B(n15299), .Z(n15301) );
  XOR U15163 ( .A(n15307), .B(n15308), .Z(n1124) );
  AND U15164 ( .A(n1048), .B(n15309), .Z(n15308) );
  XOR U15165 ( .A(n15310), .B(n15307), .Z(n15309) );
  XOR U15166 ( .A(n15311), .B(n15312), .Z(n15299) );
  AND U15167 ( .A(n15313), .B(n15314), .Z(n15312) );
  XOR U15168 ( .A(n15311), .B(n1139), .Z(n15314) );
  XOR U15169 ( .A(n15315), .B(n15316), .Z(n1139) );
  AND U15170 ( .A(n1051), .B(n15317), .Z(n15316) );
  XOR U15171 ( .A(n15318), .B(n15315), .Z(n15317) );
  XNOR U15172 ( .A(n1136), .B(n15311), .Z(n15313) );
  XOR U15173 ( .A(n15319), .B(n15320), .Z(n1136) );
  AND U15174 ( .A(n1048), .B(n15321), .Z(n15320) );
  XOR U15175 ( .A(n15322), .B(n15319), .Z(n15321) );
  XOR U15176 ( .A(n15323), .B(n15324), .Z(n15311) );
  AND U15177 ( .A(n15325), .B(n15326), .Z(n15324) );
  XOR U15178 ( .A(n15323), .B(n1151), .Z(n15326) );
  XOR U15179 ( .A(n15327), .B(n15328), .Z(n1151) );
  AND U15180 ( .A(n1051), .B(n15329), .Z(n15328) );
  XOR U15181 ( .A(n15330), .B(n15327), .Z(n15329) );
  XNOR U15182 ( .A(n1148), .B(n15323), .Z(n15325) );
  XOR U15183 ( .A(n15331), .B(n15332), .Z(n1148) );
  AND U15184 ( .A(n1048), .B(n15333), .Z(n15332) );
  XOR U15185 ( .A(n15334), .B(n15331), .Z(n15333) );
  XOR U15186 ( .A(n15335), .B(n15336), .Z(n15323) );
  AND U15187 ( .A(n15337), .B(n15338), .Z(n15336) );
  XOR U15188 ( .A(n15335), .B(n1163), .Z(n15338) );
  XOR U15189 ( .A(n15339), .B(n15340), .Z(n1163) );
  AND U15190 ( .A(n1051), .B(n15341), .Z(n15340) );
  XOR U15191 ( .A(n15342), .B(n15339), .Z(n15341) );
  XNOR U15192 ( .A(n1160), .B(n15335), .Z(n15337) );
  XOR U15193 ( .A(n15343), .B(n15344), .Z(n1160) );
  AND U15194 ( .A(n1048), .B(n15345), .Z(n15344) );
  XOR U15195 ( .A(n15346), .B(n15343), .Z(n15345) );
  XOR U15196 ( .A(n15347), .B(n15348), .Z(n15335) );
  AND U15197 ( .A(n15349), .B(n15350), .Z(n15348) );
  XOR U15198 ( .A(n15347), .B(n1175), .Z(n15350) );
  XOR U15199 ( .A(n15351), .B(n15352), .Z(n1175) );
  AND U15200 ( .A(n1051), .B(n15353), .Z(n15352) );
  XOR U15201 ( .A(n15354), .B(n15351), .Z(n15353) );
  XNOR U15202 ( .A(n1172), .B(n15347), .Z(n15349) );
  XOR U15203 ( .A(n15355), .B(n15356), .Z(n1172) );
  AND U15204 ( .A(n1048), .B(n15357), .Z(n15356) );
  XOR U15205 ( .A(n15358), .B(n15355), .Z(n15357) );
  XOR U15206 ( .A(n15359), .B(n15360), .Z(n15347) );
  AND U15207 ( .A(n15361), .B(n15362), .Z(n15360) );
  XOR U15208 ( .A(n15359), .B(n1187), .Z(n15362) );
  XOR U15209 ( .A(n15363), .B(n15364), .Z(n1187) );
  AND U15210 ( .A(n1051), .B(n15365), .Z(n15364) );
  XOR U15211 ( .A(n15366), .B(n15363), .Z(n15365) );
  XNOR U15212 ( .A(n1184), .B(n15359), .Z(n15361) );
  XOR U15213 ( .A(n15367), .B(n15368), .Z(n1184) );
  AND U15214 ( .A(n1048), .B(n15369), .Z(n15368) );
  XOR U15215 ( .A(n15370), .B(n15367), .Z(n15369) );
  XOR U15216 ( .A(n15371), .B(n15372), .Z(n15359) );
  AND U15217 ( .A(n15373), .B(n15374), .Z(n15372) );
  XOR U15218 ( .A(n15371), .B(n1199), .Z(n15374) );
  XOR U15219 ( .A(n15375), .B(n15376), .Z(n1199) );
  AND U15220 ( .A(n1051), .B(n15377), .Z(n15376) );
  XOR U15221 ( .A(n15378), .B(n15375), .Z(n15377) );
  XNOR U15222 ( .A(n1196), .B(n15371), .Z(n15373) );
  XOR U15223 ( .A(n15379), .B(n15380), .Z(n1196) );
  AND U15224 ( .A(n1048), .B(n15381), .Z(n15380) );
  XOR U15225 ( .A(n15382), .B(n15379), .Z(n15381) );
  XOR U15226 ( .A(n15383), .B(n15384), .Z(n15371) );
  AND U15227 ( .A(n15385), .B(n15386), .Z(n15384) );
  XOR U15228 ( .A(n15383), .B(n1211), .Z(n15386) );
  XOR U15229 ( .A(n15387), .B(n15388), .Z(n1211) );
  AND U15230 ( .A(n1051), .B(n15389), .Z(n15388) );
  XOR U15231 ( .A(n15390), .B(n15387), .Z(n15389) );
  XNOR U15232 ( .A(n1208), .B(n15383), .Z(n15385) );
  XOR U15233 ( .A(n15391), .B(n15392), .Z(n1208) );
  AND U15234 ( .A(n1048), .B(n15393), .Z(n15392) );
  XOR U15235 ( .A(n15394), .B(n15391), .Z(n15393) );
  XOR U15236 ( .A(n15395), .B(n15396), .Z(n15383) );
  AND U15237 ( .A(n15397), .B(n15398), .Z(n15396) );
  XOR U15238 ( .A(n15395), .B(n1223), .Z(n15398) );
  XOR U15239 ( .A(n15399), .B(n15400), .Z(n1223) );
  AND U15240 ( .A(n1051), .B(n15401), .Z(n15400) );
  XOR U15241 ( .A(n15402), .B(n15399), .Z(n15401) );
  XNOR U15242 ( .A(n1220), .B(n15395), .Z(n15397) );
  XOR U15243 ( .A(n15403), .B(n15404), .Z(n1220) );
  AND U15244 ( .A(n1048), .B(n15405), .Z(n15404) );
  XOR U15245 ( .A(n15406), .B(n15403), .Z(n15405) );
  XOR U15246 ( .A(n15407), .B(n15408), .Z(n15395) );
  AND U15247 ( .A(n15409), .B(n15410), .Z(n15408) );
  XOR U15248 ( .A(n15407), .B(n1235), .Z(n15410) );
  XOR U15249 ( .A(n15411), .B(n15412), .Z(n1235) );
  AND U15250 ( .A(n1051), .B(n15413), .Z(n15412) );
  XOR U15251 ( .A(n15414), .B(n15411), .Z(n15413) );
  XNOR U15252 ( .A(n1232), .B(n15407), .Z(n15409) );
  XOR U15253 ( .A(n15415), .B(n15416), .Z(n1232) );
  AND U15254 ( .A(n1048), .B(n15417), .Z(n15416) );
  XOR U15255 ( .A(n15418), .B(n15415), .Z(n15417) );
  XOR U15256 ( .A(n15419), .B(n15420), .Z(n15407) );
  AND U15257 ( .A(n15421), .B(n15422), .Z(n15420) );
  XNOR U15258 ( .A(n15423), .B(n1247), .Z(n15422) );
  XOR U15259 ( .A(n15424), .B(n15425), .Z(n1247) );
  AND U15260 ( .A(n1051), .B(n15426), .Z(n15425) );
  XOR U15261 ( .A(n15424), .B(n15427), .Z(n15426) );
  XNOR U15262 ( .A(n1244), .B(n15419), .Z(n15421) );
  XOR U15263 ( .A(n15428), .B(n15429), .Z(n1244) );
  AND U15264 ( .A(n1048), .B(n15430), .Z(n15429) );
  XOR U15265 ( .A(n15428), .B(n15431), .Z(n15430) );
  IV U15266 ( .A(n15423), .Z(n15419) );
  AND U15267 ( .A(n15247), .B(n15250), .Z(n15423) );
  XNOR U15268 ( .A(n15432), .B(n15433), .Z(n15250) );
  AND U15269 ( .A(n1051), .B(n15434), .Z(n15433) );
  XNOR U15270 ( .A(n15435), .B(n15432), .Z(n15434) );
  XOR U15271 ( .A(n15436), .B(n15437), .Z(n1051) );
  AND U15272 ( .A(n15438), .B(n15439), .Z(n15437) );
  XOR U15273 ( .A(n15436), .B(n15258), .Z(n15439) );
  XOR U15274 ( .A(n15440), .B(n15441), .Z(n15258) );
  AND U15275 ( .A(n1019), .B(n15442), .Z(n15441) );
  XOR U15276 ( .A(n15443), .B(n15440), .Z(n15442) );
  XNOR U15277 ( .A(n15255), .B(n15436), .Z(n15438) );
  XOR U15278 ( .A(n15444), .B(n15445), .Z(n15255) );
  AND U15279 ( .A(n1017), .B(n15446), .Z(n15445) );
  XOR U15280 ( .A(n15447), .B(n15444), .Z(n15446) );
  XOR U15281 ( .A(n15448), .B(n15449), .Z(n15436) );
  AND U15282 ( .A(n15450), .B(n15451), .Z(n15449) );
  XOR U15283 ( .A(n15448), .B(n15270), .Z(n15451) );
  XOR U15284 ( .A(n15452), .B(n15453), .Z(n15270) );
  AND U15285 ( .A(n1019), .B(n15454), .Z(n15453) );
  XOR U15286 ( .A(n15455), .B(n15452), .Z(n15454) );
  XNOR U15287 ( .A(n15267), .B(n15448), .Z(n15450) );
  XOR U15288 ( .A(n15456), .B(n15457), .Z(n15267) );
  AND U15289 ( .A(n1017), .B(n15458), .Z(n15457) );
  XOR U15290 ( .A(n15459), .B(n15456), .Z(n15458) );
  XOR U15291 ( .A(n15460), .B(n15461), .Z(n15448) );
  AND U15292 ( .A(n15462), .B(n15463), .Z(n15461) );
  XOR U15293 ( .A(n15460), .B(n15282), .Z(n15463) );
  XOR U15294 ( .A(n15464), .B(n15465), .Z(n15282) );
  AND U15295 ( .A(n1019), .B(n15466), .Z(n15465) );
  XOR U15296 ( .A(n15467), .B(n15464), .Z(n15466) );
  XNOR U15297 ( .A(n15279), .B(n15460), .Z(n15462) );
  XOR U15298 ( .A(n15468), .B(n15469), .Z(n15279) );
  AND U15299 ( .A(n1017), .B(n15470), .Z(n15469) );
  XOR U15300 ( .A(n15471), .B(n15468), .Z(n15470) );
  XOR U15301 ( .A(n15472), .B(n15473), .Z(n15460) );
  AND U15302 ( .A(n15474), .B(n15475), .Z(n15473) );
  XOR U15303 ( .A(n15472), .B(n15294), .Z(n15475) );
  XOR U15304 ( .A(n15476), .B(n15477), .Z(n15294) );
  AND U15305 ( .A(n1019), .B(n15478), .Z(n15477) );
  XOR U15306 ( .A(n15479), .B(n15476), .Z(n15478) );
  XNOR U15307 ( .A(n15291), .B(n15472), .Z(n15474) );
  XOR U15308 ( .A(n15480), .B(n15481), .Z(n15291) );
  AND U15309 ( .A(n1017), .B(n15482), .Z(n15481) );
  XOR U15310 ( .A(n15483), .B(n15480), .Z(n15482) );
  XOR U15311 ( .A(n15484), .B(n15485), .Z(n15472) );
  AND U15312 ( .A(n15486), .B(n15487), .Z(n15485) );
  XOR U15313 ( .A(n15484), .B(n15306), .Z(n15487) );
  XOR U15314 ( .A(n15488), .B(n15489), .Z(n15306) );
  AND U15315 ( .A(n1019), .B(n15490), .Z(n15489) );
  XOR U15316 ( .A(n15491), .B(n15488), .Z(n15490) );
  XNOR U15317 ( .A(n15303), .B(n15484), .Z(n15486) );
  XOR U15318 ( .A(n15492), .B(n15493), .Z(n15303) );
  AND U15319 ( .A(n1017), .B(n15494), .Z(n15493) );
  XOR U15320 ( .A(n15495), .B(n15492), .Z(n15494) );
  XOR U15321 ( .A(n15496), .B(n15497), .Z(n15484) );
  AND U15322 ( .A(n15498), .B(n15499), .Z(n15497) );
  XOR U15323 ( .A(n15496), .B(n15318), .Z(n15499) );
  XOR U15324 ( .A(n15500), .B(n15501), .Z(n15318) );
  AND U15325 ( .A(n1019), .B(n15502), .Z(n15501) );
  XOR U15326 ( .A(n15503), .B(n15500), .Z(n15502) );
  XNOR U15327 ( .A(n15315), .B(n15496), .Z(n15498) );
  XOR U15328 ( .A(n15504), .B(n15505), .Z(n15315) );
  AND U15329 ( .A(n1017), .B(n15506), .Z(n15505) );
  XOR U15330 ( .A(n15507), .B(n15504), .Z(n15506) );
  XOR U15331 ( .A(n15508), .B(n15509), .Z(n15496) );
  AND U15332 ( .A(n15510), .B(n15511), .Z(n15509) );
  XOR U15333 ( .A(n15508), .B(n15330), .Z(n15511) );
  XOR U15334 ( .A(n15512), .B(n15513), .Z(n15330) );
  AND U15335 ( .A(n1019), .B(n15514), .Z(n15513) );
  XOR U15336 ( .A(n15515), .B(n15512), .Z(n15514) );
  XNOR U15337 ( .A(n15327), .B(n15508), .Z(n15510) );
  XOR U15338 ( .A(n15516), .B(n15517), .Z(n15327) );
  AND U15339 ( .A(n1017), .B(n15518), .Z(n15517) );
  XOR U15340 ( .A(n15519), .B(n15516), .Z(n15518) );
  XOR U15341 ( .A(n15520), .B(n15521), .Z(n15508) );
  AND U15342 ( .A(n15522), .B(n15523), .Z(n15521) );
  XOR U15343 ( .A(n15520), .B(n15342), .Z(n15523) );
  XOR U15344 ( .A(n15524), .B(n15525), .Z(n15342) );
  AND U15345 ( .A(n1019), .B(n15526), .Z(n15525) );
  XOR U15346 ( .A(n15527), .B(n15524), .Z(n15526) );
  XNOR U15347 ( .A(n15339), .B(n15520), .Z(n15522) );
  XOR U15348 ( .A(n15528), .B(n15529), .Z(n15339) );
  AND U15349 ( .A(n1017), .B(n15530), .Z(n15529) );
  XOR U15350 ( .A(n15531), .B(n15528), .Z(n15530) );
  XOR U15351 ( .A(n15532), .B(n15533), .Z(n15520) );
  AND U15352 ( .A(n15534), .B(n15535), .Z(n15533) );
  XOR U15353 ( .A(n15532), .B(n15354), .Z(n15535) );
  XOR U15354 ( .A(n15536), .B(n15537), .Z(n15354) );
  AND U15355 ( .A(n1019), .B(n15538), .Z(n15537) );
  XOR U15356 ( .A(n15539), .B(n15536), .Z(n15538) );
  XNOR U15357 ( .A(n15351), .B(n15532), .Z(n15534) );
  XOR U15358 ( .A(n15540), .B(n15541), .Z(n15351) );
  AND U15359 ( .A(n1017), .B(n15542), .Z(n15541) );
  XOR U15360 ( .A(n15543), .B(n15540), .Z(n15542) );
  XOR U15361 ( .A(n15544), .B(n15545), .Z(n15532) );
  AND U15362 ( .A(n15546), .B(n15547), .Z(n15545) );
  XOR U15363 ( .A(n15544), .B(n15366), .Z(n15547) );
  XOR U15364 ( .A(n15548), .B(n15549), .Z(n15366) );
  AND U15365 ( .A(n1019), .B(n15550), .Z(n15549) );
  XOR U15366 ( .A(n15551), .B(n15548), .Z(n15550) );
  XNOR U15367 ( .A(n15363), .B(n15544), .Z(n15546) );
  XOR U15368 ( .A(n15552), .B(n15553), .Z(n15363) );
  AND U15369 ( .A(n1017), .B(n15554), .Z(n15553) );
  XOR U15370 ( .A(n15555), .B(n15552), .Z(n15554) );
  XOR U15371 ( .A(n15556), .B(n15557), .Z(n15544) );
  AND U15372 ( .A(n15558), .B(n15559), .Z(n15557) );
  XOR U15373 ( .A(n15556), .B(n15378), .Z(n15559) );
  XOR U15374 ( .A(n15560), .B(n15561), .Z(n15378) );
  AND U15375 ( .A(n1019), .B(n15562), .Z(n15561) );
  XOR U15376 ( .A(n15563), .B(n15560), .Z(n15562) );
  XNOR U15377 ( .A(n15375), .B(n15556), .Z(n15558) );
  XOR U15378 ( .A(n15564), .B(n15565), .Z(n15375) );
  AND U15379 ( .A(n1017), .B(n15566), .Z(n15565) );
  XOR U15380 ( .A(n15567), .B(n15564), .Z(n15566) );
  XOR U15381 ( .A(n15568), .B(n15569), .Z(n15556) );
  AND U15382 ( .A(n15570), .B(n15571), .Z(n15569) );
  XOR U15383 ( .A(n15568), .B(n15390), .Z(n15571) );
  XOR U15384 ( .A(n15572), .B(n15573), .Z(n15390) );
  AND U15385 ( .A(n1019), .B(n15574), .Z(n15573) );
  XOR U15386 ( .A(n15575), .B(n15572), .Z(n15574) );
  XNOR U15387 ( .A(n15387), .B(n15568), .Z(n15570) );
  XOR U15388 ( .A(n15576), .B(n15577), .Z(n15387) );
  AND U15389 ( .A(n1017), .B(n15578), .Z(n15577) );
  XOR U15390 ( .A(n15579), .B(n15576), .Z(n15578) );
  XOR U15391 ( .A(n15580), .B(n15581), .Z(n15568) );
  AND U15392 ( .A(n15582), .B(n15583), .Z(n15581) );
  XOR U15393 ( .A(n15580), .B(n15402), .Z(n15583) );
  XOR U15394 ( .A(n15584), .B(n15585), .Z(n15402) );
  AND U15395 ( .A(n1019), .B(n15586), .Z(n15585) );
  XOR U15396 ( .A(n15587), .B(n15584), .Z(n15586) );
  XNOR U15397 ( .A(n15399), .B(n15580), .Z(n15582) );
  XOR U15398 ( .A(n15588), .B(n15589), .Z(n15399) );
  AND U15399 ( .A(n1017), .B(n15590), .Z(n15589) );
  XOR U15400 ( .A(n15591), .B(n15588), .Z(n15590) );
  XOR U15401 ( .A(n15592), .B(n15593), .Z(n15580) );
  AND U15402 ( .A(n15594), .B(n15595), .Z(n15593) );
  XOR U15403 ( .A(n15592), .B(n15414), .Z(n15595) );
  XOR U15404 ( .A(n15596), .B(n15597), .Z(n15414) );
  AND U15405 ( .A(n1019), .B(n15598), .Z(n15597) );
  XOR U15406 ( .A(n15599), .B(n15596), .Z(n15598) );
  XNOR U15407 ( .A(n15411), .B(n15592), .Z(n15594) );
  XOR U15408 ( .A(n15600), .B(n15601), .Z(n15411) );
  AND U15409 ( .A(n1017), .B(n15602), .Z(n15601) );
  XOR U15410 ( .A(n15603), .B(n15600), .Z(n15602) );
  XOR U15411 ( .A(n15604), .B(n15605), .Z(n15592) );
  AND U15412 ( .A(n15606), .B(n15607), .Z(n15605) );
  XNOR U15413 ( .A(n15608), .B(n15427), .Z(n15607) );
  XOR U15414 ( .A(n15609), .B(n15610), .Z(n15427) );
  AND U15415 ( .A(n1019), .B(n15611), .Z(n15610) );
  XOR U15416 ( .A(n15609), .B(n15612), .Z(n15611) );
  XNOR U15417 ( .A(n15424), .B(n15604), .Z(n15606) );
  XOR U15418 ( .A(n15613), .B(n15614), .Z(n15424) );
  AND U15419 ( .A(n1017), .B(n15615), .Z(n15614) );
  XOR U15420 ( .A(n15613), .B(n15616), .Z(n15615) );
  IV U15421 ( .A(n15608), .Z(n15604) );
  AND U15422 ( .A(n15432), .B(n15435), .Z(n15608) );
  XNOR U15423 ( .A(n15617), .B(n15618), .Z(n15435) );
  AND U15424 ( .A(n1019), .B(n15619), .Z(n15618) );
  XNOR U15425 ( .A(n15620), .B(n15617), .Z(n15619) );
  XOR U15426 ( .A(n15621), .B(n15622), .Z(n1019) );
  AND U15427 ( .A(n15623), .B(n15624), .Z(n15622) );
  XOR U15428 ( .A(n15621), .B(n15443), .Z(n15624) );
  XNOR U15429 ( .A(n15625), .B(n15626), .Z(n15443) );
  AND U15430 ( .A(n15627), .B(n947), .Z(n15626) );
  AND U15431 ( .A(n15625), .B(n15628), .Z(n15627) );
  XNOR U15432 ( .A(n15440), .B(n15621), .Z(n15623) );
  XOR U15433 ( .A(n15629), .B(n15630), .Z(n15440) );
  AND U15434 ( .A(n15631), .B(n945), .Z(n15630) );
  NOR U15435 ( .A(n15629), .B(n15632), .Z(n15631) );
  XOR U15436 ( .A(n15633), .B(n15634), .Z(n15621) );
  AND U15437 ( .A(n15635), .B(n15636), .Z(n15634) );
  XOR U15438 ( .A(n15633), .B(n15455), .Z(n15636) );
  XOR U15439 ( .A(n15637), .B(n15638), .Z(n15455) );
  AND U15440 ( .A(n947), .B(n15639), .Z(n15638) );
  XOR U15441 ( .A(n15640), .B(n15637), .Z(n15639) );
  XNOR U15442 ( .A(n15452), .B(n15633), .Z(n15635) );
  XOR U15443 ( .A(n15641), .B(n15642), .Z(n15452) );
  AND U15444 ( .A(n945), .B(n15643), .Z(n15642) );
  XOR U15445 ( .A(n15644), .B(n15641), .Z(n15643) );
  XOR U15446 ( .A(n15645), .B(n15646), .Z(n15633) );
  AND U15447 ( .A(n15647), .B(n15648), .Z(n15646) );
  XOR U15448 ( .A(n15645), .B(n15467), .Z(n15648) );
  XOR U15449 ( .A(n15649), .B(n15650), .Z(n15467) );
  AND U15450 ( .A(n947), .B(n15651), .Z(n15650) );
  XOR U15451 ( .A(n15652), .B(n15649), .Z(n15651) );
  XNOR U15452 ( .A(n15464), .B(n15645), .Z(n15647) );
  XOR U15453 ( .A(n15653), .B(n15654), .Z(n15464) );
  AND U15454 ( .A(n945), .B(n15655), .Z(n15654) );
  XOR U15455 ( .A(n15656), .B(n15653), .Z(n15655) );
  XOR U15456 ( .A(n15657), .B(n15658), .Z(n15645) );
  AND U15457 ( .A(n15659), .B(n15660), .Z(n15658) );
  XOR U15458 ( .A(n15657), .B(n15479), .Z(n15660) );
  XOR U15459 ( .A(n15661), .B(n15662), .Z(n15479) );
  AND U15460 ( .A(n947), .B(n15663), .Z(n15662) );
  XOR U15461 ( .A(n15664), .B(n15661), .Z(n15663) );
  XNOR U15462 ( .A(n15476), .B(n15657), .Z(n15659) );
  XOR U15463 ( .A(n15665), .B(n15666), .Z(n15476) );
  AND U15464 ( .A(n945), .B(n15667), .Z(n15666) );
  XOR U15465 ( .A(n15668), .B(n15665), .Z(n15667) );
  XOR U15466 ( .A(n15669), .B(n15670), .Z(n15657) );
  AND U15467 ( .A(n15671), .B(n15672), .Z(n15670) );
  XOR U15468 ( .A(n15669), .B(n15491), .Z(n15672) );
  XOR U15469 ( .A(n15673), .B(n15674), .Z(n15491) );
  AND U15470 ( .A(n947), .B(n15675), .Z(n15674) );
  XOR U15471 ( .A(n15676), .B(n15673), .Z(n15675) );
  XNOR U15472 ( .A(n15488), .B(n15669), .Z(n15671) );
  XOR U15473 ( .A(n15677), .B(n15678), .Z(n15488) );
  AND U15474 ( .A(n945), .B(n15679), .Z(n15678) );
  XOR U15475 ( .A(n15680), .B(n15677), .Z(n15679) );
  XOR U15476 ( .A(n15681), .B(n15682), .Z(n15669) );
  AND U15477 ( .A(n15683), .B(n15684), .Z(n15682) );
  XOR U15478 ( .A(n15681), .B(n15503), .Z(n15684) );
  XOR U15479 ( .A(n15685), .B(n15686), .Z(n15503) );
  AND U15480 ( .A(n947), .B(n15687), .Z(n15686) );
  XOR U15481 ( .A(n15688), .B(n15685), .Z(n15687) );
  XNOR U15482 ( .A(n15500), .B(n15681), .Z(n15683) );
  XOR U15483 ( .A(n15689), .B(n15690), .Z(n15500) );
  AND U15484 ( .A(n945), .B(n15691), .Z(n15690) );
  XOR U15485 ( .A(n15692), .B(n15689), .Z(n15691) );
  XOR U15486 ( .A(n15693), .B(n15694), .Z(n15681) );
  AND U15487 ( .A(n15695), .B(n15696), .Z(n15694) );
  XOR U15488 ( .A(n15693), .B(n15515), .Z(n15696) );
  XOR U15489 ( .A(n15697), .B(n15698), .Z(n15515) );
  AND U15490 ( .A(n947), .B(n15699), .Z(n15698) );
  XOR U15491 ( .A(n15700), .B(n15697), .Z(n15699) );
  XNOR U15492 ( .A(n15512), .B(n15693), .Z(n15695) );
  XOR U15493 ( .A(n15701), .B(n15702), .Z(n15512) );
  AND U15494 ( .A(n945), .B(n15703), .Z(n15702) );
  XOR U15495 ( .A(n15704), .B(n15701), .Z(n15703) );
  XOR U15496 ( .A(n15705), .B(n15706), .Z(n15693) );
  AND U15497 ( .A(n15707), .B(n15708), .Z(n15706) );
  XOR U15498 ( .A(n15705), .B(n15527), .Z(n15708) );
  XOR U15499 ( .A(n15709), .B(n15710), .Z(n15527) );
  AND U15500 ( .A(n947), .B(n15711), .Z(n15710) );
  XOR U15501 ( .A(n15712), .B(n15709), .Z(n15711) );
  XNOR U15502 ( .A(n15524), .B(n15705), .Z(n15707) );
  XOR U15503 ( .A(n15713), .B(n15714), .Z(n15524) );
  AND U15504 ( .A(n945), .B(n15715), .Z(n15714) );
  XOR U15505 ( .A(n15716), .B(n15713), .Z(n15715) );
  XOR U15506 ( .A(n15717), .B(n15718), .Z(n15705) );
  AND U15507 ( .A(n15719), .B(n15720), .Z(n15718) );
  XOR U15508 ( .A(n15717), .B(n15539), .Z(n15720) );
  XOR U15509 ( .A(n15721), .B(n15722), .Z(n15539) );
  AND U15510 ( .A(n947), .B(n15723), .Z(n15722) );
  XOR U15511 ( .A(n15724), .B(n15721), .Z(n15723) );
  XNOR U15512 ( .A(n15536), .B(n15717), .Z(n15719) );
  XOR U15513 ( .A(n15725), .B(n15726), .Z(n15536) );
  AND U15514 ( .A(n945), .B(n15727), .Z(n15726) );
  XOR U15515 ( .A(n15728), .B(n15725), .Z(n15727) );
  XOR U15516 ( .A(n15729), .B(n15730), .Z(n15717) );
  AND U15517 ( .A(n15731), .B(n15732), .Z(n15730) );
  XOR U15518 ( .A(n15729), .B(n15551), .Z(n15732) );
  XOR U15519 ( .A(n15733), .B(n15734), .Z(n15551) );
  AND U15520 ( .A(n947), .B(n15735), .Z(n15734) );
  XOR U15521 ( .A(n15736), .B(n15733), .Z(n15735) );
  XNOR U15522 ( .A(n15548), .B(n15729), .Z(n15731) );
  XOR U15523 ( .A(n15737), .B(n15738), .Z(n15548) );
  AND U15524 ( .A(n945), .B(n15739), .Z(n15738) );
  XOR U15525 ( .A(n15740), .B(n15737), .Z(n15739) );
  XOR U15526 ( .A(n15741), .B(n15742), .Z(n15729) );
  AND U15527 ( .A(n15743), .B(n15744), .Z(n15742) );
  XOR U15528 ( .A(n15741), .B(n15563), .Z(n15744) );
  XOR U15529 ( .A(n15745), .B(n15746), .Z(n15563) );
  AND U15530 ( .A(n947), .B(n15747), .Z(n15746) );
  XOR U15531 ( .A(n15748), .B(n15745), .Z(n15747) );
  XNOR U15532 ( .A(n15560), .B(n15741), .Z(n15743) );
  XOR U15533 ( .A(n15749), .B(n15750), .Z(n15560) );
  AND U15534 ( .A(n945), .B(n15751), .Z(n15750) );
  XOR U15535 ( .A(n15752), .B(n15749), .Z(n15751) );
  XOR U15536 ( .A(n15753), .B(n15754), .Z(n15741) );
  AND U15537 ( .A(n15755), .B(n15756), .Z(n15754) );
  XOR U15538 ( .A(n15753), .B(n15575), .Z(n15756) );
  XOR U15539 ( .A(n15757), .B(n15758), .Z(n15575) );
  AND U15540 ( .A(n947), .B(n15759), .Z(n15758) );
  XOR U15541 ( .A(n15760), .B(n15757), .Z(n15759) );
  XNOR U15542 ( .A(n15572), .B(n15753), .Z(n15755) );
  XOR U15543 ( .A(n15761), .B(n15762), .Z(n15572) );
  AND U15544 ( .A(n945), .B(n15763), .Z(n15762) );
  XOR U15545 ( .A(n15764), .B(n15761), .Z(n15763) );
  XOR U15546 ( .A(n15765), .B(n15766), .Z(n15753) );
  AND U15547 ( .A(n15767), .B(n15768), .Z(n15766) );
  XOR U15548 ( .A(n15765), .B(n15587), .Z(n15768) );
  XOR U15549 ( .A(n15769), .B(n15770), .Z(n15587) );
  AND U15550 ( .A(n947), .B(n15771), .Z(n15770) );
  XOR U15551 ( .A(n15772), .B(n15769), .Z(n15771) );
  XNOR U15552 ( .A(n15584), .B(n15765), .Z(n15767) );
  XOR U15553 ( .A(n15773), .B(n15774), .Z(n15584) );
  AND U15554 ( .A(n945), .B(n15775), .Z(n15774) );
  XOR U15555 ( .A(n15776), .B(n15773), .Z(n15775) );
  XOR U15556 ( .A(n15777), .B(n15778), .Z(n15765) );
  AND U15557 ( .A(n15779), .B(n15780), .Z(n15778) );
  XOR U15558 ( .A(n15777), .B(n15599), .Z(n15780) );
  XOR U15559 ( .A(n15781), .B(n15782), .Z(n15599) );
  AND U15560 ( .A(n947), .B(n15783), .Z(n15782) );
  XOR U15561 ( .A(n15784), .B(n15781), .Z(n15783) );
  XNOR U15562 ( .A(n15596), .B(n15777), .Z(n15779) );
  XOR U15563 ( .A(n15785), .B(n15786), .Z(n15596) );
  AND U15564 ( .A(n945), .B(n15787), .Z(n15786) );
  XOR U15565 ( .A(n15788), .B(n15785), .Z(n15787) );
  XOR U15566 ( .A(n15789), .B(n15790), .Z(n15777) );
  AND U15567 ( .A(n15791), .B(n15792), .Z(n15790) );
  XNOR U15568 ( .A(n15793), .B(n15612), .Z(n15792) );
  XOR U15569 ( .A(n15794), .B(n15795), .Z(n15612) );
  AND U15570 ( .A(n947), .B(n15796), .Z(n15795) );
  XOR U15571 ( .A(n15794), .B(n15797), .Z(n15796) );
  XNOR U15572 ( .A(n15609), .B(n15789), .Z(n15791) );
  XOR U15573 ( .A(n15798), .B(n15799), .Z(n15609) );
  AND U15574 ( .A(n945), .B(n15800), .Z(n15799) );
  XOR U15575 ( .A(n15798), .B(n15801), .Z(n15800) );
  IV U15576 ( .A(n15793), .Z(n15789) );
  AND U15577 ( .A(n15617), .B(n15620), .Z(n15793) );
  XNOR U15578 ( .A(n15802), .B(n15803), .Z(n15620) );
  AND U15579 ( .A(n947), .B(n15804), .Z(n15803) );
  XNOR U15580 ( .A(n15805), .B(n15802), .Z(n15804) );
  XOR U15581 ( .A(n15806), .B(n15807), .Z(n947) );
  AND U15582 ( .A(n15808), .B(n15809), .Z(n15807) );
  XOR U15583 ( .A(n15628), .B(n15806), .Z(n15809) );
  IV U15584 ( .A(n15810), .Z(n15628) );
  AND U15585 ( .A(n15811), .B(n15812), .Z(n15810) );
  XOR U15586 ( .A(n15806), .B(n15625), .Z(n15808) );
  AND U15587 ( .A(n15813), .B(n15814), .Z(n15625) );
  XOR U15588 ( .A(n15815), .B(n15816), .Z(n15806) );
  AND U15589 ( .A(n15817), .B(n15818), .Z(n15816) );
  XOR U15590 ( .A(n15815), .B(n15640), .Z(n15818) );
  XOR U15591 ( .A(n15819), .B(n15820), .Z(n15640) );
  AND U15592 ( .A(n795), .B(n15821), .Z(n15820) );
  XOR U15593 ( .A(n15822), .B(n15819), .Z(n15821) );
  XNOR U15594 ( .A(n15637), .B(n15815), .Z(n15817) );
  XOR U15595 ( .A(n15823), .B(n15824), .Z(n15637) );
  AND U15596 ( .A(n793), .B(n15825), .Z(n15824) );
  XOR U15597 ( .A(n15826), .B(n15823), .Z(n15825) );
  XOR U15598 ( .A(n15827), .B(n15828), .Z(n15815) );
  AND U15599 ( .A(n15829), .B(n15830), .Z(n15828) );
  XOR U15600 ( .A(n15827), .B(n15652), .Z(n15830) );
  XOR U15601 ( .A(n15831), .B(n15832), .Z(n15652) );
  AND U15602 ( .A(n795), .B(n15833), .Z(n15832) );
  XOR U15603 ( .A(n15834), .B(n15831), .Z(n15833) );
  XNOR U15604 ( .A(n15649), .B(n15827), .Z(n15829) );
  XOR U15605 ( .A(n15835), .B(n15836), .Z(n15649) );
  AND U15606 ( .A(n793), .B(n15837), .Z(n15836) );
  XOR U15607 ( .A(n15838), .B(n15835), .Z(n15837) );
  XOR U15608 ( .A(n15839), .B(n15840), .Z(n15827) );
  AND U15609 ( .A(n15841), .B(n15842), .Z(n15840) );
  XOR U15610 ( .A(n15839), .B(n15664), .Z(n15842) );
  XOR U15611 ( .A(n15843), .B(n15844), .Z(n15664) );
  AND U15612 ( .A(n795), .B(n15845), .Z(n15844) );
  XOR U15613 ( .A(n15846), .B(n15843), .Z(n15845) );
  XNOR U15614 ( .A(n15661), .B(n15839), .Z(n15841) );
  XOR U15615 ( .A(n15847), .B(n15848), .Z(n15661) );
  AND U15616 ( .A(n793), .B(n15849), .Z(n15848) );
  XOR U15617 ( .A(n15850), .B(n15847), .Z(n15849) );
  XOR U15618 ( .A(n15851), .B(n15852), .Z(n15839) );
  AND U15619 ( .A(n15853), .B(n15854), .Z(n15852) );
  XOR U15620 ( .A(n15851), .B(n15676), .Z(n15854) );
  XOR U15621 ( .A(n15855), .B(n15856), .Z(n15676) );
  AND U15622 ( .A(n795), .B(n15857), .Z(n15856) );
  XOR U15623 ( .A(n15858), .B(n15855), .Z(n15857) );
  XNOR U15624 ( .A(n15673), .B(n15851), .Z(n15853) );
  XOR U15625 ( .A(n15859), .B(n15860), .Z(n15673) );
  AND U15626 ( .A(n793), .B(n15861), .Z(n15860) );
  XOR U15627 ( .A(n15862), .B(n15859), .Z(n15861) );
  XOR U15628 ( .A(n15863), .B(n15864), .Z(n15851) );
  AND U15629 ( .A(n15865), .B(n15866), .Z(n15864) );
  XOR U15630 ( .A(n15863), .B(n15688), .Z(n15866) );
  XOR U15631 ( .A(n15867), .B(n15868), .Z(n15688) );
  AND U15632 ( .A(n795), .B(n15869), .Z(n15868) );
  XOR U15633 ( .A(n15870), .B(n15867), .Z(n15869) );
  XNOR U15634 ( .A(n15685), .B(n15863), .Z(n15865) );
  XOR U15635 ( .A(n15871), .B(n15872), .Z(n15685) );
  AND U15636 ( .A(n793), .B(n15873), .Z(n15872) );
  XOR U15637 ( .A(n15874), .B(n15871), .Z(n15873) );
  XOR U15638 ( .A(n15875), .B(n15876), .Z(n15863) );
  AND U15639 ( .A(n15877), .B(n15878), .Z(n15876) );
  XOR U15640 ( .A(n15875), .B(n15700), .Z(n15878) );
  XOR U15641 ( .A(n15879), .B(n15880), .Z(n15700) );
  AND U15642 ( .A(n795), .B(n15881), .Z(n15880) );
  XOR U15643 ( .A(n15882), .B(n15879), .Z(n15881) );
  XNOR U15644 ( .A(n15697), .B(n15875), .Z(n15877) );
  XOR U15645 ( .A(n15883), .B(n15884), .Z(n15697) );
  AND U15646 ( .A(n793), .B(n15885), .Z(n15884) );
  XOR U15647 ( .A(n15886), .B(n15883), .Z(n15885) );
  XOR U15648 ( .A(n15887), .B(n15888), .Z(n15875) );
  AND U15649 ( .A(n15889), .B(n15890), .Z(n15888) );
  XOR U15650 ( .A(n15887), .B(n15712), .Z(n15890) );
  XOR U15651 ( .A(n15891), .B(n15892), .Z(n15712) );
  AND U15652 ( .A(n795), .B(n15893), .Z(n15892) );
  XOR U15653 ( .A(n15894), .B(n15891), .Z(n15893) );
  XNOR U15654 ( .A(n15709), .B(n15887), .Z(n15889) );
  XOR U15655 ( .A(n15895), .B(n15896), .Z(n15709) );
  AND U15656 ( .A(n793), .B(n15897), .Z(n15896) );
  XOR U15657 ( .A(n15898), .B(n15895), .Z(n15897) );
  XOR U15658 ( .A(n15899), .B(n15900), .Z(n15887) );
  AND U15659 ( .A(n15901), .B(n15902), .Z(n15900) );
  XOR U15660 ( .A(n15899), .B(n15724), .Z(n15902) );
  XOR U15661 ( .A(n15903), .B(n15904), .Z(n15724) );
  AND U15662 ( .A(n795), .B(n15905), .Z(n15904) );
  XOR U15663 ( .A(n15906), .B(n15903), .Z(n15905) );
  XNOR U15664 ( .A(n15721), .B(n15899), .Z(n15901) );
  XOR U15665 ( .A(n15907), .B(n15908), .Z(n15721) );
  AND U15666 ( .A(n793), .B(n15909), .Z(n15908) );
  XOR U15667 ( .A(n15910), .B(n15907), .Z(n15909) );
  XOR U15668 ( .A(n15911), .B(n15912), .Z(n15899) );
  AND U15669 ( .A(n15913), .B(n15914), .Z(n15912) );
  XOR U15670 ( .A(n15911), .B(n15736), .Z(n15914) );
  XOR U15671 ( .A(n15915), .B(n15916), .Z(n15736) );
  AND U15672 ( .A(n795), .B(n15917), .Z(n15916) );
  XOR U15673 ( .A(n15918), .B(n15915), .Z(n15917) );
  XNOR U15674 ( .A(n15733), .B(n15911), .Z(n15913) );
  XOR U15675 ( .A(n15919), .B(n15920), .Z(n15733) );
  AND U15676 ( .A(n793), .B(n15921), .Z(n15920) );
  XOR U15677 ( .A(n15922), .B(n15919), .Z(n15921) );
  XOR U15678 ( .A(n15923), .B(n15924), .Z(n15911) );
  AND U15679 ( .A(n15925), .B(n15926), .Z(n15924) );
  XOR U15680 ( .A(n15923), .B(n15748), .Z(n15926) );
  XOR U15681 ( .A(n15927), .B(n15928), .Z(n15748) );
  AND U15682 ( .A(n795), .B(n15929), .Z(n15928) );
  XOR U15683 ( .A(n15930), .B(n15927), .Z(n15929) );
  XNOR U15684 ( .A(n15745), .B(n15923), .Z(n15925) );
  XOR U15685 ( .A(n15931), .B(n15932), .Z(n15745) );
  AND U15686 ( .A(n793), .B(n15933), .Z(n15932) );
  XOR U15687 ( .A(n15934), .B(n15931), .Z(n15933) );
  XOR U15688 ( .A(n15935), .B(n15936), .Z(n15923) );
  AND U15689 ( .A(n15937), .B(n15938), .Z(n15936) );
  XOR U15690 ( .A(n15935), .B(n15760), .Z(n15938) );
  XOR U15691 ( .A(n15939), .B(n15940), .Z(n15760) );
  AND U15692 ( .A(n795), .B(n15941), .Z(n15940) );
  XOR U15693 ( .A(n15942), .B(n15939), .Z(n15941) );
  XNOR U15694 ( .A(n15757), .B(n15935), .Z(n15937) );
  XOR U15695 ( .A(n15943), .B(n15944), .Z(n15757) );
  AND U15696 ( .A(n793), .B(n15945), .Z(n15944) );
  XOR U15697 ( .A(n15946), .B(n15943), .Z(n15945) );
  XOR U15698 ( .A(n15947), .B(n15948), .Z(n15935) );
  AND U15699 ( .A(n15949), .B(n15950), .Z(n15948) );
  XOR U15700 ( .A(n15947), .B(n15772), .Z(n15950) );
  XOR U15701 ( .A(n15951), .B(n15952), .Z(n15772) );
  AND U15702 ( .A(n795), .B(n15953), .Z(n15952) );
  XOR U15703 ( .A(n15954), .B(n15951), .Z(n15953) );
  XNOR U15704 ( .A(n15769), .B(n15947), .Z(n15949) );
  XOR U15705 ( .A(n15955), .B(n15956), .Z(n15769) );
  AND U15706 ( .A(n793), .B(n15957), .Z(n15956) );
  XOR U15707 ( .A(n15958), .B(n15955), .Z(n15957) );
  XOR U15708 ( .A(n15959), .B(n15960), .Z(n15947) );
  AND U15709 ( .A(n15961), .B(n15962), .Z(n15960) );
  XOR U15710 ( .A(n15959), .B(n15784), .Z(n15962) );
  XOR U15711 ( .A(n15963), .B(n15964), .Z(n15784) );
  AND U15712 ( .A(n795), .B(n15965), .Z(n15964) );
  XOR U15713 ( .A(n15966), .B(n15963), .Z(n15965) );
  XNOR U15714 ( .A(n15781), .B(n15959), .Z(n15961) );
  XOR U15715 ( .A(n15967), .B(n15968), .Z(n15781) );
  AND U15716 ( .A(n793), .B(n15969), .Z(n15968) );
  XOR U15717 ( .A(n15970), .B(n15967), .Z(n15969) );
  XOR U15718 ( .A(n15971), .B(n15972), .Z(n15959) );
  AND U15719 ( .A(n15973), .B(n15974), .Z(n15972) );
  XNOR U15720 ( .A(n15975), .B(n15797), .Z(n15974) );
  XOR U15721 ( .A(n15976), .B(n15977), .Z(n15797) );
  AND U15722 ( .A(n795), .B(n15978), .Z(n15977) );
  XOR U15723 ( .A(n15976), .B(n15979), .Z(n15978) );
  XNOR U15724 ( .A(n15794), .B(n15971), .Z(n15973) );
  XOR U15725 ( .A(n15980), .B(n15981), .Z(n15794) );
  AND U15726 ( .A(n793), .B(n15982), .Z(n15981) );
  XOR U15727 ( .A(n15980), .B(n15983), .Z(n15982) );
  IV U15728 ( .A(n15975), .Z(n15971) );
  AND U15729 ( .A(n15802), .B(n15805), .Z(n15975) );
  XNOR U15730 ( .A(n15984), .B(n15985), .Z(n15805) );
  AND U15731 ( .A(n795), .B(n15986), .Z(n15985) );
  XNOR U15732 ( .A(n15987), .B(n15984), .Z(n15986) );
  XOR U15733 ( .A(n15988), .B(n15989), .Z(n795) );
  AND U15734 ( .A(n15990), .B(n15991), .Z(n15989) );
  XNOR U15735 ( .A(n15811), .B(n15988), .Z(n15991) );
  AND U15736 ( .A(n15992), .B(n15993), .Z(n15811) );
  XOR U15737 ( .A(n15988), .B(n15812), .Z(n15990) );
  AND U15738 ( .A(n15994), .B(n15995), .Z(n15812) );
  XOR U15739 ( .A(n15996), .B(n15997), .Z(n15988) );
  AND U15740 ( .A(n15998), .B(n15999), .Z(n15997) );
  XOR U15741 ( .A(n15996), .B(n15822), .Z(n15999) );
  XOR U15742 ( .A(n16000), .B(n16001), .Z(n15822) );
  AND U15743 ( .A(n483), .B(n16002), .Z(n16001) );
  XOR U15744 ( .A(n16003), .B(n16000), .Z(n16002) );
  XNOR U15745 ( .A(n15819), .B(n15996), .Z(n15998) );
  XOR U15746 ( .A(n16004), .B(n16005), .Z(n15819) );
  AND U15747 ( .A(n481), .B(n16006), .Z(n16005) );
  XOR U15748 ( .A(n16007), .B(n16004), .Z(n16006) );
  XOR U15749 ( .A(n16008), .B(n16009), .Z(n15996) );
  AND U15750 ( .A(n16010), .B(n16011), .Z(n16009) );
  XOR U15751 ( .A(n16008), .B(n15834), .Z(n16011) );
  XOR U15752 ( .A(n16012), .B(n16013), .Z(n15834) );
  AND U15753 ( .A(n483), .B(n16014), .Z(n16013) );
  XOR U15754 ( .A(n16015), .B(n16012), .Z(n16014) );
  XNOR U15755 ( .A(n15831), .B(n16008), .Z(n16010) );
  XOR U15756 ( .A(n16016), .B(n16017), .Z(n15831) );
  AND U15757 ( .A(n481), .B(n16018), .Z(n16017) );
  XOR U15758 ( .A(n16019), .B(n16016), .Z(n16018) );
  XOR U15759 ( .A(n16020), .B(n16021), .Z(n16008) );
  AND U15760 ( .A(n16022), .B(n16023), .Z(n16021) );
  XOR U15761 ( .A(n16020), .B(n15846), .Z(n16023) );
  XOR U15762 ( .A(n16024), .B(n16025), .Z(n15846) );
  AND U15763 ( .A(n483), .B(n16026), .Z(n16025) );
  XOR U15764 ( .A(n16027), .B(n16024), .Z(n16026) );
  XNOR U15765 ( .A(n15843), .B(n16020), .Z(n16022) );
  XOR U15766 ( .A(n16028), .B(n16029), .Z(n15843) );
  AND U15767 ( .A(n481), .B(n16030), .Z(n16029) );
  XOR U15768 ( .A(n16031), .B(n16028), .Z(n16030) );
  XOR U15769 ( .A(n16032), .B(n16033), .Z(n16020) );
  AND U15770 ( .A(n16034), .B(n16035), .Z(n16033) );
  XOR U15771 ( .A(n16032), .B(n15858), .Z(n16035) );
  XOR U15772 ( .A(n16036), .B(n16037), .Z(n15858) );
  AND U15773 ( .A(n483), .B(n16038), .Z(n16037) );
  XOR U15774 ( .A(n16039), .B(n16036), .Z(n16038) );
  XNOR U15775 ( .A(n15855), .B(n16032), .Z(n16034) );
  XOR U15776 ( .A(n16040), .B(n16041), .Z(n15855) );
  AND U15777 ( .A(n481), .B(n16042), .Z(n16041) );
  XOR U15778 ( .A(n16043), .B(n16040), .Z(n16042) );
  XOR U15779 ( .A(n16044), .B(n16045), .Z(n16032) );
  AND U15780 ( .A(n16046), .B(n16047), .Z(n16045) );
  XOR U15781 ( .A(n16044), .B(n15870), .Z(n16047) );
  XOR U15782 ( .A(n16048), .B(n16049), .Z(n15870) );
  AND U15783 ( .A(n483), .B(n16050), .Z(n16049) );
  XOR U15784 ( .A(n16051), .B(n16048), .Z(n16050) );
  XNOR U15785 ( .A(n15867), .B(n16044), .Z(n16046) );
  XOR U15786 ( .A(n16052), .B(n16053), .Z(n15867) );
  AND U15787 ( .A(n481), .B(n16054), .Z(n16053) );
  XOR U15788 ( .A(n16055), .B(n16052), .Z(n16054) );
  XOR U15789 ( .A(n16056), .B(n16057), .Z(n16044) );
  AND U15790 ( .A(n16058), .B(n16059), .Z(n16057) );
  XOR U15791 ( .A(n16056), .B(n15882), .Z(n16059) );
  XOR U15792 ( .A(n16060), .B(n16061), .Z(n15882) );
  AND U15793 ( .A(n483), .B(n16062), .Z(n16061) );
  XOR U15794 ( .A(n16063), .B(n16060), .Z(n16062) );
  XNOR U15795 ( .A(n15879), .B(n16056), .Z(n16058) );
  XOR U15796 ( .A(n16064), .B(n16065), .Z(n15879) );
  AND U15797 ( .A(n481), .B(n16066), .Z(n16065) );
  XOR U15798 ( .A(n16067), .B(n16064), .Z(n16066) );
  XOR U15799 ( .A(n16068), .B(n16069), .Z(n16056) );
  AND U15800 ( .A(n16070), .B(n16071), .Z(n16069) );
  XOR U15801 ( .A(n16068), .B(n15894), .Z(n16071) );
  XOR U15802 ( .A(n16072), .B(n16073), .Z(n15894) );
  AND U15803 ( .A(n483), .B(n16074), .Z(n16073) );
  XOR U15804 ( .A(n16075), .B(n16072), .Z(n16074) );
  XNOR U15805 ( .A(n15891), .B(n16068), .Z(n16070) );
  XOR U15806 ( .A(n16076), .B(n16077), .Z(n15891) );
  AND U15807 ( .A(n481), .B(n16078), .Z(n16077) );
  XOR U15808 ( .A(n16079), .B(n16076), .Z(n16078) );
  XOR U15809 ( .A(n16080), .B(n16081), .Z(n16068) );
  AND U15810 ( .A(n16082), .B(n16083), .Z(n16081) );
  XOR U15811 ( .A(n16080), .B(n15906), .Z(n16083) );
  XOR U15812 ( .A(n16084), .B(n16085), .Z(n15906) );
  AND U15813 ( .A(n483), .B(n16086), .Z(n16085) );
  XOR U15814 ( .A(n16087), .B(n16084), .Z(n16086) );
  XNOR U15815 ( .A(n15903), .B(n16080), .Z(n16082) );
  XOR U15816 ( .A(n16088), .B(n16089), .Z(n15903) );
  AND U15817 ( .A(n481), .B(n16090), .Z(n16089) );
  XOR U15818 ( .A(n16091), .B(n16088), .Z(n16090) );
  XOR U15819 ( .A(n16092), .B(n16093), .Z(n16080) );
  AND U15820 ( .A(n16094), .B(n16095), .Z(n16093) );
  XOR U15821 ( .A(n16092), .B(n15918), .Z(n16095) );
  XOR U15822 ( .A(n16096), .B(n16097), .Z(n15918) );
  AND U15823 ( .A(n483), .B(n16098), .Z(n16097) );
  XOR U15824 ( .A(n16099), .B(n16096), .Z(n16098) );
  XNOR U15825 ( .A(n15915), .B(n16092), .Z(n16094) );
  XOR U15826 ( .A(n16100), .B(n16101), .Z(n15915) );
  AND U15827 ( .A(n481), .B(n16102), .Z(n16101) );
  XOR U15828 ( .A(n16103), .B(n16100), .Z(n16102) );
  XOR U15829 ( .A(n16104), .B(n16105), .Z(n16092) );
  AND U15830 ( .A(n16106), .B(n16107), .Z(n16105) );
  XOR U15831 ( .A(n16104), .B(n15930), .Z(n16107) );
  XOR U15832 ( .A(n16108), .B(n16109), .Z(n15930) );
  AND U15833 ( .A(n483), .B(n16110), .Z(n16109) );
  XOR U15834 ( .A(n16111), .B(n16108), .Z(n16110) );
  XNOR U15835 ( .A(n15927), .B(n16104), .Z(n16106) );
  XOR U15836 ( .A(n16112), .B(n16113), .Z(n15927) );
  AND U15837 ( .A(n481), .B(n16114), .Z(n16113) );
  XOR U15838 ( .A(n16115), .B(n16112), .Z(n16114) );
  XOR U15839 ( .A(n16116), .B(n16117), .Z(n16104) );
  AND U15840 ( .A(n16118), .B(n16119), .Z(n16117) );
  XOR U15841 ( .A(n16116), .B(n15942), .Z(n16119) );
  XOR U15842 ( .A(n16120), .B(n16121), .Z(n15942) );
  AND U15843 ( .A(n483), .B(n16122), .Z(n16121) );
  XOR U15844 ( .A(n16123), .B(n16120), .Z(n16122) );
  XNOR U15845 ( .A(n15939), .B(n16116), .Z(n16118) );
  XOR U15846 ( .A(n16124), .B(n16125), .Z(n15939) );
  AND U15847 ( .A(n481), .B(n16126), .Z(n16125) );
  XOR U15848 ( .A(n16127), .B(n16124), .Z(n16126) );
  XOR U15849 ( .A(n16128), .B(n16129), .Z(n16116) );
  AND U15850 ( .A(n16130), .B(n16131), .Z(n16129) );
  XOR U15851 ( .A(n16128), .B(n15954), .Z(n16131) );
  XOR U15852 ( .A(n16132), .B(n16133), .Z(n15954) );
  AND U15853 ( .A(n483), .B(n16134), .Z(n16133) );
  XOR U15854 ( .A(n16135), .B(n16132), .Z(n16134) );
  XNOR U15855 ( .A(n15951), .B(n16128), .Z(n16130) );
  XOR U15856 ( .A(n16136), .B(n16137), .Z(n15951) );
  AND U15857 ( .A(n481), .B(n16138), .Z(n16137) );
  XOR U15858 ( .A(n16139), .B(n16136), .Z(n16138) );
  XOR U15859 ( .A(n16140), .B(n16141), .Z(n16128) );
  AND U15860 ( .A(n16142), .B(n16143), .Z(n16141) );
  XOR U15861 ( .A(n16140), .B(n15966), .Z(n16143) );
  XOR U15862 ( .A(n16144), .B(n16145), .Z(n15966) );
  AND U15863 ( .A(n483), .B(n16146), .Z(n16145) );
  XOR U15864 ( .A(n16147), .B(n16144), .Z(n16146) );
  XNOR U15865 ( .A(n15963), .B(n16140), .Z(n16142) );
  XOR U15866 ( .A(n16148), .B(n16149), .Z(n15963) );
  AND U15867 ( .A(n481), .B(n16150), .Z(n16149) );
  XOR U15868 ( .A(n16151), .B(n16148), .Z(n16150) );
  XOR U15869 ( .A(n16152), .B(n16153), .Z(n16140) );
  AND U15870 ( .A(n16154), .B(n16155), .Z(n16153) );
  XNOR U15871 ( .A(n16156), .B(n15979), .Z(n16155) );
  XOR U15872 ( .A(n16157), .B(n16158), .Z(n15979) );
  AND U15873 ( .A(n483), .B(n16159), .Z(n16158) );
  XOR U15874 ( .A(n16157), .B(n16160), .Z(n16159) );
  XNOR U15875 ( .A(n15976), .B(n16152), .Z(n16154) );
  XOR U15876 ( .A(n16161), .B(n16162), .Z(n15976) );
  AND U15877 ( .A(n481), .B(n16163), .Z(n16162) );
  XOR U15878 ( .A(n16161), .B(n16164), .Z(n16163) );
  IV U15879 ( .A(n16156), .Z(n16152) );
  AND U15880 ( .A(n15984), .B(n15987), .Z(n16156) );
  XNOR U15881 ( .A(n16165), .B(n16166), .Z(n15987) );
  AND U15882 ( .A(n483), .B(n16167), .Z(n16166) );
  XNOR U15883 ( .A(n16168), .B(n16165), .Z(n16167) );
  XOR U15884 ( .A(n16169), .B(n16170), .Z(n483) );
  AND U15885 ( .A(n16171), .B(n16172), .Z(n16170) );
  XNOR U15886 ( .A(n15992), .B(n16169), .Z(n16172) );
  AND U15887 ( .A(p_input[2047]), .B(p_input[2031]), .Z(n15992) );
  XOR U15888 ( .A(n16169), .B(n15993), .Z(n16171) );
  AND U15889 ( .A(p_input[2015]), .B(p_input[1999]), .Z(n15993) );
  XOR U15890 ( .A(n16173), .B(n16174), .Z(n16169) );
  AND U15891 ( .A(n16175), .B(n16176), .Z(n16174) );
  XOR U15892 ( .A(n16173), .B(n16003), .Z(n16176) );
  XNOR U15893 ( .A(p_input[2030]), .B(n16177), .Z(n16003) );
  AND U15894 ( .A(n611), .B(n16178), .Z(n16177) );
  XOR U15895 ( .A(p_input[2046]), .B(p_input[2030]), .Z(n16178) );
  XNOR U15896 ( .A(n16000), .B(n16173), .Z(n16175) );
  XOR U15897 ( .A(n16179), .B(n16180), .Z(n16000) );
  AND U15898 ( .A(n609), .B(n16181), .Z(n16180) );
  XOR U15899 ( .A(p_input[2014]), .B(p_input[1998]), .Z(n16181) );
  XOR U15900 ( .A(n16182), .B(n16183), .Z(n16173) );
  AND U15901 ( .A(n16184), .B(n16185), .Z(n16183) );
  XOR U15902 ( .A(n16182), .B(n16015), .Z(n16185) );
  XNOR U15903 ( .A(p_input[2029]), .B(n16186), .Z(n16015) );
  AND U15904 ( .A(n611), .B(n16187), .Z(n16186) );
  XOR U15905 ( .A(p_input[2045]), .B(p_input[2029]), .Z(n16187) );
  XNOR U15906 ( .A(n16012), .B(n16182), .Z(n16184) );
  XOR U15907 ( .A(n16188), .B(n16189), .Z(n16012) );
  AND U15908 ( .A(n609), .B(n16190), .Z(n16189) );
  XOR U15909 ( .A(p_input[2013]), .B(p_input[1997]), .Z(n16190) );
  XOR U15910 ( .A(n16191), .B(n16192), .Z(n16182) );
  AND U15911 ( .A(n16193), .B(n16194), .Z(n16192) );
  XOR U15912 ( .A(n16191), .B(n16027), .Z(n16194) );
  XNOR U15913 ( .A(p_input[2028]), .B(n16195), .Z(n16027) );
  AND U15914 ( .A(n611), .B(n16196), .Z(n16195) );
  XOR U15915 ( .A(p_input[2044]), .B(p_input[2028]), .Z(n16196) );
  XNOR U15916 ( .A(n16024), .B(n16191), .Z(n16193) );
  XOR U15917 ( .A(n16197), .B(n16198), .Z(n16024) );
  AND U15918 ( .A(n609), .B(n16199), .Z(n16198) );
  XOR U15919 ( .A(p_input[2012]), .B(p_input[1996]), .Z(n16199) );
  XOR U15920 ( .A(n16200), .B(n16201), .Z(n16191) );
  AND U15921 ( .A(n16202), .B(n16203), .Z(n16201) );
  XOR U15922 ( .A(n16200), .B(n16039), .Z(n16203) );
  XNOR U15923 ( .A(p_input[2027]), .B(n16204), .Z(n16039) );
  AND U15924 ( .A(n611), .B(n16205), .Z(n16204) );
  XOR U15925 ( .A(p_input[2043]), .B(p_input[2027]), .Z(n16205) );
  XNOR U15926 ( .A(n16036), .B(n16200), .Z(n16202) );
  XOR U15927 ( .A(n16206), .B(n16207), .Z(n16036) );
  AND U15928 ( .A(n609), .B(n16208), .Z(n16207) );
  XOR U15929 ( .A(p_input[2011]), .B(p_input[1995]), .Z(n16208) );
  XOR U15930 ( .A(n16209), .B(n16210), .Z(n16200) );
  AND U15931 ( .A(n16211), .B(n16212), .Z(n16210) );
  XOR U15932 ( .A(n16209), .B(n16051), .Z(n16212) );
  XNOR U15933 ( .A(p_input[2026]), .B(n16213), .Z(n16051) );
  AND U15934 ( .A(n611), .B(n16214), .Z(n16213) );
  XOR U15935 ( .A(p_input[2042]), .B(p_input[2026]), .Z(n16214) );
  XNOR U15936 ( .A(n16048), .B(n16209), .Z(n16211) );
  XOR U15937 ( .A(n16215), .B(n16216), .Z(n16048) );
  AND U15938 ( .A(n609), .B(n16217), .Z(n16216) );
  XOR U15939 ( .A(p_input[2010]), .B(p_input[1994]), .Z(n16217) );
  XOR U15940 ( .A(n16218), .B(n16219), .Z(n16209) );
  AND U15941 ( .A(n16220), .B(n16221), .Z(n16219) );
  XOR U15942 ( .A(n16218), .B(n16063), .Z(n16221) );
  XNOR U15943 ( .A(p_input[2025]), .B(n16222), .Z(n16063) );
  AND U15944 ( .A(n611), .B(n16223), .Z(n16222) );
  XOR U15945 ( .A(p_input[2041]), .B(p_input[2025]), .Z(n16223) );
  XNOR U15946 ( .A(n16060), .B(n16218), .Z(n16220) );
  XOR U15947 ( .A(n16224), .B(n16225), .Z(n16060) );
  AND U15948 ( .A(n609), .B(n16226), .Z(n16225) );
  XOR U15949 ( .A(p_input[2009]), .B(p_input[1993]), .Z(n16226) );
  XOR U15950 ( .A(n16227), .B(n16228), .Z(n16218) );
  AND U15951 ( .A(n16229), .B(n16230), .Z(n16228) );
  XOR U15952 ( .A(n16227), .B(n16075), .Z(n16230) );
  XNOR U15953 ( .A(p_input[2024]), .B(n16231), .Z(n16075) );
  AND U15954 ( .A(n611), .B(n16232), .Z(n16231) );
  XOR U15955 ( .A(p_input[2040]), .B(p_input[2024]), .Z(n16232) );
  XNOR U15956 ( .A(n16072), .B(n16227), .Z(n16229) );
  XOR U15957 ( .A(n16233), .B(n16234), .Z(n16072) );
  AND U15958 ( .A(n609), .B(n16235), .Z(n16234) );
  XOR U15959 ( .A(p_input[2008]), .B(p_input[1992]), .Z(n16235) );
  XOR U15960 ( .A(n16236), .B(n16237), .Z(n16227) );
  AND U15961 ( .A(n16238), .B(n16239), .Z(n16237) );
  XOR U15962 ( .A(n16236), .B(n16087), .Z(n16239) );
  XNOR U15963 ( .A(p_input[2023]), .B(n16240), .Z(n16087) );
  AND U15964 ( .A(n611), .B(n16241), .Z(n16240) );
  XOR U15965 ( .A(p_input[2039]), .B(p_input[2023]), .Z(n16241) );
  XNOR U15966 ( .A(n16084), .B(n16236), .Z(n16238) );
  XOR U15967 ( .A(n16242), .B(n16243), .Z(n16084) );
  AND U15968 ( .A(n609), .B(n16244), .Z(n16243) );
  XOR U15969 ( .A(p_input[2007]), .B(p_input[1991]), .Z(n16244) );
  XOR U15970 ( .A(n16245), .B(n16246), .Z(n16236) );
  AND U15971 ( .A(n16247), .B(n16248), .Z(n16246) );
  XOR U15972 ( .A(n16245), .B(n16099), .Z(n16248) );
  XNOR U15973 ( .A(p_input[2022]), .B(n16249), .Z(n16099) );
  AND U15974 ( .A(n611), .B(n16250), .Z(n16249) );
  XOR U15975 ( .A(p_input[2038]), .B(p_input[2022]), .Z(n16250) );
  XNOR U15976 ( .A(n16096), .B(n16245), .Z(n16247) );
  XOR U15977 ( .A(n16251), .B(n16252), .Z(n16096) );
  AND U15978 ( .A(n609), .B(n16253), .Z(n16252) );
  XOR U15979 ( .A(p_input[2006]), .B(p_input[1990]), .Z(n16253) );
  XOR U15980 ( .A(n16254), .B(n16255), .Z(n16245) );
  AND U15981 ( .A(n16256), .B(n16257), .Z(n16255) );
  XOR U15982 ( .A(n16254), .B(n16111), .Z(n16257) );
  XNOR U15983 ( .A(p_input[2021]), .B(n16258), .Z(n16111) );
  AND U15984 ( .A(n611), .B(n16259), .Z(n16258) );
  XOR U15985 ( .A(p_input[2037]), .B(p_input[2021]), .Z(n16259) );
  XNOR U15986 ( .A(n16108), .B(n16254), .Z(n16256) );
  XOR U15987 ( .A(n16260), .B(n16261), .Z(n16108) );
  AND U15988 ( .A(n609), .B(n16262), .Z(n16261) );
  XOR U15989 ( .A(p_input[2005]), .B(p_input[1989]), .Z(n16262) );
  XOR U15990 ( .A(n16263), .B(n16264), .Z(n16254) );
  AND U15991 ( .A(n16265), .B(n16266), .Z(n16264) );
  XOR U15992 ( .A(n16263), .B(n16123), .Z(n16266) );
  XNOR U15993 ( .A(p_input[2020]), .B(n16267), .Z(n16123) );
  AND U15994 ( .A(n611), .B(n16268), .Z(n16267) );
  XOR U15995 ( .A(p_input[2036]), .B(p_input[2020]), .Z(n16268) );
  XNOR U15996 ( .A(n16120), .B(n16263), .Z(n16265) );
  XOR U15997 ( .A(n16269), .B(n16270), .Z(n16120) );
  AND U15998 ( .A(n609), .B(n16271), .Z(n16270) );
  XOR U15999 ( .A(p_input[2004]), .B(p_input[1988]), .Z(n16271) );
  XOR U16000 ( .A(n16272), .B(n16273), .Z(n16263) );
  AND U16001 ( .A(n16274), .B(n16275), .Z(n16273) );
  XOR U16002 ( .A(n16272), .B(n16135), .Z(n16275) );
  XNOR U16003 ( .A(p_input[2019]), .B(n16276), .Z(n16135) );
  AND U16004 ( .A(n611), .B(n16277), .Z(n16276) );
  XOR U16005 ( .A(p_input[2035]), .B(p_input[2019]), .Z(n16277) );
  XNOR U16006 ( .A(n16132), .B(n16272), .Z(n16274) );
  XOR U16007 ( .A(n16278), .B(n16279), .Z(n16132) );
  AND U16008 ( .A(n609), .B(n16280), .Z(n16279) );
  XOR U16009 ( .A(p_input[2003]), .B(p_input[1987]), .Z(n16280) );
  XOR U16010 ( .A(n16281), .B(n16282), .Z(n16272) );
  AND U16011 ( .A(n16283), .B(n16284), .Z(n16282) );
  XOR U16012 ( .A(n16281), .B(n16147), .Z(n16284) );
  XNOR U16013 ( .A(p_input[2018]), .B(n16285), .Z(n16147) );
  AND U16014 ( .A(n611), .B(n16286), .Z(n16285) );
  XOR U16015 ( .A(p_input[2034]), .B(p_input[2018]), .Z(n16286) );
  XNOR U16016 ( .A(n16144), .B(n16281), .Z(n16283) );
  XOR U16017 ( .A(n16287), .B(n16288), .Z(n16144) );
  AND U16018 ( .A(n609), .B(n16289), .Z(n16288) );
  XOR U16019 ( .A(p_input[2002]), .B(p_input[1986]), .Z(n16289) );
  XOR U16020 ( .A(n16290), .B(n16291), .Z(n16281) );
  AND U16021 ( .A(n16292), .B(n16293), .Z(n16291) );
  XNOR U16022 ( .A(n16294), .B(n16160), .Z(n16293) );
  XNOR U16023 ( .A(p_input[2017]), .B(n16295), .Z(n16160) );
  AND U16024 ( .A(n611), .B(n16296), .Z(n16295) );
  XNOR U16025 ( .A(p_input[2033]), .B(n16297), .Z(n16296) );
  IV U16026 ( .A(p_input[2017]), .Z(n16297) );
  XNOR U16027 ( .A(n16157), .B(n16290), .Z(n16292) );
  XNOR U16028 ( .A(p_input[1985]), .B(n16298), .Z(n16157) );
  AND U16029 ( .A(n609), .B(n16299), .Z(n16298) );
  XOR U16030 ( .A(p_input[2001]), .B(p_input[1985]), .Z(n16299) );
  IV U16031 ( .A(n16294), .Z(n16290) );
  AND U16032 ( .A(n16165), .B(n16168), .Z(n16294) );
  XOR U16033 ( .A(p_input[2016]), .B(n16300), .Z(n16168) );
  AND U16034 ( .A(n611), .B(n16301), .Z(n16300) );
  XOR U16035 ( .A(p_input[2032]), .B(p_input[2016]), .Z(n16301) );
  XOR U16036 ( .A(n16302), .B(n16303), .Z(n611) );
  AND U16037 ( .A(n16304), .B(n16305), .Z(n16303) );
  XNOR U16038 ( .A(p_input[2047]), .B(n16302), .Z(n16305) );
  XOR U16039 ( .A(n16302), .B(p_input[2031]), .Z(n16304) );
  XOR U16040 ( .A(n16306), .B(n16307), .Z(n16302) );
  AND U16041 ( .A(n16308), .B(n16309), .Z(n16307) );
  XNOR U16042 ( .A(p_input[2046]), .B(n16306), .Z(n16309) );
  XOR U16043 ( .A(n16306), .B(p_input[2030]), .Z(n16308) );
  XOR U16044 ( .A(n16310), .B(n16311), .Z(n16306) );
  AND U16045 ( .A(n16312), .B(n16313), .Z(n16311) );
  XNOR U16046 ( .A(p_input[2045]), .B(n16310), .Z(n16313) );
  XOR U16047 ( .A(n16310), .B(p_input[2029]), .Z(n16312) );
  XOR U16048 ( .A(n16314), .B(n16315), .Z(n16310) );
  AND U16049 ( .A(n16316), .B(n16317), .Z(n16315) );
  XNOR U16050 ( .A(p_input[2044]), .B(n16314), .Z(n16317) );
  XOR U16051 ( .A(n16314), .B(p_input[2028]), .Z(n16316) );
  XOR U16052 ( .A(n16318), .B(n16319), .Z(n16314) );
  AND U16053 ( .A(n16320), .B(n16321), .Z(n16319) );
  XNOR U16054 ( .A(p_input[2043]), .B(n16318), .Z(n16321) );
  XOR U16055 ( .A(n16318), .B(p_input[2027]), .Z(n16320) );
  XOR U16056 ( .A(n16322), .B(n16323), .Z(n16318) );
  AND U16057 ( .A(n16324), .B(n16325), .Z(n16323) );
  XNOR U16058 ( .A(p_input[2042]), .B(n16322), .Z(n16325) );
  XOR U16059 ( .A(n16322), .B(p_input[2026]), .Z(n16324) );
  XOR U16060 ( .A(n16326), .B(n16327), .Z(n16322) );
  AND U16061 ( .A(n16328), .B(n16329), .Z(n16327) );
  XNOR U16062 ( .A(p_input[2041]), .B(n16326), .Z(n16329) );
  XOR U16063 ( .A(n16326), .B(p_input[2025]), .Z(n16328) );
  XOR U16064 ( .A(n16330), .B(n16331), .Z(n16326) );
  AND U16065 ( .A(n16332), .B(n16333), .Z(n16331) );
  XNOR U16066 ( .A(p_input[2040]), .B(n16330), .Z(n16333) );
  XOR U16067 ( .A(n16330), .B(p_input[2024]), .Z(n16332) );
  XOR U16068 ( .A(n16334), .B(n16335), .Z(n16330) );
  AND U16069 ( .A(n16336), .B(n16337), .Z(n16335) );
  XNOR U16070 ( .A(p_input[2039]), .B(n16334), .Z(n16337) );
  XOR U16071 ( .A(n16334), .B(p_input[2023]), .Z(n16336) );
  XOR U16072 ( .A(n16338), .B(n16339), .Z(n16334) );
  AND U16073 ( .A(n16340), .B(n16341), .Z(n16339) );
  XNOR U16074 ( .A(p_input[2038]), .B(n16338), .Z(n16341) );
  XOR U16075 ( .A(n16338), .B(p_input[2022]), .Z(n16340) );
  XOR U16076 ( .A(n16342), .B(n16343), .Z(n16338) );
  AND U16077 ( .A(n16344), .B(n16345), .Z(n16343) );
  XNOR U16078 ( .A(p_input[2037]), .B(n16342), .Z(n16345) );
  XOR U16079 ( .A(n16342), .B(p_input[2021]), .Z(n16344) );
  XOR U16080 ( .A(n16346), .B(n16347), .Z(n16342) );
  AND U16081 ( .A(n16348), .B(n16349), .Z(n16347) );
  XNOR U16082 ( .A(p_input[2036]), .B(n16346), .Z(n16349) );
  XOR U16083 ( .A(n16346), .B(p_input[2020]), .Z(n16348) );
  XOR U16084 ( .A(n16350), .B(n16351), .Z(n16346) );
  AND U16085 ( .A(n16352), .B(n16353), .Z(n16351) );
  XNOR U16086 ( .A(p_input[2035]), .B(n16350), .Z(n16353) );
  XOR U16087 ( .A(n16350), .B(p_input[2019]), .Z(n16352) );
  XOR U16088 ( .A(n16354), .B(n16355), .Z(n16350) );
  AND U16089 ( .A(n16356), .B(n16357), .Z(n16355) );
  XNOR U16090 ( .A(p_input[2034]), .B(n16354), .Z(n16357) );
  XOR U16091 ( .A(n16354), .B(p_input[2018]), .Z(n16356) );
  XNOR U16092 ( .A(n16358), .B(n16359), .Z(n16354) );
  AND U16093 ( .A(n16360), .B(n16361), .Z(n16359) );
  XOR U16094 ( .A(p_input[2033]), .B(n16358), .Z(n16361) );
  XNOR U16095 ( .A(p_input[2017]), .B(n16358), .Z(n16360) );
  AND U16096 ( .A(p_input[2032]), .B(n16362), .Z(n16358) );
  IV U16097 ( .A(p_input[2016]), .Z(n16362) );
  XNOR U16098 ( .A(p_input[1984]), .B(n16363), .Z(n16165) );
  AND U16099 ( .A(n609), .B(n16364), .Z(n16363) );
  XOR U16100 ( .A(p_input[2000]), .B(p_input[1984]), .Z(n16364) );
  XOR U16101 ( .A(n16365), .B(n16366), .Z(n609) );
  AND U16102 ( .A(n16367), .B(n16368), .Z(n16366) );
  XNOR U16103 ( .A(p_input[2015]), .B(n16365), .Z(n16368) );
  XOR U16104 ( .A(n16365), .B(p_input[1999]), .Z(n16367) );
  XOR U16105 ( .A(n16369), .B(n16370), .Z(n16365) );
  AND U16106 ( .A(n16371), .B(n16372), .Z(n16370) );
  XNOR U16107 ( .A(p_input[2014]), .B(n16369), .Z(n16372) );
  XNOR U16108 ( .A(n16369), .B(n16179), .Z(n16371) );
  IV U16109 ( .A(p_input[1998]), .Z(n16179) );
  XOR U16110 ( .A(n16373), .B(n16374), .Z(n16369) );
  AND U16111 ( .A(n16375), .B(n16376), .Z(n16374) );
  XNOR U16112 ( .A(p_input[2013]), .B(n16373), .Z(n16376) );
  XNOR U16113 ( .A(n16373), .B(n16188), .Z(n16375) );
  IV U16114 ( .A(p_input[1997]), .Z(n16188) );
  XOR U16115 ( .A(n16377), .B(n16378), .Z(n16373) );
  AND U16116 ( .A(n16379), .B(n16380), .Z(n16378) );
  XNOR U16117 ( .A(p_input[2012]), .B(n16377), .Z(n16380) );
  XNOR U16118 ( .A(n16377), .B(n16197), .Z(n16379) );
  IV U16119 ( .A(p_input[1996]), .Z(n16197) );
  XOR U16120 ( .A(n16381), .B(n16382), .Z(n16377) );
  AND U16121 ( .A(n16383), .B(n16384), .Z(n16382) );
  XNOR U16122 ( .A(p_input[2011]), .B(n16381), .Z(n16384) );
  XNOR U16123 ( .A(n16381), .B(n16206), .Z(n16383) );
  IV U16124 ( .A(p_input[1995]), .Z(n16206) );
  XOR U16125 ( .A(n16385), .B(n16386), .Z(n16381) );
  AND U16126 ( .A(n16387), .B(n16388), .Z(n16386) );
  XNOR U16127 ( .A(p_input[2010]), .B(n16385), .Z(n16388) );
  XNOR U16128 ( .A(n16385), .B(n16215), .Z(n16387) );
  IV U16129 ( .A(p_input[1994]), .Z(n16215) );
  XOR U16130 ( .A(n16389), .B(n16390), .Z(n16385) );
  AND U16131 ( .A(n16391), .B(n16392), .Z(n16390) );
  XNOR U16132 ( .A(p_input[2009]), .B(n16389), .Z(n16392) );
  XNOR U16133 ( .A(n16389), .B(n16224), .Z(n16391) );
  IV U16134 ( .A(p_input[1993]), .Z(n16224) );
  XOR U16135 ( .A(n16393), .B(n16394), .Z(n16389) );
  AND U16136 ( .A(n16395), .B(n16396), .Z(n16394) );
  XNOR U16137 ( .A(p_input[2008]), .B(n16393), .Z(n16396) );
  XNOR U16138 ( .A(n16393), .B(n16233), .Z(n16395) );
  IV U16139 ( .A(p_input[1992]), .Z(n16233) );
  XOR U16140 ( .A(n16397), .B(n16398), .Z(n16393) );
  AND U16141 ( .A(n16399), .B(n16400), .Z(n16398) );
  XNOR U16142 ( .A(p_input[2007]), .B(n16397), .Z(n16400) );
  XNOR U16143 ( .A(n16397), .B(n16242), .Z(n16399) );
  IV U16144 ( .A(p_input[1991]), .Z(n16242) );
  XOR U16145 ( .A(n16401), .B(n16402), .Z(n16397) );
  AND U16146 ( .A(n16403), .B(n16404), .Z(n16402) );
  XNOR U16147 ( .A(p_input[2006]), .B(n16401), .Z(n16404) );
  XNOR U16148 ( .A(n16401), .B(n16251), .Z(n16403) );
  IV U16149 ( .A(p_input[1990]), .Z(n16251) );
  XOR U16150 ( .A(n16405), .B(n16406), .Z(n16401) );
  AND U16151 ( .A(n16407), .B(n16408), .Z(n16406) );
  XNOR U16152 ( .A(p_input[2005]), .B(n16405), .Z(n16408) );
  XNOR U16153 ( .A(n16405), .B(n16260), .Z(n16407) );
  IV U16154 ( .A(p_input[1989]), .Z(n16260) );
  XOR U16155 ( .A(n16409), .B(n16410), .Z(n16405) );
  AND U16156 ( .A(n16411), .B(n16412), .Z(n16410) );
  XNOR U16157 ( .A(p_input[2004]), .B(n16409), .Z(n16412) );
  XNOR U16158 ( .A(n16409), .B(n16269), .Z(n16411) );
  IV U16159 ( .A(p_input[1988]), .Z(n16269) );
  XOR U16160 ( .A(n16413), .B(n16414), .Z(n16409) );
  AND U16161 ( .A(n16415), .B(n16416), .Z(n16414) );
  XNOR U16162 ( .A(p_input[2003]), .B(n16413), .Z(n16416) );
  XNOR U16163 ( .A(n16413), .B(n16278), .Z(n16415) );
  IV U16164 ( .A(p_input[1987]), .Z(n16278) );
  XOR U16165 ( .A(n16417), .B(n16418), .Z(n16413) );
  AND U16166 ( .A(n16419), .B(n16420), .Z(n16418) );
  XNOR U16167 ( .A(p_input[2002]), .B(n16417), .Z(n16420) );
  XNOR U16168 ( .A(n16417), .B(n16287), .Z(n16419) );
  IV U16169 ( .A(p_input[1986]), .Z(n16287) );
  XNOR U16170 ( .A(n16421), .B(n16422), .Z(n16417) );
  AND U16171 ( .A(n16423), .B(n16424), .Z(n16422) );
  XOR U16172 ( .A(p_input[2001]), .B(n16421), .Z(n16424) );
  XNOR U16173 ( .A(p_input[1985]), .B(n16421), .Z(n16423) );
  AND U16174 ( .A(p_input[2000]), .B(n16425), .Z(n16421) );
  IV U16175 ( .A(p_input[1984]), .Z(n16425) );
  XOR U16176 ( .A(n16426), .B(n16427), .Z(n15984) );
  AND U16177 ( .A(n481), .B(n16428), .Z(n16427) );
  XNOR U16178 ( .A(n16429), .B(n16426), .Z(n16428) );
  XOR U16179 ( .A(n16430), .B(n16431), .Z(n481) );
  AND U16180 ( .A(n16432), .B(n16433), .Z(n16431) );
  XNOR U16181 ( .A(n15994), .B(n16430), .Z(n16433) );
  AND U16182 ( .A(p_input[1983]), .B(p_input[1967]), .Z(n15994) );
  XOR U16183 ( .A(n16430), .B(n15995), .Z(n16432) );
  AND U16184 ( .A(p_input[1951]), .B(p_input[1935]), .Z(n15995) );
  XOR U16185 ( .A(n16434), .B(n16435), .Z(n16430) );
  AND U16186 ( .A(n16436), .B(n16437), .Z(n16435) );
  XOR U16187 ( .A(n16434), .B(n16007), .Z(n16437) );
  XNOR U16188 ( .A(p_input[1966]), .B(n16438), .Z(n16007) );
  AND U16189 ( .A(n615), .B(n16439), .Z(n16438) );
  XOR U16190 ( .A(p_input[1982]), .B(p_input[1966]), .Z(n16439) );
  XNOR U16191 ( .A(n16004), .B(n16434), .Z(n16436) );
  XOR U16192 ( .A(n16440), .B(n16441), .Z(n16004) );
  AND U16193 ( .A(n612), .B(n16442), .Z(n16441) );
  XOR U16194 ( .A(p_input[1950]), .B(p_input[1934]), .Z(n16442) );
  XOR U16195 ( .A(n16443), .B(n16444), .Z(n16434) );
  AND U16196 ( .A(n16445), .B(n16446), .Z(n16444) );
  XOR U16197 ( .A(n16443), .B(n16019), .Z(n16446) );
  XNOR U16198 ( .A(p_input[1965]), .B(n16447), .Z(n16019) );
  AND U16199 ( .A(n615), .B(n16448), .Z(n16447) );
  XOR U16200 ( .A(p_input[1981]), .B(p_input[1965]), .Z(n16448) );
  XNOR U16201 ( .A(n16016), .B(n16443), .Z(n16445) );
  XOR U16202 ( .A(n16449), .B(n16450), .Z(n16016) );
  AND U16203 ( .A(n612), .B(n16451), .Z(n16450) );
  XOR U16204 ( .A(p_input[1949]), .B(p_input[1933]), .Z(n16451) );
  XOR U16205 ( .A(n16452), .B(n16453), .Z(n16443) );
  AND U16206 ( .A(n16454), .B(n16455), .Z(n16453) );
  XOR U16207 ( .A(n16452), .B(n16031), .Z(n16455) );
  XNOR U16208 ( .A(p_input[1964]), .B(n16456), .Z(n16031) );
  AND U16209 ( .A(n615), .B(n16457), .Z(n16456) );
  XOR U16210 ( .A(p_input[1980]), .B(p_input[1964]), .Z(n16457) );
  XNOR U16211 ( .A(n16028), .B(n16452), .Z(n16454) );
  XOR U16212 ( .A(n16458), .B(n16459), .Z(n16028) );
  AND U16213 ( .A(n612), .B(n16460), .Z(n16459) );
  XOR U16214 ( .A(p_input[1948]), .B(p_input[1932]), .Z(n16460) );
  XOR U16215 ( .A(n16461), .B(n16462), .Z(n16452) );
  AND U16216 ( .A(n16463), .B(n16464), .Z(n16462) );
  XOR U16217 ( .A(n16461), .B(n16043), .Z(n16464) );
  XNOR U16218 ( .A(p_input[1963]), .B(n16465), .Z(n16043) );
  AND U16219 ( .A(n615), .B(n16466), .Z(n16465) );
  XOR U16220 ( .A(p_input[1979]), .B(p_input[1963]), .Z(n16466) );
  XNOR U16221 ( .A(n16040), .B(n16461), .Z(n16463) );
  XOR U16222 ( .A(n16467), .B(n16468), .Z(n16040) );
  AND U16223 ( .A(n612), .B(n16469), .Z(n16468) );
  XOR U16224 ( .A(p_input[1947]), .B(p_input[1931]), .Z(n16469) );
  XOR U16225 ( .A(n16470), .B(n16471), .Z(n16461) );
  AND U16226 ( .A(n16472), .B(n16473), .Z(n16471) );
  XOR U16227 ( .A(n16470), .B(n16055), .Z(n16473) );
  XNOR U16228 ( .A(p_input[1962]), .B(n16474), .Z(n16055) );
  AND U16229 ( .A(n615), .B(n16475), .Z(n16474) );
  XOR U16230 ( .A(p_input[1978]), .B(p_input[1962]), .Z(n16475) );
  XNOR U16231 ( .A(n16052), .B(n16470), .Z(n16472) );
  XOR U16232 ( .A(n16476), .B(n16477), .Z(n16052) );
  AND U16233 ( .A(n612), .B(n16478), .Z(n16477) );
  XOR U16234 ( .A(p_input[1946]), .B(p_input[1930]), .Z(n16478) );
  XOR U16235 ( .A(n16479), .B(n16480), .Z(n16470) );
  AND U16236 ( .A(n16481), .B(n16482), .Z(n16480) );
  XOR U16237 ( .A(n16479), .B(n16067), .Z(n16482) );
  XNOR U16238 ( .A(p_input[1961]), .B(n16483), .Z(n16067) );
  AND U16239 ( .A(n615), .B(n16484), .Z(n16483) );
  XOR U16240 ( .A(p_input[1977]), .B(p_input[1961]), .Z(n16484) );
  XNOR U16241 ( .A(n16064), .B(n16479), .Z(n16481) );
  XOR U16242 ( .A(n16485), .B(n16486), .Z(n16064) );
  AND U16243 ( .A(n612), .B(n16487), .Z(n16486) );
  XOR U16244 ( .A(p_input[1945]), .B(p_input[1929]), .Z(n16487) );
  XOR U16245 ( .A(n16488), .B(n16489), .Z(n16479) );
  AND U16246 ( .A(n16490), .B(n16491), .Z(n16489) );
  XOR U16247 ( .A(n16488), .B(n16079), .Z(n16491) );
  XNOR U16248 ( .A(p_input[1960]), .B(n16492), .Z(n16079) );
  AND U16249 ( .A(n615), .B(n16493), .Z(n16492) );
  XOR U16250 ( .A(p_input[1976]), .B(p_input[1960]), .Z(n16493) );
  XNOR U16251 ( .A(n16076), .B(n16488), .Z(n16490) );
  XOR U16252 ( .A(n16494), .B(n16495), .Z(n16076) );
  AND U16253 ( .A(n612), .B(n16496), .Z(n16495) );
  XOR U16254 ( .A(p_input[1944]), .B(p_input[1928]), .Z(n16496) );
  XOR U16255 ( .A(n16497), .B(n16498), .Z(n16488) );
  AND U16256 ( .A(n16499), .B(n16500), .Z(n16498) );
  XOR U16257 ( .A(n16497), .B(n16091), .Z(n16500) );
  XNOR U16258 ( .A(p_input[1959]), .B(n16501), .Z(n16091) );
  AND U16259 ( .A(n615), .B(n16502), .Z(n16501) );
  XOR U16260 ( .A(p_input[1975]), .B(p_input[1959]), .Z(n16502) );
  XNOR U16261 ( .A(n16088), .B(n16497), .Z(n16499) );
  XOR U16262 ( .A(n16503), .B(n16504), .Z(n16088) );
  AND U16263 ( .A(n612), .B(n16505), .Z(n16504) );
  XOR U16264 ( .A(p_input[1943]), .B(p_input[1927]), .Z(n16505) );
  XOR U16265 ( .A(n16506), .B(n16507), .Z(n16497) );
  AND U16266 ( .A(n16508), .B(n16509), .Z(n16507) );
  XOR U16267 ( .A(n16506), .B(n16103), .Z(n16509) );
  XNOR U16268 ( .A(p_input[1958]), .B(n16510), .Z(n16103) );
  AND U16269 ( .A(n615), .B(n16511), .Z(n16510) );
  XOR U16270 ( .A(p_input[1974]), .B(p_input[1958]), .Z(n16511) );
  XNOR U16271 ( .A(n16100), .B(n16506), .Z(n16508) );
  XOR U16272 ( .A(n16512), .B(n16513), .Z(n16100) );
  AND U16273 ( .A(n612), .B(n16514), .Z(n16513) );
  XOR U16274 ( .A(p_input[1942]), .B(p_input[1926]), .Z(n16514) );
  XOR U16275 ( .A(n16515), .B(n16516), .Z(n16506) );
  AND U16276 ( .A(n16517), .B(n16518), .Z(n16516) );
  XOR U16277 ( .A(n16515), .B(n16115), .Z(n16518) );
  XNOR U16278 ( .A(p_input[1957]), .B(n16519), .Z(n16115) );
  AND U16279 ( .A(n615), .B(n16520), .Z(n16519) );
  XOR U16280 ( .A(p_input[1973]), .B(p_input[1957]), .Z(n16520) );
  XNOR U16281 ( .A(n16112), .B(n16515), .Z(n16517) );
  XOR U16282 ( .A(n16521), .B(n16522), .Z(n16112) );
  AND U16283 ( .A(n612), .B(n16523), .Z(n16522) );
  XOR U16284 ( .A(p_input[1941]), .B(p_input[1925]), .Z(n16523) );
  XOR U16285 ( .A(n16524), .B(n16525), .Z(n16515) );
  AND U16286 ( .A(n16526), .B(n16527), .Z(n16525) );
  XOR U16287 ( .A(n16524), .B(n16127), .Z(n16527) );
  XNOR U16288 ( .A(p_input[1956]), .B(n16528), .Z(n16127) );
  AND U16289 ( .A(n615), .B(n16529), .Z(n16528) );
  XOR U16290 ( .A(p_input[1972]), .B(p_input[1956]), .Z(n16529) );
  XNOR U16291 ( .A(n16124), .B(n16524), .Z(n16526) );
  XOR U16292 ( .A(n16530), .B(n16531), .Z(n16124) );
  AND U16293 ( .A(n612), .B(n16532), .Z(n16531) );
  XOR U16294 ( .A(p_input[1940]), .B(p_input[1924]), .Z(n16532) );
  XOR U16295 ( .A(n16533), .B(n16534), .Z(n16524) );
  AND U16296 ( .A(n16535), .B(n16536), .Z(n16534) );
  XOR U16297 ( .A(n16533), .B(n16139), .Z(n16536) );
  XNOR U16298 ( .A(p_input[1955]), .B(n16537), .Z(n16139) );
  AND U16299 ( .A(n615), .B(n16538), .Z(n16537) );
  XOR U16300 ( .A(p_input[1971]), .B(p_input[1955]), .Z(n16538) );
  XNOR U16301 ( .A(n16136), .B(n16533), .Z(n16535) );
  XOR U16302 ( .A(n16539), .B(n16540), .Z(n16136) );
  AND U16303 ( .A(n612), .B(n16541), .Z(n16540) );
  XOR U16304 ( .A(p_input[1939]), .B(p_input[1923]), .Z(n16541) );
  XOR U16305 ( .A(n16542), .B(n16543), .Z(n16533) );
  AND U16306 ( .A(n16544), .B(n16545), .Z(n16543) );
  XOR U16307 ( .A(n16542), .B(n16151), .Z(n16545) );
  XNOR U16308 ( .A(p_input[1954]), .B(n16546), .Z(n16151) );
  AND U16309 ( .A(n615), .B(n16547), .Z(n16546) );
  XOR U16310 ( .A(p_input[1970]), .B(p_input[1954]), .Z(n16547) );
  XNOR U16311 ( .A(n16148), .B(n16542), .Z(n16544) );
  XOR U16312 ( .A(n16548), .B(n16549), .Z(n16148) );
  AND U16313 ( .A(n612), .B(n16550), .Z(n16549) );
  XOR U16314 ( .A(p_input[1938]), .B(p_input[1922]), .Z(n16550) );
  XOR U16315 ( .A(n16551), .B(n16552), .Z(n16542) );
  AND U16316 ( .A(n16553), .B(n16554), .Z(n16552) );
  XNOR U16317 ( .A(n16555), .B(n16164), .Z(n16554) );
  XNOR U16318 ( .A(p_input[1953]), .B(n16556), .Z(n16164) );
  AND U16319 ( .A(n615), .B(n16557), .Z(n16556) );
  XNOR U16320 ( .A(p_input[1969]), .B(n16558), .Z(n16557) );
  IV U16321 ( .A(p_input[1953]), .Z(n16558) );
  XNOR U16322 ( .A(n16161), .B(n16551), .Z(n16553) );
  XNOR U16323 ( .A(p_input[1921]), .B(n16559), .Z(n16161) );
  AND U16324 ( .A(n612), .B(n16560), .Z(n16559) );
  XOR U16325 ( .A(p_input[1937]), .B(p_input[1921]), .Z(n16560) );
  IV U16326 ( .A(n16555), .Z(n16551) );
  AND U16327 ( .A(n16426), .B(n16429), .Z(n16555) );
  XOR U16328 ( .A(p_input[1952]), .B(n16561), .Z(n16429) );
  AND U16329 ( .A(n615), .B(n16562), .Z(n16561) );
  XOR U16330 ( .A(p_input[1968]), .B(p_input[1952]), .Z(n16562) );
  XOR U16331 ( .A(n16563), .B(n16564), .Z(n615) );
  AND U16332 ( .A(n16565), .B(n16566), .Z(n16564) );
  XNOR U16333 ( .A(p_input[1983]), .B(n16563), .Z(n16566) );
  XOR U16334 ( .A(n16563), .B(p_input[1967]), .Z(n16565) );
  XOR U16335 ( .A(n16567), .B(n16568), .Z(n16563) );
  AND U16336 ( .A(n16569), .B(n16570), .Z(n16568) );
  XNOR U16337 ( .A(p_input[1982]), .B(n16567), .Z(n16570) );
  XOR U16338 ( .A(n16567), .B(p_input[1966]), .Z(n16569) );
  XOR U16339 ( .A(n16571), .B(n16572), .Z(n16567) );
  AND U16340 ( .A(n16573), .B(n16574), .Z(n16572) );
  XNOR U16341 ( .A(p_input[1981]), .B(n16571), .Z(n16574) );
  XOR U16342 ( .A(n16571), .B(p_input[1965]), .Z(n16573) );
  XOR U16343 ( .A(n16575), .B(n16576), .Z(n16571) );
  AND U16344 ( .A(n16577), .B(n16578), .Z(n16576) );
  XNOR U16345 ( .A(p_input[1980]), .B(n16575), .Z(n16578) );
  XOR U16346 ( .A(n16575), .B(p_input[1964]), .Z(n16577) );
  XOR U16347 ( .A(n16579), .B(n16580), .Z(n16575) );
  AND U16348 ( .A(n16581), .B(n16582), .Z(n16580) );
  XNOR U16349 ( .A(p_input[1979]), .B(n16579), .Z(n16582) );
  XOR U16350 ( .A(n16579), .B(p_input[1963]), .Z(n16581) );
  XOR U16351 ( .A(n16583), .B(n16584), .Z(n16579) );
  AND U16352 ( .A(n16585), .B(n16586), .Z(n16584) );
  XNOR U16353 ( .A(p_input[1978]), .B(n16583), .Z(n16586) );
  XOR U16354 ( .A(n16583), .B(p_input[1962]), .Z(n16585) );
  XOR U16355 ( .A(n16587), .B(n16588), .Z(n16583) );
  AND U16356 ( .A(n16589), .B(n16590), .Z(n16588) );
  XNOR U16357 ( .A(p_input[1977]), .B(n16587), .Z(n16590) );
  XOR U16358 ( .A(n16587), .B(p_input[1961]), .Z(n16589) );
  XOR U16359 ( .A(n16591), .B(n16592), .Z(n16587) );
  AND U16360 ( .A(n16593), .B(n16594), .Z(n16592) );
  XNOR U16361 ( .A(p_input[1976]), .B(n16591), .Z(n16594) );
  XOR U16362 ( .A(n16591), .B(p_input[1960]), .Z(n16593) );
  XOR U16363 ( .A(n16595), .B(n16596), .Z(n16591) );
  AND U16364 ( .A(n16597), .B(n16598), .Z(n16596) );
  XNOR U16365 ( .A(p_input[1975]), .B(n16595), .Z(n16598) );
  XOR U16366 ( .A(n16595), .B(p_input[1959]), .Z(n16597) );
  XOR U16367 ( .A(n16599), .B(n16600), .Z(n16595) );
  AND U16368 ( .A(n16601), .B(n16602), .Z(n16600) );
  XNOR U16369 ( .A(p_input[1974]), .B(n16599), .Z(n16602) );
  XOR U16370 ( .A(n16599), .B(p_input[1958]), .Z(n16601) );
  XOR U16371 ( .A(n16603), .B(n16604), .Z(n16599) );
  AND U16372 ( .A(n16605), .B(n16606), .Z(n16604) );
  XNOR U16373 ( .A(p_input[1973]), .B(n16603), .Z(n16606) );
  XOR U16374 ( .A(n16603), .B(p_input[1957]), .Z(n16605) );
  XOR U16375 ( .A(n16607), .B(n16608), .Z(n16603) );
  AND U16376 ( .A(n16609), .B(n16610), .Z(n16608) );
  XNOR U16377 ( .A(p_input[1972]), .B(n16607), .Z(n16610) );
  XOR U16378 ( .A(n16607), .B(p_input[1956]), .Z(n16609) );
  XOR U16379 ( .A(n16611), .B(n16612), .Z(n16607) );
  AND U16380 ( .A(n16613), .B(n16614), .Z(n16612) );
  XNOR U16381 ( .A(p_input[1971]), .B(n16611), .Z(n16614) );
  XOR U16382 ( .A(n16611), .B(p_input[1955]), .Z(n16613) );
  XOR U16383 ( .A(n16615), .B(n16616), .Z(n16611) );
  AND U16384 ( .A(n16617), .B(n16618), .Z(n16616) );
  XNOR U16385 ( .A(p_input[1970]), .B(n16615), .Z(n16618) );
  XOR U16386 ( .A(n16615), .B(p_input[1954]), .Z(n16617) );
  XNOR U16387 ( .A(n16619), .B(n16620), .Z(n16615) );
  AND U16388 ( .A(n16621), .B(n16622), .Z(n16620) );
  XOR U16389 ( .A(p_input[1969]), .B(n16619), .Z(n16622) );
  XNOR U16390 ( .A(p_input[1953]), .B(n16619), .Z(n16621) );
  AND U16391 ( .A(p_input[1968]), .B(n16623), .Z(n16619) );
  IV U16392 ( .A(p_input[1952]), .Z(n16623) );
  XNOR U16393 ( .A(p_input[1920]), .B(n16624), .Z(n16426) );
  AND U16394 ( .A(n612), .B(n16625), .Z(n16624) );
  XOR U16395 ( .A(p_input[1936]), .B(p_input[1920]), .Z(n16625) );
  XOR U16396 ( .A(n16626), .B(n16627), .Z(n612) );
  AND U16397 ( .A(n16628), .B(n16629), .Z(n16627) );
  XNOR U16398 ( .A(p_input[1951]), .B(n16626), .Z(n16629) );
  XOR U16399 ( .A(n16626), .B(p_input[1935]), .Z(n16628) );
  XOR U16400 ( .A(n16630), .B(n16631), .Z(n16626) );
  AND U16401 ( .A(n16632), .B(n16633), .Z(n16631) );
  XNOR U16402 ( .A(p_input[1950]), .B(n16630), .Z(n16633) );
  XNOR U16403 ( .A(n16630), .B(n16440), .Z(n16632) );
  IV U16404 ( .A(p_input[1934]), .Z(n16440) );
  XOR U16405 ( .A(n16634), .B(n16635), .Z(n16630) );
  AND U16406 ( .A(n16636), .B(n16637), .Z(n16635) );
  XNOR U16407 ( .A(p_input[1949]), .B(n16634), .Z(n16637) );
  XNOR U16408 ( .A(n16634), .B(n16449), .Z(n16636) );
  IV U16409 ( .A(p_input[1933]), .Z(n16449) );
  XOR U16410 ( .A(n16638), .B(n16639), .Z(n16634) );
  AND U16411 ( .A(n16640), .B(n16641), .Z(n16639) );
  XNOR U16412 ( .A(p_input[1948]), .B(n16638), .Z(n16641) );
  XNOR U16413 ( .A(n16638), .B(n16458), .Z(n16640) );
  IV U16414 ( .A(p_input[1932]), .Z(n16458) );
  XOR U16415 ( .A(n16642), .B(n16643), .Z(n16638) );
  AND U16416 ( .A(n16644), .B(n16645), .Z(n16643) );
  XNOR U16417 ( .A(p_input[1947]), .B(n16642), .Z(n16645) );
  XNOR U16418 ( .A(n16642), .B(n16467), .Z(n16644) );
  IV U16419 ( .A(p_input[1931]), .Z(n16467) );
  XOR U16420 ( .A(n16646), .B(n16647), .Z(n16642) );
  AND U16421 ( .A(n16648), .B(n16649), .Z(n16647) );
  XNOR U16422 ( .A(p_input[1946]), .B(n16646), .Z(n16649) );
  XNOR U16423 ( .A(n16646), .B(n16476), .Z(n16648) );
  IV U16424 ( .A(p_input[1930]), .Z(n16476) );
  XOR U16425 ( .A(n16650), .B(n16651), .Z(n16646) );
  AND U16426 ( .A(n16652), .B(n16653), .Z(n16651) );
  XNOR U16427 ( .A(p_input[1945]), .B(n16650), .Z(n16653) );
  XNOR U16428 ( .A(n16650), .B(n16485), .Z(n16652) );
  IV U16429 ( .A(p_input[1929]), .Z(n16485) );
  XOR U16430 ( .A(n16654), .B(n16655), .Z(n16650) );
  AND U16431 ( .A(n16656), .B(n16657), .Z(n16655) );
  XNOR U16432 ( .A(p_input[1944]), .B(n16654), .Z(n16657) );
  XNOR U16433 ( .A(n16654), .B(n16494), .Z(n16656) );
  IV U16434 ( .A(p_input[1928]), .Z(n16494) );
  XOR U16435 ( .A(n16658), .B(n16659), .Z(n16654) );
  AND U16436 ( .A(n16660), .B(n16661), .Z(n16659) );
  XNOR U16437 ( .A(p_input[1943]), .B(n16658), .Z(n16661) );
  XNOR U16438 ( .A(n16658), .B(n16503), .Z(n16660) );
  IV U16439 ( .A(p_input[1927]), .Z(n16503) );
  XOR U16440 ( .A(n16662), .B(n16663), .Z(n16658) );
  AND U16441 ( .A(n16664), .B(n16665), .Z(n16663) );
  XNOR U16442 ( .A(p_input[1942]), .B(n16662), .Z(n16665) );
  XNOR U16443 ( .A(n16662), .B(n16512), .Z(n16664) );
  IV U16444 ( .A(p_input[1926]), .Z(n16512) );
  XOR U16445 ( .A(n16666), .B(n16667), .Z(n16662) );
  AND U16446 ( .A(n16668), .B(n16669), .Z(n16667) );
  XNOR U16447 ( .A(p_input[1941]), .B(n16666), .Z(n16669) );
  XNOR U16448 ( .A(n16666), .B(n16521), .Z(n16668) );
  IV U16449 ( .A(p_input[1925]), .Z(n16521) );
  XOR U16450 ( .A(n16670), .B(n16671), .Z(n16666) );
  AND U16451 ( .A(n16672), .B(n16673), .Z(n16671) );
  XNOR U16452 ( .A(p_input[1940]), .B(n16670), .Z(n16673) );
  XNOR U16453 ( .A(n16670), .B(n16530), .Z(n16672) );
  IV U16454 ( .A(p_input[1924]), .Z(n16530) );
  XOR U16455 ( .A(n16674), .B(n16675), .Z(n16670) );
  AND U16456 ( .A(n16676), .B(n16677), .Z(n16675) );
  XNOR U16457 ( .A(p_input[1939]), .B(n16674), .Z(n16677) );
  XNOR U16458 ( .A(n16674), .B(n16539), .Z(n16676) );
  IV U16459 ( .A(p_input[1923]), .Z(n16539) );
  XOR U16460 ( .A(n16678), .B(n16679), .Z(n16674) );
  AND U16461 ( .A(n16680), .B(n16681), .Z(n16679) );
  XNOR U16462 ( .A(p_input[1938]), .B(n16678), .Z(n16681) );
  XNOR U16463 ( .A(n16678), .B(n16548), .Z(n16680) );
  IV U16464 ( .A(p_input[1922]), .Z(n16548) );
  XNOR U16465 ( .A(n16682), .B(n16683), .Z(n16678) );
  AND U16466 ( .A(n16684), .B(n16685), .Z(n16683) );
  XOR U16467 ( .A(p_input[1937]), .B(n16682), .Z(n16685) );
  XNOR U16468 ( .A(p_input[1921]), .B(n16682), .Z(n16684) );
  AND U16469 ( .A(p_input[1936]), .B(n16686), .Z(n16682) );
  IV U16470 ( .A(p_input[1920]), .Z(n16686) );
  XOR U16471 ( .A(n16687), .B(n16688), .Z(n15802) );
  AND U16472 ( .A(n793), .B(n16689), .Z(n16688) );
  XNOR U16473 ( .A(n16690), .B(n16687), .Z(n16689) );
  XOR U16474 ( .A(n16691), .B(n16692), .Z(n793) );
  AND U16475 ( .A(n16693), .B(n16694), .Z(n16692) );
  XNOR U16476 ( .A(n15814), .B(n16691), .Z(n16694) );
  AND U16477 ( .A(n16695), .B(n16696), .Z(n15814) );
  XOR U16478 ( .A(n16691), .B(n15813), .Z(n16693) );
  AND U16479 ( .A(n16697), .B(n16698), .Z(n15813) );
  XOR U16480 ( .A(n16699), .B(n16700), .Z(n16691) );
  AND U16481 ( .A(n16701), .B(n16702), .Z(n16700) );
  XOR U16482 ( .A(n16699), .B(n15826), .Z(n16702) );
  XOR U16483 ( .A(n16703), .B(n16704), .Z(n15826) );
  AND U16484 ( .A(n487), .B(n16705), .Z(n16704) );
  XOR U16485 ( .A(n16706), .B(n16703), .Z(n16705) );
  XNOR U16486 ( .A(n15823), .B(n16699), .Z(n16701) );
  XOR U16487 ( .A(n16707), .B(n16708), .Z(n15823) );
  AND U16488 ( .A(n484), .B(n16709), .Z(n16708) );
  XOR U16489 ( .A(n16710), .B(n16707), .Z(n16709) );
  XOR U16490 ( .A(n16711), .B(n16712), .Z(n16699) );
  AND U16491 ( .A(n16713), .B(n16714), .Z(n16712) );
  XOR U16492 ( .A(n16711), .B(n15838), .Z(n16714) );
  XOR U16493 ( .A(n16715), .B(n16716), .Z(n15838) );
  AND U16494 ( .A(n487), .B(n16717), .Z(n16716) );
  XOR U16495 ( .A(n16718), .B(n16715), .Z(n16717) );
  XNOR U16496 ( .A(n15835), .B(n16711), .Z(n16713) );
  XOR U16497 ( .A(n16719), .B(n16720), .Z(n15835) );
  AND U16498 ( .A(n484), .B(n16721), .Z(n16720) );
  XOR U16499 ( .A(n16722), .B(n16719), .Z(n16721) );
  XOR U16500 ( .A(n16723), .B(n16724), .Z(n16711) );
  AND U16501 ( .A(n16725), .B(n16726), .Z(n16724) );
  XOR U16502 ( .A(n16723), .B(n15850), .Z(n16726) );
  XOR U16503 ( .A(n16727), .B(n16728), .Z(n15850) );
  AND U16504 ( .A(n487), .B(n16729), .Z(n16728) );
  XOR U16505 ( .A(n16730), .B(n16727), .Z(n16729) );
  XNOR U16506 ( .A(n15847), .B(n16723), .Z(n16725) );
  XOR U16507 ( .A(n16731), .B(n16732), .Z(n15847) );
  AND U16508 ( .A(n484), .B(n16733), .Z(n16732) );
  XOR U16509 ( .A(n16734), .B(n16731), .Z(n16733) );
  XOR U16510 ( .A(n16735), .B(n16736), .Z(n16723) );
  AND U16511 ( .A(n16737), .B(n16738), .Z(n16736) );
  XOR U16512 ( .A(n16735), .B(n15862), .Z(n16738) );
  XOR U16513 ( .A(n16739), .B(n16740), .Z(n15862) );
  AND U16514 ( .A(n487), .B(n16741), .Z(n16740) );
  XOR U16515 ( .A(n16742), .B(n16739), .Z(n16741) );
  XNOR U16516 ( .A(n15859), .B(n16735), .Z(n16737) );
  XOR U16517 ( .A(n16743), .B(n16744), .Z(n15859) );
  AND U16518 ( .A(n484), .B(n16745), .Z(n16744) );
  XOR U16519 ( .A(n16746), .B(n16743), .Z(n16745) );
  XOR U16520 ( .A(n16747), .B(n16748), .Z(n16735) );
  AND U16521 ( .A(n16749), .B(n16750), .Z(n16748) );
  XOR U16522 ( .A(n16747), .B(n15874), .Z(n16750) );
  XOR U16523 ( .A(n16751), .B(n16752), .Z(n15874) );
  AND U16524 ( .A(n487), .B(n16753), .Z(n16752) );
  XOR U16525 ( .A(n16754), .B(n16751), .Z(n16753) );
  XNOR U16526 ( .A(n15871), .B(n16747), .Z(n16749) );
  XOR U16527 ( .A(n16755), .B(n16756), .Z(n15871) );
  AND U16528 ( .A(n484), .B(n16757), .Z(n16756) );
  XOR U16529 ( .A(n16758), .B(n16755), .Z(n16757) );
  XOR U16530 ( .A(n16759), .B(n16760), .Z(n16747) );
  AND U16531 ( .A(n16761), .B(n16762), .Z(n16760) );
  XOR U16532 ( .A(n16759), .B(n15886), .Z(n16762) );
  XOR U16533 ( .A(n16763), .B(n16764), .Z(n15886) );
  AND U16534 ( .A(n487), .B(n16765), .Z(n16764) );
  XOR U16535 ( .A(n16766), .B(n16763), .Z(n16765) );
  XNOR U16536 ( .A(n15883), .B(n16759), .Z(n16761) );
  XOR U16537 ( .A(n16767), .B(n16768), .Z(n15883) );
  AND U16538 ( .A(n484), .B(n16769), .Z(n16768) );
  XOR U16539 ( .A(n16770), .B(n16767), .Z(n16769) );
  XOR U16540 ( .A(n16771), .B(n16772), .Z(n16759) );
  AND U16541 ( .A(n16773), .B(n16774), .Z(n16772) );
  XOR U16542 ( .A(n16771), .B(n15898), .Z(n16774) );
  XOR U16543 ( .A(n16775), .B(n16776), .Z(n15898) );
  AND U16544 ( .A(n487), .B(n16777), .Z(n16776) );
  XOR U16545 ( .A(n16778), .B(n16775), .Z(n16777) );
  XNOR U16546 ( .A(n15895), .B(n16771), .Z(n16773) );
  XOR U16547 ( .A(n16779), .B(n16780), .Z(n15895) );
  AND U16548 ( .A(n484), .B(n16781), .Z(n16780) );
  XOR U16549 ( .A(n16782), .B(n16779), .Z(n16781) );
  XOR U16550 ( .A(n16783), .B(n16784), .Z(n16771) );
  AND U16551 ( .A(n16785), .B(n16786), .Z(n16784) );
  XOR U16552 ( .A(n16783), .B(n15910), .Z(n16786) );
  XOR U16553 ( .A(n16787), .B(n16788), .Z(n15910) );
  AND U16554 ( .A(n487), .B(n16789), .Z(n16788) );
  XOR U16555 ( .A(n16790), .B(n16787), .Z(n16789) );
  XNOR U16556 ( .A(n15907), .B(n16783), .Z(n16785) );
  XOR U16557 ( .A(n16791), .B(n16792), .Z(n15907) );
  AND U16558 ( .A(n484), .B(n16793), .Z(n16792) );
  XOR U16559 ( .A(n16794), .B(n16791), .Z(n16793) );
  XOR U16560 ( .A(n16795), .B(n16796), .Z(n16783) );
  AND U16561 ( .A(n16797), .B(n16798), .Z(n16796) );
  XOR U16562 ( .A(n16795), .B(n15922), .Z(n16798) );
  XOR U16563 ( .A(n16799), .B(n16800), .Z(n15922) );
  AND U16564 ( .A(n487), .B(n16801), .Z(n16800) );
  XOR U16565 ( .A(n16802), .B(n16799), .Z(n16801) );
  XNOR U16566 ( .A(n15919), .B(n16795), .Z(n16797) );
  XOR U16567 ( .A(n16803), .B(n16804), .Z(n15919) );
  AND U16568 ( .A(n484), .B(n16805), .Z(n16804) );
  XOR U16569 ( .A(n16806), .B(n16803), .Z(n16805) );
  XOR U16570 ( .A(n16807), .B(n16808), .Z(n16795) );
  AND U16571 ( .A(n16809), .B(n16810), .Z(n16808) );
  XOR U16572 ( .A(n16807), .B(n15934), .Z(n16810) );
  XOR U16573 ( .A(n16811), .B(n16812), .Z(n15934) );
  AND U16574 ( .A(n487), .B(n16813), .Z(n16812) );
  XOR U16575 ( .A(n16814), .B(n16811), .Z(n16813) );
  XNOR U16576 ( .A(n15931), .B(n16807), .Z(n16809) );
  XOR U16577 ( .A(n16815), .B(n16816), .Z(n15931) );
  AND U16578 ( .A(n484), .B(n16817), .Z(n16816) );
  XOR U16579 ( .A(n16818), .B(n16815), .Z(n16817) );
  XOR U16580 ( .A(n16819), .B(n16820), .Z(n16807) );
  AND U16581 ( .A(n16821), .B(n16822), .Z(n16820) );
  XOR U16582 ( .A(n16819), .B(n15946), .Z(n16822) );
  XOR U16583 ( .A(n16823), .B(n16824), .Z(n15946) );
  AND U16584 ( .A(n487), .B(n16825), .Z(n16824) );
  XOR U16585 ( .A(n16826), .B(n16823), .Z(n16825) );
  XNOR U16586 ( .A(n15943), .B(n16819), .Z(n16821) );
  XOR U16587 ( .A(n16827), .B(n16828), .Z(n15943) );
  AND U16588 ( .A(n484), .B(n16829), .Z(n16828) );
  XOR U16589 ( .A(n16830), .B(n16827), .Z(n16829) );
  XOR U16590 ( .A(n16831), .B(n16832), .Z(n16819) );
  AND U16591 ( .A(n16833), .B(n16834), .Z(n16832) );
  XOR U16592 ( .A(n16831), .B(n15958), .Z(n16834) );
  XOR U16593 ( .A(n16835), .B(n16836), .Z(n15958) );
  AND U16594 ( .A(n487), .B(n16837), .Z(n16836) );
  XOR U16595 ( .A(n16838), .B(n16835), .Z(n16837) );
  XNOR U16596 ( .A(n15955), .B(n16831), .Z(n16833) );
  XOR U16597 ( .A(n16839), .B(n16840), .Z(n15955) );
  AND U16598 ( .A(n484), .B(n16841), .Z(n16840) );
  XOR U16599 ( .A(n16842), .B(n16839), .Z(n16841) );
  XOR U16600 ( .A(n16843), .B(n16844), .Z(n16831) );
  AND U16601 ( .A(n16845), .B(n16846), .Z(n16844) );
  XOR U16602 ( .A(n16843), .B(n15970), .Z(n16846) );
  XOR U16603 ( .A(n16847), .B(n16848), .Z(n15970) );
  AND U16604 ( .A(n487), .B(n16849), .Z(n16848) );
  XOR U16605 ( .A(n16850), .B(n16847), .Z(n16849) );
  XNOR U16606 ( .A(n15967), .B(n16843), .Z(n16845) );
  XOR U16607 ( .A(n16851), .B(n16852), .Z(n15967) );
  AND U16608 ( .A(n484), .B(n16853), .Z(n16852) );
  XOR U16609 ( .A(n16854), .B(n16851), .Z(n16853) );
  XOR U16610 ( .A(n16855), .B(n16856), .Z(n16843) );
  AND U16611 ( .A(n16857), .B(n16858), .Z(n16856) );
  XNOR U16612 ( .A(n16859), .B(n15983), .Z(n16858) );
  XOR U16613 ( .A(n16860), .B(n16861), .Z(n15983) );
  AND U16614 ( .A(n487), .B(n16862), .Z(n16861) );
  XOR U16615 ( .A(n16860), .B(n16863), .Z(n16862) );
  XNOR U16616 ( .A(n15980), .B(n16855), .Z(n16857) );
  XOR U16617 ( .A(n16864), .B(n16865), .Z(n15980) );
  AND U16618 ( .A(n484), .B(n16866), .Z(n16865) );
  XOR U16619 ( .A(n16864), .B(n16867), .Z(n16866) );
  IV U16620 ( .A(n16859), .Z(n16855) );
  AND U16621 ( .A(n16687), .B(n16690), .Z(n16859) );
  XNOR U16622 ( .A(n16868), .B(n16869), .Z(n16690) );
  AND U16623 ( .A(n487), .B(n16870), .Z(n16869) );
  XNOR U16624 ( .A(n16871), .B(n16868), .Z(n16870) );
  XOR U16625 ( .A(n16872), .B(n16873), .Z(n487) );
  AND U16626 ( .A(n16874), .B(n16875), .Z(n16873) );
  XNOR U16627 ( .A(n16695), .B(n16872), .Z(n16875) );
  AND U16628 ( .A(p_input[1919]), .B(p_input[1903]), .Z(n16695) );
  XOR U16629 ( .A(n16872), .B(n16696), .Z(n16874) );
  AND U16630 ( .A(p_input[1887]), .B(p_input[1871]), .Z(n16696) );
  XOR U16631 ( .A(n16876), .B(n16877), .Z(n16872) );
  AND U16632 ( .A(n16878), .B(n16879), .Z(n16877) );
  XOR U16633 ( .A(n16876), .B(n16706), .Z(n16879) );
  XNOR U16634 ( .A(p_input[1902]), .B(n16880), .Z(n16706) );
  AND U16635 ( .A(n623), .B(n16881), .Z(n16880) );
  XOR U16636 ( .A(p_input[1918]), .B(p_input[1902]), .Z(n16881) );
  XNOR U16637 ( .A(n16703), .B(n16876), .Z(n16878) );
  XOR U16638 ( .A(n16882), .B(n16883), .Z(n16703) );
  AND U16639 ( .A(n621), .B(n16884), .Z(n16883) );
  XOR U16640 ( .A(p_input[1886]), .B(p_input[1870]), .Z(n16884) );
  XOR U16641 ( .A(n16885), .B(n16886), .Z(n16876) );
  AND U16642 ( .A(n16887), .B(n16888), .Z(n16886) );
  XOR U16643 ( .A(n16885), .B(n16718), .Z(n16888) );
  XNOR U16644 ( .A(p_input[1901]), .B(n16889), .Z(n16718) );
  AND U16645 ( .A(n623), .B(n16890), .Z(n16889) );
  XOR U16646 ( .A(p_input[1917]), .B(p_input[1901]), .Z(n16890) );
  XNOR U16647 ( .A(n16715), .B(n16885), .Z(n16887) );
  XOR U16648 ( .A(n16891), .B(n16892), .Z(n16715) );
  AND U16649 ( .A(n621), .B(n16893), .Z(n16892) );
  XOR U16650 ( .A(p_input[1885]), .B(p_input[1869]), .Z(n16893) );
  XOR U16651 ( .A(n16894), .B(n16895), .Z(n16885) );
  AND U16652 ( .A(n16896), .B(n16897), .Z(n16895) );
  XOR U16653 ( .A(n16894), .B(n16730), .Z(n16897) );
  XNOR U16654 ( .A(p_input[1900]), .B(n16898), .Z(n16730) );
  AND U16655 ( .A(n623), .B(n16899), .Z(n16898) );
  XOR U16656 ( .A(p_input[1916]), .B(p_input[1900]), .Z(n16899) );
  XNOR U16657 ( .A(n16727), .B(n16894), .Z(n16896) );
  XOR U16658 ( .A(n16900), .B(n16901), .Z(n16727) );
  AND U16659 ( .A(n621), .B(n16902), .Z(n16901) );
  XOR U16660 ( .A(p_input[1884]), .B(p_input[1868]), .Z(n16902) );
  XOR U16661 ( .A(n16903), .B(n16904), .Z(n16894) );
  AND U16662 ( .A(n16905), .B(n16906), .Z(n16904) );
  XOR U16663 ( .A(n16903), .B(n16742), .Z(n16906) );
  XNOR U16664 ( .A(p_input[1899]), .B(n16907), .Z(n16742) );
  AND U16665 ( .A(n623), .B(n16908), .Z(n16907) );
  XOR U16666 ( .A(p_input[1915]), .B(p_input[1899]), .Z(n16908) );
  XNOR U16667 ( .A(n16739), .B(n16903), .Z(n16905) );
  XOR U16668 ( .A(n16909), .B(n16910), .Z(n16739) );
  AND U16669 ( .A(n621), .B(n16911), .Z(n16910) );
  XOR U16670 ( .A(p_input[1883]), .B(p_input[1867]), .Z(n16911) );
  XOR U16671 ( .A(n16912), .B(n16913), .Z(n16903) );
  AND U16672 ( .A(n16914), .B(n16915), .Z(n16913) );
  XOR U16673 ( .A(n16912), .B(n16754), .Z(n16915) );
  XNOR U16674 ( .A(p_input[1898]), .B(n16916), .Z(n16754) );
  AND U16675 ( .A(n623), .B(n16917), .Z(n16916) );
  XOR U16676 ( .A(p_input[1914]), .B(p_input[1898]), .Z(n16917) );
  XNOR U16677 ( .A(n16751), .B(n16912), .Z(n16914) );
  XOR U16678 ( .A(n16918), .B(n16919), .Z(n16751) );
  AND U16679 ( .A(n621), .B(n16920), .Z(n16919) );
  XOR U16680 ( .A(p_input[1882]), .B(p_input[1866]), .Z(n16920) );
  XOR U16681 ( .A(n16921), .B(n16922), .Z(n16912) );
  AND U16682 ( .A(n16923), .B(n16924), .Z(n16922) );
  XOR U16683 ( .A(n16921), .B(n16766), .Z(n16924) );
  XNOR U16684 ( .A(p_input[1897]), .B(n16925), .Z(n16766) );
  AND U16685 ( .A(n623), .B(n16926), .Z(n16925) );
  XOR U16686 ( .A(p_input[1913]), .B(p_input[1897]), .Z(n16926) );
  XNOR U16687 ( .A(n16763), .B(n16921), .Z(n16923) );
  XOR U16688 ( .A(n16927), .B(n16928), .Z(n16763) );
  AND U16689 ( .A(n621), .B(n16929), .Z(n16928) );
  XOR U16690 ( .A(p_input[1881]), .B(p_input[1865]), .Z(n16929) );
  XOR U16691 ( .A(n16930), .B(n16931), .Z(n16921) );
  AND U16692 ( .A(n16932), .B(n16933), .Z(n16931) );
  XOR U16693 ( .A(n16930), .B(n16778), .Z(n16933) );
  XNOR U16694 ( .A(p_input[1896]), .B(n16934), .Z(n16778) );
  AND U16695 ( .A(n623), .B(n16935), .Z(n16934) );
  XOR U16696 ( .A(p_input[1912]), .B(p_input[1896]), .Z(n16935) );
  XNOR U16697 ( .A(n16775), .B(n16930), .Z(n16932) );
  XOR U16698 ( .A(n16936), .B(n16937), .Z(n16775) );
  AND U16699 ( .A(n621), .B(n16938), .Z(n16937) );
  XOR U16700 ( .A(p_input[1880]), .B(p_input[1864]), .Z(n16938) );
  XOR U16701 ( .A(n16939), .B(n16940), .Z(n16930) );
  AND U16702 ( .A(n16941), .B(n16942), .Z(n16940) );
  XOR U16703 ( .A(n16939), .B(n16790), .Z(n16942) );
  XNOR U16704 ( .A(p_input[1895]), .B(n16943), .Z(n16790) );
  AND U16705 ( .A(n623), .B(n16944), .Z(n16943) );
  XOR U16706 ( .A(p_input[1911]), .B(p_input[1895]), .Z(n16944) );
  XNOR U16707 ( .A(n16787), .B(n16939), .Z(n16941) );
  XOR U16708 ( .A(n16945), .B(n16946), .Z(n16787) );
  AND U16709 ( .A(n621), .B(n16947), .Z(n16946) );
  XOR U16710 ( .A(p_input[1879]), .B(p_input[1863]), .Z(n16947) );
  XOR U16711 ( .A(n16948), .B(n16949), .Z(n16939) );
  AND U16712 ( .A(n16950), .B(n16951), .Z(n16949) );
  XOR U16713 ( .A(n16948), .B(n16802), .Z(n16951) );
  XNOR U16714 ( .A(p_input[1894]), .B(n16952), .Z(n16802) );
  AND U16715 ( .A(n623), .B(n16953), .Z(n16952) );
  XOR U16716 ( .A(p_input[1910]), .B(p_input[1894]), .Z(n16953) );
  XNOR U16717 ( .A(n16799), .B(n16948), .Z(n16950) );
  XOR U16718 ( .A(n16954), .B(n16955), .Z(n16799) );
  AND U16719 ( .A(n621), .B(n16956), .Z(n16955) );
  XOR U16720 ( .A(p_input[1878]), .B(p_input[1862]), .Z(n16956) );
  XOR U16721 ( .A(n16957), .B(n16958), .Z(n16948) );
  AND U16722 ( .A(n16959), .B(n16960), .Z(n16958) );
  XOR U16723 ( .A(n16957), .B(n16814), .Z(n16960) );
  XNOR U16724 ( .A(p_input[1893]), .B(n16961), .Z(n16814) );
  AND U16725 ( .A(n623), .B(n16962), .Z(n16961) );
  XOR U16726 ( .A(p_input[1909]), .B(p_input[1893]), .Z(n16962) );
  XNOR U16727 ( .A(n16811), .B(n16957), .Z(n16959) );
  XOR U16728 ( .A(n16963), .B(n16964), .Z(n16811) );
  AND U16729 ( .A(n621), .B(n16965), .Z(n16964) );
  XOR U16730 ( .A(p_input[1877]), .B(p_input[1861]), .Z(n16965) );
  XOR U16731 ( .A(n16966), .B(n16967), .Z(n16957) );
  AND U16732 ( .A(n16968), .B(n16969), .Z(n16967) );
  XOR U16733 ( .A(n16966), .B(n16826), .Z(n16969) );
  XNOR U16734 ( .A(p_input[1892]), .B(n16970), .Z(n16826) );
  AND U16735 ( .A(n623), .B(n16971), .Z(n16970) );
  XOR U16736 ( .A(p_input[1908]), .B(p_input[1892]), .Z(n16971) );
  XNOR U16737 ( .A(n16823), .B(n16966), .Z(n16968) );
  XOR U16738 ( .A(n16972), .B(n16973), .Z(n16823) );
  AND U16739 ( .A(n621), .B(n16974), .Z(n16973) );
  XOR U16740 ( .A(p_input[1876]), .B(p_input[1860]), .Z(n16974) );
  XOR U16741 ( .A(n16975), .B(n16976), .Z(n16966) );
  AND U16742 ( .A(n16977), .B(n16978), .Z(n16976) );
  XOR U16743 ( .A(n16975), .B(n16838), .Z(n16978) );
  XNOR U16744 ( .A(p_input[1891]), .B(n16979), .Z(n16838) );
  AND U16745 ( .A(n623), .B(n16980), .Z(n16979) );
  XOR U16746 ( .A(p_input[1907]), .B(p_input[1891]), .Z(n16980) );
  XNOR U16747 ( .A(n16835), .B(n16975), .Z(n16977) );
  XOR U16748 ( .A(n16981), .B(n16982), .Z(n16835) );
  AND U16749 ( .A(n621), .B(n16983), .Z(n16982) );
  XOR U16750 ( .A(p_input[1875]), .B(p_input[1859]), .Z(n16983) );
  XOR U16751 ( .A(n16984), .B(n16985), .Z(n16975) );
  AND U16752 ( .A(n16986), .B(n16987), .Z(n16985) );
  XOR U16753 ( .A(n16984), .B(n16850), .Z(n16987) );
  XNOR U16754 ( .A(p_input[1890]), .B(n16988), .Z(n16850) );
  AND U16755 ( .A(n623), .B(n16989), .Z(n16988) );
  XOR U16756 ( .A(p_input[1906]), .B(p_input[1890]), .Z(n16989) );
  XNOR U16757 ( .A(n16847), .B(n16984), .Z(n16986) );
  XOR U16758 ( .A(n16990), .B(n16991), .Z(n16847) );
  AND U16759 ( .A(n621), .B(n16992), .Z(n16991) );
  XOR U16760 ( .A(p_input[1874]), .B(p_input[1858]), .Z(n16992) );
  XOR U16761 ( .A(n16993), .B(n16994), .Z(n16984) );
  AND U16762 ( .A(n16995), .B(n16996), .Z(n16994) );
  XNOR U16763 ( .A(n16997), .B(n16863), .Z(n16996) );
  XNOR U16764 ( .A(p_input[1889]), .B(n16998), .Z(n16863) );
  AND U16765 ( .A(n623), .B(n16999), .Z(n16998) );
  XNOR U16766 ( .A(p_input[1905]), .B(n17000), .Z(n16999) );
  IV U16767 ( .A(p_input[1889]), .Z(n17000) );
  XNOR U16768 ( .A(n16860), .B(n16993), .Z(n16995) );
  XNOR U16769 ( .A(p_input[1857]), .B(n17001), .Z(n16860) );
  AND U16770 ( .A(n621), .B(n17002), .Z(n17001) );
  XOR U16771 ( .A(p_input[1873]), .B(p_input[1857]), .Z(n17002) );
  IV U16772 ( .A(n16997), .Z(n16993) );
  AND U16773 ( .A(n16868), .B(n16871), .Z(n16997) );
  XOR U16774 ( .A(p_input[1888]), .B(n17003), .Z(n16871) );
  AND U16775 ( .A(n623), .B(n17004), .Z(n17003) );
  XOR U16776 ( .A(p_input[1904]), .B(p_input[1888]), .Z(n17004) );
  XOR U16777 ( .A(n17005), .B(n17006), .Z(n623) );
  AND U16778 ( .A(n17007), .B(n17008), .Z(n17006) );
  XNOR U16779 ( .A(p_input[1919]), .B(n17005), .Z(n17008) );
  XOR U16780 ( .A(n17005), .B(p_input[1903]), .Z(n17007) );
  XOR U16781 ( .A(n17009), .B(n17010), .Z(n17005) );
  AND U16782 ( .A(n17011), .B(n17012), .Z(n17010) );
  XNOR U16783 ( .A(p_input[1918]), .B(n17009), .Z(n17012) );
  XOR U16784 ( .A(n17009), .B(p_input[1902]), .Z(n17011) );
  XOR U16785 ( .A(n17013), .B(n17014), .Z(n17009) );
  AND U16786 ( .A(n17015), .B(n17016), .Z(n17014) );
  XNOR U16787 ( .A(p_input[1917]), .B(n17013), .Z(n17016) );
  XOR U16788 ( .A(n17013), .B(p_input[1901]), .Z(n17015) );
  XOR U16789 ( .A(n17017), .B(n17018), .Z(n17013) );
  AND U16790 ( .A(n17019), .B(n17020), .Z(n17018) );
  XNOR U16791 ( .A(p_input[1916]), .B(n17017), .Z(n17020) );
  XOR U16792 ( .A(n17017), .B(p_input[1900]), .Z(n17019) );
  XOR U16793 ( .A(n17021), .B(n17022), .Z(n17017) );
  AND U16794 ( .A(n17023), .B(n17024), .Z(n17022) );
  XNOR U16795 ( .A(p_input[1915]), .B(n17021), .Z(n17024) );
  XOR U16796 ( .A(n17021), .B(p_input[1899]), .Z(n17023) );
  XOR U16797 ( .A(n17025), .B(n17026), .Z(n17021) );
  AND U16798 ( .A(n17027), .B(n17028), .Z(n17026) );
  XNOR U16799 ( .A(p_input[1914]), .B(n17025), .Z(n17028) );
  XOR U16800 ( .A(n17025), .B(p_input[1898]), .Z(n17027) );
  XOR U16801 ( .A(n17029), .B(n17030), .Z(n17025) );
  AND U16802 ( .A(n17031), .B(n17032), .Z(n17030) );
  XNOR U16803 ( .A(p_input[1913]), .B(n17029), .Z(n17032) );
  XOR U16804 ( .A(n17029), .B(p_input[1897]), .Z(n17031) );
  XOR U16805 ( .A(n17033), .B(n17034), .Z(n17029) );
  AND U16806 ( .A(n17035), .B(n17036), .Z(n17034) );
  XNOR U16807 ( .A(p_input[1912]), .B(n17033), .Z(n17036) );
  XOR U16808 ( .A(n17033), .B(p_input[1896]), .Z(n17035) );
  XOR U16809 ( .A(n17037), .B(n17038), .Z(n17033) );
  AND U16810 ( .A(n17039), .B(n17040), .Z(n17038) );
  XNOR U16811 ( .A(p_input[1911]), .B(n17037), .Z(n17040) );
  XOR U16812 ( .A(n17037), .B(p_input[1895]), .Z(n17039) );
  XOR U16813 ( .A(n17041), .B(n17042), .Z(n17037) );
  AND U16814 ( .A(n17043), .B(n17044), .Z(n17042) );
  XNOR U16815 ( .A(p_input[1910]), .B(n17041), .Z(n17044) );
  XOR U16816 ( .A(n17041), .B(p_input[1894]), .Z(n17043) );
  XOR U16817 ( .A(n17045), .B(n17046), .Z(n17041) );
  AND U16818 ( .A(n17047), .B(n17048), .Z(n17046) );
  XNOR U16819 ( .A(p_input[1909]), .B(n17045), .Z(n17048) );
  XOR U16820 ( .A(n17045), .B(p_input[1893]), .Z(n17047) );
  XOR U16821 ( .A(n17049), .B(n17050), .Z(n17045) );
  AND U16822 ( .A(n17051), .B(n17052), .Z(n17050) );
  XNOR U16823 ( .A(p_input[1908]), .B(n17049), .Z(n17052) );
  XOR U16824 ( .A(n17049), .B(p_input[1892]), .Z(n17051) );
  XOR U16825 ( .A(n17053), .B(n17054), .Z(n17049) );
  AND U16826 ( .A(n17055), .B(n17056), .Z(n17054) );
  XNOR U16827 ( .A(p_input[1907]), .B(n17053), .Z(n17056) );
  XOR U16828 ( .A(n17053), .B(p_input[1891]), .Z(n17055) );
  XOR U16829 ( .A(n17057), .B(n17058), .Z(n17053) );
  AND U16830 ( .A(n17059), .B(n17060), .Z(n17058) );
  XNOR U16831 ( .A(p_input[1906]), .B(n17057), .Z(n17060) );
  XOR U16832 ( .A(n17057), .B(p_input[1890]), .Z(n17059) );
  XNOR U16833 ( .A(n17061), .B(n17062), .Z(n17057) );
  AND U16834 ( .A(n17063), .B(n17064), .Z(n17062) );
  XOR U16835 ( .A(p_input[1905]), .B(n17061), .Z(n17064) );
  XNOR U16836 ( .A(p_input[1889]), .B(n17061), .Z(n17063) );
  AND U16837 ( .A(p_input[1904]), .B(n17065), .Z(n17061) );
  IV U16838 ( .A(p_input[1888]), .Z(n17065) );
  XNOR U16839 ( .A(p_input[1856]), .B(n17066), .Z(n16868) );
  AND U16840 ( .A(n621), .B(n17067), .Z(n17066) );
  XOR U16841 ( .A(p_input[1872]), .B(p_input[1856]), .Z(n17067) );
  XOR U16842 ( .A(n17068), .B(n17069), .Z(n621) );
  AND U16843 ( .A(n17070), .B(n17071), .Z(n17069) );
  XNOR U16844 ( .A(p_input[1887]), .B(n17068), .Z(n17071) );
  XOR U16845 ( .A(n17068), .B(p_input[1871]), .Z(n17070) );
  XOR U16846 ( .A(n17072), .B(n17073), .Z(n17068) );
  AND U16847 ( .A(n17074), .B(n17075), .Z(n17073) );
  XNOR U16848 ( .A(p_input[1886]), .B(n17072), .Z(n17075) );
  XNOR U16849 ( .A(n17072), .B(n16882), .Z(n17074) );
  IV U16850 ( .A(p_input[1870]), .Z(n16882) );
  XOR U16851 ( .A(n17076), .B(n17077), .Z(n17072) );
  AND U16852 ( .A(n17078), .B(n17079), .Z(n17077) );
  XNOR U16853 ( .A(p_input[1885]), .B(n17076), .Z(n17079) );
  XNOR U16854 ( .A(n17076), .B(n16891), .Z(n17078) );
  IV U16855 ( .A(p_input[1869]), .Z(n16891) );
  XOR U16856 ( .A(n17080), .B(n17081), .Z(n17076) );
  AND U16857 ( .A(n17082), .B(n17083), .Z(n17081) );
  XNOR U16858 ( .A(p_input[1884]), .B(n17080), .Z(n17083) );
  XNOR U16859 ( .A(n17080), .B(n16900), .Z(n17082) );
  IV U16860 ( .A(p_input[1868]), .Z(n16900) );
  XOR U16861 ( .A(n17084), .B(n17085), .Z(n17080) );
  AND U16862 ( .A(n17086), .B(n17087), .Z(n17085) );
  XNOR U16863 ( .A(p_input[1883]), .B(n17084), .Z(n17087) );
  XNOR U16864 ( .A(n17084), .B(n16909), .Z(n17086) );
  IV U16865 ( .A(p_input[1867]), .Z(n16909) );
  XOR U16866 ( .A(n17088), .B(n17089), .Z(n17084) );
  AND U16867 ( .A(n17090), .B(n17091), .Z(n17089) );
  XNOR U16868 ( .A(p_input[1882]), .B(n17088), .Z(n17091) );
  XNOR U16869 ( .A(n17088), .B(n16918), .Z(n17090) );
  IV U16870 ( .A(p_input[1866]), .Z(n16918) );
  XOR U16871 ( .A(n17092), .B(n17093), .Z(n17088) );
  AND U16872 ( .A(n17094), .B(n17095), .Z(n17093) );
  XNOR U16873 ( .A(p_input[1881]), .B(n17092), .Z(n17095) );
  XNOR U16874 ( .A(n17092), .B(n16927), .Z(n17094) );
  IV U16875 ( .A(p_input[1865]), .Z(n16927) );
  XOR U16876 ( .A(n17096), .B(n17097), .Z(n17092) );
  AND U16877 ( .A(n17098), .B(n17099), .Z(n17097) );
  XNOR U16878 ( .A(p_input[1880]), .B(n17096), .Z(n17099) );
  XNOR U16879 ( .A(n17096), .B(n16936), .Z(n17098) );
  IV U16880 ( .A(p_input[1864]), .Z(n16936) );
  XOR U16881 ( .A(n17100), .B(n17101), .Z(n17096) );
  AND U16882 ( .A(n17102), .B(n17103), .Z(n17101) );
  XNOR U16883 ( .A(p_input[1879]), .B(n17100), .Z(n17103) );
  XNOR U16884 ( .A(n17100), .B(n16945), .Z(n17102) );
  IV U16885 ( .A(p_input[1863]), .Z(n16945) );
  XOR U16886 ( .A(n17104), .B(n17105), .Z(n17100) );
  AND U16887 ( .A(n17106), .B(n17107), .Z(n17105) );
  XNOR U16888 ( .A(p_input[1878]), .B(n17104), .Z(n17107) );
  XNOR U16889 ( .A(n17104), .B(n16954), .Z(n17106) );
  IV U16890 ( .A(p_input[1862]), .Z(n16954) );
  XOR U16891 ( .A(n17108), .B(n17109), .Z(n17104) );
  AND U16892 ( .A(n17110), .B(n17111), .Z(n17109) );
  XNOR U16893 ( .A(p_input[1877]), .B(n17108), .Z(n17111) );
  XNOR U16894 ( .A(n17108), .B(n16963), .Z(n17110) );
  IV U16895 ( .A(p_input[1861]), .Z(n16963) );
  XOR U16896 ( .A(n17112), .B(n17113), .Z(n17108) );
  AND U16897 ( .A(n17114), .B(n17115), .Z(n17113) );
  XNOR U16898 ( .A(p_input[1876]), .B(n17112), .Z(n17115) );
  XNOR U16899 ( .A(n17112), .B(n16972), .Z(n17114) );
  IV U16900 ( .A(p_input[1860]), .Z(n16972) );
  XOR U16901 ( .A(n17116), .B(n17117), .Z(n17112) );
  AND U16902 ( .A(n17118), .B(n17119), .Z(n17117) );
  XNOR U16903 ( .A(p_input[1875]), .B(n17116), .Z(n17119) );
  XNOR U16904 ( .A(n17116), .B(n16981), .Z(n17118) );
  IV U16905 ( .A(p_input[1859]), .Z(n16981) );
  XOR U16906 ( .A(n17120), .B(n17121), .Z(n17116) );
  AND U16907 ( .A(n17122), .B(n17123), .Z(n17121) );
  XNOR U16908 ( .A(p_input[1874]), .B(n17120), .Z(n17123) );
  XNOR U16909 ( .A(n17120), .B(n16990), .Z(n17122) );
  IV U16910 ( .A(p_input[1858]), .Z(n16990) );
  XNOR U16911 ( .A(n17124), .B(n17125), .Z(n17120) );
  AND U16912 ( .A(n17126), .B(n17127), .Z(n17125) );
  XOR U16913 ( .A(p_input[1873]), .B(n17124), .Z(n17127) );
  XNOR U16914 ( .A(p_input[1857]), .B(n17124), .Z(n17126) );
  AND U16915 ( .A(p_input[1872]), .B(n17128), .Z(n17124) );
  IV U16916 ( .A(p_input[1856]), .Z(n17128) );
  XOR U16917 ( .A(n17129), .B(n17130), .Z(n16687) );
  AND U16918 ( .A(n484), .B(n17131), .Z(n17130) );
  XNOR U16919 ( .A(n17132), .B(n17129), .Z(n17131) );
  XOR U16920 ( .A(n17133), .B(n17134), .Z(n484) );
  AND U16921 ( .A(n17135), .B(n17136), .Z(n17134) );
  XNOR U16922 ( .A(n16698), .B(n17133), .Z(n17136) );
  AND U16923 ( .A(p_input[1855]), .B(p_input[1839]), .Z(n16698) );
  XOR U16924 ( .A(n17133), .B(n16697), .Z(n17135) );
  AND U16925 ( .A(p_input[1807]), .B(p_input[1823]), .Z(n16697) );
  XOR U16926 ( .A(n17137), .B(n17138), .Z(n17133) );
  AND U16927 ( .A(n17139), .B(n17140), .Z(n17138) );
  XOR U16928 ( .A(n17137), .B(n16710), .Z(n17140) );
  XNOR U16929 ( .A(p_input[1838]), .B(n17141), .Z(n16710) );
  AND U16930 ( .A(n627), .B(n17142), .Z(n17141) );
  XOR U16931 ( .A(p_input[1854]), .B(p_input[1838]), .Z(n17142) );
  XNOR U16932 ( .A(n16707), .B(n17137), .Z(n17139) );
  XOR U16933 ( .A(n17143), .B(n17144), .Z(n16707) );
  AND U16934 ( .A(n624), .B(n17145), .Z(n17144) );
  XOR U16935 ( .A(p_input[1822]), .B(p_input[1806]), .Z(n17145) );
  XOR U16936 ( .A(n17146), .B(n17147), .Z(n17137) );
  AND U16937 ( .A(n17148), .B(n17149), .Z(n17147) );
  XOR U16938 ( .A(n17146), .B(n16722), .Z(n17149) );
  XNOR U16939 ( .A(p_input[1837]), .B(n17150), .Z(n16722) );
  AND U16940 ( .A(n627), .B(n17151), .Z(n17150) );
  XOR U16941 ( .A(p_input[1853]), .B(p_input[1837]), .Z(n17151) );
  XNOR U16942 ( .A(n16719), .B(n17146), .Z(n17148) );
  XOR U16943 ( .A(n17152), .B(n17153), .Z(n16719) );
  AND U16944 ( .A(n624), .B(n17154), .Z(n17153) );
  XOR U16945 ( .A(p_input[1821]), .B(p_input[1805]), .Z(n17154) );
  XOR U16946 ( .A(n17155), .B(n17156), .Z(n17146) );
  AND U16947 ( .A(n17157), .B(n17158), .Z(n17156) );
  XOR U16948 ( .A(n17155), .B(n16734), .Z(n17158) );
  XNOR U16949 ( .A(p_input[1836]), .B(n17159), .Z(n16734) );
  AND U16950 ( .A(n627), .B(n17160), .Z(n17159) );
  XOR U16951 ( .A(p_input[1852]), .B(p_input[1836]), .Z(n17160) );
  XNOR U16952 ( .A(n16731), .B(n17155), .Z(n17157) );
  XOR U16953 ( .A(n17161), .B(n17162), .Z(n16731) );
  AND U16954 ( .A(n624), .B(n17163), .Z(n17162) );
  XOR U16955 ( .A(p_input[1820]), .B(p_input[1804]), .Z(n17163) );
  XOR U16956 ( .A(n17164), .B(n17165), .Z(n17155) );
  AND U16957 ( .A(n17166), .B(n17167), .Z(n17165) );
  XOR U16958 ( .A(n17164), .B(n16746), .Z(n17167) );
  XNOR U16959 ( .A(p_input[1835]), .B(n17168), .Z(n16746) );
  AND U16960 ( .A(n627), .B(n17169), .Z(n17168) );
  XOR U16961 ( .A(p_input[1851]), .B(p_input[1835]), .Z(n17169) );
  XNOR U16962 ( .A(n16743), .B(n17164), .Z(n17166) );
  XOR U16963 ( .A(n17170), .B(n17171), .Z(n16743) );
  AND U16964 ( .A(n624), .B(n17172), .Z(n17171) );
  XOR U16965 ( .A(p_input[1819]), .B(p_input[1803]), .Z(n17172) );
  XOR U16966 ( .A(n17173), .B(n17174), .Z(n17164) );
  AND U16967 ( .A(n17175), .B(n17176), .Z(n17174) );
  XOR U16968 ( .A(n17173), .B(n16758), .Z(n17176) );
  XNOR U16969 ( .A(p_input[1834]), .B(n17177), .Z(n16758) );
  AND U16970 ( .A(n627), .B(n17178), .Z(n17177) );
  XOR U16971 ( .A(p_input[1850]), .B(p_input[1834]), .Z(n17178) );
  XNOR U16972 ( .A(n16755), .B(n17173), .Z(n17175) );
  XOR U16973 ( .A(n17179), .B(n17180), .Z(n16755) );
  AND U16974 ( .A(n624), .B(n17181), .Z(n17180) );
  XOR U16975 ( .A(p_input[1818]), .B(p_input[1802]), .Z(n17181) );
  XOR U16976 ( .A(n17182), .B(n17183), .Z(n17173) );
  AND U16977 ( .A(n17184), .B(n17185), .Z(n17183) );
  XOR U16978 ( .A(n17182), .B(n16770), .Z(n17185) );
  XNOR U16979 ( .A(p_input[1833]), .B(n17186), .Z(n16770) );
  AND U16980 ( .A(n627), .B(n17187), .Z(n17186) );
  XOR U16981 ( .A(p_input[1849]), .B(p_input[1833]), .Z(n17187) );
  XNOR U16982 ( .A(n16767), .B(n17182), .Z(n17184) );
  XOR U16983 ( .A(n17188), .B(n17189), .Z(n16767) );
  AND U16984 ( .A(n624), .B(n17190), .Z(n17189) );
  XOR U16985 ( .A(p_input[1817]), .B(p_input[1801]), .Z(n17190) );
  XOR U16986 ( .A(n17191), .B(n17192), .Z(n17182) );
  AND U16987 ( .A(n17193), .B(n17194), .Z(n17192) );
  XOR U16988 ( .A(n17191), .B(n16782), .Z(n17194) );
  XNOR U16989 ( .A(p_input[1832]), .B(n17195), .Z(n16782) );
  AND U16990 ( .A(n627), .B(n17196), .Z(n17195) );
  XOR U16991 ( .A(p_input[1848]), .B(p_input[1832]), .Z(n17196) );
  XNOR U16992 ( .A(n16779), .B(n17191), .Z(n17193) );
  XOR U16993 ( .A(n17197), .B(n17198), .Z(n16779) );
  AND U16994 ( .A(n624), .B(n17199), .Z(n17198) );
  XOR U16995 ( .A(p_input[1816]), .B(p_input[1800]), .Z(n17199) );
  XOR U16996 ( .A(n17200), .B(n17201), .Z(n17191) );
  AND U16997 ( .A(n17202), .B(n17203), .Z(n17201) );
  XOR U16998 ( .A(n17200), .B(n16794), .Z(n17203) );
  XNOR U16999 ( .A(p_input[1831]), .B(n17204), .Z(n16794) );
  AND U17000 ( .A(n627), .B(n17205), .Z(n17204) );
  XOR U17001 ( .A(p_input[1847]), .B(p_input[1831]), .Z(n17205) );
  XNOR U17002 ( .A(n16791), .B(n17200), .Z(n17202) );
  XOR U17003 ( .A(n17206), .B(n17207), .Z(n16791) );
  AND U17004 ( .A(n624), .B(n17208), .Z(n17207) );
  XOR U17005 ( .A(p_input[1815]), .B(p_input[1799]), .Z(n17208) );
  XOR U17006 ( .A(n17209), .B(n17210), .Z(n17200) );
  AND U17007 ( .A(n17211), .B(n17212), .Z(n17210) );
  XOR U17008 ( .A(n17209), .B(n16806), .Z(n17212) );
  XNOR U17009 ( .A(p_input[1830]), .B(n17213), .Z(n16806) );
  AND U17010 ( .A(n627), .B(n17214), .Z(n17213) );
  XOR U17011 ( .A(p_input[1846]), .B(p_input[1830]), .Z(n17214) );
  XNOR U17012 ( .A(n16803), .B(n17209), .Z(n17211) );
  XOR U17013 ( .A(n17215), .B(n17216), .Z(n16803) );
  AND U17014 ( .A(n624), .B(n17217), .Z(n17216) );
  XOR U17015 ( .A(p_input[1814]), .B(p_input[1798]), .Z(n17217) );
  XOR U17016 ( .A(n17218), .B(n17219), .Z(n17209) );
  AND U17017 ( .A(n17220), .B(n17221), .Z(n17219) );
  XOR U17018 ( .A(n17218), .B(n16818), .Z(n17221) );
  XNOR U17019 ( .A(p_input[1829]), .B(n17222), .Z(n16818) );
  AND U17020 ( .A(n627), .B(n17223), .Z(n17222) );
  XOR U17021 ( .A(p_input[1845]), .B(p_input[1829]), .Z(n17223) );
  XNOR U17022 ( .A(n16815), .B(n17218), .Z(n17220) );
  XOR U17023 ( .A(n17224), .B(n17225), .Z(n16815) );
  AND U17024 ( .A(n624), .B(n17226), .Z(n17225) );
  XOR U17025 ( .A(p_input[1813]), .B(p_input[1797]), .Z(n17226) );
  XOR U17026 ( .A(n17227), .B(n17228), .Z(n17218) );
  AND U17027 ( .A(n17229), .B(n17230), .Z(n17228) );
  XOR U17028 ( .A(n17227), .B(n16830), .Z(n17230) );
  XNOR U17029 ( .A(p_input[1828]), .B(n17231), .Z(n16830) );
  AND U17030 ( .A(n627), .B(n17232), .Z(n17231) );
  XOR U17031 ( .A(p_input[1844]), .B(p_input[1828]), .Z(n17232) );
  XNOR U17032 ( .A(n16827), .B(n17227), .Z(n17229) );
  XOR U17033 ( .A(n17233), .B(n17234), .Z(n16827) );
  AND U17034 ( .A(n624), .B(n17235), .Z(n17234) );
  XOR U17035 ( .A(p_input[1812]), .B(p_input[1796]), .Z(n17235) );
  XOR U17036 ( .A(n17236), .B(n17237), .Z(n17227) );
  AND U17037 ( .A(n17238), .B(n17239), .Z(n17237) );
  XOR U17038 ( .A(n17236), .B(n16842), .Z(n17239) );
  XNOR U17039 ( .A(p_input[1827]), .B(n17240), .Z(n16842) );
  AND U17040 ( .A(n627), .B(n17241), .Z(n17240) );
  XOR U17041 ( .A(p_input[1843]), .B(p_input[1827]), .Z(n17241) );
  XNOR U17042 ( .A(n16839), .B(n17236), .Z(n17238) );
  XOR U17043 ( .A(n17242), .B(n17243), .Z(n16839) );
  AND U17044 ( .A(n624), .B(n17244), .Z(n17243) );
  XOR U17045 ( .A(p_input[1811]), .B(p_input[1795]), .Z(n17244) );
  XOR U17046 ( .A(n17245), .B(n17246), .Z(n17236) );
  AND U17047 ( .A(n17247), .B(n17248), .Z(n17246) );
  XOR U17048 ( .A(n17245), .B(n16854), .Z(n17248) );
  XNOR U17049 ( .A(p_input[1826]), .B(n17249), .Z(n16854) );
  AND U17050 ( .A(n627), .B(n17250), .Z(n17249) );
  XOR U17051 ( .A(p_input[1842]), .B(p_input[1826]), .Z(n17250) );
  XNOR U17052 ( .A(n16851), .B(n17245), .Z(n17247) );
  XOR U17053 ( .A(n17251), .B(n17252), .Z(n16851) );
  AND U17054 ( .A(n624), .B(n17253), .Z(n17252) );
  XOR U17055 ( .A(p_input[1810]), .B(p_input[1794]), .Z(n17253) );
  XOR U17056 ( .A(n17254), .B(n17255), .Z(n17245) );
  AND U17057 ( .A(n17256), .B(n17257), .Z(n17255) );
  XNOR U17058 ( .A(n17258), .B(n16867), .Z(n17257) );
  XNOR U17059 ( .A(p_input[1825]), .B(n17259), .Z(n16867) );
  AND U17060 ( .A(n627), .B(n17260), .Z(n17259) );
  XNOR U17061 ( .A(p_input[1841]), .B(n17261), .Z(n17260) );
  IV U17062 ( .A(p_input[1825]), .Z(n17261) );
  XNOR U17063 ( .A(n16864), .B(n17254), .Z(n17256) );
  XNOR U17064 ( .A(p_input[1793]), .B(n17262), .Z(n16864) );
  AND U17065 ( .A(n624), .B(n17263), .Z(n17262) );
  XOR U17066 ( .A(p_input[1809]), .B(p_input[1793]), .Z(n17263) );
  IV U17067 ( .A(n17258), .Z(n17254) );
  AND U17068 ( .A(n17129), .B(n17132), .Z(n17258) );
  XOR U17069 ( .A(p_input[1824]), .B(n17264), .Z(n17132) );
  AND U17070 ( .A(n627), .B(n17265), .Z(n17264) );
  XOR U17071 ( .A(p_input[1840]), .B(p_input[1824]), .Z(n17265) );
  XOR U17072 ( .A(n17266), .B(n17267), .Z(n627) );
  AND U17073 ( .A(n17268), .B(n17269), .Z(n17267) );
  XNOR U17074 ( .A(p_input[1855]), .B(n17266), .Z(n17269) );
  XOR U17075 ( .A(n17266), .B(p_input[1839]), .Z(n17268) );
  XOR U17076 ( .A(n17270), .B(n17271), .Z(n17266) );
  AND U17077 ( .A(n17272), .B(n17273), .Z(n17271) );
  XNOR U17078 ( .A(p_input[1854]), .B(n17270), .Z(n17273) );
  XOR U17079 ( .A(n17270), .B(p_input[1838]), .Z(n17272) );
  XOR U17080 ( .A(n17274), .B(n17275), .Z(n17270) );
  AND U17081 ( .A(n17276), .B(n17277), .Z(n17275) );
  XNOR U17082 ( .A(p_input[1853]), .B(n17274), .Z(n17277) );
  XOR U17083 ( .A(n17274), .B(p_input[1837]), .Z(n17276) );
  XOR U17084 ( .A(n17278), .B(n17279), .Z(n17274) );
  AND U17085 ( .A(n17280), .B(n17281), .Z(n17279) );
  XNOR U17086 ( .A(p_input[1852]), .B(n17278), .Z(n17281) );
  XOR U17087 ( .A(n17278), .B(p_input[1836]), .Z(n17280) );
  XOR U17088 ( .A(n17282), .B(n17283), .Z(n17278) );
  AND U17089 ( .A(n17284), .B(n17285), .Z(n17283) );
  XNOR U17090 ( .A(p_input[1851]), .B(n17282), .Z(n17285) );
  XOR U17091 ( .A(n17282), .B(p_input[1835]), .Z(n17284) );
  XOR U17092 ( .A(n17286), .B(n17287), .Z(n17282) );
  AND U17093 ( .A(n17288), .B(n17289), .Z(n17287) );
  XNOR U17094 ( .A(p_input[1850]), .B(n17286), .Z(n17289) );
  XOR U17095 ( .A(n17286), .B(p_input[1834]), .Z(n17288) );
  XOR U17096 ( .A(n17290), .B(n17291), .Z(n17286) );
  AND U17097 ( .A(n17292), .B(n17293), .Z(n17291) );
  XNOR U17098 ( .A(p_input[1849]), .B(n17290), .Z(n17293) );
  XOR U17099 ( .A(n17290), .B(p_input[1833]), .Z(n17292) );
  XOR U17100 ( .A(n17294), .B(n17295), .Z(n17290) );
  AND U17101 ( .A(n17296), .B(n17297), .Z(n17295) );
  XNOR U17102 ( .A(p_input[1848]), .B(n17294), .Z(n17297) );
  XOR U17103 ( .A(n17294), .B(p_input[1832]), .Z(n17296) );
  XOR U17104 ( .A(n17298), .B(n17299), .Z(n17294) );
  AND U17105 ( .A(n17300), .B(n17301), .Z(n17299) );
  XNOR U17106 ( .A(p_input[1847]), .B(n17298), .Z(n17301) );
  XOR U17107 ( .A(n17298), .B(p_input[1831]), .Z(n17300) );
  XOR U17108 ( .A(n17302), .B(n17303), .Z(n17298) );
  AND U17109 ( .A(n17304), .B(n17305), .Z(n17303) );
  XNOR U17110 ( .A(p_input[1846]), .B(n17302), .Z(n17305) );
  XOR U17111 ( .A(n17302), .B(p_input[1830]), .Z(n17304) );
  XOR U17112 ( .A(n17306), .B(n17307), .Z(n17302) );
  AND U17113 ( .A(n17308), .B(n17309), .Z(n17307) );
  XNOR U17114 ( .A(p_input[1845]), .B(n17306), .Z(n17309) );
  XOR U17115 ( .A(n17306), .B(p_input[1829]), .Z(n17308) );
  XOR U17116 ( .A(n17310), .B(n17311), .Z(n17306) );
  AND U17117 ( .A(n17312), .B(n17313), .Z(n17311) );
  XNOR U17118 ( .A(p_input[1844]), .B(n17310), .Z(n17313) );
  XOR U17119 ( .A(n17310), .B(p_input[1828]), .Z(n17312) );
  XOR U17120 ( .A(n17314), .B(n17315), .Z(n17310) );
  AND U17121 ( .A(n17316), .B(n17317), .Z(n17315) );
  XNOR U17122 ( .A(p_input[1843]), .B(n17314), .Z(n17317) );
  XOR U17123 ( .A(n17314), .B(p_input[1827]), .Z(n17316) );
  XOR U17124 ( .A(n17318), .B(n17319), .Z(n17314) );
  AND U17125 ( .A(n17320), .B(n17321), .Z(n17319) );
  XNOR U17126 ( .A(p_input[1842]), .B(n17318), .Z(n17321) );
  XOR U17127 ( .A(n17318), .B(p_input[1826]), .Z(n17320) );
  XNOR U17128 ( .A(n17322), .B(n17323), .Z(n17318) );
  AND U17129 ( .A(n17324), .B(n17325), .Z(n17323) );
  XOR U17130 ( .A(p_input[1841]), .B(n17322), .Z(n17325) );
  XNOR U17131 ( .A(p_input[1825]), .B(n17322), .Z(n17324) );
  AND U17132 ( .A(p_input[1840]), .B(n17326), .Z(n17322) );
  IV U17133 ( .A(p_input[1824]), .Z(n17326) );
  XNOR U17134 ( .A(p_input[1792]), .B(n17327), .Z(n17129) );
  AND U17135 ( .A(n624), .B(n17328), .Z(n17327) );
  XOR U17136 ( .A(p_input[1808]), .B(p_input[1792]), .Z(n17328) );
  XOR U17137 ( .A(n17329), .B(n17330), .Z(n624) );
  AND U17138 ( .A(n17331), .B(n17332), .Z(n17330) );
  XNOR U17139 ( .A(p_input[1823]), .B(n17329), .Z(n17332) );
  XOR U17140 ( .A(n17329), .B(p_input[1807]), .Z(n17331) );
  XOR U17141 ( .A(n17333), .B(n17334), .Z(n17329) );
  AND U17142 ( .A(n17335), .B(n17336), .Z(n17334) );
  XNOR U17143 ( .A(p_input[1822]), .B(n17333), .Z(n17336) );
  XNOR U17144 ( .A(n17333), .B(n17143), .Z(n17335) );
  IV U17145 ( .A(p_input[1806]), .Z(n17143) );
  XOR U17146 ( .A(n17337), .B(n17338), .Z(n17333) );
  AND U17147 ( .A(n17339), .B(n17340), .Z(n17338) );
  XNOR U17148 ( .A(p_input[1821]), .B(n17337), .Z(n17340) );
  XNOR U17149 ( .A(n17337), .B(n17152), .Z(n17339) );
  IV U17150 ( .A(p_input[1805]), .Z(n17152) );
  XOR U17151 ( .A(n17341), .B(n17342), .Z(n17337) );
  AND U17152 ( .A(n17343), .B(n17344), .Z(n17342) );
  XNOR U17153 ( .A(p_input[1820]), .B(n17341), .Z(n17344) );
  XNOR U17154 ( .A(n17341), .B(n17161), .Z(n17343) );
  IV U17155 ( .A(p_input[1804]), .Z(n17161) );
  XOR U17156 ( .A(n17345), .B(n17346), .Z(n17341) );
  AND U17157 ( .A(n17347), .B(n17348), .Z(n17346) );
  XNOR U17158 ( .A(p_input[1819]), .B(n17345), .Z(n17348) );
  XNOR U17159 ( .A(n17345), .B(n17170), .Z(n17347) );
  IV U17160 ( .A(p_input[1803]), .Z(n17170) );
  XOR U17161 ( .A(n17349), .B(n17350), .Z(n17345) );
  AND U17162 ( .A(n17351), .B(n17352), .Z(n17350) );
  XNOR U17163 ( .A(p_input[1818]), .B(n17349), .Z(n17352) );
  XNOR U17164 ( .A(n17349), .B(n17179), .Z(n17351) );
  IV U17165 ( .A(p_input[1802]), .Z(n17179) );
  XOR U17166 ( .A(n17353), .B(n17354), .Z(n17349) );
  AND U17167 ( .A(n17355), .B(n17356), .Z(n17354) );
  XNOR U17168 ( .A(p_input[1817]), .B(n17353), .Z(n17356) );
  XNOR U17169 ( .A(n17353), .B(n17188), .Z(n17355) );
  IV U17170 ( .A(p_input[1801]), .Z(n17188) );
  XOR U17171 ( .A(n17357), .B(n17358), .Z(n17353) );
  AND U17172 ( .A(n17359), .B(n17360), .Z(n17358) );
  XNOR U17173 ( .A(p_input[1816]), .B(n17357), .Z(n17360) );
  XNOR U17174 ( .A(n17357), .B(n17197), .Z(n17359) );
  IV U17175 ( .A(p_input[1800]), .Z(n17197) );
  XOR U17176 ( .A(n17361), .B(n17362), .Z(n17357) );
  AND U17177 ( .A(n17363), .B(n17364), .Z(n17362) );
  XNOR U17178 ( .A(p_input[1815]), .B(n17361), .Z(n17364) );
  XNOR U17179 ( .A(n17361), .B(n17206), .Z(n17363) );
  IV U17180 ( .A(p_input[1799]), .Z(n17206) );
  XOR U17181 ( .A(n17365), .B(n17366), .Z(n17361) );
  AND U17182 ( .A(n17367), .B(n17368), .Z(n17366) );
  XNOR U17183 ( .A(p_input[1814]), .B(n17365), .Z(n17368) );
  XNOR U17184 ( .A(n17365), .B(n17215), .Z(n17367) );
  IV U17185 ( .A(p_input[1798]), .Z(n17215) );
  XOR U17186 ( .A(n17369), .B(n17370), .Z(n17365) );
  AND U17187 ( .A(n17371), .B(n17372), .Z(n17370) );
  XNOR U17188 ( .A(p_input[1813]), .B(n17369), .Z(n17372) );
  XNOR U17189 ( .A(n17369), .B(n17224), .Z(n17371) );
  IV U17190 ( .A(p_input[1797]), .Z(n17224) );
  XOR U17191 ( .A(n17373), .B(n17374), .Z(n17369) );
  AND U17192 ( .A(n17375), .B(n17376), .Z(n17374) );
  XNOR U17193 ( .A(p_input[1812]), .B(n17373), .Z(n17376) );
  XNOR U17194 ( .A(n17373), .B(n17233), .Z(n17375) );
  IV U17195 ( .A(p_input[1796]), .Z(n17233) );
  XOR U17196 ( .A(n17377), .B(n17378), .Z(n17373) );
  AND U17197 ( .A(n17379), .B(n17380), .Z(n17378) );
  XNOR U17198 ( .A(p_input[1811]), .B(n17377), .Z(n17380) );
  XNOR U17199 ( .A(n17377), .B(n17242), .Z(n17379) );
  IV U17200 ( .A(p_input[1795]), .Z(n17242) );
  XOR U17201 ( .A(n17381), .B(n17382), .Z(n17377) );
  AND U17202 ( .A(n17383), .B(n17384), .Z(n17382) );
  XNOR U17203 ( .A(p_input[1810]), .B(n17381), .Z(n17384) );
  XNOR U17204 ( .A(n17381), .B(n17251), .Z(n17383) );
  IV U17205 ( .A(p_input[1794]), .Z(n17251) );
  XNOR U17206 ( .A(n17385), .B(n17386), .Z(n17381) );
  AND U17207 ( .A(n17387), .B(n17388), .Z(n17386) );
  XOR U17208 ( .A(p_input[1809]), .B(n17385), .Z(n17388) );
  XNOR U17209 ( .A(p_input[1793]), .B(n17385), .Z(n17387) );
  AND U17210 ( .A(p_input[1808]), .B(n17389), .Z(n17385) );
  IV U17211 ( .A(p_input[1792]), .Z(n17389) );
  XOR U17212 ( .A(n17390), .B(n17391), .Z(n15617) );
  AND U17213 ( .A(n945), .B(n17392), .Z(n17391) );
  XNOR U17214 ( .A(n17393), .B(n17390), .Z(n17392) );
  XOR U17215 ( .A(n17394), .B(n17395), .Z(n945) );
  AND U17216 ( .A(n17396), .B(n17397), .Z(n17395) );
  XNOR U17217 ( .A(n15632), .B(n17394), .Z(n17397) );
  AND U17218 ( .A(n17398), .B(n17399), .Z(n15632) );
  XNOR U17219 ( .A(n17394), .B(n15629), .Z(n17396) );
  IV U17220 ( .A(n17400), .Z(n15629) );
  AND U17221 ( .A(n17401), .B(n17402), .Z(n17400) );
  XOR U17222 ( .A(n17403), .B(n17404), .Z(n17394) );
  AND U17223 ( .A(n17405), .B(n17406), .Z(n17404) );
  XOR U17224 ( .A(n17403), .B(n15644), .Z(n17406) );
  XOR U17225 ( .A(n17407), .B(n17408), .Z(n15644) );
  AND U17226 ( .A(n799), .B(n17409), .Z(n17408) );
  XOR U17227 ( .A(n17410), .B(n17407), .Z(n17409) );
  XNOR U17228 ( .A(n15641), .B(n17403), .Z(n17405) );
  XOR U17229 ( .A(n17411), .B(n17412), .Z(n15641) );
  AND U17230 ( .A(n796), .B(n17413), .Z(n17412) );
  XOR U17231 ( .A(n17414), .B(n17411), .Z(n17413) );
  XOR U17232 ( .A(n17415), .B(n17416), .Z(n17403) );
  AND U17233 ( .A(n17417), .B(n17418), .Z(n17416) );
  XOR U17234 ( .A(n17415), .B(n15656), .Z(n17418) );
  XOR U17235 ( .A(n17419), .B(n17420), .Z(n15656) );
  AND U17236 ( .A(n799), .B(n17421), .Z(n17420) );
  XOR U17237 ( .A(n17422), .B(n17419), .Z(n17421) );
  XNOR U17238 ( .A(n15653), .B(n17415), .Z(n17417) );
  XOR U17239 ( .A(n17423), .B(n17424), .Z(n15653) );
  AND U17240 ( .A(n796), .B(n17425), .Z(n17424) );
  XOR U17241 ( .A(n17426), .B(n17423), .Z(n17425) );
  XOR U17242 ( .A(n17427), .B(n17428), .Z(n17415) );
  AND U17243 ( .A(n17429), .B(n17430), .Z(n17428) );
  XOR U17244 ( .A(n17427), .B(n15668), .Z(n17430) );
  XOR U17245 ( .A(n17431), .B(n17432), .Z(n15668) );
  AND U17246 ( .A(n799), .B(n17433), .Z(n17432) );
  XOR U17247 ( .A(n17434), .B(n17431), .Z(n17433) );
  XNOR U17248 ( .A(n15665), .B(n17427), .Z(n17429) );
  XOR U17249 ( .A(n17435), .B(n17436), .Z(n15665) );
  AND U17250 ( .A(n796), .B(n17437), .Z(n17436) );
  XOR U17251 ( .A(n17438), .B(n17435), .Z(n17437) );
  XOR U17252 ( .A(n17439), .B(n17440), .Z(n17427) );
  AND U17253 ( .A(n17441), .B(n17442), .Z(n17440) );
  XOR U17254 ( .A(n17439), .B(n15680), .Z(n17442) );
  XOR U17255 ( .A(n17443), .B(n17444), .Z(n15680) );
  AND U17256 ( .A(n799), .B(n17445), .Z(n17444) );
  XOR U17257 ( .A(n17446), .B(n17443), .Z(n17445) );
  XNOR U17258 ( .A(n15677), .B(n17439), .Z(n17441) );
  XOR U17259 ( .A(n17447), .B(n17448), .Z(n15677) );
  AND U17260 ( .A(n796), .B(n17449), .Z(n17448) );
  XOR U17261 ( .A(n17450), .B(n17447), .Z(n17449) );
  XOR U17262 ( .A(n17451), .B(n17452), .Z(n17439) );
  AND U17263 ( .A(n17453), .B(n17454), .Z(n17452) );
  XOR U17264 ( .A(n17451), .B(n15692), .Z(n17454) );
  XOR U17265 ( .A(n17455), .B(n17456), .Z(n15692) );
  AND U17266 ( .A(n799), .B(n17457), .Z(n17456) );
  XOR U17267 ( .A(n17458), .B(n17455), .Z(n17457) );
  XNOR U17268 ( .A(n15689), .B(n17451), .Z(n17453) );
  XOR U17269 ( .A(n17459), .B(n17460), .Z(n15689) );
  AND U17270 ( .A(n796), .B(n17461), .Z(n17460) );
  XOR U17271 ( .A(n17462), .B(n17459), .Z(n17461) );
  XOR U17272 ( .A(n17463), .B(n17464), .Z(n17451) );
  AND U17273 ( .A(n17465), .B(n17466), .Z(n17464) );
  XOR U17274 ( .A(n17463), .B(n15704), .Z(n17466) );
  XOR U17275 ( .A(n17467), .B(n17468), .Z(n15704) );
  AND U17276 ( .A(n799), .B(n17469), .Z(n17468) );
  XOR U17277 ( .A(n17470), .B(n17467), .Z(n17469) );
  XNOR U17278 ( .A(n15701), .B(n17463), .Z(n17465) );
  XOR U17279 ( .A(n17471), .B(n17472), .Z(n15701) );
  AND U17280 ( .A(n796), .B(n17473), .Z(n17472) );
  XOR U17281 ( .A(n17474), .B(n17471), .Z(n17473) );
  XOR U17282 ( .A(n17475), .B(n17476), .Z(n17463) );
  AND U17283 ( .A(n17477), .B(n17478), .Z(n17476) );
  XOR U17284 ( .A(n17475), .B(n15716), .Z(n17478) );
  XOR U17285 ( .A(n17479), .B(n17480), .Z(n15716) );
  AND U17286 ( .A(n799), .B(n17481), .Z(n17480) );
  XOR U17287 ( .A(n17482), .B(n17479), .Z(n17481) );
  XNOR U17288 ( .A(n15713), .B(n17475), .Z(n17477) );
  XOR U17289 ( .A(n17483), .B(n17484), .Z(n15713) );
  AND U17290 ( .A(n796), .B(n17485), .Z(n17484) );
  XOR U17291 ( .A(n17486), .B(n17483), .Z(n17485) );
  XOR U17292 ( .A(n17487), .B(n17488), .Z(n17475) );
  AND U17293 ( .A(n17489), .B(n17490), .Z(n17488) );
  XOR U17294 ( .A(n17487), .B(n15728), .Z(n17490) );
  XOR U17295 ( .A(n17491), .B(n17492), .Z(n15728) );
  AND U17296 ( .A(n799), .B(n17493), .Z(n17492) );
  XOR U17297 ( .A(n17494), .B(n17491), .Z(n17493) );
  XNOR U17298 ( .A(n15725), .B(n17487), .Z(n17489) );
  XOR U17299 ( .A(n17495), .B(n17496), .Z(n15725) );
  AND U17300 ( .A(n796), .B(n17497), .Z(n17496) );
  XOR U17301 ( .A(n17498), .B(n17495), .Z(n17497) );
  XOR U17302 ( .A(n17499), .B(n17500), .Z(n17487) );
  AND U17303 ( .A(n17501), .B(n17502), .Z(n17500) );
  XOR U17304 ( .A(n17499), .B(n15740), .Z(n17502) );
  XOR U17305 ( .A(n17503), .B(n17504), .Z(n15740) );
  AND U17306 ( .A(n799), .B(n17505), .Z(n17504) );
  XOR U17307 ( .A(n17506), .B(n17503), .Z(n17505) );
  XNOR U17308 ( .A(n15737), .B(n17499), .Z(n17501) );
  XOR U17309 ( .A(n17507), .B(n17508), .Z(n15737) );
  AND U17310 ( .A(n796), .B(n17509), .Z(n17508) );
  XOR U17311 ( .A(n17510), .B(n17507), .Z(n17509) );
  XOR U17312 ( .A(n17511), .B(n17512), .Z(n17499) );
  AND U17313 ( .A(n17513), .B(n17514), .Z(n17512) );
  XOR U17314 ( .A(n17511), .B(n15752), .Z(n17514) );
  XOR U17315 ( .A(n17515), .B(n17516), .Z(n15752) );
  AND U17316 ( .A(n799), .B(n17517), .Z(n17516) );
  XOR U17317 ( .A(n17518), .B(n17515), .Z(n17517) );
  XNOR U17318 ( .A(n15749), .B(n17511), .Z(n17513) );
  XOR U17319 ( .A(n17519), .B(n17520), .Z(n15749) );
  AND U17320 ( .A(n796), .B(n17521), .Z(n17520) );
  XOR U17321 ( .A(n17522), .B(n17519), .Z(n17521) );
  XOR U17322 ( .A(n17523), .B(n17524), .Z(n17511) );
  AND U17323 ( .A(n17525), .B(n17526), .Z(n17524) );
  XOR U17324 ( .A(n17523), .B(n15764), .Z(n17526) );
  XOR U17325 ( .A(n17527), .B(n17528), .Z(n15764) );
  AND U17326 ( .A(n799), .B(n17529), .Z(n17528) );
  XOR U17327 ( .A(n17530), .B(n17527), .Z(n17529) );
  XNOR U17328 ( .A(n15761), .B(n17523), .Z(n17525) );
  XOR U17329 ( .A(n17531), .B(n17532), .Z(n15761) );
  AND U17330 ( .A(n796), .B(n17533), .Z(n17532) );
  XOR U17331 ( .A(n17534), .B(n17531), .Z(n17533) );
  XOR U17332 ( .A(n17535), .B(n17536), .Z(n17523) );
  AND U17333 ( .A(n17537), .B(n17538), .Z(n17536) );
  XOR U17334 ( .A(n17535), .B(n15776), .Z(n17538) );
  XOR U17335 ( .A(n17539), .B(n17540), .Z(n15776) );
  AND U17336 ( .A(n799), .B(n17541), .Z(n17540) );
  XOR U17337 ( .A(n17542), .B(n17539), .Z(n17541) );
  XNOR U17338 ( .A(n15773), .B(n17535), .Z(n17537) );
  XOR U17339 ( .A(n17543), .B(n17544), .Z(n15773) );
  AND U17340 ( .A(n796), .B(n17545), .Z(n17544) );
  XOR U17341 ( .A(n17546), .B(n17543), .Z(n17545) );
  XOR U17342 ( .A(n17547), .B(n17548), .Z(n17535) );
  AND U17343 ( .A(n17549), .B(n17550), .Z(n17548) );
  XOR U17344 ( .A(n17547), .B(n15788), .Z(n17550) );
  XOR U17345 ( .A(n17551), .B(n17552), .Z(n15788) );
  AND U17346 ( .A(n799), .B(n17553), .Z(n17552) );
  XOR U17347 ( .A(n17554), .B(n17551), .Z(n17553) );
  XNOR U17348 ( .A(n15785), .B(n17547), .Z(n17549) );
  XOR U17349 ( .A(n17555), .B(n17556), .Z(n15785) );
  AND U17350 ( .A(n796), .B(n17557), .Z(n17556) );
  XOR U17351 ( .A(n17558), .B(n17555), .Z(n17557) );
  XOR U17352 ( .A(n17559), .B(n17560), .Z(n17547) );
  AND U17353 ( .A(n17561), .B(n17562), .Z(n17560) );
  XNOR U17354 ( .A(n17563), .B(n15801), .Z(n17562) );
  XOR U17355 ( .A(n17564), .B(n17565), .Z(n15801) );
  AND U17356 ( .A(n799), .B(n17566), .Z(n17565) );
  XOR U17357 ( .A(n17564), .B(n17567), .Z(n17566) );
  XNOR U17358 ( .A(n15798), .B(n17559), .Z(n17561) );
  XOR U17359 ( .A(n17568), .B(n17569), .Z(n15798) );
  AND U17360 ( .A(n796), .B(n17570), .Z(n17569) );
  XOR U17361 ( .A(n17568), .B(n17571), .Z(n17570) );
  IV U17362 ( .A(n17563), .Z(n17559) );
  AND U17363 ( .A(n17390), .B(n17393), .Z(n17563) );
  XNOR U17364 ( .A(n17572), .B(n17573), .Z(n17393) );
  AND U17365 ( .A(n799), .B(n17574), .Z(n17573) );
  XNOR U17366 ( .A(n17575), .B(n17572), .Z(n17574) );
  XOR U17367 ( .A(n17576), .B(n17577), .Z(n799) );
  AND U17368 ( .A(n17578), .B(n17579), .Z(n17577) );
  XNOR U17369 ( .A(n17398), .B(n17576), .Z(n17579) );
  AND U17370 ( .A(n17580), .B(n17581), .Z(n17398) );
  XOR U17371 ( .A(n17576), .B(n17399), .Z(n17578) );
  AND U17372 ( .A(n17582), .B(n17583), .Z(n17399) );
  XOR U17373 ( .A(n17584), .B(n17585), .Z(n17576) );
  AND U17374 ( .A(n17586), .B(n17587), .Z(n17585) );
  XOR U17375 ( .A(n17584), .B(n17410), .Z(n17587) );
  XOR U17376 ( .A(n17588), .B(n17589), .Z(n17410) );
  AND U17377 ( .A(n495), .B(n17590), .Z(n17589) );
  XOR U17378 ( .A(n17591), .B(n17588), .Z(n17590) );
  XNOR U17379 ( .A(n17407), .B(n17584), .Z(n17586) );
  XOR U17380 ( .A(n17592), .B(n17593), .Z(n17407) );
  AND U17381 ( .A(n493), .B(n17594), .Z(n17593) );
  XOR U17382 ( .A(n17595), .B(n17592), .Z(n17594) );
  XOR U17383 ( .A(n17596), .B(n17597), .Z(n17584) );
  AND U17384 ( .A(n17598), .B(n17599), .Z(n17597) );
  XOR U17385 ( .A(n17596), .B(n17422), .Z(n17599) );
  XOR U17386 ( .A(n17600), .B(n17601), .Z(n17422) );
  AND U17387 ( .A(n495), .B(n17602), .Z(n17601) );
  XOR U17388 ( .A(n17603), .B(n17600), .Z(n17602) );
  XNOR U17389 ( .A(n17419), .B(n17596), .Z(n17598) );
  XOR U17390 ( .A(n17604), .B(n17605), .Z(n17419) );
  AND U17391 ( .A(n493), .B(n17606), .Z(n17605) );
  XOR U17392 ( .A(n17607), .B(n17604), .Z(n17606) );
  XOR U17393 ( .A(n17608), .B(n17609), .Z(n17596) );
  AND U17394 ( .A(n17610), .B(n17611), .Z(n17609) );
  XOR U17395 ( .A(n17608), .B(n17434), .Z(n17611) );
  XOR U17396 ( .A(n17612), .B(n17613), .Z(n17434) );
  AND U17397 ( .A(n495), .B(n17614), .Z(n17613) );
  XOR U17398 ( .A(n17615), .B(n17612), .Z(n17614) );
  XNOR U17399 ( .A(n17431), .B(n17608), .Z(n17610) );
  XOR U17400 ( .A(n17616), .B(n17617), .Z(n17431) );
  AND U17401 ( .A(n493), .B(n17618), .Z(n17617) );
  XOR U17402 ( .A(n17619), .B(n17616), .Z(n17618) );
  XOR U17403 ( .A(n17620), .B(n17621), .Z(n17608) );
  AND U17404 ( .A(n17622), .B(n17623), .Z(n17621) );
  XOR U17405 ( .A(n17620), .B(n17446), .Z(n17623) );
  XOR U17406 ( .A(n17624), .B(n17625), .Z(n17446) );
  AND U17407 ( .A(n495), .B(n17626), .Z(n17625) );
  XOR U17408 ( .A(n17627), .B(n17624), .Z(n17626) );
  XNOR U17409 ( .A(n17443), .B(n17620), .Z(n17622) );
  XOR U17410 ( .A(n17628), .B(n17629), .Z(n17443) );
  AND U17411 ( .A(n493), .B(n17630), .Z(n17629) );
  XOR U17412 ( .A(n17631), .B(n17628), .Z(n17630) );
  XOR U17413 ( .A(n17632), .B(n17633), .Z(n17620) );
  AND U17414 ( .A(n17634), .B(n17635), .Z(n17633) );
  XOR U17415 ( .A(n17632), .B(n17458), .Z(n17635) );
  XOR U17416 ( .A(n17636), .B(n17637), .Z(n17458) );
  AND U17417 ( .A(n495), .B(n17638), .Z(n17637) );
  XOR U17418 ( .A(n17639), .B(n17636), .Z(n17638) );
  XNOR U17419 ( .A(n17455), .B(n17632), .Z(n17634) );
  XOR U17420 ( .A(n17640), .B(n17641), .Z(n17455) );
  AND U17421 ( .A(n493), .B(n17642), .Z(n17641) );
  XOR U17422 ( .A(n17643), .B(n17640), .Z(n17642) );
  XOR U17423 ( .A(n17644), .B(n17645), .Z(n17632) );
  AND U17424 ( .A(n17646), .B(n17647), .Z(n17645) );
  XOR U17425 ( .A(n17644), .B(n17470), .Z(n17647) );
  XOR U17426 ( .A(n17648), .B(n17649), .Z(n17470) );
  AND U17427 ( .A(n495), .B(n17650), .Z(n17649) );
  XOR U17428 ( .A(n17651), .B(n17648), .Z(n17650) );
  XNOR U17429 ( .A(n17467), .B(n17644), .Z(n17646) );
  XOR U17430 ( .A(n17652), .B(n17653), .Z(n17467) );
  AND U17431 ( .A(n493), .B(n17654), .Z(n17653) );
  XOR U17432 ( .A(n17655), .B(n17652), .Z(n17654) );
  XOR U17433 ( .A(n17656), .B(n17657), .Z(n17644) );
  AND U17434 ( .A(n17658), .B(n17659), .Z(n17657) );
  XOR U17435 ( .A(n17656), .B(n17482), .Z(n17659) );
  XOR U17436 ( .A(n17660), .B(n17661), .Z(n17482) );
  AND U17437 ( .A(n495), .B(n17662), .Z(n17661) );
  XOR U17438 ( .A(n17663), .B(n17660), .Z(n17662) );
  XNOR U17439 ( .A(n17479), .B(n17656), .Z(n17658) );
  XOR U17440 ( .A(n17664), .B(n17665), .Z(n17479) );
  AND U17441 ( .A(n493), .B(n17666), .Z(n17665) );
  XOR U17442 ( .A(n17667), .B(n17664), .Z(n17666) );
  XOR U17443 ( .A(n17668), .B(n17669), .Z(n17656) );
  AND U17444 ( .A(n17670), .B(n17671), .Z(n17669) );
  XOR U17445 ( .A(n17668), .B(n17494), .Z(n17671) );
  XOR U17446 ( .A(n17672), .B(n17673), .Z(n17494) );
  AND U17447 ( .A(n495), .B(n17674), .Z(n17673) );
  XOR U17448 ( .A(n17675), .B(n17672), .Z(n17674) );
  XNOR U17449 ( .A(n17491), .B(n17668), .Z(n17670) );
  XOR U17450 ( .A(n17676), .B(n17677), .Z(n17491) );
  AND U17451 ( .A(n493), .B(n17678), .Z(n17677) );
  XOR U17452 ( .A(n17679), .B(n17676), .Z(n17678) );
  XOR U17453 ( .A(n17680), .B(n17681), .Z(n17668) );
  AND U17454 ( .A(n17682), .B(n17683), .Z(n17681) );
  XOR U17455 ( .A(n17680), .B(n17506), .Z(n17683) );
  XOR U17456 ( .A(n17684), .B(n17685), .Z(n17506) );
  AND U17457 ( .A(n495), .B(n17686), .Z(n17685) );
  XOR U17458 ( .A(n17687), .B(n17684), .Z(n17686) );
  XNOR U17459 ( .A(n17503), .B(n17680), .Z(n17682) );
  XOR U17460 ( .A(n17688), .B(n17689), .Z(n17503) );
  AND U17461 ( .A(n493), .B(n17690), .Z(n17689) );
  XOR U17462 ( .A(n17691), .B(n17688), .Z(n17690) );
  XOR U17463 ( .A(n17692), .B(n17693), .Z(n17680) );
  AND U17464 ( .A(n17694), .B(n17695), .Z(n17693) );
  XOR U17465 ( .A(n17692), .B(n17518), .Z(n17695) );
  XOR U17466 ( .A(n17696), .B(n17697), .Z(n17518) );
  AND U17467 ( .A(n495), .B(n17698), .Z(n17697) );
  XOR U17468 ( .A(n17699), .B(n17696), .Z(n17698) );
  XNOR U17469 ( .A(n17515), .B(n17692), .Z(n17694) );
  XOR U17470 ( .A(n17700), .B(n17701), .Z(n17515) );
  AND U17471 ( .A(n493), .B(n17702), .Z(n17701) );
  XOR U17472 ( .A(n17703), .B(n17700), .Z(n17702) );
  XOR U17473 ( .A(n17704), .B(n17705), .Z(n17692) );
  AND U17474 ( .A(n17706), .B(n17707), .Z(n17705) );
  XOR U17475 ( .A(n17704), .B(n17530), .Z(n17707) );
  XOR U17476 ( .A(n17708), .B(n17709), .Z(n17530) );
  AND U17477 ( .A(n495), .B(n17710), .Z(n17709) );
  XOR U17478 ( .A(n17711), .B(n17708), .Z(n17710) );
  XNOR U17479 ( .A(n17527), .B(n17704), .Z(n17706) );
  XOR U17480 ( .A(n17712), .B(n17713), .Z(n17527) );
  AND U17481 ( .A(n493), .B(n17714), .Z(n17713) );
  XOR U17482 ( .A(n17715), .B(n17712), .Z(n17714) );
  XOR U17483 ( .A(n17716), .B(n17717), .Z(n17704) );
  AND U17484 ( .A(n17718), .B(n17719), .Z(n17717) );
  XOR U17485 ( .A(n17716), .B(n17542), .Z(n17719) );
  XOR U17486 ( .A(n17720), .B(n17721), .Z(n17542) );
  AND U17487 ( .A(n495), .B(n17722), .Z(n17721) );
  XOR U17488 ( .A(n17723), .B(n17720), .Z(n17722) );
  XNOR U17489 ( .A(n17539), .B(n17716), .Z(n17718) );
  XOR U17490 ( .A(n17724), .B(n17725), .Z(n17539) );
  AND U17491 ( .A(n493), .B(n17726), .Z(n17725) );
  XOR U17492 ( .A(n17727), .B(n17724), .Z(n17726) );
  XOR U17493 ( .A(n17728), .B(n17729), .Z(n17716) );
  AND U17494 ( .A(n17730), .B(n17731), .Z(n17729) );
  XOR U17495 ( .A(n17728), .B(n17554), .Z(n17731) );
  XOR U17496 ( .A(n17732), .B(n17733), .Z(n17554) );
  AND U17497 ( .A(n495), .B(n17734), .Z(n17733) );
  XOR U17498 ( .A(n17735), .B(n17732), .Z(n17734) );
  XNOR U17499 ( .A(n17551), .B(n17728), .Z(n17730) );
  XOR U17500 ( .A(n17736), .B(n17737), .Z(n17551) );
  AND U17501 ( .A(n493), .B(n17738), .Z(n17737) );
  XOR U17502 ( .A(n17739), .B(n17736), .Z(n17738) );
  XOR U17503 ( .A(n17740), .B(n17741), .Z(n17728) );
  AND U17504 ( .A(n17742), .B(n17743), .Z(n17741) );
  XNOR U17505 ( .A(n17744), .B(n17567), .Z(n17743) );
  XOR U17506 ( .A(n17745), .B(n17746), .Z(n17567) );
  AND U17507 ( .A(n495), .B(n17747), .Z(n17746) );
  XOR U17508 ( .A(n17745), .B(n17748), .Z(n17747) );
  XNOR U17509 ( .A(n17564), .B(n17740), .Z(n17742) );
  XOR U17510 ( .A(n17749), .B(n17750), .Z(n17564) );
  AND U17511 ( .A(n493), .B(n17751), .Z(n17750) );
  XOR U17512 ( .A(n17749), .B(n17752), .Z(n17751) );
  IV U17513 ( .A(n17744), .Z(n17740) );
  AND U17514 ( .A(n17572), .B(n17575), .Z(n17744) );
  XNOR U17515 ( .A(n17753), .B(n17754), .Z(n17575) );
  AND U17516 ( .A(n495), .B(n17755), .Z(n17754) );
  XNOR U17517 ( .A(n17756), .B(n17753), .Z(n17755) );
  XOR U17518 ( .A(n17757), .B(n17758), .Z(n495) );
  AND U17519 ( .A(n17759), .B(n17760), .Z(n17758) );
  XNOR U17520 ( .A(n17580), .B(n17757), .Z(n17760) );
  AND U17521 ( .A(p_input[1791]), .B(p_input[1775]), .Z(n17580) );
  XOR U17522 ( .A(n17757), .B(n17581), .Z(n17759) );
  AND U17523 ( .A(p_input[1759]), .B(p_input[1743]), .Z(n17581) );
  XOR U17524 ( .A(n17761), .B(n17762), .Z(n17757) );
  AND U17525 ( .A(n17763), .B(n17764), .Z(n17762) );
  XOR U17526 ( .A(n17761), .B(n17591), .Z(n17764) );
  XNOR U17527 ( .A(p_input[1774]), .B(n17765), .Z(n17591) );
  AND U17528 ( .A(n639), .B(n17766), .Z(n17765) );
  XOR U17529 ( .A(p_input[1790]), .B(p_input[1774]), .Z(n17766) );
  XNOR U17530 ( .A(n17588), .B(n17761), .Z(n17763) );
  XOR U17531 ( .A(n17767), .B(n17768), .Z(n17588) );
  AND U17532 ( .A(n637), .B(n17769), .Z(n17768) );
  XOR U17533 ( .A(p_input[1758]), .B(p_input[1742]), .Z(n17769) );
  XOR U17534 ( .A(n17770), .B(n17771), .Z(n17761) );
  AND U17535 ( .A(n17772), .B(n17773), .Z(n17771) );
  XOR U17536 ( .A(n17770), .B(n17603), .Z(n17773) );
  XNOR U17537 ( .A(p_input[1773]), .B(n17774), .Z(n17603) );
  AND U17538 ( .A(n639), .B(n17775), .Z(n17774) );
  XOR U17539 ( .A(p_input[1789]), .B(p_input[1773]), .Z(n17775) );
  XNOR U17540 ( .A(n17600), .B(n17770), .Z(n17772) );
  XOR U17541 ( .A(n17776), .B(n17777), .Z(n17600) );
  AND U17542 ( .A(n637), .B(n17778), .Z(n17777) );
  XOR U17543 ( .A(p_input[1757]), .B(p_input[1741]), .Z(n17778) );
  XOR U17544 ( .A(n17779), .B(n17780), .Z(n17770) );
  AND U17545 ( .A(n17781), .B(n17782), .Z(n17780) );
  XOR U17546 ( .A(n17779), .B(n17615), .Z(n17782) );
  XNOR U17547 ( .A(p_input[1772]), .B(n17783), .Z(n17615) );
  AND U17548 ( .A(n639), .B(n17784), .Z(n17783) );
  XOR U17549 ( .A(p_input[1788]), .B(p_input[1772]), .Z(n17784) );
  XNOR U17550 ( .A(n17612), .B(n17779), .Z(n17781) );
  XOR U17551 ( .A(n17785), .B(n17786), .Z(n17612) );
  AND U17552 ( .A(n637), .B(n17787), .Z(n17786) );
  XOR U17553 ( .A(p_input[1756]), .B(p_input[1740]), .Z(n17787) );
  XOR U17554 ( .A(n17788), .B(n17789), .Z(n17779) );
  AND U17555 ( .A(n17790), .B(n17791), .Z(n17789) );
  XOR U17556 ( .A(n17788), .B(n17627), .Z(n17791) );
  XNOR U17557 ( .A(p_input[1771]), .B(n17792), .Z(n17627) );
  AND U17558 ( .A(n639), .B(n17793), .Z(n17792) );
  XOR U17559 ( .A(p_input[1787]), .B(p_input[1771]), .Z(n17793) );
  XNOR U17560 ( .A(n17624), .B(n17788), .Z(n17790) );
  XOR U17561 ( .A(n17794), .B(n17795), .Z(n17624) );
  AND U17562 ( .A(n637), .B(n17796), .Z(n17795) );
  XOR U17563 ( .A(p_input[1755]), .B(p_input[1739]), .Z(n17796) );
  XOR U17564 ( .A(n17797), .B(n17798), .Z(n17788) );
  AND U17565 ( .A(n17799), .B(n17800), .Z(n17798) );
  XOR U17566 ( .A(n17797), .B(n17639), .Z(n17800) );
  XNOR U17567 ( .A(p_input[1770]), .B(n17801), .Z(n17639) );
  AND U17568 ( .A(n639), .B(n17802), .Z(n17801) );
  XOR U17569 ( .A(p_input[1786]), .B(p_input[1770]), .Z(n17802) );
  XNOR U17570 ( .A(n17636), .B(n17797), .Z(n17799) );
  XOR U17571 ( .A(n17803), .B(n17804), .Z(n17636) );
  AND U17572 ( .A(n637), .B(n17805), .Z(n17804) );
  XOR U17573 ( .A(p_input[1754]), .B(p_input[1738]), .Z(n17805) );
  XOR U17574 ( .A(n17806), .B(n17807), .Z(n17797) );
  AND U17575 ( .A(n17808), .B(n17809), .Z(n17807) );
  XOR U17576 ( .A(n17806), .B(n17651), .Z(n17809) );
  XNOR U17577 ( .A(p_input[1769]), .B(n17810), .Z(n17651) );
  AND U17578 ( .A(n639), .B(n17811), .Z(n17810) );
  XOR U17579 ( .A(p_input[1785]), .B(p_input[1769]), .Z(n17811) );
  XNOR U17580 ( .A(n17648), .B(n17806), .Z(n17808) );
  XOR U17581 ( .A(n17812), .B(n17813), .Z(n17648) );
  AND U17582 ( .A(n637), .B(n17814), .Z(n17813) );
  XOR U17583 ( .A(p_input[1753]), .B(p_input[1737]), .Z(n17814) );
  XOR U17584 ( .A(n17815), .B(n17816), .Z(n17806) );
  AND U17585 ( .A(n17817), .B(n17818), .Z(n17816) );
  XOR U17586 ( .A(n17815), .B(n17663), .Z(n17818) );
  XNOR U17587 ( .A(p_input[1768]), .B(n17819), .Z(n17663) );
  AND U17588 ( .A(n639), .B(n17820), .Z(n17819) );
  XOR U17589 ( .A(p_input[1784]), .B(p_input[1768]), .Z(n17820) );
  XNOR U17590 ( .A(n17660), .B(n17815), .Z(n17817) );
  XOR U17591 ( .A(n17821), .B(n17822), .Z(n17660) );
  AND U17592 ( .A(n637), .B(n17823), .Z(n17822) );
  XOR U17593 ( .A(p_input[1752]), .B(p_input[1736]), .Z(n17823) );
  XOR U17594 ( .A(n17824), .B(n17825), .Z(n17815) );
  AND U17595 ( .A(n17826), .B(n17827), .Z(n17825) );
  XOR U17596 ( .A(n17824), .B(n17675), .Z(n17827) );
  XNOR U17597 ( .A(p_input[1767]), .B(n17828), .Z(n17675) );
  AND U17598 ( .A(n639), .B(n17829), .Z(n17828) );
  XOR U17599 ( .A(p_input[1783]), .B(p_input[1767]), .Z(n17829) );
  XNOR U17600 ( .A(n17672), .B(n17824), .Z(n17826) );
  XOR U17601 ( .A(n17830), .B(n17831), .Z(n17672) );
  AND U17602 ( .A(n637), .B(n17832), .Z(n17831) );
  XOR U17603 ( .A(p_input[1751]), .B(p_input[1735]), .Z(n17832) );
  XOR U17604 ( .A(n17833), .B(n17834), .Z(n17824) );
  AND U17605 ( .A(n17835), .B(n17836), .Z(n17834) );
  XOR U17606 ( .A(n17833), .B(n17687), .Z(n17836) );
  XNOR U17607 ( .A(p_input[1766]), .B(n17837), .Z(n17687) );
  AND U17608 ( .A(n639), .B(n17838), .Z(n17837) );
  XOR U17609 ( .A(p_input[1782]), .B(p_input[1766]), .Z(n17838) );
  XNOR U17610 ( .A(n17684), .B(n17833), .Z(n17835) );
  XOR U17611 ( .A(n17839), .B(n17840), .Z(n17684) );
  AND U17612 ( .A(n637), .B(n17841), .Z(n17840) );
  XOR U17613 ( .A(p_input[1750]), .B(p_input[1734]), .Z(n17841) );
  XOR U17614 ( .A(n17842), .B(n17843), .Z(n17833) );
  AND U17615 ( .A(n17844), .B(n17845), .Z(n17843) );
  XOR U17616 ( .A(n17842), .B(n17699), .Z(n17845) );
  XNOR U17617 ( .A(p_input[1765]), .B(n17846), .Z(n17699) );
  AND U17618 ( .A(n639), .B(n17847), .Z(n17846) );
  XOR U17619 ( .A(p_input[1781]), .B(p_input[1765]), .Z(n17847) );
  XNOR U17620 ( .A(n17696), .B(n17842), .Z(n17844) );
  XOR U17621 ( .A(n17848), .B(n17849), .Z(n17696) );
  AND U17622 ( .A(n637), .B(n17850), .Z(n17849) );
  XOR U17623 ( .A(p_input[1749]), .B(p_input[1733]), .Z(n17850) );
  XOR U17624 ( .A(n17851), .B(n17852), .Z(n17842) );
  AND U17625 ( .A(n17853), .B(n17854), .Z(n17852) );
  XOR U17626 ( .A(n17851), .B(n17711), .Z(n17854) );
  XNOR U17627 ( .A(p_input[1764]), .B(n17855), .Z(n17711) );
  AND U17628 ( .A(n639), .B(n17856), .Z(n17855) );
  XOR U17629 ( .A(p_input[1780]), .B(p_input[1764]), .Z(n17856) );
  XNOR U17630 ( .A(n17708), .B(n17851), .Z(n17853) );
  XOR U17631 ( .A(n17857), .B(n17858), .Z(n17708) );
  AND U17632 ( .A(n637), .B(n17859), .Z(n17858) );
  XOR U17633 ( .A(p_input[1748]), .B(p_input[1732]), .Z(n17859) );
  XOR U17634 ( .A(n17860), .B(n17861), .Z(n17851) );
  AND U17635 ( .A(n17862), .B(n17863), .Z(n17861) );
  XOR U17636 ( .A(n17860), .B(n17723), .Z(n17863) );
  XNOR U17637 ( .A(p_input[1763]), .B(n17864), .Z(n17723) );
  AND U17638 ( .A(n639), .B(n17865), .Z(n17864) );
  XOR U17639 ( .A(p_input[1779]), .B(p_input[1763]), .Z(n17865) );
  XNOR U17640 ( .A(n17720), .B(n17860), .Z(n17862) );
  XOR U17641 ( .A(n17866), .B(n17867), .Z(n17720) );
  AND U17642 ( .A(n637), .B(n17868), .Z(n17867) );
  XOR U17643 ( .A(p_input[1747]), .B(p_input[1731]), .Z(n17868) );
  XOR U17644 ( .A(n17869), .B(n17870), .Z(n17860) );
  AND U17645 ( .A(n17871), .B(n17872), .Z(n17870) );
  XOR U17646 ( .A(n17869), .B(n17735), .Z(n17872) );
  XNOR U17647 ( .A(p_input[1762]), .B(n17873), .Z(n17735) );
  AND U17648 ( .A(n639), .B(n17874), .Z(n17873) );
  XOR U17649 ( .A(p_input[1778]), .B(p_input[1762]), .Z(n17874) );
  XNOR U17650 ( .A(n17732), .B(n17869), .Z(n17871) );
  XOR U17651 ( .A(n17875), .B(n17876), .Z(n17732) );
  AND U17652 ( .A(n637), .B(n17877), .Z(n17876) );
  XOR U17653 ( .A(p_input[1746]), .B(p_input[1730]), .Z(n17877) );
  XOR U17654 ( .A(n17878), .B(n17879), .Z(n17869) );
  AND U17655 ( .A(n17880), .B(n17881), .Z(n17879) );
  XNOR U17656 ( .A(n17882), .B(n17748), .Z(n17881) );
  XNOR U17657 ( .A(p_input[1761]), .B(n17883), .Z(n17748) );
  AND U17658 ( .A(n639), .B(n17884), .Z(n17883) );
  XNOR U17659 ( .A(p_input[1777]), .B(n17885), .Z(n17884) );
  IV U17660 ( .A(p_input[1761]), .Z(n17885) );
  XNOR U17661 ( .A(n17745), .B(n17878), .Z(n17880) );
  XNOR U17662 ( .A(p_input[1729]), .B(n17886), .Z(n17745) );
  AND U17663 ( .A(n637), .B(n17887), .Z(n17886) );
  XOR U17664 ( .A(p_input[1745]), .B(p_input[1729]), .Z(n17887) );
  IV U17665 ( .A(n17882), .Z(n17878) );
  AND U17666 ( .A(n17753), .B(n17756), .Z(n17882) );
  XOR U17667 ( .A(p_input[1760]), .B(n17888), .Z(n17756) );
  AND U17668 ( .A(n639), .B(n17889), .Z(n17888) );
  XOR U17669 ( .A(p_input[1776]), .B(p_input[1760]), .Z(n17889) );
  XOR U17670 ( .A(n17890), .B(n17891), .Z(n639) );
  AND U17671 ( .A(n17892), .B(n17893), .Z(n17891) );
  XNOR U17672 ( .A(p_input[1791]), .B(n17890), .Z(n17893) );
  XOR U17673 ( .A(n17890), .B(p_input[1775]), .Z(n17892) );
  XOR U17674 ( .A(n17894), .B(n17895), .Z(n17890) );
  AND U17675 ( .A(n17896), .B(n17897), .Z(n17895) );
  XNOR U17676 ( .A(p_input[1790]), .B(n17894), .Z(n17897) );
  XOR U17677 ( .A(n17894), .B(p_input[1774]), .Z(n17896) );
  XOR U17678 ( .A(n17898), .B(n17899), .Z(n17894) );
  AND U17679 ( .A(n17900), .B(n17901), .Z(n17899) );
  XNOR U17680 ( .A(p_input[1789]), .B(n17898), .Z(n17901) );
  XOR U17681 ( .A(n17898), .B(p_input[1773]), .Z(n17900) );
  XOR U17682 ( .A(n17902), .B(n17903), .Z(n17898) );
  AND U17683 ( .A(n17904), .B(n17905), .Z(n17903) );
  XNOR U17684 ( .A(p_input[1788]), .B(n17902), .Z(n17905) );
  XOR U17685 ( .A(n17902), .B(p_input[1772]), .Z(n17904) );
  XOR U17686 ( .A(n17906), .B(n17907), .Z(n17902) );
  AND U17687 ( .A(n17908), .B(n17909), .Z(n17907) );
  XNOR U17688 ( .A(p_input[1787]), .B(n17906), .Z(n17909) );
  XOR U17689 ( .A(n17906), .B(p_input[1771]), .Z(n17908) );
  XOR U17690 ( .A(n17910), .B(n17911), .Z(n17906) );
  AND U17691 ( .A(n17912), .B(n17913), .Z(n17911) );
  XNOR U17692 ( .A(p_input[1786]), .B(n17910), .Z(n17913) );
  XOR U17693 ( .A(n17910), .B(p_input[1770]), .Z(n17912) );
  XOR U17694 ( .A(n17914), .B(n17915), .Z(n17910) );
  AND U17695 ( .A(n17916), .B(n17917), .Z(n17915) );
  XNOR U17696 ( .A(p_input[1785]), .B(n17914), .Z(n17917) );
  XOR U17697 ( .A(n17914), .B(p_input[1769]), .Z(n17916) );
  XOR U17698 ( .A(n17918), .B(n17919), .Z(n17914) );
  AND U17699 ( .A(n17920), .B(n17921), .Z(n17919) );
  XNOR U17700 ( .A(p_input[1784]), .B(n17918), .Z(n17921) );
  XOR U17701 ( .A(n17918), .B(p_input[1768]), .Z(n17920) );
  XOR U17702 ( .A(n17922), .B(n17923), .Z(n17918) );
  AND U17703 ( .A(n17924), .B(n17925), .Z(n17923) );
  XNOR U17704 ( .A(p_input[1783]), .B(n17922), .Z(n17925) );
  XOR U17705 ( .A(n17922), .B(p_input[1767]), .Z(n17924) );
  XOR U17706 ( .A(n17926), .B(n17927), .Z(n17922) );
  AND U17707 ( .A(n17928), .B(n17929), .Z(n17927) );
  XNOR U17708 ( .A(p_input[1782]), .B(n17926), .Z(n17929) );
  XOR U17709 ( .A(n17926), .B(p_input[1766]), .Z(n17928) );
  XOR U17710 ( .A(n17930), .B(n17931), .Z(n17926) );
  AND U17711 ( .A(n17932), .B(n17933), .Z(n17931) );
  XNOR U17712 ( .A(p_input[1781]), .B(n17930), .Z(n17933) );
  XOR U17713 ( .A(n17930), .B(p_input[1765]), .Z(n17932) );
  XOR U17714 ( .A(n17934), .B(n17935), .Z(n17930) );
  AND U17715 ( .A(n17936), .B(n17937), .Z(n17935) );
  XNOR U17716 ( .A(p_input[1780]), .B(n17934), .Z(n17937) );
  XOR U17717 ( .A(n17934), .B(p_input[1764]), .Z(n17936) );
  XOR U17718 ( .A(n17938), .B(n17939), .Z(n17934) );
  AND U17719 ( .A(n17940), .B(n17941), .Z(n17939) );
  XNOR U17720 ( .A(p_input[1779]), .B(n17938), .Z(n17941) );
  XOR U17721 ( .A(n17938), .B(p_input[1763]), .Z(n17940) );
  XOR U17722 ( .A(n17942), .B(n17943), .Z(n17938) );
  AND U17723 ( .A(n17944), .B(n17945), .Z(n17943) );
  XNOR U17724 ( .A(p_input[1778]), .B(n17942), .Z(n17945) );
  XOR U17725 ( .A(n17942), .B(p_input[1762]), .Z(n17944) );
  XNOR U17726 ( .A(n17946), .B(n17947), .Z(n17942) );
  AND U17727 ( .A(n17948), .B(n17949), .Z(n17947) );
  XOR U17728 ( .A(p_input[1777]), .B(n17946), .Z(n17949) );
  XNOR U17729 ( .A(p_input[1761]), .B(n17946), .Z(n17948) );
  AND U17730 ( .A(p_input[1776]), .B(n17950), .Z(n17946) );
  IV U17731 ( .A(p_input[1760]), .Z(n17950) );
  XNOR U17732 ( .A(p_input[1728]), .B(n17951), .Z(n17753) );
  AND U17733 ( .A(n637), .B(n17952), .Z(n17951) );
  XOR U17734 ( .A(p_input[1744]), .B(p_input[1728]), .Z(n17952) );
  XOR U17735 ( .A(n17953), .B(n17954), .Z(n637) );
  AND U17736 ( .A(n17955), .B(n17956), .Z(n17954) );
  XNOR U17737 ( .A(p_input[1759]), .B(n17953), .Z(n17956) );
  XOR U17738 ( .A(n17953), .B(p_input[1743]), .Z(n17955) );
  XOR U17739 ( .A(n17957), .B(n17958), .Z(n17953) );
  AND U17740 ( .A(n17959), .B(n17960), .Z(n17958) );
  XNOR U17741 ( .A(p_input[1758]), .B(n17957), .Z(n17960) );
  XNOR U17742 ( .A(n17957), .B(n17767), .Z(n17959) );
  IV U17743 ( .A(p_input[1742]), .Z(n17767) );
  XOR U17744 ( .A(n17961), .B(n17962), .Z(n17957) );
  AND U17745 ( .A(n17963), .B(n17964), .Z(n17962) );
  XNOR U17746 ( .A(p_input[1757]), .B(n17961), .Z(n17964) );
  XNOR U17747 ( .A(n17961), .B(n17776), .Z(n17963) );
  IV U17748 ( .A(p_input[1741]), .Z(n17776) );
  XOR U17749 ( .A(n17965), .B(n17966), .Z(n17961) );
  AND U17750 ( .A(n17967), .B(n17968), .Z(n17966) );
  XNOR U17751 ( .A(p_input[1756]), .B(n17965), .Z(n17968) );
  XNOR U17752 ( .A(n17965), .B(n17785), .Z(n17967) );
  IV U17753 ( .A(p_input[1740]), .Z(n17785) );
  XOR U17754 ( .A(n17969), .B(n17970), .Z(n17965) );
  AND U17755 ( .A(n17971), .B(n17972), .Z(n17970) );
  XNOR U17756 ( .A(p_input[1755]), .B(n17969), .Z(n17972) );
  XNOR U17757 ( .A(n17969), .B(n17794), .Z(n17971) );
  IV U17758 ( .A(p_input[1739]), .Z(n17794) );
  XOR U17759 ( .A(n17973), .B(n17974), .Z(n17969) );
  AND U17760 ( .A(n17975), .B(n17976), .Z(n17974) );
  XNOR U17761 ( .A(p_input[1754]), .B(n17973), .Z(n17976) );
  XNOR U17762 ( .A(n17973), .B(n17803), .Z(n17975) );
  IV U17763 ( .A(p_input[1738]), .Z(n17803) );
  XOR U17764 ( .A(n17977), .B(n17978), .Z(n17973) );
  AND U17765 ( .A(n17979), .B(n17980), .Z(n17978) );
  XNOR U17766 ( .A(p_input[1753]), .B(n17977), .Z(n17980) );
  XNOR U17767 ( .A(n17977), .B(n17812), .Z(n17979) );
  IV U17768 ( .A(p_input[1737]), .Z(n17812) );
  XOR U17769 ( .A(n17981), .B(n17982), .Z(n17977) );
  AND U17770 ( .A(n17983), .B(n17984), .Z(n17982) );
  XNOR U17771 ( .A(p_input[1752]), .B(n17981), .Z(n17984) );
  XNOR U17772 ( .A(n17981), .B(n17821), .Z(n17983) );
  IV U17773 ( .A(p_input[1736]), .Z(n17821) );
  XOR U17774 ( .A(n17985), .B(n17986), .Z(n17981) );
  AND U17775 ( .A(n17987), .B(n17988), .Z(n17986) );
  XNOR U17776 ( .A(p_input[1751]), .B(n17985), .Z(n17988) );
  XNOR U17777 ( .A(n17985), .B(n17830), .Z(n17987) );
  IV U17778 ( .A(p_input[1735]), .Z(n17830) );
  XOR U17779 ( .A(n17989), .B(n17990), .Z(n17985) );
  AND U17780 ( .A(n17991), .B(n17992), .Z(n17990) );
  XNOR U17781 ( .A(p_input[1750]), .B(n17989), .Z(n17992) );
  XNOR U17782 ( .A(n17989), .B(n17839), .Z(n17991) );
  IV U17783 ( .A(p_input[1734]), .Z(n17839) );
  XOR U17784 ( .A(n17993), .B(n17994), .Z(n17989) );
  AND U17785 ( .A(n17995), .B(n17996), .Z(n17994) );
  XNOR U17786 ( .A(p_input[1749]), .B(n17993), .Z(n17996) );
  XNOR U17787 ( .A(n17993), .B(n17848), .Z(n17995) );
  IV U17788 ( .A(p_input[1733]), .Z(n17848) );
  XOR U17789 ( .A(n17997), .B(n17998), .Z(n17993) );
  AND U17790 ( .A(n17999), .B(n18000), .Z(n17998) );
  XNOR U17791 ( .A(p_input[1748]), .B(n17997), .Z(n18000) );
  XNOR U17792 ( .A(n17997), .B(n17857), .Z(n17999) );
  IV U17793 ( .A(p_input[1732]), .Z(n17857) );
  XOR U17794 ( .A(n18001), .B(n18002), .Z(n17997) );
  AND U17795 ( .A(n18003), .B(n18004), .Z(n18002) );
  XNOR U17796 ( .A(p_input[1747]), .B(n18001), .Z(n18004) );
  XNOR U17797 ( .A(n18001), .B(n17866), .Z(n18003) );
  IV U17798 ( .A(p_input[1731]), .Z(n17866) );
  XOR U17799 ( .A(n18005), .B(n18006), .Z(n18001) );
  AND U17800 ( .A(n18007), .B(n18008), .Z(n18006) );
  XNOR U17801 ( .A(p_input[1746]), .B(n18005), .Z(n18008) );
  XNOR U17802 ( .A(n18005), .B(n17875), .Z(n18007) );
  IV U17803 ( .A(p_input[1730]), .Z(n17875) );
  XNOR U17804 ( .A(n18009), .B(n18010), .Z(n18005) );
  AND U17805 ( .A(n18011), .B(n18012), .Z(n18010) );
  XOR U17806 ( .A(p_input[1745]), .B(n18009), .Z(n18012) );
  XNOR U17807 ( .A(p_input[1729]), .B(n18009), .Z(n18011) );
  AND U17808 ( .A(p_input[1744]), .B(n18013), .Z(n18009) );
  IV U17809 ( .A(p_input[1728]), .Z(n18013) );
  XOR U17810 ( .A(n18014), .B(n18015), .Z(n17572) );
  AND U17811 ( .A(n493), .B(n18016), .Z(n18015) );
  XNOR U17812 ( .A(n18017), .B(n18014), .Z(n18016) );
  XOR U17813 ( .A(n18018), .B(n18019), .Z(n493) );
  AND U17814 ( .A(n18020), .B(n18021), .Z(n18019) );
  XNOR U17815 ( .A(n17582), .B(n18018), .Z(n18021) );
  AND U17816 ( .A(p_input[1727]), .B(p_input[1711]), .Z(n17582) );
  XOR U17817 ( .A(n18018), .B(n17583), .Z(n18020) );
  AND U17818 ( .A(p_input[1695]), .B(p_input[1679]), .Z(n17583) );
  XOR U17819 ( .A(n18022), .B(n18023), .Z(n18018) );
  AND U17820 ( .A(n18024), .B(n18025), .Z(n18023) );
  XOR U17821 ( .A(n18022), .B(n17595), .Z(n18025) );
  XNOR U17822 ( .A(p_input[1710]), .B(n18026), .Z(n17595) );
  AND U17823 ( .A(n643), .B(n18027), .Z(n18026) );
  XOR U17824 ( .A(p_input[1726]), .B(p_input[1710]), .Z(n18027) );
  XNOR U17825 ( .A(n17592), .B(n18022), .Z(n18024) );
  XOR U17826 ( .A(n18028), .B(n18029), .Z(n17592) );
  AND U17827 ( .A(n640), .B(n18030), .Z(n18029) );
  XOR U17828 ( .A(p_input[1694]), .B(p_input[1678]), .Z(n18030) );
  XOR U17829 ( .A(n18031), .B(n18032), .Z(n18022) );
  AND U17830 ( .A(n18033), .B(n18034), .Z(n18032) );
  XOR U17831 ( .A(n18031), .B(n17607), .Z(n18034) );
  XNOR U17832 ( .A(p_input[1709]), .B(n18035), .Z(n17607) );
  AND U17833 ( .A(n643), .B(n18036), .Z(n18035) );
  XOR U17834 ( .A(p_input[1725]), .B(p_input[1709]), .Z(n18036) );
  XNOR U17835 ( .A(n17604), .B(n18031), .Z(n18033) );
  XOR U17836 ( .A(n18037), .B(n18038), .Z(n17604) );
  AND U17837 ( .A(n640), .B(n18039), .Z(n18038) );
  XOR U17838 ( .A(p_input[1693]), .B(p_input[1677]), .Z(n18039) );
  XOR U17839 ( .A(n18040), .B(n18041), .Z(n18031) );
  AND U17840 ( .A(n18042), .B(n18043), .Z(n18041) );
  XOR U17841 ( .A(n18040), .B(n17619), .Z(n18043) );
  XNOR U17842 ( .A(p_input[1708]), .B(n18044), .Z(n17619) );
  AND U17843 ( .A(n643), .B(n18045), .Z(n18044) );
  XOR U17844 ( .A(p_input[1724]), .B(p_input[1708]), .Z(n18045) );
  XNOR U17845 ( .A(n17616), .B(n18040), .Z(n18042) );
  XOR U17846 ( .A(n18046), .B(n18047), .Z(n17616) );
  AND U17847 ( .A(n640), .B(n18048), .Z(n18047) );
  XOR U17848 ( .A(p_input[1692]), .B(p_input[1676]), .Z(n18048) );
  XOR U17849 ( .A(n18049), .B(n18050), .Z(n18040) );
  AND U17850 ( .A(n18051), .B(n18052), .Z(n18050) );
  XOR U17851 ( .A(n18049), .B(n17631), .Z(n18052) );
  XNOR U17852 ( .A(p_input[1707]), .B(n18053), .Z(n17631) );
  AND U17853 ( .A(n643), .B(n18054), .Z(n18053) );
  XOR U17854 ( .A(p_input[1723]), .B(p_input[1707]), .Z(n18054) );
  XNOR U17855 ( .A(n17628), .B(n18049), .Z(n18051) );
  XOR U17856 ( .A(n18055), .B(n18056), .Z(n17628) );
  AND U17857 ( .A(n640), .B(n18057), .Z(n18056) );
  XOR U17858 ( .A(p_input[1691]), .B(p_input[1675]), .Z(n18057) );
  XOR U17859 ( .A(n18058), .B(n18059), .Z(n18049) );
  AND U17860 ( .A(n18060), .B(n18061), .Z(n18059) );
  XOR U17861 ( .A(n18058), .B(n17643), .Z(n18061) );
  XNOR U17862 ( .A(p_input[1706]), .B(n18062), .Z(n17643) );
  AND U17863 ( .A(n643), .B(n18063), .Z(n18062) );
  XOR U17864 ( .A(p_input[1722]), .B(p_input[1706]), .Z(n18063) );
  XNOR U17865 ( .A(n17640), .B(n18058), .Z(n18060) );
  XOR U17866 ( .A(n18064), .B(n18065), .Z(n17640) );
  AND U17867 ( .A(n640), .B(n18066), .Z(n18065) );
  XOR U17868 ( .A(p_input[1690]), .B(p_input[1674]), .Z(n18066) );
  XOR U17869 ( .A(n18067), .B(n18068), .Z(n18058) );
  AND U17870 ( .A(n18069), .B(n18070), .Z(n18068) );
  XOR U17871 ( .A(n18067), .B(n17655), .Z(n18070) );
  XNOR U17872 ( .A(p_input[1705]), .B(n18071), .Z(n17655) );
  AND U17873 ( .A(n643), .B(n18072), .Z(n18071) );
  XOR U17874 ( .A(p_input[1721]), .B(p_input[1705]), .Z(n18072) );
  XNOR U17875 ( .A(n17652), .B(n18067), .Z(n18069) );
  XOR U17876 ( .A(n18073), .B(n18074), .Z(n17652) );
  AND U17877 ( .A(n640), .B(n18075), .Z(n18074) );
  XOR U17878 ( .A(p_input[1689]), .B(p_input[1673]), .Z(n18075) );
  XOR U17879 ( .A(n18076), .B(n18077), .Z(n18067) );
  AND U17880 ( .A(n18078), .B(n18079), .Z(n18077) );
  XOR U17881 ( .A(n18076), .B(n17667), .Z(n18079) );
  XNOR U17882 ( .A(p_input[1704]), .B(n18080), .Z(n17667) );
  AND U17883 ( .A(n643), .B(n18081), .Z(n18080) );
  XOR U17884 ( .A(p_input[1720]), .B(p_input[1704]), .Z(n18081) );
  XNOR U17885 ( .A(n17664), .B(n18076), .Z(n18078) );
  XOR U17886 ( .A(n18082), .B(n18083), .Z(n17664) );
  AND U17887 ( .A(n640), .B(n18084), .Z(n18083) );
  XOR U17888 ( .A(p_input[1688]), .B(p_input[1672]), .Z(n18084) );
  XOR U17889 ( .A(n18085), .B(n18086), .Z(n18076) );
  AND U17890 ( .A(n18087), .B(n18088), .Z(n18086) );
  XOR U17891 ( .A(n18085), .B(n17679), .Z(n18088) );
  XNOR U17892 ( .A(p_input[1703]), .B(n18089), .Z(n17679) );
  AND U17893 ( .A(n643), .B(n18090), .Z(n18089) );
  XOR U17894 ( .A(p_input[1719]), .B(p_input[1703]), .Z(n18090) );
  XNOR U17895 ( .A(n17676), .B(n18085), .Z(n18087) );
  XOR U17896 ( .A(n18091), .B(n18092), .Z(n17676) );
  AND U17897 ( .A(n640), .B(n18093), .Z(n18092) );
  XOR U17898 ( .A(p_input[1687]), .B(p_input[1671]), .Z(n18093) );
  XOR U17899 ( .A(n18094), .B(n18095), .Z(n18085) );
  AND U17900 ( .A(n18096), .B(n18097), .Z(n18095) );
  XOR U17901 ( .A(n18094), .B(n17691), .Z(n18097) );
  XNOR U17902 ( .A(p_input[1702]), .B(n18098), .Z(n17691) );
  AND U17903 ( .A(n643), .B(n18099), .Z(n18098) );
  XOR U17904 ( .A(p_input[1718]), .B(p_input[1702]), .Z(n18099) );
  XNOR U17905 ( .A(n17688), .B(n18094), .Z(n18096) );
  XOR U17906 ( .A(n18100), .B(n18101), .Z(n17688) );
  AND U17907 ( .A(n640), .B(n18102), .Z(n18101) );
  XOR U17908 ( .A(p_input[1686]), .B(p_input[1670]), .Z(n18102) );
  XOR U17909 ( .A(n18103), .B(n18104), .Z(n18094) );
  AND U17910 ( .A(n18105), .B(n18106), .Z(n18104) );
  XOR U17911 ( .A(n18103), .B(n17703), .Z(n18106) );
  XNOR U17912 ( .A(p_input[1701]), .B(n18107), .Z(n17703) );
  AND U17913 ( .A(n643), .B(n18108), .Z(n18107) );
  XOR U17914 ( .A(p_input[1717]), .B(p_input[1701]), .Z(n18108) );
  XNOR U17915 ( .A(n17700), .B(n18103), .Z(n18105) );
  XOR U17916 ( .A(n18109), .B(n18110), .Z(n17700) );
  AND U17917 ( .A(n640), .B(n18111), .Z(n18110) );
  XOR U17918 ( .A(p_input[1685]), .B(p_input[1669]), .Z(n18111) );
  XOR U17919 ( .A(n18112), .B(n18113), .Z(n18103) );
  AND U17920 ( .A(n18114), .B(n18115), .Z(n18113) );
  XOR U17921 ( .A(n18112), .B(n17715), .Z(n18115) );
  XNOR U17922 ( .A(p_input[1700]), .B(n18116), .Z(n17715) );
  AND U17923 ( .A(n643), .B(n18117), .Z(n18116) );
  XOR U17924 ( .A(p_input[1716]), .B(p_input[1700]), .Z(n18117) );
  XNOR U17925 ( .A(n17712), .B(n18112), .Z(n18114) );
  XOR U17926 ( .A(n18118), .B(n18119), .Z(n17712) );
  AND U17927 ( .A(n640), .B(n18120), .Z(n18119) );
  XOR U17928 ( .A(p_input[1684]), .B(p_input[1668]), .Z(n18120) );
  XOR U17929 ( .A(n18121), .B(n18122), .Z(n18112) );
  AND U17930 ( .A(n18123), .B(n18124), .Z(n18122) );
  XOR U17931 ( .A(n18121), .B(n17727), .Z(n18124) );
  XNOR U17932 ( .A(p_input[1699]), .B(n18125), .Z(n17727) );
  AND U17933 ( .A(n643), .B(n18126), .Z(n18125) );
  XOR U17934 ( .A(p_input[1715]), .B(p_input[1699]), .Z(n18126) );
  XNOR U17935 ( .A(n17724), .B(n18121), .Z(n18123) );
  XOR U17936 ( .A(n18127), .B(n18128), .Z(n17724) );
  AND U17937 ( .A(n640), .B(n18129), .Z(n18128) );
  XOR U17938 ( .A(p_input[1683]), .B(p_input[1667]), .Z(n18129) );
  XOR U17939 ( .A(n18130), .B(n18131), .Z(n18121) );
  AND U17940 ( .A(n18132), .B(n18133), .Z(n18131) );
  XOR U17941 ( .A(n18130), .B(n17739), .Z(n18133) );
  XNOR U17942 ( .A(p_input[1698]), .B(n18134), .Z(n17739) );
  AND U17943 ( .A(n643), .B(n18135), .Z(n18134) );
  XOR U17944 ( .A(p_input[1714]), .B(p_input[1698]), .Z(n18135) );
  XNOR U17945 ( .A(n17736), .B(n18130), .Z(n18132) );
  XOR U17946 ( .A(n18136), .B(n18137), .Z(n17736) );
  AND U17947 ( .A(n640), .B(n18138), .Z(n18137) );
  XOR U17948 ( .A(p_input[1682]), .B(p_input[1666]), .Z(n18138) );
  XOR U17949 ( .A(n18139), .B(n18140), .Z(n18130) );
  AND U17950 ( .A(n18141), .B(n18142), .Z(n18140) );
  XNOR U17951 ( .A(n18143), .B(n17752), .Z(n18142) );
  XNOR U17952 ( .A(p_input[1697]), .B(n18144), .Z(n17752) );
  AND U17953 ( .A(n643), .B(n18145), .Z(n18144) );
  XNOR U17954 ( .A(p_input[1713]), .B(n18146), .Z(n18145) );
  IV U17955 ( .A(p_input[1697]), .Z(n18146) );
  XNOR U17956 ( .A(n17749), .B(n18139), .Z(n18141) );
  XNOR U17957 ( .A(p_input[1665]), .B(n18147), .Z(n17749) );
  AND U17958 ( .A(n640), .B(n18148), .Z(n18147) );
  XOR U17959 ( .A(p_input[1681]), .B(p_input[1665]), .Z(n18148) );
  IV U17960 ( .A(n18143), .Z(n18139) );
  AND U17961 ( .A(n18014), .B(n18017), .Z(n18143) );
  XOR U17962 ( .A(p_input[1696]), .B(n18149), .Z(n18017) );
  AND U17963 ( .A(n643), .B(n18150), .Z(n18149) );
  XOR U17964 ( .A(p_input[1712]), .B(p_input[1696]), .Z(n18150) );
  XOR U17965 ( .A(n18151), .B(n18152), .Z(n643) );
  AND U17966 ( .A(n18153), .B(n18154), .Z(n18152) );
  XNOR U17967 ( .A(p_input[1727]), .B(n18151), .Z(n18154) );
  XOR U17968 ( .A(n18151), .B(p_input[1711]), .Z(n18153) );
  XOR U17969 ( .A(n18155), .B(n18156), .Z(n18151) );
  AND U17970 ( .A(n18157), .B(n18158), .Z(n18156) );
  XNOR U17971 ( .A(p_input[1726]), .B(n18155), .Z(n18158) );
  XOR U17972 ( .A(n18155), .B(p_input[1710]), .Z(n18157) );
  XOR U17973 ( .A(n18159), .B(n18160), .Z(n18155) );
  AND U17974 ( .A(n18161), .B(n18162), .Z(n18160) );
  XNOR U17975 ( .A(p_input[1725]), .B(n18159), .Z(n18162) );
  XOR U17976 ( .A(n18159), .B(p_input[1709]), .Z(n18161) );
  XOR U17977 ( .A(n18163), .B(n18164), .Z(n18159) );
  AND U17978 ( .A(n18165), .B(n18166), .Z(n18164) );
  XNOR U17979 ( .A(p_input[1724]), .B(n18163), .Z(n18166) );
  XOR U17980 ( .A(n18163), .B(p_input[1708]), .Z(n18165) );
  XOR U17981 ( .A(n18167), .B(n18168), .Z(n18163) );
  AND U17982 ( .A(n18169), .B(n18170), .Z(n18168) );
  XNOR U17983 ( .A(p_input[1723]), .B(n18167), .Z(n18170) );
  XOR U17984 ( .A(n18167), .B(p_input[1707]), .Z(n18169) );
  XOR U17985 ( .A(n18171), .B(n18172), .Z(n18167) );
  AND U17986 ( .A(n18173), .B(n18174), .Z(n18172) );
  XNOR U17987 ( .A(p_input[1722]), .B(n18171), .Z(n18174) );
  XOR U17988 ( .A(n18171), .B(p_input[1706]), .Z(n18173) );
  XOR U17989 ( .A(n18175), .B(n18176), .Z(n18171) );
  AND U17990 ( .A(n18177), .B(n18178), .Z(n18176) );
  XNOR U17991 ( .A(p_input[1721]), .B(n18175), .Z(n18178) );
  XOR U17992 ( .A(n18175), .B(p_input[1705]), .Z(n18177) );
  XOR U17993 ( .A(n18179), .B(n18180), .Z(n18175) );
  AND U17994 ( .A(n18181), .B(n18182), .Z(n18180) );
  XNOR U17995 ( .A(p_input[1720]), .B(n18179), .Z(n18182) );
  XOR U17996 ( .A(n18179), .B(p_input[1704]), .Z(n18181) );
  XOR U17997 ( .A(n18183), .B(n18184), .Z(n18179) );
  AND U17998 ( .A(n18185), .B(n18186), .Z(n18184) );
  XNOR U17999 ( .A(p_input[1719]), .B(n18183), .Z(n18186) );
  XOR U18000 ( .A(n18183), .B(p_input[1703]), .Z(n18185) );
  XOR U18001 ( .A(n18187), .B(n18188), .Z(n18183) );
  AND U18002 ( .A(n18189), .B(n18190), .Z(n18188) );
  XNOR U18003 ( .A(p_input[1718]), .B(n18187), .Z(n18190) );
  XOR U18004 ( .A(n18187), .B(p_input[1702]), .Z(n18189) );
  XOR U18005 ( .A(n18191), .B(n18192), .Z(n18187) );
  AND U18006 ( .A(n18193), .B(n18194), .Z(n18192) );
  XNOR U18007 ( .A(p_input[1717]), .B(n18191), .Z(n18194) );
  XOR U18008 ( .A(n18191), .B(p_input[1701]), .Z(n18193) );
  XOR U18009 ( .A(n18195), .B(n18196), .Z(n18191) );
  AND U18010 ( .A(n18197), .B(n18198), .Z(n18196) );
  XNOR U18011 ( .A(p_input[1716]), .B(n18195), .Z(n18198) );
  XOR U18012 ( .A(n18195), .B(p_input[1700]), .Z(n18197) );
  XOR U18013 ( .A(n18199), .B(n18200), .Z(n18195) );
  AND U18014 ( .A(n18201), .B(n18202), .Z(n18200) );
  XNOR U18015 ( .A(p_input[1715]), .B(n18199), .Z(n18202) );
  XOR U18016 ( .A(n18199), .B(p_input[1699]), .Z(n18201) );
  XOR U18017 ( .A(n18203), .B(n18204), .Z(n18199) );
  AND U18018 ( .A(n18205), .B(n18206), .Z(n18204) );
  XNOR U18019 ( .A(p_input[1714]), .B(n18203), .Z(n18206) );
  XOR U18020 ( .A(n18203), .B(p_input[1698]), .Z(n18205) );
  XNOR U18021 ( .A(n18207), .B(n18208), .Z(n18203) );
  AND U18022 ( .A(n18209), .B(n18210), .Z(n18208) );
  XOR U18023 ( .A(p_input[1713]), .B(n18207), .Z(n18210) );
  XNOR U18024 ( .A(p_input[1697]), .B(n18207), .Z(n18209) );
  AND U18025 ( .A(p_input[1712]), .B(n18211), .Z(n18207) );
  IV U18026 ( .A(p_input[1696]), .Z(n18211) );
  XNOR U18027 ( .A(p_input[1664]), .B(n18212), .Z(n18014) );
  AND U18028 ( .A(n640), .B(n18213), .Z(n18212) );
  XOR U18029 ( .A(p_input[1680]), .B(p_input[1664]), .Z(n18213) );
  XOR U18030 ( .A(n18214), .B(n18215), .Z(n640) );
  AND U18031 ( .A(n18216), .B(n18217), .Z(n18215) );
  XNOR U18032 ( .A(p_input[1695]), .B(n18214), .Z(n18217) );
  XOR U18033 ( .A(n18214), .B(p_input[1679]), .Z(n18216) );
  XOR U18034 ( .A(n18218), .B(n18219), .Z(n18214) );
  AND U18035 ( .A(n18220), .B(n18221), .Z(n18219) );
  XNOR U18036 ( .A(p_input[1694]), .B(n18218), .Z(n18221) );
  XNOR U18037 ( .A(n18218), .B(n18028), .Z(n18220) );
  IV U18038 ( .A(p_input[1678]), .Z(n18028) );
  XOR U18039 ( .A(n18222), .B(n18223), .Z(n18218) );
  AND U18040 ( .A(n18224), .B(n18225), .Z(n18223) );
  XNOR U18041 ( .A(p_input[1693]), .B(n18222), .Z(n18225) );
  XNOR U18042 ( .A(n18222), .B(n18037), .Z(n18224) );
  IV U18043 ( .A(p_input[1677]), .Z(n18037) );
  XOR U18044 ( .A(n18226), .B(n18227), .Z(n18222) );
  AND U18045 ( .A(n18228), .B(n18229), .Z(n18227) );
  XNOR U18046 ( .A(p_input[1692]), .B(n18226), .Z(n18229) );
  XNOR U18047 ( .A(n18226), .B(n18046), .Z(n18228) );
  IV U18048 ( .A(p_input[1676]), .Z(n18046) );
  XOR U18049 ( .A(n18230), .B(n18231), .Z(n18226) );
  AND U18050 ( .A(n18232), .B(n18233), .Z(n18231) );
  XNOR U18051 ( .A(p_input[1691]), .B(n18230), .Z(n18233) );
  XNOR U18052 ( .A(n18230), .B(n18055), .Z(n18232) );
  IV U18053 ( .A(p_input[1675]), .Z(n18055) );
  XOR U18054 ( .A(n18234), .B(n18235), .Z(n18230) );
  AND U18055 ( .A(n18236), .B(n18237), .Z(n18235) );
  XNOR U18056 ( .A(p_input[1690]), .B(n18234), .Z(n18237) );
  XNOR U18057 ( .A(n18234), .B(n18064), .Z(n18236) );
  IV U18058 ( .A(p_input[1674]), .Z(n18064) );
  XOR U18059 ( .A(n18238), .B(n18239), .Z(n18234) );
  AND U18060 ( .A(n18240), .B(n18241), .Z(n18239) );
  XNOR U18061 ( .A(p_input[1689]), .B(n18238), .Z(n18241) );
  XNOR U18062 ( .A(n18238), .B(n18073), .Z(n18240) );
  IV U18063 ( .A(p_input[1673]), .Z(n18073) );
  XOR U18064 ( .A(n18242), .B(n18243), .Z(n18238) );
  AND U18065 ( .A(n18244), .B(n18245), .Z(n18243) );
  XNOR U18066 ( .A(p_input[1688]), .B(n18242), .Z(n18245) );
  XNOR U18067 ( .A(n18242), .B(n18082), .Z(n18244) );
  IV U18068 ( .A(p_input[1672]), .Z(n18082) );
  XOR U18069 ( .A(n18246), .B(n18247), .Z(n18242) );
  AND U18070 ( .A(n18248), .B(n18249), .Z(n18247) );
  XNOR U18071 ( .A(p_input[1687]), .B(n18246), .Z(n18249) );
  XNOR U18072 ( .A(n18246), .B(n18091), .Z(n18248) );
  IV U18073 ( .A(p_input[1671]), .Z(n18091) );
  XOR U18074 ( .A(n18250), .B(n18251), .Z(n18246) );
  AND U18075 ( .A(n18252), .B(n18253), .Z(n18251) );
  XNOR U18076 ( .A(p_input[1686]), .B(n18250), .Z(n18253) );
  XNOR U18077 ( .A(n18250), .B(n18100), .Z(n18252) );
  IV U18078 ( .A(p_input[1670]), .Z(n18100) );
  XOR U18079 ( .A(n18254), .B(n18255), .Z(n18250) );
  AND U18080 ( .A(n18256), .B(n18257), .Z(n18255) );
  XNOR U18081 ( .A(p_input[1685]), .B(n18254), .Z(n18257) );
  XNOR U18082 ( .A(n18254), .B(n18109), .Z(n18256) );
  IV U18083 ( .A(p_input[1669]), .Z(n18109) );
  XOR U18084 ( .A(n18258), .B(n18259), .Z(n18254) );
  AND U18085 ( .A(n18260), .B(n18261), .Z(n18259) );
  XNOR U18086 ( .A(p_input[1684]), .B(n18258), .Z(n18261) );
  XNOR U18087 ( .A(n18258), .B(n18118), .Z(n18260) );
  IV U18088 ( .A(p_input[1668]), .Z(n18118) );
  XOR U18089 ( .A(n18262), .B(n18263), .Z(n18258) );
  AND U18090 ( .A(n18264), .B(n18265), .Z(n18263) );
  XNOR U18091 ( .A(p_input[1683]), .B(n18262), .Z(n18265) );
  XNOR U18092 ( .A(n18262), .B(n18127), .Z(n18264) );
  IV U18093 ( .A(p_input[1667]), .Z(n18127) );
  XOR U18094 ( .A(n18266), .B(n18267), .Z(n18262) );
  AND U18095 ( .A(n18268), .B(n18269), .Z(n18267) );
  XNOR U18096 ( .A(p_input[1682]), .B(n18266), .Z(n18269) );
  XNOR U18097 ( .A(n18266), .B(n18136), .Z(n18268) );
  IV U18098 ( .A(p_input[1666]), .Z(n18136) );
  XNOR U18099 ( .A(n18270), .B(n18271), .Z(n18266) );
  AND U18100 ( .A(n18272), .B(n18273), .Z(n18271) );
  XOR U18101 ( .A(p_input[1681]), .B(n18270), .Z(n18273) );
  XNOR U18102 ( .A(p_input[1665]), .B(n18270), .Z(n18272) );
  AND U18103 ( .A(p_input[1680]), .B(n18274), .Z(n18270) );
  IV U18104 ( .A(p_input[1664]), .Z(n18274) );
  XOR U18105 ( .A(n18275), .B(n18276), .Z(n17390) );
  AND U18106 ( .A(n796), .B(n18277), .Z(n18276) );
  XNOR U18107 ( .A(n18278), .B(n18275), .Z(n18277) );
  XOR U18108 ( .A(n18279), .B(n18280), .Z(n796) );
  AND U18109 ( .A(n18281), .B(n18282), .Z(n18280) );
  XNOR U18110 ( .A(n17402), .B(n18279), .Z(n18282) );
  AND U18111 ( .A(n18283), .B(n18284), .Z(n17402) );
  XOR U18112 ( .A(n18279), .B(n17401), .Z(n18281) );
  AND U18113 ( .A(n18285), .B(n18286), .Z(n17401) );
  XOR U18114 ( .A(n18287), .B(n18288), .Z(n18279) );
  AND U18115 ( .A(n18289), .B(n18290), .Z(n18288) );
  XOR U18116 ( .A(n18287), .B(n17414), .Z(n18290) );
  XOR U18117 ( .A(n18291), .B(n18292), .Z(n17414) );
  AND U18118 ( .A(n499), .B(n18293), .Z(n18292) );
  XOR U18119 ( .A(n18294), .B(n18291), .Z(n18293) );
  XNOR U18120 ( .A(n17411), .B(n18287), .Z(n18289) );
  XOR U18121 ( .A(n18295), .B(n18296), .Z(n17411) );
  AND U18122 ( .A(n496), .B(n18297), .Z(n18296) );
  XOR U18123 ( .A(n18298), .B(n18295), .Z(n18297) );
  XOR U18124 ( .A(n18299), .B(n18300), .Z(n18287) );
  AND U18125 ( .A(n18301), .B(n18302), .Z(n18300) );
  XOR U18126 ( .A(n18299), .B(n17426), .Z(n18302) );
  XOR U18127 ( .A(n18303), .B(n18304), .Z(n17426) );
  AND U18128 ( .A(n499), .B(n18305), .Z(n18304) );
  XOR U18129 ( .A(n18306), .B(n18303), .Z(n18305) );
  XNOR U18130 ( .A(n17423), .B(n18299), .Z(n18301) );
  XOR U18131 ( .A(n18307), .B(n18308), .Z(n17423) );
  AND U18132 ( .A(n496), .B(n18309), .Z(n18308) );
  XOR U18133 ( .A(n18310), .B(n18307), .Z(n18309) );
  XOR U18134 ( .A(n18311), .B(n18312), .Z(n18299) );
  AND U18135 ( .A(n18313), .B(n18314), .Z(n18312) );
  XOR U18136 ( .A(n18311), .B(n17438), .Z(n18314) );
  XOR U18137 ( .A(n18315), .B(n18316), .Z(n17438) );
  AND U18138 ( .A(n499), .B(n18317), .Z(n18316) );
  XOR U18139 ( .A(n18318), .B(n18315), .Z(n18317) );
  XNOR U18140 ( .A(n17435), .B(n18311), .Z(n18313) );
  XOR U18141 ( .A(n18319), .B(n18320), .Z(n17435) );
  AND U18142 ( .A(n496), .B(n18321), .Z(n18320) );
  XOR U18143 ( .A(n18322), .B(n18319), .Z(n18321) );
  XOR U18144 ( .A(n18323), .B(n18324), .Z(n18311) );
  AND U18145 ( .A(n18325), .B(n18326), .Z(n18324) );
  XOR U18146 ( .A(n18323), .B(n17450), .Z(n18326) );
  XOR U18147 ( .A(n18327), .B(n18328), .Z(n17450) );
  AND U18148 ( .A(n499), .B(n18329), .Z(n18328) );
  XOR U18149 ( .A(n18330), .B(n18327), .Z(n18329) );
  XNOR U18150 ( .A(n17447), .B(n18323), .Z(n18325) );
  XOR U18151 ( .A(n18331), .B(n18332), .Z(n17447) );
  AND U18152 ( .A(n496), .B(n18333), .Z(n18332) );
  XOR U18153 ( .A(n18334), .B(n18331), .Z(n18333) );
  XOR U18154 ( .A(n18335), .B(n18336), .Z(n18323) );
  AND U18155 ( .A(n18337), .B(n18338), .Z(n18336) );
  XOR U18156 ( .A(n18335), .B(n17462), .Z(n18338) );
  XOR U18157 ( .A(n18339), .B(n18340), .Z(n17462) );
  AND U18158 ( .A(n499), .B(n18341), .Z(n18340) );
  XOR U18159 ( .A(n18342), .B(n18339), .Z(n18341) );
  XNOR U18160 ( .A(n17459), .B(n18335), .Z(n18337) );
  XOR U18161 ( .A(n18343), .B(n18344), .Z(n17459) );
  AND U18162 ( .A(n496), .B(n18345), .Z(n18344) );
  XOR U18163 ( .A(n18346), .B(n18343), .Z(n18345) );
  XOR U18164 ( .A(n18347), .B(n18348), .Z(n18335) );
  AND U18165 ( .A(n18349), .B(n18350), .Z(n18348) );
  XOR U18166 ( .A(n18347), .B(n17474), .Z(n18350) );
  XOR U18167 ( .A(n18351), .B(n18352), .Z(n17474) );
  AND U18168 ( .A(n499), .B(n18353), .Z(n18352) );
  XOR U18169 ( .A(n18354), .B(n18351), .Z(n18353) );
  XNOR U18170 ( .A(n17471), .B(n18347), .Z(n18349) );
  XOR U18171 ( .A(n18355), .B(n18356), .Z(n17471) );
  AND U18172 ( .A(n496), .B(n18357), .Z(n18356) );
  XOR U18173 ( .A(n18358), .B(n18355), .Z(n18357) );
  XOR U18174 ( .A(n18359), .B(n18360), .Z(n18347) );
  AND U18175 ( .A(n18361), .B(n18362), .Z(n18360) );
  XOR U18176 ( .A(n18359), .B(n17486), .Z(n18362) );
  XOR U18177 ( .A(n18363), .B(n18364), .Z(n17486) );
  AND U18178 ( .A(n499), .B(n18365), .Z(n18364) );
  XOR U18179 ( .A(n18366), .B(n18363), .Z(n18365) );
  XNOR U18180 ( .A(n17483), .B(n18359), .Z(n18361) );
  XOR U18181 ( .A(n18367), .B(n18368), .Z(n17483) );
  AND U18182 ( .A(n496), .B(n18369), .Z(n18368) );
  XOR U18183 ( .A(n18370), .B(n18367), .Z(n18369) );
  XOR U18184 ( .A(n18371), .B(n18372), .Z(n18359) );
  AND U18185 ( .A(n18373), .B(n18374), .Z(n18372) );
  XOR U18186 ( .A(n18371), .B(n17498), .Z(n18374) );
  XOR U18187 ( .A(n18375), .B(n18376), .Z(n17498) );
  AND U18188 ( .A(n499), .B(n18377), .Z(n18376) );
  XOR U18189 ( .A(n18378), .B(n18375), .Z(n18377) );
  XNOR U18190 ( .A(n17495), .B(n18371), .Z(n18373) );
  XOR U18191 ( .A(n18379), .B(n18380), .Z(n17495) );
  AND U18192 ( .A(n496), .B(n18381), .Z(n18380) );
  XOR U18193 ( .A(n18382), .B(n18379), .Z(n18381) );
  XOR U18194 ( .A(n18383), .B(n18384), .Z(n18371) );
  AND U18195 ( .A(n18385), .B(n18386), .Z(n18384) );
  XOR U18196 ( .A(n18383), .B(n17510), .Z(n18386) );
  XOR U18197 ( .A(n18387), .B(n18388), .Z(n17510) );
  AND U18198 ( .A(n499), .B(n18389), .Z(n18388) );
  XOR U18199 ( .A(n18390), .B(n18387), .Z(n18389) );
  XNOR U18200 ( .A(n17507), .B(n18383), .Z(n18385) );
  XOR U18201 ( .A(n18391), .B(n18392), .Z(n17507) );
  AND U18202 ( .A(n496), .B(n18393), .Z(n18392) );
  XOR U18203 ( .A(n18394), .B(n18391), .Z(n18393) );
  XOR U18204 ( .A(n18395), .B(n18396), .Z(n18383) );
  AND U18205 ( .A(n18397), .B(n18398), .Z(n18396) );
  XOR U18206 ( .A(n18395), .B(n17522), .Z(n18398) );
  XOR U18207 ( .A(n18399), .B(n18400), .Z(n17522) );
  AND U18208 ( .A(n499), .B(n18401), .Z(n18400) );
  XOR U18209 ( .A(n18402), .B(n18399), .Z(n18401) );
  XNOR U18210 ( .A(n17519), .B(n18395), .Z(n18397) );
  XOR U18211 ( .A(n18403), .B(n18404), .Z(n17519) );
  AND U18212 ( .A(n496), .B(n18405), .Z(n18404) );
  XOR U18213 ( .A(n18406), .B(n18403), .Z(n18405) );
  XOR U18214 ( .A(n18407), .B(n18408), .Z(n18395) );
  AND U18215 ( .A(n18409), .B(n18410), .Z(n18408) );
  XOR U18216 ( .A(n18407), .B(n17534), .Z(n18410) );
  XOR U18217 ( .A(n18411), .B(n18412), .Z(n17534) );
  AND U18218 ( .A(n499), .B(n18413), .Z(n18412) );
  XOR U18219 ( .A(n18414), .B(n18411), .Z(n18413) );
  XNOR U18220 ( .A(n17531), .B(n18407), .Z(n18409) );
  XOR U18221 ( .A(n18415), .B(n18416), .Z(n17531) );
  AND U18222 ( .A(n496), .B(n18417), .Z(n18416) );
  XOR U18223 ( .A(n18418), .B(n18415), .Z(n18417) );
  XOR U18224 ( .A(n18419), .B(n18420), .Z(n18407) );
  AND U18225 ( .A(n18421), .B(n18422), .Z(n18420) );
  XOR U18226 ( .A(n18419), .B(n17546), .Z(n18422) );
  XOR U18227 ( .A(n18423), .B(n18424), .Z(n17546) );
  AND U18228 ( .A(n499), .B(n18425), .Z(n18424) );
  XOR U18229 ( .A(n18426), .B(n18423), .Z(n18425) );
  XNOR U18230 ( .A(n17543), .B(n18419), .Z(n18421) );
  XOR U18231 ( .A(n18427), .B(n18428), .Z(n17543) );
  AND U18232 ( .A(n496), .B(n18429), .Z(n18428) );
  XOR U18233 ( .A(n18430), .B(n18427), .Z(n18429) );
  XOR U18234 ( .A(n18431), .B(n18432), .Z(n18419) );
  AND U18235 ( .A(n18433), .B(n18434), .Z(n18432) );
  XOR U18236 ( .A(n18431), .B(n17558), .Z(n18434) );
  XOR U18237 ( .A(n18435), .B(n18436), .Z(n17558) );
  AND U18238 ( .A(n499), .B(n18437), .Z(n18436) );
  XOR U18239 ( .A(n18438), .B(n18435), .Z(n18437) );
  XNOR U18240 ( .A(n17555), .B(n18431), .Z(n18433) );
  XOR U18241 ( .A(n18439), .B(n18440), .Z(n17555) );
  AND U18242 ( .A(n496), .B(n18441), .Z(n18440) );
  XOR U18243 ( .A(n18442), .B(n18439), .Z(n18441) );
  XOR U18244 ( .A(n18443), .B(n18444), .Z(n18431) );
  AND U18245 ( .A(n18445), .B(n18446), .Z(n18444) );
  XNOR U18246 ( .A(n18447), .B(n17571), .Z(n18446) );
  XOR U18247 ( .A(n18448), .B(n18449), .Z(n17571) );
  AND U18248 ( .A(n499), .B(n18450), .Z(n18449) );
  XOR U18249 ( .A(n18448), .B(n18451), .Z(n18450) );
  XNOR U18250 ( .A(n17568), .B(n18443), .Z(n18445) );
  XOR U18251 ( .A(n18452), .B(n18453), .Z(n17568) );
  AND U18252 ( .A(n496), .B(n18454), .Z(n18453) );
  XOR U18253 ( .A(n18452), .B(n18455), .Z(n18454) );
  IV U18254 ( .A(n18447), .Z(n18443) );
  AND U18255 ( .A(n18275), .B(n18278), .Z(n18447) );
  XNOR U18256 ( .A(n18456), .B(n18457), .Z(n18278) );
  AND U18257 ( .A(n499), .B(n18458), .Z(n18457) );
  XNOR U18258 ( .A(n18459), .B(n18456), .Z(n18458) );
  XOR U18259 ( .A(n18460), .B(n18461), .Z(n499) );
  AND U18260 ( .A(n18462), .B(n18463), .Z(n18461) );
  XNOR U18261 ( .A(n18283), .B(n18460), .Z(n18463) );
  AND U18262 ( .A(p_input[1663]), .B(p_input[1647]), .Z(n18283) );
  XOR U18263 ( .A(n18460), .B(n18284), .Z(n18462) );
  AND U18264 ( .A(p_input[1631]), .B(p_input[1615]), .Z(n18284) );
  XOR U18265 ( .A(n18464), .B(n18465), .Z(n18460) );
  AND U18266 ( .A(n18466), .B(n18467), .Z(n18465) );
  XOR U18267 ( .A(n18464), .B(n18294), .Z(n18467) );
  XNOR U18268 ( .A(p_input[1646]), .B(n18468), .Z(n18294) );
  AND U18269 ( .A(n651), .B(n18469), .Z(n18468) );
  XOR U18270 ( .A(p_input[1662]), .B(p_input[1646]), .Z(n18469) );
  XNOR U18271 ( .A(n18291), .B(n18464), .Z(n18466) );
  XOR U18272 ( .A(n18470), .B(n18471), .Z(n18291) );
  AND U18273 ( .A(n649), .B(n18472), .Z(n18471) );
  XOR U18274 ( .A(p_input[1630]), .B(p_input[1614]), .Z(n18472) );
  XOR U18275 ( .A(n18473), .B(n18474), .Z(n18464) );
  AND U18276 ( .A(n18475), .B(n18476), .Z(n18474) );
  XOR U18277 ( .A(n18473), .B(n18306), .Z(n18476) );
  XNOR U18278 ( .A(p_input[1645]), .B(n18477), .Z(n18306) );
  AND U18279 ( .A(n651), .B(n18478), .Z(n18477) );
  XOR U18280 ( .A(p_input[1661]), .B(p_input[1645]), .Z(n18478) );
  XNOR U18281 ( .A(n18303), .B(n18473), .Z(n18475) );
  XOR U18282 ( .A(n18479), .B(n18480), .Z(n18303) );
  AND U18283 ( .A(n649), .B(n18481), .Z(n18480) );
  XOR U18284 ( .A(p_input[1629]), .B(p_input[1613]), .Z(n18481) );
  XOR U18285 ( .A(n18482), .B(n18483), .Z(n18473) );
  AND U18286 ( .A(n18484), .B(n18485), .Z(n18483) );
  XOR U18287 ( .A(n18482), .B(n18318), .Z(n18485) );
  XNOR U18288 ( .A(p_input[1644]), .B(n18486), .Z(n18318) );
  AND U18289 ( .A(n651), .B(n18487), .Z(n18486) );
  XOR U18290 ( .A(p_input[1660]), .B(p_input[1644]), .Z(n18487) );
  XNOR U18291 ( .A(n18315), .B(n18482), .Z(n18484) );
  XOR U18292 ( .A(n18488), .B(n18489), .Z(n18315) );
  AND U18293 ( .A(n649), .B(n18490), .Z(n18489) );
  XOR U18294 ( .A(p_input[1628]), .B(p_input[1612]), .Z(n18490) );
  XOR U18295 ( .A(n18491), .B(n18492), .Z(n18482) );
  AND U18296 ( .A(n18493), .B(n18494), .Z(n18492) );
  XOR U18297 ( .A(n18491), .B(n18330), .Z(n18494) );
  XNOR U18298 ( .A(p_input[1643]), .B(n18495), .Z(n18330) );
  AND U18299 ( .A(n651), .B(n18496), .Z(n18495) );
  XOR U18300 ( .A(p_input[1659]), .B(p_input[1643]), .Z(n18496) );
  XNOR U18301 ( .A(n18327), .B(n18491), .Z(n18493) );
  XOR U18302 ( .A(n18497), .B(n18498), .Z(n18327) );
  AND U18303 ( .A(n649), .B(n18499), .Z(n18498) );
  XOR U18304 ( .A(p_input[1627]), .B(p_input[1611]), .Z(n18499) );
  XOR U18305 ( .A(n18500), .B(n18501), .Z(n18491) );
  AND U18306 ( .A(n18502), .B(n18503), .Z(n18501) );
  XOR U18307 ( .A(n18500), .B(n18342), .Z(n18503) );
  XNOR U18308 ( .A(p_input[1642]), .B(n18504), .Z(n18342) );
  AND U18309 ( .A(n651), .B(n18505), .Z(n18504) );
  XOR U18310 ( .A(p_input[1658]), .B(p_input[1642]), .Z(n18505) );
  XNOR U18311 ( .A(n18339), .B(n18500), .Z(n18502) );
  XOR U18312 ( .A(n18506), .B(n18507), .Z(n18339) );
  AND U18313 ( .A(n649), .B(n18508), .Z(n18507) );
  XOR U18314 ( .A(p_input[1626]), .B(p_input[1610]), .Z(n18508) );
  XOR U18315 ( .A(n18509), .B(n18510), .Z(n18500) );
  AND U18316 ( .A(n18511), .B(n18512), .Z(n18510) );
  XOR U18317 ( .A(n18509), .B(n18354), .Z(n18512) );
  XNOR U18318 ( .A(p_input[1641]), .B(n18513), .Z(n18354) );
  AND U18319 ( .A(n651), .B(n18514), .Z(n18513) );
  XOR U18320 ( .A(p_input[1657]), .B(p_input[1641]), .Z(n18514) );
  XNOR U18321 ( .A(n18351), .B(n18509), .Z(n18511) );
  XOR U18322 ( .A(n18515), .B(n18516), .Z(n18351) );
  AND U18323 ( .A(n649), .B(n18517), .Z(n18516) );
  XOR U18324 ( .A(p_input[1625]), .B(p_input[1609]), .Z(n18517) );
  XOR U18325 ( .A(n18518), .B(n18519), .Z(n18509) );
  AND U18326 ( .A(n18520), .B(n18521), .Z(n18519) );
  XOR U18327 ( .A(n18518), .B(n18366), .Z(n18521) );
  XNOR U18328 ( .A(p_input[1640]), .B(n18522), .Z(n18366) );
  AND U18329 ( .A(n651), .B(n18523), .Z(n18522) );
  XOR U18330 ( .A(p_input[1656]), .B(p_input[1640]), .Z(n18523) );
  XNOR U18331 ( .A(n18363), .B(n18518), .Z(n18520) );
  XOR U18332 ( .A(n18524), .B(n18525), .Z(n18363) );
  AND U18333 ( .A(n649), .B(n18526), .Z(n18525) );
  XOR U18334 ( .A(p_input[1624]), .B(p_input[1608]), .Z(n18526) );
  XOR U18335 ( .A(n18527), .B(n18528), .Z(n18518) );
  AND U18336 ( .A(n18529), .B(n18530), .Z(n18528) );
  XOR U18337 ( .A(n18527), .B(n18378), .Z(n18530) );
  XNOR U18338 ( .A(p_input[1639]), .B(n18531), .Z(n18378) );
  AND U18339 ( .A(n651), .B(n18532), .Z(n18531) );
  XOR U18340 ( .A(p_input[1655]), .B(p_input[1639]), .Z(n18532) );
  XNOR U18341 ( .A(n18375), .B(n18527), .Z(n18529) );
  XOR U18342 ( .A(n18533), .B(n18534), .Z(n18375) );
  AND U18343 ( .A(n649), .B(n18535), .Z(n18534) );
  XOR U18344 ( .A(p_input[1623]), .B(p_input[1607]), .Z(n18535) );
  XOR U18345 ( .A(n18536), .B(n18537), .Z(n18527) );
  AND U18346 ( .A(n18538), .B(n18539), .Z(n18537) );
  XOR U18347 ( .A(n18536), .B(n18390), .Z(n18539) );
  XNOR U18348 ( .A(p_input[1638]), .B(n18540), .Z(n18390) );
  AND U18349 ( .A(n651), .B(n18541), .Z(n18540) );
  XOR U18350 ( .A(p_input[1654]), .B(p_input[1638]), .Z(n18541) );
  XNOR U18351 ( .A(n18387), .B(n18536), .Z(n18538) );
  XOR U18352 ( .A(n18542), .B(n18543), .Z(n18387) );
  AND U18353 ( .A(n649), .B(n18544), .Z(n18543) );
  XOR U18354 ( .A(p_input[1622]), .B(p_input[1606]), .Z(n18544) );
  XOR U18355 ( .A(n18545), .B(n18546), .Z(n18536) );
  AND U18356 ( .A(n18547), .B(n18548), .Z(n18546) );
  XOR U18357 ( .A(n18545), .B(n18402), .Z(n18548) );
  XNOR U18358 ( .A(p_input[1637]), .B(n18549), .Z(n18402) );
  AND U18359 ( .A(n651), .B(n18550), .Z(n18549) );
  XOR U18360 ( .A(p_input[1653]), .B(p_input[1637]), .Z(n18550) );
  XNOR U18361 ( .A(n18399), .B(n18545), .Z(n18547) );
  XOR U18362 ( .A(n18551), .B(n18552), .Z(n18399) );
  AND U18363 ( .A(n649), .B(n18553), .Z(n18552) );
  XOR U18364 ( .A(p_input[1621]), .B(p_input[1605]), .Z(n18553) );
  XOR U18365 ( .A(n18554), .B(n18555), .Z(n18545) );
  AND U18366 ( .A(n18556), .B(n18557), .Z(n18555) );
  XOR U18367 ( .A(n18554), .B(n18414), .Z(n18557) );
  XNOR U18368 ( .A(p_input[1636]), .B(n18558), .Z(n18414) );
  AND U18369 ( .A(n651), .B(n18559), .Z(n18558) );
  XOR U18370 ( .A(p_input[1652]), .B(p_input[1636]), .Z(n18559) );
  XNOR U18371 ( .A(n18411), .B(n18554), .Z(n18556) );
  XOR U18372 ( .A(n18560), .B(n18561), .Z(n18411) );
  AND U18373 ( .A(n649), .B(n18562), .Z(n18561) );
  XOR U18374 ( .A(p_input[1620]), .B(p_input[1604]), .Z(n18562) );
  XOR U18375 ( .A(n18563), .B(n18564), .Z(n18554) );
  AND U18376 ( .A(n18565), .B(n18566), .Z(n18564) );
  XOR U18377 ( .A(n18563), .B(n18426), .Z(n18566) );
  XNOR U18378 ( .A(p_input[1635]), .B(n18567), .Z(n18426) );
  AND U18379 ( .A(n651), .B(n18568), .Z(n18567) );
  XOR U18380 ( .A(p_input[1651]), .B(p_input[1635]), .Z(n18568) );
  XNOR U18381 ( .A(n18423), .B(n18563), .Z(n18565) );
  XOR U18382 ( .A(n18569), .B(n18570), .Z(n18423) );
  AND U18383 ( .A(n649), .B(n18571), .Z(n18570) );
  XOR U18384 ( .A(p_input[1619]), .B(p_input[1603]), .Z(n18571) );
  XOR U18385 ( .A(n18572), .B(n18573), .Z(n18563) );
  AND U18386 ( .A(n18574), .B(n18575), .Z(n18573) );
  XOR U18387 ( .A(n18572), .B(n18438), .Z(n18575) );
  XNOR U18388 ( .A(p_input[1634]), .B(n18576), .Z(n18438) );
  AND U18389 ( .A(n651), .B(n18577), .Z(n18576) );
  XOR U18390 ( .A(p_input[1650]), .B(p_input[1634]), .Z(n18577) );
  XNOR U18391 ( .A(n18435), .B(n18572), .Z(n18574) );
  XOR U18392 ( .A(n18578), .B(n18579), .Z(n18435) );
  AND U18393 ( .A(n649), .B(n18580), .Z(n18579) );
  XOR U18394 ( .A(p_input[1618]), .B(p_input[1602]), .Z(n18580) );
  XOR U18395 ( .A(n18581), .B(n18582), .Z(n18572) );
  AND U18396 ( .A(n18583), .B(n18584), .Z(n18582) );
  XNOR U18397 ( .A(n18585), .B(n18451), .Z(n18584) );
  XNOR U18398 ( .A(p_input[1633]), .B(n18586), .Z(n18451) );
  AND U18399 ( .A(n651), .B(n18587), .Z(n18586) );
  XNOR U18400 ( .A(p_input[1649]), .B(n18588), .Z(n18587) );
  IV U18401 ( .A(p_input[1633]), .Z(n18588) );
  XNOR U18402 ( .A(n18448), .B(n18581), .Z(n18583) );
  XNOR U18403 ( .A(p_input[1601]), .B(n18589), .Z(n18448) );
  AND U18404 ( .A(n649), .B(n18590), .Z(n18589) );
  XOR U18405 ( .A(p_input[1617]), .B(p_input[1601]), .Z(n18590) );
  IV U18406 ( .A(n18585), .Z(n18581) );
  AND U18407 ( .A(n18456), .B(n18459), .Z(n18585) );
  XOR U18408 ( .A(p_input[1632]), .B(n18591), .Z(n18459) );
  AND U18409 ( .A(n651), .B(n18592), .Z(n18591) );
  XOR U18410 ( .A(p_input[1648]), .B(p_input[1632]), .Z(n18592) );
  XOR U18411 ( .A(n18593), .B(n18594), .Z(n651) );
  AND U18412 ( .A(n18595), .B(n18596), .Z(n18594) );
  XNOR U18413 ( .A(p_input[1663]), .B(n18593), .Z(n18596) );
  XOR U18414 ( .A(n18593), .B(p_input[1647]), .Z(n18595) );
  XOR U18415 ( .A(n18597), .B(n18598), .Z(n18593) );
  AND U18416 ( .A(n18599), .B(n18600), .Z(n18598) );
  XNOR U18417 ( .A(p_input[1662]), .B(n18597), .Z(n18600) );
  XOR U18418 ( .A(n18597), .B(p_input[1646]), .Z(n18599) );
  XOR U18419 ( .A(n18601), .B(n18602), .Z(n18597) );
  AND U18420 ( .A(n18603), .B(n18604), .Z(n18602) );
  XNOR U18421 ( .A(p_input[1661]), .B(n18601), .Z(n18604) );
  XOR U18422 ( .A(n18601), .B(p_input[1645]), .Z(n18603) );
  XOR U18423 ( .A(n18605), .B(n18606), .Z(n18601) );
  AND U18424 ( .A(n18607), .B(n18608), .Z(n18606) );
  XNOR U18425 ( .A(p_input[1660]), .B(n18605), .Z(n18608) );
  XOR U18426 ( .A(n18605), .B(p_input[1644]), .Z(n18607) );
  XOR U18427 ( .A(n18609), .B(n18610), .Z(n18605) );
  AND U18428 ( .A(n18611), .B(n18612), .Z(n18610) );
  XNOR U18429 ( .A(p_input[1659]), .B(n18609), .Z(n18612) );
  XOR U18430 ( .A(n18609), .B(p_input[1643]), .Z(n18611) );
  XOR U18431 ( .A(n18613), .B(n18614), .Z(n18609) );
  AND U18432 ( .A(n18615), .B(n18616), .Z(n18614) );
  XNOR U18433 ( .A(p_input[1658]), .B(n18613), .Z(n18616) );
  XOR U18434 ( .A(n18613), .B(p_input[1642]), .Z(n18615) );
  XOR U18435 ( .A(n18617), .B(n18618), .Z(n18613) );
  AND U18436 ( .A(n18619), .B(n18620), .Z(n18618) );
  XNOR U18437 ( .A(p_input[1657]), .B(n18617), .Z(n18620) );
  XOR U18438 ( .A(n18617), .B(p_input[1641]), .Z(n18619) );
  XOR U18439 ( .A(n18621), .B(n18622), .Z(n18617) );
  AND U18440 ( .A(n18623), .B(n18624), .Z(n18622) );
  XNOR U18441 ( .A(p_input[1656]), .B(n18621), .Z(n18624) );
  XOR U18442 ( .A(n18621), .B(p_input[1640]), .Z(n18623) );
  XOR U18443 ( .A(n18625), .B(n18626), .Z(n18621) );
  AND U18444 ( .A(n18627), .B(n18628), .Z(n18626) );
  XNOR U18445 ( .A(p_input[1655]), .B(n18625), .Z(n18628) );
  XOR U18446 ( .A(n18625), .B(p_input[1639]), .Z(n18627) );
  XOR U18447 ( .A(n18629), .B(n18630), .Z(n18625) );
  AND U18448 ( .A(n18631), .B(n18632), .Z(n18630) );
  XNOR U18449 ( .A(p_input[1654]), .B(n18629), .Z(n18632) );
  XOR U18450 ( .A(n18629), .B(p_input[1638]), .Z(n18631) );
  XOR U18451 ( .A(n18633), .B(n18634), .Z(n18629) );
  AND U18452 ( .A(n18635), .B(n18636), .Z(n18634) );
  XNOR U18453 ( .A(p_input[1653]), .B(n18633), .Z(n18636) );
  XOR U18454 ( .A(n18633), .B(p_input[1637]), .Z(n18635) );
  XOR U18455 ( .A(n18637), .B(n18638), .Z(n18633) );
  AND U18456 ( .A(n18639), .B(n18640), .Z(n18638) );
  XNOR U18457 ( .A(p_input[1652]), .B(n18637), .Z(n18640) );
  XOR U18458 ( .A(n18637), .B(p_input[1636]), .Z(n18639) );
  XOR U18459 ( .A(n18641), .B(n18642), .Z(n18637) );
  AND U18460 ( .A(n18643), .B(n18644), .Z(n18642) );
  XNOR U18461 ( .A(p_input[1651]), .B(n18641), .Z(n18644) );
  XOR U18462 ( .A(n18641), .B(p_input[1635]), .Z(n18643) );
  XOR U18463 ( .A(n18645), .B(n18646), .Z(n18641) );
  AND U18464 ( .A(n18647), .B(n18648), .Z(n18646) );
  XNOR U18465 ( .A(p_input[1650]), .B(n18645), .Z(n18648) );
  XOR U18466 ( .A(n18645), .B(p_input[1634]), .Z(n18647) );
  XNOR U18467 ( .A(n18649), .B(n18650), .Z(n18645) );
  AND U18468 ( .A(n18651), .B(n18652), .Z(n18650) );
  XOR U18469 ( .A(p_input[1649]), .B(n18649), .Z(n18652) );
  XNOR U18470 ( .A(p_input[1633]), .B(n18649), .Z(n18651) );
  AND U18471 ( .A(p_input[1648]), .B(n18653), .Z(n18649) );
  IV U18472 ( .A(p_input[1632]), .Z(n18653) );
  XNOR U18473 ( .A(p_input[1600]), .B(n18654), .Z(n18456) );
  AND U18474 ( .A(n649), .B(n18655), .Z(n18654) );
  XOR U18475 ( .A(p_input[1616]), .B(p_input[1600]), .Z(n18655) );
  XOR U18476 ( .A(n18656), .B(n18657), .Z(n649) );
  AND U18477 ( .A(n18658), .B(n18659), .Z(n18657) );
  XNOR U18478 ( .A(p_input[1631]), .B(n18656), .Z(n18659) );
  XOR U18479 ( .A(n18656), .B(p_input[1615]), .Z(n18658) );
  XOR U18480 ( .A(n18660), .B(n18661), .Z(n18656) );
  AND U18481 ( .A(n18662), .B(n18663), .Z(n18661) );
  XNOR U18482 ( .A(p_input[1630]), .B(n18660), .Z(n18663) );
  XNOR U18483 ( .A(n18660), .B(n18470), .Z(n18662) );
  IV U18484 ( .A(p_input[1614]), .Z(n18470) );
  XOR U18485 ( .A(n18664), .B(n18665), .Z(n18660) );
  AND U18486 ( .A(n18666), .B(n18667), .Z(n18665) );
  XNOR U18487 ( .A(p_input[1629]), .B(n18664), .Z(n18667) );
  XNOR U18488 ( .A(n18664), .B(n18479), .Z(n18666) );
  IV U18489 ( .A(p_input[1613]), .Z(n18479) );
  XOR U18490 ( .A(n18668), .B(n18669), .Z(n18664) );
  AND U18491 ( .A(n18670), .B(n18671), .Z(n18669) );
  XNOR U18492 ( .A(p_input[1628]), .B(n18668), .Z(n18671) );
  XNOR U18493 ( .A(n18668), .B(n18488), .Z(n18670) );
  IV U18494 ( .A(p_input[1612]), .Z(n18488) );
  XOR U18495 ( .A(n18672), .B(n18673), .Z(n18668) );
  AND U18496 ( .A(n18674), .B(n18675), .Z(n18673) );
  XNOR U18497 ( .A(p_input[1627]), .B(n18672), .Z(n18675) );
  XNOR U18498 ( .A(n18672), .B(n18497), .Z(n18674) );
  IV U18499 ( .A(p_input[1611]), .Z(n18497) );
  XOR U18500 ( .A(n18676), .B(n18677), .Z(n18672) );
  AND U18501 ( .A(n18678), .B(n18679), .Z(n18677) );
  XNOR U18502 ( .A(p_input[1626]), .B(n18676), .Z(n18679) );
  XNOR U18503 ( .A(n18676), .B(n18506), .Z(n18678) );
  IV U18504 ( .A(p_input[1610]), .Z(n18506) );
  XOR U18505 ( .A(n18680), .B(n18681), .Z(n18676) );
  AND U18506 ( .A(n18682), .B(n18683), .Z(n18681) );
  XNOR U18507 ( .A(p_input[1625]), .B(n18680), .Z(n18683) );
  XNOR U18508 ( .A(n18680), .B(n18515), .Z(n18682) );
  IV U18509 ( .A(p_input[1609]), .Z(n18515) );
  XOR U18510 ( .A(n18684), .B(n18685), .Z(n18680) );
  AND U18511 ( .A(n18686), .B(n18687), .Z(n18685) );
  XNOR U18512 ( .A(p_input[1624]), .B(n18684), .Z(n18687) );
  XNOR U18513 ( .A(n18684), .B(n18524), .Z(n18686) );
  IV U18514 ( .A(p_input[1608]), .Z(n18524) );
  XOR U18515 ( .A(n18688), .B(n18689), .Z(n18684) );
  AND U18516 ( .A(n18690), .B(n18691), .Z(n18689) );
  XNOR U18517 ( .A(p_input[1623]), .B(n18688), .Z(n18691) );
  XNOR U18518 ( .A(n18688), .B(n18533), .Z(n18690) );
  IV U18519 ( .A(p_input[1607]), .Z(n18533) );
  XOR U18520 ( .A(n18692), .B(n18693), .Z(n18688) );
  AND U18521 ( .A(n18694), .B(n18695), .Z(n18693) );
  XNOR U18522 ( .A(p_input[1622]), .B(n18692), .Z(n18695) );
  XNOR U18523 ( .A(n18692), .B(n18542), .Z(n18694) );
  IV U18524 ( .A(p_input[1606]), .Z(n18542) );
  XOR U18525 ( .A(n18696), .B(n18697), .Z(n18692) );
  AND U18526 ( .A(n18698), .B(n18699), .Z(n18697) );
  XNOR U18527 ( .A(p_input[1621]), .B(n18696), .Z(n18699) );
  XNOR U18528 ( .A(n18696), .B(n18551), .Z(n18698) );
  IV U18529 ( .A(p_input[1605]), .Z(n18551) );
  XOR U18530 ( .A(n18700), .B(n18701), .Z(n18696) );
  AND U18531 ( .A(n18702), .B(n18703), .Z(n18701) );
  XNOR U18532 ( .A(p_input[1620]), .B(n18700), .Z(n18703) );
  XNOR U18533 ( .A(n18700), .B(n18560), .Z(n18702) );
  IV U18534 ( .A(p_input[1604]), .Z(n18560) );
  XOR U18535 ( .A(n18704), .B(n18705), .Z(n18700) );
  AND U18536 ( .A(n18706), .B(n18707), .Z(n18705) );
  XNOR U18537 ( .A(p_input[1619]), .B(n18704), .Z(n18707) );
  XNOR U18538 ( .A(n18704), .B(n18569), .Z(n18706) );
  IV U18539 ( .A(p_input[1603]), .Z(n18569) );
  XOR U18540 ( .A(n18708), .B(n18709), .Z(n18704) );
  AND U18541 ( .A(n18710), .B(n18711), .Z(n18709) );
  XNOR U18542 ( .A(p_input[1618]), .B(n18708), .Z(n18711) );
  XNOR U18543 ( .A(n18708), .B(n18578), .Z(n18710) );
  IV U18544 ( .A(p_input[1602]), .Z(n18578) );
  XNOR U18545 ( .A(n18712), .B(n18713), .Z(n18708) );
  AND U18546 ( .A(n18714), .B(n18715), .Z(n18713) );
  XOR U18547 ( .A(p_input[1617]), .B(n18712), .Z(n18715) );
  XNOR U18548 ( .A(p_input[1601]), .B(n18712), .Z(n18714) );
  AND U18549 ( .A(p_input[1616]), .B(n18716), .Z(n18712) );
  IV U18550 ( .A(p_input[1600]), .Z(n18716) );
  XOR U18551 ( .A(n18717), .B(n18718), .Z(n18275) );
  AND U18552 ( .A(n496), .B(n18719), .Z(n18718) );
  XNOR U18553 ( .A(n18720), .B(n18717), .Z(n18719) );
  XOR U18554 ( .A(n18721), .B(n18722), .Z(n496) );
  AND U18555 ( .A(n18723), .B(n18724), .Z(n18722) );
  XNOR U18556 ( .A(n18286), .B(n18721), .Z(n18724) );
  AND U18557 ( .A(p_input[1599]), .B(p_input[1583]), .Z(n18286) );
  XOR U18558 ( .A(n18721), .B(n18285), .Z(n18723) );
  AND U18559 ( .A(p_input[1551]), .B(p_input[1567]), .Z(n18285) );
  XOR U18560 ( .A(n18725), .B(n18726), .Z(n18721) );
  AND U18561 ( .A(n18727), .B(n18728), .Z(n18726) );
  XOR U18562 ( .A(n18725), .B(n18298), .Z(n18728) );
  XNOR U18563 ( .A(p_input[1582]), .B(n18729), .Z(n18298) );
  AND U18564 ( .A(n655), .B(n18730), .Z(n18729) );
  XOR U18565 ( .A(p_input[1598]), .B(p_input[1582]), .Z(n18730) );
  XNOR U18566 ( .A(n18295), .B(n18725), .Z(n18727) );
  XOR U18567 ( .A(n18731), .B(n18732), .Z(n18295) );
  AND U18568 ( .A(n652), .B(n18733), .Z(n18732) );
  XOR U18569 ( .A(p_input[1566]), .B(p_input[1550]), .Z(n18733) );
  XOR U18570 ( .A(n18734), .B(n18735), .Z(n18725) );
  AND U18571 ( .A(n18736), .B(n18737), .Z(n18735) );
  XOR U18572 ( .A(n18734), .B(n18310), .Z(n18737) );
  XNOR U18573 ( .A(p_input[1581]), .B(n18738), .Z(n18310) );
  AND U18574 ( .A(n655), .B(n18739), .Z(n18738) );
  XOR U18575 ( .A(p_input[1597]), .B(p_input[1581]), .Z(n18739) );
  XNOR U18576 ( .A(n18307), .B(n18734), .Z(n18736) );
  XOR U18577 ( .A(n18740), .B(n18741), .Z(n18307) );
  AND U18578 ( .A(n652), .B(n18742), .Z(n18741) );
  XOR U18579 ( .A(p_input[1565]), .B(p_input[1549]), .Z(n18742) );
  XOR U18580 ( .A(n18743), .B(n18744), .Z(n18734) );
  AND U18581 ( .A(n18745), .B(n18746), .Z(n18744) );
  XOR U18582 ( .A(n18743), .B(n18322), .Z(n18746) );
  XNOR U18583 ( .A(p_input[1580]), .B(n18747), .Z(n18322) );
  AND U18584 ( .A(n655), .B(n18748), .Z(n18747) );
  XOR U18585 ( .A(p_input[1596]), .B(p_input[1580]), .Z(n18748) );
  XNOR U18586 ( .A(n18319), .B(n18743), .Z(n18745) );
  XOR U18587 ( .A(n18749), .B(n18750), .Z(n18319) );
  AND U18588 ( .A(n652), .B(n18751), .Z(n18750) );
  XOR U18589 ( .A(p_input[1564]), .B(p_input[1548]), .Z(n18751) );
  XOR U18590 ( .A(n18752), .B(n18753), .Z(n18743) );
  AND U18591 ( .A(n18754), .B(n18755), .Z(n18753) );
  XOR U18592 ( .A(n18752), .B(n18334), .Z(n18755) );
  XNOR U18593 ( .A(p_input[1579]), .B(n18756), .Z(n18334) );
  AND U18594 ( .A(n655), .B(n18757), .Z(n18756) );
  XOR U18595 ( .A(p_input[1595]), .B(p_input[1579]), .Z(n18757) );
  XNOR U18596 ( .A(n18331), .B(n18752), .Z(n18754) );
  XOR U18597 ( .A(n18758), .B(n18759), .Z(n18331) );
  AND U18598 ( .A(n652), .B(n18760), .Z(n18759) );
  XOR U18599 ( .A(p_input[1563]), .B(p_input[1547]), .Z(n18760) );
  XOR U18600 ( .A(n18761), .B(n18762), .Z(n18752) );
  AND U18601 ( .A(n18763), .B(n18764), .Z(n18762) );
  XOR U18602 ( .A(n18761), .B(n18346), .Z(n18764) );
  XNOR U18603 ( .A(p_input[1578]), .B(n18765), .Z(n18346) );
  AND U18604 ( .A(n655), .B(n18766), .Z(n18765) );
  XOR U18605 ( .A(p_input[1594]), .B(p_input[1578]), .Z(n18766) );
  XNOR U18606 ( .A(n18343), .B(n18761), .Z(n18763) );
  XOR U18607 ( .A(n18767), .B(n18768), .Z(n18343) );
  AND U18608 ( .A(n652), .B(n18769), .Z(n18768) );
  XOR U18609 ( .A(p_input[1562]), .B(p_input[1546]), .Z(n18769) );
  XOR U18610 ( .A(n18770), .B(n18771), .Z(n18761) );
  AND U18611 ( .A(n18772), .B(n18773), .Z(n18771) );
  XOR U18612 ( .A(n18770), .B(n18358), .Z(n18773) );
  XNOR U18613 ( .A(p_input[1577]), .B(n18774), .Z(n18358) );
  AND U18614 ( .A(n655), .B(n18775), .Z(n18774) );
  XOR U18615 ( .A(p_input[1593]), .B(p_input[1577]), .Z(n18775) );
  XNOR U18616 ( .A(n18355), .B(n18770), .Z(n18772) );
  XOR U18617 ( .A(n18776), .B(n18777), .Z(n18355) );
  AND U18618 ( .A(n652), .B(n18778), .Z(n18777) );
  XOR U18619 ( .A(p_input[1561]), .B(p_input[1545]), .Z(n18778) );
  XOR U18620 ( .A(n18779), .B(n18780), .Z(n18770) );
  AND U18621 ( .A(n18781), .B(n18782), .Z(n18780) );
  XOR U18622 ( .A(n18779), .B(n18370), .Z(n18782) );
  XNOR U18623 ( .A(p_input[1576]), .B(n18783), .Z(n18370) );
  AND U18624 ( .A(n655), .B(n18784), .Z(n18783) );
  XOR U18625 ( .A(p_input[1592]), .B(p_input[1576]), .Z(n18784) );
  XNOR U18626 ( .A(n18367), .B(n18779), .Z(n18781) );
  XOR U18627 ( .A(n18785), .B(n18786), .Z(n18367) );
  AND U18628 ( .A(n652), .B(n18787), .Z(n18786) );
  XOR U18629 ( .A(p_input[1560]), .B(p_input[1544]), .Z(n18787) );
  XOR U18630 ( .A(n18788), .B(n18789), .Z(n18779) );
  AND U18631 ( .A(n18790), .B(n18791), .Z(n18789) );
  XOR U18632 ( .A(n18788), .B(n18382), .Z(n18791) );
  XNOR U18633 ( .A(p_input[1575]), .B(n18792), .Z(n18382) );
  AND U18634 ( .A(n655), .B(n18793), .Z(n18792) );
  XOR U18635 ( .A(p_input[1591]), .B(p_input[1575]), .Z(n18793) );
  XNOR U18636 ( .A(n18379), .B(n18788), .Z(n18790) );
  XOR U18637 ( .A(n18794), .B(n18795), .Z(n18379) );
  AND U18638 ( .A(n652), .B(n18796), .Z(n18795) );
  XOR U18639 ( .A(p_input[1559]), .B(p_input[1543]), .Z(n18796) );
  XOR U18640 ( .A(n18797), .B(n18798), .Z(n18788) );
  AND U18641 ( .A(n18799), .B(n18800), .Z(n18798) );
  XOR U18642 ( .A(n18797), .B(n18394), .Z(n18800) );
  XNOR U18643 ( .A(p_input[1574]), .B(n18801), .Z(n18394) );
  AND U18644 ( .A(n655), .B(n18802), .Z(n18801) );
  XOR U18645 ( .A(p_input[1590]), .B(p_input[1574]), .Z(n18802) );
  XNOR U18646 ( .A(n18391), .B(n18797), .Z(n18799) );
  XOR U18647 ( .A(n18803), .B(n18804), .Z(n18391) );
  AND U18648 ( .A(n652), .B(n18805), .Z(n18804) );
  XOR U18649 ( .A(p_input[1558]), .B(p_input[1542]), .Z(n18805) );
  XOR U18650 ( .A(n18806), .B(n18807), .Z(n18797) );
  AND U18651 ( .A(n18808), .B(n18809), .Z(n18807) );
  XOR U18652 ( .A(n18806), .B(n18406), .Z(n18809) );
  XNOR U18653 ( .A(p_input[1573]), .B(n18810), .Z(n18406) );
  AND U18654 ( .A(n655), .B(n18811), .Z(n18810) );
  XOR U18655 ( .A(p_input[1589]), .B(p_input[1573]), .Z(n18811) );
  XNOR U18656 ( .A(n18403), .B(n18806), .Z(n18808) );
  XOR U18657 ( .A(n18812), .B(n18813), .Z(n18403) );
  AND U18658 ( .A(n652), .B(n18814), .Z(n18813) );
  XOR U18659 ( .A(p_input[1557]), .B(p_input[1541]), .Z(n18814) );
  XOR U18660 ( .A(n18815), .B(n18816), .Z(n18806) );
  AND U18661 ( .A(n18817), .B(n18818), .Z(n18816) );
  XOR U18662 ( .A(n18815), .B(n18418), .Z(n18818) );
  XNOR U18663 ( .A(p_input[1572]), .B(n18819), .Z(n18418) );
  AND U18664 ( .A(n655), .B(n18820), .Z(n18819) );
  XOR U18665 ( .A(p_input[1588]), .B(p_input[1572]), .Z(n18820) );
  XNOR U18666 ( .A(n18415), .B(n18815), .Z(n18817) );
  XOR U18667 ( .A(n18821), .B(n18822), .Z(n18415) );
  AND U18668 ( .A(n652), .B(n18823), .Z(n18822) );
  XOR U18669 ( .A(p_input[1556]), .B(p_input[1540]), .Z(n18823) );
  XOR U18670 ( .A(n18824), .B(n18825), .Z(n18815) );
  AND U18671 ( .A(n18826), .B(n18827), .Z(n18825) );
  XOR U18672 ( .A(n18824), .B(n18430), .Z(n18827) );
  XNOR U18673 ( .A(p_input[1571]), .B(n18828), .Z(n18430) );
  AND U18674 ( .A(n655), .B(n18829), .Z(n18828) );
  XOR U18675 ( .A(p_input[1587]), .B(p_input[1571]), .Z(n18829) );
  XNOR U18676 ( .A(n18427), .B(n18824), .Z(n18826) );
  XOR U18677 ( .A(n18830), .B(n18831), .Z(n18427) );
  AND U18678 ( .A(n652), .B(n18832), .Z(n18831) );
  XOR U18679 ( .A(p_input[1555]), .B(p_input[1539]), .Z(n18832) );
  XOR U18680 ( .A(n18833), .B(n18834), .Z(n18824) );
  AND U18681 ( .A(n18835), .B(n18836), .Z(n18834) );
  XOR U18682 ( .A(n18833), .B(n18442), .Z(n18836) );
  XNOR U18683 ( .A(p_input[1570]), .B(n18837), .Z(n18442) );
  AND U18684 ( .A(n655), .B(n18838), .Z(n18837) );
  XOR U18685 ( .A(p_input[1586]), .B(p_input[1570]), .Z(n18838) );
  XNOR U18686 ( .A(n18439), .B(n18833), .Z(n18835) );
  XOR U18687 ( .A(n18839), .B(n18840), .Z(n18439) );
  AND U18688 ( .A(n652), .B(n18841), .Z(n18840) );
  XOR U18689 ( .A(p_input[1554]), .B(p_input[1538]), .Z(n18841) );
  XOR U18690 ( .A(n18842), .B(n18843), .Z(n18833) );
  AND U18691 ( .A(n18844), .B(n18845), .Z(n18843) );
  XNOR U18692 ( .A(n18846), .B(n18455), .Z(n18845) );
  XNOR U18693 ( .A(p_input[1569]), .B(n18847), .Z(n18455) );
  AND U18694 ( .A(n655), .B(n18848), .Z(n18847) );
  XNOR U18695 ( .A(p_input[1585]), .B(n18849), .Z(n18848) );
  IV U18696 ( .A(p_input[1569]), .Z(n18849) );
  XNOR U18697 ( .A(n18452), .B(n18842), .Z(n18844) );
  XNOR U18698 ( .A(p_input[1537]), .B(n18850), .Z(n18452) );
  AND U18699 ( .A(n652), .B(n18851), .Z(n18850) );
  XOR U18700 ( .A(p_input[1553]), .B(p_input[1537]), .Z(n18851) );
  IV U18701 ( .A(n18846), .Z(n18842) );
  AND U18702 ( .A(n18717), .B(n18720), .Z(n18846) );
  XOR U18703 ( .A(p_input[1568]), .B(n18852), .Z(n18720) );
  AND U18704 ( .A(n655), .B(n18853), .Z(n18852) );
  XOR U18705 ( .A(p_input[1584]), .B(p_input[1568]), .Z(n18853) );
  XOR U18706 ( .A(n18854), .B(n18855), .Z(n655) );
  AND U18707 ( .A(n18856), .B(n18857), .Z(n18855) );
  XNOR U18708 ( .A(p_input[1599]), .B(n18854), .Z(n18857) );
  XOR U18709 ( .A(n18854), .B(p_input[1583]), .Z(n18856) );
  XOR U18710 ( .A(n18858), .B(n18859), .Z(n18854) );
  AND U18711 ( .A(n18860), .B(n18861), .Z(n18859) );
  XNOR U18712 ( .A(p_input[1598]), .B(n18858), .Z(n18861) );
  XOR U18713 ( .A(n18858), .B(p_input[1582]), .Z(n18860) );
  XOR U18714 ( .A(n18862), .B(n18863), .Z(n18858) );
  AND U18715 ( .A(n18864), .B(n18865), .Z(n18863) );
  XNOR U18716 ( .A(p_input[1597]), .B(n18862), .Z(n18865) );
  XOR U18717 ( .A(n18862), .B(p_input[1581]), .Z(n18864) );
  XOR U18718 ( .A(n18866), .B(n18867), .Z(n18862) );
  AND U18719 ( .A(n18868), .B(n18869), .Z(n18867) );
  XNOR U18720 ( .A(p_input[1596]), .B(n18866), .Z(n18869) );
  XOR U18721 ( .A(n18866), .B(p_input[1580]), .Z(n18868) );
  XOR U18722 ( .A(n18870), .B(n18871), .Z(n18866) );
  AND U18723 ( .A(n18872), .B(n18873), .Z(n18871) );
  XNOR U18724 ( .A(p_input[1595]), .B(n18870), .Z(n18873) );
  XOR U18725 ( .A(n18870), .B(p_input[1579]), .Z(n18872) );
  XOR U18726 ( .A(n18874), .B(n18875), .Z(n18870) );
  AND U18727 ( .A(n18876), .B(n18877), .Z(n18875) );
  XNOR U18728 ( .A(p_input[1594]), .B(n18874), .Z(n18877) );
  XOR U18729 ( .A(n18874), .B(p_input[1578]), .Z(n18876) );
  XOR U18730 ( .A(n18878), .B(n18879), .Z(n18874) );
  AND U18731 ( .A(n18880), .B(n18881), .Z(n18879) );
  XNOR U18732 ( .A(p_input[1593]), .B(n18878), .Z(n18881) );
  XOR U18733 ( .A(n18878), .B(p_input[1577]), .Z(n18880) );
  XOR U18734 ( .A(n18882), .B(n18883), .Z(n18878) );
  AND U18735 ( .A(n18884), .B(n18885), .Z(n18883) );
  XNOR U18736 ( .A(p_input[1592]), .B(n18882), .Z(n18885) );
  XOR U18737 ( .A(n18882), .B(p_input[1576]), .Z(n18884) );
  XOR U18738 ( .A(n18886), .B(n18887), .Z(n18882) );
  AND U18739 ( .A(n18888), .B(n18889), .Z(n18887) );
  XNOR U18740 ( .A(p_input[1591]), .B(n18886), .Z(n18889) );
  XOR U18741 ( .A(n18886), .B(p_input[1575]), .Z(n18888) );
  XOR U18742 ( .A(n18890), .B(n18891), .Z(n18886) );
  AND U18743 ( .A(n18892), .B(n18893), .Z(n18891) );
  XNOR U18744 ( .A(p_input[1590]), .B(n18890), .Z(n18893) );
  XOR U18745 ( .A(n18890), .B(p_input[1574]), .Z(n18892) );
  XOR U18746 ( .A(n18894), .B(n18895), .Z(n18890) );
  AND U18747 ( .A(n18896), .B(n18897), .Z(n18895) );
  XNOR U18748 ( .A(p_input[1589]), .B(n18894), .Z(n18897) );
  XOR U18749 ( .A(n18894), .B(p_input[1573]), .Z(n18896) );
  XOR U18750 ( .A(n18898), .B(n18899), .Z(n18894) );
  AND U18751 ( .A(n18900), .B(n18901), .Z(n18899) );
  XNOR U18752 ( .A(p_input[1588]), .B(n18898), .Z(n18901) );
  XOR U18753 ( .A(n18898), .B(p_input[1572]), .Z(n18900) );
  XOR U18754 ( .A(n18902), .B(n18903), .Z(n18898) );
  AND U18755 ( .A(n18904), .B(n18905), .Z(n18903) );
  XNOR U18756 ( .A(p_input[1587]), .B(n18902), .Z(n18905) );
  XOR U18757 ( .A(n18902), .B(p_input[1571]), .Z(n18904) );
  XOR U18758 ( .A(n18906), .B(n18907), .Z(n18902) );
  AND U18759 ( .A(n18908), .B(n18909), .Z(n18907) );
  XNOR U18760 ( .A(p_input[1586]), .B(n18906), .Z(n18909) );
  XOR U18761 ( .A(n18906), .B(p_input[1570]), .Z(n18908) );
  XNOR U18762 ( .A(n18910), .B(n18911), .Z(n18906) );
  AND U18763 ( .A(n18912), .B(n18913), .Z(n18911) );
  XOR U18764 ( .A(p_input[1585]), .B(n18910), .Z(n18913) );
  XNOR U18765 ( .A(p_input[1569]), .B(n18910), .Z(n18912) );
  AND U18766 ( .A(p_input[1584]), .B(n18914), .Z(n18910) );
  IV U18767 ( .A(p_input[1568]), .Z(n18914) );
  XNOR U18768 ( .A(p_input[1536]), .B(n18915), .Z(n18717) );
  AND U18769 ( .A(n652), .B(n18916), .Z(n18915) );
  XOR U18770 ( .A(p_input[1552]), .B(p_input[1536]), .Z(n18916) );
  XOR U18771 ( .A(n18917), .B(n18918), .Z(n652) );
  AND U18772 ( .A(n18919), .B(n18920), .Z(n18918) );
  XNOR U18773 ( .A(p_input[1567]), .B(n18917), .Z(n18920) );
  XOR U18774 ( .A(n18917), .B(p_input[1551]), .Z(n18919) );
  XOR U18775 ( .A(n18921), .B(n18922), .Z(n18917) );
  AND U18776 ( .A(n18923), .B(n18924), .Z(n18922) );
  XNOR U18777 ( .A(p_input[1566]), .B(n18921), .Z(n18924) );
  XNOR U18778 ( .A(n18921), .B(n18731), .Z(n18923) );
  IV U18779 ( .A(p_input[1550]), .Z(n18731) );
  XOR U18780 ( .A(n18925), .B(n18926), .Z(n18921) );
  AND U18781 ( .A(n18927), .B(n18928), .Z(n18926) );
  XNOR U18782 ( .A(p_input[1565]), .B(n18925), .Z(n18928) );
  XNOR U18783 ( .A(n18925), .B(n18740), .Z(n18927) );
  IV U18784 ( .A(p_input[1549]), .Z(n18740) );
  XOR U18785 ( .A(n18929), .B(n18930), .Z(n18925) );
  AND U18786 ( .A(n18931), .B(n18932), .Z(n18930) );
  XNOR U18787 ( .A(p_input[1564]), .B(n18929), .Z(n18932) );
  XNOR U18788 ( .A(n18929), .B(n18749), .Z(n18931) );
  IV U18789 ( .A(p_input[1548]), .Z(n18749) );
  XOR U18790 ( .A(n18933), .B(n18934), .Z(n18929) );
  AND U18791 ( .A(n18935), .B(n18936), .Z(n18934) );
  XNOR U18792 ( .A(p_input[1563]), .B(n18933), .Z(n18936) );
  XNOR U18793 ( .A(n18933), .B(n18758), .Z(n18935) );
  IV U18794 ( .A(p_input[1547]), .Z(n18758) );
  XOR U18795 ( .A(n18937), .B(n18938), .Z(n18933) );
  AND U18796 ( .A(n18939), .B(n18940), .Z(n18938) );
  XNOR U18797 ( .A(p_input[1562]), .B(n18937), .Z(n18940) );
  XNOR U18798 ( .A(n18937), .B(n18767), .Z(n18939) );
  IV U18799 ( .A(p_input[1546]), .Z(n18767) );
  XOR U18800 ( .A(n18941), .B(n18942), .Z(n18937) );
  AND U18801 ( .A(n18943), .B(n18944), .Z(n18942) );
  XNOR U18802 ( .A(p_input[1561]), .B(n18941), .Z(n18944) );
  XNOR U18803 ( .A(n18941), .B(n18776), .Z(n18943) );
  IV U18804 ( .A(p_input[1545]), .Z(n18776) );
  XOR U18805 ( .A(n18945), .B(n18946), .Z(n18941) );
  AND U18806 ( .A(n18947), .B(n18948), .Z(n18946) );
  XNOR U18807 ( .A(p_input[1560]), .B(n18945), .Z(n18948) );
  XNOR U18808 ( .A(n18945), .B(n18785), .Z(n18947) );
  IV U18809 ( .A(p_input[1544]), .Z(n18785) );
  XOR U18810 ( .A(n18949), .B(n18950), .Z(n18945) );
  AND U18811 ( .A(n18951), .B(n18952), .Z(n18950) );
  XNOR U18812 ( .A(p_input[1559]), .B(n18949), .Z(n18952) );
  XNOR U18813 ( .A(n18949), .B(n18794), .Z(n18951) );
  IV U18814 ( .A(p_input[1543]), .Z(n18794) );
  XOR U18815 ( .A(n18953), .B(n18954), .Z(n18949) );
  AND U18816 ( .A(n18955), .B(n18956), .Z(n18954) );
  XNOR U18817 ( .A(p_input[1558]), .B(n18953), .Z(n18956) );
  XNOR U18818 ( .A(n18953), .B(n18803), .Z(n18955) );
  IV U18819 ( .A(p_input[1542]), .Z(n18803) );
  XOR U18820 ( .A(n18957), .B(n18958), .Z(n18953) );
  AND U18821 ( .A(n18959), .B(n18960), .Z(n18958) );
  XNOR U18822 ( .A(p_input[1557]), .B(n18957), .Z(n18960) );
  XNOR U18823 ( .A(n18957), .B(n18812), .Z(n18959) );
  IV U18824 ( .A(p_input[1541]), .Z(n18812) );
  XOR U18825 ( .A(n18961), .B(n18962), .Z(n18957) );
  AND U18826 ( .A(n18963), .B(n18964), .Z(n18962) );
  XNOR U18827 ( .A(p_input[1556]), .B(n18961), .Z(n18964) );
  XNOR U18828 ( .A(n18961), .B(n18821), .Z(n18963) );
  IV U18829 ( .A(p_input[1540]), .Z(n18821) );
  XOR U18830 ( .A(n18965), .B(n18966), .Z(n18961) );
  AND U18831 ( .A(n18967), .B(n18968), .Z(n18966) );
  XNOR U18832 ( .A(p_input[1555]), .B(n18965), .Z(n18968) );
  XNOR U18833 ( .A(n18965), .B(n18830), .Z(n18967) );
  IV U18834 ( .A(p_input[1539]), .Z(n18830) );
  XOR U18835 ( .A(n18969), .B(n18970), .Z(n18965) );
  AND U18836 ( .A(n18971), .B(n18972), .Z(n18970) );
  XNOR U18837 ( .A(p_input[1554]), .B(n18969), .Z(n18972) );
  XNOR U18838 ( .A(n18969), .B(n18839), .Z(n18971) );
  IV U18839 ( .A(p_input[1538]), .Z(n18839) );
  XNOR U18840 ( .A(n18973), .B(n18974), .Z(n18969) );
  AND U18841 ( .A(n18975), .B(n18976), .Z(n18974) );
  XOR U18842 ( .A(p_input[1553]), .B(n18973), .Z(n18976) );
  XNOR U18843 ( .A(p_input[1537]), .B(n18973), .Z(n18975) );
  AND U18844 ( .A(p_input[1552]), .B(n18977), .Z(n18973) );
  IV U18845 ( .A(p_input[1536]), .Z(n18977) );
  XOR U18846 ( .A(n18978), .B(n18979), .Z(n15432) );
  AND U18847 ( .A(n1017), .B(n18980), .Z(n18979) );
  XNOR U18848 ( .A(n18981), .B(n18978), .Z(n18980) );
  XOR U18849 ( .A(n18982), .B(n18983), .Z(n1017) );
  AND U18850 ( .A(n18984), .B(n18985), .Z(n18983) );
  XOR U18851 ( .A(n18982), .B(n15447), .Z(n18985) );
  XNOR U18852 ( .A(n18986), .B(n18987), .Z(n15447) );
  AND U18853 ( .A(n18988), .B(n951), .Z(n18987) );
  AND U18854 ( .A(n18986), .B(n18989), .Z(n18988) );
  XNOR U18855 ( .A(n15444), .B(n18982), .Z(n18984) );
  XOR U18856 ( .A(n18990), .B(n18991), .Z(n15444) );
  AND U18857 ( .A(n18992), .B(n948), .Z(n18991) );
  NOR U18858 ( .A(n18990), .B(n18993), .Z(n18992) );
  XOR U18859 ( .A(n18994), .B(n18995), .Z(n18982) );
  AND U18860 ( .A(n18996), .B(n18997), .Z(n18995) );
  XOR U18861 ( .A(n18994), .B(n15459), .Z(n18997) );
  XOR U18862 ( .A(n18998), .B(n18999), .Z(n15459) );
  AND U18863 ( .A(n951), .B(n19000), .Z(n18999) );
  XOR U18864 ( .A(n19001), .B(n18998), .Z(n19000) );
  XNOR U18865 ( .A(n15456), .B(n18994), .Z(n18996) );
  XOR U18866 ( .A(n19002), .B(n19003), .Z(n15456) );
  AND U18867 ( .A(n948), .B(n19004), .Z(n19003) );
  XOR U18868 ( .A(n19005), .B(n19002), .Z(n19004) );
  XOR U18869 ( .A(n19006), .B(n19007), .Z(n18994) );
  AND U18870 ( .A(n19008), .B(n19009), .Z(n19007) );
  XOR U18871 ( .A(n19006), .B(n15471), .Z(n19009) );
  XOR U18872 ( .A(n19010), .B(n19011), .Z(n15471) );
  AND U18873 ( .A(n951), .B(n19012), .Z(n19011) );
  XOR U18874 ( .A(n19013), .B(n19010), .Z(n19012) );
  XNOR U18875 ( .A(n15468), .B(n19006), .Z(n19008) );
  XOR U18876 ( .A(n19014), .B(n19015), .Z(n15468) );
  AND U18877 ( .A(n948), .B(n19016), .Z(n19015) );
  XOR U18878 ( .A(n19017), .B(n19014), .Z(n19016) );
  XOR U18879 ( .A(n19018), .B(n19019), .Z(n19006) );
  AND U18880 ( .A(n19020), .B(n19021), .Z(n19019) );
  XOR U18881 ( .A(n19018), .B(n15483), .Z(n19021) );
  XOR U18882 ( .A(n19022), .B(n19023), .Z(n15483) );
  AND U18883 ( .A(n951), .B(n19024), .Z(n19023) );
  XOR U18884 ( .A(n19025), .B(n19022), .Z(n19024) );
  XNOR U18885 ( .A(n15480), .B(n19018), .Z(n19020) );
  XOR U18886 ( .A(n19026), .B(n19027), .Z(n15480) );
  AND U18887 ( .A(n948), .B(n19028), .Z(n19027) );
  XOR U18888 ( .A(n19029), .B(n19026), .Z(n19028) );
  XOR U18889 ( .A(n19030), .B(n19031), .Z(n19018) );
  AND U18890 ( .A(n19032), .B(n19033), .Z(n19031) );
  XOR U18891 ( .A(n19030), .B(n15495), .Z(n19033) );
  XOR U18892 ( .A(n19034), .B(n19035), .Z(n15495) );
  AND U18893 ( .A(n951), .B(n19036), .Z(n19035) );
  XOR U18894 ( .A(n19037), .B(n19034), .Z(n19036) );
  XNOR U18895 ( .A(n15492), .B(n19030), .Z(n19032) );
  XOR U18896 ( .A(n19038), .B(n19039), .Z(n15492) );
  AND U18897 ( .A(n948), .B(n19040), .Z(n19039) );
  XOR U18898 ( .A(n19041), .B(n19038), .Z(n19040) );
  XOR U18899 ( .A(n19042), .B(n19043), .Z(n19030) );
  AND U18900 ( .A(n19044), .B(n19045), .Z(n19043) );
  XOR U18901 ( .A(n19042), .B(n15507), .Z(n19045) );
  XOR U18902 ( .A(n19046), .B(n19047), .Z(n15507) );
  AND U18903 ( .A(n951), .B(n19048), .Z(n19047) );
  XOR U18904 ( .A(n19049), .B(n19046), .Z(n19048) );
  XNOR U18905 ( .A(n15504), .B(n19042), .Z(n19044) );
  XOR U18906 ( .A(n19050), .B(n19051), .Z(n15504) );
  AND U18907 ( .A(n948), .B(n19052), .Z(n19051) );
  XOR U18908 ( .A(n19053), .B(n19050), .Z(n19052) );
  XOR U18909 ( .A(n19054), .B(n19055), .Z(n19042) );
  AND U18910 ( .A(n19056), .B(n19057), .Z(n19055) );
  XOR U18911 ( .A(n19054), .B(n15519), .Z(n19057) );
  XOR U18912 ( .A(n19058), .B(n19059), .Z(n15519) );
  AND U18913 ( .A(n951), .B(n19060), .Z(n19059) );
  XOR U18914 ( .A(n19061), .B(n19058), .Z(n19060) );
  XNOR U18915 ( .A(n15516), .B(n19054), .Z(n19056) );
  XOR U18916 ( .A(n19062), .B(n19063), .Z(n15516) );
  AND U18917 ( .A(n948), .B(n19064), .Z(n19063) );
  XOR U18918 ( .A(n19065), .B(n19062), .Z(n19064) );
  XOR U18919 ( .A(n19066), .B(n19067), .Z(n19054) );
  AND U18920 ( .A(n19068), .B(n19069), .Z(n19067) );
  XOR U18921 ( .A(n19066), .B(n15531), .Z(n19069) );
  XOR U18922 ( .A(n19070), .B(n19071), .Z(n15531) );
  AND U18923 ( .A(n951), .B(n19072), .Z(n19071) );
  XOR U18924 ( .A(n19073), .B(n19070), .Z(n19072) );
  XNOR U18925 ( .A(n15528), .B(n19066), .Z(n19068) );
  XOR U18926 ( .A(n19074), .B(n19075), .Z(n15528) );
  AND U18927 ( .A(n948), .B(n19076), .Z(n19075) );
  XOR U18928 ( .A(n19077), .B(n19074), .Z(n19076) );
  XOR U18929 ( .A(n19078), .B(n19079), .Z(n19066) );
  AND U18930 ( .A(n19080), .B(n19081), .Z(n19079) );
  XOR U18931 ( .A(n19078), .B(n15543), .Z(n19081) );
  XOR U18932 ( .A(n19082), .B(n19083), .Z(n15543) );
  AND U18933 ( .A(n951), .B(n19084), .Z(n19083) );
  XOR U18934 ( .A(n19085), .B(n19082), .Z(n19084) );
  XNOR U18935 ( .A(n15540), .B(n19078), .Z(n19080) );
  XOR U18936 ( .A(n19086), .B(n19087), .Z(n15540) );
  AND U18937 ( .A(n948), .B(n19088), .Z(n19087) );
  XOR U18938 ( .A(n19089), .B(n19086), .Z(n19088) );
  XOR U18939 ( .A(n19090), .B(n19091), .Z(n19078) );
  AND U18940 ( .A(n19092), .B(n19093), .Z(n19091) );
  XOR U18941 ( .A(n19090), .B(n15555), .Z(n19093) );
  XOR U18942 ( .A(n19094), .B(n19095), .Z(n15555) );
  AND U18943 ( .A(n951), .B(n19096), .Z(n19095) );
  XOR U18944 ( .A(n19097), .B(n19094), .Z(n19096) );
  XNOR U18945 ( .A(n15552), .B(n19090), .Z(n19092) );
  XOR U18946 ( .A(n19098), .B(n19099), .Z(n15552) );
  AND U18947 ( .A(n948), .B(n19100), .Z(n19099) );
  XOR U18948 ( .A(n19101), .B(n19098), .Z(n19100) );
  XOR U18949 ( .A(n19102), .B(n19103), .Z(n19090) );
  AND U18950 ( .A(n19104), .B(n19105), .Z(n19103) );
  XOR U18951 ( .A(n19102), .B(n15567), .Z(n19105) );
  XOR U18952 ( .A(n19106), .B(n19107), .Z(n15567) );
  AND U18953 ( .A(n951), .B(n19108), .Z(n19107) );
  XOR U18954 ( .A(n19109), .B(n19106), .Z(n19108) );
  XNOR U18955 ( .A(n15564), .B(n19102), .Z(n19104) );
  XOR U18956 ( .A(n19110), .B(n19111), .Z(n15564) );
  AND U18957 ( .A(n948), .B(n19112), .Z(n19111) );
  XOR U18958 ( .A(n19113), .B(n19110), .Z(n19112) );
  XOR U18959 ( .A(n19114), .B(n19115), .Z(n19102) );
  AND U18960 ( .A(n19116), .B(n19117), .Z(n19115) );
  XOR U18961 ( .A(n19114), .B(n15579), .Z(n19117) );
  XOR U18962 ( .A(n19118), .B(n19119), .Z(n15579) );
  AND U18963 ( .A(n951), .B(n19120), .Z(n19119) );
  XOR U18964 ( .A(n19121), .B(n19118), .Z(n19120) );
  XNOR U18965 ( .A(n15576), .B(n19114), .Z(n19116) );
  XOR U18966 ( .A(n19122), .B(n19123), .Z(n15576) );
  AND U18967 ( .A(n948), .B(n19124), .Z(n19123) );
  XOR U18968 ( .A(n19125), .B(n19122), .Z(n19124) );
  XOR U18969 ( .A(n19126), .B(n19127), .Z(n19114) );
  AND U18970 ( .A(n19128), .B(n19129), .Z(n19127) );
  XOR U18971 ( .A(n19126), .B(n15591), .Z(n19129) );
  XOR U18972 ( .A(n19130), .B(n19131), .Z(n15591) );
  AND U18973 ( .A(n951), .B(n19132), .Z(n19131) );
  XOR U18974 ( .A(n19133), .B(n19130), .Z(n19132) );
  XNOR U18975 ( .A(n15588), .B(n19126), .Z(n19128) );
  XOR U18976 ( .A(n19134), .B(n19135), .Z(n15588) );
  AND U18977 ( .A(n948), .B(n19136), .Z(n19135) );
  XOR U18978 ( .A(n19137), .B(n19134), .Z(n19136) );
  XOR U18979 ( .A(n19138), .B(n19139), .Z(n19126) );
  AND U18980 ( .A(n19140), .B(n19141), .Z(n19139) );
  XOR U18981 ( .A(n19138), .B(n15603), .Z(n19141) );
  XOR U18982 ( .A(n19142), .B(n19143), .Z(n15603) );
  AND U18983 ( .A(n951), .B(n19144), .Z(n19143) );
  XOR U18984 ( .A(n19145), .B(n19142), .Z(n19144) );
  XNOR U18985 ( .A(n15600), .B(n19138), .Z(n19140) );
  XOR U18986 ( .A(n19146), .B(n19147), .Z(n15600) );
  AND U18987 ( .A(n948), .B(n19148), .Z(n19147) );
  XOR U18988 ( .A(n19149), .B(n19146), .Z(n19148) );
  XOR U18989 ( .A(n19150), .B(n19151), .Z(n19138) );
  AND U18990 ( .A(n19152), .B(n19153), .Z(n19151) );
  XNOR U18991 ( .A(n19154), .B(n15616), .Z(n19153) );
  XOR U18992 ( .A(n19155), .B(n19156), .Z(n15616) );
  AND U18993 ( .A(n951), .B(n19157), .Z(n19156) );
  XOR U18994 ( .A(n19155), .B(n19158), .Z(n19157) );
  XNOR U18995 ( .A(n15613), .B(n19150), .Z(n19152) );
  XOR U18996 ( .A(n19159), .B(n19160), .Z(n15613) );
  AND U18997 ( .A(n948), .B(n19161), .Z(n19160) );
  XOR U18998 ( .A(n19159), .B(n19162), .Z(n19161) );
  IV U18999 ( .A(n19154), .Z(n19150) );
  AND U19000 ( .A(n18978), .B(n18981), .Z(n19154) );
  XNOR U19001 ( .A(n19163), .B(n19164), .Z(n18981) );
  AND U19002 ( .A(n951), .B(n19165), .Z(n19164) );
  XNOR U19003 ( .A(n19166), .B(n19163), .Z(n19165) );
  XOR U19004 ( .A(n19167), .B(n19168), .Z(n951) );
  AND U19005 ( .A(n19169), .B(n19170), .Z(n19168) );
  XOR U19006 ( .A(n18989), .B(n19167), .Z(n19170) );
  IV U19007 ( .A(n19171), .Z(n18989) );
  AND U19008 ( .A(n19172), .B(n19173), .Z(n19171) );
  XOR U19009 ( .A(n19167), .B(n18986), .Z(n19169) );
  AND U19010 ( .A(n19174), .B(n19175), .Z(n18986) );
  XOR U19011 ( .A(n19176), .B(n19177), .Z(n19167) );
  AND U19012 ( .A(n19178), .B(n19179), .Z(n19177) );
  XOR U19013 ( .A(n19176), .B(n19001), .Z(n19179) );
  XOR U19014 ( .A(n19180), .B(n19181), .Z(n19001) );
  AND U19015 ( .A(n807), .B(n19182), .Z(n19181) );
  XOR U19016 ( .A(n19183), .B(n19180), .Z(n19182) );
  XNOR U19017 ( .A(n18998), .B(n19176), .Z(n19178) );
  XOR U19018 ( .A(n19184), .B(n19185), .Z(n18998) );
  AND U19019 ( .A(n805), .B(n19186), .Z(n19185) );
  XOR U19020 ( .A(n19187), .B(n19184), .Z(n19186) );
  XOR U19021 ( .A(n19188), .B(n19189), .Z(n19176) );
  AND U19022 ( .A(n19190), .B(n19191), .Z(n19189) );
  XOR U19023 ( .A(n19188), .B(n19013), .Z(n19191) );
  XOR U19024 ( .A(n19192), .B(n19193), .Z(n19013) );
  AND U19025 ( .A(n807), .B(n19194), .Z(n19193) );
  XOR U19026 ( .A(n19195), .B(n19192), .Z(n19194) );
  XNOR U19027 ( .A(n19010), .B(n19188), .Z(n19190) );
  XOR U19028 ( .A(n19196), .B(n19197), .Z(n19010) );
  AND U19029 ( .A(n805), .B(n19198), .Z(n19197) );
  XOR U19030 ( .A(n19199), .B(n19196), .Z(n19198) );
  XOR U19031 ( .A(n19200), .B(n19201), .Z(n19188) );
  AND U19032 ( .A(n19202), .B(n19203), .Z(n19201) );
  XOR U19033 ( .A(n19200), .B(n19025), .Z(n19203) );
  XOR U19034 ( .A(n19204), .B(n19205), .Z(n19025) );
  AND U19035 ( .A(n807), .B(n19206), .Z(n19205) );
  XOR U19036 ( .A(n19207), .B(n19204), .Z(n19206) );
  XNOR U19037 ( .A(n19022), .B(n19200), .Z(n19202) );
  XOR U19038 ( .A(n19208), .B(n19209), .Z(n19022) );
  AND U19039 ( .A(n805), .B(n19210), .Z(n19209) );
  XOR U19040 ( .A(n19211), .B(n19208), .Z(n19210) );
  XOR U19041 ( .A(n19212), .B(n19213), .Z(n19200) );
  AND U19042 ( .A(n19214), .B(n19215), .Z(n19213) );
  XOR U19043 ( .A(n19212), .B(n19037), .Z(n19215) );
  XOR U19044 ( .A(n19216), .B(n19217), .Z(n19037) );
  AND U19045 ( .A(n807), .B(n19218), .Z(n19217) );
  XOR U19046 ( .A(n19219), .B(n19216), .Z(n19218) );
  XNOR U19047 ( .A(n19034), .B(n19212), .Z(n19214) );
  XOR U19048 ( .A(n19220), .B(n19221), .Z(n19034) );
  AND U19049 ( .A(n805), .B(n19222), .Z(n19221) );
  XOR U19050 ( .A(n19223), .B(n19220), .Z(n19222) );
  XOR U19051 ( .A(n19224), .B(n19225), .Z(n19212) );
  AND U19052 ( .A(n19226), .B(n19227), .Z(n19225) );
  XOR U19053 ( .A(n19224), .B(n19049), .Z(n19227) );
  XOR U19054 ( .A(n19228), .B(n19229), .Z(n19049) );
  AND U19055 ( .A(n807), .B(n19230), .Z(n19229) );
  XOR U19056 ( .A(n19231), .B(n19228), .Z(n19230) );
  XNOR U19057 ( .A(n19046), .B(n19224), .Z(n19226) );
  XOR U19058 ( .A(n19232), .B(n19233), .Z(n19046) );
  AND U19059 ( .A(n805), .B(n19234), .Z(n19233) );
  XOR U19060 ( .A(n19235), .B(n19232), .Z(n19234) );
  XOR U19061 ( .A(n19236), .B(n19237), .Z(n19224) );
  AND U19062 ( .A(n19238), .B(n19239), .Z(n19237) );
  XOR U19063 ( .A(n19236), .B(n19061), .Z(n19239) );
  XOR U19064 ( .A(n19240), .B(n19241), .Z(n19061) );
  AND U19065 ( .A(n807), .B(n19242), .Z(n19241) );
  XOR U19066 ( .A(n19243), .B(n19240), .Z(n19242) );
  XNOR U19067 ( .A(n19058), .B(n19236), .Z(n19238) );
  XOR U19068 ( .A(n19244), .B(n19245), .Z(n19058) );
  AND U19069 ( .A(n805), .B(n19246), .Z(n19245) );
  XOR U19070 ( .A(n19247), .B(n19244), .Z(n19246) );
  XOR U19071 ( .A(n19248), .B(n19249), .Z(n19236) );
  AND U19072 ( .A(n19250), .B(n19251), .Z(n19249) );
  XOR U19073 ( .A(n19248), .B(n19073), .Z(n19251) );
  XOR U19074 ( .A(n19252), .B(n19253), .Z(n19073) );
  AND U19075 ( .A(n807), .B(n19254), .Z(n19253) );
  XOR U19076 ( .A(n19255), .B(n19252), .Z(n19254) );
  XNOR U19077 ( .A(n19070), .B(n19248), .Z(n19250) );
  XOR U19078 ( .A(n19256), .B(n19257), .Z(n19070) );
  AND U19079 ( .A(n805), .B(n19258), .Z(n19257) );
  XOR U19080 ( .A(n19259), .B(n19256), .Z(n19258) );
  XOR U19081 ( .A(n19260), .B(n19261), .Z(n19248) );
  AND U19082 ( .A(n19262), .B(n19263), .Z(n19261) );
  XOR U19083 ( .A(n19260), .B(n19085), .Z(n19263) );
  XOR U19084 ( .A(n19264), .B(n19265), .Z(n19085) );
  AND U19085 ( .A(n807), .B(n19266), .Z(n19265) );
  XOR U19086 ( .A(n19267), .B(n19264), .Z(n19266) );
  XNOR U19087 ( .A(n19082), .B(n19260), .Z(n19262) );
  XOR U19088 ( .A(n19268), .B(n19269), .Z(n19082) );
  AND U19089 ( .A(n805), .B(n19270), .Z(n19269) );
  XOR U19090 ( .A(n19271), .B(n19268), .Z(n19270) );
  XOR U19091 ( .A(n19272), .B(n19273), .Z(n19260) );
  AND U19092 ( .A(n19274), .B(n19275), .Z(n19273) );
  XOR U19093 ( .A(n19272), .B(n19097), .Z(n19275) );
  XOR U19094 ( .A(n19276), .B(n19277), .Z(n19097) );
  AND U19095 ( .A(n807), .B(n19278), .Z(n19277) );
  XOR U19096 ( .A(n19279), .B(n19276), .Z(n19278) );
  XNOR U19097 ( .A(n19094), .B(n19272), .Z(n19274) );
  XOR U19098 ( .A(n19280), .B(n19281), .Z(n19094) );
  AND U19099 ( .A(n805), .B(n19282), .Z(n19281) );
  XOR U19100 ( .A(n19283), .B(n19280), .Z(n19282) );
  XOR U19101 ( .A(n19284), .B(n19285), .Z(n19272) );
  AND U19102 ( .A(n19286), .B(n19287), .Z(n19285) );
  XOR U19103 ( .A(n19284), .B(n19109), .Z(n19287) );
  XOR U19104 ( .A(n19288), .B(n19289), .Z(n19109) );
  AND U19105 ( .A(n807), .B(n19290), .Z(n19289) );
  XOR U19106 ( .A(n19291), .B(n19288), .Z(n19290) );
  XNOR U19107 ( .A(n19106), .B(n19284), .Z(n19286) );
  XOR U19108 ( .A(n19292), .B(n19293), .Z(n19106) );
  AND U19109 ( .A(n805), .B(n19294), .Z(n19293) );
  XOR U19110 ( .A(n19295), .B(n19292), .Z(n19294) );
  XOR U19111 ( .A(n19296), .B(n19297), .Z(n19284) );
  AND U19112 ( .A(n19298), .B(n19299), .Z(n19297) );
  XOR U19113 ( .A(n19296), .B(n19121), .Z(n19299) );
  XOR U19114 ( .A(n19300), .B(n19301), .Z(n19121) );
  AND U19115 ( .A(n807), .B(n19302), .Z(n19301) );
  XOR U19116 ( .A(n19303), .B(n19300), .Z(n19302) );
  XNOR U19117 ( .A(n19118), .B(n19296), .Z(n19298) );
  XOR U19118 ( .A(n19304), .B(n19305), .Z(n19118) );
  AND U19119 ( .A(n805), .B(n19306), .Z(n19305) );
  XOR U19120 ( .A(n19307), .B(n19304), .Z(n19306) );
  XOR U19121 ( .A(n19308), .B(n19309), .Z(n19296) );
  AND U19122 ( .A(n19310), .B(n19311), .Z(n19309) );
  XOR U19123 ( .A(n19308), .B(n19133), .Z(n19311) );
  XOR U19124 ( .A(n19312), .B(n19313), .Z(n19133) );
  AND U19125 ( .A(n807), .B(n19314), .Z(n19313) );
  XOR U19126 ( .A(n19315), .B(n19312), .Z(n19314) );
  XNOR U19127 ( .A(n19130), .B(n19308), .Z(n19310) );
  XOR U19128 ( .A(n19316), .B(n19317), .Z(n19130) );
  AND U19129 ( .A(n805), .B(n19318), .Z(n19317) );
  XOR U19130 ( .A(n19319), .B(n19316), .Z(n19318) );
  XOR U19131 ( .A(n19320), .B(n19321), .Z(n19308) );
  AND U19132 ( .A(n19322), .B(n19323), .Z(n19321) );
  XOR U19133 ( .A(n19320), .B(n19145), .Z(n19323) );
  XOR U19134 ( .A(n19324), .B(n19325), .Z(n19145) );
  AND U19135 ( .A(n807), .B(n19326), .Z(n19325) );
  XOR U19136 ( .A(n19327), .B(n19324), .Z(n19326) );
  XNOR U19137 ( .A(n19142), .B(n19320), .Z(n19322) );
  XOR U19138 ( .A(n19328), .B(n19329), .Z(n19142) );
  AND U19139 ( .A(n805), .B(n19330), .Z(n19329) );
  XOR U19140 ( .A(n19331), .B(n19328), .Z(n19330) );
  XOR U19141 ( .A(n19332), .B(n19333), .Z(n19320) );
  AND U19142 ( .A(n19334), .B(n19335), .Z(n19333) );
  XNOR U19143 ( .A(n19336), .B(n19158), .Z(n19335) );
  XOR U19144 ( .A(n19337), .B(n19338), .Z(n19158) );
  AND U19145 ( .A(n807), .B(n19339), .Z(n19338) );
  XOR U19146 ( .A(n19337), .B(n19340), .Z(n19339) );
  XNOR U19147 ( .A(n19155), .B(n19332), .Z(n19334) );
  XOR U19148 ( .A(n19341), .B(n19342), .Z(n19155) );
  AND U19149 ( .A(n805), .B(n19343), .Z(n19342) );
  XOR U19150 ( .A(n19341), .B(n19344), .Z(n19343) );
  IV U19151 ( .A(n19336), .Z(n19332) );
  AND U19152 ( .A(n19163), .B(n19166), .Z(n19336) );
  XNOR U19153 ( .A(n19345), .B(n19346), .Z(n19166) );
  AND U19154 ( .A(n807), .B(n19347), .Z(n19346) );
  XNOR U19155 ( .A(n19348), .B(n19345), .Z(n19347) );
  XOR U19156 ( .A(n19349), .B(n19350), .Z(n807) );
  AND U19157 ( .A(n19351), .B(n19352), .Z(n19350) );
  XNOR U19158 ( .A(n19172), .B(n19349), .Z(n19352) );
  AND U19159 ( .A(n19353), .B(n19354), .Z(n19172) );
  XOR U19160 ( .A(n19349), .B(n19173), .Z(n19351) );
  AND U19161 ( .A(n19355), .B(n19356), .Z(n19173) );
  XOR U19162 ( .A(n19357), .B(n19358), .Z(n19349) );
  AND U19163 ( .A(n19359), .B(n19360), .Z(n19358) );
  XOR U19164 ( .A(n19357), .B(n19183), .Z(n19360) );
  XOR U19165 ( .A(n19361), .B(n19362), .Z(n19183) );
  AND U19166 ( .A(n511), .B(n19363), .Z(n19362) );
  XOR U19167 ( .A(n19364), .B(n19361), .Z(n19363) );
  XNOR U19168 ( .A(n19180), .B(n19357), .Z(n19359) );
  XOR U19169 ( .A(n19365), .B(n19366), .Z(n19180) );
  AND U19170 ( .A(n509), .B(n19367), .Z(n19366) );
  XOR U19171 ( .A(n19368), .B(n19365), .Z(n19367) );
  XOR U19172 ( .A(n19369), .B(n19370), .Z(n19357) );
  AND U19173 ( .A(n19371), .B(n19372), .Z(n19370) );
  XOR U19174 ( .A(n19369), .B(n19195), .Z(n19372) );
  XOR U19175 ( .A(n19373), .B(n19374), .Z(n19195) );
  AND U19176 ( .A(n511), .B(n19375), .Z(n19374) );
  XOR U19177 ( .A(n19376), .B(n19373), .Z(n19375) );
  XNOR U19178 ( .A(n19192), .B(n19369), .Z(n19371) );
  XOR U19179 ( .A(n19377), .B(n19378), .Z(n19192) );
  AND U19180 ( .A(n509), .B(n19379), .Z(n19378) );
  XOR U19181 ( .A(n19380), .B(n19377), .Z(n19379) );
  XOR U19182 ( .A(n19381), .B(n19382), .Z(n19369) );
  AND U19183 ( .A(n19383), .B(n19384), .Z(n19382) );
  XOR U19184 ( .A(n19381), .B(n19207), .Z(n19384) );
  XOR U19185 ( .A(n19385), .B(n19386), .Z(n19207) );
  AND U19186 ( .A(n511), .B(n19387), .Z(n19386) );
  XOR U19187 ( .A(n19388), .B(n19385), .Z(n19387) );
  XNOR U19188 ( .A(n19204), .B(n19381), .Z(n19383) );
  XOR U19189 ( .A(n19389), .B(n19390), .Z(n19204) );
  AND U19190 ( .A(n509), .B(n19391), .Z(n19390) );
  XOR U19191 ( .A(n19392), .B(n19389), .Z(n19391) );
  XOR U19192 ( .A(n19393), .B(n19394), .Z(n19381) );
  AND U19193 ( .A(n19395), .B(n19396), .Z(n19394) );
  XOR U19194 ( .A(n19393), .B(n19219), .Z(n19396) );
  XOR U19195 ( .A(n19397), .B(n19398), .Z(n19219) );
  AND U19196 ( .A(n511), .B(n19399), .Z(n19398) );
  XOR U19197 ( .A(n19400), .B(n19397), .Z(n19399) );
  XNOR U19198 ( .A(n19216), .B(n19393), .Z(n19395) );
  XOR U19199 ( .A(n19401), .B(n19402), .Z(n19216) );
  AND U19200 ( .A(n509), .B(n19403), .Z(n19402) );
  XOR U19201 ( .A(n19404), .B(n19401), .Z(n19403) );
  XOR U19202 ( .A(n19405), .B(n19406), .Z(n19393) );
  AND U19203 ( .A(n19407), .B(n19408), .Z(n19406) );
  XOR U19204 ( .A(n19405), .B(n19231), .Z(n19408) );
  XOR U19205 ( .A(n19409), .B(n19410), .Z(n19231) );
  AND U19206 ( .A(n511), .B(n19411), .Z(n19410) );
  XOR U19207 ( .A(n19412), .B(n19409), .Z(n19411) );
  XNOR U19208 ( .A(n19228), .B(n19405), .Z(n19407) );
  XOR U19209 ( .A(n19413), .B(n19414), .Z(n19228) );
  AND U19210 ( .A(n509), .B(n19415), .Z(n19414) );
  XOR U19211 ( .A(n19416), .B(n19413), .Z(n19415) );
  XOR U19212 ( .A(n19417), .B(n19418), .Z(n19405) );
  AND U19213 ( .A(n19419), .B(n19420), .Z(n19418) );
  XOR U19214 ( .A(n19417), .B(n19243), .Z(n19420) );
  XOR U19215 ( .A(n19421), .B(n19422), .Z(n19243) );
  AND U19216 ( .A(n511), .B(n19423), .Z(n19422) );
  XOR U19217 ( .A(n19424), .B(n19421), .Z(n19423) );
  XNOR U19218 ( .A(n19240), .B(n19417), .Z(n19419) );
  XOR U19219 ( .A(n19425), .B(n19426), .Z(n19240) );
  AND U19220 ( .A(n509), .B(n19427), .Z(n19426) );
  XOR U19221 ( .A(n19428), .B(n19425), .Z(n19427) );
  XOR U19222 ( .A(n19429), .B(n19430), .Z(n19417) );
  AND U19223 ( .A(n19431), .B(n19432), .Z(n19430) );
  XOR U19224 ( .A(n19429), .B(n19255), .Z(n19432) );
  XOR U19225 ( .A(n19433), .B(n19434), .Z(n19255) );
  AND U19226 ( .A(n511), .B(n19435), .Z(n19434) );
  XOR U19227 ( .A(n19436), .B(n19433), .Z(n19435) );
  XNOR U19228 ( .A(n19252), .B(n19429), .Z(n19431) );
  XOR U19229 ( .A(n19437), .B(n19438), .Z(n19252) );
  AND U19230 ( .A(n509), .B(n19439), .Z(n19438) );
  XOR U19231 ( .A(n19440), .B(n19437), .Z(n19439) );
  XOR U19232 ( .A(n19441), .B(n19442), .Z(n19429) );
  AND U19233 ( .A(n19443), .B(n19444), .Z(n19442) );
  XOR U19234 ( .A(n19441), .B(n19267), .Z(n19444) );
  XOR U19235 ( .A(n19445), .B(n19446), .Z(n19267) );
  AND U19236 ( .A(n511), .B(n19447), .Z(n19446) );
  XOR U19237 ( .A(n19448), .B(n19445), .Z(n19447) );
  XNOR U19238 ( .A(n19264), .B(n19441), .Z(n19443) );
  XOR U19239 ( .A(n19449), .B(n19450), .Z(n19264) );
  AND U19240 ( .A(n509), .B(n19451), .Z(n19450) );
  XOR U19241 ( .A(n19452), .B(n19449), .Z(n19451) );
  XOR U19242 ( .A(n19453), .B(n19454), .Z(n19441) );
  AND U19243 ( .A(n19455), .B(n19456), .Z(n19454) );
  XOR U19244 ( .A(n19453), .B(n19279), .Z(n19456) );
  XOR U19245 ( .A(n19457), .B(n19458), .Z(n19279) );
  AND U19246 ( .A(n511), .B(n19459), .Z(n19458) );
  XOR U19247 ( .A(n19460), .B(n19457), .Z(n19459) );
  XNOR U19248 ( .A(n19276), .B(n19453), .Z(n19455) );
  XOR U19249 ( .A(n19461), .B(n19462), .Z(n19276) );
  AND U19250 ( .A(n509), .B(n19463), .Z(n19462) );
  XOR U19251 ( .A(n19464), .B(n19461), .Z(n19463) );
  XOR U19252 ( .A(n19465), .B(n19466), .Z(n19453) );
  AND U19253 ( .A(n19467), .B(n19468), .Z(n19466) );
  XOR U19254 ( .A(n19465), .B(n19291), .Z(n19468) );
  XOR U19255 ( .A(n19469), .B(n19470), .Z(n19291) );
  AND U19256 ( .A(n511), .B(n19471), .Z(n19470) );
  XOR U19257 ( .A(n19472), .B(n19469), .Z(n19471) );
  XNOR U19258 ( .A(n19288), .B(n19465), .Z(n19467) );
  XOR U19259 ( .A(n19473), .B(n19474), .Z(n19288) );
  AND U19260 ( .A(n509), .B(n19475), .Z(n19474) );
  XOR U19261 ( .A(n19476), .B(n19473), .Z(n19475) );
  XOR U19262 ( .A(n19477), .B(n19478), .Z(n19465) );
  AND U19263 ( .A(n19479), .B(n19480), .Z(n19478) );
  XOR U19264 ( .A(n19477), .B(n19303), .Z(n19480) );
  XOR U19265 ( .A(n19481), .B(n19482), .Z(n19303) );
  AND U19266 ( .A(n511), .B(n19483), .Z(n19482) );
  XOR U19267 ( .A(n19484), .B(n19481), .Z(n19483) );
  XNOR U19268 ( .A(n19300), .B(n19477), .Z(n19479) );
  XOR U19269 ( .A(n19485), .B(n19486), .Z(n19300) );
  AND U19270 ( .A(n509), .B(n19487), .Z(n19486) );
  XOR U19271 ( .A(n19488), .B(n19485), .Z(n19487) );
  XOR U19272 ( .A(n19489), .B(n19490), .Z(n19477) );
  AND U19273 ( .A(n19491), .B(n19492), .Z(n19490) );
  XOR U19274 ( .A(n19489), .B(n19315), .Z(n19492) );
  XOR U19275 ( .A(n19493), .B(n19494), .Z(n19315) );
  AND U19276 ( .A(n511), .B(n19495), .Z(n19494) );
  XOR U19277 ( .A(n19496), .B(n19493), .Z(n19495) );
  XNOR U19278 ( .A(n19312), .B(n19489), .Z(n19491) );
  XOR U19279 ( .A(n19497), .B(n19498), .Z(n19312) );
  AND U19280 ( .A(n509), .B(n19499), .Z(n19498) );
  XOR U19281 ( .A(n19500), .B(n19497), .Z(n19499) );
  XOR U19282 ( .A(n19501), .B(n19502), .Z(n19489) );
  AND U19283 ( .A(n19503), .B(n19504), .Z(n19502) );
  XOR U19284 ( .A(n19501), .B(n19327), .Z(n19504) );
  XOR U19285 ( .A(n19505), .B(n19506), .Z(n19327) );
  AND U19286 ( .A(n511), .B(n19507), .Z(n19506) );
  XOR U19287 ( .A(n19508), .B(n19505), .Z(n19507) );
  XNOR U19288 ( .A(n19324), .B(n19501), .Z(n19503) );
  XOR U19289 ( .A(n19509), .B(n19510), .Z(n19324) );
  AND U19290 ( .A(n509), .B(n19511), .Z(n19510) );
  XOR U19291 ( .A(n19512), .B(n19509), .Z(n19511) );
  XOR U19292 ( .A(n19513), .B(n19514), .Z(n19501) );
  AND U19293 ( .A(n19515), .B(n19516), .Z(n19514) );
  XNOR U19294 ( .A(n19517), .B(n19340), .Z(n19516) );
  XOR U19295 ( .A(n19518), .B(n19519), .Z(n19340) );
  AND U19296 ( .A(n511), .B(n19520), .Z(n19519) );
  XOR U19297 ( .A(n19518), .B(n19521), .Z(n19520) );
  XNOR U19298 ( .A(n19337), .B(n19513), .Z(n19515) );
  XOR U19299 ( .A(n19522), .B(n19523), .Z(n19337) );
  AND U19300 ( .A(n509), .B(n19524), .Z(n19523) );
  XOR U19301 ( .A(n19522), .B(n19525), .Z(n19524) );
  IV U19302 ( .A(n19517), .Z(n19513) );
  AND U19303 ( .A(n19345), .B(n19348), .Z(n19517) );
  XNOR U19304 ( .A(n19526), .B(n19527), .Z(n19348) );
  AND U19305 ( .A(n511), .B(n19528), .Z(n19527) );
  XNOR U19306 ( .A(n19529), .B(n19526), .Z(n19528) );
  XOR U19307 ( .A(n19530), .B(n19531), .Z(n511) );
  AND U19308 ( .A(n19532), .B(n19533), .Z(n19531) );
  XNOR U19309 ( .A(n19353), .B(n19530), .Z(n19533) );
  AND U19310 ( .A(p_input[1535]), .B(p_input[1519]), .Z(n19353) );
  XOR U19311 ( .A(n19530), .B(n19354), .Z(n19532) );
  AND U19312 ( .A(p_input[1503]), .B(p_input[1487]), .Z(n19354) );
  XOR U19313 ( .A(n19534), .B(n19535), .Z(n19530) );
  AND U19314 ( .A(n19536), .B(n19537), .Z(n19535) );
  XOR U19315 ( .A(n19534), .B(n19364), .Z(n19537) );
  XNOR U19316 ( .A(p_input[1518]), .B(n19538), .Z(n19364) );
  AND U19317 ( .A(n671), .B(n19539), .Z(n19538) );
  XOR U19318 ( .A(p_input[1534]), .B(p_input[1518]), .Z(n19539) );
  XNOR U19319 ( .A(n19361), .B(n19534), .Z(n19536) );
  XOR U19320 ( .A(n19540), .B(n19541), .Z(n19361) );
  AND U19321 ( .A(n669), .B(n19542), .Z(n19541) );
  XOR U19322 ( .A(p_input[1502]), .B(p_input[1486]), .Z(n19542) );
  XOR U19323 ( .A(n19543), .B(n19544), .Z(n19534) );
  AND U19324 ( .A(n19545), .B(n19546), .Z(n19544) );
  XOR U19325 ( .A(n19543), .B(n19376), .Z(n19546) );
  XNOR U19326 ( .A(p_input[1517]), .B(n19547), .Z(n19376) );
  AND U19327 ( .A(n671), .B(n19548), .Z(n19547) );
  XOR U19328 ( .A(p_input[1533]), .B(p_input[1517]), .Z(n19548) );
  XNOR U19329 ( .A(n19373), .B(n19543), .Z(n19545) );
  XOR U19330 ( .A(n19549), .B(n19550), .Z(n19373) );
  AND U19331 ( .A(n669), .B(n19551), .Z(n19550) );
  XOR U19332 ( .A(p_input[1501]), .B(p_input[1485]), .Z(n19551) );
  XOR U19333 ( .A(n19552), .B(n19553), .Z(n19543) );
  AND U19334 ( .A(n19554), .B(n19555), .Z(n19553) );
  XOR U19335 ( .A(n19552), .B(n19388), .Z(n19555) );
  XNOR U19336 ( .A(p_input[1516]), .B(n19556), .Z(n19388) );
  AND U19337 ( .A(n671), .B(n19557), .Z(n19556) );
  XOR U19338 ( .A(p_input[1532]), .B(p_input[1516]), .Z(n19557) );
  XNOR U19339 ( .A(n19385), .B(n19552), .Z(n19554) );
  XOR U19340 ( .A(n19558), .B(n19559), .Z(n19385) );
  AND U19341 ( .A(n669), .B(n19560), .Z(n19559) );
  XOR U19342 ( .A(p_input[1500]), .B(p_input[1484]), .Z(n19560) );
  XOR U19343 ( .A(n19561), .B(n19562), .Z(n19552) );
  AND U19344 ( .A(n19563), .B(n19564), .Z(n19562) );
  XOR U19345 ( .A(n19561), .B(n19400), .Z(n19564) );
  XNOR U19346 ( .A(p_input[1515]), .B(n19565), .Z(n19400) );
  AND U19347 ( .A(n671), .B(n19566), .Z(n19565) );
  XOR U19348 ( .A(p_input[1531]), .B(p_input[1515]), .Z(n19566) );
  XNOR U19349 ( .A(n19397), .B(n19561), .Z(n19563) );
  XOR U19350 ( .A(n19567), .B(n19568), .Z(n19397) );
  AND U19351 ( .A(n669), .B(n19569), .Z(n19568) );
  XOR U19352 ( .A(p_input[1499]), .B(p_input[1483]), .Z(n19569) );
  XOR U19353 ( .A(n19570), .B(n19571), .Z(n19561) );
  AND U19354 ( .A(n19572), .B(n19573), .Z(n19571) );
  XOR U19355 ( .A(n19570), .B(n19412), .Z(n19573) );
  XNOR U19356 ( .A(p_input[1514]), .B(n19574), .Z(n19412) );
  AND U19357 ( .A(n671), .B(n19575), .Z(n19574) );
  XOR U19358 ( .A(p_input[1530]), .B(p_input[1514]), .Z(n19575) );
  XNOR U19359 ( .A(n19409), .B(n19570), .Z(n19572) );
  XOR U19360 ( .A(n19576), .B(n19577), .Z(n19409) );
  AND U19361 ( .A(n669), .B(n19578), .Z(n19577) );
  XOR U19362 ( .A(p_input[1498]), .B(p_input[1482]), .Z(n19578) );
  XOR U19363 ( .A(n19579), .B(n19580), .Z(n19570) );
  AND U19364 ( .A(n19581), .B(n19582), .Z(n19580) );
  XOR U19365 ( .A(n19579), .B(n19424), .Z(n19582) );
  XNOR U19366 ( .A(p_input[1513]), .B(n19583), .Z(n19424) );
  AND U19367 ( .A(n671), .B(n19584), .Z(n19583) );
  XOR U19368 ( .A(p_input[1529]), .B(p_input[1513]), .Z(n19584) );
  XNOR U19369 ( .A(n19421), .B(n19579), .Z(n19581) );
  XOR U19370 ( .A(n19585), .B(n19586), .Z(n19421) );
  AND U19371 ( .A(n669), .B(n19587), .Z(n19586) );
  XOR U19372 ( .A(p_input[1497]), .B(p_input[1481]), .Z(n19587) );
  XOR U19373 ( .A(n19588), .B(n19589), .Z(n19579) );
  AND U19374 ( .A(n19590), .B(n19591), .Z(n19589) );
  XOR U19375 ( .A(n19588), .B(n19436), .Z(n19591) );
  XNOR U19376 ( .A(p_input[1512]), .B(n19592), .Z(n19436) );
  AND U19377 ( .A(n671), .B(n19593), .Z(n19592) );
  XOR U19378 ( .A(p_input[1528]), .B(p_input[1512]), .Z(n19593) );
  XNOR U19379 ( .A(n19433), .B(n19588), .Z(n19590) );
  XOR U19380 ( .A(n19594), .B(n19595), .Z(n19433) );
  AND U19381 ( .A(n669), .B(n19596), .Z(n19595) );
  XOR U19382 ( .A(p_input[1496]), .B(p_input[1480]), .Z(n19596) );
  XOR U19383 ( .A(n19597), .B(n19598), .Z(n19588) );
  AND U19384 ( .A(n19599), .B(n19600), .Z(n19598) );
  XOR U19385 ( .A(n19597), .B(n19448), .Z(n19600) );
  XNOR U19386 ( .A(p_input[1511]), .B(n19601), .Z(n19448) );
  AND U19387 ( .A(n671), .B(n19602), .Z(n19601) );
  XOR U19388 ( .A(p_input[1527]), .B(p_input[1511]), .Z(n19602) );
  XNOR U19389 ( .A(n19445), .B(n19597), .Z(n19599) );
  XOR U19390 ( .A(n19603), .B(n19604), .Z(n19445) );
  AND U19391 ( .A(n669), .B(n19605), .Z(n19604) );
  XOR U19392 ( .A(p_input[1495]), .B(p_input[1479]), .Z(n19605) );
  XOR U19393 ( .A(n19606), .B(n19607), .Z(n19597) );
  AND U19394 ( .A(n19608), .B(n19609), .Z(n19607) );
  XOR U19395 ( .A(n19606), .B(n19460), .Z(n19609) );
  XNOR U19396 ( .A(p_input[1510]), .B(n19610), .Z(n19460) );
  AND U19397 ( .A(n671), .B(n19611), .Z(n19610) );
  XOR U19398 ( .A(p_input[1526]), .B(p_input[1510]), .Z(n19611) );
  XNOR U19399 ( .A(n19457), .B(n19606), .Z(n19608) );
  XOR U19400 ( .A(n19612), .B(n19613), .Z(n19457) );
  AND U19401 ( .A(n669), .B(n19614), .Z(n19613) );
  XOR U19402 ( .A(p_input[1494]), .B(p_input[1478]), .Z(n19614) );
  XOR U19403 ( .A(n19615), .B(n19616), .Z(n19606) );
  AND U19404 ( .A(n19617), .B(n19618), .Z(n19616) );
  XOR U19405 ( .A(n19615), .B(n19472), .Z(n19618) );
  XNOR U19406 ( .A(p_input[1509]), .B(n19619), .Z(n19472) );
  AND U19407 ( .A(n671), .B(n19620), .Z(n19619) );
  XOR U19408 ( .A(p_input[1525]), .B(p_input[1509]), .Z(n19620) );
  XNOR U19409 ( .A(n19469), .B(n19615), .Z(n19617) );
  XOR U19410 ( .A(n19621), .B(n19622), .Z(n19469) );
  AND U19411 ( .A(n669), .B(n19623), .Z(n19622) );
  XOR U19412 ( .A(p_input[1493]), .B(p_input[1477]), .Z(n19623) );
  XOR U19413 ( .A(n19624), .B(n19625), .Z(n19615) );
  AND U19414 ( .A(n19626), .B(n19627), .Z(n19625) );
  XOR U19415 ( .A(n19624), .B(n19484), .Z(n19627) );
  XNOR U19416 ( .A(p_input[1508]), .B(n19628), .Z(n19484) );
  AND U19417 ( .A(n671), .B(n19629), .Z(n19628) );
  XOR U19418 ( .A(p_input[1524]), .B(p_input[1508]), .Z(n19629) );
  XNOR U19419 ( .A(n19481), .B(n19624), .Z(n19626) );
  XOR U19420 ( .A(n19630), .B(n19631), .Z(n19481) );
  AND U19421 ( .A(n669), .B(n19632), .Z(n19631) );
  XOR U19422 ( .A(p_input[1492]), .B(p_input[1476]), .Z(n19632) );
  XOR U19423 ( .A(n19633), .B(n19634), .Z(n19624) );
  AND U19424 ( .A(n19635), .B(n19636), .Z(n19634) );
  XOR U19425 ( .A(n19633), .B(n19496), .Z(n19636) );
  XNOR U19426 ( .A(p_input[1507]), .B(n19637), .Z(n19496) );
  AND U19427 ( .A(n671), .B(n19638), .Z(n19637) );
  XOR U19428 ( .A(p_input[1523]), .B(p_input[1507]), .Z(n19638) );
  XNOR U19429 ( .A(n19493), .B(n19633), .Z(n19635) );
  XOR U19430 ( .A(n19639), .B(n19640), .Z(n19493) );
  AND U19431 ( .A(n669), .B(n19641), .Z(n19640) );
  XOR U19432 ( .A(p_input[1491]), .B(p_input[1475]), .Z(n19641) );
  XOR U19433 ( .A(n19642), .B(n19643), .Z(n19633) );
  AND U19434 ( .A(n19644), .B(n19645), .Z(n19643) );
  XOR U19435 ( .A(n19642), .B(n19508), .Z(n19645) );
  XNOR U19436 ( .A(p_input[1506]), .B(n19646), .Z(n19508) );
  AND U19437 ( .A(n671), .B(n19647), .Z(n19646) );
  XOR U19438 ( .A(p_input[1522]), .B(p_input[1506]), .Z(n19647) );
  XNOR U19439 ( .A(n19505), .B(n19642), .Z(n19644) );
  XOR U19440 ( .A(n19648), .B(n19649), .Z(n19505) );
  AND U19441 ( .A(n669), .B(n19650), .Z(n19649) );
  XOR U19442 ( .A(p_input[1490]), .B(p_input[1474]), .Z(n19650) );
  XOR U19443 ( .A(n19651), .B(n19652), .Z(n19642) );
  AND U19444 ( .A(n19653), .B(n19654), .Z(n19652) );
  XNOR U19445 ( .A(n19655), .B(n19521), .Z(n19654) );
  XNOR U19446 ( .A(p_input[1505]), .B(n19656), .Z(n19521) );
  AND U19447 ( .A(n671), .B(n19657), .Z(n19656) );
  XNOR U19448 ( .A(p_input[1521]), .B(n19658), .Z(n19657) );
  IV U19449 ( .A(p_input[1505]), .Z(n19658) );
  XNOR U19450 ( .A(n19518), .B(n19651), .Z(n19653) );
  XNOR U19451 ( .A(p_input[1473]), .B(n19659), .Z(n19518) );
  AND U19452 ( .A(n669), .B(n19660), .Z(n19659) );
  XOR U19453 ( .A(p_input[1489]), .B(p_input[1473]), .Z(n19660) );
  IV U19454 ( .A(n19655), .Z(n19651) );
  AND U19455 ( .A(n19526), .B(n19529), .Z(n19655) );
  XOR U19456 ( .A(p_input[1504]), .B(n19661), .Z(n19529) );
  AND U19457 ( .A(n671), .B(n19662), .Z(n19661) );
  XOR U19458 ( .A(p_input[1520]), .B(p_input[1504]), .Z(n19662) );
  XOR U19459 ( .A(n19663), .B(n19664), .Z(n671) );
  AND U19460 ( .A(n19665), .B(n19666), .Z(n19664) );
  XNOR U19461 ( .A(p_input[1535]), .B(n19663), .Z(n19666) );
  XOR U19462 ( .A(n19663), .B(p_input[1519]), .Z(n19665) );
  XOR U19463 ( .A(n19667), .B(n19668), .Z(n19663) );
  AND U19464 ( .A(n19669), .B(n19670), .Z(n19668) );
  XNOR U19465 ( .A(p_input[1534]), .B(n19667), .Z(n19670) );
  XOR U19466 ( .A(n19667), .B(p_input[1518]), .Z(n19669) );
  XOR U19467 ( .A(n19671), .B(n19672), .Z(n19667) );
  AND U19468 ( .A(n19673), .B(n19674), .Z(n19672) );
  XNOR U19469 ( .A(p_input[1533]), .B(n19671), .Z(n19674) );
  XOR U19470 ( .A(n19671), .B(p_input[1517]), .Z(n19673) );
  XOR U19471 ( .A(n19675), .B(n19676), .Z(n19671) );
  AND U19472 ( .A(n19677), .B(n19678), .Z(n19676) );
  XNOR U19473 ( .A(p_input[1532]), .B(n19675), .Z(n19678) );
  XOR U19474 ( .A(n19675), .B(p_input[1516]), .Z(n19677) );
  XOR U19475 ( .A(n19679), .B(n19680), .Z(n19675) );
  AND U19476 ( .A(n19681), .B(n19682), .Z(n19680) );
  XNOR U19477 ( .A(p_input[1531]), .B(n19679), .Z(n19682) );
  XOR U19478 ( .A(n19679), .B(p_input[1515]), .Z(n19681) );
  XOR U19479 ( .A(n19683), .B(n19684), .Z(n19679) );
  AND U19480 ( .A(n19685), .B(n19686), .Z(n19684) );
  XNOR U19481 ( .A(p_input[1530]), .B(n19683), .Z(n19686) );
  XOR U19482 ( .A(n19683), .B(p_input[1514]), .Z(n19685) );
  XOR U19483 ( .A(n19687), .B(n19688), .Z(n19683) );
  AND U19484 ( .A(n19689), .B(n19690), .Z(n19688) );
  XNOR U19485 ( .A(p_input[1529]), .B(n19687), .Z(n19690) );
  XOR U19486 ( .A(n19687), .B(p_input[1513]), .Z(n19689) );
  XOR U19487 ( .A(n19691), .B(n19692), .Z(n19687) );
  AND U19488 ( .A(n19693), .B(n19694), .Z(n19692) );
  XNOR U19489 ( .A(p_input[1528]), .B(n19691), .Z(n19694) );
  XOR U19490 ( .A(n19691), .B(p_input[1512]), .Z(n19693) );
  XOR U19491 ( .A(n19695), .B(n19696), .Z(n19691) );
  AND U19492 ( .A(n19697), .B(n19698), .Z(n19696) );
  XNOR U19493 ( .A(p_input[1527]), .B(n19695), .Z(n19698) );
  XOR U19494 ( .A(n19695), .B(p_input[1511]), .Z(n19697) );
  XOR U19495 ( .A(n19699), .B(n19700), .Z(n19695) );
  AND U19496 ( .A(n19701), .B(n19702), .Z(n19700) );
  XNOR U19497 ( .A(p_input[1526]), .B(n19699), .Z(n19702) );
  XOR U19498 ( .A(n19699), .B(p_input[1510]), .Z(n19701) );
  XOR U19499 ( .A(n19703), .B(n19704), .Z(n19699) );
  AND U19500 ( .A(n19705), .B(n19706), .Z(n19704) );
  XNOR U19501 ( .A(p_input[1525]), .B(n19703), .Z(n19706) );
  XOR U19502 ( .A(n19703), .B(p_input[1509]), .Z(n19705) );
  XOR U19503 ( .A(n19707), .B(n19708), .Z(n19703) );
  AND U19504 ( .A(n19709), .B(n19710), .Z(n19708) );
  XNOR U19505 ( .A(p_input[1524]), .B(n19707), .Z(n19710) );
  XOR U19506 ( .A(n19707), .B(p_input[1508]), .Z(n19709) );
  XOR U19507 ( .A(n19711), .B(n19712), .Z(n19707) );
  AND U19508 ( .A(n19713), .B(n19714), .Z(n19712) );
  XNOR U19509 ( .A(p_input[1523]), .B(n19711), .Z(n19714) );
  XOR U19510 ( .A(n19711), .B(p_input[1507]), .Z(n19713) );
  XOR U19511 ( .A(n19715), .B(n19716), .Z(n19711) );
  AND U19512 ( .A(n19717), .B(n19718), .Z(n19716) );
  XNOR U19513 ( .A(p_input[1522]), .B(n19715), .Z(n19718) );
  XOR U19514 ( .A(n19715), .B(p_input[1506]), .Z(n19717) );
  XNOR U19515 ( .A(n19719), .B(n19720), .Z(n19715) );
  AND U19516 ( .A(n19721), .B(n19722), .Z(n19720) );
  XOR U19517 ( .A(p_input[1521]), .B(n19719), .Z(n19722) );
  XNOR U19518 ( .A(p_input[1505]), .B(n19719), .Z(n19721) );
  AND U19519 ( .A(p_input[1520]), .B(n19723), .Z(n19719) );
  IV U19520 ( .A(p_input[1504]), .Z(n19723) );
  XNOR U19521 ( .A(p_input[1472]), .B(n19724), .Z(n19526) );
  AND U19522 ( .A(n669), .B(n19725), .Z(n19724) );
  XOR U19523 ( .A(p_input[1488]), .B(p_input[1472]), .Z(n19725) );
  XOR U19524 ( .A(n19726), .B(n19727), .Z(n669) );
  AND U19525 ( .A(n19728), .B(n19729), .Z(n19727) );
  XNOR U19526 ( .A(p_input[1503]), .B(n19726), .Z(n19729) );
  XOR U19527 ( .A(n19726), .B(p_input[1487]), .Z(n19728) );
  XOR U19528 ( .A(n19730), .B(n19731), .Z(n19726) );
  AND U19529 ( .A(n19732), .B(n19733), .Z(n19731) );
  XNOR U19530 ( .A(p_input[1502]), .B(n19730), .Z(n19733) );
  XNOR U19531 ( .A(n19730), .B(n19540), .Z(n19732) );
  IV U19532 ( .A(p_input[1486]), .Z(n19540) );
  XOR U19533 ( .A(n19734), .B(n19735), .Z(n19730) );
  AND U19534 ( .A(n19736), .B(n19737), .Z(n19735) );
  XNOR U19535 ( .A(p_input[1501]), .B(n19734), .Z(n19737) );
  XNOR U19536 ( .A(n19734), .B(n19549), .Z(n19736) );
  IV U19537 ( .A(p_input[1485]), .Z(n19549) );
  XOR U19538 ( .A(n19738), .B(n19739), .Z(n19734) );
  AND U19539 ( .A(n19740), .B(n19741), .Z(n19739) );
  XNOR U19540 ( .A(p_input[1500]), .B(n19738), .Z(n19741) );
  XNOR U19541 ( .A(n19738), .B(n19558), .Z(n19740) );
  IV U19542 ( .A(p_input[1484]), .Z(n19558) );
  XOR U19543 ( .A(n19742), .B(n19743), .Z(n19738) );
  AND U19544 ( .A(n19744), .B(n19745), .Z(n19743) );
  XNOR U19545 ( .A(p_input[1499]), .B(n19742), .Z(n19745) );
  XNOR U19546 ( .A(n19742), .B(n19567), .Z(n19744) );
  IV U19547 ( .A(p_input[1483]), .Z(n19567) );
  XOR U19548 ( .A(n19746), .B(n19747), .Z(n19742) );
  AND U19549 ( .A(n19748), .B(n19749), .Z(n19747) );
  XNOR U19550 ( .A(p_input[1498]), .B(n19746), .Z(n19749) );
  XNOR U19551 ( .A(n19746), .B(n19576), .Z(n19748) );
  IV U19552 ( .A(p_input[1482]), .Z(n19576) );
  XOR U19553 ( .A(n19750), .B(n19751), .Z(n19746) );
  AND U19554 ( .A(n19752), .B(n19753), .Z(n19751) );
  XNOR U19555 ( .A(p_input[1497]), .B(n19750), .Z(n19753) );
  XNOR U19556 ( .A(n19750), .B(n19585), .Z(n19752) );
  IV U19557 ( .A(p_input[1481]), .Z(n19585) );
  XOR U19558 ( .A(n19754), .B(n19755), .Z(n19750) );
  AND U19559 ( .A(n19756), .B(n19757), .Z(n19755) );
  XNOR U19560 ( .A(p_input[1496]), .B(n19754), .Z(n19757) );
  XNOR U19561 ( .A(n19754), .B(n19594), .Z(n19756) );
  IV U19562 ( .A(p_input[1480]), .Z(n19594) );
  XOR U19563 ( .A(n19758), .B(n19759), .Z(n19754) );
  AND U19564 ( .A(n19760), .B(n19761), .Z(n19759) );
  XNOR U19565 ( .A(p_input[1495]), .B(n19758), .Z(n19761) );
  XNOR U19566 ( .A(n19758), .B(n19603), .Z(n19760) );
  IV U19567 ( .A(p_input[1479]), .Z(n19603) );
  XOR U19568 ( .A(n19762), .B(n19763), .Z(n19758) );
  AND U19569 ( .A(n19764), .B(n19765), .Z(n19763) );
  XNOR U19570 ( .A(p_input[1494]), .B(n19762), .Z(n19765) );
  XNOR U19571 ( .A(n19762), .B(n19612), .Z(n19764) );
  IV U19572 ( .A(p_input[1478]), .Z(n19612) );
  XOR U19573 ( .A(n19766), .B(n19767), .Z(n19762) );
  AND U19574 ( .A(n19768), .B(n19769), .Z(n19767) );
  XNOR U19575 ( .A(p_input[1493]), .B(n19766), .Z(n19769) );
  XNOR U19576 ( .A(n19766), .B(n19621), .Z(n19768) );
  IV U19577 ( .A(p_input[1477]), .Z(n19621) );
  XOR U19578 ( .A(n19770), .B(n19771), .Z(n19766) );
  AND U19579 ( .A(n19772), .B(n19773), .Z(n19771) );
  XNOR U19580 ( .A(p_input[1492]), .B(n19770), .Z(n19773) );
  XNOR U19581 ( .A(n19770), .B(n19630), .Z(n19772) );
  IV U19582 ( .A(p_input[1476]), .Z(n19630) );
  XOR U19583 ( .A(n19774), .B(n19775), .Z(n19770) );
  AND U19584 ( .A(n19776), .B(n19777), .Z(n19775) );
  XNOR U19585 ( .A(p_input[1491]), .B(n19774), .Z(n19777) );
  XNOR U19586 ( .A(n19774), .B(n19639), .Z(n19776) );
  IV U19587 ( .A(p_input[1475]), .Z(n19639) );
  XOR U19588 ( .A(n19778), .B(n19779), .Z(n19774) );
  AND U19589 ( .A(n19780), .B(n19781), .Z(n19779) );
  XNOR U19590 ( .A(p_input[1490]), .B(n19778), .Z(n19781) );
  XNOR U19591 ( .A(n19778), .B(n19648), .Z(n19780) );
  IV U19592 ( .A(p_input[1474]), .Z(n19648) );
  XNOR U19593 ( .A(n19782), .B(n19783), .Z(n19778) );
  AND U19594 ( .A(n19784), .B(n19785), .Z(n19783) );
  XOR U19595 ( .A(p_input[1489]), .B(n19782), .Z(n19785) );
  XNOR U19596 ( .A(p_input[1473]), .B(n19782), .Z(n19784) );
  AND U19597 ( .A(p_input[1488]), .B(n19786), .Z(n19782) );
  IV U19598 ( .A(p_input[1472]), .Z(n19786) );
  XOR U19599 ( .A(n19787), .B(n19788), .Z(n19345) );
  AND U19600 ( .A(n509), .B(n19789), .Z(n19788) );
  XNOR U19601 ( .A(n19790), .B(n19787), .Z(n19789) );
  XOR U19602 ( .A(n19791), .B(n19792), .Z(n509) );
  AND U19603 ( .A(n19793), .B(n19794), .Z(n19792) );
  XNOR U19604 ( .A(n19355), .B(n19791), .Z(n19794) );
  AND U19605 ( .A(p_input[1471]), .B(p_input[1455]), .Z(n19355) );
  XOR U19606 ( .A(n19791), .B(n19356), .Z(n19793) );
  AND U19607 ( .A(p_input[1439]), .B(p_input[1423]), .Z(n19356) );
  XOR U19608 ( .A(n19795), .B(n19796), .Z(n19791) );
  AND U19609 ( .A(n19797), .B(n19798), .Z(n19796) );
  XOR U19610 ( .A(n19795), .B(n19368), .Z(n19798) );
  XNOR U19611 ( .A(p_input[1454]), .B(n19799), .Z(n19368) );
  AND U19612 ( .A(n675), .B(n19800), .Z(n19799) );
  XOR U19613 ( .A(p_input[1470]), .B(p_input[1454]), .Z(n19800) );
  XNOR U19614 ( .A(n19365), .B(n19795), .Z(n19797) );
  XOR U19615 ( .A(n19801), .B(n19802), .Z(n19365) );
  AND U19616 ( .A(n672), .B(n19803), .Z(n19802) );
  XOR U19617 ( .A(p_input[1438]), .B(p_input[1422]), .Z(n19803) );
  XOR U19618 ( .A(n19804), .B(n19805), .Z(n19795) );
  AND U19619 ( .A(n19806), .B(n19807), .Z(n19805) );
  XOR U19620 ( .A(n19804), .B(n19380), .Z(n19807) );
  XNOR U19621 ( .A(p_input[1453]), .B(n19808), .Z(n19380) );
  AND U19622 ( .A(n675), .B(n19809), .Z(n19808) );
  XOR U19623 ( .A(p_input[1469]), .B(p_input[1453]), .Z(n19809) );
  XNOR U19624 ( .A(n19377), .B(n19804), .Z(n19806) );
  XOR U19625 ( .A(n19810), .B(n19811), .Z(n19377) );
  AND U19626 ( .A(n672), .B(n19812), .Z(n19811) );
  XOR U19627 ( .A(p_input[1437]), .B(p_input[1421]), .Z(n19812) );
  XOR U19628 ( .A(n19813), .B(n19814), .Z(n19804) );
  AND U19629 ( .A(n19815), .B(n19816), .Z(n19814) );
  XOR U19630 ( .A(n19813), .B(n19392), .Z(n19816) );
  XNOR U19631 ( .A(p_input[1452]), .B(n19817), .Z(n19392) );
  AND U19632 ( .A(n675), .B(n19818), .Z(n19817) );
  XOR U19633 ( .A(p_input[1468]), .B(p_input[1452]), .Z(n19818) );
  XNOR U19634 ( .A(n19389), .B(n19813), .Z(n19815) );
  XOR U19635 ( .A(n19819), .B(n19820), .Z(n19389) );
  AND U19636 ( .A(n672), .B(n19821), .Z(n19820) );
  XOR U19637 ( .A(p_input[1436]), .B(p_input[1420]), .Z(n19821) );
  XOR U19638 ( .A(n19822), .B(n19823), .Z(n19813) );
  AND U19639 ( .A(n19824), .B(n19825), .Z(n19823) );
  XOR U19640 ( .A(n19822), .B(n19404), .Z(n19825) );
  XNOR U19641 ( .A(p_input[1451]), .B(n19826), .Z(n19404) );
  AND U19642 ( .A(n675), .B(n19827), .Z(n19826) );
  XOR U19643 ( .A(p_input[1467]), .B(p_input[1451]), .Z(n19827) );
  XNOR U19644 ( .A(n19401), .B(n19822), .Z(n19824) );
  XOR U19645 ( .A(n19828), .B(n19829), .Z(n19401) );
  AND U19646 ( .A(n672), .B(n19830), .Z(n19829) );
  XOR U19647 ( .A(p_input[1435]), .B(p_input[1419]), .Z(n19830) );
  XOR U19648 ( .A(n19831), .B(n19832), .Z(n19822) );
  AND U19649 ( .A(n19833), .B(n19834), .Z(n19832) );
  XOR U19650 ( .A(n19831), .B(n19416), .Z(n19834) );
  XNOR U19651 ( .A(p_input[1450]), .B(n19835), .Z(n19416) );
  AND U19652 ( .A(n675), .B(n19836), .Z(n19835) );
  XOR U19653 ( .A(p_input[1466]), .B(p_input[1450]), .Z(n19836) );
  XNOR U19654 ( .A(n19413), .B(n19831), .Z(n19833) );
  XOR U19655 ( .A(n19837), .B(n19838), .Z(n19413) );
  AND U19656 ( .A(n672), .B(n19839), .Z(n19838) );
  XOR U19657 ( .A(p_input[1434]), .B(p_input[1418]), .Z(n19839) );
  XOR U19658 ( .A(n19840), .B(n19841), .Z(n19831) );
  AND U19659 ( .A(n19842), .B(n19843), .Z(n19841) );
  XOR U19660 ( .A(n19840), .B(n19428), .Z(n19843) );
  XNOR U19661 ( .A(p_input[1449]), .B(n19844), .Z(n19428) );
  AND U19662 ( .A(n675), .B(n19845), .Z(n19844) );
  XOR U19663 ( .A(p_input[1465]), .B(p_input[1449]), .Z(n19845) );
  XNOR U19664 ( .A(n19425), .B(n19840), .Z(n19842) );
  XOR U19665 ( .A(n19846), .B(n19847), .Z(n19425) );
  AND U19666 ( .A(n672), .B(n19848), .Z(n19847) );
  XOR U19667 ( .A(p_input[1433]), .B(p_input[1417]), .Z(n19848) );
  XOR U19668 ( .A(n19849), .B(n19850), .Z(n19840) );
  AND U19669 ( .A(n19851), .B(n19852), .Z(n19850) );
  XOR U19670 ( .A(n19849), .B(n19440), .Z(n19852) );
  XNOR U19671 ( .A(p_input[1448]), .B(n19853), .Z(n19440) );
  AND U19672 ( .A(n675), .B(n19854), .Z(n19853) );
  XOR U19673 ( .A(p_input[1464]), .B(p_input[1448]), .Z(n19854) );
  XNOR U19674 ( .A(n19437), .B(n19849), .Z(n19851) );
  XOR U19675 ( .A(n19855), .B(n19856), .Z(n19437) );
  AND U19676 ( .A(n672), .B(n19857), .Z(n19856) );
  XOR U19677 ( .A(p_input[1432]), .B(p_input[1416]), .Z(n19857) );
  XOR U19678 ( .A(n19858), .B(n19859), .Z(n19849) );
  AND U19679 ( .A(n19860), .B(n19861), .Z(n19859) );
  XOR U19680 ( .A(n19858), .B(n19452), .Z(n19861) );
  XNOR U19681 ( .A(p_input[1447]), .B(n19862), .Z(n19452) );
  AND U19682 ( .A(n675), .B(n19863), .Z(n19862) );
  XOR U19683 ( .A(p_input[1463]), .B(p_input[1447]), .Z(n19863) );
  XNOR U19684 ( .A(n19449), .B(n19858), .Z(n19860) );
  XOR U19685 ( .A(n19864), .B(n19865), .Z(n19449) );
  AND U19686 ( .A(n672), .B(n19866), .Z(n19865) );
  XOR U19687 ( .A(p_input[1431]), .B(p_input[1415]), .Z(n19866) );
  XOR U19688 ( .A(n19867), .B(n19868), .Z(n19858) );
  AND U19689 ( .A(n19869), .B(n19870), .Z(n19868) );
  XOR U19690 ( .A(n19867), .B(n19464), .Z(n19870) );
  XNOR U19691 ( .A(p_input[1446]), .B(n19871), .Z(n19464) );
  AND U19692 ( .A(n675), .B(n19872), .Z(n19871) );
  XOR U19693 ( .A(p_input[1462]), .B(p_input[1446]), .Z(n19872) );
  XNOR U19694 ( .A(n19461), .B(n19867), .Z(n19869) );
  XOR U19695 ( .A(n19873), .B(n19874), .Z(n19461) );
  AND U19696 ( .A(n672), .B(n19875), .Z(n19874) );
  XOR U19697 ( .A(p_input[1430]), .B(p_input[1414]), .Z(n19875) );
  XOR U19698 ( .A(n19876), .B(n19877), .Z(n19867) );
  AND U19699 ( .A(n19878), .B(n19879), .Z(n19877) );
  XOR U19700 ( .A(n19876), .B(n19476), .Z(n19879) );
  XNOR U19701 ( .A(p_input[1445]), .B(n19880), .Z(n19476) );
  AND U19702 ( .A(n675), .B(n19881), .Z(n19880) );
  XOR U19703 ( .A(p_input[1461]), .B(p_input[1445]), .Z(n19881) );
  XNOR U19704 ( .A(n19473), .B(n19876), .Z(n19878) );
  XOR U19705 ( .A(n19882), .B(n19883), .Z(n19473) );
  AND U19706 ( .A(n672), .B(n19884), .Z(n19883) );
  XOR U19707 ( .A(p_input[1429]), .B(p_input[1413]), .Z(n19884) );
  XOR U19708 ( .A(n19885), .B(n19886), .Z(n19876) );
  AND U19709 ( .A(n19887), .B(n19888), .Z(n19886) );
  XOR U19710 ( .A(n19885), .B(n19488), .Z(n19888) );
  XNOR U19711 ( .A(p_input[1444]), .B(n19889), .Z(n19488) );
  AND U19712 ( .A(n675), .B(n19890), .Z(n19889) );
  XOR U19713 ( .A(p_input[1460]), .B(p_input[1444]), .Z(n19890) );
  XNOR U19714 ( .A(n19485), .B(n19885), .Z(n19887) );
  XOR U19715 ( .A(n19891), .B(n19892), .Z(n19485) );
  AND U19716 ( .A(n672), .B(n19893), .Z(n19892) );
  XOR U19717 ( .A(p_input[1428]), .B(p_input[1412]), .Z(n19893) );
  XOR U19718 ( .A(n19894), .B(n19895), .Z(n19885) );
  AND U19719 ( .A(n19896), .B(n19897), .Z(n19895) );
  XOR U19720 ( .A(n19894), .B(n19500), .Z(n19897) );
  XNOR U19721 ( .A(p_input[1443]), .B(n19898), .Z(n19500) );
  AND U19722 ( .A(n675), .B(n19899), .Z(n19898) );
  XOR U19723 ( .A(p_input[1459]), .B(p_input[1443]), .Z(n19899) );
  XNOR U19724 ( .A(n19497), .B(n19894), .Z(n19896) );
  XOR U19725 ( .A(n19900), .B(n19901), .Z(n19497) );
  AND U19726 ( .A(n672), .B(n19902), .Z(n19901) );
  XOR U19727 ( .A(p_input[1427]), .B(p_input[1411]), .Z(n19902) );
  XOR U19728 ( .A(n19903), .B(n19904), .Z(n19894) );
  AND U19729 ( .A(n19905), .B(n19906), .Z(n19904) );
  XOR U19730 ( .A(n19903), .B(n19512), .Z(n19906) );
  XNOR U19731 ( .A(p_input[1442]), .B(n19907), .Z(n19512) );
  AND U19732 ( .A(n675), .B(n19908), .Z(n19907) );
  XOR U19733 ( .A(p_input[1458]), .B(p_input[1442]), .Z(n19908) );
  XNOR U19734 ( .A(n19509), .B(n19903), .Z(n19905) );
  XOR U19735 ( .A(n19909), .B(n19910), .Z(n19509) );
  AND U19736 ( .A(n672), .B(n19911), .Z(n19910) );
  XOR U19737 ( .A(p_input[1426]), .B(p_input[1410]), .Z(n19911) );
  XOR U19738 ( .A(n19912), .B(n19913), .Z(n19903) );
  AND U19739 ( .A(n19914), .B(n19915), .Z(n19913) );
  XNOR U19740 ( .A(n19916), .B(n19525), .Z(n19915) );
  XNOR U19741 ( .A(p_input[1441]), .B(n19917), .Z(n19525) );
  AND U19742 ( .A(n675), .B(n19918), .Z(n19917) );
  XNOR U19743 ( .A(p_input[1457]), .B(n19919), .Z(n19918) );
  IV U19744 ( .A(p_input[1441]), .Z(n19919) );
  XNOR U19745 ( .A(n19522), .B(n19912), .Z(n19914) );
  XNOR U19746 ( .A(p_input[1409]), .B(n19920), .Z(n19522) );
  AND U19747 ( .A(n672), .B(n19921), .Z(n19920) );
  XOR U19748 ( .A(p_input[1425]), .B(p_input[1409]), .Z(n19921) );
  IV U19749 ( .A(n19916), .Z(n19912) );
  AND U19750 ( .A(n19787), .B(n19790), .Z(n19916) );
  XOR U19751 ( .A(p_input[1440]), .B(n19922), .Z(n19790) );
  AND U19752 ( .A(n675), .B(n19923), .Z(n19922) );
  XOR U19753 ( .A(p_input[1456]), .B(p_input[1440]), .Z(n19923) );
  XOR U19754 ( .A(n19924), .B(n19925), .Z(n675) );
  AND U19755 ( .A(n19926), .B(n19927), .Z(n19925) );
  XNOR U19756 ( .A(p_input[1471]), .B(n19924), .Z(n19927) );
  XOR U19757 ( .A(n19924), .B(p_input[1455]), .Z(n19926) );
  XOR U19758 ( .A(n19928), .B(n19929), .Z(n19924) );
  AND U19759 ( .A(n19930), .B(n19931), .Z(n19929) );
  XNOR U19760 ( .A(p_input[1470]), .B(n19928), .Z(n19931) );
  XOR U19761 ( .A(n19928), .B(p_input[1454]), .Z(n19930) );
  XOR U19762 ( .A(n19932), .B(n19933), .Z(n19928) );
  AND U19763 ( .A(n19934), .B(n19935), .Z(n19933) );
  XNOR U19764 ( .A(p_input[1469]), .B(n19932), .Z(n19935) );
  XOR U19765 ( .A(n19932), .B(p_input[1453]), .Z(n19934) );
  XOR U19766 ( .A(n19936), .B(n19937), .Z(n19932) );
  AND U19767 ( .A(n19938), .B(n19939), .Z(n19937) );
  XNOR U19768 ( .A(p_input[1468]), .B(n19936), .Z(n19939) );
  XOR U19769 ( .A(n19936), .B(p_input[1452]), .Z(n19938) );
  XOR U19770 ( .A(n19940), .B(n19941), .Z(n19936) );
  AND U19771 ( .A(n19942), .B(n19943), .Z(n19941) );
  XNOR U19772 ( .A(p_input[1467]), .B(n19940), .Z(n19943) );
  XOR U19773 ( .A(n19940), .B(p_input[1451]), .Z(n19942) );
  XOR U19774 ( .A(n19944), .B(n19945), .Z(n19940) );
  AND U19775 ( .A(n19946), .B(n19947), .Z(n19945) );
  XNOR U19776 ( .A(p_input[1466]), .B(n19944), .Z(n19947) );
  XOR U19777 ( .A(n19944), .B(p_input[1450]), .Z(n19946) );
  XOR U19778 ( .A(n19948), .B(n19949), .Z(n19944) );
  AND U19779 ( .A(n19950), .B(n19951), .Z(n19949) );
  XNOR U19780 ( .A(p_input[1465]), .B(n19948), .Z(n19951) );
  XOR U19781 ( .A(n19948), .B(p_input[1449]), .Z(n19950) );
  XOR U19782 ( .A(n19952), .B(n19953), .Z(n19948) );
  AND U19783 ( .A(n19954), .B(n19955), .Z(n19953) );
  XNOR U19784 ( .A(p_input[1464]), .B(n19952), .Z(n19955) );
  XOR U19785 ( .A(n19952), .B(p_input[1448]), .Z(n19954) );
  XOR U19786 ( .A(n19956), .B(n19957), .Z(n19952) );
  AND U19787 ( .A(n19958), .B(n19959), .Z(n19957) );
  XNOR U19788 ( .A(p_input[1463]), .B(n19956), .Z(n19959) );
  XOR U19789 ( .A(n19956), .B(p_input[1447]), .Z(n19958) );
  XOR U19790 ( .A(n19960), .B(n19961), .Z(n19956) );
  AND U19791 ( .A(n19962), .B(n19963), .Z(n19961) );
  XNOR U19792 ( .A(p_input[1462]), .B(n19960), .Z(n19963) );
  XOR U19793 ( .A(n19960), .B(p_input[1446]), .Z(n19962) );
  XOR U19794 ( .A(n19964), .B(n19965), .Z(n19960) );
  AND U19795 ( .A(n19966), .B(n19967), .Z(n19965) );
  XNOR U19796 ( .A(p_input[1461]), .B(n19964), .Z(n19967) );
  XOR U19797 ( .A(n19964), .B(p_input[1445]), .Z(n19966) );
  XOR U19798 ( .A(n19968), .B(n19969), .Z(n19964) );
  AND U19799 ( .A(n19970), .B(n19971), .Z(n19969) );
  XNOR U19800 ( .A(p_input[1460]), .B(n19968), .Z(n19971) );
  XOR U19801 ( .A(n19968), .B(p_input[1444]), .Z(n19970) );
  XOR U19802 ( .A(n19972), .B(n19973), .Z(n19968) );
  AND U19803 ( .A(n19974), .B(n19975), .Z(n19973) );
  XNOR U19804 ( .A(p_input[1459]), .B(n19972), .Z(n19975) );
  XOR U19805 ( .A(n19972), .B(p_input[1443]), .Z(n19974) );
  XOR U19806 ( .A(n19976), .B(n19977), .Z(n19972) );
  AND U19807 ( .A(n19978), .B(n19979), .Z(n19977) );
  XNOR U19808 ( .A(p_input[1458]), .B(n19976), .Z(n19979) );
  XOR U19809 ( .A(n19976), .B(p_input[1442]), .Z(n19978) );
  XNOR U19810 ( .A(n19980), .B(n19981), .Z(n19976) );
  AND U19811 ( .A(n19982), .B(n19983), .Z(n19981) );
  XOR U19812 ( .A(p_input[1457]), .B(n19980), .Z(n19983) );
  XNOR U19813 ( .A(p_input[1441]), .B(n19980), .Z(n19982) );
  AND U19814 ( .A(p_input[1456]), .B(n19984), .Z(n19980) );
  IV U19815 ( .A(p_input[1440]), .Z(n19984) );
  XNOR U19816 ( .A(p_input[1408]), .B(n19985), .Z(n19787) );
  AND U19817 ( .A(n672), .B(n19986), .Z(n19985) );
  XOR U19818 ( .A(p_input[1424]), .B(p_input[1408]), .Z(n19986) );
  XOR U19819 ( .A(n19987), .B(n19988), .Z(n672) );
  AND U19820 ( .A(n19989), .B(n19990), .Z(n19988) );
  XNOR U19821 ( .A(p_input[1439]), .B(n19987), .Z(n19990) );
  XOR U19822 ( .A(n19987), .B(p_input[1423]), .Z(n19989) );
  XOR U19823 ( .A(n19991), .B(n19992), .Z(n19987) );
  AND U19824 ( .A(n19993), .B(n19994), .Z(n19992) );
  XNOR U19825 ( .A(p_input[1438]), .B(n19991), .Z(n19994) );
  XNOR U19826 ( .A(n19991), .B(n19801), .Z(n19993) );
  IV U19827 ( .A(p_input[1422]), .Z(n19801) );
  XOR U19828 ( .A(n19995), .B(n19996), .Z(n19991) );
  AND U19829 ( .A(n19997), .B(n19998), .Z(n19996) );
  XNOR U19830 ( .A(p_input[1437]), .B(n19995), .Z(n19998) );
  XNOR U19831 ( .A(n19995), .B(n19810), .Z(n19997) );
  IV U19832 ( .A(p_input[1421]), .Z(n19810) );
  XOR U19833 ( .A(n19999), .B(n20000), .Z(n19995) );
  AND U19834 ( .A(n20001), .B(n20002), .Z(n20000) );
  XNOR U19835 ( .A(p_input[1436]), .B(n19999), .Z(n20002) );
  XNOR U19836 ( .A(n19999), .B(n19819), .Z(n20001) );
  IV U19837 ( .A(p_input[1420]), .Z(n19819) );
  XOR U19838 ( .A(n20003), .B(n20004), .Z(n19999) );
  AND U19839 ( .A(n20005), .B(n20006), .Z(n20004) );
  XNOR U19840 ( .A(p_input[1435]), .B(n20003), .Z(n20006) );
  XNOR U19841 ( .A(n20003), .B(n19828), .Z(n20005) );
  IV U19842 ( .A(p_input[1419]), .Z(n19828) );
  XOR U19843 ( .A(n20007), .B(n20008), .Z(n20003) );
  AND U19844 ( .A(n20009), .B(n20010), .Z(n20008) );
  XNOR U19845 ( .A(p_input[1434]), .B(n20007), .Z(n20010) );
  XNOR U19846 ( .A(n20007), .B(n19837), .Z(n20009) );
  IV U19847 ( .A(p_input[1418]), .Z(n19837) );
  XOR U19848 ( .A(n20011), .B(n20012), .Z(n20007) );
  AND U19849 ( .A(n20013), .B(n20014), .Z(n20012) );
  XNOR U19850 ( .A(p_input[1433]), .B(n20011), .Z(n20014) );
  XNOR U19851 ( .A(n20011), .B(n19846), .Z(n20013) );
  IV U19852 ( .A(p_input[1417]), .Z(n19846) );
  XOR U19853 ( .A(n20015), .B(n20016), .Z(n20011) );
  AND U19854 ( .A(n20017), .B(n20018), .Z(n20016) );
  XNOR U19855 ( .A(p_input[1432]), .B(n20015), .Z(n20018) );
  XNOR U19856 ( .A(n20015), .B(n19855), .Z(n20017) );
  IV U19857 ( .A(p_input[1416]), .Z(n19855) );
  XOR U19858 ( .A(n20019), .B(n20020), .Z(n20015) );
  AND U19859 ( .A(n20021), .B(n20022), .Z(n20020) );
  XNOR U19860 ( .A(p_input[1431]), .B(n20019), .Z(n20022) );
  XNOR U19861 ( .A(n20019), .B(n19864), .Z(n20021) );
  IV U19862 ( .A(p_input[1415]), .Z(n19864) );
  XOR U19863 ( .A(n20023), .B(n20024), .Z(n20019) );
  AND U19864 ( .A(n20025), .B(n20026), .Z(n20024) );
  XNOR U19865 ( .A(p_input[1430]), .B(n20023), .Z(n20026) );
  XNOR U19866 ( .A(n20023), .B(n19873), .Z(n20025) );
  IV U19867 ( .A(p_input[1414]), .Z(n19873) );
  XOR U19868 ( .A(n20027), .B(n20028), .Z(n20023) );
  AND U19869 ( .A(n20029), .B(n20030), .Z(n20028) );
  XNOR U19870 ( .A(p_input[1429]), .B(n20027), .Z(n20030) );
  XNOR U19871 ( .A(n20027), .B(n19882), .Z(n20029) );
  IV U19872 ( .A(p_input[1413]), .Z(n19882) );
  XOR U19873 ( .A(n20031), .B(n20032), .Z(n20027) );
  AND U19874 ( .A(n20033), .B(n20034), .Z(n20032) );
  XNOR U19875 ( .A(p_input[1428]), .B(n20031), .Z(n20034) );
  XNOR U19876 ( .A(n20031), .B(n19891), .Z(n20033) );
  IV U19877 ( .A(p_input[1412]), .Z(n19891) );
  XOR U19878 ( .A(n20035), .B(n20036), .Z(n20031) );
  AND U19879 ( .A(n20037), .B(n20038), .Z(n20036) );
  XNOR U19880 ( .A(p_input[1427]), .B(n20035), .Z(n20038) );
  XNOR U19881 ( .A(n20035), .B(n19900), .Z(n20037) );
  IV U19882 ( .A(p_input[1411]), .Z(n19900) );
  XOR U19883 ( .A(n20039), .B(n20040), .Z(n20035) );
  AND U19884 ( .A(n20041), .B(n20042), .Z(n20040) );
  XNOR U19885 ( .A(p_input[1426]), .B(n20039), .Z(n20042) );
  XNOR U19886 ( .A(n20039), .B(n19909), .Z(n20041) );
  IV U19887 ( .A(p_input[1410]), .Z(n19909) );
  XNOR U19888 ( .A(n20043), .B(n20044), .Z(n20039) );
  AND U19889 ( .A(n20045), .B(n20046), .Z(n20044) );
  XOR U19890 ( .A(p_input[1425]), .B(n20043), .Z(n20046) );
  XNOR U19891 ( .A(p_input[1409]), .B(n20043), .Z(n20045) );
  AND U19892 ( .A(p_input[1424]), .B(n20047), .Z(n20043) );
  IV U19893 ( .A(p_input[1408]), .Z(n20047) );
  XOR U19894 ( .A(n20048), .B(n20049), .Z(n19163) );
  AND U19895 ( .A(n805), .B(n20050), .Z(n20049) );
  XNOR U19896 ( .A(n20051), .B(n20048), .Z(n20050) );
  XOR U19897 ( .A(n20052), .B(n20053), .Z(n805) );
  AND U19898 ( .A(n20054), .B(n20055), .Z(n20053) );
  XNOR U19899 ( .A(n19175), .B(n20052), .Z(n20055) );
  AND U19900 ( .A(n20056), .B(n20057), .Z(n19175) );
  XOR U19901 ( .A(n20052), .B(n19174), .Z(n20054) );
  AND U19902 ( .A(n20058), .B(n20059), .Z(n19174) );
  XOR U19903 ( .A(n20060), .B(n20061), .Z(n20052) );
  AND U19904 ( .A(n20062), .B(n20063), .Z(n20061) );
  XOR U19905 ( .A(n20060), .B(n19187), .Z(n20063) );
  XOR U19906 ( .A(n20064), .B(n20065), .Z(n19187) );
  AND U19907 ( .A(n515), .B(n20066), .Z(n20065) );
  XOR U19908 ( .A(n20067), .B(n20064), .Z(n20066) );
  XNOR U19909 ( .A(n19184), .B(n20060), .Z(n20062) );
  XOR U19910 ( .A(n20068), .B(n20069), .Z(n19184) );
  AND U19911 ( .A(n512), .B(n20070), .Z(n20069) );
  XOR U19912 ( .A(n20071), .B(n20068), .Z(n20070) );
  XOR U19913 ( .A(n20072), .B(n20073), .Z(n20060) );
  AND U19914 ( .A(n20074), .B(n20075), .Z(n20073) );
  XOR U19915 ( .A(n20072), .B(n19199), .Z(n20075) );
  XOR U19916 ( .A(n20076), .B(n20077), .Z(n19199) );
  AND U19917 ( .A(n515), .B(n20078), .Z(n20077) );
  XOR U19918 ( .A(n20079), .B(n20076), .Z(n20078) );
  XNOR U19919 ( .A(n19196), .B(n20072), .Z(n20074) );
  XOR U19920 ( .A(n20080), .B(n20081), .Z(n19196) );
  AND U19921 ( .A(n512), .B(n20082), .Z(n20081) );
  XOR U19922 ( .A(n20083), .B(n20080), .Z(n20082) );
  XOR U19923 ( .A(n20084), .B(n20085), .Z(n20072) );
  AND U19924 ( .A(n20086), .B(n20087), .Z(n20085) );
  XOR U19925 ( .A(n20084), .B(n19211), .Z(n20087) );
  XOR U19926 ( .A(n20088), .B(n20089), .Z(n19211) );
  AND U19927 ( .A(n515), .B(n20090), .Z(n20089) );
  XOR U19928 ( .A(n20091), .B(n20088), .Z(n20090) );
  XNOR U19929 ( .A(n19208), .B(n20084), .Z(n20086) );
  XOR U19930 ( .A(n20092), .B(n20093), .Z(n19208) );
  AND U19931 ( .A(n512), .B(n20094), .Z(n20093) );
  XOR U19932 ( .A(n20095), .B(n20092), .Z(n20094) );
  XOR U19933 ( .A(n20096), .B(n20097), .Z(n20084) );
  AND U19934 ( .A(n20098), .B(n20099), .Z(n20097) );
  XOR U19935 ( .A(n20096), .B(n19223), .Z(n20099) );
  XOR U19936 ( .A(n20100), .B(n20101), .Z(n19223) );
  AND U19937 ( .A(n515), .B(n20102), .Z(n20101) );
  XOR U19938 ( .A(n20103), .B(n20100), .Z(n20102) );
  XNOR U19939 ( .A(n19220), .B(n20096), .Z(n20098) );
  XOR U19940 ( .A(n20104), .B(n20105), .Z(n19220) );
  AND U19941 ( .A(n512), .B(n20106), .Z(n20105) );
  XOR U19942 ( .A(n20107), .B(n20104), .Z(n20106) );
  XOR U19943 ( .A(n20108), .B(n20109), .Z(n20096) );
  AND U19944 ( .A(n20110), .B(n20111), .Z(n20109) );
  XOR U19945 ( .A(n20108), .B(n19235), .Z(n20111) );
  XOR U19946 ( .A(n20112), .B(n20113), .Z(n19235) );
  AND U19947 ( .A(n515), .B(n20114), .Z(n20113) );
  XOR U19948 ( .A(n20115), .B(n20112), .Z(n20114) );
  XNOR U19949 ( .A(n19232), .B(n20108), .Z(n20110) );
  XOR U19950 ( .A(n20116), .B(n20117), .Z(n19232) );
  AND U19951 ( .A(n512), .B(n20118), .Z(n20117) );
  XOR U19952 ( .A(n20119), .B(n20116), .Z(n20118) );
  XOR U19953 ( .A(n20120), .B(n20121), .Z(n20108) );
  AND U19954 ( .A(n20122), .B(n20123), .Z(n20121) );
  XOR U19955 ( .A(n20120), .B(n19247), .Z(n20123) );
  XOR U19956 ( .A(n20124), .B(n20125), .Z(n19247) );
  AND U19957 ( .A(n515), .B(n20126), .Z(n20125) );
  XOR U19958 ( .A(n20127), .B(n20124), .Z(n20126) );
  XNOR U19959 ( .A(n19244), .B(n20120), .Z(n20122) );
  XOR U19960 ( .A(n20128), .B(n20129), .Z(n19244) );
  AND U19961 ( .A(n512), .B(n20130), .Z(n20129) );
  XOR U19962 ( .A(n20131), .B(n20128), .Z(n20130) );
  XOR U19963 ( .A(n20132), .B(n20133), .Z(n20120) );
  AND U19964 ( .A(n20134), .B(n20135), .Z(n20133) );
  XOR U19965 ( .A(n20132), .B(n19259), .Z(n20135) );
  XOR U19966 ( .A(n20136), .B(n20137), .Z(n19259) );
  AND U19967 ( .A(n515), .B(n20138), .Z(n20137) );
  XOR U19968 ( .A(n20139), .B(n20136), .Z(n20138) );
  XNOR U19969 ( .A(n19256), .B(n20132), .Z(n20134) );
  XOR U19970 ( .A(n20140), .B(n20141), .Z(n19256) );
  AND U19971 ( .A(n512), .B(n20142), .Z(n20141) );
  XOR U19972 ( .A(n20143), .B(n20140), .Z(n20142) );
  XOR U19973 ( .A(n20144), .B(n20145), .Z(n20132) );
  AND U19974 ( .A(n20146), .B(n20147), .Z(n20145) );
  XOR U19975 ( .A(n20144), .B(n19271), .Z(n20147) );
  XOR U19976 ( .A(n20148), .B(n20149), .Z(n19271) );
  AND U19977 ( .A(n515), .B(n20150), .Z(n20149) );
  XOR U19978 ( .A(n20151), .B(n20148), .Z(n20150) );
  XNOR U19979 ( .A(n19268), .B(n20144), .Z(n20146) );
  XOR U19980 ( .A(n20152), .B(n20153), .Z(n19268) );
  AND U19981 ( .A(n512), .B(n20154), .Z(n20153) );
  XOR U19982 ( .A(n20155), .B(n20152), .Z(n20154) );
  XOR U19983 ( .A(n20156), .B(n20157), .Z(n20144) );
  AND U19984 ( .A(n20158), .B(n20159), .Z(n20157) );
  XOR U19985 ( .A(n20156), .B(n19283), .Z(n20159) );
  XOR U19986 ( .A(n20160), .B(n20161), .Z(n19283) );
  AND U19987 ( .A(n515), .B(n20162), .Z(n20161) );
  XOR U19988 ( .A(n20163), .B(n20160), .Z(n20162) );
  XNOR U19989 ( .A(n19280), .B(n20156), .Z(n20158) );
  XOR U19990 ( .A(n20164), .B(n20165), .Z(n19280) );
  AND U19991 ( .A(n512), .B(n20166), .Z(n20165) );
  XOR U19992 ( .A(n20167), .B(n20164), .Z(n20166) );
  XOR U19993 ( .A(n20168), .B(n20169), .Z(n20156) );
  AND U19994 ( .A(n20170), .B(n20171), .Z(n20169) );
  XOR U19995 ( .A(n20168), .B(n19295), .Z(n20171) );
  XOR U19996 ( .A(n20172), .B(n20173), .Z(n19295) );
  AND U19997 ( .A(n515), .B(n20174), .Z(n20173) );
  XOR U19998 ( .A(n20175), .B(n20172), .Z(n20174) );
  XNOR U19999 ( .A(n19292), .B(n20168), .Z(n20170) );
  XOR U20000 ( .A(n20176), .B(n20177), .Z(n19292) );
  AND U20001 ( .A(n512), .B(n20178), .Z(n20177) );
  XOR U20002 ( .A(n20179), .B(n20176), .Z(n20178) );
  XOR U20003 ( .A(n20180), .B(n20181), .Z(n20168) );
  AND U20004 ( .A(n20182), .B(n20183), .Z(n20181) );
  XOR U20005 ( .A(n20180), .B(n19307), .Z(n20183) );
  XOR U20006 ( .A(n20184), .B(n20185), .Z(n19307) );
  AND U20007 ( .A(n515), .B(n20186), .Z(n20185) );
  XOR U20008 ( .A(n20187), .B(n20184), .Z(n20186) );
  XNOR U20009 ( .A(n19304), .B(n20180), .Z(n20182) );
  XOR U20010 ( .A(n20188), .B(n20189), .Z(n19304) );
  AND U20011 ( .A(n512), .B(n20190), .Z(n20189) );
  XOR U20012 ( .A(n20191), .B(n20188), .Z(n20190) );
  XOR U20013 ( .A(n20192), .B(n20193), .Z(n20180) );
  AND U20014 ( .A(n20194), .B(n20195), .Z(n20193) );
  XOR U20015 ( .A(n20192), .B(n19319), .Z(n20195) );
  XOR U20016 ( .A(n20196), .B(n20197), .Z(n19319) );
  AND U20017 ( .A(n515), .B(n20198), .Z(n20197) );
  XOR U20018 ( .A(n20199), .B(n20196), .Z(n20198) );
  XNOR U20019 ( .A(n19316), .B(n20192), .Z(n20194) );
  XOR U20020 ( .A(n20200), .B(n20201), .Z(n19316) );
  AND U20021 ( .A(n512), .B(n20202), .Z(n20201) );
  XOR U20022 ( .A(n20203), .B(n20200), .Z(n20202) );
  XOR U20023 ( .A(n20204), .B(n20205), .Z(n20192) );
  AND U20024 ( .A(n20206), .B(n20207), .Z(n20205) );
  XOR U20025 ( .A(n20204), .B(n19331), .Z(n20207) );
  XOR U20026 ( .A(n20208), .B(n20209), .Z(n19331) );
  AND U20027 ( .A(n515), .B(n20210), .Z(n20209) );
  XOR U20028 ( .A(n20211), .B(n20208), .Z(n20210) );
  XNOR U20029 ( .A(n19328), .B(n20204), .Z(n20206) );
  XOR U20030 ( .A(n20212), .B(n20213), .Z(n19328) );
  AND U20031 ( .A(n512), .B(n20214), .Z(n20213) );
  XOR U20032 ( .A(n20215), .B(n20212), .Z(n20214) );
  XOR U20033 ( .A(n20216), .B(n20217), .Z(n20204) );
  AND U20034 ( .A(n20218), .B(n20219), .Z(n20217) );
  XNOR U20035 ( .A(n20220), .B(n19344), .Z(n20219) );
  XOR U20036 ( .A(n20221), .B(n20222), .Z(n19344) );
  AND U20037 ( .A(n515), .B(n20223), .Z(n20222) );
  XOR U20038 ( .A(n20221), .B(n20224), .Z(n20223) );
  XNOR U20039 ( .A(n19341), .B(n20216), .Z(n20218) );
  XOR U20040 ( .A(n20225), .B(n20226), .Z(n19341) );
  AND U20041 ( .A(n512), .B(n20227), .Z(n20226) );
  XOR U20042 ( .A(n20225), .B(n20228), .Z(n20227) );
  IV U20043 ( .A(n20220), .Z(n20216) );
  AND U20044 ( .A(n20048), .B(n20051), .Z(n20220) );
  XNOR U20045 ( .A(n20229), .B(n20230), .Z(n20051) );
  AND U20046 ( .A(n515), .B(n20231), .Z(n20230) );
  XNOR U20047 ( .A(n20232), .B(n20229), .Z(n20231) );
  XOR U20048 ( .A(n20233), .B(n20234), .Z(n515) );
  AND U20049 ( .A(n20235), .B(n20236), .Z(n20234) );
  XNOR U20050 ( .A(n20056), .B(n20233), .Z(n20236) );
  AND U20051 ( .A(p_input[1407]), .B(p_input[1391]), .Z(n20056) );
  XOR U20052 ( .A(n20233), .B(n20057), .Z(n20235) );
  AND U20053 ( .A(p_input[1375]), .B(p_input[1359]), .Z(n20057) );
  XOR U20054 ( .A(n20237), .B(n20238), .Z(n20233) );
  AND U20055 ( .A(n20239), .B(n20240), .Z(n20238) );
  XOR U20056 ( .A(n20237), .B(n20067), .Z(n20240) );
  XNOR U20057 ( .A(p_input[1390]), .B(n20241), .Z(n20067) );
  AND U20058 ( .A(n683), .B(n20242), .Z(n20241) );
  XOR U20059 ( .A(p_input[1406]), .B(p_input[1390]), .Z(n20242) );
  XNOR U20060 ( .A(n20064), .B(n20237), .Z(n20239) );
  XOR U20061 ( .A(n20243), .B(n20244), .Z(n20064) );
  AND U20062 ( .A(n681), .B(n20245), .Z(n20244) );
  XOR U20063 ( .A(p_input[1374]), .B(p_input[1358]), .Z(n20245) );
  XOR U20064 ( .A(n20246), .B(n20247), .Z(n20237) );
  AND U20065 ( .A(n20248), .B(n20249), .Z(n20247) );
  XOR U20066 ( .A(n20246), .B(n20079), .Z(n20249) );
  XNOR U20067 ( .A(p_input[1389]), .B(n20250), .Z(n20079) );
  AND U20068 ( .A(n683), .B(n20251), .Z(n20250) );
  XOR U20069 ( .A(p_input[1405]), .B(p_input[1389]), .Z(n20251) );
  XNOR U20070 ( .A(n20076), .B(n20246), .Z(n20248) );
  XOR U20071 ( .A(n20252), .B(n20253), .Z(n20076) );
  AND U20072 ( .A(n681), .B(n20254), .Z(n20253) );
  XOR U20073 ( .A(p_input[1373]), .B(p_input[1357]), .Z(n20254) );
  XOR U20074 ( .A(n20255), .B(n20256), .Z(n20246) );
  AND U20075 ( .A(n20257), .B(n20258), .Z(n20256) );
  XOR U20076 ( .A(n20255), .B(n20091), .Z(n20258) );
  XNOR U20077 ( .A(p_input[1388]), .B(n20259), .Z(n20091) );
  AND U20078 ( .A(n683), .B(n20260), .Z(n20259) );
  XOR U20079 ( .A(p_input[1404]), .B(p_input[1388]), .Z(n20260) );
  XNOR U20080 ( .A(n20088), .B(n20255), .Z(n20257) );
  XOR U20081 ( .A(n20261), .B(n20262), .Z(n20088) );
  AND U20082 ( .A(n681), .B(n20263), .Z(n20262) );
  XOR U20083 ( .A(p_input[1372]), .B(p_input[1356]), .Z(n20263) );
  XOR U20084 ( .A(n20264), .B(n20265), .Z(n20255) );
  AND U20085 ( .A(n20266), .B(n20267), .Z(n20265) );
  XOR U20086 ( .A(n20264), .B(n20103), .Z(n20267) );
  XNOR U20087 ( .A(p_input[1387]), .B(n20268), .Z(n20103) );
  AND U20088 ( .A(n683), .B(n20269), .Z(n20268) );
  XOR U20089 ( .A(p_input[1403]), .B(p_input[1387]), .Z(n20269) );
  XNOR U20090 ( .A(n20100), .B(n20264), .Z(n20266) );
  XOR U20091 ( .A(n20270), .B(n20271), .Z(n20100) );
  AND U20092 ( .A(n681), .B(n20272), .Z(n20271) );
  XOR U20093 ( .A(p_input[1371]), .B(p_input[1355]), .Z(n20272) );
  XOR U20094 ( .A(n20273), .B(n20274), .Z(n20264) );
  AND U20095 ( .A(n20275), .B(n20276), .Z(n20274) );
  XOR U20096 ( .A(n20273), .B(n20115), .Z(n20276) );
  XNOR U20097 ( .A(p_input[1386]), .B(n20277), .Z(n20115) );
  AND U20098 ( .A(n683), .B(n20278), .Z(n20277) );
  XOR U20099 ( .A(p_input[1402]), .B(p_input[1386]), .Z(n20278) );
  XNOR U20100 ( .A(n20112), .B(n20273), .Z(n20275) );
  XOR U20101 ( .A(n20279), .B(n20280), .Z(n20112) );
  AND U20102 ( .A(n681), .B(n20281), .Z(n20280) );
  XOR U20103 ( .A(p_input[1370]), .B(p_input[1354]), .Z(n20281) );
  XOR U20104 ( .A(n20282), .B(n20283), .Z(n20273) );
  AND U20105 ( .A(n20284), .B(n20285), .Z(n20283) );
  XOR U20106 ( .A(n20282), .B(n20127), .Z(n20285) );
  XNOR U20107 ( .A(p_input[1385]), .B(n20286), .Z(n20127) );
  AND U20108 ( .A(n683), .B(n20287), .Z(n20286) );
  XOR U20109 ( .A(p_input[1401]), .B(p_input[1385]), .Z(n20287) );
  XNOR U20110 ( .A(n20124), .B(n20282), .Z(n20284) );
  XOR U20111 ( .A(n20288), .B(n20289), .Z(n20124) );
  AND U20112 ( .A(n681), .B(n20290), .Z(n20289) );
  XOR U20113 ( .A(p_input[1369]), .B(p_input[1353]), .Z(n20290) );
  XOR U20114 ( .A(n20291), .B(n20292), .Z(n20282) );
  AND U20115 ( .A(n20293), .B(n20294), .Z(n20292) );
  XOR U20116 ( .A(n20291), .B(n20139), .Z(n20294) );
  XNOR U20117 ( .A(p_input[1384]), .B(n20295), .Z(n20139) );
  AND U20118 ( .A(n683), .B(n20296), .Z(n20295) );
  XOR U20119 ( .A(p_input[1400]), .B(p_input[1384]), .Z(n20296) );
  XNOR U20120 ( .A(n20136), .B(n20291), .Z(n20293) );
  XOR U20121 ( .A(n20297), .B(n20298), .Z(n20136) );
  AND U20122 ( .A(n681), .B(n20299), .Z(n20298) );
  XOR U20123 ( .A(p_input[1368]), .B(p_input[1352]), .Z(n20299) );
  XOR U20124 ( .A(n20300), .B(n20301), .Z(n20291) );
  AND U20125 ( .A(n20302), .B(n20303), .Z(n20301) );
  XOR U20126 ( .A(n20300), .B(n20151), .Z(n20303) );
  XNOR U20127 ( .A(p_input[1383]), .B(n20304), .Z(n20151) );
  AND U20128 ( .A(n683), .B(n20305), .Z(n20304) );
  XOR U20129 ( .A(p_input[1399]), .B(p_input[1383]), .Z(n20305) );
  XNOR U20130 ( .A(n20148), .B(n20300), .Z(n20302) );
  XOR U20131 ( .A(n20306), .B(n20307), .Z(n20148) );
  AND U20132 ( .A(n681), .B(n20308), .Z(n20307) );
  XOR U20133 ( .A(p_input[1367]), .B(p_input[1351]), .Z(n20308) );
  XOR U20134 ( .A(n20309), .B(n20310), .Z(n20300) );
  AND U20135 ( .A(n20311), .B(n20312), .Z(n20310) );
  XOR U20136 ( .A(n20309), .B(n20163), .Z(n20312) );
  XNOR U20137 ( .A(p_input[1382]), .B(n20313), .Z(n20163) );
  AND U20138 ( .A(n683), .B(n20314), .Z(n20313) );
  XOR U20139 ( .A(p_input[1398]), .B(p_input[1382]), .Z(n20314) );
  XNOR U20140 ( .A(n20160), .B(n20309), .Z(n20311) );
  XOR U20141 ( .A(n20315), .B(n20316), .Z(n20160) );
  AND U20142 ( .A(n681), .B(n20317), .Z(n20316) );
  XOR U20143 ( .A(p_input[1366]), .B(p_input[1350]), .Z(n20317) );
  XOR U20144 ( .A(n20318), .B(n20319), .Z(n20309) );
  AND U20145 ( .A(n20320), .B(n20321), .Z(n20319) );
  XOR U20146 ( .A(n20318), .B(n20175), .Z(n20321) );
  XNOR U20147 ( .A(p_input[1381]), .B(n20322), .Z(n20175) );
  AND U20148 ( .A(n683), .B(n20323), .Z(n20322) );
  XOR U20149 ( .A(p_input[1397]), .B(p_input[1381]), .Z(n20323) );
  XNOR U20150 ( .A(n20172), .B(n20318), .Z(n20320) );
  XOR U20151 ( .A(n20324), .B(n20325), .Z(n20172) );
  AND U20152 ( .A(n681), .B(n20326), .Z(n20325) );
  XOR U20153 ( .A(p_input[1365]), .B(p_input[1349]), .Z(n20326) );
  XOR U20154 ( .A(n20327), .B(n20328), .Z(n20318) );
  AND U20155 ( .A(n20329), .B(n20330), .Z(n20328) );
  XOR U20156 ( .A(n20327), .B(n20187), .Z(n20330) );
  XNOR U20157 ( .A(p_input[1380]), .B(n20331), .Z(n20187) );
  AND U20158 ( .A(n683), .B(n20332), .Z(n20331) );
  XOR U20159 ( .A(p_input[1396]), .B(p_input[1380]), .Z(n20332) );
  XNOR U20160 ( .A(n20184), .B(n20327), .Z(n20329) );
  XOR U20161 ( .A(n20333), .B(n20334), .Z(n20184) );
  AND U20162 ( .A(n681), .B(n20335), .Z(n20334) );
  XOR U20163 ( .A(p_input[1364]), .B(p_input[1348]), .Z(n20335) );
  XOR U20164 ( .A(n20336), .B(n20337), .Z(n20327) );
  AND U20165 ( .A(n20338), .B(n20339), .Z(n20337) );
  XOR U20166 ( .A(n20336), .B(n20199), .Z(n20339) );
  XNOR U20167 ( .A(p_input[1379]), .B(n20340), .Z(n20199) );
  AND U20168 ( .A(n683), .B(n20341), .Z(n20340) );
  XOR U20169 ( .A(p_input[1395]), .B(p_input[1379]), .Z(n20341) );
  XNOR U20170 ( .A(n20196), .B(n20336), .Z(n20338) );
  XOR U20171 ( .A(n20342), .B(n20343), .Z(n20196) );
  AND U20172 ( .A(n681), .B(n20344), .Z(n20343) );
  XOR U20173 ( .A(p_input[1363]), .B(p_input[1347]), .Z(n20344) );
  XOR U20174 ( .A(n20345), .B(n20346), .Z(n20336) );
  AND U20175 ( .A(n20347), .B(n20348), .Z(n20346) );
  XOR U20176 ( .A(n20345), .B(n20211), .Z(n20348) );
  XNOR U20177 ( .A(p_input[1378]), .B(n20349), .Z(n20211) );
  AND U20178 ( .A(n683), .B(n20350), .Z(n20349) );
  XOR U20179 ( .A(p_input[1394]), .B(p_input[1378]), .Z(n20350) );
  XNOR U20180 ( .A(n20208), .B(n20345), .Z(n20347) );
  XOR U20181 ( .A(n20351), .B(n20352), .Z(n20208) );
  AND U20182 ( .A(n681), .B(n20353), .Z(n20352) );
  XOR U20183 ( .A(p_input[1362]), .B(p_input[1346]), .Z(n20353) );
  XOR U20184 ( .A(n20354), .B(n20355), .Z(n20345) );
  AND U20185 ( .A(n20356), .B(n20357), .Z(n20355) );
  XNOR U20186 ( .A(n20358), .B(n20224), .Z(n20357) );
  XNOR U20187 ( .A(p_input[1377]), .B(n20359), .Z(n20224) );
  AND U20188 ( .A(n683), .B(n20360), .Z(n20359) );
  XNOR U20189 ( .A(p_input[1393]), .B(n20361), .Z(n20360) );
  IV U20190 ( .A(p_input[1377]), .Z(n20361) );
  XNOR U20191 ( .A(n20221), .B(n20354), .Z(n20356) );
  XNOR U20192 ( .A(p_input[1345]), .B(n20362), .Z(n20221) );
  AND U20193 ( .A(n681), .B(n20363), .Z(n20362) );
  XOR U20194 ( .A(p_input[1361]), .B(p_input[1345]), .Z(n20363) );
  IV U20195 ( .A(n20358), .Z(n20354) );
  AND U20196 ( .A(n20229), .B(n20232), .Z(n20358) );
  XOR U20197 ( .A(p_input[1376]), .B(n20364), .Z(n20232) );
  AND U20198 ( .A(n683), .B(n20365), .Z(n20364) );
  XOR U20199 ( .A(p_input[1392]), .B(p_input[1376]), .Z(n20365) );
  XOR U20200 ( .A(n20366), .B(n20367), .Z(n683) );
  AND U20201 ( .A(n20368), .B(n20369), .Z(n20367) );
  XNOR U20202 ( .A(p_input[1407]), .B(n20366), .Z(n20369) );
  XOR U20203 ( .A(n20366), .B(p_input[1391]), .Z(n20368) );
  XOR U20204 ( .A(n20370), .B(n20371), .Z(n20366) );
  AND U20205 ( .A(n20372), .B(n20373), .Z(n20371) );
  XNOR U20206 ( .A(p_input[1406]), .B(n20370), .Z(n20373) );
  XOR U20207 ( .A(n20370), .B(p_input[1390]), .Z(n20372) );
  XOR U20208 ( .A(n20374), .B(n20375), .Z(n20370) );
  AND U20209 ( .A(n20376), .B(n20377), .Z(n20375) );
  XNOR U20210 ( .A(p_input[1405]), .B(n20374), .Z(n20377) );
  XOR U20211 ( .A(n20374), .B(p_input[1389]), .Z(n20376) );
  XOR U20212 ( .A(n20378), .B(n20379), .Z(n20374) );
  AND U20213 ( .A(n20380), .B(n20381), .Z(n20379) );
  XNOR U20214 ( .A(p_input[1404]), .B(n20378), .Z(n20381) );
  XOR U20215 ( .A(n20378), .B(p_input[1388]), .Z(n20380) );
  XOR U20216 ( .A(n20382), .B(n20383), .Z(n20378) );
  AND U20217 ( .A(n20384), .B(n20385), .Z(n20383) );
  XNOR U20218 ( .A(p_input[1403]), .B(n20382), .Z(n20385) );
  XOR U20219 ( .A(n20382), .B(p_input[1387]), .Z(n20384) );
  XOR U20220 ( .A(n20386), .B(n20387), .Z(n20382) );
  AND U20221 ( .A(n20388), .B(n20389), .Z(n20387) );
  XNOR U20222 ( .A(p_input[1402]), .B(n20386), .Z(n20389) );
  XOR U20223 ( .A(n20386), .B(p_input[1386]), .Z(n20388) );
  XOR U20224 ( .A(n20390), .B(n20391), .Z(n20386) );
  AND U20225 ( .A(n20392), .B(n20393), .Z(n20391) );
  XNOR U20226 ( .A(p_input[1401]), .B(n20390), .Z(n20393) );
  XOR U20227 ( .A(n20390), .B(p_input[1385]), .Z(n20392) );
  XOR U20228 ( .A(n20394), .B(n20395), .Z(n20390) );
  AND U20229 ( .A(n20396), .B(n20397), .Z(n20395) );
  XNOR U20230 ( .A(p_input[1400]), .B(n20394), .Z(n20397) );
  XOR U20231 ( .A(n20394), .B(p_input[1384]), .Z(n20396) );
  XOR U20232 ( .A(n20398), .B(n20399), .Z(n20394) );
  AND U20233 ( .A(n20400), .B(n20401), .Z(n20399) );
  XNOR U20234 ( .A(p_input[1399]), .B(n20398), .Z(n20401) );
  XOR U20235 ( .A(n20398), .B(p_input[1383]), .Z(n20400) );
  XOR U20236 ( .A(n20402), .B(n20403), .Z(n20398) );
  AND U20237 ( .A(n20404), .B(n20405), .Z(n20403) );
  XNOR U20238 ( .A(p_input[1398]), .B(n20402), .Z(n20405) );
  XOR U20239 ( .A(n20402), .B(p_input[1382]), .Z(n20404) );
  XOR U20240 ( .A(n20406), .B(n20407), .Z(n20402) );
  AND U20241 ( .A(n20408), .B(n20409), .Z(n20407) );
  XNOR U20242 ( .A(p_input[1397]), .B(n20406), .Z(n20409) );
  XOR U20243 ( .A(n20406), .B(p_input[1381]), .Z(n20408) );
  XOR U20244 ( .A(n20410), .B(n20411), .Z(n20406) );
  AND U20245 ( .A(n20412), .B(n20413), .Z(n20411) );
  XNOR U20246 ( .A(p_input[1396]), .B(n20410), .Z(n20413) );
  XOR U20247 ( .A(n20410), .B(p_input[1380]), .Z(n20412) );
  XOR U20248 ( .A(n20414), .B(n20415), .Z(n20410) );
  AND U20249 ( .A(n20416), .B(n20417), .Z(n20415) );
  XNOR U20250 ( .A(p_input[1395]), .B(n20414), .Z(n20417) );
  XOR U20251 ( .A(n20414), .B(p_input[1379]), .Z(n20416) );
  XOR U20252 ( .A(n20418), .B(n20419), .Z(n20414) );
  AND U20253 ( .A(n20420), .B(n20421), .Z(n20419) );
  XNOR U20254 ( .A(p_input[1394]), .B(n20418), .Z(n20421) );
  XOR U20255 ( .A(n20418), .B(p_input[1378]), .Z(n20420) );
  XNOR U20256 ( .A(n20422), .B(n20423), .Z(n20418) );
  AND U20257 ( .A(n20424), .B(n20425), .Z(n20423) );
  XOR U20258 ( .A(p_input[1393]), .B(n20422), .Z(n20425) );
  XNOR U20259 ( .A(p_input[1377]), .B(n20422), .Z(n20424) );
  AND U20260 ( .A(p_input[1392]), .B(n20426), .Z(n20422) );
  IV U20261 ( .A(p_input[1376]), .Z(n20426) );
  XNOR U20262 ( .A(p_input[1344]), .B(n20427), .Z(n20229) );
  AND U20263 ( .A(n681), .B(n20428), .Z(n20427) );
  XOR U20264 ( .A(p_input[1360]), .B(p_input[1344]), .Z(n20428) );
  XOR U20265 ( .A(n20429), .B(n20430), .Z(n681) );
  AND U20266 ( .A(n20431), .B(n20432), .Z(n20430) );
  XNOR U20267 ( .A(p_input[1375]), .B(n20429), .Z(n20432) );
  XOR U20268 ( .A(n20429), .B(p_input[1359]), .Z(n20431) );
  XOR U20269 ( .A(n20433), .B(n20434), .Z(n20429) );
  AND U20270 ( .A(n20435), .B(n20436), .Z(n20434) );
  XNOR U20271 ( .A(p_input[1374]), .B(n20433), .Z(n20436) );
  XNOR U20272 ( .A(n20433), .B(n20243), .Z(n20435) );
  IV U20273 ( .A(p_input[1358]), .Z(n20243) );
  XOR U20274 ( .A(n20437), .B(n20438), .Z(n20433) );
  AND U20275 ( .A(n20439), .B(n20440), .Z(n20438) );
  XNOR U20276 ( .A(p_input[1373]), .B(n20437), .Z(n20440) );
  XNOR U20277 ( .A(n20437), .B(n20252), .Z(n20439) );
  IV U20278 ( .A(p_input[1357]), .Z(n20252) );
  XOR U20279 ( .A(n20441), .B(n20442), .Z(n20437) );
  AND U20280 ( .A(n20443), .B(n20444), .Z(n20442) );
  XNOR U20281 ( .A(p_input[1372]), .B(n20441), .Z(n20444) );
  XNOR U20282 ( .A(n20441), .B(n20261), .Z(n20443) );
  IV U20283 ( .A(p_input[1356]), .Z(n20261) );
  XOR U20284 ( .A(n20445), .B(n20446), .Z(n20441) );
  AND U20285 ( .A(n20447), .B(n20448), .Z(n20446) );
  XNOR U20286 ( .A(p_input[1371]), .B(n20445), .Z(n20448) );
  XNOR U20287 ( .A(n20445), .B(n20270), .Z(n20447) );
  IV U20288 ( .A(p_input[1355]), .Z(n20270) );
  XOR U20289 ( .A(n20449), .B(n20450), .Z(n20445) );
  AND U20290 ( .A(n20451), .B(n20452), .Z(n20450) );
  XNOR U20291 ( .A(p_input[1370]), .B(n20449), .Z(n20452) );
  XNOR U20292 ( .A(n20449), .B(n20279), .Z(n20451) );
  IV U20293 ( .A(p_input[1354]), .Z(n20279) );
  XOR U20294 ( .A(n20453), .B(n20454), .Z(n20449) );
  AND U20295 ( .A(n20455), .B(n20456), .Z(n20454) );
  XNOR U20296 ( .A(p_input[1369]), .B(n20453), .Z(n20456) );
  XNOR U20297 ( .A(n20453), .B(n20288), .Z(n20455) );
  IV U20298 ( .A(p_input[1353]), .Z(n20288) );
  XOR U20299 ( .A(n20457), .B(n20458), .Z(n20453) );
  AND U20300 ( .A(n20459), .B(n20460), .Z(n20458) );
  XNOR U20301 ( .A(p_input[1368]), .B(n20457), .Z(n20460) );
  XNOR U20302 ( .A(n20457), .B(n20297), .Z(n20459) );
  IV U20303 ( .A(p_input[1352]), .Z(n20297) );
  XOR U20304 ( .A(n20461), .B(n20462), .Z(n20457) );
  AND U20305 ( .A(n20463), .B(n20464), .Z(n20462) );
  XNOR U20306 ( .A(p_input[1367]), .B(n20461), .Z(n20464) );
  XNOR U20307 ( .A(n20461), .B(n20306), .Z(n20463) );
  IV U20308 ( .A(p_input[1351]), .Z(n20306) );
  XOR U20309 ( .A(n20465), .B(n20466), .Z(n20461) );
  AND U20310 ( .A(n20467), .B(n20468), .Z(n20466) );
  XNOR U20311 ( .A(p_input[1366]), .B(n20465), .Z(n20468) );
  XNOR U20312 ( .A(n20465), .B(n20315), .Z(n20467) );
  IV U20313 ( .A(p_input[1350]), .Z(n20315) );
  XOR U20314 ( .A(n20469), .B(n20470), .Z(n20465) );
  AND U20315 ( .A(n20471), .B(n20472), .Z(n20470) );
  XNOR U20316 ( .A(p_input[1365]), .B(n20469), .Z(n20472) );
  XNOR U20317 ( .A(n20469), .B(n20324), .Z(n20471) );
  IV U20318 ( .A(p_input[1349]), .Z(n20324) );
  XOR U20319 ( .A(n20473), .B(n20474), .Z(n20469) );
  AND U20320 ( .A(n20475), .B(n20476), .Z(n20474) );
  XNOR U20321 ( .A(p_input[1364]), .B(n20473), .Z(n20476) );
  XNOR U20322 ( .A(n20473), .B(n20333), .Z(n20475) );
  IV U20323 ( .A(p_input[1348]), .Z(n20333) );
  XOR U20324 ( .A(n20477), .B(n20478), .Z(n20473) );
  AND U20325 ( .A(n20479), .B(n20480), .Z(n20478) );
  XNOR U20326 ( .A(p_input[1363]), .B(n20477), .Z(n20480) );
  XNOR U20327 ( .A(n20477), .B(n20342), .Z(n20479) );
  IV U20328 ( .A(p_input[1347]), .Z(n20342) );
  XOR U20329 ( .A(n20481), .B(n20482), .Z(n20477) );
  AND U20330 ( .A(n20483), .B(n20484), .Z(n20482) );
  XNOR U20331 ( .A(p_input[1362]), .B(n20481), .Z(n20484) );
  XNOR U20332 ( .A(n20481), .B(n20351), .Z(n20483) );
  IV U20333 ( .A(p_input[1346]), .Z(n20351) );
  XNOR U20334 ( .A(n20485), .B(n20486), .Z(n20481) );
  AND U20335 ( .A(n20487), .B(n20488), .Z(n20486) );
  XOR U20336 ( .A(p_input[1361]), .B(n20485), .Z(n20488) );
  XNOR U20337 ( .A(p_input[1345]), .B(n20485), .Z(n20487) );
  AND U20338 ( .A(p_input[1360]), .B(n20489), .Z(n20485) );
  IV U20339 ( .A(p_input[1344]), .Z(n20489) );
  XOR U20340 ( .A(n20490), .B(n20491), .Z(n20048) );
  AND U20341 ( .A(n512), .B(n20492), .Z(n20491) );
  XNOR U20342 ( .A(n20493), .B(n20490), .Z(n20492) );
  XOR U20343 ( .A(n20494), .B(n20495), .Z(n512) );
  AND U20344 ( .A(n20496), .B(n20497), .Z(n20495) );
  XNOR U20345 ( .A(n20059), .B(n20494), .Z(n20497) );
  AND U20346 ( .A(p_input[1343]), .B(p_input[1327]), .Z(n20059) );
  XOR U20347 ( .A(n20494), .B(n20058), .Z(n20496) );
  AND U20348 ( .A(p_input[1295]), .B(p_input[1311]), .Z(n20058) );
  XOR U20349 ( .A(n20498), .B(n20499), .Z(n20494) );
  AND U20350 ( .A(n20500), .B(n20501), .Z(n20499) );
  XOR U20351 ( .A(n20498), .B(n20071), .Z(n20501) );
  XNOR U20352 ( .A(p_input[1326]), .B(n20502), .Z(n20071) );
  AND U20353 ( .A(n687), .B(n20503), .Z(n20502) );
  XOR U20354 ( .A(p_input[1342]), .B(p_input[1326]), .Z(n20503) );
  XNOR U20355 ( .A(n20068), .B(n20498), .Z(n20500) );
  XOR U20356 ( .A(n20504), .B(n20505), .Z(n20068) );
  AND U20357 ( .A(n684), .B(n20506), .Z(n20505) );
  XOR U20358 ( .A(p_input[1310]), .B(p_input[1294]), .Z(n20506) );
  XOR U20359 ( .A(n20507), .B(n20508), .Z(n20498) );
  AND U20360 ( .A(n20509), .B(n20510), .Z(n20508) );
  XOR U20361 ( .A(n20507), .B(n20083), .Z(n20510) );
  XNOR U20362 ( .A(p_input[1325]), .B(n20511), .Z(n20083) );
  AND U20363 ( .A(n687), .B(n20512), .Z(n20511) );
  XOR U20364 ( .A(p_input[1341]), .B(p_input[1325]), .Z(n20512) );
  XNOR U20365 ( .A(n20080), .B(n20507), .Z(n20509) );
  XOR U20366 ( .A(n20513), .B(n20514), .Z(n20080) );
  AND U20367 ( .A(n684), .B(n20515), .Z(n20514) );
  XOR U20368 ( .A(p_input[1309]), .B(p_input[1293]), .Z(n20515) );
  XOR U20369 ( .A(n20516), .B(n20517), .Z(n20507) );
  AND U20370 ( .A(n20518), .B(n20519), .Z(n20517) );
  XOR U20371 ( .A(n20516), .B(n20095), .Z(n20519) );
  XNOR U20372 ( .A(p_input[1324]), .B(n20520), .Z(n20095) );
  AND U20373 ( .A(n687), .B(n20521), .Z(n20520) );
  XOR U20374 ( .A(p_input[1340]), .B(p_input[1324]), .Z(n20521) );
  XNOR U20375 ( .A(n20092), .B(n20516), .Z(n20518) );
  XOR U20376 ( .A(n20522), .B(n20523), .Z(n20092) );
  AND U20377 ( .A(n684), .B(n20524), .Z(n20523) );
  XOR U20378 ( .A(p_input[1308]), .B(p_input[1292]), .Z(n20524) );
  XOR U20379 ( .A(n20525), .B(n20526), .Z(n20516) );
  AND U20380 ( .A(n20527), .B(n20528), .Z(n20526) );
  XOR U20381 ( .A(n20525), .B(n20107), .Z(n20528) );
  XNOR U20382 ( .A(p_input[1323]), .B(n20529), .Z(n20107) );
  AND U20383 ( .A(n687), .B(n20530), .Z(n20529) );
  XOR U20384 ( .A(p_input[1339]), .B(p_input[1323]), .Z(n20530) );
  XNOR U20385 ( .A(n20104), .B(n20525), .Z(n20527) );
  XOR U20386 ( .A(n20531), .B(n20532), .Z(n20104) );
  AND U20387 ( .A(n684), .B(n20533), .Z(n20532) );
  XOR U20388 ( .A(p_input[1307]), .B(p_input[1291]), .Z(n20533) );
  XOR U20389 ( .A(n20534), .B(n20535), .Z(n20525) );
  AND U20390 ( .A(n20536), .B(n20537), .Z(n20535) );
  XOR U20391 ( .A(n20534), .B(n20119), .Z(n20537) );
  XNOR U20392 ( .A(p_input[1322]), .B(n20538), .Z(n20119) );
  AND U20393 ( .A(n687), .B(n20539), .Z(n20538) );
  XOR U20394 ( .A(p_input[1338]), .B(p_input[1322]), .Z(n20539) );
  XNOR U20395 ( .A(n20116), .B(n20534), .Z(n20536) );
  XOR U20396 ( .A(n20540), .B(n20541), .Z(n20116) );
  AND U20397 ( .A(n684), .B(n20542), .Z(n20541) );
  XOR U20398 ( .A(p_input[1306]), .B(p_input[1290]), .Z(n20542) );
  XOR U20399 ( .A(n20543), .B(n20544), .Z(n20534) );
  AND U20400 ( .A(n20545), .B(n20546), .Z(n20544) );
  XOR U20401 ( .A(n20543), .B(n20131), .Z(n20546) );
  XNOR U20402 ( .A(p_input[1321]), .B(n20547), .Z(n20131) );
  AND U20403 ( .A(n687), .B(n20548), .Z(n20547) );
  XOR U20404 ( .A(p_input[1337]), .B(p_input[1321]), .Z(n20548) );
  XNOR U20405 ( .A(n20128), .B(n20543), .Z(n20545) );
  XOR U20406 ( .A(n20549), .B(n20550), .Z(n20128) );
  AND U20407 ( .A(n684), .B(n20551), .Z(n20550) );
  XOR U20408 ( .A(p_input[1305]), .B(p_input[1289]), .Z(n20551) );
  XOR U20409 ( .A(n20552), .B(n20553), .Z(n20543) );
  AND U20410 ( .A(n20554), .B(n20555), .Z(n20553) );
  XOR U20411 ( .A(n20552), .B(n20143), .Z(n20555) );
  XNOR U20412 ( .A(p_input[1320]), .B(n20556), .Z(n20143) );
  AND U20413 ( .A(n687), .B(n20557), .Z(n20556) );
  XOR U20414 ( .A(p_input[1336]), .B(p_input[1320]), .Z(n20557) );
  XNOR U20415 ( .A(n20140), .B(n20552), .Z(n20554) );
  XOR U20416 ( .A(n20558), .B(n20559), .Z(n20140) );
  AND U20417 ( .A(n684), .B(n20560), .Z(n20559) );
  XOR U20418 ( .A(p_input[1304]), .B(p_input[1288]), .Z(n20560) );
  XOR U20419 ( .A(n20561), .B(n20562), .Z(n20552) );
  AND U20420 ( .A(n20563), .B(n20564), .Z(n20562) );
  XOR U20421 ( .A(n20561), .B(n20155), .Z(n20564) );
  XNOR U20422 ( .A(p_input[1319]), .B(n20565), .Z(n20155) );
  AND U20423 ( .A(n687), .B(n20566), .Z(n20565) );
  XOR U20424 ( .A(p_input[1335]), .B(p_input[1319]), .Z(n20566) );
  XNOR U20425 ( .A(n20152), .B(n20561), .Z(n20563) );
  XOR U20426 ( .A(n20567), .B(n20568), .Z(n20152) );
  AND U20427 ( .A(n684), .B(n20569), .Z(n20568) );
  XOR U20428 ( .A(p_input[1303]), .B(p_input[1287]), .Z(n20569) );
  XOR U20429 ( .A(n20570), .B(n20571), .Z(n20561) );
  AND U20430 ( .A(n20572), .B(n20573), .Z(n20571) );
  XOR U20431 ( .A(n20570), .B(n20167), .Z(n20573) );
  XNOR U20432 ( .A(p_input[1318]), .B(n20574), .Z(n20167) );
  AND U20433 ( .A(n687), .B(n20575), .Z(n20574) );
  XOR U20434 ( .A(p_input[1334]), .B(p_input[1318]), .Z(n20575) );
  XNOR U20435 ( .A(n20164), .B(n20570), .Z(n20572) );
  XOR U20436 ( .A(n20576), .B(n20577), .Z(n20164) );
  AND U20437 ( .A(n684), .B(n20578), .Z(n20577) );
  XOR U20438 ( .A(p_input[1302]), .B(p_input[1286]), .Z(n20578) );
  XOR U20439 ( .A(n20579), .B(n20580), .Z(n20570) );
  AND U20440 ( .A(n20581), .B(n20582), .Z(n20580) );
  XOR U20441 ( .A(n20579), .B(n20179), .Z(n20582) );
  XNOR U20442 ( .A(p_input[1317]), .B(n20583), .Z(n20179) );
  AND U20443 ( .A(n687), .B(n20584), .Z(n20583) );
  XOR U20444 ( .A(p_input[1333]), .B(p_input[1317]), .Z(n20584) );
  XNOR U20445 ( .A(n20176), .B(n20579), .Z(n20581) );
  XOR U20446 ( .A(n20585), .B(n20586), .Z(n20176) );
  AND U20447 ( .A(n684), .B(n20587), .Z(n20586) );
  XOR U20448 ( .A(p_input[1301]), .B(p_input[1285]), .Z(n20587) );
  XOR U20449 ( .A(n20588), .B(n20589), .Z(n20579) );
  AND U20450 ( .A(n20590), .B(n20591), .Z(n20589) );
  XOR U20451 ( .A(n20588), .B(n20191), .Z(n20591) );
  XNOR U20452 ( .A(p_input[1316]), .B(n20592), .Z(n20191) );
  AND U20453 ( .A(n687), .B(n20593), .Z(n20592) );
  XOR U20454 ( .A(p_input[1332]), .B(p_input[1316]), .Z(n20593) );
  XNOR U20455 ( .A(n20188), .B(n20588), .Z(n20590) );
  XOR U20456 ( .A(n20594), .B(n20595), .Z(n20188) );
  AND U20457 ( .A(n684), .B(n20596), .Z(n20595) );
  XOR U20458 ( .A(p_input[1300]), .B(p_input[1284]), .Z(n20596) );
  XOR U20459 ( .A(n20597), .B(n20598), .Z(n20588) );
  AND U20460 ( .A(n20599), .B(n20600), .Z(n20598) );
  XOR U20461 ( .A(n20597), .B(n20203), .Z(n20600) );
  XNOR U20462 ( .A(p_input[1315]), .B(n20601), .Z(n20203) );
  AND U20463 ( .A(n687), .B(n20602), .Z(n20601) );
  XOR U20464 ( .A(p_input[1331]), .B(p_input[1315]), .Z(n20602) );
  XNOR U20465 ( .A(n20200), .B(n20597), .Z(n20599) );
  XOR U20466 ( .A(n20603), .B(n20604), .Z(n20200) );
  AND U20467 ( .A(n684), .B(n20605), .Z(n20604) );
  XOR U20468 ( .A(p_input[1299]), .B(p_input[1283]), .Z(n20605) );
  XOR U20469 ( .A(n20606), .B(n20607), .Z(n20597) );
  AND U20470 ( .A(n20608), .B(n20609), .Z(n20607) );
  XOR U20471 ( .A(n20606), .B(n20215), .Z(n20609) );
  XNOR U20472 ( .A(p_input[1314]), .B(n20610), .Z(n20215) );
  AND U20473 ( .A(n687), .B(n20611), .Z(n20610) );
  XOR U20474 ( .A(p_input[1330]), .B(p_input[1314]), .Z(n20611) );
  XNOR U20475 ( .A(n20212), .B(n20606), .Z(n20608) );
  XOR U20476 ( .A(n20612), .B(n20613), .Z(n20212) );
  AND U20477 ( .A(n684), .B(n20614), .Z(n20613) );
  XOR U20478 ( .A(p_input[1298]), .B(p_input[1282]), .Z(n20614) );
  XOR U20479 ( .A(n20615), .B(n20616), .Z(n20606) );
  AND U20480 ( .A(n20617), .B(n20618), .Z(n20616) );
  XNOR U20481 ( .A(n20619), .B(n20228), .Z(n20618) );
  XNOR U20482 ( .A(p_input[1313]), .B(n20620), .Z(n20228) );
  AND U20483 ( .A(n687), .B(n20621), .Z(n20620) );
  XNOR U20484 ( .A(p_input[1329]), .B(n20622), .Z(n20621) );
  IV U20485 ( .A(p_input[1313]), .Z(n20622) );
  XNOR U20486 ( .A(n20225), .B(n20615), .Z(n20617) );
  XNOR U20487 ( .A(p_input[1281]), .B(n20623), .Z(n20225) );
  AND U20488 ( .A(n684), .B(n20624), .Z(n20623) );
  XOR U20489 ( .A(p_input[1297]), .B(p_input[1281]), .Z(n20624) );
  IV U20490 ( .A(n20619), .Z(n20615) );
  AND U20491 ( .A(n20490), .B(n20493), .Z(n20619) );
  XOR U20492 ( .A(p_input[1312]), .B(n20625), .Z(n20493) );
  AND U20493 ( .A(n687), .B(n20626), .Z(n20625) );
  XOR U20494 ( .A(p_input[1328]), .B(p_input[1312]), .Z(n20626) );
  XOR U20495 ( .A(n20627), .B(n20628), .Z(n687) );
  AND U20496 ( .A(n20629), .B(n20630), .Z(n20628) );
  XNOR U20497 ( .A(p_input[1343]), .B(n20627), .Z(n20630) );
  XOR U20498 ( .A(n20627), .B(p_input[1327]), .Z(n20629) );
  XOR U20499 ( .A(n20631), .B(n20632), .Z(n20627) );
  AND U20500 ( .A(n20633), .B(n20634), .Z(n20632) );
  XNOR U20501 ( .A(p_input[1342]), .B(n20631), .Z(n20634) );
  XOR U20502 ( .A(n20631), .B(p_input[1326]), .Z(n20633) );
  XOR U20503 ( .A(n20635), .B(n20636), .Z(n20631) );
  AND U20504 ( .A(n20637), .B(n20638), .Z(n20636) );
  XNOR U20505 ( .A(p_input[1341]), .B(n20635), .Z(n20638) );
  XOR U20506 ( .A(n20635), .B(p_input[1325]), .Z(n20637) );
  XOR U20507 ( .A(n20639), .B(n20640), .Z(n20635) );
  AND U20508 ( .A(n20641), .B(n20642), .Z(n20640) );
  XNOR U20509 ( .A(p_input[1340]), .B(n20639), .Z(n20642) );
  XOR U20510 ( .A(n20639), .B(p_input[1324]), .Z(n20641) );
  XOR U20511 ( .A(n20643), .B(n20644), .Z(n20639) );
  AND U20512 ( .A(n20645), .B(n20646), .Z(n20644) );
  XNOR U20513 ( .A(p_input[1339]), .B(n20643), .Z(n20646) );
  XOR U20514 ( .A(n20643), .B(p_input[1323]), .Z(n20645) );
  XOR U20515 ( .A(n20647), .B(n20648), .Z(n20643) );
  AND U20516 ( .A(n20649), .B(n20650), .Z(n20648) );
  XNOR U20517 ( .A(p_input[1338]), .B(n20647), .Z(n20650) );
  XOR U20518 ( .A(n20647), .B(p_input[1322]), .Z(n20649) );
  XOR U20519 ( .A(n20651), .B(n20652), .Z(n20647) );
  AND U20520 ( .A(n20653), .B(n20654), .Z(n20652) );
  XNOR U20521 ( .A(p_input[1337]), .B(n20651), .Z(n20654) );
  XOR U20522 ( .A(n20651), .B(p_input[1321]), .Z(n20653) );
  XOR U20523 ( .A(n20655), .B(n20656), .Z(n20651) );
  AND U20524 ( .A(n20657), .B(n20658), .Z(n20656) );
  XNOR U20525 ( .A(p_input[1336]), .B(n20655), .Z(n20658) );
  XOR U20526 ( .A(n20655), .B(p_input[1320]), .Z(n20657) );
  XOR U20527 ( .A(n20659), .B(n20660), .Z(n20655) );
  AND U20528 ( .A(n20661), .B(n20662), .Z(n20660) );
  XNOR U20529 ( .A(p_input[1335]), .B(n20659), .Z(n20662) );
  XOR U20530 ( .A(n20659), .B(p_input[1319]), .Z(n20661) );
  XOR U20531 ( .A(n20663), .B(n20664), .Z(n20659) );
  AND U20532 ( .A(n20665), .B(n20666), .Z(n20664) );
  XNOR U20533 ( .A(p_input[1334]), .B(n20663), .Z(n20666) );
  XOR U20534 ( .A(n20663), .B(p_input[1318]), .Z(n20665) );
  XOR U20535 ( .A(n20667), .B(n20668), .Z(n20663) );
  AND U20536 ( .A(n20669), .B(n20670), .Z(n20668) );
  XNOR U20537 ( .A(p_input[1333]), .B(n20667), .Z(n20670) );
  XOR U20538 ( .A(n20667), .B(p_input[1317]), .Z(n20669) );
  XOR U20539 ( .A(n20671), .B(n20672), .Z(n20667) );
  AND U20540 ( .A(n20673), .B(n20674), .Z(n20672) );
  XNOR U20541 ( .A(p_input[1332]), .B(n20671), .Z(n20674) );
  XOR U20542 ( .A(n20671), .B(p_input[1316]), .Z(n20673) );
  XOR U20543 ( .A(n20675), .B(n20676), .Z(n20671) );
  AND U20544 ( .A(n20677), .B(n20678), .Z(n20676) );
  XNOR U20545 ( .A(p_input[1331]), .B(n20675), .Z(n20678) );
  XOR U20546 ( .A(n20675), .B(p_input[1315]), .Z(n20677) );
  XOR U20547 ( .A(n20679), .B(n20680), .Z(n20675) );
  AND U20548 ( .A(n20681), .B(n20682), .Z(n20680) );
  XNOR U20549 ( .A(p_input[1330]), .B(n20679), .Z(n20682) );
  XOR U20550 ( .A(n20679), .B(p_input[1314]), .Z(n20681) );
  XNOR U20551 ( .A(n20683), .B(n20684), .Z(n20679) );
  AND U20552 ( .A(n20685), .B(n20686), .Z(n20684) );
  XOR U20553 ( .A(p_input[1329]), .B(n20683), .Z(n20686) );
  XNOR U20554 ( .A(p_input[1313]), .B(n20683), .Z(n20685) );
  AND U20555 ( .A(p_input[1328]), .B(n20687), .Z(n20683) );
  IV U20556 ( .A(p_input[1312]), .Z(n20687) );
  XNOR U20557 ( .A(p_input[1280]), .B(n20688), .Z(n20490) );
  AND U20558 ( .A(n684), .B(n20689), .Z(n20688) );
  XOR U20559 ( .A(p_input[1296]), .B(p_input[1280]), .Z(n20689) );
  XOR U20560 ( .A(n20690), .B(n20691), .Z(n684) );
  AND U20561 ( .A(n20692), .B(n20693), .Z(n20691) );
  XNOR U20562 ( .A(p_input[1311]), .B(n20690), .Z(n20693) );
  XOR U20563 ( .A(n20690), .B(p_input[1295]), .Z(n20692) );
  XOR U20564 ( .A(n20694), .B(n20695), .Z(n20690) );
  AND U20565 ( .A(n20696), .B(n20697), .Z(n20695) );
  XNOR U20566 ( .A(p_input[1310]), .B(n20694), .Z(n20697) );
  XNOR U20567 ( .A(n20694), .B(n20504), .Z(n20696) );
  IV U20568 ( .A(p_input[1294]), .Z(n20504) );
  XOR U20569 ( .A(n20698), .B(n20699), .Z(n20694) );
  AND U20570 ( .A(n20700), .B(n20701), .Z(n20699) );
  XNOR U20571 ( .A(p_input[1309]), .B(n20698), .Z(n20701) );
  XNOR U20572 ( .A(n20698), .B(n20513), .Z(n20700) );
  IV U20573 ( .A(p_input[1293]), .Z(n20513) );
  XOR U20574 ( .A(n20702), .B(n20703), .Z(n20698) );
  AND U20575 ( .A(n20704), .B(n20705), .Z(n20703) );
  XNOR U20576 ( .A(p_input[1308]), .B(n20702), .Z(n20705) );
  XNOR U20577 ( .A(n20702), .B(n20522), .Z(n20704) );
  IV U20578 ( .A(p_input[1292]), .Z(n20522) );
  XOR U20579 ( .A(n20706), .B(n20707), .Z(n20702) );
  AND U20580 ( .A(n20708), .B(n20709), .Z(n20707) );
  XNOR U20581 ( .A(p_input[1307]), .B(n20706), .Z(n20709) );
  XNOR U20582 ( .A(n20706), .B(n20531), .Z(n20708) );
  IV U20583 ( .A(p_input[1291]), .Z(n20531) );
  XOR U20584 ( .A(n20710), .B(n20711), .Z(n20706) );
  AND U20585 ( .A(n20712), .B(n20713), .Z(n20711) );
  XNOR U20586 ( .A(p_input[1306]), .B(n20710), .Z(n20713) );
  XNOR U20587 ( .A(n20710), .B(n20540), .Z(n20712) );
  IV U20588 ( .A(p_input[1290]), .Z(n20540) );
  XOR U20589 ( .A(n20714), .B(n20715), .Z(n20710) );
  AND U20590 ( .A(n20716), .B(n20717), .Z(n20715) );
  XNOR U20591 ( .A(p_input[1305]), .B(n20714), .Z(n20717) );
  XNOR U20592 ( .A(n20714), .B(n20549), .Z(n20716) );
  IV U20593 ( .A(p_input[1289]), .Z(n20549) );
  XOR U20594 ( .A(n20718), .B(n20719), .Z(n20714) );
  AND U20595 ( .A(n20720), .B(n20721), .Z(n20719) );
  XNOR U20596 ( .A(p_input[1304]), .B(n20718), .Z(n20721) );
  XNOR U20597 ( .A(n20718), .B(n20558), .Z(n20720) );
  IV U20598 ( .A(p_input[1288]), .Z(n20558) );
  XOR U20599 ( .A(n20722), .B(n20723), .Z(n20718) );
  AND U20600 ( .A(n20724), .B(n20725), .Z(n20723) );
  XNOR U20601 ( .A(p_input[1303]), .B(n20722), .Z(n20725) );
  XNOR U20602 ( .A(n20722), .B(n20567), .Z(n20724) );
  IV U20603 ( .A(p_input[1287]), .Z(n20567) );
  XOR U20604 ( .A(n20726), .B(n20727), .Z(n20722) );
  AND U20605 ( .A(n20728), .B(n20729), .Z(n20727) );
  XNOR U20606 ( .A(p_input[1302]), .B(n20726), .Z(n20729) );
  XNOR U20607 ( .A(n20726), .B(n20576), .Z(n20728) );
  IV U20608 ( .A(p_input[1286]), .Z(n20576) );
  XOR U20609 ( .A(n20730), .B(n20731), .Z(n20726) );
  AND U20610 ( .A(n20732), .B(n20733), .Z(n20731) );
  XNOR U20611 ( .A(p_input[1301]), .B(n20730), .Z(n20733) );
  XNOR U20612 ( .A(n20730), .B(n20585), .Z(n20732) );
  IV U20613 ( .A(p_input[1285]), .Z(n20585) );
  XOR U20614 ( .A(n20734), .B(n20735), .Z(n20730) );
  AND U20615 ( .A(n20736), .B(n20737), .Z(n20735) );
  XNOR U20616 ( .A(p_input[1300]), .B(n20734), .Z(n20737) );
  XNOR U20617 ( .A(n20734), .B(n20594), .Z(n20736) );
  IV U20618 ( .A(p_input[1284]), .Z(n20594) );
  XOR U20619 ( .A(n20738), .B(n20739), .Z(n20734) );
  AND U20620 ( .A(n20740), .B(n20741), .Z(n20739) );
  XNOR U20621 ( .A(p_input[1299]), .B(n20738), .Z(n20741) );
  XNOR U20622 ( .A(n20738), .B(n20603), .Z(n20740) );
  IV U20623 ( .A(p_input[1283]), .Z(n20603) );
  XOR U20624 ( .A(n20742), .B(n20743), .Z(n20738) );
  AND U20625 ( .A(n20744), .B(n20745), .Z(n20743) );
  XNOR U20626 ( .A(p_input[1298]), .B(n20742), .Z(n20745) );
  XNOR U20627 ( .A(n20742), .B(n20612), .Z(n20744) );
  IV U20628 ( .A(p_input[1282]), .Z(n20612) );
  XNOR U20629 ( .A(n20746), .B(n20747), .Z(n20742) );
  AND U20630 ( .A(n20748), .B(n20749), .Z(n20747) );
  XOR U20631 ( .A(p_input[1297]), .B(n20746), .Z(n20749) );
  XNOR U20632 ( .A(p_input[1281]), .B(n20746), .Z(n20748) );
  AND U20633 ( .A(p_input[1296]), .B(n20750), .Z(n20746) );
  IV U20634 ( .A(p_input[1280]), .Z(n20750) );
  XOR U20635 ( .A(n20751), .B(n20752), .Z(n18978) );
  AND U20636 ( .A(n948), .B(n20753), .Z(n20752) );
  XNOR U20637 ( .A(n20754), .B(n20751), .Z(n20753) );
  XOR U20638 ( .A(n20755), .B(n20756), .Z(n948) );
  AND U20639 ( .A(n20757), .B(n20758), .Z(n20756) );
  XNOR U20640 ( .A(n18993), .B(n20755), .Z(n20758) );
  AND U20641 ( .A(n20759), .B(n20760), .Z(n18993) );
  XNOR U20642 ( .A(n20755), .B(n18990), .Z(n20757) );
  IV U20643 ( .A(n20761), .Z(n18990) );
  AND U20644 ( .A(n20762), .B(n20763), .Z(n20761) );
  XOR U20645 ( .A(n20764), .B(n20765), .Z(n20755) );
  AND U20646 ( .A(n20766), .B(n20767), .Z(n20765) );
  XOR U20647 ( .A(n20764), .B(n19005), .Z(n20767) );
  XOR U20648 ( .A(n20768), .B(n20769), .Z(n19005) );
  AND U20649 ( .A(n811), .B(n20770), .Z(n20769) );
  XOR U20650 ( .A(n20771), .B(n20768), .Z(n20770) );
  XNOR U20651 ( .A(n19002), .B(n20764), .Z(n20766) );
  XOR U20652 ( .A(n20772), .B(n20773), .Z(n19002) );
  AND U20653 ( .A(n808), .B(n20774), .Z(n20773) );
  XOR U20654 ( .A(n20775), .B(n20772), .Z(n20774) );
  XOR U20655 ( .A(n20776), .B(n20777), .Z(n20764) );
  AND U20656 ( .A(n20778), .B(n20779), .Z(n20777) );
  XOR U20657 ( .A(n20776), .B(n19017), .Z(n20779) );
  XOR U20658 ( .A(n20780), .B(n20781), .Z(n19017) );
  AND U20659 ( .A(n811), .B(n20782), .Z(n20781) );
  XOR U20660 ( .A(n20783), .B(n20780), .Z(n20782) );
  XNOR U20661 ( .A(n19014), .B(n20776), .Z(n20778) );
  XOR U20662 ( .A(n20784), .B(n20785), .Z(n19014) );
  AND U20663 ( .A(n808), .B(n20786), .Z(n20785) );
  XOR U20664 ( .A(n20787), .B(n20784), .Z(n20786) );
  XOR U20665 ( .A(n20788), .B(n20789), .Z(n20776) );
  AND U20666 ( .A(n20790), .B(n20791), .Z(n20789) );
  XOR U20667 ( .A(n20788), .B(n19029), .Z(n20791) );
  XOR U20668 ( .A(n20792), .B(n20793), .Z(n19029) );
  AND U20669 ( .A(n811), .B(n20794), .Z(n20793) );
  XOR U20670 ( .A(n20795), .B(n20792), .Z(n20794) );
  XNOR U20671 ( .A(n19026), .B(n20788), .Z(n20790) );
  XOR U20672 ( .A(n20796), .B(n20797), .Z(n19026) );
  AND U20673 ( .A(n808), .B(n20798), .Z(n20797) );
  XOR U20674 ( .A(n20799), .B(n20796), .Z(n20798) );
  XOR U20675 ( .A(n20800), .B(n20801), .Z(n20788) );
  AND U20676 ( .A(n20802), .B(n20803), .Z(n20801) );
  XOR U20677 ( .A(n20800), .B(n19041), .Z(n20803) );
  XOR U20678 ( .A(n20804), .B(n20805), .Z(n19041) );
  AND U20679 ( .A(n811), .B(n20806), .Z(n20805) );
  XOR U20680 ( .A(n20807), .B(n20804), .Z(n20806) );
  XNOR U20681 ( .A(n19038), .B(n20800), .Z(n20802) );
  XOR U20682 ( .A(n20808), .B(n20809), .Z(n19038) );
  AND U20683 ( .A(n808), .B(n20810), .Z(n20809) );
  XOR U20684 ( .A(n20811), .B(n20808), .Z(n20810) );
  XOR U20685 ( .A(n20812), .B(n20813), .Z(n20800) );
  AND U20686 ( .A(n20814), .B(n20815), .Z(n20813) );
  XOR U20687 ( .A(n20812), .B(n19053), .Z(n20815) );
  XOR U20688 ( .A(n20816), .B(n20817), .Z(n19053) );
  AND U20689 ( .A(n811), .B(n20818), .Z(n20817) );
  XOR U20690 ( .A(n20819), .B(n20816), .Z(n20818) );
  XNOR U20691 ( .A(n19050), .B(n20812), .Z(n20814) );
  XOR U20692 ( .A(n20820), .B(n20821), .Z(n19050) );
  AND U20693 ( .A(n808), .B(n20822), .Z(n20821) );
  XOR U20694 ( .A(n20823), .B(n20820), .Z(n20822) );
  XOR U20695 ( .A(n20824), .B(n20825), .Z(n20812) );
  AND U20696 ( .A(n20826), .B(n20827), .Z(n20825) );
  XOR U20697 ( .A(n20824), .B(n19065), .Z(n20827) );
  XOR U20698 ( .A(n20828), .B(n20829), .Z(n19065) );
  AND U20699 ( .A(n811), .B(n20830), .Z(n20829) );
  XOR U20700 ( .A(n20831), .B(n20828), .Z(n20830) );
  XNOR U20701 ( .A(n19062), .B(n20824), .Z(n20826) );
  XOR U20702 ( .A(n20832), .B(n20833), .Z(n19062) );
  AND U20703 ( .A(n808), .B(n20834), .Z(n20833) );
  XOR U20704 ( .A(n20835), .B(n20832), .Z(n20834) );
  XOR U20705 ( .A(n20836), .B(n20837), .Z(n20824) );
  AND U20706 ( .A(n20838), .B(n20839), .Z(n20837) );
  XOR U20707 ( .A(n20836), .B(n19077), .Z(n20839) );
  XOR U20708 ( .A(n20840), .B(n20841), .Z(n19077) );
  AND U20709 ( .A(n811), .B(n20842), .Z(n20841) );
  XOR U20710 ( .A(n20843), .B(n20840), .Z(n20842) );
  XNOR U20711 ( .A(n19074), .B(n20836), .Z(n20838) );
  XOR U20712 ( .A(n20844), .B(n20845), .Z(n19074) );
  AND U20713 ( .A(n808), .B(n20846), .Z(n20845) );
  XOR U20714 ( .A(n20847), .B(n20844), .Z(n20846) );
  XOR U20715 ( .A(n20848), .B(n20849), .Z(n20836) );
  AND U20716 ( .A(n20850), .B(n20851), .Z(n20849) );
  XOR U20717 ( .A(n20848), .B(n19089), .Z(n20851) );
  XOR U20718 ( .A(n20852), .B(n20853), .Z(n19089) );
  AND U20719 ( .A(n811), .B(n20854), .Z(n20853) );
  XOR U20720 ( .A(n20855), .B(n20852), .Z(n20854) );
  XNOR U20721 ( .A(n19086), .B(n20848), .Z(n20850) );
  XOR U20722 ( .A(n20856), .B(n20857), .Z(n19086) );
  AND U20723 ( .A(n808), .B(n20858), .Z(n20857) );
  XOR U20724 ( .A(n20859), .B(n20856), .Z(n20858) );
  XOR U20725 ( .A(n20860), .B(n20861), .Z(n20848) );
  AND U20726 ( .A(n20862), .B(n20863), .Z(n20861) );
  XOR U20727 ( .A(n20860), .B(n19101), .Z(n20863) );
  XOR U20728 ( .A(n20864), .B(n20865), .Z(n19101) );
  AND U20729 ( .A(n811), .B(n20866), .Z(n20865) );
  XOR U20730 ( .A(n20867), .B(n20864), .Z(n20866) );
  XNOR U20731 ( .A(n19098), .B(n20860), .Z(n20862) );
  XOR U20732 ( .A(n20868), .B(n20869), .Z(n19098) );
  AND U20733 ( .A(n808), .B(n20870), .Z(n20869) );
  XOR U20734 ( .A(n20871), .B(n20868), .Z(n20870) );
  XOR U20735 ( .A(n20872), .B(n20873), .Z(n20860) );
  AND U20736 ( .A(n20874), .B(n20875), .Z(n20873) );
  XOR U20737 ( .A(n20872), .B(n19113), .Z(n20875) );
  XOR U20738 ( .A(n20876), .B(n20877), .Z(n19113) );
  AND U20739 ( .A(n811), .B(n20878), .Z(n20877) );
  XOR U20740 ( .A(n20879), .B(n20876), .Z(n20878) );
  XNOR U20741 ( .A(n19110), .B(n20872), .Z(n20874) );
  XOR U20742 ( .A(n20880), .B(n20881), .Z(n19110) );
  AND U20743 ( .A(n808), .B(n20882), .Z(n20881) );
  XOR U20744 ( .A(n20883), .B(n20880), .Z(n20882) );
  XOR U20745 ( .A(n20884), .B(n20885), .Z(n20872) );
  AND U20746 ( .A(n20886), .B(n20887), .Z(n20885) );
  XOR U20747 ( .A(n20884), .B(n19125), .Z(n20887) );
  XOR U20748 ( .A(n20888), .B(n20889), .Z(n19125) );
  AND U20749 ( .A(n811), .B(n20890), .Z(n20889) );
  XOR U20750 ( .A(n20891), .B(n20888), .Z(n20890) );
  XNOR U20751 ( .A(n19122), .B(n20884), .Z(n20886) );
  XOR U20752 ( .A(n20892), .B(n20893), .Z(n19122) );
  AND U20753 ( .A(n808), .B(n20894), .Z(n20893) );
  XOR U20754 ( .A(n20895), .B(n20892), .Z(n20894) );
  XOR U20755 ( .A(n20896), .B(n20897), .Z(n20884) );
  AND U20756 ( .A(n20898), .B(n20899), .Z(n20897) );
  XOR U20757 ( .A(n20896), .B(n19137), .Z(n20899) );
  XOR U20758 ( .A(n20900), .B(n20901), .Z(n19137) );
  AND U20759 ( .A(n811), .B(n20902), .Z(n20901) );
  XOR U20760 ( .A(n20903), .B(n20900), .Z(n20902) );
  XNOR U20761 ( .A(n19134), .B(n20896), .Z(n20898) );
  XOR U20762 ( .A(n20904), .B(n20905), .Z(n19134) );
  AND U20763 ( .A(n808), .B(n20906), .Z(n20905) );
  XOR U20764 ( .A(n20907), .B(n20904), .Z(n20906) );
  XOR U20765 ( .A(n20908), .B(n20909), .Z(n20896) );
  AND U20766 ( .A(n20910), .B(n20911), .Z(n20909) );
  XOR U20767 ( .A(n20908), .B(n19149), .Z(n20911) );
  XOR U20768 ( .A(n20912), .B(n20913), .Z(n19149) );
  AND U20769 ( .A(n811), .B(n20914), .Z(n20913) );
  XOR U20770 ( .A(n20915), .B(n20912), .Z(n20914) );
  XNOR U20771 ( .A(n19146), .B(n20908), .Z(n20910) );
  XOR U20772 ( .A(n20916), .B(n20917), .Z(n19146) );
  AND U20773 ( .A(n808), .B(n20918), .Z(n20917) );
  XOR U20774 ( .A(n20919), .B(n20916), .Z(n20918) );
  XOR U20775 ( .A(n20920), .B(n20921), .Z(n20908) );
  AND U20776 ( .A(n20922), .B(n20923), .Z(n20921) );
  XNOR U20777 ( .A(n20924), .B(n19162), .Z(n20923) );
  XOR U20778 ( .A(n20925), .B(n20926), .Z(n19162) );
  AND U20779 ( .A(n811), .B(n20927), .Z(n20926) );
  XOR U20780 ( .A(n20925), .B(n20928), .Z(n20927) );
  XNOR U20781 ( .A(n19159), .B(n20920), .Z(n20922) );
  XOR U20782 ( .A(n20929), .B(n20930), .Z(n19159) );
  AND U20783 ( .A(n808), .B(n20931), .Z(n20930) );
  XOR U20784 ( .A(n20929), .B(n20932), .Z(n20931) );
  IV U20785 ( .A(n20924), .Z(n20920) );
  AND U20786 ( .A(n20751), .B(n20754), .Z(n20924) );
  XNOR U20787 ( .A(n20933), .B(n20934), .Z(n20754) );
  AND U20788 ( .A(n811), .B(n20935), .Z(n20934) );
  XNOR U20789 ( .A(n20936), .B(n20933), .Z(n20935) );
  XOR U20790 ( .A(n20937), .B(n20938), .Z(n811) );
  AND U20791 ( .A(n20939), .B(n20940), .Z(n20938) );
  XNOR U20792 ( .A(n20759), .B(n20937), .Z(n20940) );
  AND U20793 ( .A(n20941), .B(n20942), .Z(n20759) );
  XOR U20794 ( .A(n20937), .B(n20760), .Z(n20939) );
  AND U20795 ( .A(n20943), .B(n20944), .Z(n20760) );
  XOR U20796 ( .A(n20945), .B(n20946), .Z(n20937) );
  AND U20797 ( .A(n20947), .B(n20948), .Z(n20946) );
  XOR U20798 ( .A(n20945), .B(n20771), .Z(n20948) );
  XOR U20799 ( .A(n20949), .B(n20950), .Z(n20771) );
  AND U20800 ( .A(n523), .B(n20951), .Z(n20950) );
  XOR U20801 ( .A(n20952), .B(n20949), .Z(n20951) );
  XNOR U20802 ( .A(n20768), .B(n20945), .Z(n20947) );
  XOR U20803 ( .A(n20953), .B(n20954), .Z(n20768) );
  AND U20804 ( .A(n521), .B(n20955), .Z(n20954) );
  XOR U20805 ( .A(n20956), .B(n20953), .Z(n20955) );
  XOR U20806 ( .A(n20957), .B(n20958), .Z(n20945) );
  AND U20807 ( .A(n20959), .B(n20960), .Z(n20958) );
  XOR U20808 ( .A(n20957), .B(n20783), .Z(n20960) );
  XOR U20809 ( .A(n20961), .B(n20962), .Z(n20783) );
  AND U20810 ( .A(n523), .B(n20963), .Z(n20962) );
  XOR U20811 ( .A(n20964), .B(n20961), .Z(n20963) );
  XNOR U20812 ( .A(n20780), .B(n20957), .Z(n20959) );
  XOR U20813 ( .A(n20965), .B(n20966), .Z(n20780) );
  AND U20814 ( .A(n521), .B(n20967), .Z(n20966) );
  XOR U20815 ( .A(n20968), .B(n20965), .Z(n20967) );
  XOR U20816 ( .A(n20969), .B(n20970), .Z(n20957) );
  AND U20817 ( .A(n20971), .B(n20972), .Z(n20970) );
  XOR U20818 ( .A(n20969), .B(n20795), .Z(n20972) );
  XOR U20819 ( .A(n20973), .B(n20974), .Z(n20795) );
  AND U20820 ( .A(n523), .B(n20975), .Z(n20974) );
  XOR U20821 ( .A(n20976), .B(n20973), .Z(n20975) );
  XNOR U20822 ( .A(n20792), .B(n20969), .Z(n20971) );
  XOR U20823 ( .A(n20977), .B(n20978), .Z(n20792) );
  AND U20824 ( .A(n521), .B(n20979), .Z(n20978) );
  XOR U20825 ( .A(n20980), .B(n20977), .Z(n20979) );
  XOR U20826 ( .A(n20981), .B(n20982), .Z(n20969) );
  AND U20827 ( .A(n20983), .B(n20984), .Z(n20982) );
  XOR U20828 ( .A(n20981), .B(n20807), .Z(n20984) );
  XOR U20829 ( .A(n20985), .B(n20986), .Z(n20807) );
  AND U20830 ( .A(n523), .B(n20987), .Z(n20986) );
  XOR U20831 ( .A(n20988), .B(n20985), .Z(n20987) );
  XNOR U20832 ( .A(n20804), .B(n20981), .Z(n20983) );
  XOR U20833 ( .A(n20989), .B(n20990), .Z(n20804) );
  AND U20834 ( .A(n521), .B(n20991), .Z(n20990) );
  XOR U20835 ( .A(n20992), .B(n20989), .Z(n20991) );
  XOR U20836 ( .A(n20993), .B(n20994), .Z(n20981) );
  AND U20837 ( .A(n20995), .B(n20996), .Z(n20994) );
  XOR U20838 ( .A(n20993), .B(n20819), .Z(n20996) );
  XOR U20839 ( .A(n20997), .B(n20998), .Z(n20819) );
  AND U20840 ( .A(n523), .B(n20999), .Z(n20998) );
  XOR U20841 ( .A(n21000), .B(n20997), .Z(n20999) );
  XNOR U20842 ( .A(n20816), .B(n20993), .Z(n20995) );
  XOR U20843 ( .A(n21001), .B(n21002), .Z(n20816) );
  AND U20844 ( .A(n521), .B(n21003), .Z(n21002) );
  XOR U20845 ( .A(n21004), .B(n21001), .Z(n21003) );
  XOR U20846 ( .A(n21005), .B(n21006), .Z(n20993) );
  AND U20847 ( .A(n21007), .B(n21008), .Z(n21006) );
  XOR U20848 ( .A(n21005), .B(n20831), .Z(n21008) );
  XOR U20849 ( .A(n21009), .B(n21010), .Z(n20831) );
  AND U20850 ( .A(n523), .B(n21011), .Z(n21010) );
  XOR U20851 ( .A(n21012), .B(n21009), .Z(n21011) );
  XNOR U20852 ( .A(n20828), .B(n21005), .Z(n21007) );
  XOR U20853 ( .A(n21013), .B(n21014), .Z(n20828) );
  AND U20854 ( .A(n521), .B(n21015), .Z(n21014) );
  XOR U20855 ( .A(n21016), .B(n21013), .Z(n21015) );
  XOR U20856 ( .A(n21017), .B(n21018), .Z(n21005) );
  AND U20857 ( .A(n21019), .B(n21020), .Z(n21018) );
  XOR U20858 ( .A(n21017), .B(n20843), .Z(n21020) );
  XOR U20859 ( .A(n21021), .B(n21022), .Z(n20843) );
  AND U20860 ( .A(n523), .B(n21023), .Z(n21022) );
  XOR U20861 ( .A(n21024), .B(n21021), .Z(n21023) );
  XNOR U20862 ( .A(n20840), .B(n21017), .Z(n21019) );
  XOR U20863 ( .A(n21025), .B(n21026), .Z(n20840) );
  AND U20864 ( .A(n521), .B(n21027), .Z(n21026) );
  XOR U20865 ( .A(n21028), .B(n21025), .Z(n21027) );
  XOR U20866 ( .A(n21029), .B(n21030), .Z(n21017) );
  AND U20867 ( .A(n21031), .B(n21032), .Z(n21030) );
  XOR U20868 ( .A(n21029), .B(n20855), .Z(n21032) );
  XOR U20869 ( .A(n21033), .B(n21034), .Z(n20855) );
  AND U20870 ( .A(n523), .B(n21035), .Z(n21034) );
  XOR U20871 ( .A(n21036), .B(n21033), .Z(n21035) );
  XNOR U20872 ( .A(n20852), .B(n21029), .Z(n21031) );
  XOR U20873 ( .A(n21037), .B(n21038), .Z(n20852) );
  AND U20874 ( .A(n521), .B(n21039), .Z(n21038) );
  XOR U20875 ( .A(n21040), .B(n21037), .Z(n21039) );
  XOR U20876 ( .A(n21041), .B(n21042), .Z(n21029) );
  AND U20877 ( .A(n21043), .B(n21044), .Z(n21042) );
  XOR U20878 ( .A(n21041), .B(n20867), .Z(n21044) );
  XOR U20879 ( .A(n21045), .B(n21046), .Z(n20867) );
  AND U20880 ( .A(n523), .B(n21047), .Z(n21046) );
  XOR U20881 ( .A(n21048), .B(n21045), .Z(n21047) );
  XNOR U20882 ( .A(n20864), .B(n21041), .Z(n21043) );
  XOR U20883 ( .A(n21049), .B(n21050), .Z(n20864) );
  AND U20884 ( .A(n521), .B(n21051), .Z(n21050) );
  XOR U20885 ( .A(n21052), .B(n21049), .Z(n21051) );
  XOR U20886 ( .A(n21053), .B(n21054), .Z(n21041) );
  AND U20887 ( .A(n21055), .B(n21056), .Z(n21054) );
  XOR U20888 ( .A(n21053), .B(n20879), .Z(n21056) );
  XOR U20889 ( .A(n21057), .B(n21058), .Z(n20879) );
  AND U20890 ( .A(n523), .B(n21059), .Z(n21058) );
  XOR U20891 ( .A(n21060), .B(n21057), .Z(n21059) );
  XNOR U20892 ( .A(n20876), .B(n21053), .Z(n21055) );
  XOR U20893 ( .A(n21061), .B(n21062), .Z(n20876) );
  AND U20894 ( .A(n521), .B(n21063), .Z(n21062) );
  XOR U20895 ( .A(n21064), .B(n21061), .Z(n21063) );
  XOR U20896 ( .A(n21065), .B(n21066), .Z(n21053) );
  AND U20897 ( .A(n21067), .B(n21068), .Z(n21066) );
  XOR U20898 ( .A(n21065), .B(n20891), .Z(n21068) );
  XOR U20899 ( .A(n21069), .B(n21070), .Z(n20891) );
  AND U20900 ( .A(n523), .B(n21071), .Z(n21070) );
  XOR U20901 ( .A(n21072), .B(n21069), .Z(n21071) );
  XNOR U20902 ( .A(n20888), .B(n21065), .Z(n21067) );
  XOR U20903 ( .A(n21073), .B(n21074), .Z(n20888) );
  AND U20904 ( .A(n521), .B(n21075), .Z(n21074) );
  XOR U20905 ( .A(n21076), .B(n21073), .Z(n21075) );
  XOR U20906 ( .A(n21077), .B(n21078), .Z(n21065) );
  AND U20907 ( .A(n21079), .B(n21080), .Z(n21078) );
  XOR U20908 ( .A(n21077), .B(n20903), .Z(n21080) );
  XOR U20909 ( .A(n21081), .B(n21082), .Z(n20903) );
  AND U20910 ( .A(n523), .B(n21083), .Z(n21082) );
  XOR U20911 ( .A(n21084), .B(n21081), .Z(n21083) );
  XNOR U20912 ( .A(n20900), .B(n21077), .Z(n21079) );
  XOR U20913 ( .A(n21085), .B(n21086), .Z(n20900) );
  AND U20914 ( .A(n521), .B(n21087), .Z(n21086) );
  XOR U20915 ( .A(n21088), .B(n21085), .Z(n21087) );
  XOR U20916 ( .A(n21089), .B(n21090), .Z(n21077) );
  AND U20917 ( .A(n21091), .B(n21092), .Z(n21090) );
  XOR U20918 ( .A(n21089), .B(n20915), .Z(n21092) );
  XOR U20919 ( .A(n21093), .B(n21094), .Z(n20915) );
  AND U20920 ( .A(n523), .B(n21095), .Z(n21094) );
  XOR U20921 ( .A(n21096), .B(n21093), .Z(n21095) );
  XNOR U20922 ( .A(n20912), .B(n21089), .Z(n21091) );
  XOR U20923 ( .A(n21097), .B(n21098), .Z(n20912) );
  AND U20924 ( .A(n521), .B(n21099), .Z(n21098) );
  XOR U20925 ( .A(n21100), .B(n21097), .Z(n21099) );
  XOR U20926 ( .A(n21101), .B(n21102), .Z(n21089) );
  AND U20927 ( .A(n21103), .B(n21104), .Z(n21102) );
  XNOR U20928 ( .A(n21105), .B(n20928), .Z(n21104) );
  XOR U20929 ( .A(n21106), .B(n21107), .Z(n20928) );
  AND U20930 ( .A(n523), .B(n21108), .Z(n21107) );
  XOR U20931 ( .A(n21106), .B(n21109), .Z(n21108) );
  XNOR U20932 ( .A(n20925), .B(n21101), .Z(n21103) );
  XOR U20933 ( .A(n21110), .B(n21111), .Z(n20925) );
  AND U20934 ( .A(n521), .B(n21112), .Z(n21111) );
  XOR U20935 ( .A(n21110), .B(n21113), .Z(n21112) );
  IV U20936 ( .A(n21105), .Z(n21101) );
  AND U20937 ( .A(n20933), .B(n20936), .Z(n21105) );
  XNOR U20938 ( .A(n21114), .B(n21115), .Z(n20936) );
  AND U20939 ( .A(n523), .B(n21116), .Z(n21115) );
  XNOR U20940 ( .A(n21117), .B(n21114), .Z(n21116) );
  XOR U20941 ( .A(n21118), .B(n21119), .Z(n523) );
  AND U20942 ( .A(n21120), .B(n21121), .Z(n21119) );
  XNOR U20943 ( .A(n20941), .B(n21118), .Z(n21121) );
  AND U20944 ( .A(p_input[1279]), .B(p_input[1263]), .Z(n20941) );
  XOR U20945 ( .A(n21118), .B(n20942), .Z(n21120) );
  AND U20946 ( .A(p_input[1247]), .B(p_input[1231]), .Z(n20942) );
  XOR U20947 ( .A(n21122), .B(n21123), .Z(n21118) );
  AND U20948 ( .A(n21124), .B(n21125), .Z(n21123) );
  XOR U20949 ( .A(n21122), .B(n20952), .Z(n21125) );
  XNOR U20950 ( .A(p_input[1262]), .B(n21126), .Z(n20952) );
  AND U20951 ( .A(n699), .B(n21127), .Z(n21126) );
  XOR U20952 ( .A(p_input[1278]), .B(p_input[1262]), .Z(n21127) );
  XNOR U20953 ( .A(n20949), .B(n21122), .Z(n21124) );
  XOR U20954 ( .A(n21128), .B(n21129), .Z(n20949) );
  AND U20955 ( .A(n697), .B(n21130), .Z(n21129) );
  XOR U20956 ( .A(p_input[1246]), .B(p_input[1230]), .Z(n21130) );
  XOR U20957 ( .A(n21131), .B(n21132), .Z(n21122) );
  AND U20958 ( .A(n21133), .B(n21134), .Z(n21132) );
  XOR U20959 ( .A(n21131), .B(n20964), .Z(n21134) );
  XNOR U20960 ( .A(p_input[1261]), .B(n21135), .Z(n20964) );
  AND U20961 ( .A(n699), .B(n21136), .Z(n21135) );
  XOR U20962 ( .A(p_input[1277]), .B(p_input[1261]), .Z(n21136) );
  XNOR U20963 ( .A(n20961), .B(n21131), .Z(n21133) );
  XOR U20964 ( .A(n21137), .B(n21138), .Z(n20961) );
  AND U20965 ( .A(n697), .B(n21139), .Z(n21138) );
  XOR U20966 ( .A(p_input[1245]), .B(p_input[1229]), .Z(n21139) );
  XOR U20967 ( .A(n21140), .B(n21141), .Z(n21131) );
  AND U20968 ( .A(n21142), .B(n21143), .Z(n21141) );
  XOR U20969 ( .A(n21140), .B(n20976), .Z(n21143) );
  XNOR U20970 ( .A(p_input[1260]), .B(n21144), .Z(n20976) );
  AND U20971 ( .A(n699), .B(n21145), .Z(n21144) );
  XOR U20972 ( .A(p_input[1276]), .B(p_input[1260]), .Z(n21145) );
  XNOR U20973 ( .A(n20973), .B(n21140), .Z(n21142) );
  XOR U20974 ( .A(n21146), .B(n21147), .Z(n20973) );
  AND U20975 ( .A(n697), .B(n21148), .Z(n21147) );
  XOR U20976 ( .A(p_input[1244]), .B(p_input[1228]), .Z(n21148) );
  XOR U20977 ( .A(n21149), .B(n21150), .Z(n21140) );
  AND U20978 ( .A(n21151), .B(n21152), .Z(n21150) );
  XOR U20979 ( .A(n21149), .B(n20988), .Z(n21152) );
  XNOR U20980 ( .A(p_input[1259]), .B(n21153), .Z(n20988) );
  AND U20981 ( .A(n699), .B(n21154), .Z(n21153) );
  XOR U20982 ( .A(p_input[1275]), .B(p_input[1259]), .Z(n21154) );
  XNOR U20983 ( .A(n20985), .B(n21149), .Z(n21151) );
  XOR U20984 ( .A(n21155), .B(n21156), .Z(n20985) );
  AND U20985 ( .A(n697), .B(n21157), .Z(n21156) );
  XOR U20986 ( .A(p_input[1243]), .B(p_input[1227]), .Z(n21157) );
  XOR U20987 ( .A(n21158), .B(n21159), .Z(n21149) );
  AND U20988 ( .A(n21160), .B(n21161), .Z(n21159) );
  XOR U20989 ( .A(n21158), .B(n21000), .Z(n21161) );
  XNOR U20990 ( .A(p_input[1258]), .B(n21162), .Z(n21000) );
  AND U20991 ( .A(n699), .B(n21163), .Z(n21162) );
  XOR U20992 ( .A(p_input[1274]), .B(p_input[1258]), .Z(n21163) );
  XNOR U20993 ( .A(n20997), .B(n21158), .Z(n21160) );
  XOR U20994 ( .A(n21164), .B(n21165), .Z(n20997) );
  AND U20995 ( .A(n697), .B(n21166), .Z(n21165) );
  XOR U20996 ( .A(p_input[1242]), .B(p_input[1226]), .Z(n21166) );
  XOR U20997 ( .A(n21167), .B(n21168), .Z(n21158) );
  AND U20998 ( .A(n21169), .B(n21170), .Z(n21168) );
  XOR U20999 ( .A(n21167), .B(n21012), .Z(n21170) );
  XNOR U21000 ( .A(p_input[1257]), .B(n21171), .Z(n21012) );
  AND U21001 ( .A(n699), .B(n21172), .Z(n21171) );
  XOR U21002 ( .A(p_input[1273]), .B(p_input[1257]), .Z(n21172) );
  XNOR U21003 ( .A(n21009), .B(n21167), .Z(n21169) );
  XOR U21004 ( .A(n21173), .B(n21174), .Z(n21009) );
  AND U21005 ( .A(n697), .B(n21175), .Z(n21174) );
  XOR U21006 ( .A(p_input[1241]), .B(p_input[1225]), .Z(n21175) );
  XOR U21007 ( .A(n21176), .B(n21177), .Z(n21167) );
  AND U21008 ( .A(n21178), .B(n21179), .Z(n21177) );
  XOR U21009 ( .A(n21176), .B(n21024), .Z(n21179) );
  XNOR U21010 ( .A(p_input[1256]), .B(n21180), .Z(n21024) );
  AND U21011 ( .A(n699), .B(n21181), .Z(n21180) );
  XOR U21012 ( .A(p_input[1272]), .B(p_input[1256]), .Z(n21181) );
  XNOR U21013 ( .A(n21021), .B(n21176), .Z(n21178) );
  XOR U21014 ( .A(n21182), .B(n21183), .Z(n21021) );
  AND U21015 ( .A(n697), .B(n21184), .Z(n21183) );
  XOR U21016 ( .A(p_input[1240]), .B(p_input[1224]), .Z(n21184) );
  XOR U21017 ( .A(n21185), .B(n21186), .Z(n21176) );
  AND U21018 ( .A(n21187), .B(n21188), .Z(n21186) );
  XOR U21019 ( .A(n21185), .B(n21036), .Z(n21188) );
  XNOR U21020 ( .A(p_input[1255]), .B(n21189), .Z(n21036) );
  AND U21021 ( .A(n699), .B(n21190), .Z(n21189) );
  XOR U21022 ( .A(p_input[1271]), .B(p_input[1255]), .Z(n21190) );
  XNOR U21023 ( .A(n21033), .B(n21185), .Z(n21187) );
  XOR U21024 ( .A(n21191), .B(n21192), .Z(n21033) );
  AND U21025 ( .A(n697), .B(n21193), .Z(n21192) );
  XOR U21026 ( .A(p_input[1239]), .B(p_input[1223]), .Z(n21193) );
  XOR U21027 ( .A(n21194), .B(n21195), .Z(n21185) );
  AND U21028 ( .A(n21196), .B(n21197), .Z(n21195) );
  XOR U21029 ( .A(n21194), .B(n21048), .Z(n21197) );
  XNOR U21030 ( .A(p_input[1254]), .B(n21198), .Z(n21048) );
  AND U21031 ( .A(n699), .B(n21199), .Z(n21198) );
  XOR U21032 ( .A(p_input[1270]), .B(p_input[1254]), .Z(n21199) );
  XNOR U21033 ( .A(n21045), .B(n21194), .Z(n21196) );
  XOR U21034 ( .A(n21200), .B(n21201), .Z(n21045) );
  AND U21035 ( .A(n697), .B(n21202), .Z(n21201) );
  XOR U21036 ( .A(p_input[1238]), .B(p_input[1222]), .Z(n21202) );
  XOR U21037 ( .A(n21203), .B(n21204), .Z(n21194) );
  AND U21038 ( .A(n21205), .B(n21206), .Z(n21204) );
  XOR U21039 ( .A(n21203), .B(n21060), .Z(n21206) );
  XNOR U21040 ( .A(p_input[1253]), .B(n21207), .Z(n21060) );
  AND U21041 ( .A(n699), .B(n21208), .Z(n21207) );
  XOR U21042 ( .A(p_input[1269]), .B(p_input[1253]), .Z(n21208) );
  XNOR U21043 ( .A(n21057), .B(n21203), .Z(n21205) );
  XOR U21044 ( .A(n21209), .B(n21210), .Z(n21057) );
  AND U21045 ( .A(n697), .B(n21211), .Z(n21210) );
  XOR U21046 ( .A(p_input[1237]), .B(p_input[1221]), .Z(n21211) );
  XOR U21047 ( .A(n21212), .B(n21213), .Z(n21203) );
  AND U21048 ( .A(n21214), .B(n21215), .Z(n21213) );
  XOR U21049 ( .A(n21212), .B(n21072), .Z(n21215) );
  XNOR U21050 ( .A(p_input[1252]), .B(n21216), .Z(n21072) );
  AND U21051 ( .A(n699), .B(n21217), .Z(n21216) );
  XOR U21052 ( .A(p_input[1268]), .B(p_input[1252]), .Z(n21217) );
  XNOR U21053 ( .A(n21069), .B(n21212), .Z(n21214) );
  XOR U21054 ( .A(n21218), .B(n21219), .Z(n21069) );
  AND U21055 ( .A(n697), .B(n21220), .Z(n21219) );
  XOR U21056 ( .A(p_input[1236]), .B(p_input[1220]), .Z(n21220) );
  XOR U21057 ( .A(n21221), .B(n21222), .Z(n21212) );
  AND U21058 ( .A(n21223), .B(n21224), .Z(n21222) );
  XOR U21059 ( .A(n21221), .B(n21084), .Z(n21224) );
  XNOR U21060 ( .A(p_input[1251]), .B(n21225), .Z(n21084) );
  AND U21061 ( .A(n699), .B(n21226), .Z(n21225) );
  XOR U21062 ( .A(p_input[1267]), .B(p_input[1251]), .Z(n21226) );
  XNOR U21063 ( .A(n21081), .B(n21221), .Z(n21223) );
  XOR U21064 ( .A(n21227), .B(n21228), .Z(n21081) );
  AND U21065 ( .A(n697), .B(n21229), .Z(n21228) );
  XOR U21066 ( .A(p_input[1235]), .B(p_input[1219]), .Z(n21229) );
  XOR U21067 ( .A(n21230), .B(n21231), .Z(n21221) );
  AND U21068 ( .A(n21232), .B(n21233), .Z(n21231) );
  XOR U21069 ( .A(n21230), .B(n21096), .Z(n21233) );
  XNOR U21070 ( .A(p_input[1250]), .B(n21234), .Z(n21096) );
  AND U21071 ( .A(n699), .B(n21235), .Z(n21234) );
  XOR U21072 ( .A(p_input[1266]), .B(p_input[1250]), .Z(n21235) );
  XNOR U21073 ( .A(n21093), .B(n21230), .Z(n21232) );
  XOR U21074 ( .A(n21236), .B(n21237), .Z(n21093) );
  AND U21075 ( .A(n697), .B(n21238), .Z(n21237) );
  XOR U21076 ( .A(p_input[1234]), .B(p_input[1218]), .Z(n21238) );
  XOR U21077 ( .A(n21239), .B(n21240), .Z(n21230) );
  AND U21078 ( .A(n21241), .B(n21242), .Z(n21240) );
  XNOR U21079 ( .A(n21243), .B(n21109), .Z(n21242) );
  XNOR U21080 ( .A(p_input[1249]), .B(n21244), .Z(n21109) );
  AND U21081 ( .A(n699), .B(n21245), .Z(n21244) );
  XNOR U21082 ( .A(p_input[1265]), .B(n21246), .Z(n21245) );
  IV U21083 ( .A(p_input[1249]), .Z(n21246) );
  XNOR U21084 ( .A(n21106), .B(n21239), .Z(n21241) );
  XNOR U21085 ( .A(p_input[1217]), .B(n21247), .Z(n21106) );
  AND U21086 ( .A(n697), .B(n21248), .Z(n21247) );
  XOR U21087 ( .A(p_input[1233]), .B(p_input[1217]), .Z(n21248) );
  IV U21088 ( .A(n21243), .Z(n21239) );
  AND U21089 ( .A(n21114), .B(n21117), .Z(n21243) );
  XOR U21090 ( .A(p_input[1248]), .B(n21249), .Z(n21117) );
  AND U21091 ( .A(n699), .B(n21250), .Z(n21249) );
  XOR U21092 ( .A(p_input[1264]), .B(p_input[1248]), .Z(n21250) );
  XOR U21093 ( .A(n21251), .B(n21252), .Z(n699) );
  AND U21094 ( .A(n21253), .B(n21254), .Z(n21252) );
  XNOR U21095 ( .A(p_input[1279]), .B(n21251), .Z(n21254) );
  XOR U21096 ( .A(n21251), .B(p_input[1263]), .Z(n21253) );
  XOR U21097 ( .A(n21255), .B(n21256), .Z(n21251) );
  AND U21098 ( .A(n21257), .B(n21258), .Z(n21256) );
  XNOR U21099 ( .A(p_input[1278]), .B(n21255), .Z(n21258) );
  XOR U21100 ( .A(n21255), .B(p_input[1262]), .Z(n21257) );
  XOR U21101 ( .A(n21259), .B(n21260), .Z(n21255) );
  AND U21102 ( .A(n21261), .B(n21262), .Z(n21260) );
  XNOR U21103 ( .A(p_input[1277]), .B(n21259), .Z(n21262) );
  XOR U21104 ( .A(n21259), .B(p_input[1261]), .Z(n21261) );
  XOR U21105 ( .A(n21263), .B(n21264), .Z(n21259) );
  AND U21106 ( .A(n21265), .B(n21266), .Z(n21264) );
  XNOR U21107 ( .A(p_input[1276]), .B(n21263), .Z(n21266) );
  XOR U21108 ( .A(n21263), .B(p_input[1260]), .Z(n21265) );
  XOR U21109 ( .A(n21267), .B(n21268), .Z(n21263) );
  AND U21110 ( .A(n21269), .B(n21270), .Z(n21268) );
  XNOR U21111 ( .A(p_input[1275]), .B(n21267), .Z(n21270) );
  XOR U21112 ( .A(n21267), .B(p_input[1259]), .Z(n21269) );
  XOR U21113 ( .A(n21271), .B(n21272), .Z(n21267) );
  AND U21114 ( .A(n21273), .B(n21274), .Z(n21272) );
  XNOR U21115 ( .A(p_input[1274]), .B(n21271), .Z(n21274) );
  XOR U21116 ( .A(n21271), .B(p_input[1258]), .Z(n21273) );
  XOR U21117 ( .A(n21275), .B(n21276), .Z(n21271) );
  AND U21118 ( .A(n21277), .B(n21278), .Z(n21276) );
  XNOR U21119 ( .A(p_input[1273]), .B(n21275), .Z(n21278) );
  XOR U21120 ( .A(n21275), .B(p_input[1257]), .Z(n21277) );
  XOR U21121 ( .A(n21279), .B(n21280), .Z(n21275) );
  AND U21122 ( .A(n21281), .B(n21282), .Z(n21280) );
  XNOR U21123 ( .A(p_input[1272]), .B(n21279), .Z(n21282) );
  XOR U21124 ( .A(n21279), .B(p_input[1256]), .Z(n21281) );
  XOR U21125 ( .A(n21283), .B(n21284), .Z(n21279) );
  AND U21126 ( .A(n21285), .B(n21286), .Z(n21284) );
  XNOR U21127 ( .A(p_input[1271]), .B(n21283), .Z(n21286) );
  XOR U21128 ( .A(n21283), .B(p_input[1255]), .Z(n21285) );
  XOR U21129 ( .A(n21287), .B(n21288), .Z(n21283) );
  AND U21130 ( .A(n21289), .B(n21290), .Z(n21288) );
  XNOR U21131 ( .A(p_input[1270]), .B(n21287), .Z(n21290) );
  XOR U21132 ( .A(n21287), .B(p_input[1254]), .Z(n21289) );
  XOR U21133 ( .A(n21291), .B(n21292), .Z(n21287) );
  AND U21134 ( .A(n21293), .B(n21294), .Z(n21292) );
  XNOR U21135 ( .A(p_input[1269]), .B(n21291), .Z(n21294) );
  XOR U21136 ( .A(n21291), .B(p_input[1253]), .Z(n21293) );
  XOR U21137 ( .A(n21295), .B(n21296), .Z(n21291) );
  AND U21138 ( .A(n21297), .B(n21298), .Z(n21296) );
  XNOR U21139 ( .A(p_input[1268]), .B(n21295), .Z(n21298) );
  XOR U21140 ( .A(n21295), .B(p_input[1252]), .Z(n21297) );
  XOR U21141 ( .A(n21299), .B(n21300), .Z(n21295) );
  AND U21142 ( .A(n21301), .B(n21302), .Z(n21300) );
  XNOR U21143 ( .A(p_input[1267]), .B(n21299), .Z(n21302) );
  XOR U21144 ( .A(n21299), .B(p_input[1251]), .Z(n21301) );
  XOR U21145 ( .A(n21303), .B(n21304), .Z(n21299) );
  AND U21146 ( .A(n21305), .B(n21306), .Z(n21304) );
  XNOR U21147 ( .A(p_input[1266]), .B(n21303), .Z(n21306) );
  XOR U21148 ( .A(n21303), .B(p_input[1250]), .Z(n21305) );
  XNOR U21149 ( .A(n21307), .B(n21308), .Z(n21303) );
  AND U21150 ( .A(n21309), .B(n21310), .Z(n21308) );
  XOR U21151 ( .A(p_input[1265]), .B(n21307), .Z(n21310) );
  XNOR U21152 ( .A(p_input[1249]), .B(n21307), .Z(n21309) );
  AND U21153 ( .A(p_input[1264]), .B(n21311), .Z(n21307) );
  IV U21154 ( .A(p_input[1248]), .Z(n21311) );
  XNOR U21155 ( .A(p_input[1216]), .B(n21312), .Z(n21114) );
  AND U21156 ( .A(n697), .B(n21313), .Z(n21312) );
  XOR U21157 ( .A(p_input[1232]), .B(p_input[1216]), .Z(n21313) );
  XOR U21158 ( .A(n21314), .B(n21315), .Z(n697) );
  AND U21159 ( .A(n21316), .B(n21317), .Z(n21315) );
  XNOR U21160 ( .A(p_input[1247]), .B(n21314), .Z(n21317) );
  XOR U21161 ( .A(n21314), .B(p_input[1231]), .Z(n21316) );
  XOR U21162 ( .A(n21318), .B(n21319), .Z(n21314) );
  AND U21163 ( .A(n21320), .B(n21321), .Z(n21319) );
  XNOR U21164 ( .A(p_input[1246]), .B(n21318), .Z(n21321) );
  XNOR U21165 ( .A(n21318), .B(n21128), .Z(n21320) );
  IV U21166 ( .A(p_input[1230]), .Z(n21128) );
  XOR U21167 ( .A(n21322), .B(n21323), .Z(n21318) );
  AND U21168 ( .A(n21324), .B(n21325), .Z(n21323) );
  XNOR U21169 ( .A(p_input[1245]), .B(n21322), .Z(n21325) );
  XNOR U21170 ( .A(n21322), .B(n21137), .Z(n21324) );
  IV U21171 ( .A(p_input[1229]), .Z(n21137) );
  XOR U21172 ( .A(n21326), .B(n21327), .Z(n21322) );
  AND U21173 ( .A(n21328), .B(n21329), .Z(n21327) );
  XNOR U21174 ( .A(p_input[1244]), .B(n21326), .Z(n21329) );
  XNOR U21175 ( .A(n21326), .B(n21146), .Z(n21328) );
  IV U21176 ( .A(p_input[1228]), .Z(n21146) );
  XOR U21177 ( .A(n21330), .B(n21331), .Z(n21326) );
  AND U21178 ( .A(n21332), .B(n21333), .Z(n21331) );
  XNOR U21179 ( .A(p_input[1243]), .B(n21330), .Z(n21333) );
  XNOR U21180 ( .A(n21330), .B(n21155), .Z(n21332) );
  IV U21181 ( .A(p_input[1227]), .Z(n21155) );
  XOR U21182 ( .A(n21334), .B(n21335), .Z(n21330) );
  AND U21183 ( .A(n21336), .B(n21337), .Z(n21335) );
  XNOR U21184 ( .A(p_input[1242]), .B(n21334), .Z(n21337) );
  XNOR U21185 ( .A(n21334), .B(n21164), .Z(n21336) );
  IV U21186 ( .A(p_input[1226]), .Z(n21164) );
  XOR U21187 ( .A(n21338), .B(n21339), .Z(n21334) );
  AND U21188 ( .A(n21340), .B(n21341), .Z(n21339) );
  XNOR U21189 ( .A(p_input[1241]), .B(n21338), .Z(n21341) );
  XNOR U21190 ( .A(n21338), .B(n21173), .Z(n21340) );
  IV U21191 ( .A(p_input[1225]), .Z(n21173) );
  XOR U21192 ( .A(n21342), .B(n21343), .Z(n21338) );
  AND U21193 ( .A(n21344), .B(n21345), .Z(n21343) );
  XNOR U21194 ( .A(p_input[1240]), .B(n21342), .Z(n21345) );
  XNOR U21195 ( .A(n21342), .B(n21182), .Z(n21344) );
  IV U21196 ( .A(p_input[1224]), .Z(n21182) );
  XOR U21197 ( .A(n21346), .B(n21347), .Z(n21342) );
  AND U21198 ( .A(n21348), .B(n21349), .Z(n21347) );
  XNOR U21199 ( .A(p_input[1239]), .B(n21346), .Z(n21349) );
  XNOR U21200 ( .A(n21346), .B(n21191), .Z(n21348) );
  IV U21201 ( .A(p_input[1223]), .Z(n21191) );
  XOR U21202 ( .A(n21350), .B(n21351), .Z(n21346) );
  AND U21203 ( .A(n21352), .B(n21353), .Z(n21351) );
  XNOR U21204 ( .A(p_input[1238]), .B(n21350), .Z(n21353) );
  XNOR U21205 ( .A(n21350), .B(n21200), .Z(n21352) );
  IV U21206 ( .A(p_input[1222]), .Z(n21200) );
  XOR U21207 ( .A(n21354), .B(n21355), .Z(n21350) );
  AND U21208 ( .A(n21356), .B(n21357), .Z(n21355) );
  XNOR U21209 ( .A(p_input[1237]), .B(n21354), .Z(n21357) );
  XNOR U21210 ( .A(n21354), .B(n21209), .Z(n21356) );
  IV U21211 ( .A(p_input[1221]), .Z(n21209) );
  XOR U21212 ( .A(n21358), .B(n21359), .Z(n21354) );
  AND U21213 ( .A(n21360), .B(n21361), .Z(n21359) );
  XNOR U21214 ( .A(p_input[1236]), .B(n21358), .Z(n21361) );
  XNOR U21215 ( .A(n21358), .B(n21218), .Z(n21360) );
  IV U21216 ( .A(p_input[1220]), .Z(n21218) );
  XOR U21217 ( .A(n21362), .B(n21363), .Z(n21358) );
  AND U21218 ( .A(n21364), .B(n21365), .Z(n21363) );
  XNOR U21219 ( .A(p_input[1235]), .B(n21362), .Z(n21365) );
  XNOR U21220 ( .A(n21362), .B(n21227), .Z(n21364) );
  IV U21221 ( .A(p_input[1219]), .Z(n21227) );
  XOR U21222 ( .A(n21366), .B(n21367), .Z(n21362) );
  AND U21223 ( .A(n21368), .B(n21369), .Z(n21367) );
  XNOR U21224 ( .A(p_input[1234]), .B(n21366), .Z(n21369) );
  XNOR U21225 ( .A(n21366), .B(n21236), .Z(n21368) );
  IV U21226 ( .A(p_input[1218]), .Z(n21236) );
  XNOR U21227 ( .A(n21370), .B(n21371), .Z(n21366) );
  AND U21228 ( .A(n21372), .B(n21373), .Z(n21371) );
  XOR U21229 ( .A(p_input[1233]), .B(n21370), .Z(n21373) );
  XNOR U21230 ( .A(p_input[1217]), .B(n21370), .Z(n21372) );
  AND U21231 ( .A(p_input[1232]), .B(n21374), .Z(n21370) );
  IV U21232 ( .A(p_input[1216]), .Z(n21374) );
  XOR U21233 ( .A(n21375), .B(n21376), .Z(n20933) );
  AND U21234 ( .A(n521), .B(n21377), .Z(n21376) );
  XNOR U21235 ( .A(n21378), .B(n21375), .Z(n21377) );
  XOR U21236 ( .A(n21379), .B(n21380), .Z(n521) );
  AND U21237 ( .A(n21381), .B(n21382), .Z(n21380) );
  XNOR U21238 ( .A(n20943), .B(n21379), .Z(n21382) );
  AND U21239 ( .A(p_input[1215]), .B(p_input[1199]), .Z(n20943) );
  XOR U21240 ( .A(n21379), .B(n20944), .Z(n21381) );
  AND U21241 ( .A(p_input[1183]), .B(p_input[1167]), .Z(n20944) );
  XOR U21242 ( .A(n21383), .B(n21384), .Z(n21379) );
  AND U21243 ( .A(n21385), .B(n21386), .Z(n21384) );
  XOR U21244 ( .A(n21383), .B(n20956), .Z(n21386) );
  XNOR U21245 ( .A(p_input[1198]), .B(n21387), .Z(n20956) );
  AND U21246 ( .A(n703), .B(n21388), .Z(n21387) );
  XOR U21247 ( .A(p_input[1214]), .B(p_input[1198]), .Z(n21388) );
  XNOR U21248 ( .A(n20953), .B(n21383), .Z(n21385) );
  XOR U21249 ( .A(n21389), .B(n21390), .Z(n20953) );
  AND U21250 ( .A(n700), .B(n21391), .Z(n21390) );
  XOR U21251 ( .A(p_input[1182]), .B(p_input[1166]), .Z(n21391) );
  XOR U21252 ( .A(n21392), .B(n21393), .Z(n21383) );
  AND U21253 ( .A(n21394), .B(n21395), .Z(n21393) );
  XOR U21254 ( .A(n21392), .B(n20968), .Z(n21395) );
  XNOR U21255 ( .A(p_input[1197]), .B(n21396), .Z(n20968) );
  AND U21256 ( .A(n703), .B(n21397), .Z(n21396) );
  XOR U21257 ( .A(p_input[1213]), .B(p_input[1197]), .Z(n21397) );
  XNOR U21258 ( .A(n20965), .B(n21392), .Z(n21394) );
  XOR U21259 ( .A(n21398), .B(n21399), .Z(n20965) );
  AND U21260 ( .A(n700), .B(n21400), .Z(n21399) );
  XOR U21261 ( .A(p_input[1181]), .B(p_input[1165]), .Z(n21400) );
  XOR U21262 ( .A(n21401), .B(n21402), .Z(n21392) );
  AND U21263 ( .A(n21403), .B(n21404), .Z(n21402) );
  XOR U21264 ( .A(n21401), .B(n20980), .Z(n21404) );
  XNOR U21265 ( .A(p_input[1196]), .B(n21405), .Z(n20980) );
  AND U21266 ( .A(n703), .B(n21406), .Z(n21405) );
  XOR U21267 ( .A(p_input[1212]), .B(p_input[1196]), .Z(n21406) );
  XNOR U21268 ( .A(n20977), .B(n21401), .Z(n21403) );
  XOR U21269 ( .A(n21407), .B(n21408), .Z(n20977) );
  AND U21270 ( .A(n700), .B(n21409), .Z(n21408) );
  XOR U21271 ( .A(p_input[1180]), .B(p_input[1164]), .Z(n21409) );
  XOR U21272 ( .A(n21410), .B(n21411), .Z(n21401) );
  AND U21273 ( .A(n21412), .B(n21413), .Z(n21411) );
  XOR U21274 ( .A(n21410), .B(n20992), .Z(n21413) );
  XNOR U21275 ( .A(p_input[1195]), .B(n21414), .Z(n20992) );
  AND U21276 ( .A(n703), .B(n21415), .Z(n21414) );
  XOR U21277 ( .A(p_input[1211]), .B(p_input[1195]), .Z(n21415) );
  XNOR U21278 ( .A(n20989), .B(n21410), .Z(n21412) );
  XOR U21279 ( .A(n21416), .B(n21417), .Z(n20989) );
  AND U21280 ( .A(n700), .B(n21418), .Z(n21417) );
  XOR U21281 ( .A(p_input[1179]), .B(p_input[1163]), .Z(n21418) );
  XOR U21282 ( .A(n21419), .B(n21420), .Z(n21410) );
  AND U21283 ( .A(n21421), .B(n21422), .Z(n21420) );
  XOR U21284 ( .A(n21419), .B(n21004), .Z(n21422) );
  XNOR U21285 ( .A(p_input[1194]), .B(n21423), .Z(n21004) );
  AND U21286 ( .A(n703), .B(n21424), .Z(n21423) );
  XOR U21287 ( .A(p_input[1210]), .B(p_input[1194]), .Z(n21424) );
  XNOR U21288 ( .A(n21001), .B(n21419), .Z(n21421) );
  XOR U21289 ( .A(n21425), .B(n21426), .Z(n21001) );
  AND U21290 ( .A(n700), .B(n21427), .Z(n21426) );
  XOR U21291 ( .A(p_input[1178]), .B(p_input[1162]), .Z(n21427) );
  XOR U21292 ( .A(n21428), .B(n21429), .Z(n21419) );
  AND U21293 ( .A(n21430), .B(n21431), .Z(n21429) );
  XOR U21294 ( .A(n21428), .B(n21016), .Z(n21431) );
  XNOR U21295 ( .A(p_input[1193]), .B(n21432), .Z(n21016) );
  AND U21296 ( .A(n703), .B(n21433), .Z(n21432) );
  XOR U21297 ( .A(p_input[1209]), .B(p_input[1193]), .Z(n21433) );
  XNOR U21298 ( .A(n21013), .B(n21428), .Z(n21430) );
  XOR U21299 ( .A(n21434), .B(n21435), .Z(n21013) );
  AND U21300 ( .A(n700), .B(n21436), .Z(n21435) );
  XOR U21301 ( .A(p_input[1177]), .B(p_input[1161]), .Z(n21436) );
  XOR U21302 ( .A(n21437), .B(n21438), .Z(n21428) );
  AND U21303 ( .A(n21439), .B(n21440), .Z(n21438) );
  XOR U21304 ( .A(n21437), .B(n21028), .Z(n21440) );
  XNOR U21305 ( .A(p_input[1192]), .B(n21441), .Z(n21028) );
  AND U21306 ( .A(n703), .B(n21442), .Z(n21441) );
  XOR U21307 ( .A(p_input[1208]), .B(p_input[1192]), .Z(n21442) );
  XNOR U21308 ( .A(n21025), .B(n21437), .Z(n21439) );
  XOR U21309 ( .A(n21443), .B(n21444), .Z(n21025) );
  AND U21310 ( .A(n700), .B(n21445), .Z(n21444) );
  XOR U21311 ( .A(p_input[1176]), .B(p_input[1160]), .Z(n21445) );
  XOR U21312 ( .A(n21446), .B(n21447), .Z(n21437) );
  AND U21313 ( .A(n21448), .B(n21449), .Z(n21447) );
  XOR U21314 ( .A(n21446), .B(n21040), .Z(n21449) );
  XNOR U21315 ( .A(p_input[1191]), .B(n21450), .Z(n21040) );
  AND U21316 ( .A(n703), .B(n21451), .Z(n21450) );
  XOR U21317 ( .A(p_input[1207]), .B(p_input[1191]), .Z(n21451) );
  XNOR U21318 ( .A(n21037), .B(n21446), .Z(n21448) );
  XOR U21319 ( .A(n21452), .B(n21453), .Z(n21037) );
  AND U21320 ( .A(n700), .B(n21454), .Z(n21453) );
  XOR U21321 ( .A(p_input[1175]), .B(p_input[1159]), .Z(n21454) );
  XOR U21322 ( .A(n21455), .B(n21456), .Z(n21446) );
  AND U21323 ( .A(n21457), .B(n21458), .Z(n21456) );
  XOR U21324 ( .A(n21455), .B(n21052), .Z(n21458) );
  XNOR U21325 ( .A(p_input[1190]), .B(n21459), .Z(n21052) );
  AND U21326 ( .A(n703), .B(n21460), .Z(n21459) );
  XOR U21327 ( .A(p_input[1206]), .B(p_input[1190]), .Z(n21460) );
  XNOR U21328 ( .A(n21049), .B(n21455), .Z(n21457) );
  XOR U21329 ( .A(n21461), .B(n21462), .Z(n21049) );
  AND U21330 ( .A(n700), .B(n21463), .Z(n21462) );
  XOR U21331 ( .A(p_input[1174]), .B(p_input[1158]), .Z(n21463) );
  XOR U21332 ( .A(n21464), .B(n21465), .Z(n21455) );
  AND U21333 ( .A(n21466), .B(n21467), .Z(n21465) );
  XOR U21334 ( .A(n21464), .B(n21064), .Z(n21467) );
  XNOR U21335 ( .A(p_input[1189]), .B(n21468), .Z(n21064) );
  AND U21336 ( .A(n703), .B(n21469), .Z(n21468) );
  XOR U21337 ( .A(p_input[1205]), .B(p_input[1189]), .Z(n21469) );
  XNOR U21338 ( .A(n21061), .B(n21464), .Z(n21466) );
  XOR U21339 ( .A(n21470), .B(n21471), .Z(n21061) );
  AND U21340 ( .A(n700), .B(n21472), .Z(n21471) );
  XOR U21341 ( .A(p_input[1173]), .B(p_input[1157]), .Z(n21472) );
  XOR U21342 ( .A(n21473), .B(n21474), .Z(n21464) );
  AND U21343 ( .A(n21475), .B(n21476), .Z(n21474) );
  XOR U21344 ( .A(n21473), .B(n21076), .Z(n21476) );
  XNOR U21345 ( .A(p_input[1188]), .B(n21477), .Z(n21076) );
  AND U21346 ( .A(n703), .B(n21478), .Z(n21477) );
  XOR U21347 ( .A(p_input[1204]), .B(p_input[1188]), .Z(n21478) );
  XNOR U21348 ( .A(n21073), .B(n21473), .Z(n21475) );
  XOR U21349 ( .A(n21479), .B(n21480), .Z(n21073) );
  AND U21350 ( .A(n700), .B(n21481), .Z(n21480) );
  XOR U21351 ( .A(p_input[1172]), .B(p_input[1156]), .Z(n21481) );
  XOR U21352 ( .A(n21482), .B(n21483), .Z(n21473) );
  AND U21353 ( .A(n21484), .B(n21485), .Z(n21483) );
  XOR U21354 ( .A(n21482), .B(n21088), .Z(n21485) );
  XNOR U21355 ( .A(p_input[1187]), .B(n21486), .Z(n21088) );
  AND U21356 ( .A(n703), .B(n21487), .Z(n21486) );
  XOR U21357 ( .A(p_input[1203]), .B(p_input[1187]), .Z(n21487) );
  XNOR U21358 ( .A(n21085), .B(n21482), .Z(n21484) );
  XOR U21359 ( .A(n21488), .B(n21489), .Z(n21085) );
  AND U21360 ( .A(n700), .B(n21490), .Z(n21489) );
  XOR U21361 ( .A(p_input[1171]), .B(p_input[1155]), .Z(n21490) );
  XOR U21362 ( .A(n21491), .B(n21492), .Z(n21482) );
  AND U21363 ( .A(n21493), .B(n21494), .Z(n21492) );
  XOR U21364 ( .A(n21491), .B(n21100), .Z(n21494) );
  XNOR U21365 ( .A(p_input[1186]), .B(n21495), .Z(n21100) );
  AND U21366 ( .A(n703), .B(n21496), .Z(n21495) );
  XOR U21367 ( .A(p_input[1202]), .B(p_input[1186]), .Z(n21496) );
  XNOR U21368 ( .A(n21097), .B(n21491), .Z(n21493) );
  XOR U21369 ( .A(n21497), .B(n21498), .Z(n21097) );
  AND U21370 ( .A(n700), .B(n21499), .Z(n21498) );
  XOR U21371 ( .A(p_input[1170]), .B(p_input[1154]), .Z(n21499) );
  XOR U21372 ( .A(n21500), .B(n21501), .Z(n21491) );
  AND U21373 ( .A(n21502), .B(n21503), .Z(n21501) );
  XNOR U21374 ( .A(n21504), .B(n21113), .Z(n21503) );
  XNOR U21375 ( .A(p_input[1185]), .B(n21505), .Z(n21113) );
  AND U21376 ( .A(n703), .B(n21506), .Z(n21505) );
  XNOR U21377 ( .A(p_input[1201]), .B(n21507), .Z(n21506) );
  IV U21378 ( .A(p_input[1185]), .Z(n21507) );
  XNOR U21379 ( .A(n21110), .B(n21500), .Z(n21502) );
  XNOR U21380 ( .A(p_input[1153]), .B(n21508), .Z(n21110) );
  AND U21381 ( .A(n700), .B(n21509), .Z(n21508) );
  XOR U21382 ( .A(p_input[1169]), .B(p_input[1153]), .Z(n21509) );
  IV U21383 ( .A(n21504), .Z(n21500) );
  AND U21384 ( .A(n21375), .B(n21378), .Z(n21504) );
  XOR U21385 ( .A(p_input[1184]), .B(n21510), .Z(n21378) );
  AND U21386 ( .A(n703), .B(n21511), .Z(n21510) );
  XOR U21387 ( .A(p_input[1200]), .B(p_input[1184]), .Z(n21511) );
  XOR U21388 ( .A(n21512), .B(n21513), .Z(n703) );
  AND U21389 ( .A(n21514), .B(n21515), .Z(n21513) );
  XNOR U21390 ( .A(p_input[1215]), .B(n21512), .Z(n21515) );
  XOR U21391 ( .A(n21512), .B(p_input[1199]), .Z(n21514) );
  XOR U21392 ( .A(n21516), .B(n21517), .Z(n21512) );
  AND U21393 ( .A(n21518), .B(n21519), .Z(n21517) );
  XNOR U21394 ( .A(p_input[1214]), .B(n21516), .Z(n21519) );
  XOR U21395 ( .A(n21516), .B(p_input[1198]), .Z(n21518) );
  XOR U21396 ( .A(n21520), .B(n21521), .Z(n21516) );
  AND U21397 ( .A(n21522), .B(n21523), .Z(n21521) );
  XNOR U21398 ( .A(p_input[1213]), .B(n21520), .Z(n21523) );
  XOR U21399 ( .A(n21520), .B(p_input[1197]), .Z(n21522) );
  XOR U21400 ( .A(n21524), .B(n21525), .Z(n21520) );
  AND U21401 ( .A(n21526), .B(n21527), .Z(n21525) );
  XNOR U21402 ( .A(p_input[1212]), .B(n21524), .Z(n21527) );
  XOR U21403 ( .A(n21524), .B(p_input[1196]), .Z(n21526) );
  XOR U21404 ( .A(n21528), .B(n21529), .Z(n21524) );
  AND U21405 ( .A(n21530), .B(n21531), .Z(n21529) );
  XNOR U21406 ( .A(p_input[1211]), .B(n21528), .Z(n21531) );
  XOR U21407 ( .A(n21528), .B(p_input[1195]), .Z(n21530) );
  XOR U21408 ( .A(n21532), .B(n21533), .Z(n21528) );
  AND U21409 ( .A(n21534), .B(n21535), .Z(n21533) );
  XNOR U21410 ( .A(p_input[1210]), .B(n21532), .Z(n21535) );
  XOR U21411 ( .A(n21532), .B(p_input[1194]), .Z(n21534) );
  XOR U21412 ( .A(n21536), .B(n21537), .Z(n21532) );
  AND U21413 ( .A(n21538), .B(n21539), .Z(n21537) );
  XNOR U21414 ( .A(p_input[1209]), .B(n21536), .Z(n21539) );
  XOR U21415 ( .A(n21536), .B(p_input[1193]), .Z(n21538) );
  XOR U21416 ( .A(n21540), .B(n21541), .Z(n21536) );
  AND U21417 ( .A(n21542), .B(n21543), .Z(n21541) );
  XNOR U21418 ( .A(p_input[1208]), .B(n21540), .Z(n21543) );
  XOR U21419 ( .A(n21540), .B(p_input[1192]), .Z(n21542) );
  XOR U21420 ( .A(n21544), .B(n21545), .Z(n21540) );
  AND U21421 ( .A(n21546), .B(n21547), .Z(n21545) );
  XNOR U21422 ( .A(p_input[1207]), .B(n21544), .Z(n21547) );
  XOR U21423 ( .A(n21544), .B(p_input[1191]), .Z(n21546) );
  XOR U21424 ( .A(n21548), .B(n21549), .Z(n21544) );
  AND U21425 ( .A(n21550), .B(n21551), .Z(n21549) );
  XNOR U21426 ( .A(p_input[1206]), .B(n21548), .Z(n21551) );
  XOR U21427 ( .A(n21548), .B(p_input[1190]), .Z(n21550) );
  XOR U21428 ( .A(n21552), .B(n21553), .Z(n21548) );
  AND U21429 ( .A(n21554), .B(n21555), .Z(n21553) );
  XNOR U21430 ( .A(p_input[1205]), .B(n21552), .Z(n21555) );
  XOR U21431 ( .A(n21552), .B(p_input[1189]), .Z(n21554) );
  XOR U21432 ( .A(n21556), .B(n21557), .Z(n21552) );
  AND U21433 ( .A(n21558), .B(n21559), .Z(n21557) );
  XNOR U21434 ( .A(p_input[1204]), .B(n21556), .Z(n21559) );
  XOR U21435 ( .A(n21556), .B(p_input[1188]), .Z(n21558) );
  XOR U21436 ( .A(n21560), .B(n21561), .Z(n21556) );
  AND U21437 ( .A(n21562), .B(n21563), .Z(n21561) );
  XNOR U21438 ( .A(p_input[1203]), .B(n21560), .Z(n21563) );
  XOR U21439 ( .A(n21560), .B(p_input[1187]), .Z(n21562) );
  XOR U21440 ( .A(n21564), .B(n21565), .Z(n21560) );
  AND U21441 ( .A(n21566), .B(n21567), .Z(n21565) );
  XNOR U21442 ( .A(p_input[1202]), .B(n21564), .Z(n21567) );
  XOR U21443 ( .A(n21564), .B(p_input[1186]), .Z(n21566) );
  XNOR U21444 ( .A(n21568), .B(n21569), .Z(n21564) );
  AND U21445 ( .A(n21570), .B(n21571), .Z(n21569) );
  XOR U21446 ( .A(p_input[1201]), .B(n21568), .Z(n21571) );
  XNOR U21447 ( .A(p_input[1185]), .B(n21568), .Z(n21570) );
  AND U21448 ( .A(p_input[1200]), .B(n21572), .Z(n21568) );
  IV U21449 ( .A(p_input[1184]), .Z(n21572) );
  XNOR U21450 ( .A(p_input[1152]), .B(n21573), .Z(n21375) );
  AND U21451 ( .A(n700), .B(n21574), .Z(n21573) );
  XOR U21452 ( .A(p_input[1168]), .B(p_input[1152]), .Z(n21574) );
  XOR U21453 ( .A(n21575), .B(n21576), .Z(n700) );
  AND U21454 ( .A(n21577), .B(n21578), .Z(n21576) );
  XNOR U21455 ( .A(p_input[1183]), .B(n21575), .Z(n21578) );
  XOR U21456 ( .A(n21575), .B(p_input[1167]), .Z(n21577) );
  XOR U21457 ( .A(n21579), .B(n21580), .Z(n21575) );
  AND U21458 ( .A(n21581), .B(n21582), .Z(n21580) );
  XNOR U21459 ( .A(p_input[1182]), .B(n21579), .Z(n21582) );
  XNOR U21460 ( .A(n21579), .B(n21389), .Z(n21581) );
  IV U21461 ( .A(p_input[1166]), .Z(n21389) );
  XOR U21462 ( .A(n21583), .B(n21584), .Z(n21579) );
  AND U21463 ( .A(n21585), .B(n21586), .Z(n21584) );
  XNOR U21464 ( .A(p_input[1181]), .B(n21583), .Z(n21586) );
  XNOR U21465 ( .A(n21583), .B(n21398), .Z(n21585) );
  IV U21466 ( .A(p_input[1165]), .Z(n21398) );
  XOR U21467 ( .A(n21587), .B(n21588), .Z(n21583) );
  AND U21468 ( .A(n21589), .B(n21590), .Z(n21588) );
  XNOR U21469 ( .A(p_input[1180]), .B(n21587), .Z(n21590) );
  XNOR U21470 ( .A(n21587), .B(n21407), .Z(n21589) );
  IV U21471 ( .A(p_input[1164]), .Z(n21407) );
  XOR U21472 ( .A(n21591), .B(n21592), .Z(n21587) );
  AND U21473 ( .A(n21593), .B(n21594), .Z(n21592) );
  XNOR U21474 ( .A(p_input[1179]), .B(n21591), .Z(n21594) );
  XNOR U21475 ( .A(n21591), .B(n21416), .Z(n21593) );
  IV U21476 ( .A(p_input[1163]), .Z(n21416) );
  XOR U21477 ( .A(n21595), .B(n21596), .Z(n21591) );
  AND U21478 ( .A(n21597), .B(n21598), .Z(n21596) );
  XNOR U21479 ( .A(p_input[1178]), .B(n21595), .Z(n21598) );
  XNOR U21480 ( .A(n21595), .B(n21425), .Z(n21597) );
  IV U21481 ( .A(p_input[1162]), .Z(n21425) );
  XOR U21482 ( .A(n21599), .B(n21600), .Z(n21595) );
  AND U21483 ( .A(n21601), .B(n21602), .Z(n21600) );
  XNOR U21484 ( .A(p_input[1177]), .B(n21599), .Z(n21602) );
  XNOR U21485 ( .A(n21599), .B(n21434), .Z(n21601) );
  IV U21486 ( .A(p_input[1161]), .Z(n21434) );
  XOR U21487 ( .A(n21603), .B(n21604), .Z(n21599) );
  AND U21488 ( .A(n21605), .B(n21606), .Z(n21604) );
  XNOR U21489 ( .A(p_input[1176]), .B(n21603), .Z(n21606) );
  XNOR U21490 ( .A(n21603), .B(n21443), .Z(n21605) );
  IV U21491 ( .A(p_input[1160]), .Z(n21443) );
  XOR U21492 ( .A(n21607), .B(n21608), .Z(n21603) );
  AND U21493 ( .A(n21609), .B(n21610), .Z(n21608) );
  XNOR U21494 ( .A(p_input[1175]), .B(n21607), .Z(n21610) );
  XNOR U21495 ( .A(n21607), .B(n21452), .Z(n21609) );
  IV U21496 ( .A(p_input[1159]), .Z(n21452) );
  XOR U21497 ( .A(n21611), .B(n21612), .Z(n21607) );
  AND U21498 ( .A(n21613), .B(n21614), .Z(n21612) );
  XNOR U21499 ( .A(p_input[1174]), .B(n21611), .Z(n21614) );
  XNOR U21500 ( .A(n21611), .B(n21461), .Z(n21613) );
  IV U21501 ( .A(p_input[1158]), .Z(n21461) );
  XOR U21502 ( .A(n21615), .B(n21616), .Z(n21611) );
  AND U21503 ( .A(n21617), .B(n21618), .Z(n21616) );
  XNOR U21504 ( .A(p_input[1173]), .B(n21615), .Z(n21618) );
  XNOR U21505 ( .A(n21615), .B(n21470), .Z(n21617) );
  IV U21506 ( .A(p_input[1157]), .Z(n21470) );
  XOR U21507 ( .A(n21619), .B(n21620), .Z(n21615) );
  AND U21508 ( .A(n21621), .B(n21622), .Z(n21620) );
  XNOR U21509 ( .A(p_input[1172]), .B(n21619), .Z(n21622) );
  XNOR U21510 ( .A(n21619), .B(n21479), .Z(n21621) );
  IV U21511 ( .A(p_input[1156]), .Z(n21479) );
  XOR U21512 ( .A(n21623), .B(n21624), .Z(n21619) );
  AND U21513 ( .A(n21625), .B(n21626), .Z(n21624) );
  XNOR U21514 ( .A(p_input[1171]), .B(n21623), .Z(n21626) );
  XNOR U21515 ( .A(n21623), .B(n21488), .Z(n21625) );
  IV U21516 ( .A(p_input[1155]), .Z(n21488) );
  XOR U21517 ( .A(n21627), .B(n21628), .Z(n21623) );
  AND U21518 ( .A(n21629), .B(n21630), .Z(n21628) );
  XNOR U21519 ( .A(p_input[1170]), .B(n21627), .Z(n21630) );
  XNOR U21520 ( .A(n21627), .B(n21497), .Z(n21629) );
  IV U21521 ( .A(p_input[1154]), .Z(n21497) );
  XNOR U21522 ( .A(n21631), .B(n21632), .Z(n21627) );
  AND U21523 ( .A(n21633), .B(n21634), .Z(n21632) );
  XOR U21524 ( .A(p_input[1169]), .B(n21631), .Z(n21634) );
  XNOR U21525 ( .A(p_input[1153]), .B(n21631), .Z(n21633) );
  AND U21526 ( .A(p_input[1168]), .B(n21635), .Z(n21631) );
  IV U21527 ( .A(p_input[1152]), .Z(n21635) );
  XOR U21528 ( .A(n21636), .B(n21637), .Z(n20751) );
  AND U21529 ( .A(n808), .B(n21638), .Z(n21637) );
  XNOR U21530 ( .A(n21639), .B(n21636), .Z(n21638) );
  XOR U21531 ( .A(n21640), .B(n21641), .Z(n808) );
  AND U21532 ( .A(n21642), .B(n21643), .Z(n21641) );
  XNOR U21533 ( .A(n20763), .B(n21640), .Z(n21643) );
  AND U21534 ( .A(n21644), .B(n21645), .Z(n20763) );
  XOR U21535 ( .A(n21640), .B(n20762), .Z(n21642) );
  AND U21536 ( .A(n21646), .B(n21647), .Z(n20762) );
  XOR U21537 ( .A(n21648), .B(n21649), .Z(n21640) );
  AND U21538 ( .A(n21650), .B(n21651), .Z(n21649) );
  XOR U21539 ( .A(n21648), .B(n20775), .Z(n21651) );
  XOR U21540 ( .A(n21652), .B(n21653), .Z(n20775) );
  AND U21541 ( .A(n527), .B(n21654), .Z(n21653) );
  XOR U21542 ( .A(n21655), .B(n21652), .Z(n21654) );
  XNOR U21543 ( .A(n20772), .B(n21648), .Z(n21650) );
  XOR U21544 ( .A(n21656), .B(n21657), .Z(n20772) );
  AND U21545 ( .A(n524), .B(n21658), .Z(n21657) );
  XOR U21546 ( .A(n21659), .B(n21656), .Z(n21658) );
  XOR U21547 ( .A(n21660), .B(n21661), .Z(n21648) );
  AND U21548 ( .A(n21662), .B(n21663), .Z(n21661) );
  XOR U21549 ( .A(n21660), .B(n20787), .Z(n21663) );
  XOR U21550 ( .A(n21664), .B(n21665), .Z(n20787) );
  AND U21551 ( .A(n527), .B(n21666), .Z(n21665) );
  XOR U21552 ( .A(n21667), .B(n21664), .Z(n21666) );
  XNOR U21553 ( .A(n20784), .B(n21660), .Z(n21662) );
  XOR U21554 ( .A(n21668), .B(n21669), .Z(n20784) );
  AND U21555 ( .A(n524), .B(n21670), .Z(n21669) );
  XOR U21556 ( .A(n21671), .B(n21668), .Z(n21670) );
  XOR U21557 ( .A(n21672), .B(n21673), .Z(n21660) );
  AND U21558 ( .A(n21674), .B(n21675), .Z(n21673) );
  XOR U21559 ( .A(n21672), .B(n20799), .Z(n21675) );
  XOR U21560 ( .A(n21676), .B(n21677), .Z(n20799) );
  AND U21561 ( .A(n527), .B(n21678), .Z(n21677) );
  XOR U21562 ( .A(n21679), .B(n21676), .Z(n21678) );
  XNOR U21563 ( .A(n20796), .B(n21672), .Z(n21674) );
  XOR U21564 ( .A(n21680), .B(n21681), .Z(n20796) );
  AND U21565 ( .A(n524), .B(n21682), .Z(n21681) );
  XOR U21566 ( .A(n21683), .B(n21680), .Z(n21682) );
  XOR U21567 ( .A(n21684), .B(n21685), .Z(n21672) );
  AND U21568 ( .A(n21686), .B(n21687), .Z(n21685) );
  XOR U21569 ( .A(n21684), .B(n20811), .Z(n21687) );
  XOR U21570 ( .A(n21688), .B(n21689), .Z(n20811) );
  AND U21571 ( .A(n527), .B(n21690), .Z(n21689) );
  XOR U21572 ( .A(n21691), .B(n21688), .Z(n21690) );
  XNOR U21573 ( .A(n20808), .B(n21684), .Z(n21686) );
  XOR U21574 ( .A(n21692), .B(n21693), .Z(n20808) );
  AND U21575 ( .A(n524), .B(n21694), .Z(n21693) );
  XOR U21576 ( .A(n21695), .B(n21692), .Z(n21694) );
  XOR U21577 ( .A(n21696), .B(n21697), .Z(n21684) );
  AND U21578 ( .A(n21698), .B(n21699), .Z(n21697) );
  XOR U21579 ( .A(n21696), .B(n20823), .Z(n21699) );
  XOR U21580 ( .A(n21700), .B(n21701), .Z(n20823) );
  AND U21581 ( .A(n527), .B(n21702), .Z(n21701) );
  XOR U21582 ( .A(n21703), .B(n21700), .Z(n21702) );
  XNOR U21583 ( .A(n20820), .B(n21696), .Z(n21698) );
  XOR U21584 ( .A(n21704), .B(n21705), .Z(n20820) );
  AND U21585 ( .A(n524), .B(n21706), .Z(n21705) );
  XOR U21586 ( .A(n21707), .B(n21704), .Z(n21706) );
  XOR U21587 ( .A(n21708), .B(n21709), .Z(n21696) );
  AND U21588 ( .A(n21710), .B(n21711), .Z(n21709) );
  XOR U21589 ( .A(n21708), .B(n20835), .Z(n21711) );
  XOR U21590 ( .A(n21712), .B(n21713), .Z(n20835) );
  AND U21591 ( .A(n527), .B(n21714), .Z(n21713) );
  XOR U21592 ( .A(n21715), .B(n21712), .Z(n21714) );
  XNOR U21593 ( .A(n20832), .B(n21708), .Z(n21710) );
  XOR U21594 ( .A(n21716), .B(n21717), .Z(n20832) );
  AND U21595 ( .A(n524), .B(n21718), .Z(n21717) );
  XOR U21596 ( .A(n21719), .B(n21716), .Z(n21718) );
  XOR U21597 ( .A(n21720), .B(n21721), .Z(n21708) );
  AND U21598 ( .A(n21722), .B(n21723), .Z(n21721) );
  XOR U21599 ( .A(n21720), .B(n20847), .Z(n21723) );
  XOR U21600 ( .A(n21724), .B(n21725), .Z(n20847) );
  AND U21601 ( .A(n527), .B(n21726), .Z(n21725) );
  XOR U21602 ( .A(n21727), .B(n21724), .Z(n21726) );
  XNOR U21603 ( .A(n20844), .B(n21720), .Z(n21722) );
  XOR U21604 ( .A(n21728), .B(n21729), .Z(n20844) );
  AND U21605 ( .A(n524), .B(n21730), .Z(n21729) );
  XOR U21606 ( .A(n21731), .B(n21728), .Z(n21730) );
  XOR U21607 ( .A(n21732), .B(n21733), .Z(n21720) );
  AND U21608 ( .A(n21734), .B(n21735), .Z(n21733) );
  XOR U21609 ( .A(n21732), .B(n20859), .Z(n21735) );
  XOR U21610 ( .A(n21736), .B(n21737), .Z(n20859) );
  AND U21611 ( .A(n527), .B(n21738), .Z(n21737) );
  XOR U21612 ( .A(n21739), .B(n21736), .Z(n21738) );
  XNOR U21613 ( .A(n20856), .B(n21732), .Z(n21734) );
  XOR U21614 ( .A(n21740), .B(n21741), .Z(n20856) );
  AND U21615 ( .A(n524), .B(n21742), .Z(n21741) );
  XOR U21616 ( .A(n21743), .B(n21740), .Z(n21742) );
  XOR U21617 ( .A(n21744), .B(n21745), .Z(n21732) );
  AND U21618 ( .A(n21746), .B(n21747), .Z(n21745) );
  XOR U21619 ( .A(n21744), .B(n20871), .Z(n21747) );
  XOR U21620 ( .A(n21748), .B(n21749), .Z(n20871) );
  AND U21621 ( .A(n527), .B(n21750), .Z(n21749) );
  XOR U21622 ( .A(n21751), .B(n21748), .Z(n21750) );
  XNOR U21623 ( .A(n20868), .B(n21744), .Z(n21746) );
  XOR U21624 ( .A(n21752), .B(n21753), .Z(n20868) );
  AND U21625 ( .A(n524), .B(n21754), .Z(n21753) );
  XOR U21626 ( .A(n21755), .B(n21752), .Z(n21754) );
  XOR U21627 ( .A(n21756), .B(n21757), .Z(n21744) );
  AND U21628 ( .A(n21758), .B(n21759), .Z(n21757) );
  XOR U21629 ( .A(n21756), .B(n20883), .Z(n21759) );
  XOR U21630 ( .A(n21760), .B(n21761), .Z(n20883) );
  AND U21631 ( .A(n527), .B(n21762), .Z(n21761) );
  XOR U21632 ( .A(n21763), .B(n21760), .Z(n21762) );
  XNOR U21633 ( .A(n20880), .B(n21756), .Z(n21758) );
  XOR U21634 ( .A(n21764), .B(n21765), .Z(n20880) );
  AND U21635 ( .A(n524), .B(n21766), .Z(n21765) );
  XOR U21636 ( .A(n21767), .B(n21764), .Z(n21766) );
  XOR U21637 ( .A(n21768), .B(n21769), .Z(n21756) );
  AND U21638 ( .A(n21770), .B(n21771), .Z(n21769) );
  XOR U21639 ( .A(n21768), .B(n20895), .Z(n21771) );
  XOR U21640 ( .A(n21772), .B(n21773), .Z(n20895) );
  AND U21641 ( .A(n527), .B(n21774), .Z(n21773) );
  XOR U21642 ( .A(n21775), .B(n21772), .Z(n21774) );
  XNOR U21643 ( .A(n20892), .B(n21768), .Z(n21770) );
  XOR U21644 ( .A(n21776), .B(n21777), .Z(n20892) );
  AND U21645 ( .A(n524), .B(n21778), .Z(n21777) );
  XOR U21646 ( .A(n21779), .B(n21776), .Z(n21778) );
  XOR U21647 ( .A(n21780), .B(n21781), .Z(n21768) );
  AND U21648 ( .A(n21782), .B(n21783), .Z(n21781) );
  XOR U21649 ( .A(n21780), .B(n20907), .Z(n21783) );
  XOR U21650 ( .A(n21784), .B(n21785), .Z(n20907) );
  AND U21651 ( .A(n527), .B(n21786), .Z(n21785) );
  XOR U21652 ( .A(n21787), .B(n21784), .Z(n21786) );
  XNOR U21653 ( .A(n20904), .B(n21780), .Z(n21782) );
  XOR U21654 ( .A(n21788), .B(n21789), .Z(n20904) );
  AND U21655 ( .A(n524), .B(n21790), .Z(n21789) );
  XOR U21656 ( .A(n21791), .B(n21788), .Z(n21790) );
  XOR U21657 ( .A(n21792), .B(n21793), .Z(n21780) );
  AND U21658 ( .A(n21794), .B(n21795), .Z(n21793) );
  XOR U21659 ( .A(n21792), .B(n20919), .Z(n21795) );
  XOR U21660 ( .A(n21796), .B(n21797), .Z(n20919) );
  AND U21661 ( .A(n527), .B(n21798), .Z(n21797) );
  XOR U21662 ( .A(n21799), .B(n21796), .Z(n21798) );
  XNOR U21663 ( .A(n20916), .B(n21792), .Z(n21794) );
  XOR U21664 ( .A(n21800), .B(n21801), .Z(n20916) );
  AND U21665 ( .A(n524), .B(n21802), .Z(n21801) );
  XOR U21666 ( .A(n21803), .B(n21800), .Z(n21802) );
  XOR U21667 ( .A(n21804), .B(n21805), .Z(n21792) );
  AND U21668 ( .A(n21806), .B(n21807), .Z(n21805) );
  XNOR U21669 ( .A(n21808), .B(n20932), .Z(n21807) );
  XOR U21670 ( .A(n21809), .B(n21810), .Z(n20932) );
  AND U21671 ( .A(n527), .B(n21811), .Z(n21810) );
  XOR U21672 ( .A(n21809), .B(n21812), .Z(n21811) );
  XNOR U21673 ( .A(n20929), .B(n21804), .Z(n21806) );
  XOR U21674 ( .A(n21813), .B(n21814), .Z(n20929) );
  AND U21675 ( .A(n524), .B(n21815), .Z(n21814) );
  XOR U21676 ( .A(n21813), .B(n21816), .Z(n21815) );
  IV U21677 ( .A(n21808), .Z(n21804) );
  AND U21678 ( .A(n21636), .B(n21639), .Z(n21808) );
  XNOR U21679 ( .A(n21817), .B(n21818), .Z(n21639) );
  AND U21680 ( .A(n527), .B(n21819), .Z(n21818) );
  XNOR U21681 ( .A(n21820), .B(n21817), .Z(n21819) );
  XOR U21682 ( .A(n21821), .B(n21822), .Z(n527) );
  AND U21683 ( .A(n21823), .B(n21824), .Z(n21822) );
  XNOR U21684 ( .A(n21644), .B(n21821), .Z(n21824) );
  AND U21685 ( .A(p_input[1151]), .B(p_input[1135]), .Z(n21644) );
  XOR U21686 ( .A(n21821), .B(n21645), .Z(n21823) );
  AND U21687 ( .A(p_input[1119]), .B(p_input[1103]), .Z(n21645) );
  XOR U21688 ( .A(n21825), .B(n21826), .Z(n21821) );
  AND U21689 ( .A(n21827), .B(n21828), .Z(n21826) );
  XOR U21690 ( .A(n21825), .B(n21655), .Z(n21828) );
  XNOR U21691 ( .A(p_input[1134]), .B(n21829), .Z(n21655) );
  AND U21692 ( .A(n711), .B(n21830), .Z(n21829) );
  XOR U21693 ( .A(p_input[1150]), .B(p_input[1134]), .Z(n21830) );
  XNOR U21694 ( .A(n21652), .B(n21825), .Z(n21827) );
  XOR U21695 ( .A(n21831), .B(n21832), .Z(n21652) );
  AND U21696 ( .A(n709), .B(n21833), .Z(n21832) );
  XOR U21697 ( .A(p_input[1118]), .B(p_input[1102]), .Z(n21833) );
  XOR U21698 ( .A(n21834), .B(n21835), .Z(n21825) );
  AND U21699 ( .A(n21836), .B(n21837), .Z(n21835) );
  XOR U21700 ( .A(n21834), .B(n21667), .Z(n21837) );
  XNOR U21701 ( .A(p_input[1133]), .B(n21838), .Z(n21667) );
  AND U21702 ( .A(n711), .B(n21839), .Z(n21838) );
  XOR U21703 ( .A(p_input[1149]), .B(p_input[1133]), .Z(n21839) );
  XNOR U21704 ( .A(n21664), .B(n21834), .Z(n21836) );
  XOR U21705 ( .A(n21840), .B(n21841), .Z(n21664) );
  AND U21706 ( .A(n709), .B(n21842), .Z(n21841) );
  XOR U21707 ( .A(p_input[1117]), .B(p_input[1101]), .Z(n21842) );
  XOR U21708 ( .A(n21843), .B(n21844), .Z(n21834) );
  AND U21709 ( .A(n21845), .B(n21846), .Z(n21844) );
  XOR U21710 ( .A(n21843), .B(n21679), .Z(n21846) );
  XNOR U21711 ( .A(p_input[1132]), .B(n21847), .Z(n21679) );
  AND U21712 ( .A(n711), .B(n21848), .Z(n21847) );
  XOR U21713 ( .A(p_input[1148]), .B(p_input[1132]), .Z(n21848) );
  XNOR U21714 ( .A(n21676), .B(n21843), .Z(n21845) );
  XOR U21715 ( .A(n21849), .B(n21850), .Z(n21676) );
  AND U21716 ( .A(n709), .B(n21851), .Z(n21850) );
  XOR U21717 ( .A(p_input[1116]), .B(p_input[1100]), .Z(n21851) );
  XOR U21718 ( .A(n21852), .B(n21853), .Z(n21843) );
  AND U21719 ( .A(n21854), .B(n21855), .Z(n21853) );
  XOR U21720 ( .A(n21852), .B(n21691), .Z(n21855) );
  XNOR U21721 ( .A(p_input[1131]), .B(n21856), .Z(n21691) );
  AND U21722 ( .A(n711), .B(n21857), .Z(n21856) );
  XOR U21723 ( .A(p_input[1147]), .B(p_input[1131]), .Z(n21857) );
  XNOR U21724 ( .A(n21688), .B(n21852), .Z(n21854) );
  XOR U21725 ( .A(n21858), .B(n21859), .Z(n21688) );
  AND U21726 ( .A(n709), .B(n21860), .Z(n21859) );
  XOR U21727 ( .A(p_input[1115]), .B(p_input[1099]), .Z(n21860) );
  XOR U21728 ( .A(n21861), .B(n21862), .Z(n21852) );
  AND U21729 ( .A(n21863), .B(n21864), .Z(n21862) );
  XOR U21730 ( .A(n21861), .B(n21703), .Z(n21864) );
  XNOR U21731 ( .A(p_input[1130]), .B(n21865), .Z(n21703) );
  AND U21732 ( .A(n711), .B(n21866), .Z(n21865) );
  XOR U21733 ( .A(p_input[1146]), .B(p_input[1130]), .Z(n21866) );
  XNOR U21734 ( .A(n21700), .B(n21861), .Z(n21863) );
  XOR U21735 ( .A(n21867), .B(n21868), .Z(n21700) );
  AND U21736 ( .A(n709), .B(n21869), .Z(n21868) );
  XOR U21737 ( .A(p_input[1114]), .B(p_input[1098]), .Z(n21869) );
  XOR U21738 ( .A(n21870), .B(n21871), .Z(n21861) );
  AND U21739 ( .A(n21872), .B(n21873), .Z(n21871) );
  XOR U21740 ( .A(n21870), .B(n21715), .Z(n21873) );
  XNOR U21741 ( .A(p_input[1129]), .B(n21874), .Z(n21715) );
  AND U21742 ( .A(n711), .B(n21875), .Z(n21874) );
  XOR U21743 ( .A(p_input[1145]), .B(p_input[1129]), .Z(n21875) );
  XNOR U21744 ( .A(n21712), .B(n21870), .Z(n21872) );
  XOR U21745 ( .A(n21876), .B(n21877), .Z(n21712) );
  AND U21746 ( .A(n709), .B(n21878), .Z(n21877) );
  XOR U21747 ( .A(p_input[1113]), .B(p_input[1097]), .Z(n21878) );
  XOR U21748 ( .A(n21879), .B(n21880), .Z(n21870) );
  AND U21749 ( .A(n21881), .B(n21882), .Z(n21880) );
  XOR U21750 ( .A(n21879), .B(n21727), .Z(n21882) );
  XNOR U21751 ( .A(p_input[1128]), .B(n21883), .Z(n21727) );
  AND U21752 ( .A(n711), .B(n21884), .Z(n21883) );
  XOR U21753 ( .A(p_input[1144]), .B(p_input[1128]), .Z(n21884) );
  XNOR U21754 ( .A(n21724), .B(n21879), .Z(n21881) );
  XOR U21755 ( .A(n21885), .B(n21886), .Z(n21724) );
  AND U21756 ( .A(n709), .B(n21887), .Z(n21886) );
  XOR U21757 ( .A(p_input[1112]), .B(p_input[1096]), .Z(n21887) );
  XOR U21758 ( .A(n21888), .B(n21889), .Z(n21879) );
  AND U21759 ( .A(n21890), .B(n21891), .Z(n21889) );
  XOR U21760 ( .A(n21888), .B(n21739), .Z(n21891) );
  XNOR U21761 ( .A(p_input[1127]), .B(n21892), .Z(n21739) );
  AND U21762 ( .A(n711), .B(n21893), .Z(n21892) );
  XOR U21763 ( .A(p_input[1143]), .B(p_input[1127]), .Z(n21893) );
  XNOR U21764 ( .A(n21736), .B(n21888), .Z(n21890) );
  XOR U21765 ( .A(n21894), .B(n21895), .Z(n21736) );
  AND U21766 ( .A(n709), .B(n21896), .Z(n21895) );
  XOR U21767 ( .A(p_input[1111]), .B(p_input[1095]), .Z(n21896) );
  XOR U21768 ( .A(n21897), .B(n21898), .Z(n21888) );
  AND U21769 ( .A(n21899), .B(n21900), .Z(n21898) );
  XOR U21770 ( .A(n21897), .B(n21751), .Z(n21900) );
  XNOR U21771 ( .A(p_input[1126]), .B(n21901), .Z(n21751) );
  AND U21772 ( .A(n711), .B(n21902), .Z(n21901) );
  XOR U21773 ( .A(p_input[1142]), .B(p_input[1126]), .Z(n21902) );
  XNOR U21774 ( .A(n21748), .B(n21897), .Z(n21899) );
  XOR U21775 ( .A(n21903), .B(n21904), .Z(n21748) );
  AND U21776 ( .A(n709), .B(n21905), .Z(n21904) );
  XOR U21777 ( .A(p_input[1110]), .B(p_input[1094]), .Z(n21905) );
  XOR U21778 ( .A(n21906), .B(n21907), .Z(n21897) );
  AND U21779 ( .A(n21908), .B(n21909), .Z(n21907) );
  XOR U21780 ( .A(n21906), .B(n21763), .Z(n21909) );
  XNOR U21781 ( .A(p_input[1125]), .B(n21910), .Z(n21763) );
  AND U21782 ( .A(n711), .B(n21911), .Z(n21910) );
  XOR U21783 ( .A(p_input[1141]), .B(p_input[1125]), .Z(n21911) );
  XNOR U21784 ( .A(n21760), .B(n21906), .Z(n21908) );
  XOR U21785 ( .A(n21912), .B(n21913), .Z(n21760) );
  AND U21786 ( .A(n709), .B(n21914), .Z(n21913) );
  XOR U21787 ( .A(p_input[1109]), .B(p_input[1093]), .Z(n21914) );
  XOR U21788 ( .A(n21915), .B(n21916), .Z(n21906) );
  AND U21789 ( .A(n21917), .B(n21918), .Z(n21916) );
  XOR U21790 ( .A(n21915), .B(n21775), .Z(n21918) );
  XNOR U21791 ( .A(p_input[1124]), .B(n21919), .Z(n21775) );
  AND U21792 ( .A(n711), .B(n21920), .Z(n21919) );
  XOR U21793 ( .A(p_input[1140]), .B(p_input[1124]), .Z(n21920) );
  XNOR U21794 ( .A(n21772), .B(n21915), .Z(n21917) );
  XOR U21795 ( .A(n21921), .B(n21922), .Z(n21772) );
  AND U21796 ( .A(n709), .B(n21923), .Z(n21922) );
  XOR U21797 ( .A(p_input[1108]), .B(p_input[1092]), .Z(n21923) );
  XOR U21798 ( .A(n21924), .B(n21925), .Z(n21915) );
  AND U21799 ( .A(n21926), .B(n21927), .Z(n21925) );
  XOR U21800 ( .A(n21924), .B(n21787), .Z(n21927) );
  XNOR U21801 ( .A(p_input[1123]), .B(n21928), .Z(n21787) );
  AND U21802 ( .A(n711), .B(n21929), .Z(n21928) );
  XOR U21803 ( .A(p_input[1139]), .B(p_input[1123]), .Z(n21929) );
  XNOR U21804 ( .A(n21784), .B(n21924), .Z(n21926) );
  XOR U21805 ( .A(n21930), .B(n21931), .Z(n21784) );
  AND U21806 ( .A(n709), .B(n21932), .Z(n21931) );
  XOR U21807 ( .A(p_input[1107]), .B(p_input[1091]), .Z(n21932) );
  XOR U21808 ( .A(n21933), .B(n21934), .Z(n21924) );
  AND U21809 ( .A(n21935), .B(n21936), .Z(n21934) );
  XOR U21810 ( .A(n21933), .B(n21799), .Z(n21936) );
  XNOR U21811 ( .A(p_input[1122]), .B(n21937), .Z(n21799) );
  AND U21812 ( .A(n711), .B(n21938), .Z(n21937) );
  XOR U21813 ( .A(p_input[1138]), .B(p_input[1122]), .Z(n21938) );
  XNOR U21814 ( .A(n21796), .B(n21933), .Z(n21935) );
  XOR U21815 ( .A(n21939), .B(n21940), .Z(n21796) );
  AND U21816 ( .A(n709), .B(n21941), .Z(n21940) );
  XOR U21817 ( .A(p_input[1106]), .B(p_input[1090]), .Z(n21941) );
  XOR U21818 ( .A(n21942), .B(n21943), .Z(n21933) );
  AND U21819 ( .A(n21944), .B(n21945), .Z(n21943) );
  XNOR U21820 ( .A(n21946), .B(n21812), .Z(n21945) );
  XNOR U21821 ( .A(p_input[1121]), .B(n21947), .Z(n21812) );
  AND U21822 ( .A(n711), .B(n21948), .Z(n21947) );
  XNOR U21823 ( .A(p_input[1137]), .B(n21949), .Z(n21948) );
  IV U21824 ( .A(p_input[1121]), .Z(n21949) );
  XNOR U21825 ( .A(n21809), .B(n21942), .Z(n21944) );
  XNOR U21826 ( .A(p_input[1089]), .B(n21950), .Z(n21809) );
  AND U21827 ( .A(n709), .B(n21951), .Z(n21950) );
  XOR U21828 ( .A(p_input[1105]), .B(p_input[1089]), .Z(n21951) );
  IV U21829 ( .A(n21946), .Z(n21942) );
  AND U21830 ( .A(n21817), .B(n21820), .Z(n21946) );
  XOR U21831 ( .A(p_input[1120]), .B(n21952), .Z(n21820) );
  AND U21832 ( .A(n711), .B(n21953), .Z(n21952) );
  XOR U21833 ( .A(p_input[1136]), .B(p_input[1120]), .Z(n21953) );
  XOR U21834 ( .A(n21954), .B(n21955), .Z(n711) );
  AND U21835 ( .A(n21956), .B(n21957), .Z(n21955) );
  XNOR U21836 ( .A(p_input[1151]), .B(n21954), .Z(n21957) );
  XOR U21837 ( .A(n21954), .B(p_input[1135]), .Z(n21956) );
  XOR U21838 ( .A(n21958), .B(n21959), .Z(n21954) );
  AND U21839 ( .A(n21960), .B(n21961), .Z(n21959) );
  XNOR U21840 ( .A(p_input[1150]), .B(n21958), .Z(n21961) );
  XOR U21841 ( .A(n21958), .B(p_input[1134]), .Z(n21960) );
  XOR U21842 ( .A(n21962), .B(n21963), .Z(n21958) );
  AND U21843 ( .A(n21964), .B(n21965), .Z(n21963) );
  XNOR U21844 ( .A(p_input[1149]), .B(n21962), .Z(n21965) );
  XOR U21845 ( .A(n21962), .B(p_input[1133]), .Z(n21964) );
  XOR U21846 ( .A(n21966), .B(n21967), .Z(n21962) );
  AND U21847 ( .A(n21968), .B(n21969), .Z(n21967) );
  XNOR U21848 ( .A(p_input[1148]), .B(n21966), .Z(n21969) );
  XOR U21849 ( .A(n21966), .B(p_input[1132]), .Z(n21968) );
  XOR U21850 ( .A(n21970), .B(n21971), .Z(n21966) );
  AND U21851 ( .A(n21972), .B(n21973), .Z(n21971) );
  XNOR U21852 ( .A(p_input[1147]), .B(n21970), .Z(n21973) );
  XOR U21853 ( .A(n21970), .B(p_input[1131]), .Z(n21972) );
  XOR U21854 ( .A(n21974), .B(n21975), .Z(n21970) );
  AND U21855 ( .A(n21976), .B(n21977), .Z(n21975) );
  XNOR U21856 ( .A(p_input[1146]), .B(n21974), .Z(n21977) );
  XOR U21857 ( .A(n21974), .B(p_input[1130]), .Z(n21976) );
  XOR U21858 ( .A(n21978), .B(n21979), .Z(n21974) );
  AND U21859 ( .A(n21980), .B(n21981), .Z(n21979) );
  XNOR U21860 ( .A(p_input[1145]), .B(n21978), .Z(n21981) );
  XOR U21861 ( .A(n21978), .B(p_input[1129]), .Z(n21980) );
  XOR U21862 ( .A(n21982), .B(n21983), .Z(n21978) );
  AND U21863 ( .A(n21984), .B(n21985), .Z(n21983) );
  XNOR U21864 ( .A(p_input[1144]), .B(n21982), .Z(n21985) );
  XOR U21865 ( .A(n21982), .B(p_input[1128]), .Z(n21984) );
  XOR U21866 ( .A(n21986), .B(n21987), .Z(n21982) );
  AND U21867 ( .A(n21988), .B(n21989), .Z(n21987) );
  XNOR U21868 ( .A(p_input[1143]), .B(n21986), .Z(n21989) );
  XOR U21869 ( .A(n21986), .B(p_input[1127]), .Z(n21988) );
  XOR U21870 ( .A(n21990), .B(n21991), .Z(n21986) );
  AND U21871 ( .A(n21992), .B(n21993), .Z(n21991) );
  XNOR U21872 ( .A(p_input[1142]), .B(n21990), .Z(n21993) );
  XOR U21873 ( .A(n21990), .B(p_input[1126]), .Z(n21992) );
  XOR U21874 ( .A(n21994), .B(n21995), .Z(n21990) );
  AND U21875 ( .A(n21996), .B(n21997), .Z(n21995) );
  XNOR U21876 ( .A(p_input[1141]), .B(n21994), .Z(n21997) );
  XOR U21877 ( .A(n21994), .B(p_input[1125]), .Z(n21996) );
  XOR U21878 ( .A(n21998), .B(n21999), .Z(n21994) );
  AND U21879 ( .A(n22000), .B(n22001), .Z(n21999) );
  XNOR U21880 ( .A(p_input[1140]), .B(n21998), .Z(n22001) );
  XOR U21881 ( .A(n21998), .B(p_input[1124]), .Z(n22000) );
  XOR U21882 ( .A(n22002), .B(n22003), .Z(n21998) );
  AND U21883 ( .A(n22004), .B(n22005), .Z(n22003) );
  XNOR U21884 ( .A(p_input[1139]), .B(n22002), .Z(n22005) );
  XOR U21885 ( .A(n22002), .B(p_input[1123]), .Z(n22004) );
  XOR U21886 ( .A(n22006), .B(n22007), .Z(n22002) );
  AND U21887 ( .A(n22008), .B(n22009), .Z(n22007) );
  XNOR U21888 ( .A(p_input[1138]), .B(n22006), .Z(n22009) );
  XOR U21889 ( .A(n22006), .B(p_input[1122]), .Z(n22008) );
  XNOR U21890 ( .A(n22010), .B(n22011), .Z(n22006) );
  AND U21891 ( .A(n22012), .B(n22013), .Z(n22011) );
  XOR U21892 ( .A(p_input[1137]), .B(n22010), .Z(n22013) );
  XNOR U21893 ( .A(p_input[1121]), .B(n22010), .Z(n22012) );
  AND U21894 ( .A(p_input[1136]), .B(n22014), .Z(n22010) );
  IV U21895 ( .A(p_input[1120]), .Z(n22014) );
  XNOR U21896 ( .A(p_input[1088]), .B(n22015), .Z(n21817) );
  AND U21897 ( .A(n709), .B(n22016), .Z(n22015) );
  XOR U21898 ( .A(p_input[1104]), .B(p_input[1088]), .Z(n22016) );
  XOR U21899 ( .A(n22017), .B(n22018), .Z(n709) );
  AND U21900 ( .A(n22019), .B(n22020), .Z(n22018) );
  XNOR U21901 ( .A(p_input[1119]), .B(n22017), .Z(n22020) );
  XOR U21902 ( .A(n22017), .B(p_input[1103]), .Z(n22019) );
  XOR U21903 ( .A(n22021), .B(n22022), .Z(n22017) );
  AND U21904 ( .A(n22023), .B(n22024), .Z(n22022) );
  XNOR U21905 ( .A(p_input[1118]), .B(n22021), .Z(n22024) );
  XNOR U21906 ( .A(n22021), .B(n21831), .Z(n22023) );
  IV U21907 ( .A(p_input[1102]), .Z(n21831) );
  XOR U21908 ( .A(n22025), .B(n22026), .Z(n22021) );
  AND U21909 ( .A(n22027), .B(n22028), .Z(n22026) );
  XNOR U21910 ( .A(p_input[1117]), .B(n22025), .Z(n22028) );
  XNOR U21911 ( .A(n22025), .B(n21840), .Z(n22027) );
  IV U21912 ( .A(p_input[1101]), .Z(n21840) );
  XOR U21913 ( .A(n22029), .B(n22030), .Z(n22025) );
  AND U21914 ( .A(n22031), .B(n22032), .Z(n22030) );
  XNOR U21915 ( .A(p_input[1116]), .B(n22029), .Z(n22032) );
  XNOR U21916 ( .A(n22029), .B(n21849), .Z(n22031) );
  IV U21917 ( .A(p_input[1100]), .Z(n21849) );
  XOR U21918 ( .A(n22033), .B(n22034), .Z(n22029) );
  AND U21919 ( .A(n22035), .B(n22036), .Z(n22034) );
  XNOR U21920 ( .A(p_input[1115]), .B(n22033), .Z(n22036) );
  XNOR U21921 ( .A(n22033), .B(n21858), .Z(n22035) );
  IV U21922 ( .A(p_input[1099]), .Z(n21858) );
  XOR U21923 ( .A(n22037), .B(n22038), .Z(n22033) );
  AND U21924 ( .A(n22039), .B(n22040), .Z(n22038) );
  XNOR U21925 ( .A(p_input[1114]), .B(n22037), .Z(n22040) );
  XNOR U21926 ( .A(n22037), .B(n21867), .Z(n22039) );
  IV U21927 ( .A(p_input[1098]), .Z(n21867) );
  XOR U21928 ( .A(n22041), .B(n22042), .Z(n22037) );
  AND U21929 ( .A(n22043), .B(n22044), .Z(n22042) );
  XNOR U21930 ( .A(p_input[1113]), .B(n22041), .Z(n22044) );
  XNOR U21931 ( .A(n22041), .B(n21876), .Z(n22043) );
  IV U21932 ( .A(p_input[1097]), .Z(n21876) );
  XOR U21933 ( .A(n22045), .B(n22046), .Z(n22041) );
  AND U21934 ( .A(n22047), .B(n22048), .Z(n22046) );
  XNOR U21935 ( .A(p_input[1112]), .B(n22045), .Z(n22048) );
  XNOR U21936 ( .A(n22045), .B(n21885), .Z(n22047) );
  IV U21937 ( .A(p_input[1096]), .Z(n21885) );
  XOR U21938 ( .A(n22049), .B(n22050), .Z(n22045) );
  AND U21939 ( .A(n22051), .B(n22052), .Z(n22050) );
  XNOR U21940 ( .A(p_input[1111]), .B(n22049), .Z(n22052) );
  XNOR U21941 ( .A(n22049), .B(n21894), .Z(n22051) );
  IV U21942 ( .A(p_input[1095]), .Z(n21894) );
  XOR U21943 ( .A(n22053), .B(n22054), .Z(n22049) );
  AND U21944 ( .A(n22055), .B(n22056), .Z(n22054) );
  XNOR U21945 ( .A(p_input[1110]), .B(n22053), .Z(n22056) );
  XNOR U21946 ( .A(n22053), .B(n21903), .Z(n22055) );
  IV U21947 ( .A(p_input[1094]), .Z(n21903) );
  XOR U21948 ( .A(n22057), .B(n22058), .Z(n22053) );
  AND U21949 ( .A(n22059), .B(n22060), .Z(n22058) );
  XNOR U21950 ( .A(p_input[1109]), .B(n22057), .Z(n22060) );
  XNOR U21951 ( .A(n22057), .B(n21912), .Z(n22059) );
  IV U21952 ( .A(p_input[1093]), .Z(n21912) );
  XOR U21953 ( .A(n22061), .B(n22062), .Z(n22057) );
  AND U21954 ( .A(n22063), .B(n22064), .Z(n22062) );
  XNOR U21955 ( .A(p_input[1108]), .B(n22061), .Z(n22064) );
  XNOR U21956 ( .A(n22061), .B(n21921), .Z(n22063) );
  IV U21957 ( .A(p_input[1092]), .Z(n21921) );
  XOR U21958 ( .A(n22065), .B(n22066), .Z(n22061) );
  AND U21959 ( .A(n22067), .B(n22068), .Z(n22066) );
  XNOR U21960 ( .A(p_input[1107]), .B(n22065), .Z(n22068) );
  XNOR U21961 ( .A(n22065), .B(n21930), .Z(n22067) );
  IV U21962 ( .A(p_input[1091]), .Z(n21930) );
  XOR U21963 ( .A(n22069), .B(n22070), .Z(n22065) );
  AND U21964 ( .A(n22071), .B(n22072), .Z(n22070) );
  XNOR U21965 ( .A(p_input[1106]), .B(n22069), .Z(n22072) );
  XNOR U21966 ( .A(n22069), .B(n21939), .Z(n22071) );
  IV U21967 ( .A(p_input[1090]), .Z(n21939) );
  XNOR U21968 ( .A(n22073), .B(n22074), .Z(n22069) );
  AND U21969 ( .A(n22075), .B(n22076), .Z(n22074) );
  XOR U21970 ( .A(p_input[1105]), .B(n22073), .Z(n22076) );
  XNOR U21971 ( .A(p_input[1089]), .B(n22073), .Z(n22075) );
  AND U21972 ( .A(p_input[1104]), .B(n22077), .Z(n22073) );
  IV U21973 ( .A(p_input[1088]), .Z(n22077) );
  XOR U21974 ( .A(n22078), .B(n22079), .Z(n21636) );
  AND U21975 ( .A(n524), .B(n22080), .Z(n22079) );
  XNOR U21976 ( .A(n22081), .B(n22078), .Z(n22080) );
  XOR U21977 ( .A(n22082), .B(n22083), .Z(n524) );
  AND U21978 ( .A(n22084), .B(n22085), .Z(n22083) );
  XNOR U21979 ( .A(n21647), .B(n22082), .Z(n22085) );
  AND U21980 ( .A(p_input[1087]), .B(p_input[1071]), .Z(n21647) );
  XOR U21981 ( .A(n22082), .B(n21646), .Z(n22084) );
  AND U21982 ( .A(p_input[1039]), .B(p_input[1055]), .Z(n21646) );
  XOR U21983 ( .A(n22086), .B(n22087), .Z(n22082) );
  AND U21984 ( .A(n22088), .B(n22089), .Z(n22087) );
  XOR U21985 ( .A(n22086), .B(n21659), .Z(n22089) );
  XNOR U21986 ( .A(p_input[1070]), .B(n22090), .Z(n21659) );
  AND U21987 ( .A(n715), .B(n22091), .Z(n22090) );
  XOR U21988 ( .A(p_input[1086]), .B(p_input[1070]), .Z(n22091) );
  XNOR U21989 ( .A(n21656), .B(n22086), .Z(n22088) );
  XOR U21990 ( .A(n22092), .B(n22093), .Z(n21656) );
  AND U21991 ( .A(n712), .B(n22094), .Z(n22093) );
  XOR U21992 ( .A(p_input[1054]), .B(p_input[1038]), .Z(n22094) );
  XOR U21993 ( .A(n22095), .B(n22096), .Z(n22086) );
  AND U21994 ( .A(n22097), .B(n22098), .Z(n22096) );
  XOR U21995 ( .A(n22095), .B(n21671), .Z(n22098) );
  XNOR U21996 ( .A(p_input[1069]), .B(n22099), .Z(n21671) );
  AND U21997 ( .A(n715), .B(n22100), .Z(n22099) );
  XOR U21998 ( .A(p_input[1085]), .B(p_input[1069]), .Z(n22100) );
  XNOR U21999 ( .A(n21668), .B(n22095), .Z(n22097) );
  XOR U22000 ( .A(n22101), .B(n22102), .Z(n21668) );
  AND U22001 ( .A(n712), .B(n22103), .Z(n22102) );
  XOR U22002 ( .A(p_input[1053]), .B(p_input[1037]), .Z(n22103) );
  XOR U22003 ( .A(n22104), .B(n22105), .Z(n22095) );
  AND U22004 ( .A(n22106), .B(n22107), .Z(n22105) );
  XOR U22005 ( .A(n22104), .B(n21683), .Z(n22107) );
  XNOR U22006 ( .A(p_input[1068]), .B(n22108), .Z(n21683) );
  AND U22007 ( .A(n715), .B(n22109), .Z(n22108) );
  XOR U22008 ( .A(p_input[1084]), .B(p_input[1068]), .Z(n22109) );
  XNOR U22009 ( .A(n21680), .B(n22104), .Z(n22106) );
  XOR U22010 ( .A(n22110), .B(n22111), .Z(n21680) );
  AND U22011 ( .A(n712), .B(n22112), .Z(n22111) );
  XOR U22012 ( .A(p_input[1052]), .B(p_input[1036]), .Z(n22112) );
  XOR U22013 ( .A(n22113), .B(n22114), .Z(n22104) );
  AND U22014 ( .A(n22115), .B(n22116), .Z(n22114) );
  XOR U22015 ( .A(n22113), .B(n21695), .Z(n22116) );
  XNOR U22016 ( .A(p_input[1067]), .B(n22117), .Z(n21695) );
  AND U22017 ( .A(n715), .B(n22118), .Z(n22117) );
  XOR U22018 ( .A(p_input[1083]), .B(p_input[1067]), .Z(n22118) );
  XNOR U22019 ( .A(n21692), .B(n22113), .Z(n22115) );
  XOR U22020 ( .A(n22119), .B(n22120), .Z(n21692) );
  AND U22021 ( .A(n712), .B(n22121), .Z(n22120) );
  XOR U22022 ( .A(p_input[1051]), .B(p_input[1035]), .Z(n22121) );
  XOR U22023 ( .A(n22122), .B(n22123), .Z(n22113) );
  AND U22024 ( .A(n22124), .B(n22125), .Z(n22123) );
  XOR U22025 ( .A(n22122), .B(n21707), .Z(n22125) );
  XNOR U22026 ( .A(p_input[1066]), .B(n22126), .Z(n21707) );
  AND U22027 ( .A(n715), .B(n22127), .Z(n22126) );
  XOR U22028 ( .A(p_input[1082]), .B(p_input[1066]), .Z(n22127) );
  XNOR U22029 ( .A(n21704), .B(n22122), .Z(n22124) );
  XOR U22030 ( .A(n22128), .B(n22129), .Z(n21704) );
  AND U22031 ( .A(n712), .B(n22130), .Z(n22129) );
  XOR U22032 ( .A(p_input[1050]), .B(p_input[1034]), .Z(n22130) );
  XOR U22033 ( .A(n22131), .B(n22132), .Z(n22122) );
  AND U22034 ( .A(n22133), .B(n22134), .Z(n22132) );
  XOR U22035 ( .A(n22131), .B(n21719), .Z(n22134) );
  XNOR U22036 ( .A(p_input[1065]), .B(n22135), .Z(n21719) );
  AND U22037 ( .A(n715), .B(n22136), .Z(n22135) );
  XOR U22038 ( .A(p_input[1081]), .B(p_input[1065]), .Z(n22136) );
  XNOR U22039 ( .A(n21716), .B(n22131), .Z(n22133) );
  XOR U22040 ( .A(n22137), .B(n22138), .Z(n21716) );
  AND U22041 ( .A(n712), .B(n22139), .Z(n22138) );
  XOR U22042 ( .A(p_input[1049]), .B(p_input[1033]), .Z(n22139) );
  XOR U22043 ( .A(n22140), .B(n22141), .Z(n22131) );
  AND U22044 ( .A(n22142), .B(n22143), .Z(n22141) );
  XOR U22045 ( .A(n22140), .B(n21731), .Z(n22143) );
  XNOR U22046 ( .A(p_input[1064]), .B(n22144), .Z(n21731) );
  AND U22047 ( .A(n715), .B(n22145), .Z(n22144) );
  XOR U22048 ( .A(p_input[1080]), .B(p_input[1064]), .Z(n22145) );
  XNOR U22049 ( .A(n21728), .B(n22140), .Z(n22142) );
  XOR U22050 ( .A(n22146), .B(n22147), .Z(n21728) );
  AND U22051 ( .A(n712), .B(n22148), .Z(n22147) );
  XOR U22052 ( .A(p_input[1048]), .B(p_input[1032]), .Z(n22148) );
  XOR U22053 ( .A(n22149), .B(n22150), .Z(n22140) );
  AND U22054 ( .A(n22151), .B(n22152), .Z(n22150) );
  XOR U22055 ( .A(n22149), .B(n21743), .Z(n22152) );
  XNOR U22056 ( .A(p_input[1063]), .B(n22153), .Z(n21743) );
  AND U22057 ( .A(n715), .B(n22154), .Z(n22153) );
  XOR U22058 ( .A(p_input[1079]), .B(p_input[1063]), .Z(n22154) );
  XNOR U22059 ( .A(n21740), .B(n22149), .Z(n22151) );
  XOR U22060 ( .A(n22155), .B(n22156), .Z(n21740) );
  AND U22061 ( .A(n712), .B(n22157), .Z(n22156) );
  XOR U22062 ( .A(p_input[1047]), .B(p_input[1031]), .Z(n22157) );
  XOR U22063 ( .A(n22158), .B(n22159), .Z(n22149) );
  AND U22064 ( .A(n22160), .B(n22161), .Z(n22159) );
  XOR U22065 ( .A(n22158), .B(n21755), .Z(n22161) );
  XNOR U22066 ( .A(p_input[1062]), .B(n22162), .Z(n21755) );
  AND U22067 ( .A(n715), .B(n22163), .Z(n22162) );
  XOR U22068 ( .A(p_input[1078]), .B(p_input[1062]), .Z(n22163) );
  XNOR U22069 ( .A(n21752), .B(n22158), .Z(n22160) );
  XOR U22070 ( .A(n22164), .B(n22165), .Z(n21752) );
  AND U22071 ( .A(n712), .B(n22166), .Z(n22165) );
  XOR U22072 ( .A(p_input[1046]), .B(p_input[1030]), .Z(n22166) );
  XOR U22073 ( .A(n22167), .B(n22168), .Z(n22158) );
  AND U22074 ( .A(n22169), .B(n22170), .Z(n22168) );
  XOR U22075 ( .A(n22167), .B(n21767), .Z(n22170) );
  XNOR U22076 ( .A(p_input[1061]), .B(n22171), .Z(n21767) );
  AND U22077 ( .A(n715), .B(n22172), .Z(n22171) );
  XOR U22078 ( .A(p_input[1077]), .B(p_input[1061]), .Z(n22172) );
  XNOR U22079 ( .A(n21764), .B(n22167), .Z(n22169) );
  XOR U22080 ( .A(n22173), .B(n22174), .Z(n21764) );
  AND U22081 ( .A(n712), .B(n22175), .Z(n22174) );
  XOR U22082 ( .A(p_input[1045]), .B(p_input[1029]), .Z(n22175) );
  XOR U22083 ( .A(n22176), .B(n22177), .Z(n22167) );
  AND U22084 ( .A(n22178), .B(n22179), .Z(n22177) );
  XOR U22085 ( .A(n22176), .B(n21779), .Z(n22179) );
  XNOR U22086 ( .A(p_input[1060]), .B(n22180), .Z(n21779) );
  AND U22087 ( .A(n715), .B(n22181), .Z(n22180) );
  XOR U22088 ( .A(p_input[1076]), .B(p_input[1060]), .Z(n22181) );
  XNOR U22089 ( .A(n21776), .B(n22176), .Z(n22178) );
  XOR U22090 ( .A(n22182), .B(n22183), .Z(n21776) );
  AND U22091 ( .A(n712), .B(n22184), .Z(n22183) );
  XOR U22092 ( .A(p_input[1044]), .B(p_input[1028]), .Z(n22184) );
  XOR U22093 ( .A(n22185), .B(n22186), .Z(n22176) );
  AND U22094 ( .A(n22187), .B(n22188), .Z(n22186) );
  XOR U22095 ( .A(n22185), .B(n21791), .Z(n22188) );
  XNOR U22096 ( .A(p_input[1059]), .B(n22189), .Z(n21791) );
  AND U22097 ( .A(n715), .B(n22190), .Z(n22189) );
  XOR U22098 ( .A(p_input[1075]), .B(p_input[1059]), .Z(n22190) );
  XNOR U22099 ( .A(n21788), .B(n22185), .Z(n22187) );
  XOR U22100 ( .A(n22191), .B(n22192), .Z(n21788) );
  AND U22101 ( .A(n712), .B(n22193), .Z(n22192) );
  XOR U22102 ( .A(p_input[1043]), .B(p_input[1027]), .Z(n22193) );
  XOR U22103 ( .A(n22194), .B(n22195), .Z(n22185) );
  AND U22104 ( .A(n22196), .B(n22197), .Z(n22195) );
  XOR U22105 ( .A(n22194), .B(n21803), .Z(n22197) );
  XNOR U22106 ( .A(p_input[1058]), .B(n22198), .Z(n21803) );
  AND U22107 ( .A(n715), .B(n22199), .Z(n22198) );
  XOR U22108 ( .A(p_input[1074]), .B(p_input[1058]), .Z(n22199) );
  XNOR U22109 ( .A(n21800), .B(n22194), .Z(n22196) );
  XOR U22110 ( .A(n22200), .B(n22201), .Z(n21800) );
  AND U22111 ( .A(n712), .B(n22202), .Z(n22201) );
  XOR U22112 ( .A(p_input[1042]), .B(p_input[1026]), .Z(n22202) );
  XOR U22113 ( .A(n22203), .B(n22204), .Z(n22194) );
  AND U22114 ( .A(n22205), .B(n22206), .Z(n22204) );
  XNOR U22115 ( .A(n22207), .B(n21816), .Z(n22206) );
  XNOR U22116 ( .A(p_input[1057]), .B(n22208), .Z(n21816) );
  AND U22117 ( .A(n715), .B(n22209), .Z(n22208) );
  XNOR U22118 ( .A(p_input[1073]), .B(n22210), .Z(n22209) );
  IV U22119 ( .A(p_input[1057]), .Z(n22210) );
  XNOR U22120 ( .A(n21813), .B(n22203), .Z(n22205) );
  XNOR U22121 ( .A(p_input[1025]), .B(n22211), .Z(n21813) );
  AND U22122 ( .A(n712), .B(n22212), .Z(n22211) );
  XOR U22123 ( .A(p_input[1041]), .B(p_input[1025]), .Z(n22212) );
  IV U22124 ( .A(n22207), .Z(n22203) );
  AND U22125 ( .A(n22078), .B(n22081), .Z(n22207) );
  XOR U22126 ( .A(p_input[1056]), .B(n22213), .Z(n22081) );
  AND U22127 ( .A(n715), .B(n22214), .Z(n22213) );
  XOR U22128 ( .A(p_input[1072]), .B(p_input[1056]), .Z(n22214) );
  XOR U22129 ( .A(n22215), .B(n22216), .Z(n715) );
  AND U22130 ( .A(n22217), .B(n22218), .Z(n22216) );
  XNOR U22131 ( .A(p_input[1087]), .B(n22215), .Z(n22218) );
  XOR U22132 ( .A(n22215), .B(p_input[1071]), .Z(n22217) );
  XOR U22133 ( .A(n22219), .B(n22220), .Z(n22215) );
  AND U22134 ( .A(n22221), .B(n22222), .Z(n22220) );
  XNOR U22135 ( .A(p_input[1086]), .B(n22219), .Z(n22222) );
  XOR U22136 ( .A(n22219), .B(p_input[1070]), .Z(n22221) );
  XOR U22137 ( .A(n22223), .B(n22224), .Z(n22219) );
  AND U22138 ( .A(n22225), .B(n22226), .Z(n22224) );
  XNOR U22139 ( .A(p_input[1085]), .B(n22223), .Z(n22226) );
  XOR U22140 ( .A(n22223), .B(p_input[1069]), .Z(n22225) );
  XOR U22141 ( .A(n22227), .B(n22228), .Z(n22223) );
  AND U22142 ( .A(n22229), .B(n22230), .Z(n22228) );
  XNOR U22143 ( .A(p_input[1084]), .B(n22227), .Z(n22230) );
  XOR U22144 ( .A(n22227), .B(p_input[1068]), .Z(n22229) );
  XOR U22145 ( .A(n22231), .B(n22232), .Z(n22227) );
  AND U22146 ( .A(n22233), .B(n22234), .Z(n22232) );
  XNOR U22147 ( .A(p_input[1083]), .B(n22231), .Z(n22234) );
  XOR U22148 ( .A(n22231), .B(p_input[1067]), .Z(n22233) );
  XOR U22149 ( .A(n22235), .B(n22236), .Z(n22231) );
  AND U22150 ( .A(n22237), .B(n22238), .Z(n22236) );
  XNOR U22151 ( .A(p_input[1082]), .B(n22235), .Z(n22238) );
  XOR U22152 ( .A(n22235), .B(p_input[1066]), .Z(n22237) );
  XOR U22153 ( .A(n22239), .B(n22240), .Z(n22235) );
  AND U22154 ( .A(n22241), .B(n22242), .Z(n22240) );
  XNOR U22155 ( .A(p_input[1081]), .B(n22239), .Z(n22242) );
  XOR U22156 ( .A(n22239), .B(p_input[1065]), .Z(n22241) );
  XOR U22157 ( .A(n22243), .B(n22244), .Z(n22239) );
  AND U22158 ( .A(n22245), .B(n22246), .Z(n22244) );
  XNOR U22159 ( .A(p_input[1080]), .B(n22243), .Z(n22246) );
  XOR U22160 ( .A(n22243), .B(p_input[1064]), .Z(n22245) );
  XOR U22161 ( .A(n22247), .B(n22248), .Z(n22243) );
  AND U22162 ( .A(n22249), .B(n22250), .Z(n22248) );
  XNOR U22163 ( .A(p_input[1079]), .B(n22247), .Z(n22250) );
  XOR U22164 ( .A(n22247), .B(p_input[1063]), .Z(n22249) );
  XOR U22165 ( .A(n22251), .B(n22252), .Z(n22247) );
  AND U22166 ( .A(n22253), .B(n22254), .Z(n22252) );
  XNOR U22167 ( .A(p_input[1078]), .B(n22251), .Z(n22254) );
  XOR U22168 ( .A(n22251), .B(p_input[1062]), .Z(n22253) );
  XOR U22169 ( .A(n22255), .B(n22256), .Z(n22251) );
  AND U22170 ( .A(n22257), .B(n22258), .Z(n22256) );
  XNOR U22171 ( .A(p_input[1077]), .B(n22255), .Z(n22258) );
  XOR U22172 ( .A(n22255), .B(p_input[1061]), .Z(n22257) );
  XOR U22173 ( .A(n22259), .B(n22260), .Z(n22255) );
  AND U22174 ( .A(n22261), .B(n22262), .Z(n22260) );
  XNOR U22175 ( .A(p_input[1076]), .B(n22259), .Z(n22262) );
  XOR U22176 ( .A(n22259), .B(p_input[1060]), .Z(n22261) );
  XOR U22177 ( .A(n22263), .B(n22264), .Z(n22259) );
  AND U22178 ( .A(n22265), .B(n22266), .Z(n22264) );
  XNOR U22179 ( .A(p_input[1075]), .B(n22263), .Z(n22266) );
  XOR U22180 ( .A(n22263), .B(p_input[1059]), .Z(n22265) );
  XOR U22181 ( .A(n22267), .B(n22268), .Z(n22263) );
  AND U22182 ( .A(n22269), .B(n22270), .Z(n22268) );
  XNOR U22183 ( .A(p_input[1074]), .B(n22267), .Z(n22270) );
  XOR U22184 ( .A(n22267), .B(p_input[1058]), .Z(n22269) );
  XNOR U22185 ( .A(n22271), .B(n22272), .Z(n22267) );
  AND U22186 ( .A(n22273), .B(n22274), .Z(n22272) );
  XOR U22187 ( .A(p_input[1073]), .B(n22271), .Z(n22274) );
  XNOR U22188 ( .A(p_input[1057]), .B(n22271), .Z(n22273) );
  AND U22189 ( .A(p_input[1072]), .B(n22275), .Z(n22271) );
  IV U22190 ( .A(p_input[1056]), .Z(n22275) );
  XNOR U22191 ( .A(p_input[1024]), .B(n22276), .Z(n22078) );
  AND U22192 ( .A(n712), .B(n22277), .Z(n22276) );
  XOR U22193 ( .A(p_input[1040]), .B(p_input[1024]), .Z(n22277) );
  XOR U22194 ( .A(n22278), .B(n22279), .Z(n712) );
  AND U22195 ( .A(n22280), .B(n22281), .Z(n22279) );
  XNOR U22196 ( .A(p_input[1055]), .B(n22278), .Z(n22281) );
  XOR U22197 ( .A(n22278), .B(p_input[1039]), .Z(n22280) );
  XOR U22198 ( .A(n22282), .B(n22283), .Z(n22278) );
  AND U22199 ( .A(n22284), .B(n22285), .Z(n22283) );
  XNOR U22200 ( .A(p_input[1054]), .B(n22282), .Z(n22285) );
  XNOR U22201 ( .A(n22282), .B(n22092), .Z(n22284) );
  IV U22202 ( .A(p_input[1038]), .Z(n22092) );
  XOR U22203 ( .A(n22286), .B(n22287), .Z(n22282) );
  AND U22204 ( .A(n22288), .B(n22289), .Z(n22287) );
  XNOR U22205 ( .A(p_input[1053]), .B(n22286), .Z(n22289) );
  XNOR U22206 ( .A(n22286), .B(n22101), .Z(n22288) );
  IV U22207 ( .A(p_input[1037]), .Z(n22101) );
  XOR U22208 ( .A(n22290), .B(n22291), .Z(n22286) );
  AND U22209 ( .A(n22292), .B(n22293), .Z(n22291) );
  XNOR U22210 ( .A(p_input[1052]), .B(n22290), .Z(n22293) );
  XNOR U22211 ( .A(n22290), .B(n22110), .Z(n22292) );
  IV U22212 ( .A(p_input[1036]), .Z(n22110) );
  XOR U22213 ( .A(n22294), .B(n22295), .Z(n22290) );
  AND U22214 ( .A(n22296), .B(n22297), .Z(n22295) );
  XNOR U22215 ( .A(p_input[1051]), .B(n22294), .Z(n22297) );
  XNOR U22216 ( .A(n22294), .B(n22119), .Z(n22296) );
  IV U22217 ( .A(p_input[1035]), .Z(n22119) );
  XOR U22218 ( .A(n22298), .B(n22299), .Z(n22294) );
  AND U22219 ( .A(n22300), .B(n22301), .Z(n22299) );
  XNOR U22220 ( .A(p_input[1050]), .B(n22298), .Z(n22301) );
  XNOR U22221 ( .A(n22298), .B(n22128), .Z(n22300) );
  IV U22222 ( .A(p_input[1034]), .Z(n22128) );
  XOR U22223 ( .A(n22302), .B(n22303), .Z(n22298) );
  AND U22224 ( .A(n22304), .B(n22305), .Z(n22303) );
  XNOR U22225 ( .A(p_input[1049]), .B(n22302), .Z(n22305) );
  XNOR U22226 ( .A(n22302), .B(n22137), .Z(n22304) );
  IV U22227 ( .A(p_input[1033]), .Z(n22137) );
  XOR U22228 ( .A(n22306), .B(n22307), .Z(n22302) );
  AND U22229 ( .A(n22308), .B(n22309), .Z(n22307) );
  XNOR U22230 ( .A(p_input[1048]), .B(n22306), .Z(n22309) );
  XNOR U22231 ( .A(n22306), .B(n22146), .Z(n22308) );
  IV U22232 ( .A(p_input[1032]), .Z(n22146) );
  XOR U22233 ( .A(n22310), .B(n22311), .Z(n22306) );
  AND U22234 ( .A(n22312), .B(n22313), .Z(n22311) );
  XNOR U22235 ( .A(p_input[1047]), .B(n22310), .Z(n22313) );
  XNOR U22236 ( .A(n22310), .B(n22155), .Z(n22312) );
  IV U22237 ( .A(p_input[1031]), .Z(n22155) );
  XOR U22238 ( .A(n22314), .B(n22315), .Z(n22310) );
  AND U22239 ( .A(n22316), .B(n22317), .Z(n22315) );
  XNOR U22240 ( .A(p_input[1046]), .B(n22314), .Z(n22317) );
  XNOR U22241 ( .A(n22314), .B(n22164), .Z(n22316) );
  IV U22242 ( .A(p_input[1030]), .Z(n22164) );
  XOR U22243 ( .A(n22318), .B(n22319), .Z(n22314) );
  AND U22244 ( .A(n22320), .B(n22321), .Z(n22319) );
  XNOR U22245 ( .A(p_input[1045]), .B(n22318), .Z(n22321) );
  XNOR U22246 ( .A(n22318), .B(n22173), .Z(n22320) );
  IV U22247 ( .A(p_input[1029]), .Z(n22173) );
  XOR U22248 ( .A(n22322), .B(n22323), .Z(n22318) );
  AND U22249 ( .A(n22324), .B(n22325), .Z(n22323) );
  XNOR U22250 ( .A(p_input[1044]), .B(n22322), .Z(n22325) );
  XNOR U22251 ( .A(n22322), .B(n22182), .Z(n22324) );
  IV U22252 ( .A(p_input[1028]), .Z(n22182) );
  XOR U22253 ( .A(n22326), .B(n22327), .Z(n22322) );
  AND U22254 ( .A(n22328), .B(n22329), .Z(n22327) );
  XNOR U22255 ( .A(p_input[1043]), .B(n22326), .Z(n22329) );
  XNOR U22256 ( .A(n22326), .B(n22191), .Z(n22328) );
  IV U22257 ( .A(p_input[1027]), .Z(n22191) );
  XOR U22258 ( .A(n22330), .B(n22331), .Z(n22326) );
  AND U22259 ( .A(n22332), .B(n22333), .Z(n22331) );
  XNOR U22260 ( .A(p_input[1042]), .B(n22330), .Z(n22333) );
  XNOR U22261 ( .A(n22330), .B(n22200), .Z(n22332) );
  IV U22262 ( .A(p_input[1026]), .Z(n22200) );
  XNOR U22263 ( .A(n22334), .B(n22335), .Z(n22330) );
  AND U22264 ( .A(n22336), .B(n22337), .Z(n22335) );
  XOR U22265 ( .A(p_input[1041]), .B(n22334), .Z(n22337) );
  XNOR U22266 ( .A(p_input[1025]), .B(n22334), .Z(n22336) );
  AND U22267 ( .A(p_input[1040]), .B(n22338), .Z(n22334) );
  IV U22268 ( .A(p_input[1024]), .Z(n22338) );
  XOR U22269 ( .A(n22339), .B(n22340), .Z(n15247) );
  AND U22270 ( .A(n1048), .B(n22341), .Z(n22340) );
  XNOR U22271 ( .A(n22342), .B(n22339), .Z(n22341) );
  XOR U22272 ( .A(n22343), .B(n22344), .Z(n1048) );
  AND U22273 ( .A(n22345), .B(n22346), .Z(n22344) );
  XOR U22274 ( .A(n22343), .B(n15262), .Z(n22346) );
  XOR U22275 ( .A(n22347), .B(n22348), .Z(n15262) );
  AND U22276 ( .A(n1023), .B(n22349), .Z(n22348) );
  XOR U22277 ( .A(n22350), .B(n22347), .Z(n22349) );
  XNOR U22278 ( .A(n15259), .B(n22343), .Z(n22345) );
  XOR U22279 ( .A(n22351), .B(n22352), .Z(n15259) );
  AND U22280 ( .A(n1020), .B(n22353), .Z(n22352) );
  XOR U22281 ( .A(n22354), .B(n22351), .Z(n22353) );
  XOR U22282 ( .A(n22355), .B(n22356), .Z(n22343) );
  AND U22283 ( .A(n22357), .B(n22358), .Z(n22356) );
  XOR U22284 ( .A(n22355), .B(n15274), .Z(n22358) );
  XOR U22285 ( .A(n22359), .B(n22360), .Z(n15274) );
  AND U22286 ( .A(n1023), .B(n22361), .Z(n22360) );
  XOR U22287 ( .A(n22362), .B(n22359), .Z(n22361) );
  XNOR U22288 ( .A(n15271), .B(n22355), .Z(n22357) );
  XOR U22289 ( .A(n22363), .B(n22364), .Z(n15271) );
  AND U22290 ( .A(n1020), .B(n22365), .Z(n22364) );
  XOR U22291 ( .A(n22366), .B(n22363), .Z(n22365) );
  XOR U22292 ( .A(n22367), .B(n22368), .Z(n22355) );
  AND U22293 ( .A(n22369), .B(n22370), .Z(n22368) );
  XOR U22294 ( .A(n22367), .B(n15286), .Z(n22370) );
  XOR U22295 ( .A(n22371), .B(n22372), .Z(n15286) );
  AND U22296 ( .A(n1023), .B(n22373), .Z(n22372) );
  XOR U22297 ( .A(n22374), .B(n22371), .Z(n22373) );
  XNOR U22298 ( .A(n15283), .B(n22367), .Z(n22369) );
  XOR U22299 ( .A(n22375), .B(n22376), .Z(n15283) );
  AND U22300 ( .A(n1020), .B(n22377), .Z(n22376) );
  XOR U22301 ( .A(n22378), .B(n22375), .Z(n22377) );
  XOR U22302 ( .A(n22379), .B(n22380), .Z(n22367) );
  AND U22303 ( .A(n22381), .B(n22382), .Z(n22380) );
  XOR U22304 ( .A(n22379), .B(n15298), .Z(n22382) );
  XOR U22305 ( .A(n22383), .B(n22384), .Z(n15298) );
  AND U22306 ( .A(n1023), .B(n22385), .Z(n22384) );
  XOR U22307 ( .A(n22386), .B(n22383), .Z(n22385) );
  XNOR U22308 ( .A(n15295), .B(n22379), .Z(n22381) );
  XOR U22309 ( .A(n22387), .B(n22388), .Z(n15295) );
  AND U22310 ( .A(n1020), .B(n22389), .Z(n22388) );
  XOR U22311 ( .A(n22390), .B(n22387), .Z(n22389) );
  XOR U22312 ( .A(n22391), .B(n22392), .Z(n22379) );
  AND U22313 ( .A(n22393), .B(n22394), .Z(n22392) );
  XOR U22314 ( .A(n22391), .B(n15310), .Z(n22394) );
  XOR U22315 ( .A(n22395), .B(n22396), .Z(n15310) );
  AND U22316 ( .A(n1023), .B(n22397), .Z(n22396) );
  XOR U22317 ( .A(n22398), .B(n22395), .Z(n22397) );
  XNOR U22318 ( .A(n15307), .B(n22391), .Z(n22393) );
  XOR U22319 ( .A(n22399), .B(n22400), .Z(n15307) );
  AND U22320 ( .A(n1020), .B(n22401), .Z(n22400) );
  XOR U22321 ( .A(n22402), .B(n22399), .Z(n22401) );
  XOR U22322 ( .A(n22403), .B(n22404), .Z(n22391) );
  AND U22323 ( .A(n22405), .B(n22406), .Z(n22404) );
  XOR U22324 ( .A(n22403), .B(n15322), .Z(n22406) );
  XOR U22325 ( .A(n22407), .B(n22408), .Z(n15322) );
  AND U22326 ( .A(n1023), .B(n22409), .Z(n22408) );
  XOR U22327 ( .A(n22410), .B(n22407), .Z(n22409) );
  XNOR U22328 ( .A(n15319), .B(n22403), .Z(n22405) );
  XOR U22329 ( .A(n22411), .B(n22412), .Z(n15319) );
  AND U22330 ( .A(n1020), .B(n22413), .Z(n22412) );
  XOR U22331 ( .A(n22414), .B(n22411), .Z(n22413) );
  XOR U22332 ( .A(n22415), .B(n22416), .Z(n22403) );
  AND U22333 ( .A(n22417), .B(n22418), .Z(n22416) );
  XOR U22334 ( .A(n22415), .B(n15334), .Z(n22418) );
  XOR U22335 ( .A(n22419), .B(n22420), .Z(n15334) );
  AND U22336 ( .A(n1023), .B(n22421), .Z(n22420) );
  XOR U22337 ( .A(n22422), .B(n22419), .Z(n22421) );
  XNOR U22338 ( .A(n15331), .B(n22415), .Z(n22417) );
  XOR U22339 ( .A(n22423), .B(n22424), .Z(n15331) );
  AND U22340 ( .A(n1020), .B(n22425), .Z(n22424) );
  XOR U22341 ( .A(n22426), .B(n22423), .Z(n22425) );
  XOR U22342 ( .A(n22427), .B(n22428), .Z(n22415) );
  AND U22343 ( .A(n22429), .B(n22430), .Z(n22428) );
  XOR U22344 ( .A(n22427), .B(n15346), .Z(n22430) );
  XOR U22345 ( .A(n22431), .B(n22432), .Z(n15346) );
  AND U22346 ( .A(n1023), .B(n22433), .Z(n22432) );
  XOR U22347 ( .A(n22434), .B(n22431), .Z(n22433) );
  XNOR U22348 ( .A(n15343), .B(n22427), .Z(n22429) );
  XOR U22349 ( .A(n22435), .B(n22436), .Z(n15343) );
  AND U22350 ( .A(n1020), .B(n22437), .Z(n22436) );
  XOR U22351 ( .A(n22438), .B(n22435), .Z(n22437) );
  XOR U22352 ( .A(n22439), .B(n22440), .Z(n22427) );
  AND U22353 ( .A(n22441), .B(n22442), .Z(n22440) );
  XOR U22354 ( .A(n22439), .B(n15358), .Z(n22442) );
  XOR U22355 ( .A(n22443), .B(n22444), .Z(n15358) );
  AND U22356 ( .A(n1023), .B(n22445), .Z(n22444) );
  XOR U22357 ( .A(n22446), .B(n22443), .Z(n22445) );
  XNOR U22358 ( .A(n15355), .B(n22439), .Z(n22441) );
  XOR U22359 ( .A(n22447), .B(n22448), .Z(n15355) );
  AND U22360 ( .A(n1020), .B(n22449), .Z(n22448) );
  XOR U22361 ( .A(n22450), .B(n22447), .Z(n22449) );
  XOR U22362 ( .A(n22451), .B(n22452), .Z(n22439) );
  AND U22363 ( .A(n22453), .B(n22454), .Z(n22452) );
  XOR U22364 ( .A(n22451), .B(n15370), .Z(n22454) );
  XOR U22365 ( .A(n22455), .B(n22456), .Z(n15370) );
  AND U22366 ( .A(n1023), .B(n22457), .Z(n22456) );
  XOR U22367 ( .A(n22458), .B(n22455), .Z(n22457) );
  XNOR U22368 ( .A(n15367), .B(n22451), .Z(n22453) );
  XOR U22369 ( .A(n22459), .B(n22460), .Z(n15367) );
  AND U22370 ( .A(n1020), .B(n22461), .Z(n22460) );
  XOR U22371 ( .A(n22462), .B(n22459), .Z(n22461) );
  XOR U22372 ( .A(n22463), .B(n22464), .Z(n22451) );
  AND U22373 ( .A(n22465), .B(n22466), .Z(n22464) );
  XOR U22374 ( .A(n22463), .B(n15382), .Z(n22466) );
  XOR U22375 ( .A(n22467), .B(n22468), .Z(n15382) );
  AND U22376 ( .A(n1023), .B(n22469), .Z(n22468) );
  XOR U22377 ( .A(n22470), .B(n22467), .Z(n22469) );
  XNOR U22378 ( .A(n15379), .B(n22463), .Z(n22465) );
  XOR U22379 ( .A(n22471), .B(n22472), .Z(n15379) );
  AND U22380 ( .A(n1020), .B(n22473), .Z(n22472) );
  XOR U22381 ( .A(n22474), .B(n22471), .Z(n22473) );
  XOR U22382 ( .A(n22475), .B(n22476), .Z(n22463) );
  AND U22383 ( .A(n22477), .B(n22478), .Z(n22476) );
  XOR U22384 ( .A(n22475), .B(n15394), .Z(n22478) );
  XOR U22385 ( .A(n22479), .B(n22480), .Z(n15394) );
  AND U22386 ( .A(n1023), .B(n22481), .Z(n22480) );
  XOR U22387 ( .A(n22482), .B(n22479), .Z(n22481) );
  XNOR U22388 ( .A(n15391), .B(n22475), .Z(n22477) );
  XOR U22389 ( .A(n22483), .B(n22484), .Z(n15391) );
  AND U22390 ( .A(n1020), .B(n22485), .Z(n22484) );
  XOR U22391 ( .A(n22486), .B(n22483), .Z(n22485) );
  XOR U22392 ( .A(n22487), .B(n22488), .Z(n22475) );
  AND U22393 ( .A(n22489), .B(n22490), .Z(n22488) );
  XOR U22394 ( .A(n22487), .B(n15406), .Z(n22490) );
  XOR U22395 ( .A(n22491), .B(n22492), .Z(n15406) );
  AND U22396 ( .A(n1023), .B(n22493), .Z(n22492) );
  XOR U22397 ( .A(n22494), .B(n22491), .Z(n22493) );
  XNOR U22398 ( .A(n15403), .B(n22487), .Z(n22489) );
  XOR U22399 ( .A(n22495), .B(n22496), .Z(n15403) );
  AND U22400 ( .A(n1020), .B(n22497), .Z(n22496) );
  XOR U22401 ( .A(n22498), .B(n22495), .Z(n22497) );
  XOR U22402 ( .A(n22499), .B(n22500), .Z(n22487) );
  AND U22403 ( .A(n22501), .B(n22502), .Z(n22500) );
  XOR U22404 ( .A(n22499), .B(n15418), .Z(n22502) );
  XOR U22405 ( .A(n22503), .B(n22504), .Z(n15418) );
  AND U22406 ( .A(n1023), .B(n22505), .Z(n22504) );
  XOR U22407 ( .A(n22506), .B(n22503), .Z(n22505) );
  XNOR U22408 ( .A(n15415), .B(n22499), .Z(n22501) );
  XOR U22409 ( .A(n22507), .B(n22508), .Z(n15415) );
  AND U22410 ( .A(n1020), .B(n22509), .Z(n22508) );
  XOR U22411 ( .A(n22510), .B(n22507), .Z(n22509) );
  XOR U22412 ( .A(n22511), .B(n22512), .Z(n22499) );
  AND U22413 ( .A(n22513), .B(n22514), .Z(n22512) );
  XNOR U22414 ( .A(n22515), .B(n15431), .Z(n22514) );
  XOR U22415 ( .A(n22516), .B(n22517), .Z(n15431) );
  AND U22416 ( .A(n1023), .B(n22518), .Z(n22517) );
  XOR U22417 ( .A(n22516), .B(n22519), .Z(n22518) );
  XNOR U22418 ( .A(n15428), .B(n22511), .Z(n22513) );
  XOR U22419 ( .A(n22520), .B(n22521), .Z(n15428) );
  AND U22420 ( .A(n1020), .B(n22522), .Z(n22521) );
  XOR U22421 ( .A(n22520), .B(n22523), .Z(n22522) );
  IV U22422 ( .A(n22515), .Z(n22511) );
  AND U22423 ( .A(n22339), .B(n22342), .Z(n22515) );
  XNOR U22424 ( .A(n22524), .B(n22525), .Z(n22342) );
  AND U22425 ( .A(n1023), .B(n22526), .Z(n22525) );
  XNOR U22426 ( .A(n22527), .B(n22524), .Z(n22526) );
  XOR U22427 ( .A(n22528), .B(n22529), .Z(n1023) );
  AND U22428 ( .A(n22530), .B(n22531), .Z(n22529) );
  XOR U22429 ( .A(n22528), .B(n22350), .Z(n22531) );
  XNOR U22430 ( .A(n22532), .B(n22533), .Z(n22350) );
  AND U22431 ( .A(n22534), .B(n959), .Z(n22533) );
  AND U22432 ( .A(n22532), .B(n22535), .Z(n22534) );
  XNOR U22433 ( .A(n22347), .B(n22528), .Z(n22530) );
  XOR U22434 ( .A(n22536), .B(n22537), .Z(n22347) );
  AND U22435 ( .A(n22538), .B(n957), .Z(n22537) );
  NOR U22436 ( .A(n22536), .B(n22539), .Z(n22538) );
  XOR U22437 ( .A(n22540), .B(n22541), .Z(n22528) );
  AND U22438 ( .A(n22542), .B(n22543), .Z(n22541) );
  XOR U22439 ( .A(n22540), .B(n22362), .Z(n22543) );
  XOR U22440 ( .A(n22544), .B(n22545), .Z(n22362) );
  AND U22441 ( .A(n959), .B(n22546), .Z(n22545) );
  XOR U22442 ( .A(n22547), .B(n22544), .Z(n22546) );
  XNOR U22443 ( .A(n22359), .B(n22540), .Z(n22542) );
  XOR U22444 ( .A(n22548), .B(n22549), .Z(n22359) );
  AND U22445 ( .A(n957), .B(n22550), .Z(n22549) );
  XOR U22446 ( .A(n22551), .B(n22548), .Z(n22550) );
  XOR U22447 ( .A(n22552), .B(n22553), .Z(n22540) );
  AND U22448 ( .A(n22554), .B(n22555), .Z(n22553) );
  XOR U22449 ( .A(n22552), .B(n22374), .Z(n22555) );
  XOR U22450 ( .A(n22556), .B(n22557), .Z(n22374) );
  AND U22451 ( .A(n959), .B(n22558), .Z(n22557) );
  XOR U22452 ( .A(n22559), .B(n22556), .Z(n22558) );
  XNOR U22453 ( .A(n22371), .B(n22552), .Z(n22554) );
  XOR U22454 ( .A(n22560), .B(n22561), .Z(n22371) );
  AND U22455 ( .A(n957), .B(n22562), .Z(n22561) );
  XOR U22456 ( .A(n22563), .B(n22560), .Z(n22562) );
  XOR U22457 ( .A(n22564), .B(n22565), .Z(n22552) );
  AND U22458 ( .A(n22566), .B(n22567), .Z(n22565) );
  XOR U22459 ( .A(n22564), .B(n22386), .Z(n22567) );
  XOR U22460 ( .A(n22568), .B(n22569), .Z(n22386) );
  AND U22461 ( .A(n959), .B(n22570), .Z(n22569) );
  XOR U22462 ( .A(n22571), .B(n22568), .Z(n22570) );
  XNOR U22463 ( .A(n22383), .B(n22564), .Z(n22566) );
  XOR U22464 ( .A(n22572), .B(n22573), .Z(n22383) );
  AND U22465 ( .A(n957), .B(n22574), .Z(n22573) );
  XOR U22466 ( .A(n22575), .B(n22572), .Z(n22574) );
  XOR U22467 ( .A(n22576), .B(n22577), .Z(n22564) );
  AND U22468 ( .A(n22578), .B(n22579), .Z(n22577) );
  XOR U22469 ( .A(n22576), .B(n22398), .Z(n22579) );
  XOR U22470 ( .A(n22580), .B(n22581), .Z(n22398) );
  AND U22471 ( .A(n959), .B(n22582), .Z(n22581) );
  XOR U22472 ( .A(n22583), .B(n22580), .Z(n22582) );
  XNOR U22473 ( .A(n22395), .B(n22576), .Z(n22578) );
  XOR U22474 ( .A(n22584), .B(n22585), .Z(n22395) );
  AND U22475 ( .A(n957), .B(n22586), .Z(n22585) );
  XOR U22476 ( .A(n22587), .B(n22584), .Z(n22586) );
  XOR U22477 ( .A(n22588), .B(n22589), .Z(n22576) );
  AND U22478 ( .A(n22590), .B(n22591), .Z(n22589) );
  XOR U22479 ( .A(n22588), .B(n22410), .Z(n22591) );
  XOR U22480 ( .A(n22592), .B(n22593), .Z(n22410) );
  AND U22481 ( .A(n959), .B(n22594), .Z(n22593) );
  XOR U22482 ( .A(n22595), .B(n22592), .Z(n22594) );
  XNOR U22483 ( .A(n22407), .B(n22588), .Z(n22590) );
  XOR U22484 ( .A(n22596), .B(n22597), .Z(n22407) );
  AND U22485 ( .A(n957), .B(n22598), .Z(n22597) );
  XOR U22486 ( .A(n22599), .B(n22596), .Z(n22598) );
  XOR U22487 ( .A(n22600), .B(n22601), .Z(n22588) );
  AND U22488 ( .A(n22602), .B(n22603), .Z(n22601) );
  XOR U22489 ( .A(n22600), .B(n22422), .Z(n22603) );
  XOR U22490 ( .A(n22604), .B(n22605), .Z(n22422) );
  AND U22491 ( .A(n959), .B(n22606), .Z(n22605) );
  XOR U22492 ( .A(n22607), .B(n22604), .Z(n22606) );
  XNOR U22493 ( .A(n22419), .B(n22600), .Z(n22602) );
  XOR U22494 ( .A(n22608), .B(n22609), .Z(n22419) );
  AND U22495 ( .A(n957), .B(n22610), .Z(n22609) );
  XOR U22496 ( .A(n22611), .B(n22608), .Z(n22610) );
  XOR U22497 ( .A(n22612), .B(n22613), .Z(n22600) );
  AND U22498 ( .A(n22614), .B(n22615), .Z(n22613) );
  XOR U22499 ( .A(n22612), .B(n22434), .Z(n22615) );
  XOR U22500 ( .A(n22616), .B(n22617), .Z(n22434) );
  AND U22501 ( .A(n959), .B(n22618), .Z(n22617) );
  XOR U22502 ( .A(n22619), .B(n22616), .Z(n22618) );
  XNOR U22503 ( .A(n22431), .B(n22612), .Z(n22614) );
  XOR U22504 ( .A(n22620), .B(n22621), .Z(n22431) );
  AND U22505 ( .A(n957), .B(n22622), .Z(n22621) );
  XOR U22506 ( .A(n22623), .B(n22620), .Z(n22622) );
  XOR U22507 ( .A(n22624), .B(n22625), .Z(n22612) );
  AND U22508 ( .A(n22626), .B(n22627), .Z(n22625) );
  XOR U22509 ( .A(n22624), .B(n22446), .Z(n22627) );
  XOR U22510 ( .A(n22628), .B(n22629), .Z(n22446) );
  AND U22511 ( .A(n959), .B(n22630), .Z(n22629) );
  XOR U22512 ( .A(n22631), .B(n22628), .Z(n22630) );
  XNOR U22513 ( .A(n22443), .B(n22624), .Z(n22626) );
  XOR U22514 ( .A(n22632), .B(n22633), .Z(n22443) );
  AND U22515 ( .A(n957), .B(n22634), .Z(n22633) );
  XOR U22516 ( .A(n22635), .B(n22632), .Z(n22634) );
  XOR U22517 ( .A(n22636), .B(n22637), .Z(n22624) );
  AND U22518 ( .A(n22638), .B(n22639), .Z(n22637) );
  XOR U22519 ( .A(n22636), .B(n22458), .Z(n22639) );
  XOR U22520 ( .A(n22640), .B(n22641), .Z(n22458) );
  AND U22521 ( .A(n959), .B(n22642), .Z(n22641) );
  XOR U22522 ( .A(n22643), .B(n22640), .Z(n22642) );
  XNOR U22523 ( .A(n22455), .B(n22636), .Z(n22638) );
  XOR U22524 ( .A(n22644), .B(n22645), .Z(n22455) );
  AND U22525 ( .A(n957), .B(n22646), .Z(n22645) );
  XOR U22526 ( .A(n22647), .B(n22644), .Z(n22646) );
  XOR U22527 ( .A(n22648), .B(n22649), .Z(n22636) );
  AND U22528 ( .A(n22650), .B(n22651), .Z(n22649) );
  XOR U22529 ( .A(n22648), .B(n22470), .Z(n22651) );
  XOR U22530 ( .A(n22652), .B(n22653), .Z(n22470) );
  AND U22531 ( .A(n959), .B(n22654), .Z(n22653) );
  XOR U22532 ( .A(n22655), .B(n22652), .Z(n22654) );
  XNOR U22533 ( .A(n22467), .B(n22648), .Z(n22650) );
  XOR U22534 ( .A(n22656), .B(n22657), .Z(n22467) );
  AND U22535 ( .A(n957), .B(n22658), .Z(n22657) );
  XOR U22536 ( .A(n22659), .B(n22656), .Z(n22658) );
  XOR U22537 ( .A(n22660), .B(n22661), .Z(n22648) );
  AND U22538 ( .A(n22662), .B(n22663), .Z(n22661) );
  XOR U22539 ( .A(n22660), .B(n22482), .Z(n22663) );
  XOR U22540 ( .A(n22664), .B(n22665), .Z(n22482) );
  AND U22541 ( .A(n959), .B(n22666), .Z(n22665) );
  XOR U22542 ( .A(n22667), .B(n22664), .Z(n22666) );
  XNOR U22543 ( .A(n22479), .B(n22660), .Z(n22662) );
  XOR U22544 ( .A(n22668), .B(n22669), .Z(n22479) );
  AND U22545 ( .A(n957), .B(n22670), .Z(n22669) );
  XOR U22546 ( .A(n22671), .B(n22668), .Z(n22670) );
  XOR U22547 ( .A(n22672), .B(n22673), .Z(n22660) );
  AND U22548 ( .A(n22674), .B(n22675), .Z(n22673) );
  XOR U22549 ( .A(n22672), .B(n22494), .Z(n22675) );
  XOR U22550 ( .A(n22676), .B(n22677), .Z(n22494) );
  AND U22551 ( .A(n959), .B(n22678), .Z(n22677) );
  XOR U22552 ( .A(n22679), .B(n22676), .Z(n22678) );
  XNOR U22553 ( .A(n22491), .B(n22672), .Z(n22674) );
  XOR U22554 ( .A(n22680), .B(n22681), .Z(n22491) );
  AND U22555 ( .A(n957), .B(n22682), .Z(n22681) );
  XOR U22556 ( .A(n22683), .B(n22680), .Z(n22682) );
  XOR U22557 ( .A(n22684), .B(n22685), .Z(n22672) );
  AND U22558 ( .A(n22686), .B(n22687), .Z(n22685) );
  XOR U22559 ( .A(n22684), .B(n22506), .Z(n22687) );
  XOR U22560 ( .A(n22688), .B(n22689), .Z(n22506) );
  AND U22561 ( .A(n959), .B(n22690), .Z(n22689) );
  XOR U22562 ( .A(n22691), .B(n22688), .Z(n22690) );
  XNOR U22563 ( .A(n22503), .B(n22684), .Z(n22686) );
  XOR U22564 ( .A(n22692), .B(n22693), .Z(n22503) );
  AND U22565 ( .A(n957), .B(n22694), .Z(n22693) );
  XOR U22566 ( .A(n22695), .B(n22692), .Z(n22694) );
  XOR U22567 ( .A(n22696), .B(n22697), .Z(n22684) );
  AND U22568 ( .A(n22698), .B(n22699), .Z(n22697) );
  XNOR U22569 ( .A(n22700), .B(n22519), .Z(n22699) );
  XOR U22570 ( .A(n22701), .B(n22702), .Z(n22519) );
  AND U22571 ( .A(n959), .B(n22703), .Z(n22702) );
  XOR U22572 ( .A(n22701), .B(n22704), .Z(n22703) );
  XNOR U22573 ( .A(n22516), .B(n22696), .Z(n22698) );
  XOR U22574 ( .A(n22705), .B(n22706), .Z(n22516) );
  AND U22575 ( .A(n957), .B(n22707), .Z(n22706) );
  XOR U22576 ( .A(n22705), .B(n22708), .Z(n22707) );
  IV U22577 ( .A(n22700), .Z(n22696) );
  AND U22578 ( .A(n22524), .B(n22527), .Z(n22700) );
  XNOR U22579 ( .A(n22709), .B(n22710), .Z(n22527) );
  AND U22580 ( .A(n959), .B(n22711), .Z(n22710) );
  XNOR U22581 ( .A(n22712), .B(n22709), .Z(n22711) );
  XOR U22582 ( .A(n22713), .B(n22714), .Z(n959) );
  AND U22583 ( .A(n22715), .B(n22716), .Z(n22714) );
  XOR U22584 ( .A(n22535), .B(n22713), .Z(n22716) );
  IV U22585 ( .A(n22717), .Z(n22535) );
  AND U22586 ( .A(n22718), .B(n22719), .Z(n22717) );
  XOR U22587 ( .A(n22713), .B(n22532), .Z(n22715) );
  AND U22588 ( .A(n22720), .B(n22721), .Z(n22532) );
  XOR U22589 ( .A(n22722), .B(n22723), .Z(n22713) );
  AND U22590 ( .A(n22724), .B(n22725), .Z(n22723) );
  XOR U22591 ( .A(n22722), .B(n22547), .Z(n22725) );
  XOR U22592 ( .A(n22726), .B(n22727), .Z(n22547) );
  AND U22593 ( .A(n823), .B(n22728), .Z(n22727) );
  XOR U22594 ( .A(n22729), .B(n22726), .Z(n22728) );
  XNOR U22595 ( .A(n22544), .B(n22722), .Z(n22724) );
  XOR U22596 ( .A(n22730), .B(n22731), .Z(n22544) );
  AND U22597 ( .A(n821), .B(n22732), .Z(n22731) );
  XOR U22598 ( .A(n22733), .B(n22730), .Z(n22732) );
  XOR U22599 ( .A(n22734), .B(n22735), .Z(n22722) );
  AND U22600 ( .A(n22736), .B(n22737), .Z(n22735) );
  XOR U22601 ( .A(n22734), .B(n22559), .Z(n22737) );
  XOR U22602 ( .A(n22738), .B(n22739), .Z(n22559) );
  AND U22603 ( .A(n823), .B(n22740), .Z(n22739) );
  XOR U22604 ( .A(n22741), .B(n22738), .Z(n22740) );
  XNOR U22605 ( .A(n22556), .B(n22734), .Z(n22736) );
  XOR U22606 ( .A(n22742), .B(n22743), .Z(n22556) );
  AND U22607 ( .A(n821), .B(n22744), .Z(n22743) );
  XOR U22608 ( .A(n22745), .B(n22742), .Z(n22744) );
  XOR U22609 ( .A(n22746), .B(n22747), .Z(n22734) );
  AND U22610 ( .A(n22748), .B(n22749), .Z(n22747) );
  XOR U22611 ( .A(n22746), .B(n22571), .Z(n22749) );
  XOR U22612 ( .A(n22750), .B(n22751), .Z(n22571) );
  AND U22613 ( .A(n823), .B(n22752), .Z(n22751) );
  XOR U22614 ( .A(n22753), .B(n22750), .Z(n22752) );
  XNOR U22615 ( .A(n22568), .B(n22746), .Z(n22748) );
  XOR U22616 ( .A(n22754), .B(n22755), .Z(n22568) );
  AND U22617 ( .A(n821), .B(n22756), .Z(n22755) );
  XOR U22618 ( .A(n22757), .B(n22754), .Z(n22756) );
  XOR U22619 ( .A(n22758), .B(n22759), .Z(n22746) );
  AND U22620 ( .A(n22760), .B(n22761), .Z(n22759) );
  XOR U22621 ( .A(n22758), .B(n22583), .Z(n22761) );
  XOR U22622 ( .A(n22762), .B(n22763), .Z(n22583) );
  AND U22623 ( .A(n823), .B(n22764), .Z(n22763) );
  XOR U22624 ( .A(n22765), .B(n22762), .Z(n22764) );
  XNOR U22625 ( .A(n22580), .B(n22758), .Z(n22760) );
  XOR U22626 ( .A(n22766), .B(n22767), .Z(n22580) );
  AND U22627 ( .A(n821), .B(n22768), .Z(n22767) );
  XOR U22628 ( .A(n22769), .B(n22766), .Z(n22768) );
  XOR U22629 ( .A(n22770), .B(n22771), .Z(n22758) );
  AND U22630 ( .A(n22772), .B(n22773), .Z(n22771) );
  XOR U22631 ( .A(n22770), .B(n22595), .Z(n22773) );
  XOR U22632 ( .A(n22774), .B(n22775), .Z(n22595) );
  AND U22633 ( .A(n823), .B(n22776), .Z(n22775) );
  XOR U22634 ( .A(n22777), .B(n22774), .Z(n22776) );
  XNOR U22635 ( .A(n22592), .B(n22770), .Z(n22772) );
  XOR U22636 ( .A(n22778), .B(n22779), .Z(n22592) );
  AND U22637 ( .A(n821), .B(n22780), .Z(n22779) );
  XOR U22638 ( .A(n22781), .B(n22778), .Z(n22780) );
  XOR U22639 ( .A(n22782), .B(n22783), .Z(n22770) );
  AND U22640 ( .A(n22784), .B(n22785), .Z(n22783) );
  XOR U22641 ( .A(n22782), .B(n22607), .Z(n22785) );
  XOR U22642 ( .A(n22786), .B(n22787), .Z(n22607) );
  AND U22643 ( .A(n823), .B(n22788), .Z(n22787) );
  XOR U22644 ( .A(n22789), .B(n22786), .Z(n22788) );
  XNOR U22645 ( .A(n22604), .B(n22782), .Z(n22784) );
  XOR U22646 ( .A(n22790), .B(n22791), .Z(n22604) );
  AND U22647 ( .A(n821), .B(n22792), .Z(n22791) );
  XOR U22648 ( .A(n22793), .B(n22790), .Z(n22792) );
  XOR U22649 ( .A(n22794), .B(n22795), .Z(n22782) );
  AND U22650 ( .A(n22796), .B(n22797), .Z(n22795) );
  XOR U22651 ( .A(n22794), .B(n22619), .Z(n22797) );
  XOR U22652 ( .A(n22798), .B(n22799), .Z(n22619) );
  AND U22653 ( .A(n823), .B(n22800), .Z(n22799) );
  XOR U22654 ( .A(n22801), .B(n22798), .Z(n22800) );
  XNOR U22655 ( .A(n22616), .B(n22794), .Z(n22796) );
  XOR U22656 ( .A(n22802), .B(n22803), .Z(n22616) );
  AND U22657 ( .A(n821), .B(n22804), .Z(n22803) );
  XOR U22658 ( .A(n22805), .B(n22802), .Z(n22804) );
  XOR U22659 ( .A(n22806), .B(n22807), .Z(n22794) );
  AND U22660 ( .A(n22808), .B(n22809), .Z(n22807) );
  XOR U22661 ( .A(n22806), .B(n22631), .Z(n22809) );
  XOR U22662 ( .A(n22810), .B(n22811), .Z(n22631) );
  AND U22663 ( .A(n823), .B(n22812), .Z(n22811) );
  XOR U22664 ( .A(n22813), .B(n22810), .Z(n22812) );
  XNOR U22665 ( .A(n22628), .B(n22806), .Z(n22808) );
  XOR U22666 ( .A(n22814), .B(n22815), .Z(n22628) );
  AND U22667 ( .A(n821), .B(n22816), .Z(n22815) );
  XOR U22668 ( .A(n22817), .B(n22814), .Z(n22816) );
  XOR U22669 ( .A(n22818), .B(n22819), .Z(n22806) );
  AND U22670 ( .A(n22820), .B(n22821), .Z(n22819) );
  XOR U22671 ( .A(n22818), .B(n22643), .Z(n22821) );
  XOR U22672 ( .A(n22822), .B(n22823), .Z(n22643) );
  AND U22673 ( .A(n823), .B(n22824), .Z(n22823) );
  XOR U22674 ( .A(n22825), .B(n22822), .Z(n22824) );
  XNOR U22675 ( .A(n22640), .B(n22818), .Z(n22820) );
  XOR U22676 ( .A(n22826), .B(n22827), .Z(n22640) );
  AND U22677 ( .A(n821), .B(n22828), .Z(n22827) );
  XOR U22678 ( .A(n22829), .B(n22826), .Z(n22828) );
  XOR U22679 ( .A(n22830), .B(n22831), .Z(n22818) );
  AND U22680 ( .A(n22832), .B(n22833), .Z(n22831) );
  XOR U22681 ( .A(n22830), .B(n22655), .Z(n22833) );
  XOR U22682 ( .A(n22834), .B(n22835), .Z(n22655) );
  AND U22683 ( .A(n823), .B(n22836), .Z(n22835) );
  XOR U22684 ( .A(n22837), .B(n22834), .Z(n22836) );
  XNOR U22685 ( .A(n22652), .B(n22830), .Z(n22832) );
  XOR U22686 ( .A(n22838), .B(n22839), .Z(n22652) );
  AND U22687 ( .A(n821), .B(n22840), .Z(n22839) );
  XOR U22688 ( .A(n22841), .B(n22838), .Z(n22840) );
  XOR U22689 ( .A(n22842), .B(n22843), .Z(n22830) );
  AND U22690 ( .A(n22844), .B(n22845), .Z(n22843) );
  XOR U22691 ( .A(n22842), .B(n22667), .Z(n22845) );
  XOR U22692 ( .A(n22846), .B(n22847), .Z(n22667) );
  AND U22693 ( .A(n823), .B(n22848), .Z(n22847) );
  XOR U22694 ( .A(n22849), .B(n22846), .Z(n22848) );
  XNOR U22695 ( .A(n22664), .B(n22842), .Z(n22844) );
  XOR U22696 ( .A(n22850), .B(n22851), .Z(n22664) );
  AND U22697 ( .A(n821), .B(n22852), .Z(n22851) );
  XOR U22698 ( .A(n22853), .B(n22850), .Z(n22852) );
  XOR U22699 ( .A(n22854), .B(n22855), .Z(n22842) );
  AND U22700 ( .A(n22856), .B(n22857), .Z(n22855) );
  XOR U22701 ( .A(n22854), .B(n22679), .Z(n22857) );
  XOR U22702 ( .A(n22858), .B(n22859), .Z(n22679) );
  AND U22703 ( .A(n823), .B(n22860), .Z(n22859) );
  XOR U22704 ( .A(n22861), .B(n22858), .Z(n22860) );
  XNOR U22705 ( .A(n22676), .B(n22854), .Z(n22856) );
  XOR U22706 ( .A(n22862), .B(n22863), .Z(n22676) );
  AND U22707 ( .A(n821), .B(n22864), .Z(n22863) );
  XOR U22708 ( .A(n22865), .B(n22862), .Z(n22864) );
  XOR U22709 ( .A(n22866), .B(n22867), .Z(n22854) );
  AND U22710 ( .A(n22868), .B(n22869), .Z(n22867) );
  XOR U22711 ( .A(n22866), .B(n22691), .Z(n22869) );
  XOR U22712 ( .A(n22870), .B(n22871), .Z(n22691) );
  AND U22713 ( .A(n823), .B(n22872), .Z(n22871) );
  XOR U22714 ( .A(n22873), .B(n22870), .Z(n22872) );
  XNOR U22715 ( .A(n22688), .B(n22866), .Z(n22868) );
  XOR U22716 ( .A(n22874), .B(n22875), .Z(n22688) );
  AND U22717 ( .A(n821), .B(n22876), .Z(n22875) );
  XOR U22718 ( .A(n22877), .B(n22874), .Z(n22876) );
  XOR U22719 ( .A(n22878), .B(n22879), .Z(n22866) );
  AND U22720 ( .A(n22880), .B(n22881), .Z(n22879) );
  XNOR U22721 ( .A(n22882), .B(n22704), .Z(n22881) );
  XOR U22722 ( .A(n22883), .B(n22884), .Z(n22704) );
  AND U22723 ( .A(n823), .B(n22885), .Z(n22884) );
  XOR U22724 ( .A(n22883), .B(n22886), .Z(n22885) );
  XNOR U22725 ( .A(n22701), .B(n22878), .Z(n22880) );
  XOR U22726 ( .A(n22887), .B(n22888), .Z(n22701) );
  AND U22727 ( .A(n821), .B(n22889), .Z(n22888) );
  XOR U22728 ( .A(n22887), .B(n22890), .Z(n22889) );
  IV U22729 ( .A(n22882), .Z(n22878) );
  AND U22730 ( .A(n22709), .B(n22712), .Z(n22882) );
  XNOR U22731 ( .A(n22891), .B(n22892), .Z(n22712) );
  AND U22732 ( .A(n823), .B(n22893), .Z(n22892) );
  XNOR U22733 ( .A(n22894), .B(n22891), .Z(n22893) );
  XOR U22734 ( .A(n22895), .B(n22896), .Z(n823) );
  AND U22735 ( .A(n22897), .B(n22898), .Z(n22896) );
  XNOR U22736 ( .A(n22718), .B(n22895), .Z(n22898) );
  AND U22737 ( .A(n22899), .B(n22900), .Z(n22718) );
  XOR U22738 ( .A(n22895), .B(n22719), .Z(n22897) );
  AND U22739 ( .A(n22901), .B(n22902), .Z(n22719) );
  XOR U22740 ( .A(n22903), .B(n22904), .Z(n22895) );
  AND U22741 ( .A(n22905), .B(n22906), .Z(n22904) );
  XOR U22742 ( .A(n22903), .B(n22729), .Z(n22906) );
  XOR U22743 ( .A(n22907), .B(n22908), .Z(n22729) );
  AND U22744 ( .A(n543), .B(n22909), .Z(n22908) );
  XOR U22745 ( .A(n22910), .B(n22907), .Z(n22909) );
  XNOR U22746 ( .A(n22726), .B(n22903), .Z(n22905) );
  XOR U22747 ( .A(n22911), .B(n22912), .Z(n22726) );
  AND U22748 ( .A(n541), .B(n22913), .Z(n22912) );
  XOR U22749 ( .A(n22914), .B(n22911), .Z(n22913) );
  XOR U22750 ( .A(n22915), .B(n22916), .Z(n22903) );
  AND U22751 ( .A(n22917), .B(n22918), .Z(n22916) );
  XOR U22752 ( .A(n22915), .B(n22741), .Z(n22918) );
  XOR U22753 ( .A(n22919), .B(n22920), .Z(n22741) );
  AND U22754 ( .A(n543), .B(n22921), .Z(n22920) );
  XOR U22755 ( .A(n22922), .B(n22919), .Z(n22921) );
  XNOR U22756 ( .A(n22738), .B(n22915), .Z(n22917) );
  XOR U22757 ( .A(n22923), .B(n22924), .Z(n22738) );
  AND U22758 ( .A(n541), .B(n22925), .Z(n22924) );
  XOR U22759 ( .A(n22926), .B(n22923), .Z(n22925) );
  XOR U22760 ( .A(n22927), .B(n22928), .Z(n22915) );
  AND U22761 ( .A(n22929), .B(n22930), .Z(n22928) );
  XOR U22762 ( .A(n22927), .B(n22753), .Z(n22930) );
  XOR U22763 ( .A(n22931), .B(n22932), .Z(n22753) );
  AND U22764 ( .A(n543), .B(n22933), .Z(n22932) );
  XOR U22765 ( .A(n22934), .B(n22931), .Z(n22933) );
  XNOR U22766 ( .A(n22750), .B(n22927), .Z(n22929) );
  XOR U22767 ( .A(n22935), .B(n22936), .Z(n22750) );
  AND U22768 ( .A(n541), .B(n22937), .Z(n22936) );
  XOR U22769 ( .A(n22938), .B(n22935), .Z(n22937) );
  XOR U22770 ( .A(n22939), .B(n22940), .Z(n22927) );
  AND U22771 ( .A(n22941), .B(n22942), .Z(n22940) );
  XOR U22772 ( .A(n22939), .B(n22765), .Z(n22942) );
  XOR U22773 ( .A(n22943), .B(n22944), .Z(n22765) );
  AND U22774 ( .A(n543), .B(n22945), .Z(n22944) );
  XOR U22775 ( .A(n22946), .B(n22943), .Z(n22945) );
  XNOR U22776 ( .A(n22762), .B(n22939), .Z(n22941) );
  XOR U22777 ( .A(n22947), .B(n22948), .Z(n22762) );
  AND U22778 ( .A(n541), .B(n22949), .Z(n22948) );
  XOR U22779 ( .A(n22950), .B(n22947), .Z(n22949) );
  XOR U22780 ( .A(n22951), .B(n22952), .Z(n22939) );
  AND U22781 ( .A(n22953), .B(n22954), .Z(n22952) );
  XOR U22782 ( .A(n22951), .B(n22777), .Z(n22954) );
  XOR U22783 ( .A(n22955), .B(n22956), .Z(n22777) );
  AND U22784 ( .A(n543), .B(n22957), .Z(n22956) );
  XOR U22785 ( .A(n22958), .B(n22955), .Z(n22957) );
  XNOR U22786 ( .A(n22774), .B(n22951), .Z(n22953) );
  XOR U22787 ( .A(n22959), .B(n22960), .Z(n22774) );
  AND U22788 ( .A(n541), .B(n22961), .Z(n22960) );
  XOR U22789 ( .A(n22962), .B(n22959), .Z(n22961) );
  XOR U22790 ( .A(n22963), .B(n22964), .Z(n22951) );
  AND U22791 ( .A(n22965), .B(n22966), .Z(n22964) );
  XOR U22792 ( .A(n22963), .B(n22789), .Z(n22966) );
  XOR U22793 ( .A(n22967), .B(n22968), .Z(n22789) );
  AND U22794 ( .A(n543), .B(n22969), .Z(n22968) );
  XOR U22795 ( .A(n22970), .B(n22967), .Z(n22969) );
  XNOR U22796 ( .A(n22786), .B(n22963), .Z(n22965) );
  XOR U22797 ( .A(n22971), .B(n22972), .Z(n22786) );
  AND U22798 ( .A(n541), .B(n22973), .Z(n22972) );
  XOR U22799 ( .A(n22974), .B(n22971), .Z(n22973) );
  XOR U22800 ( .A(n22975), .B(n22976), .Z(n22963) );
  AND U22801 ( .A(n22977), .B(n22978), .Z(n22976) );
  XOR U22802 ( .A(n22975), .B(n22801), .Z(n22978) );
  XOR U22803 ( .A(n22979), .B(n22980), .Z(n22801) );
  AND U22804 ( .A(n543), .B(n22981), .Z(n22980) );
  XOR U22805 ( .A(n22982), .B(n22979), .Z(n22981) );
  XNOR U22806 ( .A(n22798), .B(n22975), .Z(n22977) );
  XOR U22807 ( .A(n22983), .B(n22984), .Z(n22798) );
  AND U22808 ( .A(n541), .B(n22985), .Z(n22984) );
  XOR U22809 ( .A(n22986), .B(n22983), .Z(n22985) );
  XOR U22810 ( .A(n22987), .B(n22988), .Z(n22975) );
  AND U22811 ( .A(n22989), .B(n22990), .Z(n22988) );
  XOR U22812 ( .A(n22987), .B(n22813), .Z(n22990) );
  XOR U22813 ( .A(n22991), .B(n22992), .Z(n22813) );
  AND U22814 ( .A(n543), .B(n22993), .Z(n22992) );
  XOR U22815 ( .A(n22994), .B(n22991), .Z(n22993) );
  XNOR U22816 ( .A(n22810), .B(n22987), .Z(n22989) );
  XOR U22817 ( .A(n22995), .B(n22996), .Z(n22810) );
  AND U22818 ( .A(n541), .B(n22997), .Z(n22996) );
  XOR U22819 ( .A(n22998), .B(n22995), .Z(n22997) );
  XOR U22820 ( .A(n22999), .B(n23000), .Z(n22987) );
  AND U22821 ( .A(n23001), .B(n23002), .Z(n23000) );
  XOR U22822 ( .A(n22999), .B(n22825), .Z(n23002) );
  XOR U22823 ( .A(n23003), .B(n23004), .Z(n22825) );
  AND U22824 ( .A(n543), .B(n23005), .Z(n23004) );
  XOR U22825 ( .A(n23006), .B(n23003), .Z(n23005) );
  XNOR U22826 ( .A(n22822), .B(n22999), .Z(n23001) );
  XOR U22827 ( .A(n23007), .B(n23008), .Z(n22822) );
  AND U22828 ( .A(n541), .B(n23009), .Z(n23008) );
  XOR U22829 ( .A(n23010), .B(n23007), .Z(n23009) );
  XOR U22830 ( .A(n23011), .B(n23012), .Z(n22999) );
  AND U22831 ( .A(n23013), .B(n23014), .Z(n23012) );
  XOR U22832 ( .A(n23011), .B(n22837), .Z(n23014) );
  XOR U22833 ( .A(n23015), .B(n23016), .Z(n22837) );
  AND U22834 ( .A(n543), .B(n23017), .Z(n23016) );
  XOR U22835 ( .A(n23018), .B(n23015), .Z(n23017) );
  XNOR U22836 ( .A(n22834), .B(n23011), .Z(n23013) );
  XOR U22837 ( .A(n23019), .B(n23020), .Z(n22834) );
  AND U22838 ( .A(n541), .B(n23021), .Z(n23020) );
  XOR U22839 ( .A(n23022), .B(n23019), .Z(n23021) );
  XOR U22840 ( .A(n23023), .B(n23024), .Z(n23011) );
  AND U22841 ( .A(n23025), .B(n23026), .Z(n23024) );
  XOR U22842 ( .A(n23023), .B(n22849), .Z(n23026) );
  XOR U22843 ( .A(n23027), .B(n23028), .Z(n22849) );
  AND U22844 ( .A(n543), .B(n23029), .Z(n23028) );
  XOR U22845 ( .A(n23030), .B(n23027), .Z(n23029) );
  XNOR U22846 ( .A(n22846), .B(n23023), .Z(n23025) );
  XOR U22847 ( .A(n23031), .B(n23032), .Z(n22846) );
  AND U22848 ( .A(n541), .B(n23033), .Z(n23032) );
  XOR U22849 ( .A(n23034), .B(n23031), .Z(n23033) );
  XOR U22850 ( .A(n23035), .B(n23036), .Z(n23023) );
  AND U22851 ( .A(n23037), .B(n23038), .Z(n23036) );
  XOR U22852 ( .A(n23035), .B(n22861), .Z(n23038) );
  XOR U22853 ( .A(n23039), .B(n23040), .Z(n22861) );
  AND U22854 ( .A(n543), .B(n23041), .Z(n23040) );
  XOR U22855 ( .A(n23042), .B(n23039), .Z(n23041) );
  XNOR U22856 ( .A(n22858), .B(n23035), .Z(n23037) );
  XOR U22857 ( .A(n23043), .B(n23044), .Z(n22858) );
  AND U22858 ( .A(n541), .B(n23045), .Z(n23044) );
  XOR U22859 ( .A(n23046), .B(n23043), .Z(n23045) );
  XOR U22860 ( .A(n23047), .B(n23048), .Z(n23035) );
  AND U22861 ( .A(n23049), .B(n23050), .Z(n23048) );
  XOR U22862 ( .A(n23047), .B(n22873), .Z(n23050) );
  XOR U22863 ( .A(n23051), .B(n23052), .Z(n22873) );
  AND U22864 ( .A(n543), .B(n23053), .Z(n23052) );
  XOR U22865 ( .A(n23054), .B(n23051), .Z(n23053) );
  XNOR U22866 ( .A(n22870), .B(n23047), .Z(n23049) );
  XOR U22867 ( .A(n23055), .B(n23056), .Z(n22870) );
  AND U22868 ( .A(n541), .B(n23057), .Z(n23056) );
  XOR U22869 ( .A(n23058), .B(n23055), .Z(n23057) );
  XOR U22870 ( .A(n23059), .B(n23060), .Z(n23047) );
  AND U22871 ( .A(n23061), .B(n23062), .Z(n23060) );
  XNOR U22872 ( .A(n23063), .B(n22886), .Z(n23062) );
  XOR U22873 ( .A(n23064), .B(n23065), .Z(n22886) );
  AND U22874 ( .A(n543), .B(n23066), .Z(n23065) );
  XOR U22875 ( .A(n23064), .B(n23067), .Z(n23066) );
  XNOR U22876 ( .A(n22883), .B(n23059), .Z(n23061) );
  XOR U22877 ( .A(n23068), .B(n23069), .Z(n22883) );
  AND U22878 ( .A(n541), .B(n23070), .Z(n23069) );
  XOR U22879 ( .A(n23068), .B(n23071), .Z(n23070) );
  IV U22880 ( .A(n23063), .Z(n23059) );
  AND U22881 ( .A(n22891), .B(n22894), .Z(n23063) );
  XNOR U22882 ( .A(n23072), .B(n23073), .Z(n22894) );
  AND U22883 ( .A(n543), .B(n23074), .Z(n23073) );
  XNOR U22884 ( .A(n23075), .B(n23072), .Z(n23074) );
  XOR U22885 ( .A(n23076), .B(n23077), .Z(n543) );
  AND U22886 ( .A(n23078), .B(n23079), .Z(n23077) );
  XNOR U22887 ( .A(n22899), .B(n23076), .Z(n23079) );
  AND U22888 ( .A(p_input[1023]), .B(p_input[1007]), .Z(n22899) );
  XOR U22889 ( .A(n23076), .B(n22900), .Z(n23078) );
  AND U22890 ( .A(p_input[991]), .B(p_input[975]), .Z(n22900) );
  XOR U22891 ( .A(n23080), .B(n23081), .Z(n23076) );
  AND U22892 ( .A(n23082), .B(n23083), .Z(n23081) );
  XOR U22893 ( .A(n23080), .B(n22910), .Z(n23083) );
  XNOR U22894 ( .A(p_input[1006]), .B(n23084), .Z(n22910) );
  AND U22895 ( .A(n859), .B(n23085), .Z(n23084) );
  XOR U22896 ( .A(p_input[1022]), .B(p_input[1006]), .Z(n23085) );
  XNOR U22897 ( .A(n22907), .B(n23080), .Z(n23082) );
  XOR U22898 ( .A(n23086), .B(n23087), .Z(n22907) );
  AND U22899 ( .A(n857), .B(n23088), .Z(n23087) );
  XOR U22900 ( .A(p_input[990]), .B(p_input[974]), .Z(n23088) );
  XOR U22901 ( .A(n23089), .B(n23090), .Z(n23080) );
  AND U22902 ( .A(n23091), .B(n23092), .Z(n23090) );
  XOR U22903 ( .A(n23089), .B(n22922), .Z(n23092) );
  XNOR U22904 ( .A(p_input[1005]), .B(n23093), .Z(n22922) );
  AND U22905 ( .A(n859), .B(n23094), .Z(n23093) );
  XOR U22906 ( .A(p_input[1021]), .B(p_input[1005]), .Z(n23094) );
  XNOR U22907 ( .A(n22919), .B(n23089), .Z(n23091) );
  XOR U22908 ( .A(n23095), .B(n23096), .Z(n22919) );
  AND U22909 ( .A(n857), .B(n23097), .Z(n23096) );
  XOR U22910 ( .A(p_input[989]), .B(p_input[973]), .Z(n23097) );
  XOR U22911 ( .A(n23098), .B(n23099), .Z(n23089) );
  AND U22912 ( .A(n23100), .B(n23101), .Z(n23099) );
  XOR U22913 ( .A(n23098), .B(n22934), .Z(n23101) );
  XNOR U22914 ( .A(p_input[1004]), .B(n23102), .Z(n22934) );
  AND U22915 ( .A(n859), .B(n23103), .Z(n23102) );
  XOR U22916 ( .A(p_input[1020]), .B(p_input[1004]), .Z(n23103) );
  XNOR U22917 ( .A(n22931), .B(n23098), .Z(n23100) );
  XOR U22918 ( .A(n23104), .B(n23105), .Z(n22931) );
  AND U22919 ( .A(n857), .B(n23106), .Z(n23105) );
  XOR U22920 ( .A(p_input[988]), .B(p_input[972]), .Z(n23106) );
  XOR U22921 ( .A(n23107), .B(n23108), .Z(n23098) );
  AND U22922 ( .A(n23109), .B(n23110), .Z(n23108) );
  XOR U22923 ( .A(n23107), .B(n22946), .Z(n23110) );
  XNOR U22924 ( .A(p_input[1003]), .B(n23111), .Z(n22946) );
  AND U22925 ( .A(n859), .B(n23112), .Z(n23111) );
  XOR U22926 ( .A(p_input[1019]), .B(p_input[1003]), .Z(n23112) );
  XNOR U22927 ( .A(n22943), .B(n23107), .Z(n23109) );
  XOR U22928 ( .A(n23113), .B(n23114), .Z(n22943) );
  AND U22929 ( .A(n857), .B(n23115), .Z(n23114) );
  XOR U22930 ( .A(p_input[987]), .B(p_input[971]), .Z(n23115) );
  XOR U22931 ( .A(n23116), .B(n23117), .Z(n23107) );
  AND U22932 ( .A(n23118), .B(n23119), .Z(n23117) );
  XOR U22933 ( .A(n23116), .B(n22958), .Z(n23119) );
  XNOR U22934 ( .A(p_input[1002]), .B(n23120), .Z(n22958) );
  AND U22935 ( .A(n859), .B(n23121), .Z(n23120) );
  XOR U22936 ( .A(p_input[1018]), .B(p_input[1002]), .Z(n23121) );
  XNOR U22937 ( .A(n22955), .B(n23116), .Z(n23118) );
  XOR U22938 ( .A(n23122), .B(n23123), .Z(n22955) );
  AND U22939 ( .A(n857), .B(n23124), .Z(n23123) );
  XOR U22940 ( .A(p_input[986]), .B(p_input[970]), .Z(n23124) );
  XOR U22941 ( .A(n23125), .B(n23126), .Z(n23116) );
  AND U22942 ( .A(n23127), .B(n23128), .Z(n23126) );
  XOR U22943 ( .A(n23125), .B(n22970), .Z(n23128) );
  XNOR U22944 ( .A(p_input[1001]), .B(n23129), .Z(n22970) );
  AND U22945 ( .A(n859), .B(n23130), .Z(n23129) );
  XOR U22946 ( .A(p_input[1017]), .B(p_input[1001]), .Z(n23130) );
  XNOR U22947 ( .A(n22967), .B(n23125), .Z(n23127) );
  XOR U22948 ( .A(n23131), .B(n23132), .Z(n22967) );
  AND U22949 ( .A(n857), .B(n23133), .Z(n23132) );
  XOR U22950 ( .A(p_input[985]), .B(p_input[969]), .Z(n23133) );
  XOR U22951 ( .A(n23134), .B(n23135), .Z(n23125) );
  AND U22952 ( .A(n23136), .B(n23137), .Z(n23135) );
  XOR U22953 ( .A(n23134), .B(n22982), .Z(n23137) );
  XNOR U22954 ( .A(p_input[1000]), .B(n23138), .Z(n22982) );
  AND U22955 ( .A(n859), .B(n23139), .Z(n23138) );
  XOR U22956 ( .A(p_input[1016]), .B(p_input[1000]), .Z(n23139) );
  XNOR U22957 ( .A(n22979), .B(n23134), .Z(n23136) );
  XOR U22958 ( .A(n23140), .B(n23141), .Z(n22979) );
  AND U22959 ( .A(n857), .B(n23142), .Z(n23141) );
  XOR U22960 ( .A(p_input[984]), .B(p_input[968]), .Z(n23142) );
  XOR U22961 ( .A(n23143), .B(n23144), .Z(n23134) );
  AND U22962 ( .A(n23145), .B(n23146), .Z(n23144) );
  XOR U22963 ( .A(n23143), .B(n22994), .Z(n23146) );
  XNOR U22964 ( .A(p_input[999]), .B(n23147), .Z(n22994) );
  AND U22965 ( .A(n859), .B(n23148), .Z(n23147) );
  XOR U22966 ( .A(p_input[999]), .B(p_input[1015]), .Z(n23148) );
  XNOR U22967 ( .A(n22991), .B(n23143), .Z(n23145) );
  XOR U22968 ( .A(n23149), .B(n23150), .Z(n22991) );
  AND U22969 ( .A(n857), .B(n23151), .Z(n23150) );
  XOR U22970 ( .A(p_input[983]), .B(p_input[967]), .Z(n23151) );
  XOR U22971 ( .A(n23152), .B(n23153), .Z(n23143) );
  AND U22972 ( .A(n23154), .B(n23155), .Z(n23153) );
  XOR U22973 ( .A(n23152), .B(n23006), .Z(n23155) );
  XNOR U22974 ( .A(p_input[998]), .B(n23156), .Z(n23006) );
  AND U22975 ( .A(n859), .B(n23157), .Z(n23156) );
  XOR U22976 ( .A(p_input[998]), .B(p_input[1014]), .Z(n23157) );
  XNOR U22977 ( .A(n23003), .B(n23152), .Z(n23154) );
  XOR U22978 ( .A(n23158), .B(n23159), .Z(n23003) );
  AND U22979 ( .A(n857), .B(n23160), .Z(n23159) );
  XOR U22980 ( .A(p_input[982]), .B(p_input[966]), .Z(n23160) );
  XOR U22981 ( .A(n23161), .B(n23162), .Z(n23152) );
  AND U22982 ( .A(n23163), .B(n23164), .Z(n23162) );
  XOR U22983 ( .A(n23161), .B(n23018), .Z(n23164) );
  XNOR U22984 ( .A(p_input[997]), .B(n23165), .Z(n23018) );
  AND U22985 ( .A(n859), .B(n23166), .Z(n23165) );
  XOR U22986 ( .A(p_input[997]), .B(p_input[1013]), .Z(n23166) );
  XNOR U22987 ( .A(n23015), .B(n23161), .Z(n23163) );
  XOR U22988 ( .A(n23167), .B(n23168), .Z(n23015) );
  AND U22989 ( .A(n857), .B(n23169), .Z(n23168) );
  XOR U22990 ( .A(p_input[981]), .B(p_input[965]), .Z(n23169) );
  XOR U22991 ( .A(n23170), .B(n23171), .Z(n23161) );
  AND U22992 ( .A(n23172), .B(n23173), .Z(n23171) );
  XOR U22993 ( .A(n23170), .B(n23030), .Z(n23173) );
  XNOR U22994 ( .A(p_input[996]), .B(n23174), .Z(n23030) );
  AND U22995 ( .A(n859), .B(n23175), .Z(n23174) );
  XOR U22996 ( .A(p_input[996]), .B(p_input[1012]), .Z(n23175) );
  XNOR U22997 ( .A(n23027), .B(n23170), .Z(n23172) );
  XOR U22998 ( .A(n23176), .B(n23177), .Z(n23027) );
  AND U22999 ( .A(n857), .B(n23178), .Z(n23177) );
  XOR U23000 ( .A(p_input[980]), .B(p_input[964]), .Z(n23178) );
  XOR U23001 ( .A(n23179), .B(n23180), .Z(n23170) );
  AND U23002 ( .A(n23181), .B(n23182), .Z(n23180) );
  XOR U23003 ( .A(n23179), .B(n23042), .Z(n23182) );
  XNOR U23004 ( .A(p_input[995]), .B(n23183), .Z(n23042) );
  AND U23005 ( .A(n859), .B(n23184), .Z(n23183) );
  XOR U23006 ( .A(p_input[995]), .B(p_input[1011]), .Z(n23184) );
  XNOR U23007 ( .A(n23039), .B(n23179), .Z(n23181) );
  XOR U23008 ( .A(n23185), .B(n23186), .Z(n23039) );
  AND U23009 ( .A(n857), .B(n23187), .Z(n23186) );
  XOR U23010 ( .A(p_input[979]), .B(p_input[963]), .Z(n23187) );
  XOR U23011 ( .A(n23188), .B(n23189), .Z(n23179) );
  AND U23012 ( .A(n23190), .B(n23191), .Z(n23189) );
  XOR U23013 ( .A(n23188), .B(n23054), .Z(n23191) );
  XNOR U23014 ( .A(p_input[994]), .B(n23192), .Z(n23054) );
  AND U23015 ( .A(n859), .B(n23193), .Z(n23192) );
  XOR U23016 ( .A(p_input[994]), .B(p_input[1010]), .Z(n23193) );
  XNOR U23017 ( .A(n23051), .B(n23188), .Z(n23190) );
  XOR U23018 ( .A(n23194), .B(n23195), .Z(n23051) );
  AND U23019 ( .A(n857), .B(n23196), .Z(n23195) );
  XOR U23020 ( .A(p_input[978]), .B(p_input[962]), .Z(n23196) );
  XOR U23021 ( .A(n23197), .B(n23198), .Z(n23188) );
  AND U23022 ( .A(n23199), .B(n23200), .Z(n23198) );
  XNOR U23023 ( .A(n23201), .B(n23067), .Z(n23200) );
  XNOR U23024 ( .A(p_input[993]), .B(n23202), .Z(n23067) );
  AND U23025 ( .A(n859), .B(n23203), .Z(n23202) );
  XNOR U23026 ( .A(n23204), .B(p_input[1009]), .Z(n23203) );
  IV U23027 ( .A(p_input[993]), .Z(n23204) );
  XNOR U23028 ( .A(n23064), .B(n23197), .Z(n23199) );
  XNOR U23029 ( .A(p_input[961]), .B(n23205), .Z(n23064) );
  AND U23030 ( .A(n857), .B(n23206), .Z(n23205) );
  XOR U23031 ( .A(p_input[977]), .B(p_input[961]), .Z(n23206) );
  IV U23032 ( .A(n23201), .Z(n23197) );
  AND U23033 ( .A(n23072), .B(n23075), .Z(n23201) );
  XOR U23034 ( .A(p_input[992]), .B(n23207), .Z(n23075) );
  AND U23035 ( .A(n859), .B(n23208), .Z(n23207) );
  XOR U23036 ( .A(p_input[992]), .B(p_input[1008]), .Z(n23208) );
  XOR U23037 ( .A(n23209), .B(n23210), .Z(n859) );
  AND U23038 ( .A(n23211), .B(n23212), .Z(n23210) );
  XNOR U23039 ( .A(p_input[1023]), .B(n23209), .Z(n23212) );
  XOR U23040 ( .A(n23209), .B(p_input[1007]), .Z(n23211) );
  XOR U23041 ( .A(n23213), .B(n23214), .Z(n23209) );
  AND U23042 ( .A(n23215), .B(n23216), .Z(n23214) );
  XNOR U23043 ( .A(p_input[1022]), .B(n23213), .Z(n23216) );
  XOR U23044 ( .A(n23213), .B(p_input[1006]), .Z(n23215) );
  XOR U23045 ( .A(n23217), .B(n23218), .Z(n23213) );
  AND U23046 ( .A(n23219), .B(n23220), .Z(n23218) );
  XNOR U23047 ( .A(p_input[1021]), .B(n23217), .Z(n23220) );
  XOR U23048 ( .A(n23217), .B(p_input[1005]), .Z(n23219) );
  XOR U23049 ( .A(n23221), .B(n23222), .Z(n23217) );
  AND U23050 ( .A(n23223), .B(n23224), .Z(n23222) );
  XNOR U23051 ( .A(p_input[1020]), .B(n23221), .Z(n23224) );
  XOR U23052 ( .A(n23221), .B(p_input[1004]), .Z(n23223) );
  XOR U23053 ( .A(n23225), .B(n23226), .Z(n23221) );
  AND U23054 ( .A(n23227), .B(n23228), .Z(n23226) );
  XNOR U23055 ( .A(p_input[1019]), .B(n23225), .Z(n23228) );
  XOR U23056 ( .A(n23225), .B(p_input[1003]), .Z(n23227) );
  XOR U23057 ( .A(n23229), .B(n23230), .Z(n23225) );
  AND U23058 ( .A(n23231), .B(n23232), .Z(n23230) );
  XNOR U23059 ( .A(p_input[1018]), .B(n23229), .Z(n23232) );
  XOR U23060 ( .A(n23229), .B(p_input[1002]), .Z(n23231) );
  XOR U23061 ( .A(n23233), .B(n23234), .Z(n23229) );
  AND U23062 ( .A(n23235), .B(n23236), .Z(n23234) );
  XNOR U23063 ( .A(p_input[1017]), .B(n23233), .Z(n23236) );
  XOR U23064 ( .A(n23233), .B(p_input[1001]), .Z(n23235) );
  XOR U23065 ( .A(n23237), .B(n23238), .Z(n23233) );
  AND U23066 ( .A(n23239), .B(n23240), .Z(n23238) );
  XNOR U23067 ( .A(p_input[1016]), .B(n23237), .Z(n23240) );
  XOR U23068 ( .A(n23237), .B(p_input[1000]), .Z(n23239) );
  XOR U23069 ( .A(n23241), .B(n23242), .Z(n23237) );
  AND U23070 ( .A(n23243), .B(n23244), .Z(n23242) );
  XNOR U23071 ( .A(p_input[1015]), .B(n23241), .Z(n23244) );
  XOR U23072 ( .A(n23241), .B(p_input[999]), .Z(n23243) );
  XOR U23073 ( .A(n23245), .B(n23246), .Z(n23241) );
  AND U23074 ( .A(n23247), .B(n23248), .Z(n23246) );
  XNOR U23075 ( .A(p_input[1014]), .B(n23245), .Z(n23248) );
  XOR U23076 ( .A(n23245), .B(p_input[998]), .Z(n23247) );
  XOR U23077 ( .A(n23249), .B(n23250), .Z(n23245) );
  AND U23078 ( .A(n23251), .B(n23252), .Z(n23250) );
  XNOR U23079 ( .A(p_input[1013]), .B(n23249), .Z(n23252) );
  XOR U23080 ( .A(n23249), .B(p_input[997]), .Z(n23251) );
  XOR U23081 ( .A(n23253), .B(n23254), .Z(n23249) );
  AND U23082 ( .A(n23255), .B(n23256), .Z(n23254) );
  XNOR U23083 ( .A(p_input[1012]), .B(n23253), .Z(n23256) );
  XOR U23084 ( .A(n23253), .B(p_input[996]), .Z(n23255) );
  XOR U23085 ( .A(n23257), .B(n23258), .Z(n23253) );
  AND U23086 ( .A(n23259), .B(n23260), .Z(n23258) );
  XNOR U23087 ( .A(p_input[1011]), .B(n23257), .Z(n23260) );
  XOR U23088 ( .A(n23257), .B(p_input[995]), .Z(n23259) );
  XOR U23089 ( .A(n23261), .B(n23262), .Z(n23257) );
  AND U23090 ( .A(n23263), .B(n23264), .Z(n23262) );
  XNOR U23091 ( .A(p_input[1010]), .B(n23261), .Z(n23264) );
  XOR U23092 ( .A(n23261), .B(p_input[994]), .Z(n23263) );
  XNOR U23093 ( .A(n23265), .B(n23266), .Z(n23261) );
  AND U23094 ( .A(n23267), .B(n23268), .Z(n23266) );
  XOR U23095 ( .A(p_input[1009]), .B(n23265), .Z(n23268) );
  XNOR U23096 ( .A(p_input[993]), .B(n23265), .Z(n23267) );
  AND U23097 ( .A(p_input[1008]), .B(n23269), .Z(n23265) );
  IV U23098 ( .A(p_input[992]), .Z(n23269) );
  XNOR U23099 ( .A(p_input[960]), .B(n23270), .Z(n23072) );
  AND U23100 ( .A(n857), .B(n23271), .Z(n23270) );
  XOR U23101 ( .A(p_input[976]), .B(p_input[960]), .Z(n23271) );
  XOR U23102 ( .A(n23272), .B(n23273), .Z(n857) );
  AND U23103 ( .A(n23274), .B(n23275), .Z(n23273) );
  XNOR U23104 ( .A(p_input[991]), .B(n23272), .Z(n23275) );
  XOR U23105 ( .A(n23272), .B(p_input[975]), .Z(n23274) );
  XOR U23106 ( .A(n23276), .B(n23277), .Z(n23272) );
  AND U23107 ( .A(n23278), .B(n23279), .Z(n23277) );
  XNOR U23108 ( .A(p_input[990]), .B(n23276), .Z(n23279) );
  XNOR U23109 ( .A(n23276), .B(n23086), .Z(n23278) );
  IV U23110 ( .A(p_input[974]), .Z(n23086) );
  XOR U23111 ( .A(n23280), .B(n23281), .Z(n23276) );
  AND U23112 ( .A(n23282), .B(n23283), .Z(n23281) );
  XNOR U23113 ( .A(p_input[989]), .B(n23280), .Z(n23283) );
  XNOR U23114 ( .A(n23280), .B(n23095), .Z(n23282) );
  IV U23115 ( .A(p_input[973]), .Z(n23095) );
  XOR U23116 ( .A(n23284), .B(n23285), .Z(n23280) );
  AND U23117 ( .A(n23286), .B(n23287), .Z(n23285) );
  XNOR U23118 ( .A(p_input[988]), .B(n23284), .Z(n23287) );
  XNOR U23119 ( .A(n23284), .B(n23104), .Z(n23286) );
  IV U23120 ( .A(p_input[972]), .Z(n23104) );
  XOR U23121 ( .A(n23288), .B(n23289), .Z(n23284) );
  AND U23122 ( .A(n23290), .B(n23291), .Z(n23289) );
  XNOR U23123 ( .A(p_input[987]), .B(n23288), .Z(n23291) );
  XNOR U23124 ( .A(n23288), .B(n23113), .Z(n23290) );
  IV U23125 ( .A(p_input[971]), .Z(n23113) );
  XOR U23126 ( .A(n23292), .B(n23293), .Z(n23288) );
  AND U23127 ( .A(n23294), .B(n23295), .Z(n23293) );
  XNOR U23128 ( .A(p_input[986]), .B(n23292), .Z(n23295) );
  XNOR U23129 ( .A(n23292), .B(n23122), .Z(n23294) );
  IV U23130 ( .A(p_input[970]), .Z(n23122) );
  XOR U23131 ( .A(n23296), .B(n23297), .Z(n23292) );
  AND U23132 ( .A(n23298), .B(n23299), .Z(n23297) );
  XNOR U23133 ( .A(p_input[985]), .B(n23296), .Z(n23299) );
  XNOR U23134 ( .A(n23296), .B(n23131), .Z(n23298) );
  IV U23135 ( .A(p_input[969]), .Z(n23131) );
  XOR U23136 ( .A(n23300), .B(n23301), .Z(n23296) );
  AND U23137 ( .A(n23302), .B(n23303), .Z(n23301) );
  XNOR U23138 ( .A(p_input[984]), .B(n23300), .Z(n23303) );
  XNOR U23139 ( .A(n23300), .B(n23140), .Z(n23302) );
  IV U23140 ( .A(p_input[968]), .Z(n23140) );
  XOR U23141 ( .A(n23304), .B(n23305), .Z(n23300) );
  AND U23142 ( .A(n23306), .B(n23307), .Z(n23305) );
  XNOR U23143 ( .A(p_input[983]), .B(n23304), .Z(n23307) );
  XNOR U23144 ( .A(n23304), .B(n23149), .Z(n23306) );
  IV U23145 ( .A(p_input[967]), .Z(n23149) );
  XOR U23146 ( .A(n23308), .B(n23309), .Z(n23304) );
  AND U23147 ( .A(n23310), .B(n23311), .Z(n23309) );
  XNOR U23148 ( .A(p_input[982]), .B(n23308), .Z(n23311) );
  XNOR U23149 ( .A(n23308), .B(n23158), .Z(n23310) );
  IV U23150 ( .A(p_input[966]), .Z(n23158) );
  XOR U23151 ( .A(n23312), .B(n23313), .Z(n23308) );
  AND U23152 ( .A(n23314), .B(n23315), .Z(n23313) );
  XNOR U23153 ( .A(p_input[981]), .B(n23312), .Z(n23315) );
  XNOR U23154 ( .A(n23312), .B(n23167), .Z(n23314) );
  IV U23155 ( .A(p_input[965]), .Z(n23167) );
  XOR U23156 ( .A(n23316), .B(n23317), .Z(n23312) );
  AND U23157 ( .A(n23318), .B(n23319), .Z(n23317) );
  XNOR U23158 ( .A(p_input[980]), .B(n23316), .Z(n23319) );
  XNOR U23159 ( .A(n23316), .B(n23176), .Z(n23318) );
  IV U23160 ( .A(p_input[964]), .Z(n23176) );
  XOR U23161 ( .A(n23320), .B(n23321), .Z(n23316) );
  AND U23162 ( .A(n23322), .B(n23323), .Z(n23321) );
  XNOR U23163 ( .A(p_input[979]), .B(n23320), .Z(n23323) );
  XNOR U23164 ( .A(n23320), .B(n23185), .Z(n23322) );
  IV U23165 ( .A(p_input[963]), .Z(n23185) );
  XOR U23166 ( .A(n23324), .B(n23325), .Z(n23320) );
  AND U23167 ( .A(n23326), .B(n23327), .Z(n23325) );
  XNOR U23168 ( .A(p_input[978]), .B(n23324), .Z(n23327) );
  XNOR U23169 ( .A(n23324), .B(n23194), .Z(n23326) );
  IV U23170 ( .A(p_input[962]), .Z(n23194) );
  XNOR U23171 ( .A(n23328), .B(n23329), .Z(n23324) );
  AND U23172 ( .A(n23330), .B(n23331), .Z(n23329) );
  XOR U23173 ( .A(p_input[977]), .B(n23328), .Z(n23331) );
  XNOR U23174 ( .A(p_input[961]), .B(n23328), .Z(n23330) );
  AND U23175 ( .A(p_input[976]), .B(n23332), .Z(n23328) );
  IV U23176 ( .A(p_input[960]), .Z(n23332) );
  XOR U23177 ( .A(n23333), .B(n23334), .Z(n22891) );
  AND U23178 ( .A(n541), .B(n23335), .Z(n23334) );
  XNOR U23179 ( .A(n23336), .B(n23333), .Z(n23335) );
  XOR U23180 ( .A(n23337), .B(n23338), .Z(n541) );
  AND U23181 ( .A(n23339), .B(n23340), .Z(n23338) );
  XNOR U23182 ( .A(n22901), .B(n23337), .Z(n23340) );
  AND U23183 ( .A(p_input[959]), .B(p_input[943]), .Z(n22901) );
  XOR U23184 ( .A(n23337), .B(n22902), .Z(n23339) );
  AND U23185 ( .A(p_input[927]), .B(p_input[911]), .Z(n22902) );
  XOR U23186 ( .A(n23341), .B(n23342), .Z(n23337) );
  AND U23187 ( .A(n23343), .B(n23344), .Z(n23342) );
  XOR U23188 ( .A(n23341), .B(n22914), .Z(n23344) );
  XNOR U23189 ( .A(p_input[942]), .B(n23345), .Z(n22914) );
  AND U23190 ( .A(n863), .B(n23346), .Z(n23345) );
  XOR U23191 ( .A(p_input[958]), .B(p_input[942]), .Z(n23346) );
  XNOR U23192 ( .A(n22911), .B(n23341), .Z(n23343) );
  XOR U23193 ( .A(n23347), .B(n23348), .Z(n22911) );
  AND U23194 ( .A(n860), .B(n23349), .Z(n23348) );
  XOR U23195 ( .A(p_input[926]), .B(p_input[910]), .Z(n23349) );
  XOR U23196 ( .A(n23350), .B(n23351), .Z(n23341) );
  AND U23197 ( .A(n23352), .B(n23353), .Z(n23351) );
  XOR U23198 ( .A(n23350), .B(n22926), .Z(n23353) );
  XNOR U23199 ( .A(p_input[941]), .B(n23354), .Z(n22926) );
  AND U23200 ( .A(n863), .B(n23355), .Z(n23354) );
  XOR U23201 ( .A(p_input[957]), .B(p_input[941]), .Z(n23355) );
  XNOR U23202 ( .A(n22923), .B(n23350), .Z(n23352) );
  XOR U23203 ( .A(n23356), .B(n23357), .Z(n22923) );
  AND U23204 ( .A(n860), .B(n23358), .Z(n23357) );
  XOR U23205 ( .A(p_input[925]), .B(p_input[909]), .Z(n23358) );
  XOR U23206 ( .A(n23359), .B(n23360), .Z(n23350) );
  AND U23207 ( .A(n23361), .B(n23362), .Z(n23360) );
  XOR U23208 ( .A(n23359), .B(n22938), .Z(n23362) );
  XNOR U23209 ( .A(p_input[940]), .B(n23363), .Z(n22938) );
  AND U23210 ( .A(n863), .B(n23364), .Z(n23363) );
  XOR U23211 ( .A(p_input[956]), .B(p_input[940]), .Z(n23364) );
  XNOR U23212 ( .A(n22935), .B(n23359), .Z(n23361) );
  XOR U23213 ( .A(n23365), .B(n23366), .Z(n22935) );
  AND U23214 ( .A(n860), .B(n23367), .Z(n23366) );
  XOR U23215 ( .A(p_input[924]), .B(p_input[908]), .Z(n23367) );
  XOR U23216 ( .A(n23368), .B(n23369), .Z(n23359) );
  AND U23217 ( .A(n23370), .B(n23371), .Z(n23369) );
  XOR U23218 ( .A(n23368), .B(n22950), .Z(n23371) );
  XNOR U23219 ( .A(p_input[939]), .B(n23372), .Z(n22950) );
  AND U23220 ( .A(n863), .B(n23373), .Z(n23372) );
  XOR U23221 ( .A(p_input[955]), .B(p_input[939]), .Z(n23373) );
  XNOR U23222 ( .A(n22947), .B(n23368), .Z(n23370) );
  XOR U23223 ( .A(n23374), .B(n23375), .Z(n22947) );
  AND U23224 ( .A(n860), .B(n23376), .Z(n23375) );
  XOR U23225 ( .A(p_input[923]), .B(p_input[907]), .Z(n23376) );
  XOR U23226 ( .A(n23377), .B(n23378), .Z(n23368) );
  AND U23227 ( .A(n23379), .B(n23380), .Z(n23378) );
  XOR U23228 ( .A(n23377), .B(n22962), .Z(n23380) );
  XNOR U23229 ( .A(p_input[938]), .B(n23381), .Z(n22962) );
  AND U23230 ( .A(n863), .B(n23382), .Z(n23381) );
  XOR U23231 ( .A(p_input[954]), .B(p_input[938]), .Z(n23382) );
  XNOR U23232 ( .A(n22959), .B(n23377), .Z(n23379) );
  XOR U23233 ( .A(n23383), .B(n23384), .Z(n22959) );
  AND U23234 ( .A(n860), .B(n23385), .Z(n23384) );
  XOR U23235 ( .A(p_input[922]), .B(p_input[906]), .Z(n23385) );
  XOR U23236 ( .A(n23386), .B(n23387), .Z(n23377) );
  AND U23237 ( .A(n23388), .B(n23389), .Z(n23387) );
  XOR U23238 ( .A(n23386), .B(n22974), .Z(n23389) );
  XNOR U23239 ( .A(p_input[937]), .B(n23390), .Z(n22974) );
  AND U23240 ( .A(n863), .B(n23391), .Z(n23390) );
  XOR U23241 ( .A(p_input[953]), .B(p_input[937]), .Z(n23391) );
  XNOR U23242 ( .A(n22971), .B(n23386), .Z(n23388) );
  XOR U23243 ( .A(n23392), .B(n23393), .Z(n22971) );
  AND U23244 ( .A(n860), .B(n23394), .Z(n23393) );
  XOR U23245 ( .A(p_input[921]), .B(p_input[905]), .Z(n23394) );
  XOR U23246 ( .A(n23395), .B(n23396), .Z(n23386) );
  AND U23247 ( .A(n23397), .B(n23398), .Z(n23396) );
  XOR U23248 ( .A(n23395), .B(n22986), .Z(n23398) );
  XNOR U23249 ( .A(p_input[936]), .B(n23399), .Z(n22986) );
  AND U23250 ( .A(n863), .B(n23400), .Z(n23399) );
  XOR U23251 ( .A(p_input[952]), .B(p_input[936]), .Z(n23400) );
  XNOR U23252 ( .A(n22983), .B(n23395), .Z(n23397) );
  XOR U23253 ( .A(n23401), .B(n23402), .Z(n22983) );
  AND U23254 ( .A(n860), .B(n23403), .Z(n23402) );
  XOR U23255 ( .A(p_input[920]), .B(p_input[904]), .Z(n23403) );
  XOR U23256 ( .A(n23404), .B(n23405), .Z(n23395) );
  AND U23257 ( .A(n23406), .B(n23407), .Z(n23405) );
  XOR U23258 ( .A(n23404), .B(n22998), .Z(n23407) );
  XNOR U23259 ( .A(p_input[935]), .B(n23408), .Z(n22998) );
  AND U23260 ( .A(n863), .B(n23409), .Z(n23408) );
  XOR U23261 ( .A(p_input[951]), .B(p_input[935]), .Z(n23409) );
  XNOR U23262 ( .A(n22995), .B(n23404), .Z(n23406) );
  XOR U23263 ( .A(n23410), .B(n23411), .Z(n22995) );
  AND U23264 ( .A(n860), .B(n23412), .Z(n23411) );
  XOR U23265 ( .A(p_input[919]), .B(p_input[903]), .Z(n23412) );
  XOR U23266 ( .A(n23413), .B(n23414), .Z(n23404) );
  AND U23267 ( .A(n23415), .B(n23416), .Z(n23414) );
  XOR U23268 ( .A(n23413), .B(n23010), .Z(n23416) );
  XNOR U23269 ( .A(p_input[934]), .B(n23417), .Z(n23010) );
  AND U23270 ( .A(n863), .B(n23418), .Z(n23417) );
  XOR U23271 ( .A(p_input[950]), .B(p_input[934]), .Z(n23418) );
  XNOR U23272 ( .A(n23007), .B(n23413), .Z(n23415) );
  XOR U23273 ( .A(n23419), .B(n23420), .Z(n23007) );
  AND U23274 ( .A(n860), .B(n23421), .Z(n23420) );
  XOR U23275 ( .A(p_input[918]), .B(p_input[902]), .Z(n23421) );
  XOR U23276 ( .A(n23422), .B(n23423), .Z(n23413) );
  AND U23277 ( .A(n23424), .B(n23425), .Z(n23423) );
  XOR U23278 ( .A(n23422), .B(n23022), .Z(n23425) );
  XNOR U23279 ( .A(p_input[933]), .B(n23426), .Z(n23022) );
  AND U23280 ( .A(n863), .B(n23427), .Z(n23426) );
  XOR U23281 ( .A(p_input[949]), .B(p_input[933]), .Z(n23427) );
  XNOR U23282 ( .A(n23019), .B(n23422), .Z(n23424) );
  XOR U23283 ( .A(n23428), .B(n23429), .Z(n23019) );
  AND U23284 ( .A(n860), .B(n23430), .Z(n23429) );
  XOR U23285 ( .A(p_input[917]), .B(p_input[901]), .Z(n23430) );
  XOR U23286 ( .A(n23431), .B(n23432), .Z(n23422) );
  AND U23287 ( .A(n23433), .B(n23434), .Z(n23432) );
  XOR U23288 ( .A(n23431), .B(n23034), .Z(n23434) );
  XNOR U23289 ( .A(p_input[932]), .B(n23435), .Z(n23034) );
  AND U23290 ( .A(n863), .B(n23436), .Z(n23435) );
  XOR U23291 ( .A(p_input[948]), .B(p_input[932]), .Z(n23436) );
  XNOR U23292 ( .A(n23031), .B(n23431), .Z(n23433) );
  XOR U23293 ( .A(n23437), .B(n23438), .Z(n23031) );
  AND U23294 ( .A(n860), .B(n23439), .Z(n23438) );
  XOR U23295 ( .A(p_input[916]), .B(p_input[900]), .Z(n23439) );
  XOR U23296 ( .A(n23440), .B(n23441), .Z(n23431) );
  AND U23297 ( .A(n23442), .B(n23443), .Z(n23441) );
  XOR U23298 ( .A(n23440), .B(n23046), .Z(n23443) );
  XNOR U23299 ( .A(p_input[931]), .B(n23444), .Z(n23046) );
  AND U23300 ( .A(n863), .B(n23445), .Z(n23444) );
  XOR U23301 ( .A(p_input[947]), .B(p_input[931]), .Z(n23445) );
  XNOR U23302 ( .A(n23043), .B(n23440), .Z(n23442) );
  XOR U23303 ( .A(n23446), .B(n23447), .Z(n23043) );
  AND U23304 ( .A(n860), .B(n23448), .Z(n23447) );
  XOR U23305 ( .A(p_input[915]), .B(p_input[899]), .Z(n23448) );
  XOR U23306 ( .A(n23449), .B(n23450), .Z(n23440) );
  AND U23307 ( .A(n23451), .B(n23452), .Z(n23450) );
  XOR U23308 ( .A(n23449), .B(n23058), .Z(n23452) );
  XNOR U23309 ( .A(p_input[930]), .B(n23453), .Z(n23058) );
  AND U23310 ( .A(n863), .B(n23454), .Z(n23453) );
  XOR U23311 ( .A(p_input[946]), .B(p_input[930]), .Z(n23454) );
  XNOR U23312 ( .A(n23055), .B(n23449), .Z(n23451) );
  XOR U23313 ( .A(n23455), .B(n23456), .Z(n23055) );
  AND U23314 ( .A(n860), .B(n23457), .Z(n23456) );
  XOR U23315 ( .A(p_input[914]), .B(p_input[898]), .Z(n23457) );
  XOR U23316 ( .A(n23458), .B(n23459), .Z(n23449) );
  AND U23317 ( .A(n23460), .B(n23461), .Z(n23459) );
  XNOR U23318 ( .A(n23462), .B(n23071), .Z(n23461) );
  XNOR U23319 ( .A(p_input[929]), .B(n23463), .Z(n23071) );
  AND U23320 ( .A(n863), .B(n23464), .Z(n23463) );
  XNOR U23321 ( .A(p_input[945]), .B(n23465), .Z(n23464) );
  IV U23322 ( .A(p_input[929]), .Z(n23465) );
  XNOR U23323 ( .A(n23068), .B(n23458), .Z(n23460) );
  XNOR U23324 ( .A(p_input[897]), .B(n23466), .Z(n23068) );
  AND U23325 ( .A(n860), .B(n23467), .Z(n23466) );
  XOR U23326 ( .A(p_input[913]), .B(p_input[897]), .Z(n23467) );
  IV U23327 ( .A(n23462), .Z(n23458) );
  AND U23328 ( .A(n23333), .B(n23336), .Z(n23462) );
  XOR U23329 ( .A(p_input[928]), .B(n23468), .Z(n23336) );
  AND U23330 ( .A(n863), .B(n23469), .Z(n23468) );
  XOR U23331 ( .A(p_input[944]), .B(p_input[928]), .Z(n23469) );
  XOR U23332 ( .A(n23470), .B(n23471), .Z(n863) );
  AND U23333 ( .A(n23472), .B(n23473), .Z(n23471) );
  XNOR U23334 ( .A(p_input[959]), .B(n23470), .Z(n23473) );
  XOR U23335 ( .A(n23470), .B(p_input[943]), .Z(n23472) );
  XOR U23336 ( .A(n23474), .B(n23475), .Z(n23470) );
  AND U23337 ( .A(n23476), .B(n23477), .Z(n23475) );
  XNOR U23338 ( .A(p_input[958]), .B(n23474), .Z(n23477) );
  XOR U23339 ( .A(n23474), .B(p_input[942]), .Z(n23476) );
  XOR U23340 ( .A(n23478), .B(n23479), .Z(n23474) );
  AND U23341 ( .A(n23480), .B(n23481), .Z(n23479) );
  XNOR U23342 ( .A(p_input[957]), .B(n23478), .Z(n23481) );
  XOR U23343 ( .A(n23478), .B(p_input[941]), .Z(n23480) );
  XOR U23344 ( .A(n23482), .B(n23483), .Z(n23478) );
  AND U23345 ( .A(n23484), .B(n23485), .Z(n23483) );
  XNOR U23346 ( .A(p_input[956]), .B(n23482), .Z(n23485) );
  XOR U23347 ( .A(n23482), .B(p_input[940]), .Z(n23484) );
  XOR U23348 ( .A(n23486), .B(n23487), .Z(n23482) );
  AND U23349 ( .A(n23488), .B(n23489), .Z(n23487) );
  XNOR U23350 ( .A(p_input[955]), .B(n23486), .Z(n23489) );
  XOR U23351 ( .A(n23486), .B(p_input[939]), .Z(n23488) );
  XOR U23352 ( .A(n23490), .B(n23491), .Z(n23486) );
  AND U23353 ( .A(n23492), .B(n23493), .Z(n23491) );
  XNOR U23354 ( .A(p_input[954]), .B(n23490), .Z(n23493) );
  XOR U23355 ( .A(n23490), .B(p_input[938]), .Z(n23492) );
  XOR U23356 ( .A(n23494), .B(n23495), .Z(n23490) );
  AND U23357 ( .A(n23496), .B(n23497), .Z(n23495) );
  XNOR U23358 ( .A(p_input[953]), .B(n23494), .Z(n23497) );
  XOR U23359 ( .A(n23494), .B(p_input[937]), .Z(n23496) );
  XOR U23360 ( .A(n23498), .B(n23499), .Z(n23494) );
  AND U23361 ( .A(n23500), .B(n23501), .Z(n23499) );
  XNOR U23362 ( .A(p_input[952]), .B(n23498), .Z(n23501) );
  XOR U23363 ( .A(n23498), .B(p_input[936]), .Z(n23500) );
  XOR U23364 ( .A(n23502), .B(n23503), .Z(n23498) );
  AND U23365 ( .A(n23504), .B(n23505), .Z(n23503) );
  XNOR U23366 ( .A(p_input[951]), .B(n23502), .Z(n23505) );
  XOR U23367 ( .A(n23502), .B(p_input[935]), .Z(n23504) );
  XOR U23368 ( .A(n23506), .B(n23507), .Z(n23502) );
  AND U23369 ( .A(n23508), .B(n23509), .Z(n23507) );
  XNOR U23370 ( .A(p_input[950]), .B(n23506), .Z(n23509) );
  XOR U23371 ( .A(n23506), .B(p_input[934]), .Z(n23508) );
  XOR U23372 ( .A(n23510), .B(n23511), .Z(n23506) );
  AND U23373 ( .A(n23512), .B(n23513), .Z(n23511) );
  XNOR U23374 ( .A(p_input[949]), .B(n23510), .Z(n23513) );
  XOR U23375 ( .A(n23510), .B(p_input[933]), .Z(n23512) );
  XOR U23376 ( .A(n23514), .B(n23515), .Z(n23510) );
  AND U23377 ( .A(n23516), .B(n23517), .Z(n23515) );
  XNOR U23378 ( .A(p_input[948]), .B(n23514), .Z(n23517) );
  XOR U23379 ( .A(n23514), .B(p_input[932]), .Z(n23516) );
  XOR U23380 ( .A(n23518), .B(n23519), .Z(n23514) );
  AND U23381 ( .A(n23520), .B(n23521), .Z(n23519) );
  XNOR U23382 ( .A(p_input[947]), .B(n23518), .Z(n23521) );
  XOR U23383 ( .A(n23518), .B(p_input[931]), .Z(n23520) );
  XOR U23384 ( .A(n23522), .B(n23523), .Z(n23518) );
  AND U23385 ( .A(n23524), .B(n23525), .Z(n23523) );
  XNOR U23386 ( .A(p_input[946]), .B(n23522), .Z(n23525) );
  XOR U23387 ( .A(n23522), .B(p_input[930]), .Z(n23524) );
  XNOR U23388 ( .A(n23526), .B(n23527), .Z(n23522) );
  AND U23389 ( .A(n23528), .B(n23529), .Z(n23527) );
  XOR U23390 ( .A(p_input[945]), .B(n23526), .Z(n23529) );
  XNOR U23391 ( .A(p_input[929]), .B(n23526), .Z(n23528) );
  AND U23392 ( .A(p_input[944]), .B(n23530), .Z(n23526) );
  IV U23393 ( .A(p_input[928]), .Z(n23530) );
  XNOR U23394 ( .A(p_input[896]), .B(n23531), .Z(n23333) );
  AND U23395 ( .A(n860), .B(n23532), .Z(n23531) );
  XOR U23396 ( .A(p_input[912]), .B(p_input[896]), .Z(n23532) );
  XOR U23397 ( .A(n23533), .B(n23534), .Z(n860) );
  AND U23398 ( .A(n23535), .B(n23536), .Z(n23534) );
  XNOR U23399 ( .A(p_input[927]), .B(n23533), .Z(n23536) );
  XOR U23400 ( .A(n23533), .B(p_input[911]), .Z(n23535) );
  XOR U23401 ( .A(n23537), .B(n23538), .Z(n23533) );
  AND U23402 ( .A(n23539), .B(n23540), .Z(n23538) );
  XNOR U23403 ( .A(p_input[926]), .B(n23537), .Z(n23540) );
  XNOR U23404 ( .A(n23537), .B(n23347), .Z(n23539) );
  IV U23405 ( .A(p_input[910]), .Z(n23347) );
  XOR U23406 ( .A(n23541), .B(n23542), .Z(n23537) );
  AND U23407 ( .A(n23543), .B(n23544), .Z(n23542) );
  XNOR U23408 ( .A(p_input[925]), .B(n23541), .Z(n23544) );
  XNOR U23409 ( .A(n23541), .B(n23356), .Z(n23543) );
  IV U23410 ( .A(p_input[909]), .Z(n23356) );
  XOR U23411 ( .A(n23545), .B(n23546), .Z(n23541) );
  AND U23412 ( .A(n23547), .B(n23548), .Z(n23546) );
  XNOR U23413 ( .A(p_input[924]), .B(n23545), .Z(n23548) );
  XNOR U23414 ( .A(n23545), .B(n23365), .Z(n23547) );
  IV U23415 ( .A(p_input[908]), .Z(n23365) );
  XOR U23416 ( .A(n23549), .B(n23550), .Z(n23545) );
  AND U23417 ( .A(n23551), .B(n23552), .Z(n23550) );
  XNOR U23418 ( .A(p_input[923]), .B(n23549), .Z(n23552) );
  XNOR U23419 ( .A(n23549), .B(n23374), .Z(n23551) );
  IV U23420 ( .A(p_input[907]), .Z(n23374) );
  XOR U23421 ( .A(n23553), .B(n23554), .Z(n23549) );
  AND U23422 ( .A(n23555), .B(n23556), .Z(n23554) );
  XNOR U23423 ( .A(p_input[922]), .B(n23553), .Z(n23556) );
  XNOR U23424 ( .A(n23553), .B(n23383), .Z(n23555) );
  IV U23425 ( .A(p_input[906]), .Z(n23383) );
  XOR U23426 ( .A(n23557), .B(n23558), .Z(n23553) );
  AND U23427 ( .A(n23559), .B(n23560), .Z(n23558) );
  XNOR U23428 ( .A(p_input[921]), .B(n23557), .Z(n23560) );
  XNOR U23429 ( .A(n23557), .B(n23392), .Z(n23559) );
  IV U23430 ( .A(p_input[905]), .Z(n23392) );
  XOR U23431 ( .A(n23561), .B(n23562), .Z(n23557) );
  AND U23432 ( .A(n23563), .B(n23564), .Z(n23562) );
  XNOR U23433 ( .A(p_input[920]), .B(n23561), .Z(n23564) );
  XNOR U23434 ( .A(n23561), .B(n23401), .Z(n23563) );
  IV U23435 ( .A(p_input[904]), .Z(n23401) );
  XOR U23436 ( .A(n23565), .B(n23566), .Z(n23561) );
  AND U23437 ( .A(n23567), .B(n23568), .Z(n23566) );
  XNOR U23438 ( .A(p_input[919]), .B(n23565), .Z(n23568) );
  XNOR U23439 ( .A(n23565), .B(n23410), .Z(n23567) );
  IV U23440 ( .A(p_input[903]), .Z(n23410) );
  XOR U23441 ( .A(n23569), .B(n23570), .Z(n23565) );
  AND U23442 ( .A(n23571), .B(n23572), .Z(n23570) );
  XNOR U23443 ( .A(p_input[918]), .B(n23569), .Z(n23572) );
  XNOR U23444 ( .A(n23569), .B(n23419), .Z(n23571) );
  IV U23445 ( .A(p_input[902]), .Z(n23419) );
  XOR U23446 ( .A(n23573), .B(n23574), .Z(n23569) );
  AND U23447 ( .A(n23575), .B(n23576), .Z(n23574) );
  XNOR U23448 ( .A(p_input[917]), .B(n23573), .Z(n23576) );
  XNOR U23449 ( .A(n23573), .B(n23428), .Z(n23575) );
  IV U23450 ( .A(p_input[901]), .Z(n23428) );
  XOR U23451 ( .A(n23577), .B(n23578), .Z(n23573) );
  AND U23452 ( .A(n23579), .B(n23580), .Z(n23578) );
  XNOR U23453 ( .A(p_input[916]), .B(n23577), .Z(n23580) );
  XNOR U23454 ( .A(n23577), .B(n23437), .Z(n23579) );
  IV U23455 ( .A(p_input[900]), .Z(n23437) );
  XOR U23456 ( .A(n23581), .B(n23582), .Z(n23577) );
  AND U23457 ( .A(n23583), .B(n23584), .Z(n23582) );
  XNOR U23458 ( .A(p_input[915]), .B(n23581), .Z(n23584) );
  XNOR U23459 ( .A(n23581), .B(n23446), .Z(n23583) );
  IV U23460 ( .A(p_input[899]), .Z(n23446) );
  XOR U23461 ( .A(n23585), .B(n23586), .Z(n23581) );
  AND U23462 ( .A(n23587), .B(n23588), .Z(n23586) );
  XNOR U23463 ( .A(p_input[914]), .B(n23585), .Z(n23588) );
  XNOR U23464 ( .A(n23585), .B(n23455), .Z(n23587) );
  IV U23465 ( .A(p_input[898]), .Z(n23455) );
  XNOR U23466 ( .A(n23589), .B(n23590), .Z(n23585) );
  AND U23467 ( .A(n23591), .B(n23592), .Z(n23590) );
  XOR U23468 ( .A(p_input[913]), .B(n23589), .Z(n23592) );
  XNOR U23469 ( .A(p_input[897]), .B(n23589), .Z(n23591) );
  AND U23470 ( .A(p_input[912]), .B(n23593), .Z(n23589) );
  IV U23471 ( .A(p_input[896]), .Z(n23593) );
  XOR U23472 ( .A(n23594), .B(n23595), .Z(n22709) );
  AND U23473 ( .A(n821), .B(n23596), .Z(n23595) );
  XNOR U23474 ( .A(n23597), .B(n23594), .Z(n23596) );
  XOR U23475 ( .A(n23598), .B(n23599), .Z(n821) );
  AND U23476 ( .A(n23600), .B(n23601), .Z(n23599) );
  XNOR U23477 ( .A(n22721), .B(n23598), .Z(n23601) );
  AND U23478 ( .A(n23602), .B(n23603), .Z(n22721) );
  XOR U23479 ( .A(n23598), .B(n22720), .Z(n23600) );
  AND U23480 ( .A(n23604), .B(n23605), .Z(n22720) );
  XOR U23481 ( .A(n23606), .B(n23607), .Z(n23598) );
  AND U23482 ( .A(n23608), .B(n23609), .Z(n23607) );
  XOR U23483 ( .A(n23606), .B(n22733), .Z(n23609) );
  XOR U23484 ( .A(n23610), .B(n23611), .Z(n22733) );
  AND U23485 ( .A(n547), .B(n23612), .Z(n23611) );
  XOR U23486 ( .A(n23613), .B(n23610), .Z(n23612) );
  XNOR U23487 ( .A(n22730), .B(n23606), .Z(n23608) );
  XOR U23488 ( .A(n23614), .B(n23615), .Z(n22730) );
  AND U23489 ( .A(n544), .B(n23616), .Z(n23615) );
  XOR U23490 ( .A(n23617), .B(n23614), .Z(n23616) );
  XOR U23491 ( .A(n23618), .B(n23619), .Z(n23606) );
  AND U23492 ( .A(n23620), .B(n23621), .Z(n23619) );
  XOR U23493 ( .A(n23618), .B(n22745), .Z(n23621) );
  XOR U23494 ( .A(n23622), .B(n23623), .Z(n22745) );
  AND U23495 ( .A(n547), .B(n23624), .Z(n23623) );
  XOR U23496 ( .A(n23625), .B(n23622), .Z(n23624) );
  XNOR U23497 ( .A(n22742), .B(n23618), .Z(n23620) );
  XOR U23498 ( .A(n23626), .B(n23627), .Z(n22742) );
  AND U23499 ( .A(n544), .B(n23628), .Z(n23627) );
  XOR U23500 ( .A(n23629), .B(n23626), .Z(n23628) );
  XOR U23501 ( .A(n23630), .B(n23631), .Z(n23618) );
  AND U23502 ( .A(n23632), .B(n23633), .Z(n23631) );
  XOR U23503 ( .A(n23630), .B(n22757), .Z(n23633) );
  XOR U23504 ( .A(n23634), .B(n23635), .Z(n22757) );
  AND U23505 ( .A(n547), .B(n23636), .Z(n23635) );
  XOR U23506 ( .A(n23637), .B(n23634), .Z(n23636) );
  XNOR U23507 ( .A(n22754), .B(n23630), .Z(n23632) );
  XOR U23508 ( .A(n23638), .B(n23639), .Z(n22754) );
  AND U23509 ( .A(n544), .B(n23640), .Z(n23639) );
  XOR U23510 ( .A(n23641), .B(n23638), .Z(n23640) );
  XOR U23511 ( .A(n23642), .B(n23643), .Z(n23630) );
  AND U23512 ( .A(n23644), .B(n23645), .Z(n23643) );
  XOR U23513 ( .A(n23642), .B(n22769), .Z(n23645) );
  XOR U23514 ( .A(n23646), .B(n23647), .Z(n22769) );
  AND U23515 ( .A(n547), .B(n23648), .Z(n23647) );
  XOR U23516 ( .A(n23649), .B(n23646), .Z(n23648) );
  XNOR U23517 ( .A(n22766), .B(n23642), .Z(n23644) );
  XOR U23518 ( .A(n23650), .B(n23651), .Z(n22766) );
  AND U23519 ( .A(n544), .B(n23652), .Z(n23651) );
  XOR U23520 ( .A(n23653), .B(n23650), .Z(n23652) );
  XOR U23521 ( .A(n23654), .B(n23655), .Z(n23642) );
  AND U23522 ( .A(n23656), .B(n23657), .Z(n23655) );
  XOR U23523 ( .A(n23654), .B(n22781), .Z(n23657) );
  XOR U23524 ( .A(n23658), .B(n23659), .Z(n22781) );
  AND U23525 ( .A(n547), .B(n23660), .Z(n23659) );
  XOR U23526 ( .A(n23661), .B(n23658), .Z(n23660) );
  XNOR U23527 ( .A(n22778), .B(n23654), .Z(n23656) );
  XOR U23528 ( .A(n23662), .B(n23663), .Z(n22778) );
  AND U23529 ( .A(n544), .B(n23664), .Z(n23663) );
  XOR U23530 ( .A(n23665), .B(n23662), .Z(n23664) );
  XOR U23531 ( .A(n23666), .B(n23667), .Z(n23654) );
  AND U23532 ( .A(n23668), .B(n23669), .Z(n23667) );
  XOR U23533 ( .A(n23666), .B(n22793), .Z(n23669) );
  XOR U23534 ( .A(n23670), .B(n23671), .Z(n22793) );
  AND U23535 ( .A(n547), .B(n23672), .Z(n23671) );
  XOR U23536 ( .A(n23673), .B(n23670), .Z(n23672) );
  XNOR U23537 ( .A(n22790), .B(n23666), .Z(n23668) );
  XOR U23538 ( .A(n23674), .B(n23675), .Z(n22790) );
  AND U23539 ( .A(n544), .B(n23676), .Z(n23675) );
  XOR U23540 ( .A(n23677), .B(n23674), .Z(n23676) );
  XOR U23541 ( .A(n23678), .B(n23679), .Z(n23666) );
  AND U23542 ( .A(n23680), .B(n23681), .Z(n23679) );
  XOR U23543 ( .A(n23678), .B(n22805), .Z(n23681) );
  XOR U23544 ( .A(n23682), .B(n23683), .Z(n22805) );
  AND U23545 ( .A(n547), .B(n23684), .Z(n23683) );
  XOR U23546 ( .A(n23685), .B(n23682), .Z(n23684) );
  XNOR U23547 ( .A(n22802), .B(n23678), .Z(n23680) );
  XOR U23548 ( .A(n23686), .B(n23687), .Z(n22802) );
  AND U23549 ( .A(n544), .B(n23688), .Z(n23687) );
  XOR U23550 ( .A(n23689), .B(n23686), .Z(n23688) );
  XOR U23551 ( .A(n23690), .B(n23691), .Z(n23678) );
  AND U23552 ( .A(n23692), .B(n23693), .Z(n23691) );
  XOR U23553 ( .A(n23690), .B(n22817), .Z(n23693) );
  XOR U23554 ( .A(n23694), .B(n23695), .Z(n22817) );
  AND U23555 ( .A(n547), .B(n23696), .Z(n23695) );
  XOR U23556 ( .A(n23697), .B(n23694), .Z(n23696) );
  XNOR U23557 ( .A(n22814), .B(n23690), .Z(n23692) );
  XOR U23558 ( .A(n23698), .B(n23699), .Z(n22814) );
  AND U23559 ( .A(n544), .B(n23700), .Z(n23699) );
  XOR U23560 ( .A(n23701), .B(n23698), .Z(n23700) );
  XOR U23561 ( .A(n23702), .B(n23703), .Z(n23690) );
  AND U23562 ( .A(n23704), .B(n23705), .Z(n23703) );
  XOR U23563 ( .A(n23702), .B(n22829), .Z(n23705) );
  XOR U23564 ( .A(n23706), .B(n23707), .Z(n22829) );
  AND U23565 ( .A(n547), .B(n23708), .Z(n23707) );
  XOR U23566 ( .A(n23709), .B(n23706), .Z(n23708) );
  XNOR U23567 ( .A(n22826), .B(n23702), .Z(n23704) );
  XOR U23568 ( .A(n23710), .B(n23711), .Z(n22826) );
  AND U23569 ( .A(n544), .B(n23712), .Z(n23711) );
  XOR U23570 ( .A(n23713), .B(n23710), .Z(n23712) );
  XOR U23571 ( .A(n23714), .B(n23715), .Z(n23702) );
  AND U23572 ( .A(n23716), .B(n23717), .Z(n23715) );
  XOR U23573 ( .A(n23714), .B(n22841), .Z(n23717) );
  XOR U23574 ( .A(n23718), .B(n23719), .Z(n22841) );
  AND U23575 ( .A(n547), .B(n23720), .Z(n23719) );
  XOR U23576 ( .A(n23721), .B(n23718), .Z(n23720) );
  XNOR U23577 ( .A(n22838), .B(n23714), .Z(n23716) );
  XOR U23578 ( .A(n23722), .B(n23723), .Z(n22838) );
  AND U23579 ( .A(n544), .B(n23724), .Z(n23723) );
  XOR U23580 ( .A(n23725), .B(n23722), .Z(n23724) );
  XOR U23581 ( .A(n23726), .B(n23727), .Z(n23714) );
  AND U23582 ( .A(n23728), .B(n23729), .Z(n23727) );
  XOR U23583 ( .A(n23726), .B(n22853), .Z(n23729) );
  XOR U23584 ( .A(n23730), .B(n23731), .Z(n22853) );
  AND U23585 ( .A(n547), .B(n23732), .Z(n23731) );
  XOR U23586 ( .A(n23733), .B(n23730), .Z(n23732) );
  XNOR U23587 ( .A(n22850), .B(n23726), .Z(n23728) );
  XOR U23588 ( .A(n23734), .B(n23735), .Z(n22850) );
  AND U23589 ( .A(n544), .B(n23736), .Z(n23735) );
  XOR U23590 ( .A(n23737), .B(n23734), .Z(n23736) );
  XOR U23591 ( .A(n23738), .B(n23739), .Z(n23726) );
  AND U23592 ( .A(n23740), .B(n23741), .Z(n23739) );
  XOR U23593 ( .A(n23738), .B(n22865), .Z(n23741) );
  XOR U23594 ( .A(n23742), .B(n23743), .Z(n22865) );
  AND U23595 ( .A(n547), .B(n23744), .Z(n23743) );
  XOR U23596 ( .A(n23745), .B(n23742), .Z(n23744) );
  XNOR U23597 ( .A(n22862), .B(n23738), .Z(n23740) );
  XOR U23598 ( .A(n23746), .B(n23747), .Z(n22862) );
  AND U23599 ( .A(n544), .B(n23748), .Z(n23747) );
  XOR U23600 ( .A(n23749), .B(n23746), .Z(n23748) );
  XOR U23601 ( .A(n23750), .B(n23751), .Z(n23738) );
  AND U23602 ( .A(n23752), .B(n23753), .Z(n23751) );
  XOR U23603 ( .A(n23750), .B(n22877), .Z(n23753) );
  XOR U23604 ( .A(n23754), .B(n23755), .Z(n22877) );
  AND U23605 ( .A(n547), .B(n23756), .Z(n23755) );
  XOR U23606 ( .A(n23757), .B(n23754), .Z(n23756) );
  XNOR U23607 ( .A(n22874), .B(n23750), .Z(n23752) );
  XOR U23608 ( .A(n23758), .B(n23759), .Z(n22874) );
  AND U23609 ( .A(n544), .B(n23760), .Z(n23759) );
  XOR U23610 ( .A(n23761), .B(n23758), .Z(n23760) );
  XOR U23611 ( .A(n23762), .B(n23763), .Z(n23750) );
  AND U23612 ( .A(n23764), .B(n23765), .Z(n23763) );
  XNOR U23613 ( .A(n23766), .B(n22890), .Z(n23765) );
  XOR U23614 ( .A(n23767), .B(n23768), .Z(n22890) );
  AND U23615 ( .A(n547), .B(n23769), .Z(n23768) );
  XOR U23616 ( .A(n23767), .B(n23770), .Z(n23769) );
  XNOR U23617 ( .A(n22887), .B(n23762), .Z(n23764) );
  XOR U23618 ( .A(n23771), .B(n23772), .Z(n22887) );
  AND U23619 ( .A(n544), .B(n23773), .Z(n23772) );
  XOR U23620 ( .A(n23771), .B(n23774), .Z(n23773) );
  IV U23621 ( .A(n23766), .Z(n23762) );
  AND U23622 ( .A(n23594), .B(n23597), .Z(n23766) );
  XNOR U23623 ( .A(n23775), .B(n23776), .Z(n23597) );
  AND U23624 ( .A(n547), .B(n23777), .Z(n23776) );
  XNOR U23625 ( .A(n23778), .B(n23775), .Z(n23777) );
  XOR U23626 ( .A(n23779), .B(n23780), .Z(n547) );
  AND U23627 ( .A(n23781), .B(n23782), .Z(n23780) );
  XNOR U23628 ( .A(n23602), .B(n23779), .Z(n23782) );
  AND U23629 ( .A(p_input[895]), .B(p_input[879]), .Z(n23602) );
  XOR U23630 ( .A(n23779), .B(n23603), .Z(n23781) );
  AND U23631 ( .A(p_input[863]), .B(p_input[847]), .Z(n23603) );
  XOR U23632 ( .A(n23783), .B(n23784), .Z(n23779) );
  AND U23633 ( .A(n23785), .B(n23786), .Z(n23784) );
  XOR U23634 ( .A(n23783), .B(n23613), .Z(n23786) );
  XNOR U23635 ( .A(p_input[878]), .B(n23787), .Z(n23613) );
  AND U23636 ( .A(n871), .B(n23788), .Z(n23787) );
  XOR U23637 ( .A(p_input[894]), .B(p_input[878]), .Z(n23788) );
  XNOR U23638 ( .A(n23610), .B(n23783), .Z(n23785) );
  XOR U23639 ( .A(n23789), .B(n23790), .Z(n23610) );
  AND U23640 ( .A(n869), .B(n23791), .Z(n23790) );
  XOR U23641 ( .A(p_input[862]), .B(p_input[846]), .Z(n23791) );
  XOR U23642 ( .A(n23792), .B(n23793), .Z(n23783) );
  AND U23643 ( .A(n23794), .B(n23795), .Z(n23793) );
  XOR U23644 ( .A(n23792), .B(n23625), .Z(n23795) );
  XNOR U23645 ( .A(p_input[877]), .B(n23796), .Z(n23625) );
  AND U23646 ( .A(n871), .B(n23797), .Z(n23796) );
  XOR U23647 ( .A(p_input[893]), .B(p_input[877]), .Z(n23797) );
  XNOR U23648 ( .A(n23622), .B(n23792), .Z(n23794) );
  XOR U23649 ( .A(n23798), .B(n23799), .Z(n23622) );
  AND U23650 ( .A(n869), .B(n23800), .Z(n23799) );
  XOR U23651 ( .A(p_input[861]), .B(p_input[845]), .Z(n23800) );
  XOR U23652 ( .A(n23801), .B(n23802), .Z(n23792) );
  AND U23653 ( .A(n23803), .B(n23804), .Z(n23802) );
  XOR U23654 ( .A(n23801), .B(n23637), .Z(n23804) );
  XNOR U23655 ( .A(p_input[876]), .B(n23805), .Z(n23637) );
  AND U23656 ( .A(n871), .B(n23806), .Z(n23805) );
  XOR U23657 ( .A(p_input[892]), .B(p_input[876]), .Z(n23806) );
  XNOR U23658 ( .A(n23634), .B(n23801), .Z(n23803) );
  XOR U23659 ( .A(n23807), .B(n23808), .Z(n23634) );
  AND U23660 ( .A(n869), .B(n23809), .Z(n23808) );
  XOR U23661 ( .A(p_input[860]), .B(p_input[844]), .Z(n23809) );
  XOR U23662 ( .A(n23810), .B(n23811), .Z(n23801) );
  AND U23663 ( .A(n23812), .B(n23813), .Z(n23811) );
  XOR U23664 ( .A(n23810), .B(n23649), .Z(n23813) );
  XNOR U23665 ( .A(p_input[875]), .B(n23814), .Z(n23649) );
  AND U23666 ( .A(n871), .B(n23815), .Z(n23814) );
  XOR U23667 ( .A(p_input[891]), .B(p_input[875]), .Z(n23815) );
  XNOR U23668 ( .A(n23646), .B(n23810), .Z(n23812) );
  XOR U23669 ( .A(n23816), .B(n23817), .Z(n23646) );
  AND U23670 ( .A(n869), .B(n23818), .Z(n23817) );
  XOR U23671 ( .A(p_input[859]), .B(p_input[843]), .Z(n23818) );
  XOR U23672 ( .A(n23819), .B(n23820), .Z(n23810) );
  AND U23673 ( .A(n23821), .B(n23822), .Z(n23820) );
  XOR U23674 ( .A(n23819), .B(n23661), .Z(n23822) );
  XNOR U23675 ( .A(p_input[874]), .B(n23823), .Z(n23661) );
  AND U23676 ( .A(n871), .B(n23824), .Z(n23823) );
  XOR U23677 ( .A(p_input[890]), .B(p_input[874]), .Z(n23824) );
  XNOR U23678 ( .A(n23658), .B(n23819), .Z(n23821) );
  XOR U23679 ( .A(n23825), .B(n23826), .Z(n23658) );
  AND U23680 ( .A(n869), .B(n23827), .Z(n23826) );
  XOR U23681 ( .A(p_input[858]), .B(p_input[842]), .Z(n23827) );
  XOR U23682 ( .A(n23828), .B(n23829), .Z(n23819) );
  AND U23683 ( .A(n23830), .B(n23831), .Z(n23829) );
  XOR U23684 ( .A(n23828), .B(n23673), .Z(n23831) );
  XNOR U23685 ( .A(p_input[873]), .B(n23832), .Z(n23673) );
  AND U23686 ( .A(n871), .B(n23833), .Z(n23832) );
  XOR U23687 ( .A(p_input[889]), .B(p_input[873]), .Z(n23833) );
  XNOR U23688 ( .A(n23670), .B(n23828), .Z(n23830) );
  XOR U23689 ( .A(n23834), .B(n23835), .Z(n23670) );
  AND U23690 ( .A(n869), .B(n23836), .Z(n23835) );
  XOR U23691 ( .A(p_input[857]), .B(p_input[841]), .Z(n23836) );
  XOR U23692 ( .A(n23837), .B(n23838), .Z(n23828) );
  AND U23693 ( .A(n23839), .B(n23840), .Z(n23838) );
  XOR U23694 ( .A(n23837), .B(n23685), .Z(n23840) );
  XNOR U23695 ( .A(p_input[872]), .B(n23841), .Z(n23685) );
  AND U23696 ( .A(n871), .B(n23842), .Z(n23841) );
  XOR U23697 ( .A(p_input[888]), .B(p_input[872]), .Z(n23842) );
  XNOR U23698 ( .A(n23682), .B(n23837), .Z(n23839) );
  XOR U23699 ( .A(n23843), .B(n23844), .Z(n23682) );
  AND U23700 ( .A(n869), .B(n23845), .Z(n23844) );
  XOR U23701 ( .A(p_input[856]), .B(p_input[840]), .Z(n23845) );
  XOR U23702 ( .A(n23846), .B(n23847), .Z(n23837) );
  AND U23703 ( .A(n23848), .B(n23849), .Z(n23847) );
  XOR U23704 ( .A(n23846), .B(n23697), .Z(n23849) );
  XNOR U23705 ( .A(p_input[871]), .B(n23850), .Z(n23697) );
  AND U23706 ( .A(n871), .B(n23851), .Z(n23850) );
  XOR U23707 ( .A(p_input[887]), .B(p_input[871]), .Z(n23851) );
  XNOR U23708 ( .A(n23694), .B(n23846), .Z(n23848) );
  XOR U23709 ( .A(n23852), .B(n23853), .Z(n23694) );
  AND U23710 ( .A(n869), .B(n23854), .Z(n23853) );
  XOR U23711 ( .A(p_input[855]), .B(p_input[839]), .Z(n23854) );
  XOR U23712 ( .A(n23855), .B(n23856), .Z(n23846) );
  AND U23713 ( .A(n23857), .B(n23858), .Z(n23856) );
  XOR U23714 ( .A(n23855), .B(n23709), .Z(n23858) );
  XNOR U23715 ( .A(p_input[870]), .B(n23859), .Z(n23709) );
  AND U23716 ( .A(n871), .B(n23860), .Z(n23859) );
  XOR U23717 ( .A(p_input[886]), .B(p_input[870]), .Z(n23860) );
  XNOR U23718 ( .A(n23706), .B(n23855), .Z(n23857) );
  XOR U23719 ( .A(n23861), .B(n23862), .Z(n23706) );
  AND U23720 ( .A(n869), .B(n23863), .Z(n23862) );
  XOR U23721 ( .A(p_input[854]), .B(p_input[838]), .Z(n23863) );
  XOR U23722 ( .A(n23864), .B(n23865), .Z(n23855) );
  AND U23723 ( .A(n23866), .B(n23867), .Z(n23865) );
  XOR U23724 ( .A(n23864), .B(n23721), .Z(n23867) );
  XNOR U23725 ( .A(p_input[869]), .B(n23868), .Z(n23721) );
  AND U23726 ( .A(n871), .B(n23869), .Z(n23868) );
  XOR U23727 ( .A(p_input[885]), .B(p_input[869]), .Z(n23869) );
  XNOR U23728 ( .A(n23718), .B(n23864), .Z(n23866) );
  XOR U23729 ( .A(n23870), .B(n23871), .Z(n23718) );
  AND U23730 ( .A(n869), .B(n23872), .Z(n23871) );
  XOR U23731 ( .A(p_input[853]), .B(p_input[837]), .Z(n23872) );
  XOR U23732 ( .A(n23873), .B(n23874), .Z(n23864) );
  AND U23733 ( .A(n23875), .B(n23876), .Z(n23874) );
  XOR U23734 ( .A(n23873), .B(n23733), .Z(n23876) );
  XNOR U23735 ( .A(p_input[868]), .B(n23877), .Z(n23733) );
  AND U23736 ( .A(n871), .B(n23878), .Z(n23877) );
  XOR U23737 ( .A(p_input[884]), .B(p_input[868]), .Z(n23878) );
  XNOR U23738 ( .A(n23730), .B(n23873), .Z(n23875) );
  XOR U23739 ( .A(n23879), .B(n23880), .Z(n23730) );
  AND U23740 ( .A(n869), .B(n23881), .Z(n23880) );
  XOR U23741 ( .A(p_input[852]), .B(p_input[836]), .Z(n23881) );
  XOR U23742 ( .A(n23882), .B(n23883), .Z(n23873) );
  AND U23743 ( .A(n23884), .B(n23885), .Z(n23883) );
  XOR U23744 ( .A(n23882), .B(n23745), .Z(n23885) );
  XNOR U23745 ( .A(p_input[867]), .B(n23886), .Z(n23745) );
  AND U23746 ( .A(n871), .B(n23887), .Z(n23886) );
  XOR U23747 ( .A(p_input[883]), .B(p_input[867]), .Z(n23887) );
  XNOR U23748 ( .A(n23742), .B(n23882), .Z(n23884) );
  XOR U23749 ( .A(n23888), .B(n23889), .Z(n23742) );
  AND U23750 ( .A(n869), .B(n23890), .Z(n23889) );
  XOR U23751 ( .A(p_input[851]), .B(p_input[835]), .Z(n23890) );
  XOR U23752 ( .A(n23891), .B(n23892), .Z(n23882) );
  AND U23753 ( .A(n23893), .B(n23894), .Z(n23892) );
  XOR U23754 ( .A(n23891), .B(n23757), .Z(n23894) );
  XNOR U23755 ( .A(p_input[866]), .B(n23895), .Z(n23757) );
  AND U23756 ( .A(n871), .B(n23896), .Z(n23895) );
  XOR U23757 ( .A(p_input[882]), .B(p_input[866]), .Z(n23896) );
  XNOR U23758 ( .A(n23754), .B(n23891), .Z(n23893) );
  XOR U23759 ( .A(n23897), .B(n23898), .Z(n23754) );
  AND U23760 ( .A(n869), .B(n23899), .Z(n23898) );
  XOR U23761 ( .A(p_input[850]), .B(p_input[834]), .Z(n23899) );
  XOR U23762 ( .A(n23900), .B(n23901), .Z(n23891) );
  AND U23763 ( .A(n23902), .B(n23903), .Z(n23901) );
  XNOR U23764 ( .A(n23904), .B(n23770), .Z(n23903) );
  XNOR U23765 ( .A(p_input[865]), .B(n23905), .Z(n23770) );
  AND U23766 ( .A(n871), .B(n23906), .Z(n23905) );
  XNOR U23767 ( .A(p_input[881]), .B(n23907), .Z(n23906) );
  IV U23768 ( .A(p_input[865]), .Z(n23907) );
  XNOR U23769 ( .A(n23767), .B(n23900), .Z(n23902) );
  XNOR U23770 ( .A(p_input[833]), .B(n23908), .Z(n23767) );
  AND U23771 ( .A(n869), .B(n23909), .Z(n23908) );
  XOR U23772 ( .A(p_input[849]), .B(p_input[833]), .Z(n23909) );
  IV U23773 ( .A(n23904), .Z(n23900) );
  AND U23774 ( .A(n23775), .B(n23778), .Z(n23904) );
  XOR U23775 ( .A(p_input[864]), .B(n23910), .Z(n23778) );
  AND U23776 ( .A(n871), .B(n23911), .Z(n23910) );
  XOR U23777 ( .A(p_input[880]), .B(p_input[864]), .Z(n23911) );
  XOR U23778 ( .A(n23912), .B(n23913), .Z(n871) );
  AND U23779 ( .A(n23914), .B(n23915), .Z(n23913) );
  XNOR U23780 ( .A(p_input[895]), .B(n23912), .Z(n23915) );
  XOR U23781 ( .A(n23912), .B(p_input[879]), .Z(n23914) );
  XOR U23782 ( .A(n23916), .B(n23917), .Z(n23912) );
  AND U23783 ( .A(n23918), .B(n23919), .Z(n23917) );
  XNOR U23784 ( .A(p_input[894]), .B(n23916), .Z(n23919) );
  XOR U23785 ( .A(n23916), .B(p_input[878]), .Z(n23918) );
  XOR U23786 ( .A(n23920), .B(n23921), .Z(n23916) );
  AND U23787 ( .A(n23922), .B(n23923), .Z(n23921) );
  XNOR U23788 ( .A(p_input[893]), .B(n23920), .Z(n23923) );
  XOR U23789 ( .A(n23920), .B(p_input[877]), .Z(n23922) );
  XOR U23790 ( .A(n23924), .B(n23925), .Z(n23920) );
  AND U23791 ( .A(n23926), .B(n23927), .Z(n23925) );
  XNOR U23792 ( .A(p_input[892]), .B(n23924), .Z(n23927) );
  XOR U23793 ( .A(n23924), .B(p_input[876]), .Z(n23926) );
  XOR U23794 ( .A(n23928), .B(n23929), .Z(n23924) );
  AND U23795 ( .A(n23930), .B(n23931), .Z(n23929) );
  XNOR U23796 ( .A(p_input[891]), .B(n23928), .Z(n23931) );
  XOR U23797 ( .A(n23928), .B(p_input[875]), .Z(n23930) );
  XOR U23798 ( .A(n23932), .B(n23933), .Z(n23928) );
  AND U23799 ( .A(n23934), .B(n23935), .Z(n23933) );
  XNOR U23800 ( .A(p_input[890]), .B(n23932), .Z(n23935) );
  XOR U23801 ( .A(n23932), .B(p_input[874]), .Z(n23934) );
  XOR U23802 ( .A(n23936), .B(n23937), .Z(n23932) );
  AND U23803 ( .A(n23938), .B(n23939), .Z(n23937) );
  XNOR U23804 ( .A(p_input[889]), .B(n23936), .Z(n23939) );
  XOR U23805 ( .A(n23936), .B(p_input[873]), .Z(n23938) );
  XOR U23806 ( .A(n23940), .B(n23941), .Z(n23936) );
  AND U23807 ( .A(n23942), .B(n23943), .Z(n23941) );
  XNOR U23808 ( .A(p_input[888]), .B(n23940), .Z(n23943) );
  XOR U23809 ( .A(n23940), .B(p_input[872]), .Z(n23942) );
  XOR U23810 ( .A(n23944), .B(n23945), .Z(n23940) );
  AND U23811 ( .A(n23946), .B(n23947), .Z(n23945) );
  XNOR U23812 ( .A(p_input[887]), .B(n23944), .Z(n23947) );
  XOR U23813 ( .A(n23944), .B(p_input[871]), .Z(n23946) );
  XOR U23814 ( .A(n23948), .B(n23949), .Z(n23944) );
  AND U23815 ( .A(n23950), .B(n23951), .Z(n23949) );
  XNOR U23816 ( .A(p_input[886]), .B(n23948), .Z(n23951) );
  XOR U23817 ( .A(n23948), .B(p_input[870]), .Z(n23950) );
  XOR U23818 ( .A(n23952), .B(n23953), .Z(n23948) );
  AND U23819 ( .A(n23954), .B(n23955), .Z(n23953) );
  XNOR U23820 ( .A(p_input[885]), .B(n23952), .Z(n23955) );
  XOR U23821 ( .A(n23952), .B(p_input[869]), .Z(n23954) );
  XOR U23822 ( .A(n23956), .B(n23957), .Z(n23952) );
  AND U23823 ( .A(n23958), .B(n23959), .Z(n23957) );
  XNOR U23824 ( .A(p_input[884]), .B(n23956), .Z(n23959) );
  XOR U23825 ( .A(n23956), .B(p_input[868]), .Z(n23958) );
  XOR U23826 ( .A(n23960), .B(n23961), .Z(n23956) );
  AND U23827 ( .A(n23962), .B(n23963), .Z(n23961) );
  XNOR U23828 ( .A(p_input[883]), .B(n23960), .Z(n23963) );
  XOR U23829 ( .A(n23960), .B(p_input[867]), .Z(n23962) );
  XOR U23830 ( .A(n23964), .B(n23965), .Z(n23960) );
  AND U23831 ( .A(n23966), .B(n23967), .Z(n23965) );
  XNOR U23832 ( .A(p_input[882]), .B(n23964), .Z(n23967) );
  XOR U23833 ( .A(n23964), .B(p_input[866]), .Z(n23966) );
  XNOR U23834 ( .A(n23968), .B(n23969), .Z(n23964) );
  AND U23835 ( .A(n23970), .B(n23971), .Z(n23969) );
  XOR U23836 ( .A(p_input[881]), .B(n23968), .Z(n23971) );
  XNOR U23837 ( .A(p_input[865]), .B(n23968), .Z(n23970) );
  AND U23838 ( .A(p_input[880]), .B(n23972), .Z(n23968) );
  IV U23839 ( .A(p_input[864]), .Z(n23972) );
  XNOR U23840 ( .A(p_input[832]), .B(n23973), .Z(n23775) );
  AND U23841 ( .A(n869), .B(n23974), .Z(n23973) );
  XOR U23842 ( .A(p_input[848]), .B(p_input[832]), .Z(n23974) );
  XOR U23843 ( .A(n23975), .B(n23976), .Z(n869) );
  AND U23844 ( .A(n23977), .B(n23978), .Z(n23976) );
  XNOR U23845 ( .A(p_input[863]), .B(n23975), .Z(n23978) );
  XOR U23846 ( .A(n23975), .B(p_input[847]), .Z(n23977) );
  XOR U23847 ( .A(n23979), .B(n23980), .Z(n23975) );
  AND U23848 ( .A(n23981), .B(n23982), .Z(n23980) );
  XNOR U23849 ( .A(p_input[862]), .B(n23979), .Z(n23982) );
  XNOR U23850 ( .A(n23979), .B(n23789), .Z(n23981) );
  IV U23851 ( .A(p_input[846]), .Z(n23789) );
  XOR U23852 ( .A(n23983), .B(n23984), .Z(n23979) );
  AND U23853 ( .A(n23985), .B(n23986), .Z(n23984) );
  XNOR U23854 ( .A(p_input[861]), .B(n23983), .Z(n23986) );
  XNOR U23855 ( .A(n23983), .B(n23798), .Z(n23985) );
  IV U23856 ( .A(p_input[845]), .Z(n23798) );
  XOR U23857 ( .A(n23987), .B(n23988), .Z(n23983) );
  AND U23858 ( .A(n23989), .B(n23990), .Z(n23988) );
  XNOR U23859 ( .A(p_input[860]), .B(n23987), .Z(n23990) );
  XNOR U23860 ( .A(n23987), .B(n23807), .Z(n23989) );
  IV U23861 ( .A(p_input[844]), .Z(n23807) );
  XOR U23862 ( .A(n23991), .B(n23992), .Z(n23987) );
  AND U23863 ( .A(n23993), .B(n23994), .Z(n23992) );
  XNOR U23864 ( .A(p_input[859]), .B(n23991), .Z(n23994) );
  XNOR U23865 ( .A(n23991), .B(n23816), .Z(n23993) );
  IV U23866 ( .A(p_input[843]), .Z(n23816) );
  XOR U23867 ( .A(n23995), .B(n23996), .Z(n23991) );
  AND U23868 ( .A(n23997), .B(n23998), .Z(n23996) );
  XNOR U23869 ( .A(p_input[858]), .B(n23995), .Z(n23998) );
  XNOR U23870 ( .A(n23995), .B(n23825), .Z(n23997) );
  IV U23871 ( .A(p_input[842]), .Z(n23825) );
  XOR U23872 ( .A(n23999), .B(n24000), .Z(n23995) );
  AND U23873 ( .A(n24001), .B(n24002), .Z(n24000) );
  XNOR U23874 ( .A(p_input[857]), .B(n23999), .Z(n24002) );
  XNOR U23875 ( .A(n23999), .B(n23834), .Z(n24001) );
  IV U23876 ( .A(p_input[841]), .Z(n23834) );
  XOR U23877 ( .A(n24003), .B(n24004), .Z(n23999) );
  AND U23878 ( .A(n24005), .B(n24006), .Z(n24004) );
  XNOR U23879 ( .A(p_input[856]), .B(n24003), .Z(n24006) );
  XNOR U23880 ( .A(n24003), .B(n23843), .Z(n24005) );
  IV U23881 ( .A(p_input[840]), .Z(n23843) );
  XOR U23882 ( .A(n24007), .B(n24008), .Z(n24003) );
  AND U23883 ( .A(n24009), .B(n24010), .Z(n24008) );
  XNOR U23884 ( .A(p_input[855]), .B(n24007), .Z(n24010) );
  XNOR U23885 ( .A(n24007), .B(n23852), .Z(n24009) );
  IV U23886 ( .A(p_input[839]), .Z(n23852) );
  XOR U23887 ( .A(n24011), .B(n24012), .Z(n24007) );
  AND U23888 ( .A(n24013), .B(n24014), .Z(n24012) );
  XNOR U23889 ( .A(p_input[854]), .B(n24011), .Z(n24014) );
  XNOR U23890 ( .A(n24011), .B(n23861), .Z(n24013) );
  IV U23891 ( .A(p_input[838]), .Z(n23861) );
  XOR U23892 ( .A(n24015), .B(n24016), .Z(n24011) );
  AND U23893 ( .A(n24017), .B(n24018), .Z(n24016) );
  XNOR U23894 ( .A(p_input[853]), .B(n24015), .Z(n24018) );
  XNOR U23895 ( .A(n24015), .B(n23870), .Z(n24017) );
  IV U23896 ( .A(p_input[837]), .Z(n23870) );
  XOR U23897 ( .A(n24019), .B(n24020), .Z(n24015) );
  AND U23898 ( .A(n24021), .B(n24022), .Z(n24020) );
  XNOR U23899 ( .A(p_input[852]), .B(n24019), .Z(n24022) );
  XNOR U23900 ( .A(n24019), .B(n23879), .Z(n24021) );
  IV U23901 ( .A(p_input[836]), .Z(n23879) );
  XOR U23902 ( .A(n24023), .B(n24024), .Z(n24019) );
  AND U23903 ( .A(n24025), .B(n24026), .Z(n24024) );
  XNOR U23904 ( .A(p_input[851]), .B(n24023), .Z(n24026) );
  XNOR U23905 ( .A(n24023), .B(n23888), .Z(n24025) );
  IV U23906 ( .A(p_input[835]), .Z(n23888) );
  XOR U23907 ( .A(n24027), .B(n24028), .Z(n24023) );
  AND U23908 ( .A(n24029), .B(n24030), .Z(n24028) );
  XNOR U23909 ( .A(p_input[850]), .B(n24027), .Z(n24030) );
  XNOR U23910 ( .A(n24027), .B(n23897), .Z(n24029) );
  IV U23911 ( .A(p_input[834]), .Z(n23897) );
  XNOR U23912 ( .A(n24031), .B(n24032), .Z(n24027) );
  AND U23913 ( .A(n24033), .B(n24034), .Z(n24032) );
  XOR U23914 ( .A(p_input[849]), .B(n24031), .Z(n24034) );
  XNOR U23915 ( .A(p_input[833]), .B(n24031), .Z(n24033) );
  AND U23916 ( .A(p_input[848]), .B(n24035), .Z(n24031) );
  IV U23917 ( .A(p_input[832]), .Z(n24035) );
  XOR U23918 ( .A(n24036), .B(n24037), .Z(n23594) );
  AND U23919 ( .A(n544), .B(n24038), .Z(n24037) );
  XNOR U23920 ( .A(n24039), .B(n24036), .Z(n24038) );
  XOR U23921 ( .A(n24040), .B(n24041), .Z(n544) );
  AND U23922 ( .A(n24042), .B(n24043), .Z(n24041) );
  XNOR U23923 ( .A(n23605), .B(n24040), .Z(n24043) );
  AND U23924 ( .A(p_input[831]), .B(p_input[815]), .Z(n23605) );
  XOR U23925 ( .A(n24040), .B(n23604), .Z(n24042) );
  AND U23926 ( .A(p_input[783]), .B(p_input[799]), .Z(n23604) );
  XOR U23927 ( .A(n24044), .B(n24045), .Z(n24040) );
  AND U23928 ( .A(n24046), .B(n24047), .Z(n24045) );
  XOR U23929 ( .A(n24044), .B(n23617), .Z(n24047) );
  XNOR U23930 ( .A(p_input[814]), .B(n24048), .Z(n23617) );
  AND U23931 ( .A(n875), .B(n24049), .Z(n24048) );
  XOR U23932 ( .A(p_input[830]), .B(p_input[814]), .Z(n24049) );
  XNOR U23933 ( .A(n23614), .B(n24044), .Z(n24046) );
  XOR U23934 ( .A(n24050), .B(n24051), .Z(n23614) );
  AND U23935 ( .A(n872), .B(n24052), .Z(n24051) );
  XOR U23936 ( .A(p_input[798]), .B(p_input[782]), .Z(n24052) );
  XOR U23937 ( .A(n24053), .B(n24054), .Z(n24044) );
  AND U23938 ( .A(n24055), .B(n24056), .Z(n24054) );
  XOR U23939 ( .A(n24053), .B(n23629), .Z(n24056) );
  XNOR U23940 ( .A(p_input[813]), .B(n24057), .Z(n23629) );
  AND U23941 ( .A(n875), .B(n24058), .Z(n24057) );
  XOR U23942 ( .A(p_input[829]), .B(p_input[813]), .Z(n24058) );
  XNOR U23943 ( .A(n23626), .B(n24053), .Z(n24055) );
  XOR U23944 ( .A(n24059), .B(n24060), .Z(n23626) );
  AND U23945 ( .A(n872), .B(n24061), .Z(n24060) );
  XOR U23946 ( .A(p_input[797]), .B(p_input[781]), .Z(n24061) );
  XOR U23947 ( .A(n24062), .B(n24063), .Z(n24053) );
  AND U23948 ( .A(n24064), .B(n24065), .Z(n24063) );
  XOR U23949 ( .A(n24062), .B(n23641), .Z(n24065) );
  XNOR U23950 ( .A(p_input[812]), .B(n24066), .Z(n23641) );
  AND U23951 ( .A(n875), .B(n24067), .Z(n24066) );
  XOR U23952 ( .A(p_input[828]), .B(p_input[812]), .Z(n24067) );
  XNOR U23953 ( .A(n23638), .B(n24062), .Z(n24064) );
  XOR U23954 ( .A(n24068), .B(n24069), .Z(n23638) );
  AND U23955 ( .A(n872), .B(n24070), .Z(n24069) );
  XOR U23956 ( .A(p_input[796]), .B(p_input[780]), .Z(n24070) );
  XOR U23957 ( .A(n24071), .B(n24072), .Z(n24062) );
  AND U23958 ( .A(n24073), .B(n24074), .Z(n24072) );
  XOR U23959 ( .A(n24071), .B(n23653), .Z(n24074) );
  XNOR U23960 ( .A(p_input[811]), .B(n24075), .Z(n23653) );
  AND U23961 ( .A(n875), .B(n24076), .Z(n24075) );
  XOR U23962 ( .A(p_input[827]), .B(p_input[811]), .Z(n24076) );
  XNOR U23963 ( .A(n23650), .B(n24071), .Z(n24073) );
  XOR U23964 ( .A(n24077), .B(n24078), .Z(n23650) );
  AND U23965 ( .A(n872), .B(n24079), .Z(n24078) );
  XOR U23966 ( .A(p_input[795]), .B(p_input[779]), .Z(n24079) );
  XOR U23967 ( .A(n24080), .B(n24081), .Z(n24071) );
  AND U23968 ( .A(n24082), .B(n24083), .Z(n24081) );
  XOR U23969 ( .A(n24080), .B(n23665), .Z(n24083) );
  XNOR U23970 ( .A(p_input[810]), .B(n24084), .Z(n23665) );
  AND U23971 ( .A(n875), .B(n24085), .Z(n24084) );
  XOR U23972 ( .A(p_input[826]), .B(p_input[810]), .Z(n24085) );
  XNOR U23973 ( .A(n23662), .B(n24080), .Z(n24082) );
  XOR U23974 ( .A(n24086), .B(n24087), .Z(n23662) );
  AND U23975 ( .A(n872), .B(n24088), .Z(n24087) );
  XOR U23976 ( .A(p_input[794]), .B(p_input[778]), .Z(n24088) );
  XOR U23977 ( .A(n24089), .B(n24090), .Z(n24080) );
  AND U23978 ( .A(n24091), .B(n24092), .Z(n24090) );
  XOR U23979 ( .A(n24089), .B(n23677), .Z(n24092) );
  XNOR U23980 ( .A(p_input[809]), .B(n24093), .Z(n23677) );
  AND U23981 ( .A(n875), .B(n24094), .Z(n24093) );
  XOR U23982 ( .A(p_input[825]), .B(p_input[809]), .Z(n24094) );
  XNOR U23983 ( .A(n23674), .B(n24089), .Z(n24091) );
  XOR U23984 ( .A(n24095), .B(n24096), .Z(n23674) );
  AND U23985 ( .A(n872), .B(n24097), .Z(n24096) );
  XOR U23986 ( .A(p_input[793]), .B(p_input[777]), .Z(n24097) );
  XOR U23987 ( .A(n24098), .B(n24099), .Z(n24089) );
  AND U23988 ( .A(n24100), .B(n24101), .Z(n24099) );
  XOR U23989 ( .A(n24098), .B(n23689), .Z(n24101) );
  XNOR U23990 ( .A(p_input[808]), .B(n24102), .Z(n23689) );
  AND U23991 ( .A(n875), .B(n24103), .Z(n24102) );
  XOR U23992 ( .A(p_input[824]), .B(p_input[808]), .Z(n24103) );
  XNOR U23993 ( .A(n23686), .B(n24098), .Z(n24100) );
  XOR U23994 ( .A(n24104), .B(n24105), .Z(n23686) );
  AND U23995 ( .A(n872), .B(n24106), .Z(n24105) );
  XOR U23996 ( .A(p_input[792]), .B(p_input[776]), .Z(n24106) );
  XOR U23997 ( .A(n24107), .B(n24108), .Z(n24098) );
  AND U23998 ( .A(n24109), .B(n24110), .Z(n24108) );
  XOR U23999 ( .A(n24107), .B(n23701), .Z(n24110) );
  XNOR U24000 ( .A(p_input[807]), .B(n24111), .Z(n23701) );
  AND U24001 ( .A(n875), .B(n24112), .Z(n24111) );
  XOR U24002 ( .A(p_input[823]), .B(p_input[807]), .Z(n24112) );
  XNOR U24003 ( .A(n23698), .B(n24107), .Z(n24109) );
  XOR U24004 ( .A(n24113), .B(n24114), .Z(n23698) );
  AND U24005 ( .A(n872), .B(n24115), .Z(n24114) );
  XOR U24006 ( .A(p_input[791]), .B(p_input[775]), .Z(n24115) );
  XOR U24007 ( .A(n24116), .B(n24117), .Z(n24107) );
  AND U24008 ( .A(n24118), .B(n24119), .Z(n24117) );
  XOR U24009 ( .A(n24116), .B(n23713), .Z(n24119) );
  XNOR U24010 ( .A(p_input[806]), .B(n24120), .Z(n23713) );
  AND U24011 ( .A(n875), .B(n24121), .Z(n24120) );
  XOR U24012 ( .A(p_input[822]), .B(p_input[806]), .Z(n24121) );
  XNOR U24013 ( .A(n23710), .B(n24116), .Z(n24118) );
  XOR U24014 ( .A(n24122), .B(n24123), .Z(n23710) );
  AND U24015 ( .A(n872), .B(n24124), .Z(n24123) );
  XOR U24016 ( .A(p_input[790]), .B(p_input[774]), .Z(n24124) );
  XOR U24017 ( .A(n24125), .B(n24126), .Z(n24116) );
  AND U24018 ( .A(n24127), .B(n24128), .Z(n24126) );
  XOR U24019 ( .A(n24125), .B(n23725), .Z(n24128) );
  XNOR U24020 ( .A(p_input[805]), .B(n24129), .Z(n23725) );
  AND U24021 ( .A(n875), .B(n24130), .Z(n24129) );
  XOR U24022 ( .A(p_input[821]), .B(p_input[805]), .Z(n24130) );
  XNOR U24023 ( .A(n23722), .B(n24125), .Z(n24127) );
  XOR U24024 ( .A(n24131), .B(n24132), .Z(n23722) );
  AND U24025 ( .A(n872), .B(n24133), .Z(n24132) );
  XOR U24026 ( .A(p_input[789]), .B(p_input[773]), .Z(n24133) );
  XOR U24027 ( .A(n24134), .B(n24135), .Z(n24125) );
  AND U24028 ( .A(n24136), .B(n24137), .Z(n24135) );
  XOR U24029 ( .A(n24134), .B(n23737), .Z(n24137) );
  XNOR U24030 ( .A(p_input[804]), .B(n24138), .Z(n23737) );
  AND U24031 ( .A(n875), .B(n24139), .Z(n24138) );
  XOR U24032 ( .A(p_input[820]), .B(p_input[804]), .Z(n24139) );
  XNOR U24033 ( .A(n23734), .B(n24134), .Z(n24136) );
  XOR U24034 ( .A(n24140), .B(n24141), .Z(n23734) );
  AND U24035 ( .A(n872), .B(n24142), .Z(n24141) );
  XOR U24036 ( .A(p_input[788]), .B(p_input[772]), .Z(n24142) );
  XOR U24037 ( .A(n24143), .B(n24144), .Z(n24134) );
  AND U24038 ( .A(n24145), .B(n24146), .Z(n24144) );
  XOR U24039 ( .A(n24143), .B(n23749), .Z(n24146) );
  XNOR U24040 ( .A(p_input[803]), .B(n24147), .Z(n23749) );
  AND U24041 ( .A(n875), .B(n24148), .Z(n24147) );
  XOR U24042 ( .A(p_input[819]), .B(p_input[803]), .Z(n24148) );
  XNOR U24043 ( .A(n23746), .B(n24143), .Z(n24145) );
  XOR U24044 ( .A(n24149), .B(n24150), .Z(n23746) );
  AND U24045 ( .A(n872), .B(n24151), .Z(n24150) );
  XOR U24046 ( .A(p_input[787]), .B(p_input[771]), .Z(n24151) );
  XOR U24047 ( .A(n24152), .B(n24153), .Z(n24143) );
  AND U24048 ( .A(n24154), .B(n24155), .Z(n24153) );
  XOR U24049 ( .A(n24152), .B(n23761), .Z(n24155) );
  XNOR U24050 ( .A(p_input[802]), .B(n24156), .Z(n23761) );
  AND U24051 ( .A(n875), .B(n24157), .Z(n24156) );
  XOR U24052 ( .A(p_input[818]), .B(p_input[802]), .Z(n24157) );
  XNOR U24053 ( .A(n23758), .B(n24152), .Z(n24154) );
  XOR U24054 ( .A(n24158), .B(n24159), .Z(n23758) );
  AND U24055 ( .A(n872), .B(n24160), .Z(n24159) );
  XOR U24056 ( .A(p_input[786]), .B(p_input[770]), .Z(n24160) );
  XOR U24057 ( .A(n24161), .B(n24162), .Z(n24152) );
  AND U24058 ( .A(n24163), .B(n24164), .Z(n24162) );
  XNOR U24059 ( .A(n24165), .B(n23774), .Z(n24164) );
  XNOR U24060 ( .A(p_input[801]), .B(n24166), .Z(n23774) );
  AND U24061 ( .A(n875), .B(n24167), .Z(n24166) );
  XNOR U24062 ( .A(p_input[817]), .B(n24168), .Z(n24167) );
  IV U24063 ( .A(p_input[801]), .Z(n24168) );
  XNOR U24064 ( .A(n23771), .B(n24161), .Z(n24163) );
  XNOR U24065 ( .A(p_input[769]), .B(n24169), .Z(n23771) );
  AND U24066 ( .A(n872), .B(n24170), .Z(n24169) );
  XOR U24067 ( .A(p_input[785]), .B(p_input[769]), .Z(n24170) );
  IV U24068 ( .A(n24165), .Z(n24161) );
  AND U24069 ( .A(n24036), .B(n24039), .Z(n24165) );
  XOR U24070 ( .A(p_input[800]), .B(n24171), .Z(n24039) );
  AND U24071 ( .A(n875), .B(n24172), .Z(n24171) );
  XOR U24072 ( .A(p_input[816]), .B(p_input[800]), .Z(n24172) );
  XOR U24073 ( .A(n24173), .B(n24174), .Z(n875) );
  AND U24074 ( .A(n24175), .B(n24176), .Z(n24174) );
  XNOR U24075 ( .A(p_input[831]), .B(n24173), .Z(n24176) );
  XOR U24076 ( .A(n24173), .B(p_input[815]), .Z(n24175) );
  XOR U24077 ( .A(n24177), .B(n24178), .Z(n24173) );
  AND U24078 ( .A(n24179), .B(n24180), .Z(n24178) );
  XNOR U24079 ( .A(p_input[830]), .B(n24177), .Z(n24180) );
  XOR U24080 ( .A(n24177), .B(p_input[814]), .Z(n24179) );
  XOR U24081 ( .A(n24181), .B(n24182), .Z(n24177) );
  AND U24082 ( .A(n24183), .B(n24184), .Z(n24182) );
  XNOR U24083 ( .A(p_input[829]), .B(n24181), .Z(n24184) );
  XOR U24084 ( .A(n24181), .B(p_input[813]), .Z(n24183) );
  XOR U24085 ( .A(n24185), .B(n24186), .Z(n24181) );
  AND U24086 ( .A(n24187), .B(n24188), .Z(n24186) );
  XNOR U24087 ( .A(p_input[828]), .B(n24185), .Z(n24188) );
  XOR U24088 ( .A(n24185), .B(p_input[812]), .Z(n24187) );
  XOR U24089 ( .A(n24189), .B(n24190), .Z(n24185) );
  AND U24090 ( .A(n24191), .B(n24192), .Z(n24190) );
  XNOR U24091 ( .A(p_input[827]), .B(n24189), .Z(n24192) );
  XOR U24092 ( .A(n24189), .B(p_input[811]), .Z(n24191) );
  XOR U24093 ( .A(n24193), .B(n24194), .Z(n24189) );
  AND U24094 ( .A(n24195), .B(n24196), .Z(n24194) );
  XNOR U24095 ( .A(p_input[826]), .B(n24193), .Z(n24196) );
  XOR U24096 ( .A(n24193), .B(p_input[810]), .Z(n24195) );
  XOR U24097 ( .A(n24197), .B(n24198), .Z(n24193) );
  AND U24098 ( .A(n24199), .B(n24200), .Z(n24198) );
  XNOR U24099 ( .A(p_input[825]), .B(n24197), .Z(n24200) );
  XOR U24100 ( .A(n24197), .B(p_input[809]), .Z(n24199) );
  XOR U24101 ( .A(n24201), .B(n24202), .Z(n24197) );
  AND U24102 ( .A(n24203), .B(n24204), .Z(n24202) );
  XNOR U24103 ( .A(p_input[824]), .B(n24201), .Z(n24204) );
  XOR U24104 ( .A(n24201), .B(p_input[808]), .Z(n24203) );
  XOR U24105 ( .A(n24205), .B(n24206), .Z(n24201) );
  AND U24106 ( .A(n24207), .B(n24208), .Z(n24206) );
  XNOR U24107 ( .A(p_input[823]), .B(n24205), .Z(n24208) );
  XOR U24108 ( .A(n24205), .B(p_input[807]), .Z(n24207) );
  XOR U24109 ( .A(n24209), .B(n24210), .Z(n24205) );
  AND U24110 ( .A(n24211), .B(n24212), .Z(n24210) );
  XNOR U24111 ( .A(p_input[822]), .B(n24209), .Z(n24212) );
  XOR U24112 ( .A(n24209), .B(p_input[806]), .Z(n24211) );
  XOR U24113 ( .A(n24213), .B(n24214), .Z(n24209) );
  AND U24114 ( .A(n24215), .B(n24216), .Z(n24214) );
  XNOR U24115 ( .A(p_input[821]), .B(n24213), .Z(n24216) );
  XOR U24116 ( .A(n24213), .B(p_input[805]), .Z(n24215) );
  XOR U24117 ( .A(n24217), .B(n24218), .Z(n24213) );
  AND U24118 ( .A(n24219), .B(n24220), .Z(n24218) );
  XNOR U24119 ( .A(p_input[820]), .B(n24217), .Z(n24220) );
  XOR U24120 ( .A(n24217), .B(p_input[804]), .Z(n24219) );
  XOR U24121 ( .A(n24221), .B(n24222), .Z(n24217) );
  AND U24122 ( .A(n24223), .B(n24224), .Z(n24222) );
  XNOR U24123 ( .A(p_input[819]), .B(n24221), .Z(n24224) );
  XOR U24124 ( .A(n24221), .B(p_input[803]), .Z(n24223) );
  XOR U24125 ( .A(n24225), .B(n24226), .Z(n24221) );
  AND U24126 ( .A(n24227), .B(n24228), .Z(n24226) );
  XNOR U24127 ( .A(p_input[818]), .B(n24225), .Z(n24228) );
  XOR U24128 ( .A(n24225), .B(p_input[802]), .Z(n24227) );
  XNOR U24129 ( .A(n24229), .B(n24230), .Z(n24225) );
  AND U24130 ( .A(n24231), .B(n24232), .Z(n24230) );
  XOR U24131 ( .A(p_input[817]), .B(n24229), .Z(n24232) );
  XNOR U24132 ( .A(p_input[801]), .B(n24229), .Z(n24231) );
  AND U24133 ( .A(p_input[816]), .B(n24233), .Z(n24229) );
  IV U24134 ( .A(p_input[800]), .Z(n24233) );
  XNOR U24135 ( .A(p_input[768]), .B(n24234), .Z(n24036) );
  AND U24136 ( .A(n872), .B(n24235), .Z(n24234) );
  XOR U24137 ( .A(p_input[784]), .B(p_input[768]), .Z(n24235) );
  XOR U24138 ( .A(n24236), .B(n24237), .Z(n872) );
  AND U24139 ( .A(n24238), .B(n24239), .Z(n24237) );
  XNOR U24140 ( .A(p_input[799]), .B(n24236), .Z(n24239) );
  XOR U24141 ( .A(n24236), .B(p_input[783]), .Z(n24238) );
  XOR U24142 ( .A(n24240), .B(n24241), .Z(n24236) );
  AND U24143 ( .A(n24242), .B(n24243), .Z(n24241) );
  XNOR U24144 ( .A(p_input[798]), .B(n24240), .Z(n24243) );
  XNOR U24145 ( .A(n24240), .B(n24050), .Z(n24242) );
  IV U24146 ( .A(p_input[782]), .Z(n24050) );
  XOR U24147 ( .A(n24244), .B(n24245), .Z(n24240) );
  AND U24148 ( .A(n24246), .B(n24247), .Z(n24245) );
  XNOR U24149 ( .A(p_input[797]), .B(n24244), .Z(n24247) );
  XNOR U24150 ( .A(n24244), .B(n24059), .Z(n24246) );
  IV U24151 ( .A(p_input[781]), .Z(n24059) );
  XOR U24152 ( .A(n24248), .B(n24249), .Z(n24244) );
  AND U24153 ( .A(n24250), .B(n24251), .Z(n24249) );
  XNOR U24154 ( .A(p_input[796]), .B(n24248), .Z(n24251) );
  XNOR U24155 ( .A(n24248), .B(n24068), .Z(n24250) );
  IV U24156 ( .A(p_input[780]), .Z(n24068) );
  XOR U24157 ( .A(n24252), .B(n24253), .Z(n24248) );
  AND U24158 ( .A(n24254), .B(n24255), .Z(n24253) );
  XNOR U24159 ( .A(p_input[795]), .B(n24252), .Z(n24255) );
  XNOR U24160 ( .A(n24252), .B(n24077), .Z(n24254) );
  IV U24161 ( .A(p_input[779]), .Z(n24077) );
  XOR U24162 ( .A(n24256), .B(n24257), .Z(n24252) );
  AND U24163 ( .A(n24258), .B(n24259), .Z(n24257) );
  XNOR U24164 ( .A(p_input[794]), .B(n24256), .Z(n24259) );
  XNOR U24165 ( .A(n24256), .B(n24086), .Z(n24258) );
  IV U24166 ( .A(p_input[778]), .Z(n24086) );
  XOR U24167 ( .A(n24260), .B(n24261), .Z(n24256) );
  AND U24168 ( .A(n24262), .B(n24263), .Z(n24261) );
  XNOR U24169 ( .A(p_input[793]), .B(n24260), .Z(n24263) );
  XNOR U24170 ( .A(n24260), .B(n24095), .Z(n24262) );
  IV U24171 ( .A(p_input[777]), .Z(n24095) );
  XOR U24172 ( .A(n24264), .B(n24265), .Z(n24260) );
  AND U24173 ( .A(n24266), .B(n24267), .Z(n24265) );
  XNOR U24174 ( .A(p_input[792]), .B(n24264), .Z(n24267) );
  XNOR U24175 ( .A(n24264), .B(n24104), .Z(n24266) );
  IV U24176 ( .A(p_input[776]), .Z(n24104) );
  XOR U24177 ( .A(n24268), .B(n24269), .Z(n24264) );
  AND U24178 ( .A(n24270), .B(n24271), .Z(n24269) );
  XNOR U24179 ( .A(p_input[791]), .B(n24268), .Z(n24271) );
  XNOR U24180 ( .A(n24268), .B(n24113), .Z(n24270) );
  IV U24181 ( .A(p_input[775]), .Z(n24113) );
  XOR U24182 ( .A(n24272), .B(n24273), .Z(n24268) );
  AND U24183 ( .A(n24274), .B(n24275), .Z(n24273) );
  XNOR U24184 ( .A(p_input[790]), .B(n24272), .Z(n24275) );
  XNOR U24185 ( .A(n24272), .B(n24122), .Z(n24274) );
  IV U24186 ( .A(p_input[774]), .Z(n24122) );
  XOR U24187 ( .A(n24276), .B(n24277), .Z(n24272) );
  AND U24188 ( .A(n24278), .B(n24279), .Z(n24277) );
  XNOR U24189 ( .A(p_input[789]), .B(n24276), .Z(n24279) );
  XNOR U24190 ( .A(n24276), .B(n24131), .Z(n24278) );
  IV U24191 ( .A(p_input[773]), .Z(n24131) );
  XOR U24192 ( .A(n24280), .B(n24281), .Z(n24276) );
  AND U24193 ( .A(n24282), .B(n24283), .Z(n24281) );
  XNOR U24194 ( .A(p_input[788]), .B(n24280), .Z(n24283) );
  XNOR U24195 ( .A(n24280), .B(n24140), .Z(n24282) );
  IV U24196 ( .A(p_input[772]), .Z(n24140) );
  XOR U24197 ( .A(n24284), .B(n24285), .Z(n24280) );
  AND U24198 ( .A(n24286), .B(n24287), .Z(n24285) );
  XNOR U24199 ( .A(p_input[787]), .B(n24284), .Z(n24287) );
  XNOR U24200 ( .A(n24284), .B(n24149), .Z(n24286) );
  IV U24201 ( .A(p_input[771]), .Z(n24149) );
  XOR U24202 ( .A(n24288), .B(n24289), .Z(n24284) );
  AND U24203 ( .A(n24290), .B(n24291), .Z(n24289) );
  XNOR U24204 ( .A(p_input[786]), .B(n24288), .Z(n24291) );
  XNOR U24205 ( .A(n24288), .B(n24158), .Z(n24290) );
  IV U24206 ( .A(p_input[770]), .Z(n24158) );
  XNOR U24207 ( .A(n24292), .B(n24293), .Z(n24288) );
  AND U24208 ( .A(n24294), .B(n24295), .Z(n24293) );
  XOR U24209 ( .A(p_input[785]), .B(n24292), .Z(n24295) );
  XNOR U24210 ( .A(p_input[769]), .B(n24292), .Z(n24294) );
  AND U24211 ( .A(p_input[784]), .B(n24296), .Z(n24292) );
  IV U24212 ( .A(p_input[768]), .Z(n24296) );
  XOR U24213 ( .A(n24297), .B(n24298), .Z(n22524) );
  AND U24214 ( .A(n957), .B(n24299), .Z(n24298) );
  XNOR U24215 ( .A(n24300), .B(n24297), .Z(n24299) );
  XOR U24216 ( .A(n24301), .B(n24302), .Z(n957) );
  AND U24217 ( .A(n24303), .B(n24304), .Z(n24302) );
  XNOR U24218 ( .A(n22539), .B(n24301), .Z(n24304) );
  AND U24219 ( .A(n24305), .B(n24306), .Z(n22539) );
  XNOR U24220 ( .A(n24301), .B(n22536), .Z(n24303) );
  IV U24221 ( .A(n24307), .Z(n22536) );
  AND U24222 ( .A(n24308), .B(n24309), .Z(n24307) );
  XOR U24223 ( .A(n24310), .B(n24311), .Z(n24301) );
  AND U24224 ( .A(n24312), .B(n24313), .Z(n24311) );
  XOR U24225 ( .A(n24310), .B(n22551), .Z(n24313) );
  XOR U24226 ( .A(n24314), .B(n24315), .Z(n22551) );
  AND U24227 ( .A(n827), .B(n24316), .Z(n24315) );
  XOR U24228 ( .A(n24317), .B(n24314), .Z(n24316) );
  XNOR U24229 ( .A(n22548), .B(n24310), .Z(n24312) );
  XOR U24230 ( .A(n24318), .B(n24319), .Z(n22548) );
  AND U24231 ( .A(n824), .B(n24320), .Z(n24319) );
  XOR U24232 ( .A(n24321), .B(n24318), .Z(n24320) );
  XOR U24233 ( .A(n24322), .B(n24323), .Z(n24310) );
  AND U24234 ( .A(n24324), .B(n24325), .Z(n24323) );
  XOR U24235 ( .A(n24322), .B(n22563), .Z(n24325) );
  XOR U24236 ( .A(n24326), .B(n24327), .Z(n22563) );
  AND U24237 ( .A(n827), .B(n24328), .Z(n24327) );
  XOR U24238 ( .A(n24329), .B(n24326), .Z(n24328) );
  XNOR U24239 ( .A(n22560), .B(n24322), .Z(n24324) );
  XOR U24240 ( .A(n24330), .B(n24331), .Z(n22560) );
  AND U24241 ( .A(n824), .B(n24332), .Z(n24331) );
  XOR U24242 ( .A(n24333), .B(n24330), .Z(n24332) );
  XOR U24243 ( .A(n24334), .B(n24335), .Z(n24322) );
  AND U24244 ( .A(n24336), .B(n24337), .Z(n24335) );
  XOR U24245 ( .A(n24334), .B(n22575), .Z(n24337) );
  XOR U24246 ( .A(n24338), .B(n24339), .Z(n22575) );
  AND U24247 ( .A(n827), .B(n24340), .Z(n24339) );
  XOR U24248 ( .A(n24341), .B(n24338), .Z(n24340) );
  XNOR U24249 ( .A(n22572), .B(n24334), .Z(n24336) );
  XOR U24250 ( .A(n24342), .B(n24343), .Z(n22572) );
  AND U24251 ( .A(n824), .B(n24344), .Z(n24343) );
  XOR U24252 ( .A(n24345), .B(n24342), .Z(n24344) );
  XOR U24253 ( .A(n24346), .B(n24347), .Z(n24334) );
  AND U24254 ( .A(n24348), .B(n24349), .Z(n24347) );
  XOR U24255 ( .A(n24346), .B(n22587), .Z(n24349) );
  XOR U24256 ( .A(n24350), .B(n24351), .Z(n22587) );
  AND U24257 ( .A(n827), .B(n24352), .Z(n24351) );
  XOR U24258 ( .A(n24353), .B(n24350), .Z(n24352) );
  XNOR U24259 ( .A(n22584), .B(n24346), .Z(n24348) );
  XOR U24260 ( .A(n24354), .B(n24355), .Z(n22584) );
  AND U24261 ( .A(n824), .B(n24356), .Z(n24355) );
  XOR U24262 ( .A(n24357), .B(n24354), .Z(n24356) );
  XOR U24263 ( .A(n24358), .B(n24359), .Z(n24346) );
  AND U24264 ( .A(n24360), .B(n24361), .Z(n24359) );
  XOR U24265 ( .A(n24358), .B(n22599), .Z(n24361) );
  XOR U24266 ( .A(n24362), .B(n24363), .Z(n22599) );
  AND U24267 ( .A(n827), .B(n24364), .Z(n24363) );
  XOR U24268 ( .A(n24365), .B(n24362), .Z(n24364) );
  XNOR U24269 ( .A(n22596), .B(n24358), .Z(n24360) );
  XOR U24270 ( .A(n24366), .B(n24367), .Z(n22596) );
  AND U24271 ( .A(n824), .B(n24368), .Z(n24367) );
  XOR U24272 ( .A(n24369), .B(n24366), .Z(n24368) );
  XOR U24273 ( .A(n24370), .B(n24371), .Z(n24358) );
  AND U24274 ( .A(n24372), .B(n24373), .Z(n24371) );
  XOR U24275 ( .A(n24370), .B(n22611), .Z(n24373) );
  XOR U24276 ( .A(n24374), .B(n24375), .Z(n22611) );
  AND U24277 ( .A(n827), .B(n24376), .Z(n24375) );
  XOR U24278 ( .A(n24377), .B(n24374), .Z(n24376) );
  XNOR U24279 ( .A(n22608), .B(n24370), .Z(n24372) );
  XOR U24280 ( .A(n24378), .B(n24379), .Z(n22608) );
  AND U24281 ( .A(n824), .B(n24380), .Z(n24379) );
  XOR U24282 ( .A(n24381), .B(n24378), .Z(n24380) );
  XOR U24283 ( .A(n24382), .B(n24383), .Z(n24370) );
  AND U24284 ( .A(n24384), .B(n24385), .Z(n24383) );
  XOR U24285 ( .A(n24382), .B(n22623), .Z(n24385) );
  XOR U24286 ( .A(n24386), .B(n24387), .Z(n22623) );
  AND U24287 ( .A(n827), .B(n24388), .Z(n24387) );
  XOR U24288 ( .A(n24389), .B(n24386), .Z(n24388) );
  XNOR U24289 ( .A(n22620), .B(n24382), .Z(n24384) );
  XOR U24290 ( .A(n24390), .B(n24391), .Z(n22620) );
  AND U24291 ( .A(n824), .B(n24392), .Z(n24391) );
  XOR U24292 ( .A(n24393), .B(n24390), .Z(n24392) );
  XOR U24293 ( .A(n24394), .B(n24395), .Z(n24382) );
  AND U24294 ( .A(n24396), .B(n24397), .Z(n24395) );
  XOR U24295 ( .A(n24394), .B(n22635), .Z(n24397) );
  XOR U24296 ( .A(n24398), .B(n24399), .Z(n22635) );
  AND U24297 ( .A(n827), .B(n24400), .Z(n24399) );
  XOR U24298 ( .A(n24401), .B(n24398), .Z(n24400) );
  XNOR U24299 ( .A(n22632), .B(n24394), .Z(n24396) );
  XOR U24300 ( .A(n24402), .B(n24403), .Z(n22632) );
  AND U24301 ( .A(n824), .B(n24404), .Z(n24403) );
  XOR U24302 ( .A(n24405), .B(n24402), .Z(n24404) );
  XOR U24303 ( .A(n24406), .B(n24407), .Z(n24394) );
  AND U24304 ( .A(n24408), .B(n24409), .Z(n24407) );
  XOR U24305 ( .A(n24406), .B(n22647), .Z(n24409) );
  XOR U24306 ( .A(n24410), .B(n24411), .Z(n22647) );
  AND U24307 ( .A(n827), .B(n24412), .Z(n24411) );
  XOR U24308 ( .A(n24413), .B(n24410), .Z(n24412) );
  XNOR U24309 ( .A(n22644), .B(n24406), .Z(n24408) );
  XOR U24310 ( .A(n24414), .B(n24415), .Z(n22644) );
  AND U24311 ( .A(n824), .B(n24416), .Z(n24415) );
  XOR U24312 ( .A(n24417), .B(n24414), .Z(n24416) );
  XOR U24313 ( .A(n24418), .B(n24419), .Z(n24406) );
  AND U24314 ( .A(n24420), .B(n24421), .Z(n24419) );
  XOR U24315 ( .A(n24418), .B(n22659), .Z(n24421) );
  XOR U24316 ( .A(n24422), .B(n24423), .Z(n22659) );
  AND U24317 ( .A(n827), .B(n24424), .Z(n24423) );
  XOR U24318 ( .A(n24425), .B(n24422), .Z(n24424) );
  XNOR U24319 ( .A(n22656), .B(n24418), .Z(n24420) );
  XOR U24320 ( .A(n24426), .B(n24427), .Z(n22656) );
  AND U24321 ( .A(n824), .B(n24428), .Z(n24427) );
  XOR U24322 ( .A(n24429), .B(n24426), .Z(n24428) );
  XOR U24323 ( .A(n24430), .B(n24431), .Z(n24418) );
  AND U24324 ( .A(n24432), .B(n24433), .Z(n24431) );
  XOR U24325 ( .A(n24430), .B(n22671), .Z(n24433) );
  XOR U24326 ( .A(n24434), .B(n24435), .Z(n22671) );
  AND U24327 ( .A(n827), .B(n24436), .Z(n24435) );
  XOR U24328 ( .A(n24437), .B(n24434), .Z(n24436) );
  XNOR U24329 ( .A(n22668), .B(n24430), .Z(n24432) );
  XOR U24330 ( .A(n24438), .B(n24439), .Z(n22668) );
  AND U24331 ( .A(n824), .B(n24440), .Z(n24439) );
  XOR U24332 ( .A(n24441), .B(n24438), .Z(n24440) );
  XOR U24333 ( .A(n24442), .B(n24443), .Z(n24430) );
  AND U24334 ( .A(n24444), .B(n24445), .Z(n24443) );
  XOR U24335 ( .A(n24442), .B(n22683), .Z(n24445) );
  XOR U24336 ( .A(n24446), .B(n24447), .Z(n22683) );
  AND U24337 ( .A(n827), .B(n24448), .Z(n24447) );
  XOR U24338 ( .A(n24449), .B(n24446), .Z(n24448) );
  XNOR U24339 ( .A(n22680), .B(n24442), .Z(n24444) );
  XOR U24340 ( .A(n24450), .B(n24451), .Z(n22680) );
  AND U24341 ( .A(n824), .B(n24452), .Z(n24451) );
  XOR U24342 ( .A(n24453), .B(n24450), .Z(n24452) );
  XOR U24343 ( .A(n24454), .B(n24455), .Z(n24442) );
  AND U24344 ( .A(n24456), .B(n24457), .Z(n24455) );
  XOR U24345 ( .A(n24454), .B(n22695), .Z(n24457) );
  XOR U24346 ( .A(n24458), .B(n24459), .Z(n22695) );
  AND U24347 ( .A(n827), .B(n24460), .Z(n24459) );
  XOR U24348 ( .A(n24461), .B(n24458), .Z(n24460) );
  XNOR U24349 ( .A(n22692), .B(n24454), .Z(n24456) );
  XOR U24350 ( .A(n24462), .B(n24463), .Z(n22692) );
  AND U24351 ( .A(n824), .B(n24464), .Z(n24463) );
  XOR U24352 ( .A(n24465), .B(n24462), .Z(n24464) );
  XOR U24353 ( .A(n24466), .B(n24467), .Z(n24454) );
  AND U24354 ( .A(n24468), .B(n24469), .Z(n24467) );
  XNOR U24355 ( .A(n24470), .B(n22708), .Z(n24469) );
  XOR U24356 ( .A(n24471), .B(n24472), .Z(n22708) );
  AND U24357 ( .A(n827), .B(n24473), .Z(n24472) );
  XOR U24358 ( .A(n24471), .B(n24474), .Z(n24473) );
  XNOR U24359 ( .A(n22705), .B(n24466), .Z(n24468) );
  XOR U24360 ( .A(n24475), .B(n24476), .Z(n22705) );
  AND U24361 ( .A(n824), .B(n24477), .Z(n24476) );
  XOR U24362 ( .A(n24475), .B(n24478), .Z(n24477) );
  IV U24363 ( .A(n24470), .Z(n24466) );
  AND U24364 ( .A(n24297), .B(n24300), .Z(n24470) );
  XNOR U24365 ( .A(n24479), .B(n24480), .Z(n24300) );
  AND U24366 ( .A(n827), .B(n24481), .Z(n24480) );
  XNOR U24367 ( .A(n24482), .B(n24479), .Z(n24481) );
  XOR U24368 ( .A(n24483), .B(n24484), .Z(n827) );
  AND U24369 ( .A(n24485), .B(n24486), .Z(n24484) );
  XNOR U24370 ( .A(n24305), .B(n24483), .Z(n24486) );
  AND U24371 ( .A(n24487), .B(n24488), .Z(n24305) );
  XOR U24372 ( .A(n24483), .B(n24306), .Z(n24485) );
  AND U24373 ( .A(n24489), .B(n24490), .Z(n24306) );
  XOR U24374 ( .A(n24491), .B(n24492), .Z(n24483) );
  AND U24375 ( .A(n24493), .B(n24494), .Z(n24492) );
  XOR U24376 ( .A(n24491), .B(n24317), .Z(n24494) );
  XOR U24377 ( .A(n24495), .B(n24496), .Z(n24317) );
  AND U24378 ( .A(n555), .B(n24497), .Z(n24496) );
  XOR U24379 ( .A(n24498), .B(n24495), .Z(n24497) );
  XNOR U24380 ( .A(n24314), .B(n24491), .Z(n24493) );
  XOR U24381 ( .A(n24499), .B(n24500), .Z(n24314) );
  AND U24382 ( .A(n553), .B(n24501), .Z(n24500) );
  XOR U24383 ( .A(n24502), .B(n24499), .Z(n24501) );
  XOR U24384 ( .A(n24503), .B(n24504), .Z(n24491) );
  AND U24385 ( .A(n24505), .B(n24506), .Z(n24504) );
  XOR U24386 ( .A(n24503), .B(n24329), .Z(n24506) );
  XOR U24387 ( .A(n24507), .B(n24508), .Z(n24329) );
  AND U24388 ( .A(n555), .B(n24509), .Z(n24508) );
  XOR U24389 ( .A(n24510), .B(n24507), .Z(n24509) );
  XNOR U24390 ( .A(n24326), .B(n24503), .Z(n24505) );
  XOR U24391 ( .A(n24511), .B(n24512), .Z(n24326) );
  AND U24392 ( .A(n553), .B(n24513), .Z(n24512) );
  XOR U24393 ( .A(n24514), .B(n24511), .Z(n24513) );
  XOR U24394 ( .A(n24515), .B(n24516), .Z(n24503) );
  AND U24395 ( .A(n24517), .B(n24518), .Z(n24516) );
  XOR U24396 ( .A(n24515), .B(n24341), .Z(n24518) );
  XOR U24397 ( .A(n24519), .B(n24520), .Z(n24341) );
  AND U24398 ( .A(n555), .B(n24521), .Z(n24520) );
  XOR U24399 ( .A(n24522), .B(n24519), .Z(n24521) );
  XNOR U24400 ( .A(n24338), .B(n24515), .Z(n24517) );
  XOR U24401 ( .A(n24523), .B(n24524), .Z(n24338) );
  AND U24402 ( .A(n553), .B(n24525), .Z(n24524) );
  XOR U24403 ( .A(n24526), .B(n24523), .Z(n24525) );
  XOR U24404 ( .A(n24527), .B(n24528), .Z(n24515) );
  AND U24405 ( .A(n24529), .B(n24530), .Z(n24528) );
  XOR U24406 ( .A(n24527), .B(n24353), .Z(n24530) );
  XOR U24407 ( .A(n24531), .B(n24532), .Z(n24353) );
  AND U24408 ( .A(n555), .B(n24533), .Z(n24532) );
  XOR U24409 ( .A(n24534), .B(n24531), .Z(n24533) );
  XNOR U24410 ( .A(n24350), .B(n24527), .Z(n24529) );
  XOR U24411 ( .A(n24535), .B(n24536), .Z(n24350) );
  AND U24412 ( .A(n553), .B(n24537), .Z(n24536) );
  XOR U24413 ( .A(n24538), .B(n24535), .Z(n24537) );
  XOR U24414 ( .A(n24539), .B(n24540), .Z(n24527) );
  AND U24415 ( .A(n24541), .B(n24542), .Z(n24540) );
  XOR U24416 ( .A(n24539), .B(n24365), .Z(n24542) );
  XOR U24417 ( .A(n24543), .B(n24544), .Z(n24365) );
  AND U24418 ( .A(n555), .B(n24545), .Z(n24544) );
  XOR U24419 ( .A(n24546), .B(n24543), .Z(n24545) );
  XNOR U24420 ( .A(n24362), .B(n24539), .Z(n24541) );
  XOR U24421 ( .A(n24547), .B(n24548), .Z(n24362) );
  AND U24422 ( .A(n553), .B(n24549), .Z(n24548) );
  XOR U24423 ( .A(n24550), .B(n24547), .Z(n24549) );
  XOR U24424 ( .A(n24551), .B(n24552), .Z(n24539) );
  AND U24425 ( .A(n24553), .B(n24554), .Z(n24552) );
  XOR U24426 ( .A(n24551), .B(n24377), .Z(n24554) );
  XOR U24427 ( .A(n24555), .B(n24556), .Z(n24377) );
  AND U24428 ( .A(n555), .B(n24557), .Z(n24556) );
  XOR U24429 ( .A(n24558), .B(n24555), .Z(n24557) );
  XNOR U24430 ( .A(n24374), .B(n24551), .Z(n24553) );
  XOR U24431 ( .A(n24559), .B(n24560), .Z(n24374) );
  AND U24432 ( .A(n553), .B(n24561), .Z(n24560) );
  XOR U24433 ( .A(n24562), .B(n24559), .Z(n24561) );
  XOR U24434 ( .A(n24563), .B(n24564), .Z(n24551) );
  AND U24435 ( .A(n24565), .B(n24566), .Z(n24564) );
  XOR U24436 ( .A(n24563), .B(n24389), .Z(n24566) );
  XOR U24437 ( .A(n24567), .B(n24568), .Z(n24389) );
  AND U24438 ( .A(n555), .B(n24569), .Z(n24568) );
  XOR U24439 ( .A(n24570), .B(n24567), .Z(n24569) );
  XNOR U24440 ( .A(n24386), .B(n24563), .Z(n24565) );
  XOR U24441 ( .A(n24571), .B(n24572), .Z(n24386) );
  AND U24442 ( .A(n553), .B(n24573), .Z(n24572) );
  XOR U24443 ( .A(n24574), .B(n24571), .Z(n24573) );
  XOR U24444 ( .A(n24575), .B(n24576), .Z(n24563) );
  AND U24445 ( .A(n24577), .B(n24578), .Z(n24576) );
  XOR U24446 ( .A(n24575), .B(n24401), .Z(n24578) );
  XOR U24447 ( .A(n24579), .B(n24580), .Z(n24401) );
  AND U24448 ( .A(n555), .B(n24581), .Z(n24580) );
  XOR U24449 ( .A(n24582), .B(n24579), .Z(n24581) );
  XNOR U24450 ( .A(n24398), .B(n24575), .Z(n24577) );
  XOR U24451 ( .A(n24583), .B(n24584), .Z(n24398) );
  AND U24452 ( .A(n553), .B(n24585), .Z(n24584) );
  XOR U24453 ( .A(n24586), .B(n24583), .Z(n24585) );
  XOR U24454 ( .A(n24587), .B(n24588), .Z(n24575) );
  AND U24455 ( .A(n24589), .B(n24590), .Z(n24588) );
  XOR U24456 ( .A(n24587), .B(n24413), .Z(n24590) );
  XOR U24457 ( .A(n24591), .B(n24592), .Z(n24413) );
  AND U24458 ( .A(n555), .B(n24593), .Z(n24592) );
  XOR U24459 ( .A(n24594), .B(n24591), .Z(n24593) );
  XNOR U24460 ( .A(n24410), .B(n24587), .Z(n24589) );
  XOR U24461 ( .A(n24595), .B(n24596), .Z(n24410) );
  AND U24462 ( .A(n553), .B(n24597), .Z(n24596) );
  XOR U24463 ( .A(n24598), .B(n24595), .Z(n24597) );
  XOR U24464 ( .A(n24599), .B(n24600), .Z(n24587) );
  AND U24465 ( .A(n24601), .B(n24602), .Z(n24600) );
  XOR U24466 ( .A(n24599), .B(n24425), .Z(n24602) );
  XOR U24467 ( .A(n24603), .B(n24604), .Z(n24425) );
  AND U24468 ( .A(n555), .B(n24605), .Z(n24604) );
  XOR U24469 ( .A(n24606), .B(n24603), .Z(n24605) );
  XNOR U24470 ( .A(n24422), .B(n24599), .Z(n24601) );
  XOR U24471 ( .A(n24607), .B(n24608), .Z(n24422) );
  AND U24472 ( .A(n553), .B(n24609), .Z(n24608) );
  XOR U24473 ( .A(n24610), .B(n24607), .Z(n24609) );
  XOR U24474 ( .A(n24611), .B(n24612), .Z(n24599) );
  AND U24475 ( .A(n24613), .B(n24614), .Z(n24612) );
  XOR U24476 ( .A(n24611), .B(n24437), .Z(n24614) );
  XOR U24477 ( .A(n24615), .B(n24616), .Z(n24437) );
  AND U24478 ( .A(n555), .B(n24617), .Z(n24616) );
  XOR U24479 ( .A(n24618), .B(n24615), .Z(n24617) );
  XNOR U24480 ( .A(n24434), .B(n24611), .Z(n24613) );
  XOR U24481 ( .A(n24619), .B(n24620), .Z(n24434) );
  AND U24482 ( .A(n553), .B(n24621), .Z(n24620) );
  XOR U24483 ( .A(n24622), .B(n24619), .Z(n24621) );
  XOR U24484 ( .A(n24623), .B(n24624), .Z(n24611) );
  AND U24485 ( .A(n24625), .B(n24626), .Z(n24624) );
  XOR U24486 ( .A(n24623), .B(n24449), .Z(n24626) );
  XOR U24487 ( .A(n24627), .B(n24628), .Z(n24449) );
  AND U24488 ( .A(n555), .B(n24629), .Z(n24628) );
  XOR U24489 ( .A(n24630), .B(n24627), .Z(n24629) );
  XNOR U24490 ( .A(n24446), .B(n24623), .Z(n24625) );
  XOR U24491 ( .A(n24631), .B(n24632), .Z(n24446) );
  AND U24492 ( .A(n553), .B(n24633), .Z(n24632) );
  XOR U24493 ( .A(n24634), .B(n24631), .Z(n24633) );
  XOR U24494 ( .A(n24635), .B(n24636), .Z(n24623) );
  AND U24495 ( .A(n24637), .B(n24638), .Z(n24636) );
  XOR U24496 ( .A(n24635), .B(n24461), .Z(n24638) );
  XOR U24497 ( .A(n24639), .B(n24640), .Z(n24461) );
  AND U24498 ( .A(n555), .B(n24641), .Z(n24640) );
  XOR U24499 ( .A(n24642), .B(n24639), .Z(n24641) );
  XNOR U24500 ( .A(n24458), .B(n24635), .Z(n24637) );
  XOR U24501 ( .A(n24643), .B(n24644), .Z(n24458) );
  AND U24502 ( .A(n553), .B(n24645), .Z(n24644) );
  XOR U24503 ( .A(n24646), .B(n24643), .Z(n24645) );
  XOR U24504 ( .A(n24647), .B(n24648), .Z(n24635) );
  AND U24505 ( .A(n24649), .B(n24650), .Z(n24648) );
  XNOR U24506 ( .A(n24651), .B(n24474), .Z(n24650) );
  XOR U24507 ( .A(n24652), .B(n24653), .Z(n24474) );
  AND U24508 ( .A(n555), .B(n24654), .Z(n24653) );
  XOR U24509 ( .A(n24652), .B(n24655), .Z(n24654) );
  XNOR U24510 ( .A(n24471), .B(n24647), .Z(n24649) );
  XOR U24511 ( .A(n24656), .B(n24657), .Z(n24471) );
  AND U24512 ( .A(n553), .B(n24658), .Z(n24657) );
  XOR U24513 ( .A(n24656), .B(n24659), .Z(n24658) );
  IV U24514 ( .A(n24651), .Z(n24647) );
  AND U24515 ( .A(n24479), .B(n24482), .Z(n24651) );
  XNOR U24516 ( .A(n24660), .B(n24661), .Z(n24482) );
  AND U24517 ( .A(n555), .B(n24662), .Z(n24661) );
  XNOR U24518 ( .A(n24663), .B(n24660), .Z(n24662) );
  XOR U24519 ( .A(n24664), .B(n24665), .Z(n555) );
  AND U24520 ( .A(n24666), .B(n24667), .Z(n24665) );
  XNOR U24521 ( .A(n24487), .B(n24664), .Z(n24667) );
  AND U24522 ( .A(p_input[767]), .B(p_input[751]), .Z(n24487) );
  XOR U24523 ( .A(n24664), .B(n24488), .Z(n24666) );
  AND U24524 ( .A(p_input[735]), .B(p_input[719]), .Z(n24488) );
  XOR U24525 ( .A(n24668), .B(n24669), .Z(n24664) );
  AND U24526 ( .A(n24670), .B(n24671), .Z(n24669) );
  XOR U24527 ( .A(n24668), .B(n24498), .Z(n24671) );
  XNOR U24528 ( .A(p_input[750]), .B(n24672), .Z(n24498) );
  AND U24529 ( .A(n887), .B(n24673), .Z(n24672) );
  XOR U24530 ( .A(p_input[766]), .B(p_input[750]), .Z(n24673) );
  XNOR U24531 ( .A(n24495), .B(n24668), .Z(n24670) );
  XOR U24532 ( .A(n24674), .B(n24675), .Z(n24495) );
  AND U24533 ( .A(n885), .B(n24676), .Z(n24675) );
  XOR U24534 ( .A(p_input[734]), .B(p_input[718]), .Z(n24676) );
  XOR U24535 ( .A(n24677), .B(n24678), .Z(n24668) );
  AND U24536 ( .A(n24679), .B(n24680), .Z(n24678) );
  XOR U24537 ( .A(n24677), .B(n24510), .Z(n24680) );
  XNOR U24538 ( .A(p_input[749]), .B(n24681), .Z(n24510) );
  AND U24539 ( .A(n887), .B(n24682), .Z(n24681) );
  XOR U24540 ( .A(p_input[765]), .B(p_input[749]), .Z(n24682) );
  XNOR U24541 ( .A(n24507), .B(n24677), .Z(n24679) );
  XOR U24542 ( .A(n24683), .B(n24684), .Z(n24507) );
  AND U24543 ( .A(n885), .B(n24685), .Z(n24684) );
  XOR U24544 ( .A(p_input[733]), .B(p_input[717]), .Z(n24685) );
  XOR U24545 ( .A(n24686), .B(n24687), .Z(n24677) );
  AND U24546 ( .A(n24688), .B(n24689), .Z(n24687) );
  XOR U24547 ( .A(n24686), .B(n24522), .Z(n24689) );
  XNOR U24548 ( .A(p_input[748]), .B(n24690), .Z(n24522) );
  AND U24549 ( .A(n887), .B(n24691), .Z(n24690) );
  XOR U24550 ( .A(p_input[764]), .B(p_input[748]), .Z(n24691) );
  XNOR U24551 ( .A(n24519), .B(n24686), .Z(n24688) );
  XOR U24552 ( .A(n24692), .B(n24693), .Z(n24519) );
  AND U24553 ( .A(n885), .B(n24694), .Z(n24693) );
  XOR U24554 ( .A(p_input[732]), .B(p_input[716]), .Z(n24694) );
  XOR U24555 ( .A(n24695), .B(n24696), .Z(n24686) );
  AND U24556 ( .A(n24697), .B(n24698), .Z(n24696) );
  XOR U24557 ( .A(n24695), .B(n24534), .Z(n24698) );
  XNOR U24558 ( .A(p_input[747]), .B(n24699), .Z(n24534) );
  AND U24559 ( .A(n887), .B(n24700), .Z(n24699) );
  XOR U24560 ( .A(p_input[763]), .B(p_input[747]), .Z(n24700) );
  XNOR U24561 ( .A(n24531), .B(n24695), .Z(n24697) );
  XOR U24562 ( .A(n24701), .B(n24702), .Z(n24531) );
  AND U24563 ( .A(n885), .B(n24703), .Z(n24702) );
  XOR U24564 ( .A(p_input[731]), .B(p_input[715]), .Z(n24703) );
  XOR U24565 ( .A(n24704), .B(n24705), .Z(n24695) );
  AND U24566 ( .A(n24706), .B(n24707), .Z(n24705) );
  XOR U24567 ( .A(n24704), .B(n24546), .Z(n24707) );
  XNOR U24568 ( .A(p_input[746]), .B(n24708), .Z(n24546) );
  AND U24569 ( .A(n887), .B(n24709), .Z(n24708) );
  XOR U24570 ( .A(p_input[762]), .B(p_input[746]), .Z(n24709) );
  XNOR U24571 ( .A(n24543), .B(n24704), .Z(n24706) );
  XOR U24572 ( .A(n24710), .B(n24711), .Z(n24543) );
  AND U24573 ( .A(n885), .B(n24712), .Z(n24711) );
  XOR U24574 ( .A(p_input[730]), .B(p_input[714]), .Z(n24712) );
  XOR U24575 ( .A(n24713), .B(n24714), .Z(n24704) );
  AND U24576 ( .A(n24715), .B(n24716), .Z(n24714) );
  XOR U24577 ( .A(n24713), .B(n24558), .Z(n24716) );
  XNOR U24578 ( .A(p_input[745]), .B(n24717), .Z(n24558) );
  AND U24579 ( .A(n887), .B(n24718), .Z(n24717) );
  XOR U24580 ( .A(p_input[761]), .B(p_input[745]), .Z(n24718) );
  XNOR U24581 ( .A(n24555), .B(n24713), .Z(n24715) );
  XOR U24582 ( .A(n24719), .B(n24720), .Z(n24555) );
  AND U24583 ( .A(n885), .B(n24721), .Z(n24720) );
  XOR U24584 ( .A(p_input[729]), .B(p_input[713]), .Z(n24721) );
  XOR U24585 ( .A(n24722), .B(n24723), .Z(n24713) );
  AND U24586 ( .A(n24724), .B(n24725), .Z(n24723) );
  XOR U24587 ( .A(n24722), .B(n24570), .Z(n24725) );
  XNOR U24588 ( .A(p_input[744]), .B(n24726), .Z(n24570) );
  AND U24589 ( .A(n887), .B(n24727), .Z(n24726) );
  XOR U24590 ( .A(p_input[760]), .B(p_input[744]), .Z(n24727) );
  XNOR U24591 ( .A(n24567), .B(n24722), .Z(n24724) );
  XOR U24592 ( .A(n24728), .B(n24729), .Z(n24567) );
  AND U24593 ( .A(n885), .B(n24730), .Z(n24729) );
  XOR U24594 ( .A(p_input[728]), .B(p_input[712]), .Z(n24730) );
  XOR U24595 ( .A(n24731), .B(n24732), .Z(n24722) );
  AND U24596 ( .A(n24733), .B(n24734), .Z(n24732) );
  XOR U24597 ( .A(n24731), .B(n24582), .Z(n24734) );
  XNOR U24598 ( .A(p_input[743]), .B(n24735), .Z(n24582) );
  AND U24599 ( .A(n887), .B(n24736), .Z(n24735) );
  XOR U24600 ( .A(p_input[759]), .B(p_input[743]), .Z(n24736) );
  XNOR U24601 ( .A(n24579), .B(n24731), .Z(n24733) );
  XOR U24602 ( .A(n24737), .B(n24738), .Z(n24579) );
  AND U24603 ( .A(n885), .B(n24739), .Z(n24738) );
  XOR U24604 ( .A(p_input[727]), .B(p_input[711]), .Z(n24739) );
  XOR U24605 ( .A(n24740), .B(n24741), .Z(n24731) );
  AND U24606 ( .A(n24742), .B(n24743), .Z(n24741) );
  XOR U24607 ( .A(n24740), .B(n24594), .Z(n24743) );
  XNOR U24608 ( .A(p_input[742]), .B(n24744), .Z(n24594) );
  AND U24609 ( .A(n887), .B(n24745), .Z(n24744) );
  XOR U24610 ( .A(p_input[758]), .B(p_input[742]), .Z(n24745) );
  XNOR U24611 ( .A(n24591), .B(n24740), .Z(n24742) );
  XOR U24612 ( .A(n24746), .B(n24747), .Z(n24591) );
  AND U24613 ( .A(n885), .B(n24748), .Z(n24747) );
  XOR U24614 ( .A(p_input[726]), .B(p_input[710]), .Z(n24748) );
  XOR U24615 ( .A(n24749), .B(n24750), .Z(n24740) );
  AND U24616 ( .A(n24751), .B(n24752), .Z(n24750) );
  XOR U24617 ( .A(n24749), .B(n24606), .Z(n24752) );
  XNOR U24618 ( .A(p_input[741]), .B(n24753), .Z(n24606) );
  AND U24619 ( .A(n887), .B(n24754), .Z(n24753) );
  XOR U24620 ( .A(p_input[757]), .B(p_input[741]), .Z(n24754) );
  XNOR U24621 ( .A(n24603), .B(n24749), .Z(n24751) );
  XOR U24622 ( .A(n24755), .B(n24756), .Z(n24603) );
  AND U24623 ( .A(n885), .B(n24757), .Z(n24756) );
  XOR U24624 ( .A(p_input[725]), .B(p_input[709]), .Z(n24757) );
  XOR U24625 ( .A(n24758), .B(n24759), .Z(n24749) );
  AND U24626 ( .A(n24760), .B(n24761), .Z(n24759) );
  XOR U24627 ( .A(n24758), .B(n24618), .Z(n24761) );
  XNOR U24628 ( .A(p_input[740]), .B(n24762), .Z(n24618) );
  AND U24629 ( .A(n887), .B(n24763), .Z(n24762) );
  XOR U24630 ( .A(p_input[756]), .B(p_input[740]), .Z(n24763) );
  XNOR U24631 ( .A(n24615), .B(n24758), .Z(n24760) );
  XOR U24632 ( .A(n24764), .B(n24765), .Z(n24615) );
  AND U24633 ( .A(n885), .B(n24766), .Z(n24765) );
  XOR U24634 ( .A(p_input[724]), .B(p_input[708]), .Z(n24766) );
  XOR U24635 ( .A(n24767), .B(n24768), .Z(n24758) );
  AND U24636 ( .A(n24769), .B(n24770), .Z(n24768) );
  XOR U24637 ( .A(n24767), .B(n24630), .Z(n24770) );
  XNOR U24638 ( .A(p_input[739]), .B(n24771), .Z(n24630) );
  AND U24639 ( .A(n887), .B(n24772), .Z(n24771) );
  XOR U24640 ( .A(p_input[755]), .B(p_input[739]), .Z(n24772) );
  XNOR U24641 ( .A(n24627), .B(n24767), .Z(n24769) );
  XOR U24642 ( .A(n24773), .B(n24774), .Z(n24627) );
  AND U24643 ( .A(n885), .B(n24775), .Z(n24774) );
  XOR U24644 ( .A(p_input[723]), .B(p_input[707]), .Z(n24775) );
  XOR U24645 ( .A(n24776), .B(n24777), .Z(n24767) );
  AND U24646 ( .A(n24778), .B(n24779), .Z(n24777) );
  XOR U24647 ( .A(n24776), .B(n24642), .Z(n24779) );
  XNOR U24648 ( .A(p_input[738]), .B(n24780), .Z(n24642) );
  AND U24649 ( .A(n887), .B(n24781), .Z(n24780) );
  XOR U24650 ( .A(p_input[754]), .B(p_input[738]), .Z(n24781) );
  XNOR U24651 ( .A(n24639), .B(n24776), .Z(n24778) );
  XOR U24652 ( .A(n24782), .B(n24783), .Z(n24639) );
  AND U24653 ( .A(n885), .B(n24784), .Z(n24783) );
  XOR U24654 ( .A(p_input[722]), .B(p_input[706]), .Z(n24784) );
  XOR U24655 ( .A(n24785), .B(n24786), .Z(n24776) );
  AND U24656 ( .A(n24787), .B(n24788), .Z(n24786) );
  XNOR U24657 ( .A(n24789), .B(n24655), .Z(n24788) );
  XNOR U24658 ( .A(p_input[737]), .B(n24790), .Z(n24655) );
  AND U24659 ( .A(n887), .B(n24791), .Z(n24790) );
  XNOR U24660 ( .A(p_input[753]), .B(n24792), .Z(n24791) );
  IV U24661 ( .A(p_input[737]), .Z(n24792) );
  XNOR U24662 ( .A(n24652), .B(n24785), .Z(n24787) );
  XNOR U24663 ( .A(p_input[705]), .B(n24793), .Z(n24652) );
  AND U24664 ( .A(n885), .B(n24794), .Z(n24793) );
  XOR U24665 ( .A(p_input[721]), .B(p_input[705]), .Z(n24794) );
  IV U24666 ( .A(n24789), .Z(n24785) );
  AND U24667 ( .A(n24660), .B(n24663), .Z(n24789) );
  XOR U24668 ( .A(p_input[736]), .B(n24795), .Z(n24663) );
  AND U24669 ( .A(n887), .B(n24796), .Z(n24795) );
  XOR U24670 ( .A(p_input[752]), .B(p_input[736]), .Z(n24796) );
  XOR U24671 ( .A(n24797), .B(n24798), .Z(n887) );
  AND U24672 ( .A(n24799), .B(n24800), .Z(n24798) );
  XNOR U24673 ( .A(p_input[767]), .B(n24797), .Z(n24800) );
  XOR U24674 ( .A(n24797), .B(p_input[751]), .Z(n24799) );
  XOR U24675 ( .A(n24801), .B(n24802), .Z(n24797) );
  AND U24676 ( .A(n24803), .B(n24804), .Z(n24802) );
  XNOR U24677 ( .A(p_input[766]), .B(n24801), .Z(n24804) );
  XOR U24678 ( .A(n24801), .B(p_input[750]), .Z(n24803) );
  XOR U24679 ( .A(n24805), .B(n24806), .Z(n24801) );
  AND U24680 ( .A(n24807), .B(n24808), .Z(n24806) );
  XNOR U24681 ( .A(p_input[765]), .B(n24805), .Z(n24808) );
  XOR U24682 ( .A(n24805), .B(p_input[749]), .Z(n24807) );
  XOR U24683 ( .A(n24809), .B(n24810), .Z(n24805) );
  AND U24684 ( .A(n24811), .B(n24812), .Z(n24810) );
  XNOR U24685 ( .A(p_input[764]), .B(n24809), .Z(n24812) );
  XOR U24686 ( .A(n24809), .B(p_input[748]), .Z(n24811) );
  XOR U24687 ( .A(n24813), .B(n24814), .Z(n24809) );
  AND U24688 ( .A(n24815), .B(n24816), .Z(n24814) );
  XNOR U24689 ( .A(p_input[763]), .B(n24813), .Z(n24816) );
  XOR U24690 ( .A(n24813), .B(p_input[747]), .Z(n24815) );
  XOR U24691 ( .A(n24817), .B(n24818), .Z(n24813) );
  AND U24692 ( .A(n24819), .B(n24820), .Z(n24818) );
  XNOR U24693 ( .A(p_input[762]), .B(n24817), .Z(n24820) );
  XOR U24694 ( .A(n24817), .B(p_input[746]), .Z(n24819) );
  XOR U24695 ( .A(n24821), .B(n24822), .Z(n24817) );
  AND U24696 ( .A(n24823), .B(n24824), .Z(n24822) );
  XNOR U24697 ( .A(p_input[761]), .B(n24821), .Z(n24824) );
  XOR U24698 ( .A(n24821), .B(p_input[745]), .Z(n24823) );
  XOR U24699 ( .A(n24825), .B(n24826), .Z(n24821) );
  AND U24700 ( .A(n24827), .B(n24828), .Z(n24826) );
  XNOR U24701 ( .A(p_input[760]), .B(n24825), .Z(n24828) );
  XOR U24702 ( .A(n24825), .B(p_input[744]), .Z(n24827) );
  XOR U24703 ( .A(n24829), .B(n24830), .Z(n24825) );
  AND U24704 ( .A(n24831), .B(n24832), .Z(n24830) );
  XNOR U24705 ( .A(p_input[759]), .B(n24829), .Z(n24832) );
  XOR U24706 ( .A(n24829), .B(p_input[743]), .Z(n24831) );
  XOR U24707 ( .A(n24833), .B(n24834), .Z(n24829) );
  AND U24708 ( .A(n24835), .B(n24836), .Z(n24834) );
  XNOR U24709 ( .A(p_input[758]), .B(n24833), .Z(n24836) );
  XOR U24710 ( .A(n24833), .B(p_input[742]), .Z(n24835) );
  XOR U24711 ( .A(n24837), .B(n24838), .Z(n24833) );
  AND U24712 ( .A(n24839), .B(n24840), .Z(n24838) );
  XNOR U24713 ( .A(p_input[757]), .B(n24837), .Z(n24840) );
  XOR U24714 ( .A(n24837), .B(p_input[741]), .Z(n24839) );
  XOR U24715 ( .A(n24841), .B(n24842), .Z(n24837) );
  AND U24716 ( .A(n24843), .B(n24844), .Z(n24842) );
  XNOR U24717 ( .A(p_input[756]), .B(n24841), .Z(n24844) );
  XOR U24718 ( .A(n24841), .B(p_input[740]), .Z(n24843) );
  XOR U24719 ( .A(n24845), .B(n24846), .Z(n24841) );
  AND U24720 ( .A(n24847), .B(n24848), .Z(n24846) );
  XNOR U24721 ( .A(p_input[755]), .B(n24845), .Z(n24848) );
  XOR U24722 ( .A(n24845), .B(p_input[739]), .Z(n24847) );
  XOR U24723 ( .A(n24849), .B(n24850), .Z(n24845) );
  AND U24724 ( .A(n24851), .B(n24852), .Z(n24850) );
  XNOR U24725 ( .A(p_input[754]), .B(n24849), .Z(n24852) );
  XOR U24726 ( .A(n24849), .B(p_input[738]), .Z(n24851) );
  XNOR U24727 ( .A(n24853), .B(n24854), .Z(n24849) );
  AND U24728 ( .A(n24855), .B(n24856), .Z(n24854) );
  XOR U24729 ( .A(p_input[753]), .B(n24853), .Z(n24856) );
  XNOR U24730 ( .A(p_input[737]), .B(n24853), .Z(n24855) );
  AND U24731 ( .A(p_input[752]), .B(n24857), .Z(n24853) );
  IV U24732 ( .A(p_input[736]), .Z(n24857) );
  XNOR U24733 ( .A(p_input[704]), .B(n24858), .Z(n24660) );
  AND U24734 ( .A(n885), .B(n24859), .Z(n24858) );
  XOR U24735 ( .A(p_input[720]), .B(p_input[704]), .Z(n24859) );
  XOR U24736 ( .A(n24860), .B(n24861), .Z(n885) );
  AND U24737 ( .A(n24862), .B(n24863), .Z(n24861) );
  XNOR U24738 ( .A(p_input[735]), .B(n24860), .Z(n24863) );
  XOR U24739 ( .A(n24860), .B(p_input[719]), .Z(n24862) );
  XOR U24740 ( .A(n24864), .B(n24865), .Z(n24860) );
  AND U24741 ( .A(n24866), .B(n24867), .Z(n24865) );
  XNOR U24742 ( .A(p_input[734]), .B(n24864), .Z(n24867) );
  XNOR U24743 ( .A(n24864), .B(n24674), .Z(n24866) );
  IV U24744 ( .A(p_input[718]), .Z(n24674) );
  XOR U24745 ( .A(n24868), .B(n24869), .Z(n24864) );
  AND U24746 ( .A(n24870), .B(n24871), .Z(n24869) );
  XNOR U24747 ( .A(p_input[733]), .B(n24868), .Z(n24871) );
  XNOR U24748 ( .A(n24868), .B(n24683), .Z(n24870) );
  IV U24749 ( .A(p_input[717]), .Z(n24683) );
  XOR U24750 ( .A(n24872), .B(n24873), .Z(n24868) );
  AND U24751 ( .A(n24874), .B(n24875), .Z(n24873) );
  XNOR U24752 ( .A(p_input[732]), .B(n24872), .Z(n24875) );
  XNOR U24753 ( .A(n24872), .B(n24692), .Z(n24874) );
  IV U24754 ( .A(p_input[716]), .Z(n24692) );
  XOR U24755 ( .A(n24876), .B(n24877), .Z(n24872) );
  AND U24756 ( .A(n24878), .B(n24879), .Z(n24877) );
  XNOR U24757 ( .A(p_input[731]), .B(n24876), .Z(n24879) );
  XNOR U24758 ( .A(n24876), .B(n24701), .Z(n24878) );
  IV U24759 ( .A(p_input[715]), .Z(n24701) );
  XOR U24760 ( .A(n24880), .B(n24881), .Z(n24876) );
  AND U24761 ( .A(n24882), .B(n24883), .Z(n24881) );
  XNOR U24762 ( .A(p_input[730]), .B(n24880), .Z(n24883) );
  XNOR U24763 ( .A(n24880), .B(n24710), .Z(n24882) );
  IV U24764 ( .A(p_input[714]), .Z(n24710) );
  XOR U24765 ( .A(n24884), .B(n24885), .Z(n24880) );
  AND U24766 ( .A(n24886), .B(n24887), .Z(n24885) );
  XNOR U24767 ( .A(p_input[729]), .B(n24884), .Z(n24887) );
  XNOR U24768 ( .A(n24884), .B(n24719), .Z(n24886) );
  IV U24769 ( .A(p_input[713]), .Z(n24719) );
  XOR U24770 ( .A(n24888), .B(n24889), .Z(n24884) );
  AND U24771 ( .A(n24890), .B(n24891), .Z(n24889) );
  XNOR U24772 ( .A(p_input[728]), .B(n24888), .Z(n24891) );
  XNOR U24773 ( .A(n24888), .B(n24728), .Z(n24890) );
  IV U24774 ( .A(p_input[712]), .Z(n24728) );
  XOR U24775 ( .A(n24892), .B(n24893), .Z(n24888) );
  AND U24776 ( .A(n24894), .B(n24895), .Z(n24893) );
  XNOR U24777 ( .A(p_input[727]), .B(n24892), .Z(n24895) );
  XNOR U24778 ( .A(n24892), .B(n24737), .Z(n24894) );
  IV U24779 ( .A(p_input[711]), .Z(n24737) );
  XOR U24780 ( .A(n24896), .B(n24897), .Z(n24892) );
  AND U24781 ( .A(n24898), .B(n24899), .Z(n24897) );
  XNOR U24782 ( .A(p_input[726]), .B(n24896), .Z(n24899) );
  XNOR U24783 ( .A(n24896), .B(n24746), .Z(n24898) );
  IV U24784 ( .A(p_input[710]), .Z(n24746) );
  XOR U24785 ( .A(n24900), .B(n24901), .Z(n24896) );
  AND U24786 ( .A(n24902), .B(n24903), .Z(n24901) );
  XNOR U24787 ( .A(p_input[725]), .B(n24900), .Z(n24903) );
  XNOR U24788 ( .A(n24900), .B(n24755), .Z(n24902) );
  IV U24789 ( .A(p_input[709]), .Z(n24755) );
  XOR U24790 ( .A(n24904), .B(n24905), .Z(n24900) );
  AND U24791 ( .A(n24906), .B(n24907), .Z(n24905) );
  XNOR U24792 ( .A(p_input[724]), .B(n24904), .Z(n24907) );
  XNOR U24793 ( .A(n24904), .B(n24764), .Z(n24906) );
  IV U24794 ( .A(p_input[708]), .Z(n24764) );
  XOR U24795 ( .A(n24908), .B(n24909), .Z(n24904) );
  AND U24796 ( .A(n24910), .B(n24911), .Z(n24909) );
  XNOR U24797 ( .A(p_input[723]), .B(n24908), .Z(n24911) );
  XNOR U24798 ( .A(n24908), .B(n24773), .Z(n24910) );
  IV U24799 ( .A(p_input[707]), .Z(n24773) );
  XOR U24800 ( .A(n24912), .B(n24913), .Z(n24908) );
  AND U24801 ( .A(n24914), .B(n24915), .Z(n24913) );
  XNOR U24802 ( .A(p_input[722]), .B(n24912), .Z(n24915) );
  XNOR U24803 ( .A(n24912), .B(n24782), .Z(n24914) );
  IV U24804 ( .A(p_input[706]), .Z(n24782) );
  XNOR U24805 ( .A(n24916), .B(n24917), .Z(n24912) );
  AND U24806 ( .A(n24918), .B(n24919), .Z(n24917) );
  XOR U24807 ( .A(p_input[721]), .B(n24916), .Z(n24919) );
  XNOR U24808 ( .A(p_input[705]), .B(n24916), .Z(n24918) );
  AND U24809 ( .A(p_input[720]), .B(n24920), .Z(n24916) );
  IV U24810 ( .A(p_input[704]), .Z(n24920) );
  XOR U24811 ( .A(n24921), .B(n24922), .Z(n24479) );
  AND U24812 ( .A(n553), .B(n24923), .Z(n24922) );
  XNOR U24813 ( .A(n24924), .B(n24921), .Z(n24923) );
  XOR U24814 ( .A(n24925), .B(n24926), .Z(n553) );
  AND U24815 ( .A(n24927), .B(n24928), .Z(n24926) );
  XNOR U24816 ( .A(n24489), .B(n24925), .Z(n24928) );
  AND U24817 ( .A(p_input[703]), .B(p_input[687]), .Z(n24489) );
  XOR U24818 ( .A(n24925), .B(n24490), .Z(n24927) );
  AND U24819 ( .A(p_input[671]), .B(p_input[655]), .Z(n24490) );
  XOR U24820 ( .A(n24929), .B(n24930), .Z(n24925) );
  AND U24821 ( .A(n24931), .B(n24932), .Z(n24930) );
  XOR U24822 ( .A(n24929), .B(n24502), .Z(n24932) );
  XNOR U24823 ( .A(p_input[686]), .B(n24933), .Z(n24502) );
  AND U24824 ( .A(n891), .B(n24934), .Z(n24933) );
  XOR U24825 ( .A(p_input[702]), .B(p_input[686]), .Z(n24934) );
  XNOR U24826 ( .A(n24499), .B(n24929), .Z(n24931) );
  XOR U24827 ( .A(n24935), .B(n24936), .Z(n24499) );
  AND U24828 ( .A(n888), .B(n24937), .Z(n24936) );
  XOR U24829 ( .A(p_input[670]), .B(p_input[654]), .Z(n24937) );
  XOR U24830 ( .A(n24938), .B(n24939), .Z(n24929) );
  AND U24831 ( .A(n24940), .B(n24941), .Z(n24939) );
  XOR U24832 ( .A(n24938), .B(n24514), .Z(n24941) );
  XNOR U24833 ( .A(p_input[685]), .B(n24942), .Z(n24514) );
  AND U24834 ( .A(n891), .B(n24943), .Z(n24942) );
  XOR U24835 ( .A(p_input[701]), .B(p_input[685]), .Z(n24943) );
  XNOR U24836 ( .A(n24511), .B(n24938), .Z(n24940) );
  XOR U24837 ( .A(n24944), .B(n24945), .Z(n24511) );
  AND U24838 ( .A(n888), .B(n24946), .Z(n24945) );
  XOR U24839 ( .A(p_input[669]), .B(p_input[653]), .Z(n24946) );
  XOR U24840 ( .A(n24947), .B(n24948), .Z(n24938) );
  AND U24841 ( .A(n24949), .B(n24950), .Z(n24948) );
  XOR U24842 ( .A(n24947), .B(n24526), .Z(n24950) );
  XNOR U24843 ( .A(p_input[684]), .B(n24951), .Z(n24526) );
  AND U24844 ( .A(n891), .B(n24952), .Z(n24951) );
  XOR U24845 ( .A(p_input[700]), .B(p_input[684]), .Z(n24952) );
  XNOR U24846 ( .A(n24523), .B(n24947), .Z(n24949) );
  XOR U24847 ( .A(n24953), .B(n24954), .Z(n24523) );
  AND U24848 ( .A(n888), .B(n24955), .Z(n24954) );
  XOR U24849 ( .A(p_input[668]), .B(p_input[652]), .Z(n24955) );
  XOR U24850 ( .A(n24956), .B(n24957), .Z(n24947) );
  AND U24851 ( .A(n24958), .B(n24959), .Z(n24957) );
  XOR U24852 ( .A(n24956), .B(n24538), .Z(n24959) );
  XNOR U24853 ( .A(p_input[683]), .B(n24960), .Z(n24538) );
  AND U24854 ( .A(n891), .B(n24961), .Z(n24960) );
  XOR U24855 ( .A(p_input[699]), .B(p_input[683]), .Z(n24961) );
  XNOR U24856 ( .A(n24535), .B(n24956), .Z(n24958) );
  XOR U24857 ( .A(n24962), .B(n24963), .Z(n24535) );
  AND U24858 ( .A(n888), .B(n24964), .Z(n24963) );
  XOR U24859 ( .A(p_input[667]), .B(p_input[651]), .Z(n24964) );
  XOR U24860 ( .A(n24965), .B(n24966), .Z(n24956) );
  AND U24861 ( .A(n24967), .B(n24968), .Z(n24966) );
  XOR U24862 ( .A(n24965), .B(n24550), .Z(n24968) );
  XNOR U24863 ( .A(p_input[682]), .B(n24969), .Z(n24550) );
  AND U24864 ( .A(n891), .B(n24970), .Z(n24969) );
  XOR U24865 ( .A(p_input[698]), .B(p_input[682]), .Z(n24970) );
  XNOR U24866 ( .A(n24547), .B(n24965), .Z(n24967) );
  XOR U24867 ( .A(n24971), .B(n24972), .Z(n24547) );
  AND U24868 ( .A(n888), .B(n24973), .Z(n24972) );
  XOR U24869 ( .A(p_input[666]), .B(p_input[650]), .Z(n24973) );
  XOR U24870 ( .A(n24974), .B(n24975), .Z(n24965) );
  AND U24871 ( .A(n24976), .B(n24977), .Z(n24975) );
  XOR U24872 ( .A(n24974), .B(n24562), .Z(n24977) );
  XNOR U24873 ( .A(p_input[681]), .B(n24978), .Z(n24562) );
  AND U24874 ( .A(n891), .B(n24979), .Z(n24978) );
  XOR U24875 ( .A(p_input[697]), .B(p_input[681]), .Z(n24979) );
  XNOR U24876 ( .A(n24559), .B(n24974), .Z(n24976) );
  XOR U24877 ( .A(n24980), .B(n24981), .Z(n24559) );
  AND U24878 ( .A(n888), .B(n24982), .Z(n24981) );
  XOR U24879 ( .A(p_input[665]), .B(p_input[649]), .Z(n24982) );
  XOR U24880 ( .A(n24983), .B(n24984), .Z(n24974) );
  AND U24881 ( .A(n24985), .B(n24986), .Z(n24984) );
  XOR U24882 ( .A(n24983), .B(n24574), .Z(n24986) );
  XNOR U24883 ( .A(p_input[680]), .B(n24987), .Z(n24574) );
  AND U24884 ( .A(n891), .B(n24988), .Z(n24987) );
  XOR U24885 ( .A(p_input[696]), .B(p_input[680]), .Z(n24988) );
  XNOR U24886 ( .A(n24571), .B(n24983), .Z(n24985) );
  XOR U24887 ( .A(n24989), .B(n24990), .Z(n24571) );
  AND U24888 ( .A(n888), .B(n24991), .Z(n24990) );
  XOR U24889 ( .A(p_input[664]), .B(p_input[648]), .Z(n24991) );
  XOR U24890 ( .A(n24992), .B(n24993), .Z(n24983) );
  AND U24891 ( .A(n24994), .B(n24995), .Z(n24993) );
  XOR U24892 ( .A(n24992), .B(n24586), .Z(n24995) );
  XNOR U24893 ( .A(p_input[679]), .B(n24996), .Z(n24586) );
  AND U24894 ( .A(n891), .B(n24997), .Z(n24996) );
  XOR U24895 ( .A(p_input[695]), .B(p_input[679]), .Z(n24997) );
  XNOR U24896 ( .A(n24583), .B(n24992), .Z(n24994) );
  XOR U24897 ( .A(n24998), .B(n24999), .Z(n24583) );
  AND U24898 ( .A(n888), .B(n25000), .Z(n24999) );
  XOR U24899 ( .A(p_input[663]), .B(p_input[647]), .Z(n25000) );
  XOR U24900 ( .A(n25001), .B(n25002), .Z(n24992) );
  AND U24901 ( .A(n25003), .B(n25004), .Z(n25002) );
  XOR U24902 ( .A(n25001), .B(n24598), .Z(n25004) );
  XNOR U24903 ( .A(p_input[678]), .B(n25005), .Z(n24598) );
  AND U24904 ( .A(n891), .B(n25006), .Z(n25005) );
  XOR U24905 ( .A(p_input[694]), .B(p_input[678]), .Z(n25006) );
  XNOR U24906 ( .A(n24595), .B(n25001), .Z(n25003) );
  XOR U24907 ( .A(n25007), .B(n25008), .Z(n24595) );
  AND U24908 ( .A(n888), .B(n25009), .Z(n25008) );
  XOR U24909 ( .A(p_input[662]), .B(p_input[646]), .Z(n25009) );
  XOR U24910 ( .A(n25010), .B(n25011), .Z(n25001) );
  AND U24911 ( .A(n25012), .B(n25013), .Z(n25011) );
  XOR U24912 ( .A(n25010), .B(n24610), .Z(n25013) );
  XNOR U24913 ( .A(p_input[677]), .B(n25014), .Z(n24610) );
  AND U24914 ( .A(n891), .B(n25015), .Z(n25014) );
  XOR U24915 ( .A(p_input[693]), .B(p_input[677]), .Z(n25015) );
  XNOR U24916 ( .A(n24607), .B(n25010), .Z(n25012) );
  XOR U24917 ( .A(n25016), .B(n25017), .Z(n24607) );
  AND U24918 ( .A(n888), .B(n25018), .Z(n25017) );
  XOR U24919 ( .A(p_input[661]), .B(p_input[645]), .Z(n25018) );
  XOR U24920 ( .A(n25019), .B(n25020), .Z(n25010) );
  AND U24921 ( .A(n25021), .B(n25022), .Z(n25020) );
  XOR U24922 ( .A(n25019), .B(n24622), .Z(n25022) );
  XNOR U24923 ( .A(p_input[676]), .B(n25023), .Z(n24622) );
  AND U24924 ( .A(n891), .B(n25024), .Z(n25023) );
  XOR U24925 ( .A(p_input[692]), .B(p_input[676]), .Z(n25024) );
  XNOR U24926 ( .A(n24619), .B(n25019), .Z(n25021) );
  XOR U24927 ( .A(n25025), .B(n25026), .Z(n24619) );
  AND U24928 ( .A(n888), .B(n25027), .Z(n25026) );
  XOR U24929 ( .A(p_input[660]), .B(p_input[644]), .Z(n25027) );
  XOR U24930 ( .A(n25028), .B(n25029), .Z(n25019) );
  AND U24931 ( .A(n25030), .B(n25031), .Z(n25029) );
  XOR U24932 ( .A(n25028), .B(n24634), .Z(n25031) );
  XNOR U24933 ( .A(p_input[675]), .B(n25032), .Z(n24634) );
  AND U24934 ( .A(n891), .B(n25033), .Z(n25032) );
  XOR U24935 ( .A(p_input[691]), .B(p_input[675]), .Z(n25033) );
  XNOR U24936 ( .A(n24631), .B(n25028), .Z(n25030) );
  XOR U24937 ( .A(n25034), .B(n25035), .Z(n24631) );
  AND U24938 ( .A(n888), .B(n25036), .Z(n25035) );
  XOR U24939 ( .A(p_input[659]), .B(p_input[643]), .Z(n25036) );
  XOR U24940 ( .A(n25037), .B(n25038), .Z(n25028) );
  AND U24941 ( .A(n25039), .B(n25040), .Z(n25038) );
  XOR U24942 ( .A(n25037), .B(n24646), .Z(n25040) );
  XNOR U24943 ( .A(p_input[674]), .B(n25041), .Z(n24646) );
  AND U24944 ( .A(n891), .B(n25042), .Z(n25041) );
  XOR U24945 ( .A(p_input[690]), .B(p_input[674]), .Z(n25042) );
  XNOR U24946 ( .A(n24643), .B(n25037), .Z(n25039) );
  XOR U24947 ( .A(n25043), .B(n25044), .Z(n24643) );
  AND U24948 ( .A(n888), .B(n25045), .Z(n25044) );
  XOR U24949 ( .A(p_input[658]), .B(p_input[642]), .Z(n25045) );
  XOR U24950 ( .A(n25046), .B(n25047), .Z(n25037) );
  AND U24951 ( .A(n25048), .B(n25049), .Z(n25047) );
  XNOR U24952 ( .A(n25050), .B(n24659), .Z(n25049) );
  XNOR U24953 ( .A(p_input[673]), .B(n25051), .Z(n24659) );
  AND U24954 ( .A(n891), .B(n25052), .Z(n25051) );
  XNOR U24955 ( .A(p_input[689]), .B(n25053), .Z(n25052) );
  IV U24956 ( .A(p_input[673]), .Z(n25053) );
  XNOR U24957 ( .A(n24656), .B(n25046), .Z(n25048) );
  XNOR U24958 ( .A(p_input[641]), .B(n25054), .Z(n24656) );
  AND U24959 ( .A(n888), .B(n25055), .Z(n25054) );
  XOR U24960 ( .A(p_input[657]), .B(p_input[641]), .Z(n25055) );
  IV U24961 ( .A(n25050), .Z(n25046) );
  AND U24962 ( .A(n24921), .B(n24924), .Z(n25050) );
  XOR U24963 ( .A(p_input[672]), .B(n25056), .Z(n24924) );
  AND U24964 ( .A(n891), .B(n25057), .Z(n25056) );
  XOR U24965 ( .A(p_input[688]), .B(p_input[672]), .Z(n25057) );
  XOR U24966 ( .A(n25058), .B(n25059), .Z(n891) );
  AND U24967 ( .A(n25060), .B(n25061), .Z(n25059) );
  XNOR U24968 ( .A(p_input[703]), .B(n25058), .Z(n25061) );
  XOR U24969 ( .A(n25058), .B(p_input[687]), .Z(n25060) );
  XOR U24970 ( .A(n25062), .B(n25063), .Z(n25058) );
  AND U24971 ( .A(n25064), .B(n25065), .Z(n25063) );
  XNOR U24972 ( .A(p_input[702]), .B(n25062), .Z(n25065) );
  XOR U24973 ( .A(n25062), .B(p_input[686]), .Z(n25064) );
  XOR U24974 ( .A(n25066), .B(n25067), .Z(n25062) );
  AND U24975 ( .A(n25068), .B(n25069), .Z(n25067) );
  XNOR U24976 ( .A(p_input[701]), .B(n25066), .Z(n25069) );
  XOR U24977 ( .A(n25066), .B(p_input[685]), .Z(n25068) );
  XOR U24978 ( .A(n25070), .B(n25071), .Z(n25066) );
  AND U24979 ( .A(n25072), .B(n25073), .Z(n25071) );
  XNOR U24980 ( .A(p_input[700]), .B(n25070), .Z(n25073) );
  XOR U24981 ( .A(n25070), .B(p_input[684]), .Z(n25072) );
  XOR U24982 ( .A(n25074), .B(n25075), .Z(n25070) );
  AND U24983 ( .A(n25076), .B(n25077), .Z(n25075) );
  XNOR U24984 ( .A(p_input[699]), .B(n25074), .Z(n25077) );
  XOR U24985 ( .A(n25074), .B(p_input[683]), .Z(n25076) );
  XOR U24986 ( .A(n25078), .B(n25079), .Z(n25074) );
  AND U24987 ( .A(n25080), .B(n25081), .Z(n25079) );
  XNOR U24988 ( .A(p_input[698]), .B(n25078), .Z(n25081) );
  XOR U24989 ( .A(n25078), .B(p_input[682]), .Z(n25080) );
  XOR U24990 ( .A(n25082), .B(n25083), .Z(n25078) );
  AND U24991 ( .A(n25084), .B(n25085), .Z(n25083) );
  XNOR U24992 ( .A(p_input[697]), .B(n25082), .Z(n25085) );
  XOR U24993 ( .A(n25082), .B(p_input[681]), .Z(n25084) );
  XOR U24994 ( .A(n25086), .B(n25087), .Z(n25082) );
  AND U24995 ( .A(n25088), .B(n25089), .Z(n25087) );
  XNOR U24996 ( .A(p_input[696]), .B(n25086), .Z(n25089) );
  XOR U24997 ( .A(n25086), .B(p_input[680]), .Z(n25088) );
  XOR U24998 ( .A(n25090), .B(n25091), .Z(n25086) );
  AND U24999 ( .A(n25092), .B(n25093), .Z(n25091) );
  XNOR U25000 ( .A(p_input[695]), .B(n25090), .Z(n25093) );
  XOR U25001 ( .A(n25090), .B(p_input[679]), .Z(n25092) );
  XOR U25002 ( .A(n25094), .B(n25095), .Z(n25090) );
  AND U25003 ( .A(n25096), .B(n25097), .Z(n25095) );
  XNOR U25004 ( .A(p_input[694]), .B(n25094), .Z(n25097) );
  XOR U25005 ( .A(n25094), .B(p_input[678]), .Z(n25096) );
  XOR U25006 ( .A(n25098), .B(n25099), .Z(n25094) );
  AND U25007 ( .A(n25100), .B(n25101), .Z(n25099) );
  XNOR U25008 ( .A(p_input[693]), .B(n25098), .Z(n25101) );
  XOR U25009 ( .A(n25098), .B(p_input[677]), .Z(n25100) );
  XOR U25010 ( .A(n25102), .B(n25103), .Z(n25098) );
  AND U25011 ( .A(n25104), .B(n25105), .Z(n25103) );
  XNOR U25012 ( .A(p_input[692]), .B(n25102), .Z(n25105) );
  XOR U25013 ( .A(n25102), .B(p_input[676]), .Z(n25104) );
  XOR U25014 ( .A(n25106), .B(n25107), .Z(n25102) );
  AND U25015 ( .A(n25108), .B(n25109), .Z(n25107) );
  XNOR U25016 ( .A(p_input[691]), .B(n25106), .Z(n25109) );
  XOR U25017 ( .A(n25106), .B(p_input[675]), .Z(n25108) );
  XOR U25018 ( .A(n25110), .B(n25111), .Z(n25106) );
  AND U25019 ( .A(n25112), .B(n25113), .Z(n25111) );
  XNOR U25020 ( .A(p_input[690]), .B(n25110), .Z(n25113) );
  XOR U25021 ( .A(n25110), .B(p_input[674]), .Z(n25112) );
  XNOR U25022 ( .A(n25114), .B(n25115), .Z(n25110) );
  AND U25023 ( .A(n25116), .B(n25117), .Z(n25115) );
  XOR U25024 ( .A(p_input[689]), .B(n25114), .Z(n25117) );
  XNOR U25025 ( .A(p_input[673]), .B(n25114), .Z(n25116) );
  AND U25026 ( .A(p_input[688]), .B(n25118), .Z(n25114) );
  IV U25027 ( .A(p_input[672]), .Z(n25118) );
  XNOR U25028 ( .A(p_input[640]), .B(n25119), .Z(n24921) );
  AND U25029 ( .A(n888), .B(n25120), .Z(n25119) );
  XOR U25030 ( .A(p_input[656]), .B(p_input[640]), .Z(n25120) );
  XOR U25031 ( .A(n25121), .B(n25122), .Z(n888) );
  AND U25032 ( .A(n25123), .B(n25124), .Z(n25122) );
  XNOR U25033 ( .A(p_input[671]), .B(n25121), .Z(n25124) );
  XOR U25034 ( .A(n25121), .B(p_input[655]), .Z(n25123) );
  XOR U25035 ( .A(n25125), .B(n25126), .Z(n25121) );
  AND U25036 ( .A(n25127), .B(n25128), .Z(n25126) );
  XNOR U25037 ( .A(p_input[670]), .B(n25125), .Z(n25128) );
  XNOR U25038 ( .A(n25125), .B(n24935), .Z(n25127) );
  IV U25039 ( .A(p_input[654]), .Z(n24935) );
  XOR U25040 ( .A(n25129), .B(n25130), .Z(n25125) );
  AND U25041 ( .A(n25131), .B(n25132), .Z(n25130) );
  XNOR U25042 ( .A(p_input[669]), .B(n25129), .Z(n25132) );
  XNOR U25043 ( .A(n25129), .B(n24944), .Z(n25131) );
  IV U25044 ( .A(p_input[653]), .Z(n24944) );
  XOR U25045 ( .A(n25133), .B(n25134), .Z(n25129) );
  AND U25046 ( .A(n25135), .B(n25136), .Z(n25134) );
  XNOR U25047 ( .A(p_input[668]), .B(n25133), .Z(n25136) );
  XNOR U25048 ( .A(n25133), .B(n24953), .Z(n25135) );
  IV U25049 ( .A(p_input[652]), .Z(n24953) );
  XOR U25050 ( .A(n25137), .B(n25138), .Z(n25133) );
  AND U25051 ( .A(n25139), .B(n25140), .Z(n25138) );
  XNOR U25052 ( .A(p_input[667]), .B(n25137), .Z(n25140) );
  XNOR U25053 ( .A(n25137), .B(n24962), .Z(n25139) );
  IV U25054 ( .A(p_input[651]), .Z(n24962) );
  XOR U25055 ( .A(n25141), .B(n25142), .Z(n25137) );
  AND U25056 ( .A(n25143), .B(n25144), .Z(n25142) );
  XNOR U25057 ( .A(p_input[666]), .B(n25141), .Z(n25144) );
  XNOR U25058 ( .A(n25141), .B(n24971), .Z(n25143) );
  IV U25059 ( .A(p_input[650]), .Z(n24971) );
  XOR U25060 ( .A(n25145), .B(n25146), .Z(n25141) );
  AND U25061 ( .A(n25147), .B(n25148), .Z(n25146) );
  XNOR U25062 ( .A(p_input[665]), .B(n25145), .Z(n25148) );
  XNOR U25063 ( .A(n25145), .B(n24980), .Z(n25147) );
  IV U25064 ( .A(p_input[649]), .Z(n24980) );
  XOR U25065 ( .A(n25149), .B(n25150), .Z(n25145) );
  AND U25066 ( .A(n25151), .B(n25152), .Z(n25150) );
  XNOR U25067 ( .A(p_input[664]), .B(n25149), .Z(n25152) );
  XNOR U25068 ( .A(n25149), .B(n24989), .Z(n25151) );
  IV U25069 ( .A(p_input[648]), .Z(n24989) );
  XOR U25070 ( .A(n25153), .B(n25154), .Z(n25149) );
  AND U25071 ( .A(n25155), .B(n25156), .Z(n25154) );
  XNOR U25072 ( .A(p_input[663]), .B(n25153), .Z(n25156) );
  XNOR U25073 ( .A(n25153), .B(n24998), .Z(n25155) );
  IV U25074 ( .A(p_input[647]), .Z(n24998) );
  XOR U25075 ( .A(n25157), .B(n25158), .Z(n25153) );
  AND U25076 ( .A(n25159), .B(n25160), .Z(n25158) );
  XNOR U25077 ( .A(p_input[662]), .B(n25157), .Z(n25160) );
  XNOR U25078 ( .A(n25157), .B(n25007), .Z(n25159) );
  IV U25079 ( .A(p_input[646]), .Z(n25007) );
  XOR U25080 ( .A(n25161), .B(n25162), .Z(n25157) );
  AND U25081 ( .A(n25163), .B(n25164), .Z(n25162) );
  XNOR U25082 ( .A(p_input[661]), .B(n25161), .Z(n25164) );
  XNOR U25083 ( .A(n25161), .B(n25016), .Z(n25163) );
  IV U25084 ( .A(p_input[645]), .Z(n25016) );
  XOR U25085 ( .A(n25165), .B(n25166), .Z(n25161) );
  AND U25086 ( .A(n25167), .B(n25168), .Z(n25166) );
  XNOR U25087 ( .A(p_input[660]), .B(n25165), .Z(n25168) );
  XNOR U25088 ( .A(n25165), .B(n25025), .Z(n25167) );
  IV U25089 ( .A(p_input[644]), .Z(n25025) );
  XOR U25090 ( .A(n25169), .B(n25170), .Z(n25165) );
  AND U25091 ( .A(n25171), .B(n25172), .Z(n25170) );
  XNOR U25092 ( .A(p_input[659]), .B(n25169), .Z(n25172) );
  XNOR U25093 ( .A(n25169), .B(n25034), .Z(n25171) );
  IV U25094 ( .A(p_input[643]), .Z(n25034) );
  XOR U25095 ( .A(n25173), .B(n25174), .Z(n25169) );
  AND U25096 ( .A(n25175), .B(n25176), .Z(n25174) );
  XNOR U25097 ( .A(p_input[658]), .B(n25173), .Z(n25176) );
  XNOR U25098 ( .A(n25173), .B(n25043), .Z(n25175) );
  IV U25099 ( .A(p_input[642]), .Z(n25043) );
  XNOR U25100 ( .A(n25177), .B(n25178), .Z(n25173) );
  AND U25101 ( .A(n25179), .B(n25180), .Z(n25178) );
  XOR U25102 ( .A(p_input[657]), .B(n25177), .Z(n25180) );
  XNOR U25103 ( .A(p_input[641]), .B(n25177), .Z(n25179) );
  AND U25104 ( .A(p_input[656]), .B(n25181), .Z(n25177) );
  IV U25105 ( .A(p_input[640]), .Z(n25181) );
  XOR U25106 ( .A(n25182), .B(n25183), .Z(n24297) );
  AND U25107 ( .A(n824), .B(n25184), .Z(n25183) );
  XNOR U25108 ( .A(n25185), .B(n25182), .Z(n25184) );
  XOR U25109 ( .A(n25186), .B(n25187), .Z(n824) );
  AND U25110 ( .A(n25188), .B(n25189), .Z(n25187) );
  XNOR U25111 ( .A(n24309), .B(n25186), .Z(n25189) );
  AND U25112 ( .A(n25190), .B(n25191), .Z(n24309) );
  XOR U25113 ( .A(n25186), .B(n24308), .Z(n25188) );
  AND U25114 ( .A(n25192), .B(n25193), .Z(n24308) );
  XOR U25115 ( .A(n25194), .B(n25195), .Z(n25186) );
  AND U25116 ( .A(n25196), .B(n25197), .Z(n25195) );
  XOR U25117 ( .A(n25194), .B(n24321), .Z(n25197) );
  XOR U25118 ( .A(n25198), .B(n25199), .Z(n24321) );
  AND U25119 ( .A(n559), .B(n25200), .Z(n25199) );
  XOR U25120 ( .A(n25201), .B(n25198), .Z(n25200) );
  XNOR U25121 ( .A(n24318), .B(n25194), .Z(n25196) );
  XOR U25122 ( .A(n25202), .B(n25203), .Z(n24318) );
  AND U25123 ( .A(n556), .B(n25204), .Z(n25203) );
  XOR U25124 ( .A(n25205), .B(n25202), .Z(n25204) );
  XOR U25125 ( .A(n25206), .B(n25207), .Z(n25194) );
  AND U25126 ( .A(n25208), .B(n25209), .Z(n25207) );
  XOR U25127 ( .A(n25206), .B(n24333), .Z(n25209) );
  XOR U25128 ( .A(n25210), .B(n25211), .Z(n24333) );
  AND U25129 ( .A(n559), .B(n25212), .Z(n25211) );
  XOR U25130 ( .A(n25213), .B(n25210), .Z(n25212) );
  XNOR U25131 ( .A(n24330), .B(n25206), .Z(n25208) );
  XOR U25132 ( .A(n25214), .B(n25215), .Z(n24330) );
  AND U25133 ( .A(n556), .B(n25216), .Z(n25215) );
  XOR U25134 ( .A(n25217), .B(n25214), .Z(n25216) );
  XOR U25135 ( .A(n25218), .B(n25219), .Z(n25206) );
  AND U25136 ( .A(n25220), .B(n25221), .Z(n25219) );
  XOR U25137 ( .A(n25218), .B(n24345), .Z(n25221) );
  XOR U25138 ( .A(n25222), .B(n25223), .Z(n24345) );
  AND U25139 ( .A(n559), .B(n25224), .Z(n25223) );
  XOR U25140 ( .A(n25225), .B(n25222), .Z(n25224) );
  XNOR U25141 ( .A(n24342), .B(n25218), .Z(n25220) );
  XOR U25142 ( .A(n25226), .B(n25227), .Z(n24342) );
  AND U25143 ( .A(n556), .B(n25228), .Z(n25227) );
  XOR U25144 ( .A(n25229), .B(n25226), .Z(n25228) );
  XOR U25145 ( .A(n25230), .B(n25231), .Z(n25218) );
  AND U25146 ( .A(n25232), .B(n25233), .Z(n25231) );
  XOR U25147 ( .A(n25230), .B(n24357), .Z(n25233) );
  XOR U25148 ( .A(n25234), .B(n25235), .Z(n24357) );
  AND U25149 ( .A(n559), .B(n25236), .Z(n25235) );
  XOR U25150 ( .A(n25237), .B(n25234), .Z(n25236) );
  XNOR U25151 ( .A(n24354), .B(n25230), .Z(n25232) );
  XOR U25152 ( .A(n25238), .B(n25239), .Z(n24354) );
  AND U25153 ( .A(n556), .B(n25240), .Z(n25239) );
  XOR U25154 ( .A(n25241), .B(n25238), .Z(n25240) );
  XOR U25155 ( .A(n25242), .B(n25243), .Z(n25230) );
  AND U25156 ( .A(n25244), .B(n25245), .Z(n25243) );
  XOR U25157 ( .A(n25242), .B(n24369), .Z(n25245) );
  XOR U25158 ( .A(n25246), .B(n25247), .Z(n24369) );
  AND U25159 ( .A(n559), .B(n25248), .Z(n25247) );
  XOR U25160 ( .A(n25249), .B(n25246), .Z(n25248) );
  XNOR U25161 ( .A(n24366), .B(n25242), .Z(n25244) );
  XOR U25162 ( .A(n25250), .B(n25251), .Z(n24366) );
  AND U25163 ( .A(n556), .B(n25252), .Z(n25251) );
  XOR U25164 ( .A(n25253), .B(n25250), .Z(n25252) );
  XOR U25165 ( .A(n25254), .B(n25255), .Z(n25242) );
  AND U25166 ( .A(n25256), .B(n25257), .Z(n25255) );
  XOR U25167 ( .A(n25254), .B(n24381), .Z(n25257) );
  XOR U25168 ( .A(n25258), .B(n25259), .Z(n24381) );
  AND U25169 ( .A(n559), .B(n25260), .Z(n25259) );
  XOR U25170 ( .A(n25261), .B(n25258), .Z(n25260) );
  XNOR U25171 ( .A(n24378), .B(n25254), .Z(n25256) );
  XOR U25172 ( .A(n25262), .B(n25263), .Z(n24378) );
  AND U25173 ( .A(n556), .B(n25264), .Z(n25263) );
  XOR U25174 ( .A(n25265), .B(n25262), .Z(n25264) );
  XOR U25175 ( .A(n25266), .B(n25267), .Z(n25254) );
  AND U25176 ( .A(n25268), .B(n25269), .Z(n25267) );
  XOR U25177 ( .A(n25266), .B(n24393), .Z(n25269) );
  XOR U25178 ( .A(n25270), .B(n25271), .Z(n24393) );
  AND U25179 ( .A(n559), .B(n25272), .Z(n25271) );
  XOR U25180 ( .A(n25273), .B(n25270), .Z(n25272) );
  XNOR U25181 ( .A(n24390), .B(n25266), .Z(n25268) );
  XOR U25182 ( .A(n25274), .B(n25275), .Z(n24390) );
  AND U25183 ( .A(n556), .B(n25276), .Z(n25275) );
  XOR U25184 ( .A(n25277), .B(n25274), .Z(n25276) );
  XOR U25185 ( .A(n25278), .B(n25279), .Z(n25266) );
  AND U25186 ( .A(n25280), .B(n25281), .Z(n25279) );
  XOR U25187 ( .A(n25278), .B(n24405), .Z(n25281) );
  XOR U25188 ( .A(n25282), .B(n25283), .Z(n24405) );
  AND U25189 ( .A(n559), .B(n25284), .Z(n25283) );
  XOR U25190 ( .A(n25285), .B(n25282), .Z(n25284) );
  XNOR U25191 ( .A(n24402), .B(n25278), .Z(n25280) );
  XOR U25192 ( .A(n25286), .B(n25287), .Z(n24402) );
  AND U25193 ( .A(n556), .B(n25288), .Z(n25287) );
  XOR U25194 ( .A(n25289), .B(n25286), .Z(n25288) );
  XOR U25195 ( .A(n25290), .B(n25291), .Z(n25278) );
  AND U25196 ( .A(n25292), .B(n25293), .Z(n25291) );
  XOR U25197 ( .A(n25290), .B(n24417), .Z(n25293) );
  XOR U25198 ( .A(n25294), .B(n25295), .Z(n24417) );
  AND U25199 ( .A(n559), .B(n25296), .Z(n25295) );
  XOR U25200 ( .A(n25297), .B(n25294), .Z(n25296) );
  XNOR U25201 ( .A(n24414), .B(n25290), .Z(n25292) );
  XOR U25202 ( .A(n25298), .B(n25299), .Z(n24414) );
  AND U25203 ( .A(n556), .B(n25300), .Z(n25299) );
  XOR U25204 ( .A(n25301), .B(n25298), .Z(n25300) );
  XOR U25205 ( .A(n25302), .B(n25303), .Z(n25290) );
  AND U25206 ( .A(n25304), .B(n25305), .Z(n25303) );
  XOR U25207 ( .A(n25302), .B(n24429), .Z(n25305) );
  XOR U25208 ( .A(n25306), .B(n25307), .Z(n24429) );
  AND U25209 ( .A(n559), .B(n25308), .Z(n25307) );
  XOR U25210 ( .A(n25309), .B(n25306), .Z(n25308) );
  XNOR U25211 ( .A(n24426), .B(n25302), .Z(n25304) );
  XOR U25212 ( .A(n25310), .B(n25311), .Z(n24426) );
  AND U25213 ( .A(n556), .B(n25312), .Z(n25311) );
  XOR U25214 ( .A(n25313), .B(n25310), .Z(n25312) );
  XOR U25215 ( .A(n25314), .B(n25315), .Z(n25302) );
  AND U25216 ( .A(n25316), .B(n25317), .Z(n25315) );
  XOR U25217 ( .A(n25314), .B(n24441), .Z(n25317) );
  XOR U25218 ( .A(n25318), .B(n25319), .Z(n24441) );
  AND U25219 ( .A(n559), .B(n25320), .Z(n25319) );
  XOR U25220 ( .A(n25321), .B(n25318), .Z(n25320) );
  XNOR U25221 ( .A(n24438), .B(n25314), .Z(n25316) );
  XOR U25222 ( .A(n25322), .B(n25323), .Z(n24438) );
  AND U25223 ( .A(n556), .B(n25324), .Z(n25323) );
  XOR U25224 ( .A(n25325), .B(n25322), .Z(n25324) );
  XOR U25225 ( .A(n25326), .B(n25327), .Z(n25314) );
  AND U25226 ( .A(n25328), .B(n25329), .Z(n25327) );
  XOR U25227 ( .A(n25326), .B(n24453), .Z(n25329) );
  XOR U25228 ( .A(n25330), .B(n25331), .Z(n24453) );
  AND U25229 ( .A(n559), .B(n25332), .Z(n25331) );
  XOR U25230 ( .A(n25333), .B(n25330), .Z(n25332) );
  XNOR U25231 ( .A(n24450), .B(n25326), .Z(n25328) );
  XOR U25232 ( .A(n25334), .B(n25335), .Z(n24450) );
  AND U25233 ( .A(n556), .B(n25336), .Z(n25335) );
  XOR U25234 ( .A(n25337), .B(n25334), .Z(n25336) );
  XOR U25235 ( .A(n25338), .B(n25339), .Z(n25326) );
  AND U25236 ( .A(n25340), .B(n25341), .Z(n25339) );
  XOR U25237 ( .A(n25338), .B(n24465), .Z(n25341) );
  XOR U25238 ( .A(n25342), .B(n25343), .Z(n24465) );
  AND U25239 ( .A(n559), .B(n25344), .Z(n25343) );
  XOR U25240 ( .A(n25345), .B(n25342), .Z(n25344) );
  XNOR U25241 ( .A(n24462), .B(n25338), .Z(n25340) );
  XOR U25242 ( .A(n25346), .B(n25347), .Z(n24462) );
  AND U25243 ( .A(n556), .B(n25348), .Z(n25347) );
  XOR U25244 ( .A(n25349), .B(n25346), .Z(n25348) );
  XOR U25245 ( .A(n25350), .B(n25351), .Z(n25338) );
  AND U25246 ( .A(n25352), .B(n25353), .Z(n25351) );
  XNOR U25247 ( .A(n25354), .B(n24478), .Z(n25353) );
  XOR U25248 ( .A(n25355), .B(n25356), .Z(n24478) );
  AND U25249 ( .A(n559), .B(n25357), .Z(n25356) );
  XOR U25250 ( .A(n25355), .B(n25358), .Z(n25357) );
  XNOR U25251 ( .A(n24475), .B(n25350), .Z(n25352) );
  XOR U25252 ( .A(n25359), .B(n25360), .Z(n24475) );
  AND U25253 ( .A(n556), .B(n25361), .Z(n25360) );
  XOR U25254 ( .A(n25359), .B(n25362), .Z(n25361) );
  IV U25255 ( .A(n25354), .Z(n25350) );
  AND U25256 ( .A(n25182), .B(n25185), .Z(n25354) );
  XNOR U25257 ( .A(n25363), .B(n25364), .Z(n25185) );
  AND U25258 ( .A(n559), .B(n25365), .Z(n25364) );
  XNOR U25259 ( .A(n25366), .B(n25363), .Z(n25365) );
  XOR U25260 ( .A(n25367), .B(n25368), .Z(n559) );
  AND U25261 ( .A(n25369), .B(n25370), .Z(n25368) );
  XNOR U25262 ( .A(n25190), .B(n25367), .Z(n25370) );
  AND U25263 ( .A(p_input[639]), .B(p_input[623]), .Z(n25190) );
  XOR U25264 ( .A(n25367), .B(n25191), .Z(n25369) );
  AND U25265 ( .A(p_input[607]), .B(p_input[591]), .Z(n25191) );
  XOR U25266 ( .A(n25371), .B(n25372), .Z(n25367) );
  AND U25267 ( .A(n25373), .B(n25374), .Z(n25372) );
  XOR U25268 ( .A(n25371), .B(n25201), .Z(n25374) );
  XNOR U25269 ( .A(p_input[622]), .B(n25375), .Z(n25201) );
  AND U25270 ( .A(n899), .B(n25376), .Z(n25375) );
  XOR U25271 ( .A(p_input[638]), .B(p_input[622]), .Z(n25376) );
  XNOR U25272 ( .A(n25198), .B(n25371), .Z(n25373) );
  XOR U25273 ( .A(n25377), .B(n25378), .Z(n25198) );
  AND U25274 ( .A(n897), .B(n25379), .Z(n25378) );
  XOR U25275 ( .A(p_input[606]), .B(p_input[590]), .Z(n25379) );
  XOR U25276 ( .A(n25380), .B(n25381), .Z(n25371) );
  AND U25277 ( .A(n25382), .B(n25383), .Z(n25381) );
  XOR U25278 ( .A(n25380), .B(n25213), .Z(n25383) );
  XNOR U25279 ( .A(p_input[621]), .B(n25384), .Z(n25213) );
  AND U25280 ( .A(n899), .B(n25385), .Z(n25384) );
  XOR U25281 ( .A(p_input[637]), .B(p_input[621]), .Z(n25385) );
  XNOR U25282 ( .A(n25210), .B(n25380), .Z(n25382) );
  XOR U25283 ( .A(n25386), .B(n25387), .Z(n25210) );
  AND U25284 ( .A(n897), .B(n25388), .Z(n25387) );
  XOR U25285 ( .A(p_input[605]), .B(p_input[589]), .Z(n25388) );
  XOR U25286 ( .A(n25389), .B(n25390), .Z(n25380) );
  AND U25287 ( .A(n25391), .B(n25392), .Z(n25390) );
  XOR U25288 ( .A(n25389), .B(n25225), .Z(n25392) );
  XNOR U25289 ( .A(p_input[620]), .B(n25393), .Z(n25225) );
  AND U25290 ( .A(n899), .B(n25394), .Z(n25393) );
  XOR U25291 ( .A(p_input[636]), .B(p_input[620]), .Z(n25394) );
  XNOR U25292 ( .A(n25222), .B(n25389), .Z(n25391) );
  XOR U25293 ( .A(n25395), .B(n25396), .Z(n25222) );
  AND U25294 ( .A(n897), .B(n25397), .Z(n25396) );
  XOR U25295 ( .A(p_input[604]), .B(p_input[588]), .Z(n25397) );
  XOR U25296 ( .A(n25398), .B(n25399), .Z(n25389) );
  AND U25297 ( .A(n25400), .B(n25401), .Z(n25399) );
  XOR U25298 ( .A(n25398), .B(n25237), .Z(n25401) );
  XNOR U25299 ( .A(p_input[619]), .B(n25402), .Z(n25237) );
  AND U25300 ( .A(n899), .B(n25403), .Z(n25402) );
  XOR U25301 ( .A(p_input[635]), .B(p_input[619]), .Z(n25403) );
  XNOR U25302 ( .A(n25234), .B(n25398), .Z(n25400) );
  XOR U25303 ( .A(n25404), .B(n25405), .Z(n25234) );
  AND U25304 ( .A(n897), .B(n25406), .Z(n25405) );
  XOR U25305 ( .A(p_input[603]), .B(p_input[587]), .Z(n25406) );
  XOR U25306 ( .A(n25407), .B(n25408), .Z(n25398) );
  AND U25307 ( .A(n25409), .B(n25410), .Z(n25408) );
  XOR U25308 ( .A(n25407), .B(n25249), .Z(n25410) );
  XNOR U25309 ( .A(p_input[618]), .B(n25411), .Z(n25249) );
  AND U25310 ( .A(n899), .B(n25412), .Z(n25411) );
  XOR U25311 ( .A(p_input[634]), .B(p_input[618]), .Z(n25412) );
  XNOR U25312 ( .A(n25246), .B(n25407), .Z(n25409) );
  XOR U25313 ( .A(n25413), .B(n25414), .Z(n25246) );
  AND U25314 ( .A(n897), .B(n25415), .Z(n25414) );
  XOR U25315 ( .A(p_input[602]), .B(p_input[586]), .Z(n25415) );
  XOR U25316 ( .A(n25416), .B(n25417), .Z(n25407) );
  AND U25317 ( .A(n25418), .B(n25419), .Z(n25417) );
  XOR U25318 ( .A(n25416), .B(n25261), .Z(n25419) );
  XNOR U25319 ( .A(p_input[617]), .B(n25420), .Z(n25261) );
  AND U25320 ( .A(n899), .B(n25421), .Z(n25420) );
  XOR U25321 ( .A(p_input[633]), .B(p_input[617]), .Z(n25421) );
  XNOR U25322 ( .A(n25258), .B(n25416), .Z(n25418) );
  XOR U25323 ( .A(n25422), .B(n25423), .Z(n25258) );
  AND U25324 ( .A(n897), .B(n25424), .Z(n25423) );
  XOR U25325 ( .A(p_input[601]), .B(p_input[585]), .Z(n25424) );
  XOR U25326 ( .A(n25425), .B(n25426), .Z(n25416) );
  AND U25327 ( .A(n25427), .B(n25428), .Z(n25426) );
  XOR U25328 ( .A(n25425), .B(n25273), .Z(n25428) );
  XNOR U25329 ( .A(p_input[616]), .B(n25429), .Z(n25273) );
  AND U25330 ( .A(n899), .B(n25430), .Z(n25429) );
  XOR U25331 ( .A(p_input[632]), .B(p_input[616]), .Z(n25430) );
  XNOR U25332 ( .A(n25270), .B(n25425), .Z(n25427) );
  XOR U25333 ( .A(n25431), .B(n25432), .Z(n25270) );
  AND U25334 ( .A(n897), .B(n25433), .Z(n25432) );
  XOR U25335 ( .A(p_input[600]), .B(p_input[584]), .Z(n25433) );
  XOR U25336 ( .A(n25434), .B(n25435), .Z(n25425) );
  AND U25337 ( .A(n25436), .B(n25437), .Z(n25435) );
  XOR U25338 ( .A(n25434), .B(n25285), .Z(n25437) );
  XNOR U25339 ( .A(p_input[615]), .B(n25438), .Z(n25285) );
  AND U25340 ( .A(n899), .B(n25439), .Z(n25438) );
  XOR U25341 ( .A(p_input[631]), .B(p_input[615]), .Z(n25439) );
  XNOR U25342 ( .A(n25282), .B(n25434), .Z(n25436) );
  XOR U25343 ( .A(n25440), .B(n25441), .Z(n25282) );
  AND U25344 ( .A(n897), .B(n25442), .Z(n25441) );
  XOR U25345 ( .A(p_input[599]), .B(p_input[583]), .Z(n25442) );
  XOR U25346 ( .A(n25443), .B(n25444), .Z(n25434) );
  AND U25347 ( .A(n25445), .B(n25446), .Z(n25444) );
  XOR U25348 ( .A(n25443), .B(n25297), .Z(n25446) );
  XNOR U25349 ( .A(p_input[614]), .B(n25447), .Z(n25297) );
  AND U25350 ( .A(n899), .B(n25448), .Z(n25447) );
  XOR U25351 ( .A(p_input[630]), .B(p_input[614]), .Z(n25448) );
  XNOR U25352 ( .A(n25294), .B(n25443), .Z(n25445) );
  XOR U25353 ( .A(n25449), .B(n25450), .Z(n25294) );
  AND U25354 ( .A(n897), .B(n25451), .Z(n25450) );
  XOR U25355 ( .A(p_input[598]), .B(p_input[582]), .Z(n25451) );
  XOR U25356 ( .A(n25452), .B(n25453), .Z(n25443) );
  AND U25357 ( .A(n25454), .B(n25455), .Z(n25453) );
  XOR U25358 ( .A(n25452), .B(n25309), .Z(n25455) );
  XNOR U25359 ( .A(p_input[613]), .B(n25456), .Z(n25309) );
  AND U25360 ( .A(n899), .B(n25457), .Z(n25456) );
  XOR U25361 ( .A(p_input[629]), .B(p_input[613]), .Z(n25457) );
  XNOR U25362 ( .A(n25306), .B(n25452), .Z(n25454) );
  XOR U25363 ( .A(n25458), .B(n25459), .Z(n25306) );
  AND U25364 ( .A(n897), .B(n25460), .Z(n25459) );
  XOR U25365 ( .A(p_input[597]), .B(p_input[581]), .Z(n25460) );
  XOR U25366 ( .A(n25461), .B(n25462), .Z(n25452) );
  AND U25367 ( .A(n25463), .B(n25464), .Z(n25462) );
  XOR U25368 ( .A(n25461), .B(n25321), .Z(n25464) );
  XNOR U25369 ( .A(p_input[612]), .B(n25465), .Z(n25321) );
  AND U25370 ( .A(n899), .B(n25466), .Z(n25465) );
  XOR U25371 ( .A(p_input[628]), .B(p_input[612]), .Z(n25466) );
  XNOR U25372 ( .A(n25318), .B(n25461), .Z(n25463) );
  XOR U25373 ( .A(n25467), .B(n25468), .Z(n25318) );
  AND U25374 ( .A(n897), .B(n25469), .Z(n25468) );
  XOR U25375 ( .A(p_input[596]), .B(p_input[580]), .Z(n25469) );
  XOR U25376 ( .A(n25470), .B(n25471), .Z(n25461) );
  AND U25377 ( .A(n25472), .B(n25473), .Z(n25471) );
  XOR U25378 ( .A(n25470), .B(n25333), .Z(n25473) );
  XNOR U25379 ( .A(p_input[611]), .B(n25474), .Z(n25333) );
  AND U25380 ( .A(n899), .B(n25475), .Z(n25474) );
  XOR U25381 ( .A(p_input[627]), .B(p_input[611]), .Z(n25475) );
  XNOR U25382 ( .A(n25330), .B(n25470), .Z(n25472) );
  XOR U25383 ( .A(n25476), .B(n25477), .Z(n25330) );
  AND U25384 ( .A(n897), .B(n25478), .Z(n25477) );
  XOR U25385 ( .A(p_input[595]), .B(p_input[579]), .Z(n25478) );
  XOR U25386 ( .A(n25479), .B(n25480), .Z(n25470) );
  AND U25387 ( .A(n25481), .B(n25482), .Z(n25480) );
  XOR U25388 ( .A(n25479), .B(n25345), .Z(n25482) );
  XNOR U25389 ( .A(p_input[610]), .B(n25483), .Z(n25345) );
  AND U25390 ( .A(n899), .B(n25484), .Z(n25483) );
  XOR U25391 ( .A(p_input[626]), .B(p_input[610]), .Z(n25484) );
  XNOR U25392 ( .A(n25342), .B(n25479), .Z(n25481) );
  XOR U25393 ( .A(n25485), .B(n25486), .Z(n25342) );
  AND U25394 ( .A(n897), .B(n25487), .Z(n25486) );
  XOR U25395 ( .A(p_input[594]), .B(p_input[578]), .Z(n25487) );
  XOR U25396 ( .A(n25488), .B(n25489), .Z(n25479) );
  AND U25397 ( .A(n25490), .B(n25491), .Z(n25489) );
  XNOR U25398 ( .A(n25492), .B(n25358), .Z(n25491) );
  XNOR U25399 ( .A(p_input[609]), .B(n25493), .Z(n25358) );
  AND U25400 ( .A(n899), .B(n25494), .Z(n25493) );
  XNOR U25401 ( .A(p_input[625]), .B(n25495), .Z(n25494) );
  IV U25402 ( .A(p_input[609]), .Z(n25495) );
  XNOR U25403 ( .A(n25355), .B(n25488), .Z(n25490) );
  XNOR U25404 ( .A(p_input[577]), .B(n25496), .Z(n25355) );
  AND U25405 ( .A(n897), .B(n25497), .Z(n25496) );
  XOR U25406 ( .A(p_input[593]), .B(p_input[577]), .Z(n25497) );
  IV U25407 ( .A(n25492), .Z(n25488) );
  AND U25408 ( .A(n25363), .B(n25366), .Z(n25492) );
  XOR U25409 ( .A(p_input[608]), .B(n25498), .Z(n25366) );
  AND U25410 ( .A(n899), .B(n25499), .Z(n25498) );
  XOR U25411 ( .A(p_input[624]), .B(p_input[608]), .Z(n25499) );
  XOR U25412 ( .A(n25500), .B(n25501), .Z(n899) );
  AND U25413 ( .A(n25502), .B(n25503), .Z(n25501) );
  XNOR U25414 ( .A(p_input[639]), .B(n25500), .Z(n25503) );
  XOR U25415 ( .A(n25500), .B(p_input[623]), .Z(n25502) );
  XOR U25416 ( .A(n25504), .B(n25505), .Z(n25500) );
  AND U25417 ( .A(n25506), .B(n25507), .Z(n25505) );
  XNOR U25418 ( .A(p_input[638]), .B(n25504), .Z(n25507) );
  XOR U25419 ( .A(n25504), .B(p_input[622]), .Z(n25506) );
  XOR U25420 ( .A(n25508), .B(n25509), .Z(n25504) );
  AND U25421 ( .A(n25510), .B(n25511), .Z(n25509) );
  XNOR U25422 ( .A(p_input[637]), .B(n25508), .Z(n25511) );
  XOR U25423 ( .A(n25508), .B(p_input[621]), .Z(n25510) );
  XOR U25424 ( .A(n25512), .B(n25513), .Z(n25508) );
  AND U25425 ( .A(n25514), .B(n25515), .Z(n25513) );
  XNOR U25426 ( .A(p_input[636]), .B(n25512), .Z(n25515) );
  XOR U25427 ( .A(n25512), .B(p_input[620]), .Z(n25514) );
  XOR U25428 ( .A(n25516), .B(n25517), .Z(n25512) );
  AND U25429 ( .A(n25518), .B(n25519), .Z(n25517) );
  XNOR U25430 ( .A(p_input[635]), .B(n25516), .Z(n25519) );
  XOR U25431 ( .A(n25516), .B(p_input[619]), .Z(n25518) );
  XOR U25432 ( .A(n25520), .B(n25521), .Z(n25516) );
  AND U25433 ( .A(n25522), .B(n25523), .Z(n25521) );
  XNOR U25434 ( .A(p_input[634]), .B(n25520), .Z(n25523) );
  XOR U25435 ( .A(n25520), .B(p_input[618]), .Z(n25522) );
  XOR U25436 ( .A(n25524), .B(n25525), .Z(n25520) );
  AND U25437 ( .A(n25526), .B(n25527), .Z(n25525) );
  XNOR U25438 ( .A(p_input[633]), .B(n25524), .Z(n25527) );
  XOR U25439 ( .A(n25524), .B(p_input[617]), .Z(n25526) );
  XOR U25440 ( .A(n25528), .B(n25529), .Z(n25524) );
  AND U25441 ( .A(n25530), .B(n25531), .Z(n25529) );
  XNOR U25442 ( .A(p_input[632]), .B(n25528), .Z(n25531) );
  XOR U25443 ( .A(n25528), .B(p_input[616]), .Z(n25530) );
  XOR U25444 ( .A(n25532), .B(n25533), .Z(n25528) );
  AND U25445 ( .A(n25534), .B(n25535), .Z(n25533) );
  XNOR U25446 ( .A(p_input[631]), .B(n25532), .Z(n25535) );
  XOR U25447 ( .A(n25532), .B(p_input[615]), .Z(n25534) );
  XOR U25448 ( .A(n25536), .B(n25537), .Z(n25532) );
  AND U25449 ( .A(n25538), .B(n25539), .Z(n25537) );
  XNOR U25450 ( .A(p_input[630]), .B(n25536), .Z(n25539) );
  XOR U25451 ( .A(n25536), .B(p_input[614]), .Z(n25538) );
  XOR U25452 ( .A(n25540), .B(n25541), .Z(n25536) );
  AND U25453 ( .A(n25542), .B(n25543), .Z(n25541) );
  XNOR U25454 ( .A(p_input[629]), .B(n25540), .Z(n25543) );
  XOR U25455 ( .A(n25540), .B(p_input[613]), .Z(n25542) );
  XOR U25456 ( .A(n25544), .B(n25545), .Z(n25540) );
  AND U25457 ( .A(n25546), .B(n25547), .Z(n25545) );
  XNOR U25458 ( .A(p_input[628]), .B(n25544), .Z(n25547) );
  XOR U25459 ( .A(n25544), .B(p_input[612]), .Z(n25546) );
  XOR U25460 ( .A(n25548), .B(n25549), .Z(n25544) );
  AND U25461 ( .A(n25550), .B(n25551), .Z(n25549) );
  XNOR U25462 ( .A(p_input[627]), .B(n25548), .Z(n25551) );
  XOR U25463 ( .A(n25548), .B(p_input[611]), .Z(n25550) );
  XOR U25464 ( .A(n25552), .B(n25553), .Z(n25548) );
  AND U25465 ( .A(n25554), .B(n25555), .Z(n25553) );
  XNOR U25466 ( .A(p_input[626]), .B(n25552), .Z(n25555) );
  XOR U25467 ( .A(n25552), .B(p_input[610]), .Z(n25554) );
  XNOR U25468 ( .A(n25556), .B(n25557), .Z(n25552) );
  AND U25469 ( .A(n25558), .B(n25559), .Z(n25557) );
  XOR U25470 ( .A(p_input[625]), .B(n25556), .Z(n25559) );
  XNOR U25471 ( .A(p_input[609]), .B(n25556), .Z(n25558) );
  AND U25472 ( .A(p_input[624]), .B(n25560), .Z(n25556) );
  IV U25473 ( .A(p_input[608]), .Z(n25560) );
  XNOR U25474 ( .A(p_input[576]), .B(n25561), .Z(n25363) );
  AND U25475 ( .A(n897), .B(n25562), .Z(n25561) );
  XOR U25476 ( .A(p_input[592]), .B(p_input[576]), .Z(n25562) );
  XOR U25477 ( .A(n25563), .B(n25564), .Z(n897) );
  AND U25478 ( .A(n25565), .B(n25566), .Z(n25564) );
  XNOR U25479 ( .A(p_input[607]), .B(n25563), .Z(n25566) );
  XOR U25480 ( .A(n25563), .B(p_input[591]), .Z(n25565) );
  XOR U25481 ( .A(n25567), .B(n25568), .Z(n25563) );
  AND U25482 ( .A(n25569), .B(n25570), .Z(n25568) );
  XNOR U25483 ( .A(p_input[606]), .B(n25567), .Z(n25570) );
  XNOR U25484 ( .A(n25567), .B(n25377), .Z(n25569) );
  IV U25485 ( .A(p_input[590]), .Z(n25377) );
  XOR U25486 ( .A(n25571), .B(n25572), .Z(n25567) );
  AND U25487 ( .A(n25573), .B(n25574), .Z(n25572) );
  XNOR U25488 ( .A(p_input[605]), .B(n25571), .Z(n25574) );
  XNOR U25489 ( .A(n25571), .B(n25386), .Z(n25573) );
  IV U25490 ( .A(p_input[589]), .Z(n25386) );
  XOR U25491 ( .A(n25575), .B(n25576), .Z(n25571) );
  AND U25492 ( .A(n25577), .B(n25578), .Z(n25576) );
  XNOR U25493 ( .A(p_input[604]), .B(n25575), .Z(n25578) );
  XNOR U25494 ( .A(n25575), .B(n25395), .Z(n25577) );
  IV U25495 ( .A(p_input[588]), .Z(n25395) );
  XOR U25496 ( .A(n25579), .B(n25580), .Z(n25575) );
  AND U25497 ( .A(n25581), .B(n25582), .Z(n25580) );
  XNOR U25498 ( .A(p_input[603]), .B(n25579), .Z(n25582) );
  XNOR U25499 ( .A(n25579), .B(n25404), .Z(n25581) );
  IV U25500 ( .A(p_input[587]), .Z(n25404) );
  XOR U25501 ( .A(n25583), .B(n25584), .Z(n25579) );
  AND U25502 ( .A(n25585), .B(n25586), .Z(n25584) );
  XNOR U25503 ( .A(p_input[602]), .B(n25583), .Z(n25586) );
  XNOR U25504 ( .A(n25583), .B(n25413), .Z(n25585) );
  IV U25505 ( .A(p_input[586]), .Z(n25413) );
  XOR U25506 ( .A(n25587), .B(n25588), .Z(n25583) );
  AND U25507 ( .A(n25589), .B(n25590), .Z(n25588) );
  XNOR U25508 ( .A(p_input[601]), .B(n25587), .Z(n25590) );
  XNOR U25509 ( .A(n25587), .B(n25422), .Z(n25589) );
  IV U25510 ( .A(p_input[585]), .Z(n25422) );
  XOR U25511 ( .A(n25591), .B(n25592), .Z(n25587) );
  AND U25512 ( .A(n25593), .B(n25594), .Z(n25592) );
  XNOR U25513 ( .A(p_input[600]), .B(n25591), .Z(n25594) );
  XNOR U25514 ( .A(n25591), .B(n25431), .Z(n25593) );
  IV U25515 ( .A(p_input[584]), .Z(n25431) );
  XOR U25516 ( .A(n25595), .B(n25596), .Z(n25591) );
  AND U25517 ( .A(n25597), .B(n25598), .Z(n25596) );
  XNOR U25518 ( .A(p_input[599]), .B(n25595), .Z(n25598) );
  XNOR U25519 ( .A(n25595), .B(n25440), .Z(n25597) );
  IV U25520 ( .A(p_input[583]), .Z(n25440) );
  XOR U25521 ( .A(n25599), .B(n25600), .Z(n25595) );
  AND U25522 ( .A(n25601), .B(n25602), .Z(n25600) );
  XNOR U25523 ( .A(p_input[598]), .B(n25599), .Z(n25602) );
  XNOR U25524 ( .A(n25599), .B(n25449), .Z(n25601) );
  IV U25525 ( .A(p_input[582]), .Z(n25449) );
  XOR U25526 ( .A(n25603), .B(n25604), .Z(n25599) );
  AND U25527 ( .A(n25605), .B(n25606), .Z(n25604) );
  XNOR U25528 ( .A(p_input[597]), .B(n25603), .Z(n25606) );
  XNOR U25529 ( .A(n25603), .B(n25458), .Z(n25605) );
  IV U25530 ( .A(p_input[581]), .Z(n25458) );
  XOR U25531 ( .A(n25607), .B(n25608), .Z(n25603) );
  AND U25532 ( .A(n25609), .B(n25610), .Z(n25608) );
  XNOR U25533 ( .A(p_input[596]), .B(n25607), .Z(n25610) );
  XNOR U25534 ( .A(n25607), .B(n25467), .Z(n25609) );
  IV U25535 ( .A(p_input[580]), .Z(n25467) );
  XOR U25536 ( .A(n25611), .B(n25612), .Z(n25607) );
  AND U25537 ( .A(n25613), .B(n25614), .Z(n25612) );
  XNOR U25538 ( .A(p_input[595]), .B(n25611), .Z(n25614) );
  XNOR U25539 ( .A(n25611), .B(n25476), .Z(n25613) );
  IV U25540 ( .A(p_input[579]), .Z(n25476) );
  XOR U25541 ( .A(n25615), .B(n25616), .Z(n25611) );
  AND U25542 ( .A(n25617), .B(n25618), .Z(n25616) );
  XNOR U25543 ( .A(p_input[594]), .B(n25615), .Z(n25618) );
  XNOR U25544 ( .A(n25615), .B(n25485), .Z(n25617) );
  IV U25545 ( .A(p_input[578]), .Z(n25485) );
  XNOR U25546 ( .A(n25619), .B(n25620), .Z(n25615) );
  AND U25547 ( .A(n25621), .B(n25622), .Z(n25620) );
  XOR U25548 ( .A(p_input[593]), .B(n25619), .Z(n25622) );
  XNOR U25549 ( .A(p_input[577]), .B(n25619), .Z(n25621) );
  AND U25550 ( .A(p_input[592]), .B(n25623), .Z(n25619) );
  IV U25551 ( .A(p_input[576]), .Z(n25623) );
  XOR U25552 ( .A(n25624), .B(n25625), .Z(n25182) );
  AND U25553 ( .A(n556), .B(n25626), .Z(n25625) );
  XNOR U25554 ( .A(n25627), .B(n25624), .Z(n25626) );
  XOR U25555 ( .A(n25628), .B(n25629), .Z(n556) );
  AND U25556 ( .A(n25630), .B(n25631), .Z(n25629) );
  XNOR U25557 ( .A(n25193), .B(n25628), .Z(n25631) );
  AND U25558 ( .A(p_input[575]), .B(p_input[559]), .Z(n25193) );
  XOR U25559 ( .A(n25628), .B(n25192), .Z(n25630) );
  AND U25560 ( .A(p_input[527]), .B(p_input[543]), .Z(n25192) );
  XOR U25561 ( .A(n25632), .B(n25633), .Z(n25628) );
  AND U25562 ( .A(n25634), .B(n25635), .Z(n25633) );
  XOR U25563 ( .A(n25632), .B(n25205), .Z(n25635) );
  XNOR U25564 ( .A(p_input[558]), .B(n25636), .Z(n25205) );
  AND U25565 ( .A(n903), .B(n25637), .Z(n25636) );
  XOR U25566 ( .A(p_input[574]), .B(p_input[558]), .Z(n25637) );
  XNOR U25567 ( .A(n25202), .B(n25632), .Z(n25634) );
  XOR U25568 ( .A(n25638), .B(n25639), .Z(n25202) );
  AND U25569 ( .A(n900), .B(n25640), .Z(n25639) );
  XOR U25570 ( .A(p_input[542]), .B(p_input[526]), .Z(n25640) );
  XOR U25571 ( .A(n25641), .B(n25642), .Z(n25632) );
  AND U25572 ( .A(n25643), .B(n25644), .Z(n25642) );
  XOR U25573 ( .A(n25641), .B(n25217), .Z(n25644) );
  XNOR U25574 ( .A(p_input[557]), .B(n25645), .Z(n25217) );
  AND U25575 ( .A(n903), .B(n25646), .Z(n25645) );
  XOR U25576 ( .A(p_input[573]), .B(p_input[557]), .Z(n25646) );
  XNOR U25577 ( .A(n25214), .B(n25641), .Z(n25643) );
  XOR U25578 ( .A(n25647), .B(n25648), .Z(n25214) );
  AND U25579 ( .A(n900), .B(n25649), .Z(n25648) );
  XOR U25580 ( .A(p_input[541]), .B(p_input[525]), .Z(n25649) );
  XOR U25581 ( .A(n25650), .B(n25651), .Z(n25641) );
  AND U25582 ( .A(n25652), .B(n25653), .Z(n25651) );
  XOR U25583 ( .A(n25650), .B(n25229), .Z(n25653) );
  XNOR U25584 ( .A(p_input[556]), .B(n25654), .Z(n25229) );
  AND U25585 ( .A(n903), .B(n25655), .Z(n25654) );
  XOR U25586 ( .A(p_input[572]), .B(p_input[556]), .Z(n25655) );
  XNOR U25587 ( .A(n25226), .B(n25650), .Z(n25652) );
  XOR U25588 ( .A(n25656), .B(n25657), .Z(n25226) );
  AND U25589 ( .A(n900), .B(n25658), .Z(n25657) );
  XOR U25590 ( .A(p_input[540]), .B(p_input[524]), .Z(n25658) );
  XOR U25591 ( .A(n25659), .B(n25660), .Z(n25650) );
  AND U25592 ( .A(n25661), .B(n25662), .Z(n25660) );
  XOR U25593 ( .A(n25659), .B(n25241), .Z(n25662) );
  XNOR U25594 ( .A(p_input[555]), .B(n25663), .Z(n25241) );
  AND U25595 ( .A(n903), .B(n25664), .Z(n25663) );
  XOR U25596 ( .A(p_input[571]), .B(p_input[555]), .Z(n25664) );
  XNOR U25597 ( .A(n25238), .B(n25659), .Z(n25661) );
  XOR U25598 ( .A(n25665), .B(n25666), .Z(n25238) );
  AND U25599 ( .A(n900), .B(n25667), .Z(n25666) );
  XOR U25600 ( .A(p_input[539]), .B(p_input[523]), .Z(n25667) );
  XOR U25601 ( .A(n25668), .B(n25669), .Z(n25659) );
  AND U25602 ( .A(n25670), .B(n25671), .Z(n25669) );
  XOR U25603 ( .A(n25668), .B(n25253), .Z(n25671) );
  XNOR U25604 ( .A(p_input[554]), .B(n25672), .Z(n25253) );
  AND U25605 ( .A(n903), .B(n25673), .Z(n25672) );
  XOR U25606 ( .A(p_input[570]), .B(p_input[554]), .Z(n25673) );
  XNOR U25607 ( .A(n25250), .B(n25668), .Z(n25670) );
  XOR U25608 ( .A(n25674), .B(n25675), .Z(n25250) );
  AND U25609 ( .A(n900), .B(n25676), .Z(n25675) );
  XOR U25610 ( .A(p_input[538]), .B(p_input[522]), .Z(n25676) );
  XOR U25611 ( .A(n25677), .B(n25678), .Z(n25668) );
  AND U25612 ( .A(n25679), .B(n25680), .Z(n25678) );
  XOR U25613 ( .A(n25677), .B(n25265), .Z(n25680) );
  XNOR U25614 ( .A(p_input[553]), .B(n25681), .Z(n25265) );
  AND U25615 ( .A(n903), .B(n25682), .Z(n25681) );
  XOR U25616 ( .A(p_input[569]), .B(p_input[553]), .Z(n25682) );
  XNOR U25617 ( .A(n25262), .B(n25677), .Z(n25679) );
  XOR U25618 ( .A(n25683), .B(n25684), .Z(n25262) );
  AND U25619 ( .A(n900), .B(n25685), .Z(n25684) );
  XOR U25620 ( .A(p_input[537]), .B(p_input[521]), .Z(n25685) );
  XOR U25621 ( .A(n25686), .B(n25687), .Z(n25677) );
  AND U25622 ( .A(n25688), .B(n25689), .Z(n25687) );
  XOR U25623 ( .A(n25686), .B(n25277), .Z(n25689) );
  XNOR U25624 ( .A(p_input[552]), .B(n25690), .Z(n25277) );
  AND U25625 ( .A(n903), .B(n25691), .Z(n25690) );
  XOR U25626 ( .A(p_input[568]), .B(p_input[552]), .Z(n25691) );
  XNOR U25627 ( .A(n25274), .B(n25686), .Z(n25688) );
  XOR U25628 ( .A(n25692), .B(n25693), .Z(n25274) );
  AND U25629 ( .A(n900), .B(n25694), .Z(n25693) );
  XOR U25630 ( .A(p_input[536]), .B(p_input[520]), .Z(n25694) );
  XOR U25631 ( .A(n25695), .B(n25696), .Z(n25686) );
  AND U25632 ( .A(n25697), .B(n25698), .Z(n25696) );
  XOR U25633 ( .A(n25695), .B(n25289), .Z(n25698) );
  XNOR U25634 ( .A(p_input[551]), .B(n25699), .Z(n25289) );
  AND U25635 ( .A(n903), .B(n25700), .Z(n25699) );
  XOR U25636 ( .A(p_input[567]), .B(p_input[551]), .Z(n25700) );
  XNOR U25637 ( .A(n25286), .B(n25695), .Z(n25697) );
  XOR U25638 ( .A(n25701), .B(n25702), .Z(n25286) );
  AND U25639 ( .A(n900), .B(n25703), .Z(n25702) );
  XOR U25640 ( .A(p_input[535]), .B(p_input[519]), .Z(n25703) );
  XOR U25641 ( .A(n25704), .B(n25705), .Z(n25695) );
  AND U25642 ( .A(n25706), .B(n25707), .Z(n25705) );
  XOR U25643 ( .A(n25704), .B(n25301), .Z(n25707) );
  XNOR U25644 ( .A(p_input[550]), .B(n25708), .Z(n25301) );
  AND U25645 ( .A(n903), .B(n25709), .Z(n25708) );
  XOR U25646 ( .A(p_input[566]), .B(p_input[550]), .Z(n25709) );
  XNOR U25647 ( .A(n25298), .B(n25704), .Z(n25706) );
  XOR U25648 ( .A(n25710), .B(n25711), .Z(n25298) );
  AND U25649 ( .A(n900), .B(n25712), .Z(n25711) );
  XOR U25650 ( .A(p_input[534]), .B(p_input[518]), .Z(n25712) );
  XOR U25651 ( .A(n25713), .B(n25714), .Z(n25704) );
  AND U25652 ( .A(n25715), .B(n25716), .Z(n25714) );
  XOR U25653 ( .A(n25713), .B(n25313), .Z(n25716) );
  XNOR U25654 ( .A(p_input[549]), .B(n25717), .Z(n25313) );
  AND U25655 ( .A(n903), .B(n25718), .Z(n25717) );
  XOR U25656 ( .A(p_input[565]), .B(p_input[549]), .Z(n25718) );
  XNOR U25657 ( .A(n25310), .B(n25713), .Z(n25715) );
  XOR U25658 ( .A(n25719), .B(n25720), .Z(n25310) );
  AND U25659 ( .A(n900), .B(n25721), .Z(n25720) );
  XOR U25660 ( .A(p_input[533]), .B(p_input[517]), .Z(n25721) );
  XOR U25661 ( .A(n25722), .B(n25723), .Z(n25713) );
  AND U25662 ( .A(n25724), .B(n25725), .Z(n25723) );
  XOR U25663 ( .A(n25722), .B(n25325), .Z(n25725) );
  XNOR U25664 ( .A(p_input[548]), .B(n25726), .Z(n25325) );
  AND U25665 ( .A(n903), .B(n25727), .Z(n25726) );
  XOR U25666 ( .A(p_input[564]), .B(p_input[548]), .Z(n25727) );
  XNOR U25667 ( .A(n25322), .B(n25722), .Z(n25724) );
  XOR U25668 ( .A(n25728), .B(n25729), .Z(n25322) );
  AND U25669 ( .A(n900), .B(n25730), .Z(n25729) );
  XOR U25670 ( .A(p_input[532]), .B(p_input[516]), .Z(n25730) );
  XOR U25671 ( .A(n25731), .B(n25732), .Z(n25722) );
  AND U25672 ( .A(n25733), .B(n25734), .Z(n25732) );
  XOR U25673 ( .A(n25731), .B(n25337), .Z(n25734) );
  XNOR U25674 ( .A(p_input[547]), .B(n25735), .Z(n25337) );
  AND U25675 ( .A(n903), .B(n25736), .Z(n25735) );
  XOR U25676 ( .A(p_input[563]), .B(p_input[547]), .Z(n25736) );
  XNOR U25677 ( .A(n25334), .B(n25731), .Z(n25733) );
  XOR U25678 ( .A(n25737), .B(n25738), .Z(n25334) );
  AND U25679 ( .A(n900), .B(n25739), .Z(n25738) );
  XOR U25680 ( .A(p_input[531]), .B(p_input[515]), .Z(n25739) );
  XOR U25681 ( .A(n25740), .B(n25741), .Z(n25731) );
  AND U25682 ( .A(n25742), .B(n25743), .Z(n25741) );
  XOR U25683 ( .A(n25740), .B(n25349), .Z(n25743) );
  XNOR U25684 ( .A(p_input[546]), .B(n25744), .Z(n25349) );
  AND U25685 ( .A(n903), .B(n25745), .Z(n25744) );
  XOR U25686 ( .A(p_input[562]), .B(p_input[546]), .Z(n25745) );
  XNOR U25687 ( .A(n25346), .B(n25740), .Z(n25742) );
  XOR U25688 ( .A(n25746), .B(n25747), .Z(n25346) );
  AND U25689 ( .A(n900), .B(n25748), .Z(n25747) );
  XOR U25690 ( .A(p_input[530]), .B(p_input[514]), .Z(n25748) );
  XOR U25691 ( .A(n25749), .B(n25750), .Z(n25740) );
  AND U25692 ( .A(n25751), .B(n25752), .Z(n25750) );
  XNOR U25693 ( .A(n25753), .B(n25362), .Z(n25752) );
  XNOR U25694 ( .A(p_input[545]), .B(n25754), .Z(n25362) );
  AND U25695 ( .A(n903), .B(n25755), .Z(n25754) );
  XNOR U25696 ( .A(p_input[561]), .B(n25756), .Z(n25755) );
  IV U25697 ( .A(p_input[545]), .Z(n25756) );
  XNOR U25698 ( .A(n25359), .B(n25749), .Z(n25751) );
  XNOR U25699 ( .A(p_input[513]), .B(n25757), .Z(n25359) );
  AND U25700 ( .A(n900), .B(n25758), .Z(n25757) );
  XOR U25701 ( .A(p_input[529]), .B(p_input[513]), .Z(n25758) );
  IV U25702 ( .A(n25753), .Z(n25749) );
  AND U25703 ( .A(n25624), .B(n25627), .Z(n25753) );
  XOR U25704 ( .A(p_input[544]), .B(n25759), .Z(n25627) );
  AND U25705 ( .A(n903), .B(n25760), .Z(n25759) );
  XOR U25706 ( .A(p_input[560]), .B(p_input[544]), .Z(n25760) );
  XOR U25707 ( .A(n25761), .B(n25762), .Z(n903) );
  AND U25708 ( .A(n25763), .B(n25764), .Z(n25762) );
  XNOR U25709 ( .A(p_input[575]), .B(n25761), .Z(n25764) );
  XOR U25710 ( .A(n25761), .B(p_input[559]), .Z(n25763) );
  XOR U25711 ( .A(n25765), .B(n25766), .Z(n25761) );
  AND U25712 ( .A(n25767), .B(n25768), .Z(n25766) );
  XNOR U25713 ( .A(p_input[574]), .B(n25765), .Z(n25768) );
  XOR U25714 ( .A(n25765), .B(p_input[558]), .Z(n25767) );
  XOR U25715 ( .A(n25769), .B(n25770), .Z(n25765) );
  AND U25716 ( .A(n25771), .B(n25772), .Z(n25770) );
  XNOR U25717 ( .A(p_input[573]), .B(n25769), .Z(n25772) );
  XOR U25718 ( .A(n25769), .B(p_input[557]), .Z(n25771) );
  XOR U25719 ( .A(n25773), .B(n25774), .Z(n25769) );
  AND U25720 ( .A(n25775), .B(n25776), .Z(n25774) );
  XNOR U25721 ( .A(p_input[572]), .B(n25773), .Z(n25776) );
  XOR U25722 ( .A(n25773), .B(p_input[556]), .Z(n25775) );
  XOR U25723 ( .A(n25777), .B(n25778), .Z(n25773) );
  AND U25724 ( .A(n25779), .B(n25780), .Z(n25778) );
  XNOR U25725 ( .A(p_input[571]), .B(n25777), .Z(n25780) );
  XOR U25726 ( .A(n25777), .B(p_input[555]), .Z(n25779) );
  XOR U25727 ( .A(n25781), .B(n25782), .Z(n25777) );
  AND U25728 ( .A(n25783), .B(n25784), .Z(n25782) );
  XNOR U25729 ( .A(p_input[570]), .B(n25781), .Z(n25784) );
  XOR U25730 ( .A(n25781), .B(p_input[554]), .Z(n25783) );
  XOR U25731 ( .A(n25785), .B(n25786), .Z(n25781) );
  AND U25732 ( .A(n25787), .B(n25788), .Z(n25786) );
  XNOR U25733 ( .A(p_input[569]), .B(n25785), .Z(n25788) );
  XOR U25734 ( .A(n25785), .B(p_input[553]), .Z(n25787) );
  XOR U25735 ( .A(n25789), .B(n25790), .Z(n25785) );
  AND U25736 ( .A(n25791), .B(n25792), .Z(n25790) );
  XNOR U25737 ( .A(p_input[568]), .B(n25789), .Z(n25792) );
  XOR U25738 ( .A(n25789), .B(p_input[552]), .Z(n25791) );
  XOR U25739 ( .A(n25793), .B(n25794), .Z(n25789) );
  AND U25740 ( .A(n25795), .B(n25796), .Z(n25794) );
  XNOR U25741 ( .A(p_input[567]), .B(n25793), .Z(n25796) );
  XOR U25742 ( .A(n25793), .B(p_input[551]), .Z(n25795) );
  XOR U25743 ( .A(n25797), .B(n25798), .Z(n25793) );
  AND U25744 ( .A(n25799), .B(n25800), .Z(n25798) );
  XNOR U25745 ( .A(p_input[566]), .B(n25797), .Z(n25800) );
  XOR U25746 ( .A(n25797), .B(p_input[550]), .Z(n25799) );
  XOR U25747 ( .A(n25801), .B(n25802), .Z(n25797) );
  AND U25748 ( .A(n25803), .B(n25804), .Z(n25802) );
  XNOR U25749 ( .A(p_input[565]), .B(n25801), .Z(n25804) );
  XOR U25750 ( .A(n25801), .B(p_input[549]), .Z(n25803) );
  XOR U25751 ( .A(n25805), .B(n25806), .Z(n25801) );
  AND U25752 ( .A(n25807), .B(n25808), .Z(n25806) );
  XNOR U25753 ( .A(p_input[564]), .B(n25805), .Z(n25808) );
  XOR U25754 ( .A(n25805), .B(p_input[548]), .Z(n25807) );
  XOR U25755 ( .A(n25809), .B(n25810), .Z(n25805) );
  AND U25756 ( .A(n25811), .B(n25812), .Z(n25810) );
  XNOR U25757 ( .A(p_input[563]), .B(n25809), .Z(n25812) );
  XOR U25758 ( .A(n25809), .B(p_input[547]), .Z(n25811) );
  XOR U25759 ( .A(n25813), .B(n25814), .Z(n25809) );
  AND U25760 ( .A(n25815), .B(n25816), .Z(n25814) );
  XNOR U25761 ( .A(p_input[562]), .B(n25813), .Z(n25816) );
  XOR U25762 ( .A(n25813), .B(p_input[546]), .Z(n25815) );
  XNOR U25763 ( .A(n25817), .B(n25818), .Z(n25813) );
  AND U25764 ( .A(n25819), .B(n25820), .Z(n25818) );
  XOR U25765 ( .A(p_input[561]), .B(n25817), .Z(n25820) );
  XNOR U25766 ( .A(p_input[545]), .B(n25817), .Z(n25819) );
  AND U25767 ( .A(p_input[560]), .B(n25821), .Z(n25817) );
  IV U25768 ( .A(p_input[544]), .Z(n25821) );
  XNOR U25769 ( .A(p_input[512]), .B(n25822), .Z(n25624) );
  AND U25770 ( .A(n900), .B(n25823), .Z(n25822) );
  XOR U25771 ( .A(p_input[528]), .B(p_input[512]), .Z(n25823) );
  XOR U25772 ( .A(n25824), .B(n25825), .Z(n900) );
  AND U25773 ( .A(n25826), .B(n25827), .Z(n25825) );
  XNOR U25774 ( .A(p_input[543]), .B(n25824), .Z(n25827) );
  XOR U25775 ( .A(n25824), .B(p_input[527]), .Z(n25826) );
  XOR U25776 ( .A(n25828), .B(n25829), .Z(n25824) );
  AND U25777 ( .A(n25830), .B(n25831), .Z(n25829) );
  XNOR U25778 ( .A(p_input[542]), .B(n25828), .Z(n25831) );
  XNOR U25779 ( .A(n25828), .B(n25638), .Z(n25830) );
  IV U25780 ( .A(p_input[526]), .Z(n25638) );
  XOR U25781 ( .A(n25832), .B(n25833), .Z(n25828) );
  AND U25782 ( .A(n25834), .B(n25835), .Z(n25833) );
  XNOR U25783 ( .A(p_input[541]), .B(n25832), .Z(n25835) );
  XNOR U25784 ( .A(n25832), .B(n25647), .Z(n25834) );
  IV U25785 ( .A(p_input[525]), .Z(n25647) );
  XOR U25786 ( .A(n25836), .B(n25837), .Z(n25832) );
  AND U25787 ( .A(n25838), .B(n25839), .Z(n25837) );
  XNOR U25788 ( .A(p_input[540]), .B(n25836), .Z(n25839) );
  XNOR U25789 ( .A(n25836), .B(n25656), .Z(n25838) );
  IV U25790 ( .A(p_input[524]), .Z(n25656) );
  XOR U25791 ( .A(n25840), .B(n25841), .Z(n25836) );
  AND U25792 ( .A(n25842), .B(n25843), .Z(n25841) );
  XNOR U25793 ( .A(p_input[539]), .B(n25840), .Z(n25843) );
  XNOR U25794 ( .A(n25840), .B(n25665), .Z(n25842) );
  IV U25795 ( .A(p_input[523]), .Z(n25665) );
  XOR U25796 ( .A(n25844), .B(n25845), .Z(n25840) );
  AND U25797 ( .A(n25846), .B(n25847), .Z(n25845) );
  XNOR U25798 ( .A(p_input[538]), .B(n25844), .Z(n25847) );
  XNOR U25799 ( .A(n25844), .B(n25674), .Z(n25846) );
  IV U25800 ( .A(p_input[522]), .Z(n25674) );
  XOR U25801 ( .A(n25848), .B(n25849), .Z(n25844) );
  AND U25802 ( .A(n25850), .B(n25851), .Z(n25849) );
  XNOR U25803 ( .A(p_input[537]), .B(n25848), .Z(n25851) );
  XNOR U25804 ( .A(n25848), .B(n25683), .Z(n25850) );
  IV U25805 ( .A(p_input[521]), .Z(n25683) );
  XOR U25806 ( .A(n25852), .B(n25853), .Z(n25848) );
  AND U25807 ( .A(n25854), .B(n25855), .Z(n25853) );
  XNOR U25808 ( .A(p_input[536]), .B(n25852), .Z(n25855) );
  XNOR U25809 ( .A(n25852), .B(n25692), .Z(n25854) );
  IV U25810 ( .A(p_input[520]), .Z(n25692) );
  XOR U25811 ( .A(n25856), .B(n25857), .Z(n25852) );
  AND U25812 ( .A(n25858), .B(n25859), .Z(n25857) );
  XNOR U25813 ( .A(p_input[535]), .B(n25856), .Z(n25859) );
  XNOR U25814 ( .A(n25856), .B(n25701), .Z(n25858) );
  IV U25815 ( .A(p_input[519]), .Z(n25701) );
  XOR U25816 ( .A(n25860), .B(n25861), .Z(n25856) );
  AND U25817 ( .A(n25862), .B(n25863), .Z(n25861) );
  XNOR U25818 ( .A(p_input[534]), .B(n25860), .Z(n25863) );
  XNOR U25819 ( .A(n25860), .B(n25710), .Z(n25862) );
  IV U25820 ( .A(p_input[518]), .Z(n25710) );
  XOR U25821 ( .A(n25864), .B(n25865), .Z(n25860) );
  AND U25822 ( .A(n25866), .B(n25867), .Z(n25865) );
  XNOR U25823 ( .A(p_input[533]), .B(n25864), .Z(n25867) );
  XNOR U25824 ( .A(n25864), .B(n25719), .Z(n25866) );
  IV U25825 ( .A(p_input[517]), .Z(n25719) );
  XOR U25826 ( .A(n25868), .B(n25869), .Z(n25864) );
  AND U25827 ( .A(n25870), .B(n25871), .Z(n25869) );
  XNOR U25828 ( .A(p_input[532]), .B(n25868), .Z(n25871) );
  XNOR U25829 ( .A(n25868), .B(n25728), .Z(n25870) );
  IV U25830 ( .A(p_input[516]), .Z(n25728) );
  XOR U25831 ( .A(n25872), .B(n25873), .Z(n25868) );
  AND U25832 ( .A(n25874), .B(n25875), .Z(n25873) );
  XNOR U25833 ( .A(p_input[531]), .B(n25872), .Z(n25875) );
  XNOR U25834 ( .A(n25872), .B(n25737), .Z(n25874) );
  IV U25835 ( .A(p_input[515]), .Z(n25737) );
  XOR U25836 ( .A(n25876), .B(n25877), .Z(n25872) );
  AND U25837 ( .A(n25878), .B(n25879), .Z(n25877) );
  XNOR U25838 ( .A(p_input[530]), .B(n25876), .Z(n25879) );
  XNOR U25839 ( .A(n25876), .B(n25746), .Z(n25878) );
  IV U25840 ( .A(p_input[514]), .Z(n25746) );
  XNOR U25841 ( .A(n25880), .B(n25881), .Z(n25876) );
  AND U25842 ( .A(n25882), .B(n25883), .Z(n25881) );
  XOR U25843 ( .A(p_input[529]), .B(n25880), .Z(n25883) );
  XNOR U25844 ( .A(p_input[513]), .B(n25880), .Z(n25882) );
  AND U25845 ( .A(p_input[528]), .B(n25884), .Z(n25880) );
  IV U25846 ( .A(p_input[512]), .Z(n25884) );
  XOR U25847 ( .A(n25885), .B(n25886), .Z(n22339) );
  AND U25848 ( .A(n1020), .B(n25887), .Z(n25886) );
  XNOR U25849 ( .A(n25888), .B(n25885), .Z(n25887) );
  XOR U25850 ( .A(n25889), .B(n25890), .Z(n1020) );
  AND U25851 ( .A(n25891), .B(n25892), .Z(n25890) );
  XOR U25852 ( .A(n25889), .B(n22354), .Z(n25892) );
  XNOR U25853 ( .A(n25893), .B(n25894), .Z(n22354) );
  AND U25854 ( .A(n25895), .B(n963), .Z(n25894) );
  AND U25855 ( .A(n25893), .B(n25896), .Z(n25895) );
  XNOR U25856 ( .A(n22351), .B(n25889), .Z(n25891) );
  XOR U25857 ( .A(n25897), .B(n25898), .Z(n22351) );
  AND U25858 ( .A(n25899), .B(n960), .Z(n25898) );
  NOR U25859 ( .A(n25897), .B(n25900), .Z(n25899) );
  XOR U25860 ( .A(n25901), .B(n25902), .Z(n25889) );
  AND U25861 ( .A(n25903), .B(n25904), .Z(n25902) );
  XOR U25862 ( .A(n25901), .B(n22366), .Z(n25904) );
  XOR U25863 ( .A(n25905), .B(n25906), .Z(n22366) );
  AND U25864 ( .A(n963), .B(n25907), .Z(n25906) );
  XOR U25865 ( .A(n25908), .B(n25905), .Z(n25907) );
  XNOR U25866 ( .A(n22363), .B(n25901), .Z(n25903) );
  XOR U25867 ( .A(n25909), .B(n25910), .Z(n22363) );
  AND U25868 ( .A(n960), .B(n25911), .Z(n25910) );
  XOR U25869 ( .A(n25912), .B(n25909), .Z(n25911) );
  XOR U25870 ( .A(n25913), .B(n25914), .Z(n25901) );
  AND U25871 ( .A(n25915), .B(n25916), .Z(n25914) );
  XOR U25872 ( .A(n25913), .B(n22378), .Z(n25916) );
  XOR U25873 ( .A(n25917), .B(n25918), .Z(n22378) );
  AND U25874 ( .A(n963), .B(n25919), .Z(n25918) );
  XOR U25875 ( .A(n25920), .B(n25917), .Z(n25919) );
  XNOR U25876 ( .A(n22375), .B(n25913), .Z(n25915) );
  XOR U25877 ( .A(n25921), .B(n25922), .Z(n22375) );
  AND U25878 ( .A(n960), .B(n25923), .Z(n25922) );
  XOR U25879 ( .A(n25924), .B(n25921), .Z(n25923) );
  XOR U25880 ( .A(n25925), .B(n25926), .Z(n25913) );
  AND U25881 ( .A(n25927), .B(n25928), .Z(n25926) );
  XOR U25882 ( .A(n25925), .B(n22390), .Z(n25928) );
  XOR U25883 ( .A(n25929), .B(n25930), .Z(n22390) );
  AND U25884 ( .A(n963), .B(n25931), .Z(n25930) );
  XOR U25885 ( .A(n25932), .B(n25929), .Z(n25931) );
  XNOR U25886 ( .A(n22387), .B(n25925), .Z(n25927) );
  XOR U25887 ( .A(n25933), .B(n25934), .Z(n22387) );
  AND U25888 ( .A(n960), .B(n25935), .Z(n25934) );
  XOR U25889 ( .A(n25936), .B(n25933), .Z(n25935) );
  XOR U25890 ( .A(n25937), .B(n25938), .Z(n25925) );
  AND U25891 ( .A(n25939), .B(n25940), .Z(n25938) );
  XOR U25892 ( .A(n25937), .B(n22402), .Z(n25940) );
  XOR U25893 ( .A(n25941), .B(n25942), .Z(n22402) );
  AND U25894 ( .A(n963), .B(n25943), .Z(n25942) );
  XOR U25895 ( .A(n25944), .B(n25941), .Z(n25943) );
  XNOR U25896 ( .A(n22399), .B(n25937), .Z(n25939) );
  XOR U25897 ( .A(n25945), .B(n25946), .Z(n22399) );
  AND U25898 ( .A(n960), .B(n25947), .Z(n25946) );
  XOR U25899 ( .A(n25948), .B(n25945), .Z(n25947) );
  XOR U25900 ( .A(n25949), .B(n25950), .Z(n25937) );
  AND U25901 ( .A(n25951), .B(n25952), .Z(n25950) );
  XOR U25902 ( .A(n25949), .B(n22414), .Z(n25952) );
  XOR U25903 ( .A(n25953), .B(n25954), .Z(n22414) );
  AND U25904 ( .A(n963), .B(n25955), .Z(n25954) );
  XOR U25905 ( .A(n25956), .B(n25953), .Z(n25955) );
  XNOR U25906 ( .A(n22411), .B(n25949), .Z(n25951) );
  XOR U25907 ( .A(n25957), .B(n25958), .Z(n22411) );
  AND U25908 ( .A(n960), .B(n25959), .Z(n25958) );
  XOR U25909 ( .A(n25960), .B(n25957), .Z(n25959) );
  XOR U25910 ( .A(n25961), .B(n25962), .Z(n25949) );
  AND U25911 ( .A(n25963), .B(n25964), .Z(n25962) );
  XOR U25912 ( .A(n25961), .B(n22426), .Z(n25964) );
  XOR U25913 ( .A(n25965), .B(n25966), .Z(n22426) );
  AND U25914 ( .A(n963), .B(n25967), .Z(n25966) );
  XOR U25915 ( .A(n25968), .B(n25965), .Z(n25967) );
  XNOR U25916 ( .A(n22423), .B(n25961), .Z(n25963) );
  XOR U25917 ( .A(n25969), .B(n25970), .Z(n22423) );
  AND U25918 ( .A(n960), .B(n25971), .Z(n25970) );
  XOR U25919 ( .A(n25972), .B(n25969), .Z(n25971) );
  XOR U25920 ( .A(n25973), .B(n25974), .Z(n25961) );
  AND U25921 ( .A(n25975), .B(n25976), .Z(n25974) );
  XOR U25922 ( .A(n25973), .B(n22438), .Z(n25976) );
  XOR U25923 ( .A(n25977), .B(n25978), .Z(n22438) );
  AND U25924 ( .A(n963), .B(n25979), .Z(n25978) );
  XOR U25925 ( .A(n25980), .B(n25977), .Z(n25979) );
  XNOR U25926 ( .A(n22435), .B(n25973), .Z(n25975) );
  XOR U25927 ( .A(n25981), .B(n25982), .Z(n22435) );
  AND U25928 ( .A(n960), .B(n25983), .Z(n25982) );
  XOR U25929 ( .A(n25984), .B(n25981), .Z(n25983) );
  XOR U25930 ( .A(n25985), .B(n25986), .Z(n25973) );
  AND U25931 ( .A(n25987), .B(n25988), .Z(n25986) );
  XOR U25932 ( .A(n25985), .B(n22450), .Z(n25988) );
  XOR U25933 ( .A(n25989), .B(n25990), .Z(n22450) );
  AND U25934 ( .A(n963), .B(n25991), .Z(n25990) );
  XOR U25935 ( .A(n25992), .B(n25989), .Z(n25991) );
  XNOR U25936 ( .A(n22447), .B(n25985), .Z(n25987) );
  XOR U25937 ( .A(n25993), .B(n25994), .Z(n22447) );
  AND U25938 ( .A(n960), .B(n25995), .Z(n25994) );
  XOR U25939 ( .A(n25996), .B(n25993), .Z(n25995) );
  XOR U25940 ( .A(n25997), .B(n25998), .Z(n25985) );
  AND U25941 ( .A(n25999), .B(n26000), .Z(n25998) );
  XOR U25942 ( .A(n25997), .B(n22462), .Z(n26000) );
  XOR U25943 ( .A(n26001), .B(n26002), .Z(n22462) );
  AND U25944 ( .A(n963), .B(n26003), .Z(n26002) );
  XOR U25945 ( .A(n26004), .B(n26001), .Z(n26003) );
  XNOR U25946 ( .A(n22459), .B(n25997), .Z(n25999) );
  XOR U25947 ( .A(n26005), .B(n26006), .Z(n22459) );
  AND U25948 ( .A(n960), .B(n26007), .Z(n26006) );
  XOR U25949 ( .A(n26008), .B(n26005), .Z(n26007) );
  XOR U25950 ( .A(n26009), .B(n26010), .Z(n25997) );
  AND U25951 ( .A(n26011), .B(n26012), .Z(n26010) );
  XOR U25952 ( .A(n26009), .B(n22474), .Z(n26012) );
  XOR U25953 ( .A(n26013), .B(n26014), .Z(n22474) );
  AND U25954 ( .A(n963), .B(n26015), .Z(n26014) );
  XOR U25955 ( .A(n26016), .B(n26013), .Z(n26015) );
  XNOR U25956 ( .A(n22471), .B(n26009), .Z(n26011) );
  XOR U25957 ( .A(n26017), .B(n26018), .Z(n22471) );
  AND U25958 ( .A(n960), .B(n26019), .Z(n26018) );
  XOR U25959 ( .A(n26020), .B(n26017), .Z(n26019) );
  XOR U25960 ( .A(n26021), .B(n26022), .Z(n26009) );
  AND U25961 ( .A(n26023), .B(n26024), .Z(n26022) );
  XOR U25962 ( .A(n26021), .B(n22486), .Z(n26024) );
  XOR U25963 ( .A(n26025), .B(n26026), .Z(n22486) );
  AND U25964 ( .A(n963), .B(n26027), .Z(n26026) );
  XOR U25965 ( .A(n26028), .B(n26025), .Z(n26027) );
  XNOR U25966 ( .A(n22483), .B(n26021), .Z(n26023) );
  XOR U25967 ( .A(n26029), .B(n26030), .Z(n22483) );
  AND U25968 ( .A(n960), .B(n26031), .Z(n26030) );
  XOR U25969 ( .A(n26032), .B(n26029), .Z(n26031) );
  XOR U25970 ( .A(n26033), .B(n26034), .Z(n26021) );
  AND U25971 ( .A(n26035), .B(n26036), .Z(n26034) );
  XOR U25972 ( .A(n26033), .B(n22498), .Z(n26036) );
  XOR U25973 ( .A(n26037), .B(n26038), .Z(n22498) );
  AND U25974 ( .A(n963), .B(n26039), .Z(n26038) );
  XOR U25975 ( .A(n26040), .B(n26037), .Z(n26039) );
  XNOR U25976 ( .A(n22495), .B(n26033), .Z(n26035) );
  XOR U25977 ( .A(n26041), .B(n26042), .Z(n22495) );
  AND U25978 ( .A(n960), .B(n26043), .Z(n26042) );
  XOR U25979 ( .A(n26044), .B(n26041), .Z(n26043) );
  XOR U25980 ( .A(n26045), .B(n26046), .Z(n26033) );
  AND U25981 ( .A(n26047), .B(n26048), .Z(n26046) );
  XOR U25982 ( .A(n26045), .B(n22510), .Z(n26048) );
  XOR U25983 ( .A(n26049), .B(n26050), .Z(n22510) );
  AND U25984 ( .A(n963), .B(n26051), .Z(n26050) );
  XOR U25985 ( .A(n26052), .B(n26049), .Z(n26051) );
  XNOR U25986 ( .A(n22507), .B(n26045), .Z(n26047) );
  XOR U25987 ( .A(n26053), .B(n26054), .Z(n22507) );
  AND U25988 ( .A(n960), .B(n26055), .Z(n26054) );
  XOR U25989 ( .A(n26056), .B(n26053), .Z(n26055) );
  XOR U25990 ( .A(n26057), .B(n26058), .Z(n26045) );
  AND U25991 ( .A(n26059), .B(n26060), .Z(n26058) );
  XNOR U25992 ( .A(n26061), .B(n22523), .Z(n26060) );
  XOR U25993 ( .A(n26062), .B(n26063), .Z(n22523) );
  AND U25994 ( .A(n963), .B(n26064), .Z(n26063) );
  XOR U25995 ( .A(n26062), .B(n26065), .Z(n26064) );
  XNOR U25996 ( .A(n22520), .B(n26057), .Z(n26059) );
  XOR U25997 ( .A(n26066), .B(n26067), .Z(n22520) );
  AND U25998 ( .A(n960), .B(n26068), .Z(n26067) );
  XOR U25999 ( .A(n26066), .B(n26069), .Z(n26068) );
  IV U26000 ( .A(n26061), .Z(n26057) );
  AND U26001 ( .A(n25885), .B(n25888), .Z(n26061) );
  XNOR U26002 ( .A(n26070), .B(n26071), .Z(n25888) );
  AND U26003 ( .A(n963), .B(n26072), .Z(n26071) );
  XNOR U26004 ( .A(n26073), .B(n26070), .Z(n26072) );
  XOR U26005 ( .A(n26074), .B(n26075), .Z(n963) );
  AND U26006 ( .A(n26076), .B(n26077), .Z(n26075) );
  XOR U26007 ( .A(n25896), .B(n26074), .Z(n26077) );
  IV U26008 ( .A(n26078), .Z(n25896) );
  AND U26009 ( .A(n26079), .B(n26080), .Z(n26078) );
  XOR U26010 ( .A(n26074), .B(n25893), .Z(n26076) );
  AND U26011 ( .A(n26081), .B(n26082), .Z(n25893) );
  XOR U26012 ( .A(n26083), .B(n26084), .Z(n26074) );
  AND U26013 ( .A(n26085), .B(n26086), .Z(n26084) );
  XOR U26014 ( .A(n26083), .B(n25908), .Z(n26086) );
  XOR U26015 ( .A(n26087), .B(n26088), .Z(n25908) );
  AND U26016 ( .A(n835), .B(n26089), .Z(n26088) );
  XOR U26017 ( .A(n26090), .B(n26087), .Z(n26089) );
  XNOR U26018 ( .A(n25905), .B(n26083), .Z(n26085) );
  XOR U26019 ( .A(n26091), .B(n26092), .Z(n25905) );
  AND U26020 ( .A(n833), .B(n26093), .Z(n26092) );
  XOR U26021 ( .A(n26094), .B(n26091), .Z(n26093) );
  XOR U26022 ( .A(n26095), .B(n26096), .Z(n26083) );
  AND U26023 ( .A(n26097), .B(n26098), .Z(n26096) );
  XOR U26024 ( .A(n26095), .B(n25920), .Z(n26098) );
  XOR U26025 ( .A(n26099), .B(n26100), .Z(n25920) );
  AND U26026 ( .A(n835), .B(n26101), .Z(n26100) );
  XOR U26027 ( .A(n26102), .B(n26099), .Z(n26101) );
  XNOR U26028 ( .A(n25917), .B(n26095), .Z(n26097) );
  XOR U26029 ( .A(n26103), .B(n26104), .Z(n25917) );
  AND U26030 ( .A(n833), .B(n26105), .Z(n26104) );
  XOR U26031 ( .A(n26106), .B(n26103), .Z(n26105) );
  XOR U26032 ( .A(n26107), .B(n26108), .Z(n26095) );
  AND U26033 ( .A(n26109), .B(n26110), .Z(n26108) );
  XOR U26034 ( .A(n26107), .B(n25932), .Z(n26110) );
  XOR U26035 ( .A(n26111), .B(n26112), .Z(n25932) );
  AND U26036 ( .A(n835), .B(n26113), .Z(n26112) );
  XOR U26037 ( .A(n26114), .B(n26111), .Z(n26113) );
  XNOR U26038 ( .A(n25929), .B(n26107), .Z(n26109) );
  XOR U26039 ( .A(n26115), .B(n26116), .Z(n25929) );
  AND U26040 ( .A(n833), .B(n26117), .Z(n26116) );
  XOR U26041 ( .A(n26118), .B(n26115), .Z(n26117) );
  XOR U26042 ( .A(n26119), .B(n26120), .Z(n26107) );
  AND U26043 ( .A(n26121), .B(n26122), .Z(n26120) );
  XOR U26044 ( .A(n26119), .B(n25944), .Z(n26122) );
  XOR U26045 ( .A(n26123), .B(n26124), .Z(n25944) );
  AND U26046 ( .A(n835), .B(n26125), .Z(n26124) );
  XOR U26047 ( .A(n26126), .B(n26123), .Z(n26125) );
  XNOR U26048 ( .A(n25941), .B(n26119), .Z(n26121) );
  XOR U26049 ( .A(n26127), .B(n26128), .Z(n25941) );
  AND U26050 ( .A(n833), .B(n26129), .Z(n26128) );
  XOR U26051 ( .A(n26130), .B(n26127), .Z(n26129) );
  XOR U26052 ( .A(n26131), .B(n26132), .Z(n26119) );
  AND U26053 ( .A(n26133), .B(n26134), .Z(n26132) );
  XOR U26054 ( .A(n26131), .B(n25956), .Z(n26134) );
  XOR U26055 ( .A(n26135), .B(n26136), .Z(n25956) );
  AND U26056 ( .A(n835), .B(n26137), .Z(n26136) );
  XOR U26057 ( .A(n26138), .B(n26135), .Z(n26137) );
  XNOR U26058 ( .A(n25953), .B(n26131), .Z(n26133) );
  XOR U26059 ( .A(n26139), .B(n26140), .Z(n25953) );
  AND U26060 ( .A(n833), .B(n26141), .Z(n26140) );
  XOR U26061 ( .A(n26142), .B(n26139), .Z(n26141) );
  XOR U26062 ( .A(n26143), .B(n26144), .Z(n26131) );
  AND U26063 ( .A(n26145), .B(n26146), .Z(n26144) );
  XOR U26064 ( .A(n26143), .B(n25968), .Z(n26146) );
  XOR U26065 ( .A(n26147), .B(n26148), .Z(n25968) );
  AND U26066 ( .A(n835), .B(n26149), .Z(n26148) );
  XOR U26067 ( .A(n26150), .B(n26147), .Z(n26149) );
  XNOR U26068 ( .A(n25965), .B(n26143), .Z(n26145) );
  XOR U26069 ( .A(n26151), .B(n26152), .Z(n25965) );
  AND U26070 ( .A(n833), .B(n26153), .Z(n26152) );
  XOR U26071 ( .A(n26154), .B(n26151), .Z(n26153) );
  XOR U26072 ( .A(n26155), .B(n26156), .Z(n26143) );
  AND U26073 ( .A(n26157), .B(n26158), .Z(n26156) );
  XOR U26074 ( .A(n26155), .B(n25980), .Z(n26158) );
  XOR U26075 ( .A(n26159), .B(n26160), .Z(n25980) );
  AND U26076 ( .A(n835), .B(n26161), .Z(n26160) );
  XOR U26077 ( .A(n26162), .B(n26159), .Z(n26161) );
  XNOR U26078 ( .A(n25977), .B(n26155), .Z(n26157) );
  XOR U26079 ( .A(n26163), .B(n26164), .Z(n25977) );
  AND U26080 ( .A(n833), .B(n26165), .Z(n26164) );
  XOR U26081 ( .A(n26166), .B(n26163), .Z(n26165) );
  XOR U26082 ( .A(n26167), .B(n26168), .Z(n26155) );
  AND U26083 ( .A(n26169), .B(n26170), .Z(n26168) );
  XOR U26084 ( .A(n26167), .B(n25992), .Z(n26170) );
  XOR U26085 ( .A(n26171), .B(n26172), .Z(n25992) );
  AND U26086 ( .A(n835), .B(n26173), .Z(n26172) );
  XOR U26087 ( .A(n26174), .B(n26171), .Z(n26173) );
  XNOR U26088 ( .A(n25989), .B(n26167), .Z(n26169) );
  XOR U26089 ( .A(n26175), .B(n26176), .Z(n25989) );
  AND U26090 ( .A(n833), .B(n26177), .Z(n26176) );
  XOR U26091 ( .A(n26178), .B(n26175), .Z(n26177) );
  XOR U26092 ( .A(n26179), .B(n26180), .Z(n26167) );
  AND U26093 ( .A(n26181), .B(n26182), .Z(n26180) );
  XOR U26094 ( .A(n26179), .B(n26004), .Z(n26182) );
  XOR U26095 ( .A(n26183), .B(n26184), .Z(n26004) );
  AND U26096 ( .A(n835), .B(n26185), .Z(n26184) );
  XOR U26097 ( .A(n26186), .B(n26183), .Z(n26185) );
  XNOR U26098 ( .A(n26001), .B(n26179), .Z(n26181) );
  XOR U26099 ( .A(n26187), .B(n26188), .Z(n26001) );
  AND U26100 ( .A(n833), .B(n26189), .Z(n26188) );
  XOR U26101 ( .A(n26190), .B(n26187), .Z(n26189) );
  XOR U26102 ( .A(n26191), .B(n26192), .Z(n26179) );
  AND U26103 ( .A(n26193), .B(n26194), .Z(n26192) );
  XOR U26104 ( .A(n26191), .B(n26016), .Z(n26194) );
  XOR U26105 ( .A(n26195), .B(n26196), .Z(n26016) );
  AND U26106 ( .A(n835), .B(n26197), .Z(n26196) );
  XOR U26107 ( .A(n26198), .B(n26195), .Z(n26197) );
  XNOR U26108 ( .A(n26013), .B(n26191), .Z(n26193) );
  XOR U26109 ( .A(n26199), .B(n26200), .Z(n26013) );
  AND U26110 ( .A(n833), .B(n26201), .Z(n26200) );
  XOR U26111 ( .A(n26202), .B(n26199), .Z(n26201) );
  XOR U26112 ( .A(n26203), .B(n26204), .Z(n26191) );
  AND U26113 ( .A(n26205), .B(n26206), .Z(n26204) );
  XOR U26114 ( .A(n26203), .B(n26028), .Z(n26206) );
  XOR U26115 ( .A(n26207), .B(n26208), .Z(n26028) );
  AND U26116 ( .A(n835), .B(n26209), .Z(n26208) );
  XOR U26117 ( .A(n26210), .B(n26207), .Z(n26209) );
  XNOR U26118 ( .A(n26025), .B(n26203), .Z(n26205) );
  XOR U26119 ( .A(n26211), .B(n26212), .Z(n26025) );
  AND U26120 ( .A(n833), .B(n26213), .Z(n26212) );
  XOR U26121 ( .A(n26214), .B(n26211), .Z(n26213) );
  XOR U26122 ( .A(n26215), .B(n26216), .Z(n26203) );
  AND U26123 ( .A(n26217), .B(n26218), .Z(n26216) );
  XOR U26124 ( .A(n26215), .B(n26040), .Z(n26218) );
  XOR U26125 ( .A(n26219), .B(n26220), .Z(n26040) );
  AND U26126 ( .A(n835), .B(n26221), .Z(n26220) );
  XOR U26127 ( .A(n26222), .B(n26219), .Z(n26221) );
  XNOR U26128 ( .A(n26037), .B(n26215), .Z(n26217) );
  XOR U26129 ( .A(n26223), .B(n26224), .Z(n26037) );
  AND U26130 ( .A(n833), .B(n26225), .Z(n26224) );
  XOR U26131 ( .A(n26226), .B(n26223), .Z(n26225) );
  XOR U26132 ( .A(n26227), .B(n26228), .Z(n26215) );
  AND U26133 ( .A(n26229), .B(n26230), .Z(n26228) );
  XOR U26134 ( .A(n26227), .B(n26052), .Z(n26230) );
  XOR U26135 ( .A(n26231), .B(n26232), .Z(n26052) );
  AND U26136 ( .A(n835), .B(n26233), .Z(n26232) );
  XOR U26137 ( .A(n26234), .B(n26231), .Z(n26233) );
  XNOR U26138 ( .A(n26049), .B(n26227), .Z(n26229) );
  XOR U26139 ( .A(n26235), .B(n26236), .Z(n26049) );
  AND U26140 ( .A(n833), .B(n26237), .Z(n26236) );
  XOR U26141 ( .A(n26238), .B(n26235), .Z(n26237) );
  XOR U26142 ( .A(n26239), .B(n26240), .Z(n26227) );
  AND U26143 ( .A(n26241), .B(n26242), .Z(n26240) );
  XNOR U26144 ( .A(n26243), .B(n26065), .Z(n26242) );
  XOR U26145 ( .A(n26244), .B(n26245), .Z(n26065) );
  AND U26146 ( .A(n835), .B(n26246), .Z(n26245) );
  XOR U26147 ( .A(n26244), .B(n26247), .Z(n26246) );
  XNOR U26148 ( .A(n26062), .B(n26239), .Z(n26241) );
  XOR U26149 ( .A(n26248), .B(n26249), .Z(n26062) );
  AND U26150 ( .A(n833), .B(n26250), .Z(n26249) );
  XOR U26151 ( .A(n26248), .B(n26251), .Z(n26250) );
  IV U26152 ( .A(n26243), .Z(n26239) );
  AND U26153 ( .A(n26070), .B(n26073), .Z(n26243) );
  XNOR U26154 ( .A(n26252), .B(n26253), .Z(n26073) );
  AND U26155 ( .A(n835), .B(n26254), .Z(n26253) );
  XNOR U26156 ( .A(n26255), .B(n26252), .Z(n26254) );
  XOR U26157 ( .A(n26256), .B(n26257), .Z(n835) );
  AND U26158 ( .A(n26258), .B(n26259), .Z(n26257) );
  XNOR U26159 ( .A(n26079), .B(n26256), .Z(n26259) );
  AND U26160 ( .A(n26260), .B(n26261), .Z(n26079) );
  XOR U26161 ( .A(n26256), .B(n26080), .Z(n26258) );
  AND U26162 ( .A(n26262), .B(n26263), .Z(n26080) );
  XOR U26163 ( .A(n26264), .B(n26265), .Z(n26256) );
  AND U26164 ( .A(n26266), .B(n26267), .Z(n26265) );
  XOR U26165 ( .A(n26264), .B(n26090), .Z(n26267) );
  XOR U26166 ( .A(n26268), .B(n26269), .Z(n26090) );
  AND U26167 ( .A(n571), .B(n26270), .Z(n26269) );
  XOR U26168 ( .A(n26271), .B(n26268), .Z(n26270) );
  XNOR U26169 ( .A(n26087), .B(n26264), .Z(n26266) );
  XOR U26170 ( .A(n26272), .B(n26273), .Z(n26087) );
  AND U26171 ( .A(n569), .B(n26274), .Z(n26273) );
  XOR U26172 ( .A(n26275), .B(n26272), .Z(n26274) );
  XOR U26173 ( .A(n26276), .B(n26277), .Z(n26264) );
  AND U26174 ( .A(n26278), .B(n26279), .Z(n26277) );
  XOR U26175 ( .A(n26276), .B(n26102), .Z(n26279) );
  XOR U26176 ( .A(n26280), .B(n26281), .Z(n26102) );
  AND U26177 ( .A(n571), .B(n26282), .Z(n26281) );
  XOR U26178 ( .A(n26283), .B(n26280), .Z(n26282) );
  XNOR U26179 ( .A(n26099), .B(n26276), .Z(n26278) );
  XOR U26180 ( .A(n26284), .B(n26285), .Z(n26099) );
  AND U26181 ( .A(n569), .B(n26286), .Z(n26285) );
  XOR U26182 ( .A(n26287), .B(n26284), .Z(n26286) );
  XOR U26183 ( .A(n26288), .B(n26289), .Z(n26276) );
  AND U26184 ( .A(n26290), .B(n26291), .Z(n26289) );
  XOR U26185 ( .A(n26288), .B(n26114), .Z(n26291) );
  XOR U26186 ( .A(n26292), .B(n26293), .Z(n26114) );
  AND U26187 ( .A(n571), .B(n26294), .Z(n26293) );
  XOR U26188 ( .A(n26295), .B(n26292), .Z(n26294) );
  XNOR U26189 ( .A(n26111), .B(n26288), .Z(n26290) );
  XOR U26190 ( .A(n26296), .B(n26297), .Z(n26111) );
  AND U26191 ( .A(n569), .B(n26298), .Z(n26297) );
  XOR U26192 ( .A(n26299), .B(n26296), .Z(n26298) );
  XOR U26193 ( .A(n26300), .B(n26301), .Z(n26288) );
  AND U26194 ( .A(n26302), .B(n26303), .Z(n26301) );
  XOR U26195 ( .A(n26300), .B(n26126), .Z(n26303) );
  XOR U26196 ( .A(n26304), .B(n26305), .Z(n26126) );
  AND U26197 ( .A(n571), .B(n26306), .Z(n26305) );
  XOR U26198 ( .A(n26307), .B(n26304), .Z(n26306) );
  XNOR U26199 ( .A(n26123), .B(n26300), .Z(n26302) );
  XOR U26200 ( .A(n26308), .B(n26309), .Z(n26123) );
  AND U26201 ( .A(n569), .B(n26310), .Z(n26309) );
  XOR U26202 ( .A(n26311), .B(n26308), .Z(n26310) );
  XOR U26203 ( .A(n26312), .B(n26313), .Z(n26300) );
  AND U26204 ( .A(n26314), .B(n26315), .Z(n26313) );
  XOR U26205 ( .A(n26312), .B(n26138), .Z(n26315) );
  XOR U26206 ( .A(n26316), .B(n26317), .Z(n26138) );
  AND U26207 ( .A(n571), .B(n26318), .Z(n26317) );
  XOR U26208 ( .A(n26319), .B(n26316), .Z(n26318) );
  XNOR U26209 ( .A(n26135), .B(n26312), .Z(n26314) );
  XOR U26210 ( .A(n26320), .B(n26321), .Z(n26135) );
  AND U26211 ( .A(n569), .B(n26322), .Z(n26321) );
  XOR U26212 ( .A(n26323), .B(n26320), .Z(n26322) );
  XOR U26213 ( .A(n26324), .B(n26325), .Z(n26312) );
  AND U26214 ( .A(n26326), .B(n26327), .Z(n26325) );
  XOR U26215 ( .A(n26324), .B(n26150), .Z(n26327) );
  XOR U26216 ( .A(n26328), .B(n26329), .Z(n26150) );
  AND U26217 ( .A(n571), .B(n26330), .Z(n26329) );
  XOR U26218 ( .A(n26331), .B(n26328), .Z(n26330) );
  XNOR U26219 ( .A(n26147), .B(n26324), .Z(n26326) );
  XOR U26220 ( .A(n26332), .B(n26333), .Z(n26147) );
  AND U26221 ( .A(n569), .B(n26334), .Z(n26333) );
  XOR U26222 ( .A(n26335), .B(n26332), .Z(n26334) );
  XOR U26223 ( .A(n26336), .B(n26337), .Z(n26324) );
  AND U26224 ( .A(n26338), .B(n26339), .Z(n26337) );
  XOR U26225 ( .A(n26336), .B(n26162), .Z(n26339) );
  XOR U26226 ( .A(n26340), .B(n26341), .Z(n26162) );
  AND U26227 ( .A(n571), .B(n26342), .Z(n26341) );
  XOR U26228 ( .A(n26343), .B(n26340), .Z(n26342) );
  XNOR U26229 ( .A(n26159), .B(n26336), .Z(n26338) );
  XOR U26230 ( .A(n26344), .B(n26345), .Z(n26159) );
  AND U26231 ( .A(n569), .B(n26346), .Z(n26345) );
  XOR U26232 ( .A(n26347), .B(n26344), .Z(n26346) );
  XOR U26233 ( .A(n26348), .B(n26349), .Z(n26336) );
  AND U26234 ( .A(n26350), .B(n26351), .Z(n26349) );
  XOR U26235 ( .A(n26348), .B(n26174), .Z(n26351) );
  XOR U26236 ( .A(n26352), .B(n26353), .Z(n26174) );
  AND U26237 ( .A(n571), .B(n26354), .Z(n26353) );
  XOR U26238 ( .A(n26355), .B(n26352), .Z(n26354) );
  XNOR U26239 ( .A(n26171), .B(n26348), .Z(n26350) );
  XOR U26240 ( .A(n26356), .B(n26357), .Z(n26171) );
  AND U26241 ( .A(n569), .B(n26358), .Z(n26357) );
  XOR U26242 ( .A(n26359), .B(n26356), .Z(n26358) );
  XOR U26243 ( .A(n26360), .B(n26361), .Z(n26348) );
  AND U26244 ( .A(n26362), .B(n26363), .Z(n26361) );
  XOR U26245 ( .A(n26360), .B(n26186), .Z(n26363) );
  XOR U26246 ( .A(n26364), .B(n26365), .Z(n26186) );
  AND U26247 ( .A(n571), .B(n26366), .Z(n26365) );
  XOR U26248 ( .A(n26367), .B(n26364), .Z(n26366) );
  XNOR U26249 ( .A(n26183), .B(n26360), .Z(n26362) );
  XOR U26250 ( .A(n26368), .B(n26369), .Z(n26183) );
  AND U26251 ( .A(n569), .B(n26370), .Z(n26369) );
  XOR U26252 ( .A(n26371), .B(n26368), .Z(n26370) );
  XOR U26253 ( .A(n26372), .B(n26373), .Z(n26360) );
  AND U26254 ( .A(n26374), .B(n26375), .Z(n26373) );
  XOR U26255 ( .A(n26372), .B(n26198), .Z(n26375) );
  XOR U26256 ( .A(n26376), .B(n26377), .Z(n26198) );
  AND U26257 ( .A(n571), .B(n26378), .Z(n26377) );
  XOR U26258 ( .A(n26379), .B(n26376), .Z(n26378) );
  XNOR U26259 ( .A(n26195), .B(n26372), .Z(n26374) );
  XOR U26260 ( .A(n26380), .B(n26381), .Z(n26195) );
  AND U26261 ( .A(n569), .B(n26382), .Z(n26381) );
  XOR U26262 ( .A(n26383), .B(n26380), .Z(n26382) );
  XOR U26263 ( .A(n26384), .B(n26385), .Z(n26372) );
  AND U26264 ( .A(n26386), .B(n26387), .Z(n26385) );
  XOR U26265 ( .A(n26384), .B(n26210), .Z(n26387) );
  XOR U26266 ( .A(n26388), .B(n26389), .Z(n26210) );
  AND U26267 ( .A(n571), .B(n26390), .Z(n26389) );
  XOR U26268 ( .A(n26391), .B(n26388), .Z(n26390) );
  XNOR U26269 ( .A(n26207), .B(n26384), .Z(n26386) );
  XOR U26270 ( .A(n26392), .B(n26393), .Z(n26207) );
  AND U26271 ( .A(n569), .B(n26394), .Z(n26393) );
  XOR U26272 ( .A(n26395), .B(n26392), .Z(n26394) );
  XOR U26273 ( .A(n26396), .B(n26397), .Z(n26384) );
  AND U26274 ( .A(n26398), .B(n26399), .Z(n26397) );
  XOR U26275 ( .A(n26396), .B(n26222), .Z(n26399) );
  XOR U26276 ( .A(n26400), .B(n26401), .Z(n26222) );
  AND U26277 ( .A(n571), .B(n26402), .Z(n26401) );
  XOR U26278 ( .A(n26403), .B(n26400), .Z(n26402) );
  XNOR U26279 ( .A(n26219), .B(n26396), .Z(n26398) );
  XOR U26280 ( .A(n26404), .B(n26405), .Z(n26219) );
  AND U26281 ( .A(n569), .B(n26406), .Z(n26405) );
  XOR U26282 ( .A(n26407), .B(n26404), .Z(n26406) );
  XOR U26283 ( .A(n26408), .B(n26409), .Z(n26396) );
  AND U26284 ( .A(n26410), .B(n26411), .Z(n26409) );
  XOR U26285 ( .A(n26408), .B(n26234), .Z(n26411) );
  XOR U26286 ( .A(n26412), .B(n26413), .Z(n26234) );
  AND U26287 ( .A(n571), .B(n26414), .Z(n26413) );
  XOR U26288 ( .A(n26415), .B(n26412), .Z(n26414) );
  XNOR U26289 ( .A(n26231), .B(n26408), .Z(n26410) );
  XOR U26290 ( .A(n26416), .B(n26417), .Z(n26231) );
  AND U26291 ( .A(n569), .B(n26418), .Z(n26417) );
  XOR U26292 ( .A(n26419), .B(n26416), .Z(n26418) );
  XOR U26293 ( .A(n26420), .B(n26421), .Z(n26408) );
  AND U26294 ( .A(n26422), .B(n26423), .Z(n26421) );
  XNOR U26295 ( .A(n26424), .B(n26247), .Z(n26423) );
  XOR U26296 ( .A(n26425), .B(n26426), .Z(n26247) );
  AND U26297 ( .A(n571), .B(n26427), .Z(n26426) );
  XOR U26298 ( .A(n26425), .B(n26428), .Z(n26427) );
  XNOR U26299 ( .A(n26244), .B(n26420), .Z(n26422) );
  XOR U26300 ( .A(n26429), .B(n26430), .Z(n26244) );
  AND U26301 ( .A(n569), .B(n26431), .Z(n26430) );
  XOR U26302 ( .A(n26429), .B(n26432), .Z(n26431) );
  IV U26303 ( .A(n26424), .Z(n26420) );
  AND U26304 ( .A(n26252), .B(n26255), .Z(n26424) );
  XNOR U26305 ( .A(n26433), .B(n26434), .Z(n26255) );
  AND U26306 ( .A(n571), .B(n26435), .Z(n26434) );
  XNOR U26307 ( .A(n26436), .B(n26433), .Z(n26435) );
  XOR U26308 ( .A(n26437), .B(n26438), .Z(n571) );
  AND U26309 ( .A(n26439), .B(n26440), .Z(n26438) );
  XNOR U26310 ( .A(n26260), .B(n26437), .Z(n26440) );
  AND U26311 ( .A(p_input[511]), .B(p_input[495]), .Z(n26260) );
  XOR U26312 ( .A(n26437), .B(n26261), .Z(n26439) );
  AND U26313 ( .A(p_input[479]), .B(p_input[463]), .Z(n26261) );
  XOR U26314 ( .A(n26441), .B(n26442), .Z(n26437) );
  AND U26315 ( .A(n26443), .B(n26444), .Z(n26442) );
  XOR U26316 ( .A(n26441), .B(n26271), .Z(n26444) );
  XNOR U26317 ( .A(p_input[494]), .B(n26445), .Z(n26271) );
  AND U26318 ( .A(n979), .B(n26446), .Z(n26445) );
  XOR U26319 ( .A(p_input[510]), .B(p_input[494]), .Z(n26446) );
  XNOR U26320 ( .A(n26268), .B(n26441), .Z(n26443) );
  XOR U26321 ( .A(n26447), .B(n26448), .Z(n26268) );
  AND U26322 ( .A(n977), .B(n26449), .Z(n26448) );
  XOR U26323 ( .A(p_input[478]), .B(p_input[462]), .Z(n26449) );
  XOR U26324 ( .A(n26450), .B(n26451), .Z(n26441) );
  AND U26325 ( .A(n26452), .B(n26453), .Z(n26451) );
  XOR U26326 ( .A(n26450), .B(n26283), .Z(n26453) );
  XNOR U26327 ( .A(p_input[493]), .B(n26454), .Z(n26283) );
  AND U26328 ( .A(n979), .B(n26455), .Z(n26454) );
  XOR U26329 ( .A(p_input[509]), .B(p_input[493]), .Z(n26455) );
  XNOR U26330 ( .A(n26280), .B(n26450), .Z(n26452) );
  XOR U26331 ( .A(n26456), .B(n26457), .Z(n26280) );
  AND U26332 ( .A(n977), .B(n26458), .Z(n26457) );
  XOR U26333 ( .A(p_input[477]), .B(p_input[461]), .Z(n26458) );
  XOR U26334 ( .A(n26459), .B(n26460), .Z(n26450) );
  AND U26335 ( .A(n26461), .B(n26462), .Z(n26460) );
  XOR U26336 ( .A(n26459), .B(n26295), .Z(n26462) );
  XNOR U26337 ( .A(p_input[492]), .B(n26463), .Z(n26295) );
  AND U26338 ( .A(n979), .B(n26464), .Z(n26463) );
  XOR U26339 ( .A(p_input[508]), .B(p_input[492]), .Z(n26464) );
  XNOR U26340 ( .A(n26292), .B(n26459), .Z(n26461) );
  XOR U26341 ( .A(n26465), .B(n26466), .Z(n26292) );
  AND U26342 ( .A(n977), .B(n26467), .Z(n26466) );
  XOR U26343 ( .A(p_input[476]), .B(p_input[460]), .Z(n26467) );
  XOR U26344 ( .A(n26468), .B(n26469), .Z(n26459) );
  AND U26345 ( .A(n26470), .B(n26471), .Z(n26469) );
  XOR U26346 ( .A(n26468), .B(n26307), .Z(n26471) );
  XNOR U26347 ( .A(p_input[491]), .B(n26472), .Z(n26307) );
  AND U26348 ( .A(n979), .B(n26473), .Z(n26472) );
  XOR U26349 ( .A(p_input[507]), .B(p_input[491]), .Z(n26473) );
  XNOR U26350 ( .A(n26304), .B(n26468), .Z(n26470) );
  XOR U26351 ( .A(n26474), .B(n26475), .Z(n26304) );
  AND U26352 ( .A(n977), .B(n26476), .Z(n26475) );
  XOR U26353 ( .A(p_input[475]), .B(p_input[459]), .Z(n26476) );
  XOR U26354 ( .A(n26477), .B(n26478), .Z(n26468) );
  AND U26355 ( .A(n26479), .B(n26480), .Z(n26478) );
  XOR U26356 ( .A(n26477), .B(n26319), .Z(n26480) );
  XNOR U26357 ( .A(p_input[490]), .B(n26481), .Z(n26319) );
  AND U26358 ( .A(n979), .B(n26482), .Z(n26481) );
  XOR U26359 ( .A(p_input[506]), .B(p_input[490]), .Z(n26482) );
  XNOR U26360 ( .A(n26316), .B(n26477), .Z(n26479) );
  XOR U26361 ( .A(n26483), .B(n26484), .Z(n26316) );
  AND U26362 ( .A(n977), .B(n26485), .Z(n26484) );
  XOR U26363 ( .A(p_input[474]), .B(p_input[458]), .Z(n26485) );
  XOR U26364 ( .A(n26486), .B(n26487), .Z(n26477) );
  AND U26365 ( .A(n26488), .B(n26489), .Z(n26487) );
  XOR U26366 ( .A(n26486), .B(n26331), .Z(n26489) );
  XNOR U26367 ( .A(p_input[489]), .B(n26490), .Z(n26331) );
  AND U26368 ( .A(n979), .B(n26491), .Z(n26490) );
  XOR U26369 ( .A(p_input[505]), .B(p_input[489]), .Z(n26491) );
  XNOR U26370 ( .A(n26328), .B(n26486), .Z(n26488) );
  XOR U26371 ( .A(n26492), .B(n26493), .Z(n26328) );
  AND U26372 ( .A(n977), .B(n26494), .Z(n26493) );
  XOR U26373 ( .A(p_input[473]), .B(p_input[457]), .Z(n26494) );
  XOR U26374 ( .A(n26495), .B(n26496), .Z(n26486) );
  AND U26375 ( .A(n26497), .B(n26498), .Z(n26496) );
  XOR U26376 ( .A(n26495), .B(n26343), .Z(n26498) );
  XNOR U26377 ( .A(p_input[488]), .B(n26499), .Z(n26343) );
  AND U26378 ( .A(n979), .B(n26500), .Z(n26499) );
  XOR U26379 ( .A(p_input[504]), .B(p_input[488]), .Z(n26500) );
  XNOR U26380 ( .A(n26340), .B(n26495), .Z(n26497) );
  XOR U26381 ( .A(n26501), .B(n26502), .Z(n26340) );
  AND U26382 ( .A(n977), .B(n26503), .Z(n26502) );
  XOR U26383 ( .A(p_input[472]), .B(p_input[456]), .Z(n26503) );
  XOR U26384 ( .A(n26504), .B(n26505), .Z(n26495) );
  AND U26385 ( .A(n26506), .B(n26507), .Z(n26505) );
  XOR U26386 ( .A(n26504), .B(n26355), .Z(n26507) );
  XNOR U26387 ( .A(p_input[487]), .B(n26508), .Z(n26355) );
  AND U26388 ( .A(n979), .B(n26509), .Z(n26508) );
  XOR U26389 ( .A(p_input[503]), .B(p_input[487]), .Z(n26509) );
  XNOR U26390 ( .A(n26352), .B(n26504), .Z(n26506) );
  XOR U26391 ( .A(n26510), .B(n26511), .Z(n26352) );
  AND U26392 ( .A(n977), .B(n26512), .Z(n26511) );
  XOR U26393 ( .A(p_input[471]), .B(p_input[455]), .Z(n26512) );
  XOR U26394 ( .A(n26513), .B(n26514), .Z(n26504) );
  AND U26395 ( .A(n26515), .B(n26516), .Z(n26514) );
  XOR U26396 ( .A(n26513), .B(n26367), .Z(n26516) );
  XNOR U26397 ( .A(p_input[486]), .B(n26517), .Z(n26367) );
  AND U26398 ( .A(n979), .B(n26518), .Z(n26517) );
  XOR U26399 ( .A(p_input[502]), .B(p_input[486]), .Z(n26518) );
  XNOR U26400 ( .A(n26364), .B(n26513), .Z(n26515) );
  XOR U26401 ( .A(n26519), .B(n26520), .Z(n26364) );
  AND U26402 ( .A(n977), .B(n26521), .Z(n26520) );
  XOR U26403 ( .A(p_input[470]), .B(p_input[454]), .Z(n26521) );
  XOR U26404 ( .A(n26522), .B(n26523), .Z(n26513) );
  AND U26405 ( .A(n26524), .B(n26525), .Z(n26523) );
  XOR U26406 ( .A(n26522), .B(n26379), .Z(n26525) );
  XNOR U26407 ( .A(p_input[485]), .B(n26526), .Z(n26379) );
  AND U26408 ( .A(n979), .B(n26527), .Z(n26526) );
  XOR U26409 ( .A(p_input[501]), .B(p_input[485]), .Z(n26527) );
  XNOR U26410 ( .A(n26376), .B(n26522), .Z(n26524) );
  XOR U26411 ( .A(n26528), .B(n26529), .Z(n26376) );
  AND U26412 ( .A(n977), .B(n26530), .Z(n26529) );
  XOR U26413 ( .A(p_input[469]), .B(p_input[453]), .Z(n26530) );
  XOR U26414 ( .A(n26531), .B(n26532), .Z(n26522) );
  AND U26415 ( .A(n26533), .B(n26534), .Z(n26532) );
  XOR U26416 ( .A(n26531), .B(n26391), .Z(n26534) );
  XNOR U26417 ( .A(p_input[484]), .B(n26535), .Z(n26391) );
  AND U26418 ( .A(n979), .B(n26536), .Z(n26535) );
  XOR U26419 ( .A(p_input[500]), .B(p_input[484]), .Z(n26536) );
  XNOR U26420 ( .A(n26388), .B(n26531), .Z(n26533) );
  XOR U26421 ( .A(n26537), .B(n26538), .Z(n26388) );
  AND U26422 ( .A(n977), .B(n26539), .Z(n26538) );
  XOR U26423 ( .A(p_input[468]), .B(p_input[452]), .Z(n26539) );
  XOR U26424 ( .A(n26540), .B(n26541), .Z(n26531) );
  AND U26425 ( .A(n26542), .B(n26543), .Z(n26541) );
  XOR U26426 ( .A(n26540), .B(n26403), .Z(n26543) );
  XNOR U26427 ( .A(p_input[483]), .B(n26544), .Z(n26403) );
  AND U26428 ( .A(n979), .B(n26545), .Z(n26544) );
  XOR U26429 ( .A(p_input[499]), .B(p_input[483]), .Z(n26545) );
  XNOR U26430 ( .A(n26400), .B(n26540), .Z(n26542) );
  XOR U26431 ( .A(n26546), .B(n26547), .Z(n26400) );
  AND U26432 ( .A(n977), .B(n26548), .Z(n26547) );
  XOR U26433 ( .A(p_input[467]), .B(p_input[451]), .Z(n26548) );
  XOR U26434 ( .A(n26549), .B(n26550), .Z(n26540) );
  AND U26435 ( .A(n26551), .B(n26552), .Z(n26550) );
  XOR U26436 ( .A(n26549), .B(n26415), .Z(n26552) );
  XNOR U26437 ( .A(p_input[482]), .B(n26553), .Z(n26415) );
  AND U26438 ( .A(n979), .B(n26554), .Z(n26553) );
  XOR U26439 ( .A(p_input[498]), .B(p_input[482]), .Z(n26554) );
  XNOR U26440 ( .A(n26412), .B(n26549), .Z(n26551) );
  XOR U26441 ( .A(n26555), .B(n26556), .Z(n26412) );
  AND U26442 ( .A(n977), .B(n26557), .Z(n26556) );
  XOR U26443 ( .A(p_input[466]), .B(p_input[450]), .Z(n26557) );
  XOR U26444 ( .A(n26558), .B(n26559), .Z(n26549) );
  AND U26445 ( .A(n26560), .B(n26561), .Z(n26559) );
  XNOR U26446 ( .A(n26562), .B(n26428), .Z(n26561) );
  XNOR U26447 ( .A(p_input[481]), .B(n26563), .Z(n26428) );
  AND U26448 ( .A(n979), .B(n26564), .Z(n26563) );
  XNOR U26449 ( .A(p_input[497]), .B(n26565), .Z(n26564) );
  IV U26450 ( .A(p_input[481]), .Z(n26565) );
  XNOR U26451 ( .A(n26425), .B(n26558), .Z(n26560) );
  XNOR U26452 ( .A(p_input[449]), .B(n26566), .Z(n26425) );
  AND U26453 ( .A(n977), .B(n26567), .Z(n26566) );
  XOR U26454 ( .A(p_input[465]), .B(p_input[449]), .Z(n26567) );
  IV U26455 ( .A(n26562), .Z(n26558) );
  AND U26456 ( .A(n26433), .B(n26436), .Z(n26562) );
  XOR U26457 ( .A(p_input[480]), .B(n26568), .Z(n26436) );
  AND U26458 ( .A(n979), .B(n26569), .Z(n26568) );
  XOR U26459 ( .A(p_input[496]), .B(p_input[480]), .Z(n26569) );
  XOR U26460 ( .A(n26570), .B(n26571), .Z(n979) );
  AND U26461 ( .A(n26572), .B(n26573), .Z(n26571) );
  XNOR U26462 ( .A(p_input[511]), .B(n26570), .Z(n26573) );
  XOR U26463 ( .A(n26570), .B(p_input[495]), .Z(n26572) );
  XOR U26464 ( .A(n26574), .B(n26575), .Z(n26570) );
  AND U26465 ( .A(n26576), .B(n26577), .Z(n26575) );
  XNOR U26466 ( .A(p_input[510]), .B(n26574), .Z(n26577) );
  XOR U26467 ( .A(n26574), .B(p_input[494]), .Z(n26576) );
  XOR U26468 ( .A(n26578), .B(n26579), .Z(n26574) );
  AND U26469 ( .A(n26580), .B(n26581), .Z(n26579) );
  XNOR U26470 ( .A(p_input[509]), .B(n26578), .Z(n26581) );
  XOR U26471 ( .A(n26578), .B(p_input[493]), .Z(n26580) );
  XOR U26472 ( .A(n26582), .B(n26583), .Z(n26578) );
  AND U26473 ( .A(n26584), .B(n26585), .Z(n26583) );
  XNOR U26474 ( .A(p_input[508]), .B(n26582), .Z(n26585) );
  XOR U26475 ( .A(n26582), .B(p_input[492]), .Z(n26584) );
  XOR U26476 ( .A(n26586), .B(n26587), .Z(n26582) );
  AND U26477 ( .A(n26588), .B(n26589), .Z(n26587) );
  XNOR U26478 ( .A(p_input[507]), .B(n26586), .Z(n26589) );
  XOR U26479 ( .A(n26586), .B(p_input[491]), .Z(n26588) );
  XOR U26480 ( .A(n26590), .B(n26591), .Z(n26586) );
  AND U26481 ( .A(n26592), .B(n26593), .Z(n26591) );
  XNOR U26482 ( .A(p_input[506]), .B(n26590), .Z(n26593) );
  XOR U26483 ( .A(n26590), .B(p_input[490]), .Z(n26592) );
  XOR U26484 ( .A(n26594), .B(n26595), .Z(n26590) );
  AND U26485 ( .A(n26596), .B(n26597), .Z(n26595) );
  XNOR U26486 ( .A(p_input[505]), .B(n26594), .Z(n26597) );
  XOR U26487 ( .A(n26594), .B(p_input[489]), .Z(n26596) );
  XOR U26488 ( .A(n26598), .B(n26599), .Z(n26594) );
  AND U26489 ( .A(n26600), .B(n26601), .Z(n26599) );
  XNOR U26490 ( .A(p_input[504]), .B(n26598), .Z(n26601) );
  XOR U26491 ( .A(n26598), .B(p_input[488]), .Z(n26600) );
  XOR U26492 ( .A(n26602), .B(n26603), .Z(n26598) );
  AND U26493 ( .A(n26604), .B(n26605), .Z(n26603) );
  XNOR U26494 ( .A(p_input[503]), .B(n26602), .Z(n26605) );
  XOR U26495 ( .A(n26602), .B(p_input[487]), .Z(n26604) );
  XOR U26496 ( .A(n26606), .B(n26607), .Z(n26602) );
  AND U26497 ( .A(n26608), .B(n26609), .Z(n26607) );
  XNOR U26498 ( .A(p_input[502]), .B(n26606), .Z(n26609) );
  XOR U26499 ( .A(n26606), .B(p_input[486]), .Z(n26608) );
  XOR U26500 ( .A(n26610), .B(n26611), .Z(n26606) );
  AND U26501 ( .A(n26612), .B(n26613), .Z(n26611) );
  XNOR U26502 ( .A(p_input[501]), .B(n26610), .Z(n26613) );
  XOR U26503 ( .A(n26610), .B(p_input[485]), .Z(n26612) );
  XOR U26504 ( .A(n26614), .B(n26615), .Z(n26610) );
  AND U26505 ( .A(n26616), .B(n26617), .Z(n26615) );
  XNOR U26506 ( .A(p_input[500]), .B(n26614), .Z(n26617) );
  XOR U26507 ( .A(n26614), .B(p_input[484]), .Z(n26616) );
  XOR U26508 ( .A(n26618), .B(n26619), .Z(n26614) );
  AND U26509 ( .A(n26620), .B(n26621), .Z(n26619) );
  XNOR U26510 ( .A(p_input[499]), .B(n26618), .Z(n26621) );
  XOR U26511 ( .A(n26618), .B(p_input[483]), .Z(n26620) );
  XOR U26512 ( .A(n26622), .B(n26623), .Z(n26618) );
  AND U26513 ( .A(n26624), .B(n26625), .Z(n26623) );
  XNOR U26514 ( .A(p_input[498]), .B(n26622), .Z(n26625) );
  XOR U26515 ( .A(n26622), .B(p_input[482]), .Z(n26624) );
  XNOR U26516 ( .A(n26626), .B(n26627), .Z(n26622) );
  AND U26517 ( .A(n26628), .B(n26629), .Z(n26627) );
  XOR U26518 ( .A(p_input[497]), .B(n26626), .Z(n26629) );
  XNOR U26519 ( .A(p_input[481]), .B(n26626), .Z(n26628) );
  AND U26520 ( .A(p_input[496]), .B(n26630), .Z(n26626) );
  IV U26521 ( .A(p_input[480]), .Z(n26630) );
  XNOR U26522 ( .A(p_input[448]), .B(n26631), .Z(n26433) );
  AND U26523 ( .A(n977), .B(n26632), .Z(n26631) );
  XOR U26524 ( .A(p_input[464]), .B(p_input[448]), .Z(n26632) );
  XOR U26525 ( .A(n26633), .B(n26634), .Z(n977) );
  AND U26526 ( .A(n26635), .B(n26636), .Z(n26634) );
  XNOR U26527 ( .A(p_input[479]), .B(n26633), .Z(n26636) );
  XOR U26528 ( .A(n26633), .B(p_input[463]), .Z(n26635) );
  XOR U26529 ( .A(n26637), .B(n26638), .Z(n26633) );
  AND U26530 ( .A(n26639), .B(n26640), .Z(n26638) );
  XNOR U26531 ( .A(p_input[478]), .B(n26637), .Z(n26640) );
  XNOR U26532 ( .A(n26637), .B(n26447), .Z(n26639) );
  IV U26533 ( .A(p_input[462]), .Z(n26447) );
  XOR U26534 ( .A(n26641), .B(n26642), .Z(n26637) );
  AND U26535 ( .A(n26643), .B(n26644), .Z(n26642) );
  XNOR U26536 ( .A(p_input[477]), .B(n26641), .Z(n26644) );
  XNOR U26537 ( .A(n26641), .B(n26456), .Z(n26643) );
  IV U26538 ( .A(p_input[461]), .Z(n26456) );
  XOR U26539 ( .A(n26645), .B(n26646), .Z(n26641) );
  AND U26540 ( .A(n26647), .B(n26648), .Z(n26646) );
  XNOR U26541 ( .A(p_input[476]), .B(n26645), .Z(n26648) );
  XNOR U26542 ( .A(n26645), .B(n26465), .Z(n26647) );
  IV U26543 ( .A(p_input[460]), .Z(n26465) );
  XOR U26544 ( .A(n26649), .B(n26650), .Z(n26645) );
  AND U26545 ( .A(n26651), .B(n26652), .Z(n26650) );
  XNOR U26546 ( .A(p_input[475]), .B(n26649), .Z(n26652) );
  XNOR U26547 ( .A(n26649), .B(n26474), .Z(n26651) );
  IV U26548 ( .A(p_input[459]), .Z(n26474) );
  XOR U26549 ( .A(n26653), .B(n26654), .Z(n26649) );
  AND U26550 ( .A(n26655), .B(n26656), .Z(n26654) );
  XNOR U26551 ( .A(p_input[474]), .B(n26653), .Z(n26656) );
  XNOR U26552 ( .A(n26653), .B(n26483), .Z(n26655) );
  IV U26553 ( .A(p_input[458]), .Z(n26483) );
  XOR U26554 ( .A(n26657), .B(n26658), .Z(n26653) );
  AND U26555 ( .A(n26659), .B(n26660), .Z(n26658) );
  XNOR U26556 ( .A(p_input[473]), .B(n26657), .Z(n26660) );
  XNOR U26557 ( .A(n26657), .B(n26492), .Z(n26659) );
  IV U26558 ( .A(p_input[457]), .Z(n26492) );
  XOR U26559 ( .A(n26661), .B(n26662), .Z(n26657) );
  AND U26560 ( .A(n26663), .B(n26664), .Z(n26662) );
  XNOR U26561 ( .A(p_input[472]), .B(n26661), .Z(n26664) );
  XNOR U26562 ( .A(n26661), .B(n26501), .Z(n26663) );
  IV U26563 ( .A(p_input[456]), .Z(n26501) );
  XOR U26564 ( .A(n26665), .B(n26666), .Z(n26661) );
  AND U26565 ( .A(n26667), .B(n26668), .Z(n26666) );
  XNOR U26566 ( .A(p_input[471]), .B(n26665), .Z(n26668) );
  XNOR U26567 ( .A(n26665), .B(n26510), .Z(n26667) );
  IV U26568 ( .A(p_input[455]), .Z(n26510) );
  XOR U26569 ( .A(n26669), .B(n26670), .Z(n26665) );
  AND U26570 ( .A(n26671), .B(n26672), .Z(n26670) );
  XNOR U26571 ( .A(p_input[470]), .B(n26669), .Z(n26672) );
  XNOR U26572 ( .A(n26669), .B(n26519), .Z(n26671) );
  IV U26573 ( .A(p_input[454]), .Z(n26519) );
  XOR U26574 ( .A(n26673), .B(n26674), .Z(n26669) );
  AND U26575 ( .A(n26675), .B(n26676), .Z(n26674) );
  XNOR U26576 ( .A(p_input[469]), .B(n26673), .Z(n26676) );
  XNOR U26577 ( .A(n26673), .B(n26528), .Z(n26675) );
  IV U26578 ( .A(p_input[453]), .Z(n26528) );
  XOR U26579 ( .A(n26677), .B(n26678), .Z(n26673) );
  AND U26580 ( .A(n26679), .B(n26680), .Z(n26678) );
  XNOR U26581 ( .A(p_input[468]), .B(n26677), .Z(n26680) );
  XNOR U26582 ( .A(n26677), .B(n26537), .Z(n26679) );
  IV U26583 ( .A(p_input[452]), .Z(n26537) );
  XOR U26584 ( .A(n26681), .B(n26682), .Z(n26677) );
  AND U26585 ( .A(n26683), .B(n26684), .Z(n26682) );
  XNOR U26586 ( .A(p_input[467]), .B(n26681), .Z(n26684) );
  XNOR U26587 ( .A(n26681), .B(n26546), .Z(n26683) );
  IV U26588 ( .A(p_input[451]), .Z(n26546) );
  XOR U26589 ( .A(n26685), .B(n26686), .Z(n26681) );
  AND U26590 ( .A(n26687), .B(n26688), .Z(n26686) );
  XNOR U26591 ( .A(p_input[466]), .B(n26685), .Z(n26688) );
  XNOR U26592 ( .A(n26685), .B(n26555), .Z(n26687) );
  IV U26593 ( .A(p_input[450]), .Z(n26555) );
  XNOR U26594 ( .A(n26689), .B(n26690), .Z(n26685) );
  AND U26595 ( .A(n26691), .B(n26692), .Z(n26690) );
  XOR U26596 ( .A(p_input[465]), .B(n26689), .Z(n26692) );
  XNOR U26597 ( .A(p_input[449]), .B(n26689), .Z(n26691) );
  AND U26598 ( .A(p_input[464]), .B(n26693), .Z(n26689) );
  IV U26599 ( .A(p_input[448]), .Z(n26693) );
  XOR U26600 ( .A(n26694), .B(n26695), .Z(n26252) );
  AND U26601 ( .A(n569), .B(n26696), .Z(n26695) );
  XNOR U26602 ( .A(n26697), .B(n26694), .Z(n26696) );
  XOR U26603 ( .A(n26698), .B(n26699), .Z(n569) );
  AND U26604 ( .A(n26700), .B(n26701), .Z(n26699) );
  XNOR U26605 ( .A(n26262), .B(n26698), .Z(n26701) );
  AND U26606 ( .A(p_input[447]), .B(p_input[431]), .Z(n26262) );
  XOR U26607 ( .A(n26698), .B(n26263), .Z(n26700) );
  AND U26608 ( .A(p_input[415]), .B(p_input[399]), .Z(n26263) );
  XOR U26609 ( .A(n26702), .B(n26703), .Z(n26698) );
  AND U26610 ( .A(n26704), .B(n26705), .Z(n26703) );
  XOR U26611 ( .A(n26702), .B(n26275), .Z(n26705) );
  XNOR U26612 ( .A(p_input[430]), .B(n26706), .Z(n26275) );
  AND U26613 ( .A(n983), .B(n26707), .Z(n26706) );
  XOR U26614 ( .A(p_input[446]), .B(p_input[430]), .Z(n26707) );
  XNOR U26615 ( .A(n26272), .B(n26702), .Z(n26704) );
  XOR U26616 ( .A(n26708), .B(n26709), .Z(n26272) );
  AND U26617 ( .A(n980), .B(n26710), .Z(n26709) );
  XOR U26618 ( .A(p_input[414]), .B(p_input[398]), .Z(n26710) );
  XOR U26619 ( .A(n26711), .B(n26712), .Z(n26702) );
  AND U26620 ( .A(n26713), .B(n26714), .Z(n26712) );
  XOR U26621 ( .A(n26711), .B(n26287), .Z(n26714) );
  XNOR U26622 ( .A(p_input[429]), .B(n26715), .Z(n26287) );
  AND U26623 ( .A(n983), .B(n26716), .Z(n26715) );
  XOR U26624 ( .A(p_input[445]), .B(p_input[429]), .Z(n26716) );
  XNOR U26625 ( .A(n26284), .B(n26711), .Z(n26713) );
  XOR U26626 ( .A(n26717), .B(n26718), .Z(n26284) );
  AND U26627 ( .A(n980), .B(n26719), .Z(n26718) );
  XOR U26628 ( .A(p_input[413]), .B(p_input[397]), .Z(n26719) );
  XOR U26629 ( .A(n26720), .B(n26721), .Z(n26711) );
  AND U26630 ( .A(n26722), .B(n26723), .Z(n26721) );
  XOR U26631 ( .A(n26720), .B(n26299), .Z(n26723) );
  XNOR U26632 ( .A(p_input[428]), .B(n26724), .Z(n26299) );
  AND U26633 ( .A(n983), .B(n26725), .Z(n26724) );
  XOR U26634 ( .A(p_input[444]), .B(p_input[428]), .Z(n26725) );
  XNOR U26635 ( .A(n26296), .B(n26720), .Z(n26722) );
  XOR U26636 ( .A(n26726), .B(n26727), .Z(n26296) );
  AND U26637 ( .A(n980), .B(n26728), .Z(n26727) );
  XOR U26638 ( .A(p_input[412]), .B(p_input[396]), .Z(n26728) );
  XOR U26639 ( .A(n26729), .B(n26730), .Z(n26720) );
  AND U26640 ( .A(n26731), .B(n26732), .Z(n26730) );
  XOR U26641 ( .A(n26729), .B(n26311), .Z(n26732) );
  XNOR U26642 ( .A(p_input[427]), .B(n26733), .Z(n26311) );
  AND U26643 ( .A(n983), .B(n26734), .Z(n26733) );
  XOR U26644 ( .A(p_input[443]), .B(p_input[427]), .Z(n26734) );
  XNOR U26645 ( .A(n26308), .B(n26729), .Z(n26731) );
  XOR U26646 ( .A(n26735), .B(n26736), .Z(n26308) );
  AND U26647 ( .A(n980), .B(n26737), .Z(n26736) );
  XOR U26648 ( .A(p_input[411]), .B(p_input[395]), .Z(n26737) );
  XOR U26649 ( .A(n26738), .B(n26739), .Z(n26729) );
  AND U26650 ( .A(n26740), .B(n26741), .Z(n26739) );
  XOR U26651 ( .A(n26738), .B(n26323), .Z(n26741) );
  XNOR U26652 ( .A(p_input[426]), .B(n26742), .Z(n26323) );
  AND U26653 ( .A(n983), .B(n26743), .Z(n26742) );
  XOR U26654 ( .A(p_input[442]), .B(p_input[426]), .Z(n26743) );
  XNOR U26655 ( .A(n26320), .B(n26738), .Z(n26740) );
  XOR U26656 ( .A(n26744), .B(n26745), .Z(n26320) );
  AND U26657 ( .A(n980), .B(n26746), .Z(n26745) );
  XOR U26658 ( .A(p_input[410]), .B(p_input[394]), .Z(n26746) );
  XOR U26659 ( .A(n26747), .B(n26748), .Z(n26738) );
  AND U26660 ( .A(n26749), .B(n26750), .Z(n26748) );
  XOR U26661 ( .A(n26747), .B(n26335), .Z(n26750) );
  XNOR U26662 ( .A(p_input[425]), .B(n26751), .Z(n26335) );
  AND U26663 ( .A(n983), .B(n26752), .Z(n26751) );
  XOR U26664 ( .A(p_input[441]), .B(p_input[425]), .Z(n26752) );
  XNOR U26665 ( .A(n26332), .B(n26747), .Z(n26749) );
  XOR U26666 ( .A(n26753), .B(n26754), .Z(n26332) );
  AND U26667 ( .A(n980), .B(n26755), .Z(n26754) );
  XOR U26668 ( .A(p_input[409]), .B(p_input[393]), .Z(n26755) );
  XOR U26669 ( .A(n26756), .B(n26757), .Z(n26747) );
  AND U26670 ( .A(n26758), .B(n26759), .Z(n26757) );
  XOR U26671 ( .A(n26756), .B(n26347), .Z(n26759) );
  XNOR U26672 ( .A(p_input[424]), .B(n26760), .Z(n26347) );
  AND U26673 ( .A(n983), .B(n26761), .Z(n26760) );
  XOR U26674 ( .A(p_input[440]), .B(p_input[424]), .Z(n26761) );
  XNOR U26675 ( .A(n26344), .B(n26756), .Z(n26758) );
  XOR U26676 ( .A(n26762), .B(n26763), .Z(n26344) );
  AND U26677 ( .A(n980), .B(n26764), .Z(n26763) );
  XOR U26678 ( .A(p_input[408]), .B(p_input[392]), .Z(n26764) );
  XOR U26679 ( .A(n26765), .B(n26766), .Z(n26756) );
  AND U26680 ( .A(n26767), .B(n26768), .Z(n26766) );
  XOR U26681 ( .A(n26765), .B(n26359), .Z(n26768) );
  XNOR U26682 ( .A(p_input[423]), .B(n26769), .Z(n26359) );
  AND U26683 ( .A(n983), .B(n26770), .Z(n26769) );
  XOR U26684 ( .A(p_input[439]), .B(p_input[423]), .Z(n26770) );
  XNOR U26685 ( .A(n26356), .B(n26765), .Z(n26767) );
  XOR U26686 ( .A(n26771), .B(n26772), .Z(n26356) );
  AND U26687 ( .A(n980), .B(n26773), .Z(n26772) );
  XOR U26688 ( .A(p_input[407]), .B(p_input[391]), .Z(n26773) );
  XOR U26689 ( .A(n26774), .B(n26775), .Z(n26765) );
  AND U26690 ( .A(n26776), .B(n26777), .Z(n26775) );
  XOR U26691 ( .A(n26774), .B(n26371), .Z(n26777) );
  XNOR U26692 ( .A(p_input[422]), .B(n26778), .Z(n26371) );
  AND U26693 ( .A(n983), .B(n26779), .Z(n26778) );
  XOR U26694 ( .A(p_input[438]), .B(p_input[422]), .Z(n26779) );
  XNOR U26695 ( .A(n26368), .B(n26774), .Z(n26776) );
  XOR U26696 ( .A(n26780), .B(n26781), .Z(n26368) );
  AND U26697 ( .A(n980), .B(n26782), .Z(n26781) );
  XOR U26698 ( .A(p_input[406]), .B(p_input[390]), .Z(n26782) );
  XOR U26699 ( .A(n26783), .B(n26784), .Z(n26774) );
  AND U26700 ( .A(n26785), .B(n26786), .Z(n26784) );
  XOR U26701 ( .A(n26783), .B(n26383), .Z(n26786) );
  XNOR U26702 ( .A(p_input[421]), .B(n26787), .Z(n26383) );
  AND U26703 ( .A(n983), .B(n26788), .Z(n26787) );
  XOR U26704 ( .A(p_input[437]), .B(p_input[421]), .Z(n26788) );
  XNOR U26705 ( .A(n26380), .B(n26783), .Z(n26785) );
  XOR U26706 ( .A(n26789), .B(n26790), .Z(n26380) );
  AND U26707 ( .A(n980), .B(n26791), .Z(n26790) );
  XOR U26708 ( .A(p_input[405]), .B(p_input[389]), .Z(n26791) );
  XOR U26709 ( .A(n26792), .B(n26793), .Z(n26783) );
  AND U26710 ( .A(n26794), .B(n26795), .Z(n26793) );
  XOR U26711 ( .A(n26792), .B(n26395), .Z(n26795) );
  XNOR U26712 ( .A(p_input[420]), .B(n26796), .Z(n26395) );
  AND U26713 ( .A(n983), .B(n26797), .Z(n26796) );
  XOR U26714 ( .A(p_input[436]), .B(p_input[420]), .Z(n26797) );
  XNOR U26715 ( .A(n26392), .B(n26792), .Z(n26794) );
  XOR U26716 ( .A(n26798), .B(n26799), .Z(n26392) );
  AND U26717 ( .A(n980), .B(n26800), .Z(n26799) );
  XOR U26718 ( .A(p_input[404]), .B(p_input[388]), .Z(n26800) );
  XOR U26719 ( .A(n26801), .B(n26802), .Z(n26792) );
  AND U26720 ( .A(n26803), .B(n26804), .Z(n26802) );
  XOR U26721 ( .A(n26801), .B(n26407), .Z(n26804) );
  XNOR U26722 ( .A(p_input[419]), .B(n26805), .Z(n26407) );
  AND U26723 ( .A(n983), .B(n26806), .Z(n26805) );
  XOR U26724 ( .A(p_input[435]), .B(p_input[419]), .Z(n26806) );
  XNOR U26725 ( .A(n26404), .B(n26801), .Z(n26803) );
  XOR U26726 ( .A(n26807), .B(n26808), .Z(n26404) );
  AND U26727 ( .A(n980), .B(n26809), .Z(n26808) );
  XOR U26728 ( .A(p_input[403]), .B(p_input[387]), .Z(n26809) );
  XOR U26729 ( .A(n26810), .B(n26811), .Z(n26801) );
  AND U26730 ( .A(n26812), .B(n26813), .Z(n26811) );
  XOR U26731 ( .A(n26810), .B(n26419), .Z(n26813) );
  XNOR U26732 ( .A(p_input[418]), .B(n26814), .Z(n26419) );
  AND U26733 ( .A(n983), .B(n26815), .Z(n26814) );
  XOR U26734 ( .A(p_input[434]), .B(p_input[418]), .Z(n26815) );
  XNOR U26735 ( .A(n26416), .B(n26810), .Z(n26812) );
  XOR U26736 ( .A(n26816), .B(n26817), .Z(n26416) );
  AND U26737 ( .A(n980), .B(n26818), .Z(n26817) );
  XOR U26738 ( .A(p_input[402]), .B(p_input[386]), .Z(n26818) );
  XOR U26739 ( .A(n26819), .B(n26820), .Z(n26810) );
  AND U26740 ( .A(n26821), .B(n26822), .Z(n26820) );
  XNOR U26741 ( .A(n26823), .B(n26432), .Z(n26822) );
  XNOR U26742 ( .A(p_input[417]), .B(n26824), .Z(n26432) );
  AND U26743 ( .A(n983), .B(n26825), .Z(n26824) );
  XNOR U26744 ( .A(p_input[433]), .B(n26826), .Z(n26825) );
  IV U26745 ( .A(p_input[417]), .Z(n26826) );
  XNOR U26746 ( .A(n26429), .B(n26819), .Z(n26821) );
  XNOR U26747 ( .A(p_input[385]), .B(n26827), .Z(n26429) );
  AND U26748 ( .A(n980), .B(n26828), .Z(n26827) );
  XOR U26749 ( .A(p_input[401]), .B(p_input[385]), .Z(n26828) );
  IV U26750 ( .A(n26823), .Z(n26819) );
  AND U26751 ( .A(n26694), .B(n26697), .Z(n26823) );
  XOR U26752 ( .A(p_input[416]), .B(n26829), .Z(n26697) );
  AND U26753 ( .A(n983), .B(n26830), .Z(n26829) );
  XOR U26754 ( .A(p_input[432]), .B(p_input[416]), .Z(n26830) );
  XOR U26755 ( .A(n26831), .B(n26832), .Z(n983) );
  AND U26756 ( .A(n26833), .B(n26834), .Z(n26832) );
  XNOR U26757 ( .A(p_input[447]), .B(n26831), .Z(n26834) );
  XOR U26758 ( .A(n26831), .B(p_input[431]), .Z(n26833) );
  XOR U26759 ( .A(n26835), .B(n26836), .Z(n26831) );
  AND U26760 ( .A(n26837), .B(n26838), .Z(n26836) );
  XNOR U26761 ( .A(p_input[446]), .B(n26835), .Z(n26838) );
  XOR U26762 ( .A(n26835), .B(p_input[430]), .Z(n26837) );
  XOR U26763 ( .A(n26839), .B(n26840), .Z(n26835) );
  AND U26764 ( .A(n26841), .B(n26842), .Z(n26840) );
  XNOR U26765 ( .A(p_input[445]), .B(n26839), .Z(n26842) );
  XOR U26766 ( .A(n26839), .B(p_input[429]), .Z(n26841) );
  XOR U26767 ( .A(n26843), .B(n26844), .Z(n26839) );
  AND U26768 ( .A(n26845), .B(n26846), .Z(n26844) );
  XNOR U26769 ( .A(p_input[444]), .B(n26843), .Z(n26846) );
  XOR U26770 ( .A(n26843), .B(p_input[428]), .Z(n26845) );
  XOR U26771 ( .A(n26847), .B(n26848), .Z(n26843) );
  AND U26772 ( .A(n26849), .B(n26850), .Z(n26848) );
  XNOR U26773 ( .A(p_input[443]), .B(n26847), .Z(n26850) );
  XOR U26774 ( .A(n26847), .B(p_input[427]), .Z(n26849) );
  XOR U26775 ( .A(n26851), .B(n26852), .Z(n26847) );
  AND U26776 ( .A(n26853), .B(n26854), .Z(n26852) );
  XNOR U26777 ( .A(p_input[442]), .B(n26851), .Z(n26854) );
  XOR U26778 ( .A(n26851), .B(p_input[426]), .Z(n26853) );
  XOR U26779 ( .A(n26855), .B(n26856), .Z(n26851) );
  AND U26780 ( .A(n26857), .B(n26858), .Z(n26856) );
  XNOR U26781 ( .A(p_input[441]), .B(n26855), .Z(n26858) );
  XOR U26782 ( .A(n26855), .B(p_input[425]), .Z(n26857) );
  XOR U26783 ( .A(n26859), .B(n26860), .Z(n26855) );
  AND U26784 ( .A(n26861), .B(n26862), .Z(n26860) );
  XNOR U26785 ( .A(p_input[440]), .B(n26859), .Z(n26862) );
  XOR U26786 ( .A(n26859), .B(p_input[424]), .Z(n26861) );
  XOR U26787 ( .A(n26863), .B(n26864), .Z(n26859) );
  AND U26788 ( .A(n26865), .B(n26866), .Z(n26864) );
  XNOR U26789 ( .A(p_input[439]), .B(n26863), .Z(n26866) );
  XOR U26790 ( .A(n26863), .B(p_input[423]), .Z(n26865) );
  XOR U26791 ( .A(n26867), .B(n26868), .Z(n26863) );
  AND U26792 ( .A(n26869), .B(n26870), .Z(n26868) );
  XNOR U26793 ( .A(p_input[438]), .B(n26867), .Z(n26870) );
  XOR U26794 ( .A(n26867), .B(p_input[422]), .Z(n26869) );
  XOR U26795 ( .A(n26871), .B(n26872), .Z(n26867) );
  AND U26796 ( .A(n26873), .B(n26874), .Z(n26872) );
  XNOR U26797 ( .A(p_input[437]), .B(n26871), .Z(n26874) );
  XOR U26798 ( .A(n26871), .B(p_input[421]), .Z(n26873) );
  XOR U26799 ( .A(n26875), .B(n26876), .Z(n26871) );
  AND U26800 ( .A(n26877), .B(n26878), .Z(n26876) );
  XNOR U26801 ( .A(p_input[436]), .B(n26875), .Z(n26878) );
  XOR U26802 ( .A(n26875), .B(p_input[420]), .Z(n26877) );
  XOR U26803 ( .A(n26879), .B(n26880), .Z(n26875) );
  AND U26804 ( .A(n26881), .B(n26882), .Z(n26880) );
  XNOR U26805 ( .A(p_input[435]), .B(n26879), .Z(n26882) );
  XOR U26806 ( .A(n26879), .B(p_input[419]), .Z(n26881) );
  XOR U26807 ( .A(n26883), .B(n26884), .Z(n26879) );
  AND U26808 ( .A(n26885), .B(n26886), .Z(n26884) );
  XNOR U26809 ( .A(p_input[434]), .B(n26883), .Z(n26886) );
  XOR U26810 ( .A(n26883), .B(p_input[418]), .Z(n26885) );
  XNOR U26811 ( .A(n26887), .B(n26888), .Z(n26883) );
  AND U26812 ( .A(n26889), .B(n26890), .Z(n26888) );
  XOR U26813 ( .A(p_input[433]), .B(n26887), .Z(n26890) );
  XNOR U26814 ( .A(p_input[417]), .B(n26887), .Z(n26889) );
  AND U26815 ( .A(p_input[432]), .B(n26891), .Z(n26887) );
  IV U26816 ( .A(p_input[416]), .Z(n26891) );
  XNOR U26817 ( .A(p_input[384]), .B(n26892), .Z(n26694) );
  AND U26818 ( .A(n980), .B(n26893), .Z(n26892) );
  XOR U26819 ( .A(p_input[400]), .B(p_input[384]), .Z(n26893) );
  XOR U26820 ( .A(n26894), .B(n26895), .Z(n980) );
  AND U26821 ( .A(n26896), .B(n26897), .Z(n26895) );
  XNOR U26822 ( .A(p_input[415]), .B(n26894), .Z(n26897) );
  XOR U26823 ( .A(n26894), .B(p_input[399]), .Z(n26896) );
  XOR U26824 ( .A(n26898), .B(n26899), .Z(n26894) );
  AND U26825 ( .A(n26900), .B(n26901), .Z(n26899) );
  XNOR U26826 ( .A(p_input[414]), .B(n26898), .Z(n26901) );
  XNOR U26827 ( .A(n26898), .B(n26708), .Z(n26900) );
  IV U26828 ( .A(p_input[398]), .Z(n26708) );
  XOR U26829 ( .A(n26902), .B(n26903), .Z(n26898) );
  AND U26830 ( .A(n26904), .B(n26905), .Z(n26903) );
  XNOR U26831 ( .A(p_input[413]), .B(n26902), .Z(n26905) );
  XNOR U26832 ( .A(n26902), .B(n26717), .Z(n26904) );
  IV U26833 ( .A(p_input[397]), .Z(n26717) );
  XOR U26834 ( .A(n26906), .B(n26907), .Z(n26902) );
  AND U26835 ( .A(n26908), .B(n26909), .Z(n26907) );
  XNOR U26836 ( .A(p_input[412]), .B(n26906), .Z(n26909) );
  XNOR U26837 ( .A(n26906), .B(n26726), .Z(n26908) );
  IV U26838 ( .A(p_input[396]), .Z(n26726) );
  XOR U26839 ( .A(n26910), .B(n26911), .Z(n26906) );
  AND U26840 ( .A(n26912), .B(n26913), .Z(n26911) );
  XNOR U26841 ( .A(p_input[411]), .B(n26910), .Z(n26913) );
  XNOR U26842 ( .A(n26910), .B(n26735), .Z(n26912) );
  IV U26843 ( .A(p_input[395]), .Z(n26735) );
  XOR U26844 ( .A(n26914), .B(n26915), .Z(n26910) );
  AND U26845 ( .A(n26916), .B(n26917), .Z(n26915) );
  XNOR U26846 ( .A(p_input[410]), .B(n26914), .Z(n26917) );
  XNOR U26847 ( .A(n26914), .B(n26744), .Z(n26916) );
  IV U26848 ( .A(p_input[394]), .Z(n26744) );
  XOR U26849 ( .A(n26918), .B(n26919), .Z(n26914) );
  AND U26850 ( .A(n26920), .B(n26921), .Z(n26919) );
  XNOR U26851 ( .A(p_input[409]), .B(n26918), .Z(n26921) );
  XNOR U26852 ( .A(n26918), .B(n26753), .Z(n26920) );
  IV U26853 ( .A(p_input[393]), .Z(n26753) );
  XOR U26854 ( .A(n26922), .B(n26923), .Z(n26918) );
  AND U26855 ( .A(n26924), .B(n26925), .Z(n26923) );
  XNOR U26856 ( .A(p_input[408]), .B(n26922), .Z(n26925) );
  XNOR U26857 ( .A(n26922), .B(n26762), .Z(n26924) );
  IV U26858 ( .A(p_input[392]), .Z(n26762) );
  XOR U26859 ( .A(n26926), .B(n26927), .Z(n26922) );
  AND U26860 ( .A(n26928), .B(n26929), .Z(n26927) );
  XNOR U26861 ( .A(p_input[407]), .B(n26926), .Z(n26929) );
  XNOR U26862 ( .A(n26926), .B(n26771), .Z(n26928) );
  IV U26863 ( .A(p_input[391]), .Z(n26771) );
  XOR U26864 ( .A(n26930), .B(n26931), .Z(n26926) );
  AND U26865 ( .A(n26932), .B(n26933), .Z(n26931) );
  XNOR U26866 ( .A(p_input[406]), .B(n26930), .Z(n26933) );
  XNOR U26867 ( .A(n26930), .B(n26780), .Z(n26932) );
  IV U26868 ( .A(p_input[390]), .Z(n26780) );
  XOR U26869 ( .A(n26934), .B(n26935), .Z(n26930) );
  AND U26870 ( .A(n26936), .B(n26937), .Z(n26935) );
  XNOR U26871 ( .A(p_input[405]), .B(n26934), .Z(n26937) );
  XNOR U26872 ( .A(n26934), .B(n26789), .Z(n26936) );
  IV U26873 ( .A(p_input[389]), .Z(n26789) );
  XOR U26874 ( .A(n26938), .B(n26939), .Z(n26934) );
  AND U26875 ( .A(n26940), .B(n26941), .Z(n26939) );
  XNOR U26876 ( .A(p_input[404]), .B(n26938), .Z(n26941) );
  XNOR U26877 ( .A(n26938), .B(n26798), .Z(n26940) );
  IV U26878 ( .A(p_input[388]), .Z(n26798) );
  XOR U26879 ( .A(n26942), .B(n26943), .Z(n26938) );
  AND U26880 ( .A(n26944), .B(n26945), .Z(n26943) );
  XNOR U26881 ( .A(p_input[403]), .B(n26942), .Z(n26945) );
  XNOR U26882 ( .A(n26942), .B(n26807), .Z(n26944) );
  IV U26883 ( .A(p_input[387]), .Z(n26807) );
  XOR U26884 ( .A(n26946), .B(n26947), .Z(n26942) );
  AND U26885 ( .A(n26948), .B(n26949), .Z(n26947) );
  XNOR U26886 ( .A(p_input[402]), .B(n26946), .Z(n26949) );
  XNOR U26887 ( .A(n26946), .B(n26816), .Z(n26948) );
  IV U26888 ( .A(p_input[386]), .Z(n26816) );
  XNOR U26889 ( .A(n26950), .B(n26951), .Z(n26946) );
  AND U26890 ( .A(n26952), .B(n26953), .Z(n26951) );
  XOR U26891 ( .A(p_input[401]), .B(n26950), .Z(n26953) );
  XNOR U26892 ( .A(p_input[385]), .B(n26950), .Z(n26952) );
  AND U26893 ( .A(p_input[400]), .B(n26954), .Z(n26950) );
  IV U26894 ( .A(p_input[384]), .Z(n26954) );
  XOR U26895 ( .A(n26955), .B(n26956), .Z(n26070) );
  AND U26896 ( .A(n833), .B(n26957), .Z(n26956) );
  XNOR U26897 ( .A(n26958), .B(n26955), .Z(n26957) );
  XOR U26898 ( .A(n26959), .B(n26960), .Z(n833) );
  AND U26899 ( .A(n26961), .B(n26962), .Z(n26960) );
  XNOR U26900 ( .A(n26082), .B(n26959), .Z(n26962) );
  AND U26901 ( .A(n26963), .B(n26964), .Z(n26082) );
  XOR U26902 ( .A(n26959), .B(n26081), .Z(n26961) );
  AND U26903 ( .A(n26965), .B(n26966), .Z(n26081) );
  XOR U26904 ( .A(n26967), .B(n26968), .Z(n26959) );
  AND U26905 ( .A(n26969), .B(n26970), .Z(n26968) );
  XOR U26906 ( .A(n26967), .B(n26094), .Z(n26970) );
  XOR U26907 ( .A(n26971), .B(n26972), .Z(n26094) );
  AND U26908 ( .A(n575), .B(n26973), .Z(n26972) );
  XOR U26909 ( .A(n26974), .B(n26971), .Z(n26973) );
  XNOR U26910 ( .A(n26091), .B(n26967), .Z(n26969) );
  XOR U26911 ( .A(n26975), .B(n26976), .Z(n26091) );
  AND U26912 ( .A(n572), .B(n26977), .Z(n26976) );
  XOR U26913 ( .A(n26978), .B(n26975), .Z(n26977) );
  XOR U26914 ( .A(n26979), .B(n26980), .Z(n26967) );
  AND U26915 ( .A(n26981), .B(n26982), .Z(n26980) );
  XOR U26916 ( .A(n26979), .B(n26106), .Z(n26982) );
  XOR U26917 ( .A(n26983), .B(n26984), .Z(n26106) );
  AND U26918 ( .A(n575), .B(n26985), .Z(n26984) );
  XOR U26919 ( .A(n26986), .B(n26983), .Z(n26985) );
  XNOR U26920 ( .A(n26103), .B(n26979), .Z(n26981) );
  XOR U26921 ( .A(n26987), .B(n26988), .Z(n26103) );
  AND U26922 ( .A(n572), .B(n26989), .Z(n26988) );
  XOR U26923 ( .A(n26990), .B(n26987), .Z(n26989) );
  XOR U26924 ( .A(n26991), .B(n26992), .Z(n26979) );
  AND U26925 ( .A(n26993), .B(n26994), .Z(n26992) );
  XOR U26926 ( .A(n26991), .B(n26118), .Z(n26994) );
  XOR U26927 ( .A(n26995), .B(n26996), .Z(n26118) );
  AND U26928 ( .A(n575), .B(n26997), .Z(n26996) );
  XOR U26929 ( .A(n26998), .B(n26995), .Z(n26997) );
  XNOR U26930 ( .A(n26115), .B(n26991), .Z(n26993) );
  XOR U26931 ( .A(n26999), .B(n27000), .Z(n26115) );
  AND U26932 ( .A(n572), .B(n27001), .Z(n27000) );
  XOR U26933 ( .A(n27002), .B(n26999), .Z(n27001) );
  XOR U26934 ( .A(n27003), .B(n27004), .Z(n26991) );
  AND U26935 ( .A(n27005), .B(n27006), .Z(n27004) );
  XOR U26936 ( .A(n27003), .B(n26130), .Z(n27006) );
  XOR U26937 ( .A(n27007), .B(n27008), .Z(n26130) );
  AND U26938 ( .A(n575), .B(n27009), .Z(n27008) );
  XOR U26939 ( .A(n27010), .B(n27007), .Z(n27009) );
  XNOR U26940 ( .A(n26127), .B(n27003), .Z(n27005) );
  XOR U26941 ( .A(n27011), .B(n27012), .Z(n26127) );
  AND U26942 ( .A(n572), .B(n27013), .Z(n27012) );
  XOR U26943 ( .A(n27014), .B(n27011), .Z(n27013) );
  XOR U26944 ( .A(n27015), .B(n27016), .Z(n27003) );
  AND U26945 ( .A(n27017), .B(n27018), .Z(n27016) );
  XOR U26946 ( .A(n27015), .B(n26142), .Z(n27018) );
  XOR U26947 ( .A(n27019), .B(n27020), .Z(n26142) );
  AND U26948 ( .A(n575), .B(n27021), .Z(n27020) );
  XOR U26949 ( .A(n27022), .B(n27019), .Z(n27021) );
  XNOR U26950 ( .A(n26139), .B(n27015), .Z(n27017) );
  XOR U26951 ( .A(n27023), .B(n27024), .Z(n26139) );
  AND U26952 ( .A(n572), .B(n27025), .Z(n27024) );
  XOR U26953 ( .A(n27026), .B(n27023), .Z(n27025) );
  XOR U26954 ( .A(n27027), .B(n27028), .Z(n27015) );
  AND U26955 ( .A(n27029), .B(n27030), .Z(n27028) );
  XOR U26956 ( .A(n27027), .B(n26154), .Z(n27030) );
  XOR U26957 ( .A(n27031), .B(n27032), .Z(n26154) );
  AND U26958 ( .A(n575), .B(n27033), .Z(n27032) );
  XOR U26959 ( .A(n27034), .B(n27031), .Z(n27033) );
  XNOR U26960 ( .A(n26151), .B(n27027), .Z(n27029) );
  XOR U26961 ( .A(n27035), .B(n27036), .Z(n26151) );
  AND U26962 ( .A(n572), .B(n27037), .Z(n27036) );
  XOR U26963 ( .A(n27038), .B(n27035), .Z(n27037) );
  XOR U26964 ( .A(n27039), .B(n27040), .Z(n27027) );
  AND U26965 ( .A(n27041), .B(n27042), .Z(n27040) );
  XOR U26966 ( .A(n27039), .B(n26166), .Z(n27042) );
  XOR U26967 ( .A(n27043), .B(n27044), .Z(n26166) );
  AND U26968 ( .A(n575), .B(n27045), .Z(n27044) );
  XOR U26969 ( .A(n27046), .B(n27043), .Z(n27045) );
  XNOR U26970 ( .A(n26163), .B(n27039), .Z(n27041) );
  XOR U26971 ( .A(n27047), .B(n27048), .Z(n26163) );
  AND U26972 ( .A(n572), .B(n27049), .Z(n27048) );
  XOR U26973 ( .A(n27050), .B(n27047), .Z(n27049) );
  XOR U26974 ( .A(n27051), .B(n27052), .Z(n27039) );
  AND U26975 ( .A(n27053), .B(n27054), .Z(n27052) );
  XOR U26976 ( .A(n27051), .B(n26178), .Z(n27054) );
  XOR U26977 ( .A(n27055), .B(n27056), .Z(n26178) );
  AND U26978 ( .A(n575), .B(n27057), .Z(n27056) );
  XOR U26979 ( .A(n27058), .B(n27055), .Z(n27057) );
  XNOR U26980 ( .A(n26175), .B(n27051), .Z(n27053) );
  XOR U26981 ( .A(n27059), .B(n27060), .Z(n26175) );
  AND U26982 ( .A(n572), .B(n27061), .Z(n27060) );
  XOR U26983 ( .A(n27062), .B(n27059), .Z(n27061) );
  XOR U26984 ( .A(n27063), .B(n27064), .Z(n27051) );
  AND U26985 ( .A(n27065), .B(n27066), .Z(n27064) );
  XOR U26986 ( .A(n27063), .B(n26190), .Z(n27066) );
  XOR U26987 ( .A(n27067), .B(n27068), .Z(n26190) );
  AND U26988 ( .A(n575), .B(n27069), .Z(n27068) );
  XOR U26989 ( .A(n27070), .B(n27067), .Z(n27069) );
  XNOR U26990 ( .A(n26187), .B(n27063), .Z(n27065) );
  XOR U26991 ( .A(n27071), .B(n27072), .Z(n26187) );
  AND U26992 ( .A(n572), .B(n27073), .Z(n27072) );
  XOR U26993 ( .A(n27074), .B(n27071), .Z(n27073) );
  XOR U26994 ( .A(n27075), .B(n27076), .Z(n27063) );
  AND U26995 ( .A(n27077), .B(n27078), .Z(n27076) );
  XOR U26996 ( .A(n27075), .B(n26202), .Z(n27078) );
  XOR U26997 ( .A(n27079), .B(n27080), .Z(n26202) );
  AND U26998 ( .A(n575), .B(n27081), .Z(n27080) );
  XOR U26999 ( .A(n27082), .B(n27079), .Z(n27081) );
  XNOR U27000 ( .A(n26199), .B(n27075), .Z(n27077) );
  XOR U27001 ( .A(n27083), .B(n27084), .Z(n26199) );
  AND U27002 ( .A(n572), .B(n27085), .Z(n27084) );
  XOR U27003 ( .A(n27086), .B(n27083), .Z(n27085) );
  XOR U27004 ( .A(n27087), .B(n27088), .Z(n27075) );
  AND U27005 ( .A(n27089), .B(n27090), .Z(n27088) );
  XOR U27006 ( .A(n27087), .B(n26214), .Z(n27090) );
  XOR U27007 ( .A(n27091), .B(n27092), .Z(n26214) );
  AND U27008 ( .A(n575), .B(n27093), .Z(n27092) );
  XOR U27009 ( .A(n27094), .B(n27091), .Z(n27093) );
  XNOR U27010 ( .A(n26211), .B(n27087), .Z(n27089) );
  XOR U27011 ( .A(n27095), .B(n27096), .Z(n26211) );
  AND U27012 ( .A(n572), .B(n27097), .Z(n27096) );
  XOR U27013 ( .A(n27098), .B(n27095), .Z(n27097) );
  XOR U27014 ( .A(n27099), .B(n27100), .Z(n27087) );
  AND U27015 ( .A(n27101), .B(n27102), .Z(n27100) );
  XOR U27016 ( .A(n27099), .B(n26226), .Z(n27102) );
  XOR U27017 ( .A(n27103), .B(n27104), .Z(n26226) );
  AND U27018 ( .A(n575), .B(n27105), .Z(n27104) );
  XOR U27019 ( .A(n27106), .B(n27103), .Z(n27105) );
  XNOR U27020 ( .A(n26223), .B(n27099), .Z(n27101) );
  XOR U27021 ( .A(n27107), .B(n27108), .Z(n26223) );
  AND U27022 ( .A(n572), .B(n27109), .Z(n27108) );
  XOR U27023 ( .A(n27110), .B(n27107), .Z(n27109) );
  XOR U27024 ( .A(n27111), .B(n27112), .Z(n27099) );
  AND U27025 ( .A(n27113), .B(n27114), .Z(n27112) );
  XOR U27026 ( .A(n27111), .B(n26238), .Z(n27114) );
  XOR U27027 ( .A(n27115), .B(n27116), .Z(n26238) );
  AND U27028 ( .A(n575), .B(n27117), .Z(n27116) );
  XOR U27029 ( .A(n27118), .B(n27115), .Z(n27117) );
  XNOR U27030 ( .A(n26235), .B(n27111), .Z(n27113) );
  XOR U27031 ( .A(n27119), .B(n27120), .Z(n26235) );
  AND U27032 ( .A(n572), .B(n27121), .Z(n27120) );
  XOR U27033 ( .A(n27122), .B(n27119), .Z(n27121) );
  XOR U27034 ( .A(n27123), .B(n27124), .Z(n27111) );
  AND U27035 ( .A(n27125), .B(n27126), .Z(n27124) );
  XNOR U27036 ( .A(n27127), .B(n26251), .Z(n27126) );
  XOR U27037 ( .A(n27128), .B(n27129), .Z(n26251) );
  AND U27038 ( .A(n575), .B(n27130), .Z(n27129) );
  XOR U27039 ( .A(n27128), .B(n27131), .Z(n27130) );
  XNOR U27040 ( .A(n26248), .B(n27123), .Z(n27125) );
  XOR U27041 ( .A(n27132), .B(n27133), .Z(n26248) );
  AND U27042 ( .A(n572), .B(n27134), .Z(n27133) );
  XOR U27043 ( .A(n27132), .B(n27135), .Z(n27134) );
  IV U27044 ( .A(n27127), .Z(n27123) );
  AND U27045 ( .A(n26955), .B(n26958), .Z(n27127) );
  XNOR U27046 ( .A(n27136), .B(n27137), .Z(n26958) );
  AND U27047 ( .A(n575), .B(n27138), .Z(n27137) );
  XNOR U27048 ( .A(n27139), .B(n27136), .Z(n27138) );
  XOR U27049 ( .A(n27140), .B(n27141), .Z(n575) );
  AND U27050 ( .A(n27142), .B(n27143), .Z(n27141) );
  XNOR U27051 ( .A(n26963), .B(n27140), .Z(n27143) );
  AND U27052 ( .A(p_input[383]), .B(p_input[367]), .Z(n26963) );
  XOR U27053 ( .A(n27140), .B(n26964), .Z(n27142) );
  AND U27054 ( .A(p_input[351]), .B(p_input[335]), .Z(n26964) );
  XOR U27055 ( .A(n27144), .B(n27145), .Z(n27140) );
  AND U27056 ( .A(n27146), .B(n27147), .Z(n27145) );
  XOR U27057 ( .A(n27144), .B(n26974), .Z(n27147) );
  XNOR U27058 ( .A(p_input[366]), .B(n27148), .Z(n26974) );
  AND U27059 ( .A(n991), .B(n27149), .Z(n27148) );
  XOR U27060 ( .A(p_input[382]), .B(p_input[366]), .Z(n27149) );
  XNOR U27061 ( .A(n26971), .B(n27144), .Z(n27146) );
  XOR U27062 ( .A(n27150), .B(n27151), .Z(n26971) );
  AND U27063 ( .A(n989), .B(n27152), .Z(n27151) );
  XOR U27064 ( .A(p_input[350]), .B(p_input[334]), .Z(n27152) );
  XOR U27065 ( .A(n27153), .B(n27154), .Z(n27144) );
  AND U27066 ( .A(n27155), .B(n27156), .Z(n27154) );
  XOR U27067 ( .A(n27153), .B(n26986), .Z(n27156) );
  XNOR U27068 ( .A(p_input[365]), .B(n27157), .Z(n26986) );
  AND U27069 ( .A(n991), .B(n27158), .Z(n27157) );
  XOR U27070 ( .A(p_input[381]), .B(p_input[365]), .Z(n27158) );
  XNOR U27071 ( .A(n26983), .B(n27153), .Z(n27155) );
  XOR U27072 ( .A(n27159), .B(n27160), .Z(n26983) );
  AND U27073 ( .A(n989), .B(n27161), .Z(n27160) );
  XOR U27074 ( .A(p_input[349]), .B(p_input[333]), .Z(n27161) );
  XOR U27075 ( .A(n27162), .B(n27163), .Z(n27153) );
  AND U27076 ( .A(n27164), .B(n27165), .Z(n27163) );
  XOR U27077 ( .A(n27162), .B(n26998), .Z(n27165) );
  XNOR U27078 ( .A(p_input[364]), .B(n27166), .Z(n26998) );
  AND U27079 ( .A(n991), .B(n27167), .Z(n27166) );
  XOR U27080 ( .A(p_input[380]), .B(p_input[364]), .Z(n27167) );
  XNOR U27081 ( .A(n26995), .B(n27162), .Z(n27164) );
  XOR U27082 ( .A(n27168), .B(n27169), .Z(n26995) );
  AND U27083 ( .A(n989), .B(n27170), .Z(n27169) );
  XOR U27084 ( .A(p_input[348]), .B(p_input[332]), .Z(n27170) );
  XOR U27085 ( .A(n27171), .B(n27172), .Z(n27162) );
  AND U27086 ( .A(n27173), .B(n27174), .Z(n27172) );
  XOR U27087 ( .A(n27171), .B(n27010), .Z(n27174) );
  XNOR U27088 ( .A(p_input[363]), .B(n27175), .Z(n27010) );
  AND U27089 ( .A(n991), .B(n27176), .Z(n27175) );
  XOR U27090 ( .A(p_input[379]), .B(p_input[363]), .Z(n27176) );
  XNOR U27091 ( .A(n27007), .B(n27171), .Z(n27173) );
  XOR U27092 ( .A(n27177), .B(n27178), .Z(n27007) );
  AND U27093 ( .A(n989), .B(n27179), .Z(n27178) );
  XOR U27094 ( .A(p_input[347]), .B(p_input[331]), .Z(n27179) );
  XOR U27095 ( .A(n27180), .B(n27181), .Z(n27171) );
  AND U27096 ( .A(n27182), .B(n27183), .Z(n27181) );
  XOR U27097 ( .A(n27180), .B(n27022), .Z(n27183) );
  XNOR U27098 ( .A(p_input[362]), .B(n27184), .Z(n27022) );
  AND U27099 ( .A(n991), .B(n27185), .Z(n27184) );
  XOR U27100 ( .A(p_input[378]), .B(p_input[362]), .Z(n27185) );
  XNOR U27101 ( .A(n27019), .B(n27180), .Z(n27182) );
  XOR U27102 ( .A(n27186), .B(n27187), .Z(n27019) );
  AND U27103 ( .A(n989), .B(n27188), .Z(n27187) );
  XOR U27104 ( .A(p_input[346]), .B(p_input[330]), .Z(n27188) );
  XOR U27105 ( .A(n27189), .B(n27190), .Z(n27180) );
  AND U27106 ( .A(n27191), .B(n27192), .Z(n27190) );
  XOR U27107 ( .A(n27189), .B(n27034), .Z(n27192) );
  XNOR U27108 ( .A(p_input[361]), .B(n27193), .Z(n27034) );
  AND U27109 ( .A(n991), .B(n27194), .Z(n27193) );
  XOR U27110 ( .A(p_input[377]), .B(p_input[361]), .Z(n27194) );
  XNOR U27111 ( .A(n27031), .B(n27189), .Z(n27191) );
  XOR U27112 ( .A(n27195), .B(n27196), .Z(n27031) );
  AND U27113 ( .A(n989), .B(n27197), .Z(n27196) );
  XOR U27114 ( .A(p_input[345]), .B(p_input[329]), .Z(n27197) );
  XOR U27115 ( .A(n27198), .B(n27199), .Z(n27189) );
  AND U27116 ( .A(n27200), .B(n27201), .Z(n27199) );
  XOR U27117 ( .A(n27198), .B(n27046), .Z(n27201) );
  XNOR U27118 ( .A(p_input[360]), .B(n27202), .Z(n27046) );
  AND U27119 ( .A(n991), .B(n27203), .Z(n27202) );
  XOR U27120 ( .A(p_input[376]), .B(p_input[360]), .Z(n27203) );
  XNOR U27121 ( .A(n27043), .B(n27198), .Z(n27200) );
  XOR U27122 ( .A(n27204), .B(n27205), .Z(n27043) );
  AND U27123 ( .A(n989), .B(n27206), .Z(n27205) );
  XOR U27124 ( .A(p_input[344]), .B(p_input[328]), .Z(n27206) );
  XOR U27125 ( .A(n27207), .B(n27208), .Z(n27198) );
  AND U27126 ( .A(n27209), .B(n27210), .Z(n27208) );
  XOR U27127 ( .A(n27207), .B(n27058), .Z(n27210) );
  XNOR U27128 ( .A(p_input[359]), .B(n27211), .Z(n27058) );
  AND U27129 ( .A(n991), .B(n27212), .Z(n27211) );
  XOR U27130 ( .A(p_input[375]), .B(p_input[359]), .Z(n27212) );
  XNOR U27131 ( .A(n27055), .B(n27207), .Z(n27209) );
  XOR U27132 ( .A(n27213), .B(n27214), .Z(n27055) );
  AND U27133 ( .A(n989), .B(n27215), .Z(n27214) );
  XOR U27134 ( .A(p_input[343]), .B(p_input[327]), .Z(n27215) );
  XOR U27135 ( .A(n27216), .B(n27217), .Z(n27207) );
  AND U27136 ( .A(n27218), .B(n27219), .Z(n27217) );
  XOR U27137 ( .A(n27216), .B(n27070), .Z(n27219) );
  XNOR U27138 ( .A(p_input[358]), .B(n27220), .Z(n27070) );
  AND U27139 ( .A(n991), .B(n27221), .Z(n27220) );
  XOR U27140 ( .A(p_input[374]), .B(p_input[358]), .Z(n27221) );
  XNOR U27141 ( .A(n27067), .B(n27216), .Z(n27218) );
  XOR U27142 ( .A(n27222), .B(n27223), .Z(n27067) );
  AND U27143 ( .A(n989), .B(n27224), .Z(n27223) );
  XOR U27144 ( .A(p_input[342]), .B(p_input[326]), .Z(n27224) );
  XOR U27145 ( .A(n27225), .B(n27226), .Z(n27216) );
  AND U27146 ( .A(n27227), .B(n27228), .Z(n27226) );
  XOR U27147 ( .A(n27225), .B(n27082), .Z(n27228) );
  XNOR U27148 ( .A(p_input[357]), .B(n27229), .Z(n27082) );
  AND U27149 ( .A(n991), .B(n27230), .Z(n27229) );
  XOR U27150 ( .A(p_input[373]), .B(p_input[357]), .Z(n27230) );
  XNOR U27151 ( .A(n27079), .B(n27225), .Z(n27227) );
  XOR U27152 ( .A(n27231), .B(n27232), .Z(n27079) );
  AND U27153 ( .A(n989), .B(n27233), .Z(n27232) );
  XOR U27154 ( .A(p_input[341]), .B(p_input[325]), .Z(n27233) );
  XOR U27155 ( .A(n27234), .B(n27235), .Z(n27225) );
  AND U27156 ( .A(n27236), .B(n27237), .Z(n27235) );
  XOR U27157 ( .A(n27234), .B(n27094), .Z(n27237) );
  XNOR U27158 ( .A(p_input[356]), .B(n27238), .Z(n27094) );
  AND U27159 ( .A(n991), .B(n27239), .Z(n27238) );
  XOR U27160 ( .A(p_input[372]), .B(p_input[356]), .Z(n27239) );
  XNOR U27161 ( .A(n27091), .B(n27234), .Z(n27236) );
  XOR U27162 ( .A(n27240), .B(n27241), .Z(n27091) );
  AND U27163 ( .A(n989), .B(n27242), .Z(n27241) );
  XOR U27164 ( .A(p_input[340]), .B(p_input[324]), .Z(n27242) );
  XOR U27165 ( .A(n27243), .B(n27244), .Z(n27234) );
  AND U27166 ( .A(n27245), .B(n27246), .Z(n27244) );
  XOR U27167 ( .A(n27243), .B(n27106), .Z(n27246) );
  XNOR U27168 ( .A(p_input[355]), .B(n27247), .Z(n27106) );
  AND U27169 ( .A(n991), .B(n27248), .Z(n27247) );
  XOR U27170 ( .A(p_input[371]), .B(p_input[355]), .Z(n27248) );
  XNOR U27171 ( .A(n27103), .B(n27243), .Z(n27245) );
  XOR U27172 ( .A(n27249), .B(n27250), .Z(n27103) );
  AND U27173 ( .A(n989), .B(n27251), .Z(n27250) );
  XOR U27174 ( .A(p_input[339]), .B(p_input[323]), .Z(n27251) );
  XOR U27175 ( .A(n27252), .B(n27253), .Z(n27243) );
  AND U27176 ( .A(n27254), .B(n27255), .Z(n27253) );
  XOR U27177 ( .A(n27252), .B(n27118), .Z(n27255) );
  XNOR U27178 ( .A(p_input[354]), .B(n27256), .Z(n27118) );
  AND U27179 ( .A(n991), .B(n27257), .Z(n27256) );
  XOR U27180 ( .A(p_input[370]), .B(p_input[354]), .Z(n27257) );
  XNOR U27181 ( .A(n27115), .B(n27252), .Z(n27254) );
  XOR U27182 ( .A(n27258), .B(n27259), .Z(n27115) );
  AND U27183 ( .A(n989), .B(n27260), .Z(n27259) );
  XOR U27184 ( .A(p_input[338]), .B(p_input[322]), .Z(n27260) );
  XOR U27185 ( .A(n27261), .B(n27262), .Z(n27252) );
  AND U27186 ( .A(n27263), .B(n27264), .Z(n27262) );
  XNOR U27187 ( .A(n27265), .B(n27131), .Z(n27264) );
  XNOR U27188 ( .A(p_input[353]), .B(n27266), .Z(n27131) );
  AND U27189 ( .A(n991), .B(n27267), .Z(n27266) );
  XNOR U27190 ( .A(p_input[369]), .B(n27268), .Z(n27267) );
  IV U27191 ( .A(p_input[353]), .Z(n27268) );
  XNOR U27192 ( .A(n27128), .B(n27261), .Z(n27263) );
  XNOR U27193 ( .A(p_input[321]), .B(n27269), .Z(n27128) );
  AND U27194 ( .A(n989), .B(n27270), .Z(n27269) );
  XOR U27195 ( .A(p_input[337]), .B(p_input[321]), .Z(n27270) );
  IV U27196 ( .A(n27265), .Z(n27261) );
  AND U27197 ( .A(n27136), .B(n27139), .Z(n27265) );
  XOR U27198 ( .A(p_input[352]), .B(n27271), .Z(n27139) );
  AND U27199 ( .A(n991), .B(n27272), .Z(n27271) );
  XOR U27200 ( .A(p_input[368]), .B(p_input[352]), .Z(n27272) );
  XOR U27201 ( .A(n27273), .B(n27274), .Z(n991) );
  AND U27202 ( .A(n27275), .B(n27276), .Z(n27274) );
  XNOR U27203 ( .A(p_input[383]), .B(n27273), .Z(n27276) );
  XOR U27204 ( .A(n27273), .B(p_input[367]), .Z(n27275) );
  XOR U27205 ( .A(n27277), .B(n27278), .Z(n27273) );
  AND U27206 ( .A(n27279), .B(n27280), .Z(n27278) );
  XNOR U27207 ( .A(p_input[382]), .B(n27277), .Z(n27280) );
  XOR U27208 ( .A(n27277), .B(p_input[366]), .Z(n27279) );
  XOR U27209 ( .A(n27281), .B(n27282), .Z(n27277) );
  AND U27210 ( .A(n27283), .B(n27284), .Z(n27282) );
  XNOR U27211 ( .A(p_input[381]), .B(n27281), .Z(n27284) );
  XOR U27212 ( .A(n27281), .B(p_input[365]), .Z(n27283) );
  XOR U27213 ( .A(n27285), .B(n27286), .Z(n27281) );
  AND U27214 ( .A(n27287), .B(n27288), .Z(n27286) );
  XNOR U27215 ( .A(p_input[380]), .B(n27285), .Z(n27288) );
  XOR U27216 ( .A(n27285), .B(p_input[364]), .Z(n27287) );
  XOR U27217 ( .A(n27289), .B(n27290), .Z(n27285) );
  AND U27218 ( .A(n27291), .B(n27292), .Z(n27290) );
  XNOR U27219 ( .A(p_input[379]), .B(n27289), .Z(n27292) );
  XOR U27220 ( .A(n27289), .B(p_input[363]), .Z(n27291) );
  XOR U27221 ( .A(n27293), .B(n27294), .Z(n27289) );
  AND U27222 ( .A(n27295), .B(n27296), .Z(n27294) );
  XNOR U27223 ( .A(p_input[378]), .B(n27293), .Z(n27296) );
  XOR U27224 ( .A(n27293), .B(p_input[362]), .Z(n27295) );
  XOR U27225 ( .A(n27297), .B(n27298), .Z(n27293) );
  AND U27226 ( .A(n27299), .B(n27300), .Z(n27298) );
  XNOR U27227 ( .A(p_input[377]), .B(n27297), .Z(n27300) );
  XOR U27228 ( .A(n27297), .B(p_input[361]), .Z(n27299) );
  XOR U27229 ( .A(n27301), .B(n27302), .Z(n27297) );
  AND U27230 ( .A(n27303), .B(n27304), .Z(n27302) );
  XNOR U27231 ( .A(p_input[376]), .B(n27301), .Z(n27304) );
  XOR U27232 ( .A(n27301), .B(p_input[360]), .Z(n27303) );
  XOR U27233 ( .A(n27305), .B(n27306), .Z(n27301) );
  AND U27234 ( .A(n27307), .B(n27308), .Z(n27306) );
  XNOR U27235 ( .A(p_input[375]), .B(n27305), .Z(n27308) );
  XOR U27236 ( .A(n27305), .B(p_input[359]), .Z(n27307) );
  XOR U27237 ( .A(n27309), .B(n27310), .Z(n27305) );
  AND U27238 ( .A(n27311), .B(n27312), .Z(n27310) );
  XNOR U27239 ( .A(p_input[374]), .B(n27309), .Z(n27312) );
  XOR U27240 ( .A(n27309), .B(p_input[358]), .Z(n27311) );
  XOR U27241 ( .A(n27313), .B(n27314), .Z(n27309) );
  AND U27242 ( .A(n27315), .B(n27316), .Z(n27314) );
  XNOR U27243 ( .A(p_input[373]), .B(n27313), .Z(n27316) );
  XOR U27244 ( .A(n27313), .B(p_input[357]), .Z(n27315) );
  XOR U27245 ( .A(n27317), .B(n27318), .Z(n27313) );
  AND U27246 ( .A(n27319), .B(n27320), .Z(n27318) );
  XNOR U27247 ( .A(p_input[372]), .B(n27317), .Z(n27320) );
  XOR U27248 ( .A(n27317), .B(p_input[356]), .Z(n27319) );
  XOR U27249 ( .A(n27321), .B(n27322), .Z(n27317) );
  AND U27250 ( .A(n27323), .B(n27324), .Z(n27322) );
  XNOR U27251 ( .A(p_input[371]), .B(n27321), .Z(n27324) );
  XOR U27252 ( .A(n27321), .B(p_input[355]), .Z(n27323) );
  XOR U27253 ( .A(n27325), .B(n27326), .Z(n27321) );
  AND U27254 ( .A(n27327), .B(n27328), .Z(n27326) );
  XNOR U27255 ( .A(p_input[370]), .B(n27325), .Z(n27328) );
  XOR U27256 ( .A(n27325), .B(p_input[354]), .Z(n27327) );
  XNOR U27257 ( .A(n27329), .B(n27330), .Z(n27325) );
  AND U27258 ( .A(n27331), .B(n27332), .Z(n27330) );
  XOR U27259 ( .A(p_input[369]), .B(n27329), .Z(n27332) );
  XNOR U27260 ( .A(p_input[353]), .B(n27329), .Z(n27331) );
  AND U27261 ( .A(p_input[368]), .B(n27333), .Z(n27329) );
  IV U27262 ( .A(p_input[352]), .Z(n27333) );
  XNOR U27263 ( .A(p_input[320]), .B(n27334), .Z(n27136) );
  AND U27264 ( .A(n989), .B(n27335), .Z(n27334) );
  XOR U27265 ( .A(p_input[336]), .B(p_input[320]), .Z(n27335) );
  XOR U27266 ( .A(n27336), .B(n27337), .Z(n989) );
  AND U27267 ( .A(n27338), .B(n27339), .Z(n27337) );
  XNOR U27268 ( .A(p_input[351]), .B(n27336), .Z(n27339) );
  XOR U27269 ( .A(n27336), .B(p_input[335]), .Z(n27338) );
  XOR U27270 ( .A(n27340), .B(n27341), .Z(n27336) );
  AND U27271 ( .A(n27342), .B(n27343), .Z(n27341) );
  XNOR U27272 ( .A(p_input[350]), .B(n27340), .Z(n27343) );
  XNOR U27273 ( .A(n27340), .B(n27150), .Z(n27342) );
  IV U27274 ( .A(p_input[334]), .Z(n27150) );
  XOR U27275 ( .A(n27344), .B(n27345), .Z(n27340) );
  AND U27276 ( .A(n27346), .B(n27347), .Z(n27345) );
  XNOR U27277 ( .A(p_input[349]), .B(n27344), .Z(n27347) );
  XNOR U27278 ( .A(n27344), .B(n27159), .Z(n27346) );
  IV U27279 ( .A(p_input[333]), .Z(n27159) );
  XOR U27280 ( .A(n27348), .B(n27349), .Z(n27344) );
  AND U27281 ( .A(n27350), .B(n27351), .Z(n27349) );
  XNOR U27282 ( .A(p_input[348]), .B(n27348), .Z(n27351) );
  XNOR U27283 ( .A(n27348), .B(n27168), .Z(n27350) );
  IV U27284 ( .A(p_input[332]), .Z(n27168) );
  XOR U27285 ( .A(n27352), .B(n27353), .Z(n27348) );
  AND U27286 ( .A(n27354), .B(n27355), .Z(n27353) );
  XNOR U27287 ( .A(p_input[347]), .B(n27352), .Z(n27355) );
  XNOR U27288 ( .A(n27352), .B(n27177), .Z(n27354) );
  IV U27289 ( .A(p_input[331]), .Z(n27177) );
  XOR U27290 ( .A(n27356), .B(n27357), .Z(n27352) );
  AND U27291 ( .A(n27358), .B(n27359), .Z(n27357) );
  XNOR U27292 ( .A(p_input[346]), .B(n27356), .Z(n27359) );
  XNOR U27293 ( .A(n27356), .B(n27186), .Z(n27358) );
  IV U27294 ( .A(p_input[330]), .Z(n27186) );
  XOR U27295 ( .A(n27360), .B(n27361), .Z(n27356) );
  AND U27296 ( .A(n27362), .B(n27363), .Z(n27361) );
  XNOR U27297 ( .A(p_input[345]), .B(n27360), .Z(n27363) );
  XNOR U27298 ( .A(n27360), .B(n27195), .Z(n27362) );
  IV U27299 ( .A(p_input[329]), .Z(n27195) );
  XOR U27300 ( .A(n27364), .B(n27365), .Z(n27360) );
  AND U27301 ( .A(n27366), .B(n27367), .Z(n27365) );
  XNOR U27302 ( .A(p_input[344]), .B(n27364), .Z(n27367) );
  XNOR U27303 ( .A(n27364), .B(n27204), .Z(n27366) );
  IV U27304 ( .A(p_input[328]), .Z(n27204) );
  XOR U27305 ( .A(n27368), .B(n27369), .Z(n27364) );
  AND U27306 ( .A(n27370), .B(n27371), .Z(n27369) );
  XNOR U27307 ( .A(p_input[343]), .B(n27368), .Z(n27371) );
  XNOR U27308 ( .A(n27368), .B(n27213), .Z(n27370) );
  IV U27309 ( .A(p_input[327]), .Z(n27213) );
  XOR U27310 ( .A(n27372), .B(n27373), .Z(n27368) );
  AND U27311 ( .A(n27374), .B(n27375), .Z(n27373) );
  XNOR U27312 ( .A(p_input[342]), .B(n27372), .Z(n27375) );
  XNOR U27313 ( .A(n27372), .B(n27222), .Z(n27374) );
  IV U27314 ( .A(p_input[326]), .Z(n27222) );
  XOR U27315 ( .A(n27376), .B(n27377), .Z(n27372) );
  AND U27316 ( .A(n27378), .B(n27379), .Z(n27377) );
  XNOR U27317 ( .A(p_input[341]), .B(n27376), .Z(n27379) );
  XNOR U27318 ( .A(n27376), .B(n27231), .Z(n27378) );
  IV U27319 ( .A(p_input[325]), .Z(n27231) );
  XOR U27320 ( .A(n27380), .B(n27381), .Z(n27376) );
  AND U27321 ( .A(n27382), .B(n27383), .Z(n27381) );
  XNOR U27322 ( .A(p_input[340]), .B(n27380), .Z(n27383) );
  XNOR U27323 ( .A(n27380), .B(n27240), .Z(n27382) );
  IV U27324 ( .A(p_input[324]), .Z(n27240) );
  XOR U27325 ( .A(n27384), .B(n27385), .Z(n27380) );
  AND U27326 ( .A(n27386), .B(n27387), .Z(n27385) );
  XNOR U27327 ( .A(p_input[339]), .B(n27384), .Z(n27387) );
  XNOR U27328 ( .A(n27384), .B(n27249), .Z(n27386) );
  IV U27329 ( .A(p_input[323]), .Z(n27249) );
  XOR U27330 ( .A(n27388), .B(n27389), .Z(n27384) );
  AND U27331 ( .A(n27390), .B(n27391), .Z(n27389) );
  XNOR U27332 ( .A(p_input[338]), .B(n27388), .Z(n27391) );
  XNOR U27333 ( .A(n27388), .B(n27258), .Z(n27390) );
  IV U27334 ( .A(p_input[322]), .Z(n27258) );
  XNOR U27335 ( .A(n27392), .B(n27393), .Z(n27388) );
  AND U27336 ( .A(n27394), .B(n27395), .Z(n27393) );
  XOR U27337 ( .A(p_input[337]), .B(n27392), .Z(n27395) );
  XNOR U27338 ( .A(p_input[321]), .B(n27392), .Z(n27394) );
  AND U27339 ( .A(p_input[336]), .B(n27396), .Z(n27392) );
  IV U27340 ( .A(p_input[320]), .Z(n27396) );
  XOR U27341 ( .A(n27397), .B(n27398), .Z(n26955) );
  AND U27342 ( .A(n572), .B(n27399), .Z(n27398) );
  XNOR U27343 ( .A(n27400), .B(n27397), .Z(n27399) );
  XOR U27344 ( .A(n27401), .B(n27402), .Z(n572) );
  AND U27345 ( .A(n27403), .B(n27404), .Z(n27402) );
  XNOR U27346 ( .A(n26966), .B(n27401), .Z(n27404) );
  AND U27347 ( .A(p_input[319]), .B(p_input[303]), .Z(n26966) );
  XOR U27348 ( .A(n27401), .B(n26965), .Z(n27403) );
  AND U27349 ( .A(p_input[271]), .B(p_input[287]), .Z(n26965) );
  XOR U27350 ( .A(n27405), .B(n27406), .Z(n27401) );
  AND U27351 ( .A(n27407), .B(n27408), .Z(n27406) );
  XOR U27352 ( .A(n27405), .B(n26978), .Z(n27408) );
  XNOR U27353 ( .A(p_input[302]), .B(n27409), .Z(n26978) );
  AND U27354 ( .A(n995), .B(n27410), .Z(n27409) );
  XOR U27355 ( .A(p_input[318]), .B(p_input[302]), .Z(n27410) );
  XNOR U27356 ( .A(n26975), .B(n27405), .Z(n27407) );
  XOR U27357 ( .A(n27411), .B(n27412), .Z(n26975) );
  AND U27358 ( .A(n992), .B(n27413), .Z(n27412) );
  XOR U27359 ( .A(p_input[286]), .B(p_input[270]), .Z(n27413) );
  XOR U27360 ( .A(n27414), .B(n27415), .Z(n27405) );
  AND U27361 ( .A(n27416), .B(n27417), .Z(n27415) );
  XOR U27362 ( .A(n27414), .B(n26990), .Z(n27417) );
  XNOR U27363 ( .A(p_input[301]), .B(n27418), .Z(n26990) );
  AND U27364 ( .A(n995), .B(n27419), .Z(n27418) );
  XOR U27365 ( .A(p_input[317]), .B(p_input[301]), .Z(n27419) );
  XNOR U27366 ( .A(n26987), .B(n27414), .Z(n27416) );
  XOR U27367 ( .A(n27420), .B(n27421), .Z(n26987) );
  AND U27368 ( .A(n992), .B(n27422), .Z(n27421) );
  XOR U27369 ( .A(p_input[285]), .B(p_input[269]), .Z(n27422) );
  XOR U27370 ( .A(n27423), .B(n27424), .Z(n27414) );
  AND U27371 ( .A(n27425), .B(n27426), .Z(n27424) );
  XOR U27372 ( .A(n27423), .B(n27002), .Z(n27426) );
  XNOR U27373 ( .A(p_input[300]), .B(n27427), .Z(n27002) );
  AND U27374 ( .A(n995), .B(n27428), .Z(n27427) );
  XOR U27375 ( .A(p_input[316]), .B(p_input[300]), .Z(n27428) );
  XNOR U27376 ( .A(n26999), .B(n27423), .Z(n27425) );
  XOR U27377 ( .A(n27429), .B(n27430), .Z(n26999) );
  AND U27378 ( .A(n992), .B(n27431), .Z(n27430) );
  XOR U27379 ( .A(p_input[284]), .B(p_input[268]), .Z(n27431) );
  XOR U27380 ( .A(n27432), .B(n27433), .Z(n27423) );
  AND U27381 ( .A(n27434), .B(n27435), .Z(n27433) );
  XOR U27382 ( .A(n27432), .B(n27014), .Z(n27435) );
  XNOR U27383 ( .A(p_input[299]), .B(n27436), .Z(n27014) );
  AND U27384 ( .A(n995), .B(n27437), .Z(n27436) );
  XOR U27385 ( .A(p_input[315]), .B(p_input[299]), .Z(n27437) );
  XNOR U27386 ( .A(n27011), .B(n27432), .Z(n27434) );
  XOR U27387 ( .A(n27438), .B(n27439), .Z(n27011) );
  AND U27388 ( .A(n992), .B(n27440), .Z(n27439) );
  XOR U27389 ( .A(p_input[283]), .B(p_input[267]), .Z(n27440) );
  XOR U27390 ( .A(n27441), .B(n27442), .Z(n27432) );
  AND U27391 ( .A(n27443), .B(n27444), .Z(n27442) );
  XOR U27392 ( .A(n27441), .B(n27026), .Z(n27444) );
  XNOR U27393 ( .A(p_input[298]), .B(n27445), .Z(n27026) );
  AND U27394 ( .A(n995), .B(n27446), .Z(n27445) );
  XOR U27395 ( .A(p_input[314]), .B(p_input[298]), .Z(n27446) );
  XNOR U27396 ( .A(n27023), .B(n27441), .Z(n27443) );
  XOR U27397 ( .A(n27447), .B(n27448), .Z(n27023) );
  AND U27398 ( .A(n992), .B(n27449), .Z(n27448) );
  XOR U27399 ( .A(p_input[282]), .B(p_input[266]), .Z(n27449) );
  XOR U27400 ( .A(n27450), .B(n27451), .Z(n27441) );
  AND U27401 ( .A(n27452), .B(n27453), .Z(n27451) );
  XOR U27402 ( .A(n27450), .B(n27038), .Z(n27453) );
  XNOR U27403 ( .A(p_input[297]), .B(n27454), .Z(n27038) );
  AND U27404 ( .A(n995), .B(n27455), .Z(n27454) );
  XOR U27405 ( .A(p_input[313]), .B(p_input[297]), .Z(n27455) );
  XNOR U27406 ( .A(n27035), .B(n27450), .Z(n27452) );
  XOR U27407 ( .A(n27456), .B(n27457), .Z(n27035) );
  AND U27408 ( .A(n992), .B(n27458), .Z(n27457) );
  XOR U27409 ( .A(p_input[281]), .B(p_input[265]), .Z(n27458) );
  XOR U27410 ( .A(n27459), .B(n27460), .Z(n27450) );
  AND U27411 ( .A(n27461), .B(n27462), .Z(n27460) );
  XOR U27412 ( .A(n27459), .B(n27050), .Z(n27462) );
  XNOR U27413 ( .A(p_input[296]), .B(n27463), .Z(n27050) );
  AND U27414 ( .A(n995), .B(n27464), .Z(n27463) );
  XOR U27415 ( .A(p_input[312]), .B(p_input[296]), .Z(n27464) );
  XNOR U27416 ( .A(n27047), .B(n27459), .Z(n27461) );
  XOR U27417 ( .A(n27465), .B(n27466), .Z(n27047) );
  AND U27418 ( .A(n992), .B(n27467), .Z(n27466) );
  XOR U27419 ( .A(p_input[280]), .B(p_input[264]), .Z(n27467) );
  XOR U27420 ( .A(n27468), .B(n27469), .Z(n27459) );
  AND U27421 ( .A(n27470), .B(n27471), .Z(n27469) );
  XOR U27422 ( .A(n27468), .B(n27062), .Z(n27471) );
  XNOR U27423 ( .A(p_input[295]), .B(n27472), .Z(n27062) );
  AND U27424 ( .A(n995), .B(n27473), .Z(n27472) );
  XOR U27425 ( .A(p_input[311]), .B(p_input[295]), .Z(n27473) );
  XNOR U27426 ( .A(n27059), .B(n27468), .Z(n27470) );
  XOR U27427 ( .A(n27474), .B(n27475), .Z(n27059) );
  AND U27428 ( .A(n992), .B(n27476), .Z(n27475) );
  XOR U27429 ( .A(p_input[279]), .B(p_input[263]), .Z(n27476) );
  XOR U27430 ( .A(n27477), .B(n27478), .Z(n27468) );
  AND U27431 ( .A(n27479), .B(n27480), .Z(n27478) );
  XOR U27432 ( .A(n27477), .B(n27074), .Z(n27480) );
  XNOR U27433 ( .A(p_input[294]), .B(n27481), .Z(n27074) );
  AND U27434 ( .A(n995), .B(n27482), .Z(n27481) );
  XOR U27435 ( .A(p_input[310]), .B(p_input[294]), .Z(n27482) );
  XNOR U27436 ( .A(n27071), .B(n27477), .Z(n27479) );
  XOR U27437 ( .A(n27483), .B(n27484), .Z(n27071) );
  AND U27438 ( .A(n992), .B(n27485), .Z(n27484) );
  XOR U27439 ( .A(p_input[278]), .B(p_input[262]), .Z(n27485) );
  XOR U27440 ( .A(n27486), .B(n27487), .Z(n27477) );
  AND U27441 ( .A(n27488), .B(n27489), .Z(n27487) );
  XOR U27442 ( .A(n27486), .B(n27086), .Z(n27489) );
  XNOR U27443 ( .A(p_input[293]), .B(n27490), .Z(n27086) );
  AND U27444 ( .A(n995), .B(n27491), .Z(n27490) );
  XOR U27445 ( .A(p_input[309]), .B(p_input[293]), .Z(n27491) );
  XNOR U27446 ( .A(n27083), .B(n27486), .Z(n27488) );
  XOR U27447 ( .A(n27492), .B(n27493), .Z(n27083) );
  AND U27448 ( .A(n992), .B(n27494), .Z(n27493) );
  XOR U27449 ( .A(p_input[277]), .B(p_input[261]), .Z(n27494) );
  XOR U27450 ( .A(n27495), .B(n27496), .Z(n27486) );
  AND U27451 ( .A(n27497), .B(n27498), .Z(n27496) );
  XOR U27452 ( .A(n27495), .B(n27098), .Z(n27498) );
  XNOR U27453 ( .A(p_input[292]), .B(n27499), .Z(n27098) );
  AND U27454 ( .A(n995), .B(n27500), .Z(n27499) );
  XOR U27455 ( .A(p_input[308]), .B(p_input[292]), .Z(n27500) );
  XNOR U27456 ( .A(n27095), .B(n27495), .Z(n27497) );
  XOR U27457 ( .A(n27501), .B(n27502), .Z(n27095) );
  AND U27458 ( .A(n992), .B(n27503), .Z(n27502) );
  XOR U27459 ( .A(p_input[276]), .B(p_input[260]), .Z(n27503) );
  XOR U27460 ( .A(n27504), .B(n27505), .Z(n27495) );
  AND U27461 ( .A(n27506), .B(n27507), .Z(n27505) );
  XOR U27462 ( .A(n27504), .B(n27110), .Z(n27507) );
  XNOR U27463 ( .A(p_input[291]), .B(n27508), .Z(n27110) );
  AND U27464 ( .A(n995), .B(n27509), .Z(n27508) );
  XOR U27465 ( .A(p_input[307]), .B(p_input[291]), .Z(n27509) );
  XNOR U27466 ( .A(n27107), .B(n27504), .Z(n27506) );
  XOR U27467 ( .A(n27510), .B(n27511), .Z(n27107) );
  AND U27468 ( .A(n992), .B(n27512), .Z(n27511) );
  XOR U27469 ( .A(p_input[275]), .B(p_input[259]), .Z(n27512) );
  XOR U27470 ( .A(n27513), .B(n27514), .Z(n27504) );
  AND U27471 ( .A(n27515), .B(n27516), .Z(n27514) );
  XOR U27472 ( .A(n27513), .B(n27122), .Z(n27516) );
  XNOR U27473 ( .A(p_input[290]), .B(n27517), .Z(n27122) );
  AND U27474 ( .A(n995), .B(n27518), .Z(n27517) );
  XOR U27475 ( .A(p_input[306]), .B(p_input[290]), .Z(n27518) );
  XNOR U27476 ( .A(n27119), .B(n27513), .Z(n27515) );
  XOR U27477 ( .A(n27519), .B(n27520), .Z(n27119) );
  AND U27478 ( .A(n992), .B(n27521), .Z(n27520) );
  XOR U27479 ( .A(p_input[274]), .B(p_input[258]), .Z(n27521) );
  XOR U27480 ( .A(n27522), .B(n27523), .Z(n27513) );
  AND U27481 ( .A(n27524), .B(n27525), .Z(n27523) );
  XNOR U27482 ( .A(n27526), .B(n27135), .Z(n27525) );
  XNOR U27483 ( .A(p_input[289]), .B(n27527), .Z(n27135) );
  AND U27484 ( .A(n995), .B(n27528), .Z(n27527) );
  XNOR U27485 ( .A(p_input[305]), .B(n27529), .Z(n27528) );
  IV U27486 ( .A(p_input[289]), .Z(n27529) );
  XNOR U27487 ( .A(n27132), .B(n27522), .Z(n27524) );
  XNOR U27488 ( .A(p_input[257]), .B(n27530), .Z(n27132) );
  AND U27489 ( .A(n992), .B(n27531), .Z(n27530) );
  XOR U27490 ( .A(p_input[273]), .B(p_input[257]), .Z(n27531) );
  IV U27491 ( .A(n27526), .Z(n27522) );
  AND U27492 ( .A(n27397), .B(n27400), .Z(n27526) );
  XOR U27493 ( .A(p_input[288]), .B(n27532), .Z(n27400) );
  AND U27494 ( .A(n995), .B(n27533), .Z(n27532) );
  XOR U27495 ( .A(p_input[304]), .B(p_input[288]), .Z(n27533) );
  XOR U27496 ( .A(n27534), .B(n27535), .Z(n995) );
  AND U27497 ( .A(n27536), .B(n27537), .Z(n27535) );
  XNOR U27498 ( .A(p_input[319]), .B(n27534), .Z(n27537) );
  XOR U27499 ( .A(n27534), .B(p_input[303]), .Z(n27536) );
  XOR U27500 ( .A(n27538), .B(n27539), .Z(n27534) );
  AND U27501 ( .A(n27540), .B(n27541), .Z(n27539) );
  XNOR U27502 ( .A(p_input[318]), .B(n27538), .Z(n27541) );
  XOR U27503 ( .A(n27538), .B(p_input[302]), .Z(n27540) );
  XOR U27504 ( .A(n27542), .B(n27543), .Z(n27538) );
  AND U27505 ( .A(n27544), .B(n27545), .Z(n27543) );
  XNOR U27506 ( .A(p_input[317]), .B(n27542), .Z(n27545) );
  XOR U27507 ( .A(n27542), .B(p_input[301]), .Z(n27544) );
  XOR U27508 ( .A(n27546), .B(n27547), .Z(n27542) );
  AND U27509 ( .A(n27548), .B(n27549), .Z(n27547) );
  XNOR U27510 ( .A(p_input[316]), .B(n27546), .Z(n27549) );
  XOR U27511 ( .A(n27546), .B(p_input[300]), .Z(n27548) );
  XOR U27512 ( .A(n27550), .B(n27551), .Z(n27546) );
  AND U27513 ( .A(n27552), .B(n27553), .Z(n27551) );
  XNOR U27514 ( .A(p_input[315]), .B(n27550), .Z(n27553) );
  XOR U27515 ( .A(n27550), .B(p_input[299]), .Z(n27552) );
  XOR U27516 ( .A(n27554), .B(n27555), .Z(n27550) );
  AND U27517 ( .A(n27556), .B(n27557), .Z(n27555) );
  XNOR U27518 ( .A(p_input[314]), .B(n27554), .Z(n27557) );
  XOR U27519 ( .A(n27554), .B(p_input[298]), .Z(n27556) );
  XOR U27520 ( .A(n27558), .B(n27559), .Z(n27554) );
  AND U27521 ( .A(n27560), .B(n27561), .Z(n27559) );
  XNOR U27522 ( .A(p_input[313]), .B(n27558), .Z(n27561) );
  XOR U27523 ( .A(n27558), .B(p_input[297]), .Z(n27560) );
  XOR U27524 ( .A(n27562), .B(n27563), .Z(n27558) );
  AND U27525 ( .A(n27564), .B(n27565), .Z(n27563) );
  XNOR U27526 ( .A(p_input[312]), .B(n27562), .Z(n27565) );
  XOR U27527 ( .A(n27562), .B(p_input[296]), .Z(n27564) );
  XOR U27528 ( .A(n27566), .B(n27567), .Z(n27562) );
  AND U27529 ( .A(n27568), .B(n27569), .Z(n27567) );
  XNOR U27530 ( .A(p_input[311]), .B(n27566), .Z(n27569) );
  XOR U27531 ( .A(n27566), .B(p_input[295]), .Z(n27568) );
  XOR U27532 ( .A(n27570), .B(n27571), .Z(n27566) );
  AND U27533 ( .A(n27572), .B(n27573), .Z(n27571) );
  XNOR U27534 ( .A(p_input[310]), .B(n27570), .Z(n27573) );
  XOR U27535 ( .A(n27570), .B(p_input[294]), .Z(n27572) );
  XOR U27536 ( .A(n27574), .B(n27575), .Z(n27570) );
  AND U27537 ( .A(n27576), .B(n27577), .Z(n27575) );
  XNOR U27538 ( .A(p_input[309]), .B(n27574), .Z(n27577) );
  XOR U27539 ( .A(n27574), .B(p_input[293]), .Z(n27576) );
  XOR U27540 ( .A(n27578), .B(n27579), .Z(n27574) );
  AND U27541 ( .A(n27580), .B(n27581), .Z(n27579) );
  XNOR U27542 ( .A(p_input[308]), .B(n27578), .Z(n27581) );
  XOR U27543 ( .A(n27578), .B(p_input[292]), .Z(n27580) );
  XOR U27544 ( .A(n27582), .B(n27583), .Z(n27578) );
  AND U27545 ( .A(n27584), .B(n27585), .Z(n27583) );
  XNOR U27546 ( .A(p_input[307]), .B(n27582), .Z(n27585) );
  XOR U27547 ( .A(n27582), .B(p_input[291]), .Z(n27584) );
  XOR U27548 ( .A(n27586), .B(n27587), .Z(n27582) );
  AND U27549 ( .A(n27588), .B(n27589), .Z(n27587) );
  XNOR U27550 ( .A(p_input[306]), .B(n27586), .Z(n27589) );
  XOR U27551 ( .A(n27586), .B(p_input[290]), .Z(n27588) );
  XNOR U27552 ( .A(n27590), .B(n27591), .Z(n27586) );
  AND U27553 ( .A(n27592), .B(n27593), .Z(n27591) );
  XOR U27554 ( .A(p_input[305]), .B(n27590), .Z(n27593) );
  XNOR U27555 ( .A(p_input[289]), .B(n27590), .Z(n27592) );
  AND U27556 ( .A(p_input[304]), .B(n27594), .Z(n27590) );
  IV U27557 ( .A(p_input[288]), .Z(n27594) );
  XNOR U27558 ( .A(p_input[256]), .B(n27595), .Z(n27397) );
  AND U27559 ( .A(n992), .B(n27596), .Z(n27595) );
  XOR U27560 ( .A(p_input[272]), .B(p_input[256]), .Z(n27596) );
  XOR U27561 ( .A(n27597), .B(n27598), .Z(n992) );
  AND U27562 ( .A(n27599), .B(n27600), .Z(n27598) );
  XNOR U27563 ( .A(p_input[287]), .B(n27597), .Z(n27600) );
  XOR U27564 ( .A(n27597), .B(p_input[271]), .Z(n27599) );
  XOR U27565 ( .A(n27601), .B(n27602), .Z(n27597) );
  AND U27566 ( .A(n27603), .B(n27604), .Z(n27602) );
  XNOR U27567 ( .A(p_input[286]), .B(n27601), .Z(n27604) );
  XNOR U27568 ( .A(n27601), .B(n27411), .Z(n27603) );
  IV U27569 ( .A(p_input[270]), .Z(n27411) );
  XOR U27570 ( .A(n27605), .B(n27606), .Z(n27601) );
  AND U27571 ( .A(n27607), .B(n27608), .Z(n27606) );
  XNOR U27572 ( .A(p_input[285]), .B(n27605), .Z(n27608) );
  XNOR U27573 ( .A(n27605), .B(n27420), .Z(n27607) );
  IV U27574 ( .A(p_input[269]), .Z(n27420) );
  XOR U27575 ( .A(n27609), .B(n27610), .Z(n27605) );
  AND U27576 ( .A(n27611), .B(n27612), .Z(n27610) );
  XNOR U27577 ( .A(p_input[284]), .B(n27609), .Z(n27612) );
  XNOR U27578 ( .A(n27609), .B(n27429), .Z(n27611) );
  IV U27579 ( .A(p_input[268]), .Z(n27429) );
  XOR U27580 ( .A(n27613), .B(n27614), .Z(n27609) );
  AND U27581 ( .A(n27615), .B(n27616), .Z(n27614) );
  XNOR U27582 ( .A(p_input[283]), .B(n27613), .Z(n27616) );
  XNOR U27583 ( .A(n27613), .B(n27438), .Z(n27615) );
  IV U27584 ( .A(p_input[267]), .Z(n27438) );
  XOR U27585 ( .A(n27617), .B(n27618), .Z(n27613) );
  AND U27586 ( .A(n27619), .B(n27620), .Z(n27618) );
  XNOR U27587 ( .A(p_input[282]), .B(n27617), .Z(n27620) );
  XNOR U27588 ( .A(n27617), .B(n27447), .Z(n27619) );
  IV U27589 ( .A(p_input[266]), .Z(n27447) );
  XOR U27590 ( .A(n27621), .B(n27622), .Z(n27617) );
  AND U27591 ( .A(n27623), .B(n27624), .Z(n27622) );
  XNOR U27592 ( .A(p_input[281]), .B(n27621), .Z(n27624) );
  XNOR U27593 ( .A(n27621), .B(n27456), .Z(n27623) );
  IV U27594 ( .A(p_input[265]), .Z(n27456) );
  XOR U27595 ( .A(n27625), .B(n27626), .Z(n27621) );
  AND U27596 ( .A(n27627), .B(n27628), .Z(n27626) );
  XNOR U27597 ( .A(p_input[280]), .B(n27625), .Z(n27628) );
  XNOR U27598 ( .A(n27625), .B(n27465), .Z(n27627) );
  IV U27599 ( .A(p_input[264]), .Z(n27465) );
  XOR U27600 ( .A(n27629), .B(n27630), .Z(n27625) );
  AND U27601 ( .A(n27631), .B(n27632), .Z(n27630) );
  XNOR U27602 ( .A(p_input[279]), .B(n27629), .Z(n27632) );
  XNOR U27603 ( .A(n27629), .B(n27474), .Z(n27631) );
  IV U27604 ( .A(p_input[263]), .Z(n27474) );
  XOR U27605 ( .A(n27633), .B(n27634), .Z(n27629) );
  AND U27606 ( .A(n27635), .B(n27636), .Z(n27634) );
  XNOR U27607 ( .A(p_input[278]), .B(n27633), .Z(n27636) );
  XNOR U27608 ( .A(n27633), .B(n27483), .Z(n27635) );
  IV U27609 ( .A(p_input[262]), .Z(n27483) );
  XOR U27610 ( .A(n27637), .B(n27638), .Z(n27633) );
  AND U27611 ( .A(n27639), .B(n27640), .Z(n27638) );
  XNOR U27612 ( .A(p_input[277]), .B(n27637), .Z(n27640) );
  XNOR U27613 ( .A(n27637), .B(n27492), .Z(n27639) );
  IV U27614 ( .A(p_input[261]), .Z(n27492) );
  XOR U27615 ( .A(n27641), .B(n27642), .Z(n27637) );
  AND U27616 ( .A(n27643), .B(n27644), .Z(n27642) );
  XNOR U27617 ( .A(p_input[276]), .B(n27641), .Z(n27644) );
  XNOR U27618 ( .A(n27641), .B(n27501), .Z(n27643) );
  IV U27619 ( .A(p_input[260]), .Z(n27501) );
  XOR U27620 ( .A(n27645), .B(n27646), .Z(n27641) );
  AND U27621 ( .A(n27647), .B(n27648), .Z(n27646) );
  XNOR U27622 ( .A(p_input[275]), .B(n27645), .Z(n27648) );
  XNOR U27623 ( .A(n27645), .B(n27510), .Z(n27647) );
  IV U27624 ( .A(p_input[259]), .Z(n27510) );
  XOR U27625 ( .A(n27649), .B(n27650), .Z(n27645) );
  AND U27626 ( .A(n27651), .B(n27652), .Z(n27650) );
  XNOR U27627 ( .A(p_input[274]), .B(n27649), .Z(n27652) );
  XNOR U27628 ( .A(n27649), .B(n27519), .Z(n27651) );
  IV U27629 ( .A(p_input[258]), .Z(n27519) );
  XNOR U27630 ( .A(n27653), .B(n27654), .Z(n27649) );
  AND U27631 ( .A(n27655), .B(n27656), .Z(n27654) );
  XOR U27632 ( .A(p_input[273]), .B(n27653), .Z(n27656) );
  XNOR U27633 ( .A(p_input[257]), .B(n27653), .Z(n27655) );
  AND U27634 ( .A(p_input[272]), .B(n27657), .Z(n27653) );
  IV U27635 ( .A(p_input[256]), .Z(n27657) );
  XOR U27636 ( .A(n27658), .B(n27659), .Z(n25885) );
  AND U27637 ( .A(n960), .B(n27660), .Z(n27659) );
  XNOR U27638 ( .A(n27661), .B(n27658), .Z(n27660) );
  XOR U27639 ( .A(n27662), .B(n27663), .Z(n960) );
  AND U27640 ( .A(n27664), .B(n27665), .Z(n27663) );
  XNOR U27641 ( .A(n25900), .B(n27662), .Z(n27665) );
  AND U27642 ( .A(n27666), .B(n27667), .Z(n25900) );
  XNOR U27643 ( .A(n27662), .B(n25897), .Z(n27664) );
  IV U27644 ( .A(n27668), .Z(n25897) );
  AND U27645 ( .A(n27669), .B(n27670), .Z(n27668) );
  XOR U27646 ( .A(n27671), .B(n27672), .Z(n27662) );
  AND U27647 ( .A(n27673), .B(n27674), .Z(n27672) );
  XOR U27648 ( .A(n27671), .B(n25912), .Z(n27674) );
  XOR U27649 ( .A(n27675), .B(n27676), .Z(n25912) );
  AND U27650 ( .A(n839), .B(n27677), .Z(n27676) );
  XOR U27651 ( .A(n27678), .B(n27675), .Z(n27677) );
  XNOR U27652 ( .A(n25909), .B(n27671), .Z(n27673) );
  XOR U27653 ( .A(n27679), .B(n27680), .Z(n25909) );
  AND U27654 ( .A(n836), .B(n27681), .Z(n27680) );
  XOR U27655 ( .A(n27682), .B(n27679), .Z(n27681) );
  XOR U27656 ( .A(n27683), .B(n27684), .Z(n27671) );
  AND U27657 ( .A(n27685), .B(n27686), .Z(n27684) );
  XOR U27658 ( .A(n27683), .B(n25924), .Z(n27686) );
  XOR U27659 ( .A(n27687), .B(n27688), .Z(n25924) );
  AND U27660 ( .A(n839), .B(n27689), .Z(n27688) );
  XOR U27661 ( .A(n27690), .B(n27687), .Z(n27689) );
  XNOR U27662 ( .A(n25921), .B(n27683), .Z(n27685) );
  XOR U27663 ( .A(n27691), .B(n27692), .Z(n25921) );
  AND U27664 ( .A(n836), .B(n27693), .Z(n27692) );
  XOR U27665 ( .A(n27694), .B(n27691), .Z(n27693) );
  XOR U27666 ( .A(n27695), .B(n27696), .Z(n27683) );
  AND U27667 ( .A(n27697), .B(n27698), .Z(n27696) );
  XOR U27668 ( .A(n27695), .B(n25936), .Z(n27698) );
  XOR U27669 ( .A(n27699), .B(n27700), .Z(n25936) );
  AND U27670 ( .A(n839), .B(n27701), .Z(n27700) );
  XOR U27671 ( .A(n27702), .B(n27699), .Z(n27701) );
  XNOR U27672 ( .A(n25933), .B(n27695), .Z(n27697) );
  XOR U27673 ( .A(n27703), .B(n27704), .Z(n25933) );
  AND U27674 ( .A(n836), .B(n27705), .Z(n27704) );
  XOR U27675 ( .A(n27706), .B(n27703), .Z(n27705) );
  XOR U27676 ( .A(n27707), .B(n27708), .Z(n27695) );
  AND U27677 ( .A(n27709), .B(n27710), .Z(n27708) );
  XOR U27678 ( .A(n27707), .B(n25948), .Z(n27710) );
  XOR U27679 ( .A(n27711), .B(n27712), .Z(n25948) );
  AND U27680 ( .A(n839), .B(n27713), .Z(n27712) );
  XOR U27681 ( .A(n27714), .B(n27711), .Z(n27713) );
  XNOR U27682 ( .A(n25945), .B(n27707), .Z(n27709) );
  XOR U27683 ( .A(n27715), .B(n27716), .Z(n25945) );
  AND U27684 ( .A(n836), .B(n27717), .Z(n27716) );
  XOR U27685 ( .A(n27718), .B(n27715), .Z(n27717) );
  XOR U27686 ( .A(n27719), .B(n27720), .Z(n27707) );
  AND U27687 ( .A(n27721), .B(n27722), .Z(n27720) );
  XOR U27688 ( .A(n27719), .B(n25960), .Z(n27722) );
  XOR U27689 ( .A(n27723), .B(n27724), .Z(n25960) );
  AND U27690 ( .A(n839), .B(n27725), .Z(n27724) );
  XOR U27691 ( .A(n27726), .B(n27723), .Z(n27725) );
  XNOR U27692 ( .A(n25957), .B(n27719), .Z(n27721) );
  XOR U27693 ( .A(n27727), .B(n27728), .Z(n25957) );
  AND U27694 ( .A(n836), .B(n27729), .Z(n27728) );
  XOR U27695 ( .A(n27730), .B(n27727), .Z(n27729) );
  XOR U27696 ( .A(n27731), .B(n27732), .Z(n27719) );
  AND U27697 ( .A(n27733), .B(n27734), .Z(n27732) );
  XOR U27698 ( .A(n27731), .B(n25972), .Z(n27734) );
  XOR U27699 ( .A(n27735), .B(n27736), .Z(n25972) );
  AND U27700 ( .A(n839), .B(n27737), .Z(n27736) );
  XOR U27701 ( .A(n27738), .B(n27735), .Z(n27737) );
  XNOR U27702 ( .A(n25969), .B(n27731), .Z(n27733) );
  XOR U27703 ( .A(n27739), .B(n27740), .Z(n25969) );
  AND U27704 ( .A(n836), .B(n27741), .Z(n27740) );
  XOR U27705 ( .A(n27742), .B(n27739), .Z(n27741) );
  XOR U27706 ( .A(n27743), .B(n27744), .Z(n27731) );
  AND U27707 ( .A(n27745), .B(n27746), .Z(n27744) );
  XOR U27708 ( .A(n27743), .B(n25984), .Z(n27746) );
  XOR U27709 ( .A(n27747), .B(n27748), .Z(n25984) );
  AND U27710 ( .A(n839), .B(n27749), .Z(n27748) );
  XOR U27711 ( .A(n27750), .B(n27747), .Z(n27749) );
  XNOR U27712 ( .A(n25981), .B(n27743), .Z(n27745) );
  XOR U27713 ( .A(n27751), .B(n27752), .Z(n25981) );
  AND U27714 ( .A(n836), .B(n27753), .Z(n27752) );
  XOR U27715 ( .A(n27754), .B(n27751), .Z(n27753) );
  XOR U27716 ( .A(n27755), .B(n27756), .Z(n27743) );
  AND U27717 ( .A(n27757), .B(n27758), .Z(n27756) );
  XOR U27718 ( .A(n27755), .B(n25996), .Z(n27758) );
  XOR U27719 ( .A(n27759), .B(n27760), .Z(n25996) );
  AND U27720 ( .A(n839), .B(n27761), .Z(n27760) );
  XOR U27721 ( .A(n27762), .B(n27759), .Z(n27761) );
  XNOR U27722 ( .A(n25993), .B(n27755), .Z(n27757) );
  XOR U27723 ( .A(n27763), .B(n27764), .Z(n25993) );
  AND U27724 ( .A(n836), .B(n27765), .Z(n27764) );
  XOR U27725 ( .A(n27766), .B(n27763), .Z(n27765) );
  XOR U27726 ( .A(n27767), .B(n27768), .Z(n27755) );
  AND U27727 ( .A(n27769), .B(n27770), .Z(n27768) );
  XOR U27728 ( .A(n27767), .B(n26008), .Z(n27770) );
  XOR U27729 ( .A(n27771), .B(n27772), .Z(n26008) );
  AND U27730 ( .A(n839), .B(n27773), .Z(n27772) );
  XOR U27731 ( .A(n27774), .B(n27771), .Z(n27773) );
  XNOR U27732 ( .A(n26005), .B(n27767), .Z(n27769) );
  XOR U27733 ( .A(n27775), .B(n27776), .Z(n26005) );
  AND U27734 ( .A(n836), .B(n27777), .Z(n27776) );
  XOR U27735 ( .A(n27778), .B(n27775), .Z(n27777) );
  XOR U27736 ( .A(n27779), .B(n27780), .Z(n27767) );
  AND U27737 ( .A(n27781), .B(n27782), .Z(n27780) );
  XOR U27738 ( .A(n27779), .B(n26020), .Z(n27782) );
  XOR U27739 ( .A(n27783), .B(n27784), .Z(n26020) );
  AND U27740 ( .A(n839), .B(n27785), .Z(n27784) );
  XOR U27741 ( .A(n27786), .B(n27783), .Z(n27785) );
  XNOR U27742 ( .A(n26017), .B(n27779), .Z(n27781) );
  XOR U27743 ( .A(n27787), .B(n27788), .Z(n26017) );
  AND U27744 ( .A(n836), .B(n27789), .Z(n27788) );
  XOR U27745 ( .A(n27790), .B(n27787), .Z(n27789) );
  XOR U27746 ( .A(n27791), .B(n27792), .Z(n27779) );
  AND U27747 ( .A(n27793), .B(n27794), .Z(n27792) );
  XOR U27748 ( .A(n27791), .B(n26032), .Z(n27794) );
  XOR U27749 ( .A(n27795), .B(n27796), .Z(n26032) );
  AND U27750 ( .A(n839), .B(n27797), .Z(n27796) );
  XOR U27751 ( .A(n27798), .B(n27795), .Z(n27797) );
  XNOR U27752 ( .A(n26029), .B(n27791), .Z(n27793) );
  XOR U27753 ( .A(n27799), .B(n27800), .Z(n26029) );
  AND U27754 ( .A(n836), .B(n27801), .Z(n27800) );
  XOR U27755 ( .A(n27802), .B(n27799), .Z(n27801) );
  XOR U27756 ( .A(n27803), .B(n27804), .Z(n27791) );
  AND U27757 ( .A(n27805), .B(n27806), .Z(n27804) );
  XOR U27758 ( .A(n27803), .B(n26044), .Z(n27806) );
  XOR U27759 ( .A(n27807), .B(n27808), .Z(n26044) );
  AND U27760 ( .A(n839), .B(n27809), .Z(n27808) );
  XOR U27761 ( .A(n27810), .B(n27807), .Z(n27809) );
  XNOR U27762 ( .A(n26041), .B(n27803), .Z(n27805) );
  XOR U27763 ( .A(n27811), .B(n27812), .Z(n26041) );
  AND U27764 ( .A(n836), .B(n27813), .Z(n27812) );
  XOR U27765 ( .A(n27814), .B(n27811), .Z(n27813) );
  XOR U27766 ( .A(n27815), .B(n27816), .Z(n27803) );
  AND U27767 ( .A(n27817), .B(n27818), .Z(n27816) );
  XOR U27768 ( .A(n27815), .B(n26056), .Z(n27818) );
  XOR U27769 ( .A(n27819), .B(n27820), .Z(n26056) );
  AND U27770 ( .A(n839), .B(n27821), .Z(n27820) );
  XOR U27771 ( .A(n27822), .B(n27819), .Z(n27821) );
  XNOR U27772 ( .A(n26053), .B(n27815), .Z(n27817) );
  XOR U27773 ( .A(n27823), .B(n27824), .Z(n26053) );
  AND U27774 ( .A(n836), .B(n27825), .Z(n27824) );
  XOR U27775 ( .A(n27826), .B(n27823), .Z(n27825) );
  XOR U27776 ( .A(n27827), .B(n27828), .Z(n27815) );
  AND U27777 ( .A(n27829), .B(n27830), .Z(n27828) );
  XNOR U27778 ( .A(n27831), .B(n26069), .Z(n27830) );
  XOR U27779 ( .A(n27832), .B(n27833), .Z(n26069) );
  AND U27780 ( .A(n839), .B(n27834), .Z(n27833) );
  XOR U27781 ( .A(n27832), .B(n27835), .Z(n27834) );
  XNOR U27782 ( .A(n26066), .B(n27827), .Z(n27829) );
  XOR U27783 ( .A(n27836), .B(n27837), .Z(n26066) );
  AND U27784 ( .A(n836), .B(n27838), .Z(n27837) );
  XOR U27785 ( .A(n27836), .B(n27839), .Z(n27838) );
  IV U27786 ( .A(n27831), .Z(n27827) );
  AND U27787 ( .A(n27658), .B(n27661), .Z(n27831) );
  XNOR U27788 ( .A(n27840), .B(n27841), .Z(n27661) );
  AND U27789 ( .A(n839), .B(n27842), .Z(n27841) );
  XNOR U27790 ( .A(n27843), .B(n27840), .Z(n27842) );
  XOR U27791 ( .A(n27844), .B(n27845), .Z(n839) );
  AND U27792 ( .A(n27846), .B(n27847), .Z(n27845) );
  XNOR U27793 ( .A(n27666), .B(n27844), .Z(n27847) );
  AND U27794 ( .A(n27848), .B(n27849), .Z(n27666) );
  XOR U27795 ( .A(n27844), .B(n27667), .Z(n27846) );
  AND U27796 ( .A(n27850), .B(n27851), .Z(n27667) );
  XOR U27797 ( .A(n27852), .B(n27853), .Z(n27844) );
  AND U27798 ( .A(n27854), .B(n27855), .Z(n27853) );
  XOR U27799 ( .A(n27852), .B(n27678), .Z(n27855) );
  XOR U27800 ( .A(n27856), .B(n27857), .Z(n27678) );
  AND U27801 ( .A(n583), .B(n27858), .Z(n27857) );
  XOR U27802 ( .A(n27859), .B(n27856), .Z(n27858) );
  XNOR U27803 ( .A(n27675), .B(n27852), .Z(n27854) );
  XOR U27804 ( .A(n27860), .B(n27861), .Z(n27675) );
  AND U27805 ( .A(n581), .B(n27862), .Z(n27861) );
  XOR U27806 ( .A(n27863), .B(n27860), .Z(n27862) );
  XOR U27807 ( .A(n27864), .B(n27865), .Z(n27852) );
  AND U27808 ( .A(n27866), .B(n27867), .Z(n27865) );
  XOR U27809 ( .A(n27864), .B(n27690), .Z(n27867) );
  XOR U27810 ( .A(n27868), .B(n27869), .Z(n27690) );
  AND U27811 ( .A(n583), .B(n27870), .Z(n27869) );
  XOR U27812 ( .A(n27871), .B(n27868), .Z(n27870) );
  XNOR U27813 ( .A(n27687), .B(n27864), .Z(n27866) );
  XOR U27814 ( .A(n27872), .B(n27873), .Z(n27687) );
  AND U27815 ( .A(n581), .B(n27874), .Z(n27873) );
  XOR U27816 ( .A(n27875), .B(n27872), .Z(n27874) );
  XOR U27817 ( .A(n27876), .B(n27877), .Z(n27864) );
  AND U27818 ( .A(n27878), .B(n27879), .Z(n27877) );
  XOR U27819 ( .A(n27876), .B(n27702), .Z(n27879) );
  XOR U27820 ( .A(n27880), .B(n27881), .Z(n27702) );
  AND U27821 ( .A(n583), .B(n27882), .Z(n27881) );
  XOR U27822 ( .A(n27883), .B(n27880), .Z(n27882) );
  XNOR U27823 ( .A(n27699), .B(n27876), .Z(n27878) );
  XOR U27824 ( .A(n27884), .B(n27885), .Z(n27699) );
  AND U27825 ( .A(n581), .B(n27886), .Z(n27885) );
  XOR U27826 ( .A(n27887), .B(n27884), .Z(n27886) );
  XOR U27827 ( .A(n27888), .B(n27889), .Z(n27876) );
  AND U27828 ( .A(n27890), .B(n27891), .Z(n27889) );
  XOR U27829 ( .A(n27888), .B(n27714), .Z(n27891) );
  XOR U27830 ( .A(n27892), .B(n27893), .Z(n27714) );
  AND U27831 ( .A(n583), .B(n27894), .Z(n27893) );
  XOR U27832 ( .A(n27895), .B(n27892), .Z(n27894) );
  XNOR U27833 ( .A(n27711), .B(n27888), .Z(n27890) );
  XOR U27834 ( .A(n27896), .B(n27897), .Z(n27711) );
  AND U27835 ( .A(n581), .B(n27898), .Z(n27897) );
  XOR U27836 ( .A(n27899), .B(n27896), .Z(n27898) );
  XOR U27837 ( .A(n27900), .B(n27901), .Z(n27888) );
  AND U27838 ( .A(n27902), .B(n27903), .Z(n27901) );
  XOR U27839 ( .A(n27900), .B(n27726), .Z(n27903) );
  XOR U27840 ( .A(n27904), .B(n27905), .Z(n27726) );
  AND U27841 ( .A(n583), .B(n27906), .Z(n27905) );
  XOR U27842 ( .A(n27907), .B(n27904), .Z(n27906) );
  XNOR U27843 ( .A(n27723), .B(n27900), .Z(n27902) );
  XOR U27844 ( .A(n27908), .B(n27909), .Z(n27723) );
  AND U27845 ( .A(n581), .B(n27910), .Z(n27909) );
  XOR U27846 ( .A(n27911), .B(n27908), .Z(n27910) );
  XOR U27847 ( .A(n27912), .B(n27913), .Z(n27900) );
  AND U27848 ( .A(n27914), .B(n27915), .Z(n27913) );
  XOR U27849 ( .A(n27912), .B(n27738), .Z(n27915) );
  XOR U27850 ( .A(n27916), .B(n27917), .Z(n27738) );
  AND U27851 ( .A(n583), .B(n27918), .Z(n27917) );
  XOR U27852 ( .A(n27919), .B(n27916), .Z(n27918) );
  XNOR U27853 ( .A(n27735), .B(n27912), .Z(n27914) );
  XOR U27854 ( .A(n27920), .B(n27921), .Z(n27735) );
  AND U27855 ( .A(n581), .B(n27922), .Z(n27921) );
  XOR U27856 ( .A(n27923), .B(n27920), .Z(n27922) );
  XOR U27857 ( .A(n27924), .B(n27925), .Z(n27912) );
  AND U27858 ( .A(n27926), .B(n27927), .Z(n27925) );
  XOR U27859 ( .A(n27924), .B(n27750), .Z(n27927) );
  XOR U27860 ( .A(n27928), .B(n27929), .Z(n27750) );
  AND U27861 ( .A(n583), .B(n27930), .Z(n27929) );
  XOR U27862 ( .A(n27931), .B(n27928), .Z(n27930) );
  XNOR U27863 ( .A(n27747), .B(n27924), .Z(n27926) );
  XOR U27864 ( .A(n27932), .B(n27933), .Z(n27747) );
  AND U27865 ( .A(n581), .B(n27934), .Z(n27933) );
  XOR U27866 ( .A(n27935), .B(n27932), .Z(n27934) );
  XOR U27867 ( .A(n27936), .B(n27937), .Z(n27924) );
  AND U27868 ( .A(n27938), .B(n27939), .Z(n27937) );
  XOR U27869 ( .A(n27936), .B(n27762), .Z(n27939) );
  XOR U27870 ( .A(n27940), .B(n27941), .Z(n27762) );
  AND U27871 ( .A(n583), .B(n27942), .Z(n27941) );
  XOR U27872 ( .A(n27943), .B(n27940), .Z(n27942) );
  XNOR U27873 ( .A(n27759), .B(n27936), .Z(n27938) );
  XOR U27874 ( .A(n27944), .B(n27945), .Z(n27759) );
  AND U27875 ( .A(n581), .B(n27946), .Z(n27945) );
  XOR U27876 ( .A(n27947), .B(n27944), .Z(n27946) );
  XOR U27877 ( .A(n27948), .B(n27949), .Z(n27936) );
  AND U27878 ( .A(n27950), .B(n27951), .Z(n27949) );
  XOR U27879 ( .A(n27948), .B(n27774), .Z(n27951) );
  XOR U27880 ( .A(n27952), .B(n27953), .Z(n27774) );
  AND U27881 ( .A(n583), .B(n27954), .Z(n27953) );
  XOR U27882 ( .A(n27955), .B(n27952), .Z(n27954) );
  XNOR U27883 ( .A(n27771), .B(n27948), .Z(n27950) );
  XOR U27884 ( .A(n27956), .B(n27957), .Z(n27771) );
  AND U27885 ( .A(n581), .B(n27958), .Z(n27957) );
  XOR U27886 ( .A(n27959), .B(n27956), .Z(n27958) );
  XOR U27887 ( .A(n27960), .B(n27961), .Z(n27948) );
  AND U27888 ( .A(n27962), .B(n27963), .Z(n27961) );
  XOR U27889 ( .A(n27960), .B(n27786), .Z(n27963) );
  XOR U27890 ( .A(n27964), .B(n27965), .Z(n27786) );
  AND U27891 ( .A(n583), .B(n27966), .Z(n27965) );
  XOR U27892 ( .A(n27967), .B(n27964), .Z(n27966) );
  XNOR U27893 ( .A(n27783), .B(n27960), .Z(n27962) );
  XOR U27894 ( .A(n27968), .B(n27969), .Z(n27783) );
  AND U27895 ( .A(n581), .B(n27970), .Z(n27969) );
  XOR U27896 ( .A(n27971), .B(n27968), .Z(n27970) );
  XOR U27897 ( .A(n27972), .B(n27973), .Z(n27960) );
  AND U27898 ( .A(n27974), .B(n27975), .Z(n27973) );
  XOR U27899 ( .A(n27972), .B(n27798), .Z(n27975) );
  XOR U27900 ( .A(n27976), .B(n27977), .Z(n27798) );
  AND U27901 ( .A(n583), .B(n27978), .Z(n27977) );
  XOR U27902 ( .A(n27979), .B(n27976), .Z(n27978) );
  XNOR U27903 ( .A(n27795), .B(n27972), .Z(n27974) );
  XOR U27904 ( .A(n27980), .B(n27981), .Z(n27795) );
  AND U27905 ( .A(n581), .B(n27982), .Z(n27981) );
  XOR U27906 ( .A(n27983), .B(n27980), .Z(n27982) );
  XOR U27907 ( .A(n27984), .B(n27985), .Z(n27972) );
  AND U27908 ( .A(n27986), .B(n27987), .Z(n27985) );
  XOR U27909 ( .A(n27984), .B(n27810), .Z(n27987) );
  XOR U27910 ( .A(n27988), .B(n27989), .Z(n27810) );
  AND U27911 ( .A(n583), .B(n27990), .Z(n27989) );
  XOR U27912 ( .A(n27991), .B(n27988), .Z(n27990) );
  XNOR U27913 ( .A(n27807), .B(n27984), .Z(n27986) );
  XOR U27914 ( .A(n27992), .B(n27993), .Z(n27807) );
  AND U27915 ( .A(n581), .B(n27994), .Z(n27993) );
  XOR U27916 ( .A(n27995), .B(n27992), .Z(n27994) );
  XOR U27917 ( .A(n27996), .B(n27997), .Z(n27984) );
  AND U27918 ( .A(n27998), .B(n27999), .Z(n27997) );
  XOR U27919 ( .A(n27996), .B(n27822), .Z(n27999) );
  XOR U27920 ( .A(n28000), .B(n28001), .Z(n27822) );
  AND U27921 ( .A(n583), .B(n28002), .Z(n28001) );
  XOR U27922 ( .A(n28003), .B(n28000), .Z(n28002) );
  XNOR U27923 ( .A(n27819), .B(n27996), .Z(n27998) );
  XOR U27924 ( .A(n28004), .B(n28005), .Z(n27819) );
  AND U27925 ( .A(n581), .B(n28006), .Z(n28005) );
  XOR U27926 ( .A(n28007), .B(n28004), .Z(n28006) );
  XOR U27927 ( .A(n28008), .B(n28009), .Z(n27996) );
  AND U27928 ( .A(n28010), .B(n28011), .Z(n28009) );
  XNOR U27929 ( .A(n28012), .B(n27835), .Z(n28011) );
  XOR U27930 ( .A(n28013), .B(n28014), .Z(n27835) );
  AND U27931 ( .A(n583), .B(n28015), .Z(n28014) );
  XOR U27932 ( .A(n28013), .B(n28016), .Z(n28015) );
  XNOR U27933 ( .A(n27832), .B(n28008), .Z(n28010) );
  XOR U27934 ( .A(n28017), .B(n28018), .Z(n27832) );
  AND U27935 ( .A(n581), .B(n28019), .Z(n28018) );
  XOR U27936 ( .A(n28017), .B(n28020), .Z(n28019) );
  IV U27937 ( .A(n28012), .Z(n28008) );
  AND U27938 ( .A(n27840), .B(n27843), .Z(n28012) );
  XNOR U27939 ( .A(n28021), .B(n28022), .Z(n27843) );
  AND U27940 ( .A(n583), .B(n28023), .Z(n28022) );
  XNOR U27941 ( .A(n28024), .B(n28021), .Z(n28023) );
  XOR U27942 ( .A(n28025), .B(n28026), .Z(n583) );
  AND U27943 ( .A(n28027), .B(n28028), .Z(n28026) );
  XNOR U27944 ( .A(n27848), .B(n28025), .Z(n28028) );
  AND U27945 ( .A(p_input[255]), .B(p_input[239]), .Z(n27848) );
  XOR U27946 ( .A(n28025), .B(n27849), .Z(n28027) );
  AND U27947 ( .A(p_input[223]), .B(p_input[207]), .Z(n27849) );
  XOR U27948 ( .A(n28029), .B(n28030), .Z(n28025) );
  AND U27949 ( .A(n28031), .B(n28032), .Z(n28030) );
  XOR U27950 ( .A(n28029), .B(n27859), .Z(n28032) );
  XNOR U27951 ( .A(p_input[238]), .B(n28033), .Z(n27859) );
  AND U27952 ( .A(n1035), .B(n28034), .Z(n28033) );
  XOR U27953 ( .A(p_input[254]), .B(p_input[238]), .Z(n28034) );
  XNOR U27954 ( .A(n27856), .B(n28029), .Z(n28031) );
  XOR U27955 ( .A(n28035), .B(n28036), .Z(n27856) );
  AND U27956 ( .A(n1033), .B(n28037), .Z(n28036) );
  XOR U27957 ( .A(p_input[222]), .B(p_input[206]), .Z(n28037) );
  XOR U27958 ( .A(n28038), .B(n28039), .Z(n28029) );
  AND U27959 ( .A(n28040), .B(n28041), .Z(n28039) );
  XOR U27960 ( .A(n28038), .B(n27871), .Z(n28041) );
  XNOR U27961 ( .A(p_input[237]), .B(n28042), .Z(n27871) );
  AND U27962 ( .A(n1035), .B(n28043), .Z(n28042) );
  XOR U27963 ( .A(p_input[253]), .B(p_input[237]), .Z(n28043) );
  XNOR U27964 ( .A(n27868), .B(n28038), .Z(n28040) );
  XOR U27965 ( .A(n28044), .B(n28045), .Z(n27868) );
  AND U27966 ( .A(n1033), .B(n28046), .Z(n28045) );
  XOR U27967 ( .A(p_input[221]), .B(p_input[205]), .Z(n28046) );
  XOR U27968 ( .A(n28047), .B(n28048), .Z(n28038) );
  AND U27969 ( .A(n28049), .B(n28050), .Z(n28048) );
  XOR U27970 ( .A(n28047), .B(n27883), .Z(n28050) );
  XNOR U27971 ( .A(p_input[236]), .B(n28051), .Z(n27883) );
  AND U27972 ( .A(n1035), .B(n28052), .Z(n28051) );
  XOR U27973 ( .A(p_input[252]), .B(p_input[236]), .Z(n28052) );
  XNOR U27974 ( .A(n27880), .B(n28047), .Z(n28049) );
  XOR U27975 ( .A(n28053), .B(n28054), .Z(n27880) );
  AND U27976 ( .A(n1033), .B(n28055), .Z(n28054) );
  XOR U27977 ( .A(p_input[220]), .B(p_input[204]), .Z(n28055) );
  XOR U27978 ( .A(n28056), .B(n28057), .Z(n28047) );
  AND U27979 ( .A(n28058), .B(n28059), .Z(n28057) );
  XOR U27980 ( .A(n28056), .B(n27895), .Z(n28059) );
  XNOR U27981 ( .A(p_input[235]), .B(n28060), .Z(n27895) );
  AND U27982 ( .A(n1035), .B(n28061), .Z(n28060) );
  XOR U27983 ( .A(p_input[251]), .B(p_input[235]), .Z(n28061) );
  XNOR U27984 ( .A(n27892), .B(n28056), .Z(n28058) );
  XOR U27985 ( .A(n28062), .B(n28063), .Z(n27892) );
  AND U27986 ( .A(n1033), .B(n28064), .Z(n28063) );
  XOR U27987 ( .A(p_input[219]), .B(p_input[203]), .Z(n28064) );
  XOR U27988 ( .A(n28065), .B(n28066), .Z(n28056) );
  AND U27989 ( .A(n28067), .B(n28068), .Z(n28066) );
  XOR U27990 ( .A(n28065), .B(n27907), .Z(n28068) );
  XNOR U27991 ( .A(p_input[234]), .B(n28069), .Z(n27907) );
  AND U27992 ( .A(n1035), .B(n28070), .Z(n28069) );
  XOR U27993 ( .A(p_input[250]), .B(p_input[234]), .Z(n28070) );
  XNOR U27994 ( .A(n27904), .B(n28065), .Z(n28067) );
  XOR U27995 ( .A(n28071), .B(n28072), .Z(n27904) );
  AND U27996 ( .A(n1033), .B(n28073), .Z(n28072) );
  XOR U27997 ( .A(p_input[218]), .B(p_input[202]), .Z(n28073) );
  XOR U27998 ( .A(n28074), .B(n28075), .Z(n28065) );
  AND U27999 ( .A(n28076), .B(n28077), .Z(n28075) );
  XOR U28000 ( .A(n28074), .B(n27919), .Z(n28077) );
  XNOR U28001 ( .A(p_input[233]), .B(n28078), .Z(n27919) );
  AND U28002 ( .A(n1035), .B(n28079), .Z(n28078) );
  XOR U28003 ( .A(p_input[249]), .B(p_input[233]), .Z(n28079) );
  XNOR U28004 ( .A(n27916), .B(n28074), .Z(n28076) );
  XOR U28005 ( .A(n28080), .B(n28081), .Z(n27916) );
  AND U28006 ( .A(n1033), .B(n28082), .Z(n28081) );
  XOR U28007 ( .A(p_input[217]), .B(p_input[201]), .Z(n28082) );
  XOR U28008 ( .A(n28083), .B(n28084), .Z(n28074) );
  AND U28009 ( .A(n28085), .B(n28086), .Z(n28084) );
  XOR U28010 ( .A(n28083), .B(n27931), .Z(n28086) );
  XNOR U28011 ( .A(p_input[232]), .B(n28087), .Z(n27931) );
  AND U28012 ( .A(n1035), .B(n28088), .Z(n28087) );
  XOR U28013 ( .A(p_input[248]), .B(p_input[232]), .Z(n28088) );
  XNOR U28014 ( .A(n27928), .B(n28083), .Z(n28085) );
  XOR U28015 ( .A(n28089), .B(n28090), .Z(n27928) );
  AND U28016 ( .A(n1033), .B(n28091), .Z(n28090) );
  XOR U28017 ( .A(p_input[216]), .B(p_input[200]), .Z(n28091) );
  XOR U28018 ( .A(n28092), .B(n28093), .Z(n28083) );
  AND U28019 ( .A(n28094), .B(n28095), .Z(n28093) );
  XOR U28020 ( .A(n28092), .B(n27943), .Z(n28095) );
  XNOR U28021 ( .A(p_input[231]), .B(n28096), .Z(n27943) );
  AND U28022 ( .A(n1035), .B(n28097), .Z(n28096) );
  XOR U28023 ( .A(p_input[247]), .B(p_input[231]), .Z(n28097) );
  XNOR U28024 ( .A(n27940), .B(n28092), .Z(n28094) );
  XOR U28025 ( .A(n28098), .B(n28099), .Z(n27940) );
  AND U28026 ( .A(n1033), .B(n28100), .Z(n28099) );
  XOR U28027 ( .A(p_input[215]), .B(p_input[199]), .Z(n28100) );
  XOR U28028 ( .A(n28101), .B(n28102), .Z(n28092) );
  AND U28029 ( .A(n28103), .B(n28104), .Z(n28102) );
  XOR U28030 ( .A(n28101), .B(n27955), .Z(n28104) );
  XNOR U28031 ( .A(p_input[230]), .B(n28105), .Z(n27955) );
  AND U28032 ( .A(n1035), .B(n28106), .Z(n28105) );
  XOR U28033 ( .A(p_input[246]), .B(p_input[230]), .Z(n28106) );
  XNOR U28034 ( .A(n27952), .B(n28101), .Z(n28103) );
  XOR U28035 ( .A(n28107), .B(n28108), .Z(n27952) );
  AND U28036 ( .A(n1033), .B(n28109), .Z(n28108) );
  XOR U28037 ( .A(p_input[214]), .B(p_input[198]), .Z(n28109) );
  XOR U28038 ( .A(n28110), .B(n28111), .Z(n28101) );
  AND U28039 ( .A(n28112), .B(n28113), .Z(n28111) );
  XOR U28040 ( .A(n28110), .B(n27967), .Z(n28113) );
  XNOR U28041 ( .A(p_input[229]), .B(n28114), .Z(n27967) );
  AND U28042 ( .A(n1035), .B(n28115), .Z(n28114) );
  XOR U28043 ( .A(p_input[245]), .B(p_input[229]), .Z(n28115) );
  XNOR U28044 ( .A(n27964), .B(n28110), .Z(n28112) );
  XOR U28045 ( .A(n28116), .B(n28117), .Z(n27964) );
  AND U28046 ( .A(n1033), .B(n28118), .Z(n28117) );
  XOR U28047 ( .A(p_input[213]), .B(p_input[197]), .Z(n28118) );
  XOR U28048 ( .A(n28119), .B(n28120), .Z(n28110) );
  AND U28049 ( .A(n28121), .B(n28122), .Z(n28120) );
  XOR U28050 ( .A(n28119), .B(n27979), .Z(n28122) );
  XNOR U28051 ( .A(p_input[228]), .B(n28123), .Z(n27979) );
  AND U28052 ( .A(n1035), .B(n28124), .Z(n28123) );
  XOR U28053 ( .A(p_input[244]), .B(p_input[228]), .Z(n28124) );
  XNOR U28054 ( .A(n27976), .B(n28119), .Z(n28121) );
  XOR U28055 ( .A(n28125), .B(n28126), .Z(n27976) );
  AND U28056 ( .A(n1033), .B(n28127), .Z(n28126) );
  XOR U28057 ( .A(p_input[212]), .B(p_input[196]), .Z(n28127) );
  XOR U28058 ( .A(n28128), .B(n28129), .Z(n28119) );
  AND U28059 ( .A(n28130), .B(n28131), .Z(n28129) );
  XOR U28060 ( .A(n28128), .B(n27991), .Z(n28131) );
  XNOR U28061 ( .A(p_input[227]), .B(n28132), .Z(n27991) );
  AND U28062 ( .A(n1035), .B(n28133), .Z(n28132) );
  XOR U28063 ( .A(p_input[243]), .B(p_input[227]), .Z(n28133) );
  XNOR U28064 ( .A(n27988), .B(n28128), .Z(n28130) );
  XOR U28065 ( .A(n28134), .B(n28135), .Z(n27988) );
  AND U28066 ( .A(n1033), .B(n28136), .Z(n28135) );
  XOR U28067 ( .A(p_input[211]), .B(p_input[195]), .Z(n28136) );
  XOR U28068 ( .A(n28137), .B(n28138), .Z(n28128) );
  AND U28069 ( .A(n28139), .B(n28140), .Z(n28138) );
  XOR U28070 ( .A(n28137), .B(n28003), .Z(n28140) );
  XNOR U28071 ( .A(p_input[226]), .B(n28141), .Z(n28003) );
  AND U28072 ( .A(n1035), .B(n28142), .Z(n28141) );
  XOR U28073 ( .A(p_input[242]), .B(p_input[226]), .Z(n28142) );
  XNOR U28074 ( .A(n28000), .B(n28137), .Z(n28139) );
  XOR U28075 ( .A(n28143), .B(n28144), .Z(n28000) );
  AND U28076 ( .A(n1033), .B(n28145), .Z(n28144) );
  XOR U28077 ( .A(p_input[210]), .B(p_input[194]), .Z(n28145) );
  XOR U28078 ( .A(n28146), .B(n28147), .Z(n28137) );
  AND U28079 ( .A(n28148), .B(n28149), .Z(n28147) );
  XNOR U28080 ( .A(n28150), .B(n28016), .Z(n28149) );
  XNOR U28081 ( .A(p_input[225]), .B(n28151), .Z(n28016) );
  AND U28082 ( .A(n1035), .B(n28152), .Z(n28151) );
  XNOR U28083 ( .A(p_input[241]), .B(n28153), .Z(n28152) );
  IV U28084 ( .A(p_input[225]), .Z(n28153) );
  XNOR U28085 ( .A(n28013), .B(n28146), .Z(n28148) );
  XNOR U28086 ( .A(p_input[193]), .B(n28154), .Z(n28013) );
  AND U28087 ( .A(n1033), .B(n28155), .Z(n28154) );
  XOR U28088 ( .A(p_input[209]), .B(p_input[193]), .Z(n28155) );
  IV U28089 ( .A(n28150), .Z(n28146) );
  AND U28090 ( .A(n28021), .B(n28024), .Z(n28150) );
  XOR U28091 ( .A(p_input[224]), .B(n28156), .Z(n28024) );
  AND U28092 ( .A(n1035), .B(n28157), .Z(n28156) );
  XOR U28093 ( .A(p_input[240]), .B(p_input[224]), .Z(n28157) );
  XOR U28094 ( .A(n28158), .B(n28159), .Z(n1035) );
  AND U28095 ( .A(n28160), .B(n28161), .Z(n28159) );
  XNOR U28096 ( .A(p_input[255]), .B(n28158), .Z(n28161) );
  XOR U28097 ( .A(n28158), .B(p_input[239]), .Z(n28160) );
  XOR U28098 ( .A(n28162), .B(n28163), .Z(n28158) );
  AND U28099 ( .A(n28164), .B(n28165), .Z(n28163) );
  XNOR U28100 ( .A(p_input[254]), .B(n28162), .Z(n28165) );
  XOR U28101 ( .A(n28162), .B(p_input[238]), .Z(n28164) );
  XOR U28102 ( .A(n28166), .B(n28167), .Z(n28162) );
  AND U28103 ( .A(n28168), .B(n28169), .Z(n28167) );
  XNOR U28104 ( .A(p_input[253]), .B(n28166), .Z(n28169) );
  XOR U28105 ( .A(n28166), .B(p_input[237]), .Z(n28168) );
  XOR U28106 ( .A(n28170), .B(n28171), .Z(n28166) );
  AND U28107 ( .A(n28172), .B(n28173), .Z(n28171) );
  XNOR U28108 ( .A(p_input[252]), .B(n28170), .Z(n28173) );
  XOR U28109 ( .A(n28170), .B(p_input[236]), .Z(n28172) );
  XOR U28110 ( .A(n28174), .B(n28175), .Z(n28170) );
  AND U28111 ( .A(n28176), .B(n28177), .Z(n28175) );
  XNOR U28112 ( .A(p_input[251]), .B(n28174), .Z(n28177) );
  XOR U28113 ( .A(n28174), .B(p_input[235]), .Z(n28176) );
  XOR U28114 ( .A(n28178), .B(n28179), .Z(n28174) );
  AND U28115 ( .A(n28180), .B(n28181), .Z(n28179) );
  XNOR U28116 ( .A(p_input[250]), .B(n28178), .Z(n28181) );
  XOR U28117 ( .A(n28178), .B(p_input[234]), .Z(n28180) );
  XOR U28118 ( .A(n28182), .B(n28183), .Z(n28178) );
  AND U28119 ( .A(n28184), .B(n28185), .Z(n28183) );
  XNOR U28120 ( .A(p_input[249]), .B(n28182), .Z(n28185) );
  XOR U28121 ( .A(n28182), .B(p_input[233]), .Z(n28184) );
  XOR U28122 ( .A(n28186), .B(n28187), .Z(n28182) );
  AND U28123 ( .A(n28188), .B(n28189), .Z(n28187) );
  XNOR U28124 ( .A(p_input[248]), .B(n28186), .Z(n28189) );
  XOR U28125 ( .A(n28186), .B(p_input[232]), .Z(n28188) );
  XOR U28126 ( .A(n28190), .B(n28191), .Z(n28186) );
  AND U28127 ( .A(n28192), .B(n28193), .Z(n28191) );
  XNOR U28128 ( .A(p_input[247]), .B(n28190), .Z(n28193) );
  XOR U28129 ( .A(n28190), .B(p_input[231]), .Z(n28192) );
  XOR U28130 ( .A(n28194), .B(n28195), .Z(n28190) );
  AND U28131 ( .A(n28196), .B(n28197), .Z(n28195) );
  XNOR U28132 ( .A(p_input[246]), .B(n28194), .Z(n28197) );
  XOR U28133 ( .A(n28194), .B(p_input[230]), .Z(n28196) );
  XOR U28134 ( .A(n28198), .B(n28199), .Z(n28194) );
  AND U28135 ( .A(n28200), .B(n28201), .Z(n28199) );
  XNOR U28136 ( .A(p_input[245]), .B(n28198), .Z(n28201) );
  XOR U28137 ( .A(n28198), .B(p_input[229]), .Z(n28200) );
  XOR U28138 ( .A(n28202), .B(n28203), .Z(n28198) );
  AND U28139 ( .A(n28204), .B(n28205), .Z(n28203) );
  XNOR U28140 ( .A(p_input[244]), .B(n28202), .Z(n28205) );
  XOR U28141 ( .A(n28202), .B(p_input[228]), .Z(n28204) );
  XOR U28142 ( .A(n28206), .B(n28207), .Z(n28202) );
  AND U28143 ( .A(n28208), .B(n28209), .Z(n28207) );
  XNOR U28144 ( .A(p_input[243]), .B(n28206), .Z(n28209) );
  XOR U28145 ( .A(n28206), .B(p_input[227]), .Z(n28208) );
  XOR U28146 ( .A(n28210), .B(n28211), .Z(n28206) );
  AND U28147 ( .A(n28212), .B(n28213), .Z(n28211) );
  XNOR U28148 ( .A(p_input[242]), .B(n28210), .Z(n28213) );
  XOR U28149 ( .A(n28210), .B(p_input[226]), .Z(n28212) );
  XNOR U28150 ( .A(n28214), .B(n28215), .Z(n28210) );
  AND U28151 ( .A(n28216), .B(n28217), .Z(n28215) );
  XOR U28152 ( .A(p_input[241]), .B(n28214), .Z(n28217) );
  XNOR U28153 ( .A(p_input[225]), .B(n28214), .Z(n28216) );
  AND U28154 ( .A(p_input[240]), .B(n28218), .Z(n28214) );
  IV U28155 ( .A(p_input[224]), .Z(n28218) );
  XNOR U28156 ( .A(p_input[192]), .B(n28219), .Z(n28021) );
  AND U28157 ( .A(n1033), .B(n28220), .Z(n28219) );
  XOR U28158 ( .A(p_input[208]), .B(p_input[192]), .Z(n28220) );
  XOR U28159 ( .A(n28221), .B(n28222), .Z(n1033) );
  AND U28160 ( .A(n28223), .B(n28224), .Z(n28222) );
  XNOR U28161 ( .A(p_input[223]), .B(n28221), .Z(n28224) );
  XOR U28162 ( .A(n28221), .B(p_input[207]), .Z(n28223) );
  XOR U28163 ( .A(n28225), .B(n28226), .Z(n28221) );
  AND U28164 ( .A(n28227), .B(n28228), .Z(n28226) );
  XNOR U28165 ( .A(p_input[222]), .B(n28225), .Z(n28228) );
  XNOR U28166 ( .A(n28225), .B(n28035), .Z(n28227) );
  IV U28167 ( .A(p_input[206]), .Z(n28035) );
  XOR U28168 ( .A(n28229), .B(n28230), .Z(n28225) );
  AND U28169 ( .A(n28231), .B(n28232), .Z(n28230) );
  XNOR U28170 ( .A(p_input[221]), .B(n28229), .Z(n28232) );
  XNOR U28171 ( .A(n28229), .B(n28044), .Z(n28231) );
  IV U28172 ( .A(p_input[205]), .Z(n28044) );
  XOR U28173 ( .A(n28233), .B(n28234), .Z(n28229) );
  AND U28174 ( .A(n28235), .B(n28236), .Z(n28234) );
  XNOR U28175 ( .A(p_input[220]), .B(n28233), .Z(n28236) );
  XNOR U28176 ( .A(n28233), .B(n28053), .Z(n28235) );
  IV U28177 ( .A(p_input[204]), .Z(n28053) );
  XOR U28178 ( .A(n28237), .B(n28238), .Z(n28233) );
  AND U28179 ( .A(n28239), .B(n28240), .Z(n28238) );
  XNOR U28180 ( .A(p_input[219]), .B(n28237), .Z(n28240) );
  XNOR U28181 ( .A(n28237), .B(n28062), .Z(n28239) );
  IV U28182 ( .A(p_input[203]), .Z(n28062) );
  XOR U28183 ( .A(n28241), .B(n28242), .Z(n28237) );
  AND U28184 ( .A(n28243), .B(n28244), .Z(n28242) );
  XNOR U28185 ( .A(p_input[218]), .B(n28241), .Z(n28244) );
  XNOR U28186 ( .A(n28241), .B(n28071), .Z(n28243) );
  IV U28187 ( .A(p_input[202]), .Z(n28071) );
  XOR U28188 ( .A(n28245), .B(n28246), .Z(n28241) );
  AND U28189 ( .A(n28247), .B(n28248), .Z(n28246) );
  XNOR U28190 ( .A(p_input[217]), .B(n28245), .Z(n28248) );
  XNOR U28191 ( .A(n28245), .B(n28080), .Z(n28247) );
  IV U28192 ( .A(p_input[201]), .Z(n28080) );
  XOR U28193 ( .A(n28249), .B(n28250), .Z(n28245) );
  AND U28194 ( .A(n28251), .B(n28252), .Z(n28250) );
  XNOR U28195 ( .A(p_input[216]), .B(n28249), .Z(n28252) );
  XNOR U28196 ( .A(n28249), .B(n28089), .Z(n28251) );
  IV U28197 ( .A(p_input[200]), .Z(n28089) );
  XOR U28198 ( .A(n28253), .B(n28254), .Z(n28249) );
  AND U28199 ( .A(n28255), .B(n28256), .Z(n28254) );
  XNOR U28200 ( .A(p_input[215]), .B(n28253), .Z(n28256) );
  XNOR U28201 ( .A(n28253), .B(n28098), .Z(n28255) );
  IV U28202 ( .A(p_input[199]), .Z(n28098) );
  XOR U28203 ( .A(n28257), .B(n28258), .Z(n28253) );
  AND U28204 ( .A(n28259), .B(n28260), .Z(n28258) );
  XNOR U28205 ( .A(p_input[214]), .B(n28257), .Z(n28260) );
  XNOR U28206 ( .A(n28257), .B(n28107), .Z(n28259) );
  IV U28207 ( .A(p_input[198]), .Z(n28107) );
  XOR U28208 ( .A(n28261), .B(n28262), .Z(n28257) );
  AND U28209 ( .A(n28263), .B(n28264), .Z(n28262) );
  XNOR U28210 ( .A(p_input[213]), .B(n28261), .Z(n28264) );
  XNOR U28211 ( .A(n28261), .B(n28116), .Z(n28263) );
  IV U28212 ( .A(p_input[197]), .Z(n28116) );
  XOR U28213 ( .A(n28265), .B(n28266), .Z(n28261) );
  AND U28214 ( .A(n28267), .B(n28268), .Z(n28266) );
  XNOR U28215 ( .A(p_input[212]), .B(n28265), .Z(n28268) );
  XNOR U28216 ( .A(n28265), .B(n28125), .Z(n28267) );
  IV U28217 ( .A(p_input[196]), .Z(n28125) );
  XOR U28218 ( .A(n28269), .B(n28270), .Z(n28265) );
  AND U28219 ( .A(n28271), .B(n28272), .Z(n28270) );
  XNOR U28220 ( .A(p_input[211]), .B(n28269), .Z(n28272) );
  XNOR U28221 ( .A(n28269), .B(n28134), .Z(n28271) );
  IV U28222 ( .A(p_input[195]), .Z(n28134) );
  XOR U28223 ( .A(n28273), .B(n28274), .Z(n28269) );
  AND U28224 ( .A(n28275), .B(n28276), .Z(n28274) );
  XNOR U28225 ( .A(p_input[210]), .B(n28273), .Z(n28276) );
  XNOR U28226 ( .A(n28273), .B(n28143), .Z(n28275) );
  IV U28227 ( .A(p_input[194]), .Z(n28143) );
  XNOR U28228 ( .A(n28277), .B(n28278), .Z(n28273) );
  AND U28229 ( .A(n28279), .B(n28280), .Z(n28278) );
  XOR U28230 ( .A(p_input[209]), .B(n28277), .Z(n28280) );
  XNOR U28231 ( .A(p_input[193]), .B(n28277), .Z(n28279) );
  AND U28232 ( .A(p_input[208]), .B(n28281), .Z(n28277) );
  IV U28233 ( .A(p_input[192]), .Z(n28281) );
  XOR U28234 ( .A(n28282), .B(n28283), .Z(n27840) );
  AND U28235 ( .A(n581), .B(n28284), .Z(n28283) );
  XNOR U28236 ( .A(n28285), .B(n28282), .Z(n28284) );
  XOR U28237 ( .A(n28286), .B(n28287), .Z(n581) );
  AND U28238 ( .A(n28288), .B(n28289), .Z(n28287) );
  XNOR U28239 ( .A(n27850), .B(n28286), .Z(n28289) );
  AND U28240 ( .A(p_input[191]), .B(p_input[175]), .Z(n27850) );
  XOR U28241 ( .A(n28286), .B(n27851), .Z(n28288) );
  AND U28242 ( .A(p_input[159]), .B(p_input[143]), .Z(n27851) );
  XOR U28243 ( .A(n28290), .B(n28291), .Z(n28286) );
  AND U28244 ( .A(n28292), .B(n28293), .Z(n28291) );
  XOR U28245 ( .A(n28290), .B(n27863), .Z(n28293) );
  XNOR U28246 ( .A(p_input[174]), .B(n28294), .Z(n27863) );
  AND U28247 ( .A(n1039), .B(n28295), .Z(n28294) );
  XOR U28248 ( .A(p_input[190]), .B(p_input[174]), .Z(n28295) );
  XNOR U28249 ( .A(n27860), .B(n28290), .Z(n28292) );
  XOR U28250 ( .A(n28296), .B(n28297), .Z(n27860) );
  AND U28251 ( .A(n1036), .B(n28298), .Z(n28297) );
  XOR U28252 ( .A(p_input[158]), .B(p_input[142]), .Z(n28298) );
  XOR U28253 ( .A(n28299), .B(n28300), .Z(n28290) );
  AND U28254 ( .A(n28301), .B(n28302), .Z(n28300) );
  XOR U28255 ( .A(n28299), .B(n27875), .Z(n28302) );
  XNOR U28256 ( .A(p_input[173]), .B(n28303), .Z(n27875) );
  AND U28257 ( .A(n1039), .B(n28304), .Z(n28303) );
  XOR U28258 ( .A(p_input[189]), .B(p_input[173]), .Z(n28304) );
  XNOR U28259 ( .A(n27872), .B(n28299), .Z(n28301) );
  XOR U28260 ( .A(n28305), .B(n28306), .Z(n27872) );
  AND U28261 ( .A(n1036), .B(n28307), .Z(n28306) );
  XOR U28262 ( .A(p_input[157]), .B(p_input[141]), .Z(n28307) );
  XOR U28263 ( .A(n28308), .B(n28309), .Z(n28299) );
  AND U28264 ( .A(n28310), .B(n28311), .Z(n28309) );
  XOR U28265 ( .A(n28308), .B(n27887), .Z(n28311) );
  XNOR U28266 ( .A(p_input[172]), .B(n28312), .Z(n27887) );
  AND U28267 ( .A(n1039), .B(n28313), .Z(n28312) );
  XOR U28268 ( .A(p_input[188]), .B(p_input[172]), .Z(n28313) );
  XNOR U28269 ( .A(n27884), .B(n28308), .Z(n28310) );
  XOR U28270 ( .A(n28314), .B(n28315), .Z(n27884) );
  AND U28271 ( .A(n1036), .B(n28316), .Z(n28315) );
  XOR U28272 ( .A(p_input[156]), .B(p_input[140]), .Z(n28316) );
  XOR U28273 ( .A(n28317), .B(n28318), .Z(n28308) );
  AND U28274 ( .A(n28319), .B(n28320), .Z(n28318) );
  XOR U28275 ( .A(n28317), .B(n27899), .Z(n28320) );
  XNOR U28276 ( .A(p_input[171]), .B(n28321), .Z(n27899) );
  AND U28277 ( .A(n1039), .B(n28322), .Z(n28321) );
  XOR U28278 ( .A(p_input[187]), .B(p_input[171]), .Z(n28322) );
  XNOR U28279 ( .A(n27896), .B(n28317), .Z(n28319) );
  XOR U28280 ( .A(n28323), .B(n28324), .Z(n27896) );
  AND U28281 ( .A(n1036), .B(n28325), .Z(n28324) );
  XOR U28282 ( .A(p_input[155]), .B(p_input[139]), .Z(n28325) );
  XOR U28283 ( .A(n28326), .B(n28327), .Z(n28317) );
  AND U28284 ( .A(n28328), .B(n28329), .Z(n28327) );
  XOR U28285 ( .A(n28326), .B(n27911), .Z(n28329) );
  XNOR U28286 ( .A(p_input[170]), .B(n28330), .Z(n27911) );
  AND U28287 ( .A(n1039), .B(n28331), .Z(n28330) );
  XOR U28288 ( .A(p_input[186]), .B(p_input[170]), .Z(n28331) );
  XNOR U28289 ( .A(n27908), .B(n28326), .Z(n28328) );
  XOR U28290 ( .A(n28332), .B(n28333), .Z(n27908) );
  AND U28291 ( .A(n1036), .B(n28334), .Z(n28333) );
  XOR U28292 ( .A(p_input[154]), .B(p_input[138]), .Z(n28334) );
  XOR U28293 ( .A(n28335), .B(n28336), .Z(n28326) );
  AND U28294 ( .A(n28337), .B(n28338), .Z(n28336) );
  XOR U28295 ( .A(n28335), .B(n27923), .Z(n28338) );
  XNOR U28296 ( .A(p_input[169]), .B(n28339), .Z(n27923) );
  AND U28297 ( .A(n1039), .B(n28340), .Z(n28339) );
  XOR U28298 ( .A(p_input[185]), .B(p_input[169]), .Z(n28340) );
  XNOR U28299 ( .A(n27920), .B(n28335), .Z(n28337) );
  XOR U28300 ( .A(n28341), .B(n28342), .Z(n27920) );
  AND U28301 ( .A(n1036), .B(n28343), .Z(n28342) );
  XOR U28302 ( .A(p_input[153]), .B(p_input[137]), .Z(n28343) );
  XOR U28303 ( .A(n28344), .B(n28345), .Z(n28335) );
  AND U28304 ( .A(n28346), .B(n28347), .Z(n28345) );
  XOR U28305 ( .A(n28344), .B(n27935), .Z(n28347) );
  XNOR U28306 ( .A(p_input[168]), .B(n28348), .Z(n27935) );
  AND U28307 ( .A(n1039), .B(n28349), .Z(n28348) );
  XOR U28308 ( .A(p_input[184]), .B(p_input[168]), .Z(n28349) );
  XNOR U28309 ( .A(n27932), .B(n28344), .Z(n28346) );
  XOR U28310 ( .A(n28350), .B(n28351), .Z(n27932) );
  AND U28311 ( .A(n1036), .B(n28352), .Z(n28351) );
  XOR U28312 ( .A(p_input[152]), .B(p_input[136]), .Z(n28352) );
  XOR U28313 ( .A(n28353), .B(n28354), .Z(n28344) );
  AND U28314 ( .A(n28355), .B(n28356), .Z(n28354) );
  XOR U28315 ( .A(n28353), .B(n27947), .Z(n28356) );
  XNOR U28316 ( .A(p_input[167]), .B(n28357), .Z(n27947) );
  AND U28317 ( .A(n1039), .B(n28358), .Z(n28357) );
  XOR U28318 ( .A(p_input[183]), .B(p_input[167]), .Z(n28358) );
  XNOR U28319 ( .A(n27944), .B(n28353), .Z(n28355) );
  XOR U28320 ( .A(n28359), .B(n28360), .Z(n27944) );
  AND U28321 ( .A(n1036), .B(n28361), .Z(n28360) );
  XOR U28322 ( .A(p_input[151]), .B(p_input[135]), .Z(n28361) );
  XOR U28323 ( .A(n28362), .B(n28363), .Z(n28353) );
  AND U28324 ( .A(n28364), .B(n28365), .Z(n28363) );
  XOR U28325 ( .A(n28362), .B(n27959), .Z(n28365) );
  XNOR U28326 ( .A(p_input[166]), .B(n28366), .Z(n27959) );
  AND U28327 ( .A(n1039), .B(n28367), .Z(n28366) );
  XOR U28328 ( .A(p_input[182]), .B(p_input[166]), .Z(n28367) );
  XNOR U28329 ( .A(n27956), .B(n28362), .Z(n28364) );
  XOR U28330 ( .A(n28368), .B(n28369), .Z(n27956) );
  AND U28331 ( .A(n1036), .B(n28370), .Z(n28369) );
  XOR U28332 ( .A(p_input[150]), .B(p_input[134]), .Z(n28370) );
  XOR U28333 ( .A(n28371), .B(n28372), .Z(n28362) );
  AND U28334 ( .A(n28373), .B(n28374), .Z(n28372) );
  XOR U28335 ( .A(n28371), .B(n27971), .Z(n28374) );
  XNOR U28336 ( .A(p_input[165]), .B(n28375), .Z(n27971) );
  AND U28337 ( .A(n1039), .B(n28376), .Z(n28375) );
  XOR U28338 ( .A(p_input[181]), .B(p_input[165]), .Z(n28376) );
  XNOR U28339 ( .A(n27968), .B(n28371), .Z(n28373) );
  XOR U28340 ( .A(n28377), .B(n28378), .Z(n27968) );
  AND U28341 ( .A(n1036), .B(n28379), .Z(n28378) );
  XOR U28342 ( .A(p_input[149]), .B(p_input[133]), .Z(n28379) );
  XOR U28343 ( .A(n28380), .B(n28381), .Z(n28371) );
  AND U28344 ( .A(n28382), .B(n28383), .Z(n28381) );
  XOR U28345 ( .A(n28380), .B(n27983), .Z(n28383) );
  XNOR U28346 ( .A(p_input[164]), .B(n28384), .Z(n27983) );
  AND U28347 ( .A(n1039), .B(n28385), .Z(n28384) );
  XOR U28348 ( .A(p_input[180]), .B(p_input[164]), .Z(n28385) );
  XNOR U28349 ( .A(n27980), .B(n28380), .Z(n28382) );
  XOR U28350 ( .A(n28386), .B(n28387), .Z(n27980) );
  AND U28351 ( .A(n1036), .B(n28388), .Z(n28387) );
  XOR U28352 ( .A(p_input[148]), .B(p_input[132]), .Z(n28388) );
  XOR U28353 ( .A(n28389), .B(n28390), .Z(n28380) );
  AND U28354 ( .A(n28391), .B(n28392), .Z(n28390) );
  XOR U28355 ( .A(n28389), .B(n27995), .Z(n28392) );
  XNOR U28356 ( .A(p_input[163]), .B(n28393), .Z(n27995) );
  AND U28357 ( .A(n1039), .B(n28394), .Z(n28393) );
  XOR U28358 ( .A(p_input[179]), .B(p_input[163]), .Z(n28394) );
  XNOR U28359 ( .A(n27992), .B(n28389), .Z(n28391) );
  XOR U28360 ( .A(n28395), .B(n28396), .Z(n27992) );
  AND U28361 ( .A(n1036), .B(n28397), .Z(n28396) );
  XOR U28362 ( .A(p_input[147]), .B(p_input[131]), .Z(n28397) );
  XOR U28363 ( .A(n28398), .B(n28399), .Z(n28389) );
  AND U28364 ( .A(n28400), .B(n28401), .Z(n28399) );
  XOR U28365 ( .A(n28398), .B(n28007), .Z(n28401) );
  XNOR U28366 ( .A(p_input[162]), .B(n28402), .Z(n28007) );
  AND U28367 ( .A(n1039), .B(n28403), .Z(n28402) );
  XOR U28368 ( .A(p_input[178]), .B(p_input[162]), .Z(n28403) );
  XNOR U28369 ( .A(n28004), .B(n28398), .Z(n28400) );
  XOR U28370 ( .A(n28404), .B(n28405), .Z(n28004) );
  AND U28371 ( .A(n1036), .B(n28406), .Z(n28405) );
  XOR U28372 ( .A(p_input[146]), .B(p_input[130]), .Z(n28406) );
  XOR U28373 ( .A(n28407), .B(n28408), .Z(n28398) );
  AND U28374 ( .A(n28409), .B(n28410), .Z(n28408) );
  XNOR U28375 ( .A(n28411), .B(n28020), .Z(n28410) );
  XNOR U28376 ( .A(p_input[161]), .B(n28412), .Z(n28020) );
  AND U28377 ( .A(n1039), .B(n28413), .Z(n28412) );
  XNOR U28378 ( .A(p_input[177]), .B(n28414), .Z(n28413) );
  IV U28379 ( .A(p_input[161]), .Z(n28414) );
  XNOR U28380 ( .A(n28017), .B(n28407), .Z(n28409) );
  XNOR U28381 ( .A(p_input[129]), .B(n28415), .Z(n28017) );
  AND U28382 ( .A(n1036), .B(n28416), .Z(n28415) );
  XOR U28383 ( .A(p_input[145]), .B(p_input[129]), .Z(n28416) );
  IV U28384 ( .A(n28411), .Z(n28407) );
  AND U28385 ( .A(n28282), .B(n28285), .Z(n28411) );
  XOR U28386 ( .A(p_input[160]), .B(n28417), .Z(n28285) );
  AND U28387 ( .A(n1039), .B(n28418), .Z(n28417) );
  XOR U28388 ( .A(p_input[176]), .B(p_input[160]), .Z(n28418) );
  XOR U28389 ( .A(n28419), .B(n28420), .Z(n1039) );
  AND U28390 ( .A(n28421), .B(n28422), .Z(n28420) );
  XNOR U28391 ( .A(p_input[191]), .B(n28419), .Z(n28422) );
  XOR U28392 ( .A(n28419), .B(p_input[175]), .Z(n28421) );
  XOR U28393 ( .A(n28423), .B(n28424), .Z(n28419) );
  AND U28394 ( .A(n28425), .B(n28426), .Z(n28424) );
  XNOR U28395 ( .A(p_input[190]), .B(n28423), .Z(n28426) );
  XOR U28396 ( .A(n28423), .B(p_input[174]), .Z(n28425) );
  XOR U28397 ( .A(n28427), .B(n28428), .Z(n28423) );
  AND U28398 ( .A(n28429), .B(n28430), .Z(n28428) );
  XNOR U28399 ( .A(p_input[189]), .B(n28427), .Z(n28430) );
  XOR U28400 ( .A(n28427), .B(p_input[173]), .Z(n28429) );
  XOR U28401 ( .A(n28431), .B(n28432), .Z(n28427) );
  AND U28402 ( .A(n28433), .B(n28434), .Z(n28432) );
  XNOR U28403 ( .A(p_input[188]), .B(n28431), .Z(n28434) );
  XOR U28404 ( .A(n28431), .B(p_input[172]), .Z(n28433) );
  XOR U28405 ( .A(n28435), .B(n28436), .Z(n28431) );
  AND U28406 ( .A(n28437), .B(n28438), .Z(n28436) );
  XNOR U28407 ( .A(p_input[187]), .B(n28435), .Z(n28438) );
  XOR U28408 ( .A(n28435), .B(p_input[171]), .Z(n28437) );
  XOR U28409 ( .A(n28439), .B(n28440), .Z(n28435) );
  AND U28410 ( .A(n28441), .B(n28442), .Z(n28440) );
  XNOR U28411 ( .A(p_input[186]), .B(n28439), .Z(n28442) );
  XOR U28412 ( .A(n28439), .B(p_input[170]), .Z(n28441) );
  XOR U28413 ( .A(n28443), .B(n28444), .Z(n28439) );
  AND U28414 ( .A(n28445), .B(n28446), .Z(n28444) );
  XNOR U28415 ( .A(p_input[185]), .B(n28443), .Z(n28446) );
  XOR U28416 ( .A(n28443), .B(p_input[169]), .Z(n28445) );
  XOR U28417 ( .A(n28447), .B(n28448), .Z(n28443) );
  AND U28418 ( .A(n28449), .B(n28450), .Z(n28448) );
  XNOR U28419 ( .A(p_input[184]), .B(n28447), .Z(n28450) );
  XOR U28420 ( .A(n28447), .B(p_input[168]), .Z(n28449) );
  XOR U28421 ( .A(n28451), .B(n28452), .Z(n28447) );
  AND U28422 ( .A(n28453), .B(n28454), .Z(n28452) );
  XNOR U28423 ( .A(p_input[183]), .B(n28451), .Z(n28454) );
  XOR U28424 ( .A(n28451), .B(p_input[167]), .Z(n28453) );
  XOR U28425 ( .A(n28455), .B(n28456), .Z(n28451) );
  AND U28426 ( .A(n28457), .B(n28458), .Z(n28456) );
  XNOR U28427 ( .A(p_input[182]), .B(n28455), .Z(n28458) );
  XOR U28428 ( .A(n28455), .B(p_input[166]), .Z(n28457) );
  XOR U28429 ( .A(n28459), .B(n28460), .Z(n28455) );
  AND U28430 ( .A(n28461), .B(n28462), .Z(n28460) );
  XNOR U28431 ( .A(p_input[181]), .B(n28459), .Z(n28462) );
  XOR U28432 ( .A(n28459), .B(p_input[165]), .Z(n28461) );
  XOR U28433 ( .A(n28463), .B(n28464), .Z(n28459) );
  AND U28434 ( .A(n28465), .B(n28466), .Z(n28464) );
  XNOR U28435 ( .A(p_input[180]), .B(n28463), .Z(n28466) );
  XOR U28436 ( .A(n28463), .B(p_input[164]), .Z(n28465) );
  XOR U28437 ( .A(n28467), .B(n28468), .Z(n28463) );
  AND U28438 ( .A(n28469), .B(n28470), .Z(n28468) );
  XNOR U28439 ( .A(p_input[179]), .B(n28467), .Z(n28470) );
  XOR U28440 ( .A(n28467), .B(p_input[163]), .Z(n28469) );
  XOR U28441 ( .A(n28471), .B(n28472), .Z(n28467) );
  AND U28442 ( .A(n28473), .B(n28474), .Z(n28472) );
  XNOR U28443 ( .A(p_input[178]), .B(n28471), .Z(n28474) );
  XOR U28444 ( .A(n28471), .B(p_input[162]), .Z(n28473) );
  XNOR U28445 ( .A(n28475), .B(n28476), .Z(n28471) );
  AND U28446 ( .A(n28477), .B(n28478), .Z(n28476) );
  XOR U28447 ( .A(p_input[177]), .B(n28475), .Z(n28478) );
  XNOR U28448 ( .A(p_input[161]), .B(n28475), .Z(n28477) );
  AND U28449 ( .A(p_input[176]), .B(n28479), .Z(n28475) );
  IV U28450 ( .A(p_input[160]), .Z(n28479) );
  XNOR U28451 ( .A(p_input[128]), .B(n28480), .Z(n28282) );
  AND U28452 ( .A(n1036), .B(n28481), .Z(n28480) );
  XOR U28453 ( .A(p_input[144]), .B(p_input[128]), .Z(n28481) );
  XOR U28454 ( .A(n28482), .B(n28483), .Z(n1036) );
  AND U28455 ( .A(n28484), .B(n28485), .Z(n28483) );
  XNOR U28456 ( .A(p_input[159]), .B(n28482), .Z(n28485) );
  XOR U28457 ( .A(n28482), .B(p_input[143]), .Z(n28484) );
  XOR U28458 ( .A(n28486), .B(n28487), .Z(n28482) );
  AND U28459 ( .A(n28488), .B(n28489), .Z(n28487) );
  XNOR U28460 ( .A(p_input[158]), .B(n28486), .Z(n28489) );
  XNOR U28461 ( .A(n28486), .B(n28296), .Z(n28488) );
  IV U28462 ( .A(p_input[142]), .Z(n28296) );
  XOR U28463 ( .A(n28490), .B(n28491), .Z(n28486) );
  AND U28464 ( .A(n28492), .B(n28493), .Z(n28491) );
  XNOR U28465 ( .A(p_input[157]), .B(n28490), .Z(n28493) );
  XNOR U28466 ( .A(n28490), .B(n28305), .Z(n28492) );
  IV U28467 ( .A(p_input[141]), .Z(n28305) );
  XOR U28468 ( .A(n28494), .B(n28495), .Z(n28490) );
  AND U28469 ( .A(n28496), .B(n28497), .Z(n28495) );
  XNOR U28470 ( .A(p_input[156]), .B(n28494), .Z(n28497) );
  XNOR U28471 ( .A(n28494), .B(n28314), .Z(n28496) );
  IV U28472 ( .A(p_input[140]), .Z(n28314) );
  XOR U28473 ( .A(n28498), .B(n28499), .Z(n28494) );
  AND U28474 ( .A(n28500), .B(n28501), .Z(n28499) );
  XNOR U28475 ( .A(p_input[155]), .B(n28498), .Z(n28501) );
  XNOR U28476 ( .A(n28498), .B(n28323), .Z(n28500) );
  IV U28477 ( .A(p_input[139]), .Z(n28323) );
  XOR U28478 ( .A(n28502), .B(n28503), .Z(n28498) );
  AND U28479 ( .A(n28504), .B(n28505), .Z(n28503) );
  XNOR U28480 ( .A(p_input[154]), .B(n28502), .Z(n28505) );
  XNOR U28481 ( .A(n28502), .B(n28332), .Z(n28504) );
  IV U28482 ( .A(p_input[138]), .Z(n28332) );
  XOR U28483 ( .A(n28506), .B(n28507), .Z(n28502) );
  AND U28484 ( .A(n28508), .B(n28509), .Z(n28507) );
  XNOR U28485 ( .A(p_input[153]), .B(n28506), .Z(n28509) );
  XNOR U28486 ( .A(n28506), .B(n28341), .Z(n28508) );
  IV U28487 ( .A(p_input[137]), .Z(n28341) );
  XOR U28488 ( .A(n28510), .B(n28511), .Z(n28506) );
  AND U28489 ( .A(n28512), .B(n28513), .Z(n28511) );
  XNOR U28490 ( .A(p_input[152]), .B(n28510), .Z(n28513) );
  XNOR U28491 ( .A(n28510), .B(n28350), .Z(n28512) );
  IV U28492 ( .A(p_input[136]), .Z(n28350) );
  XOR U28493 ( .A(n28514), .B(n28515), .Z(n28510) );
  AND U28494 ( .A(n28516), .B(n28517), .Z(n28515) );
  XNOR U28495 ( .A(p_input[151]), .B(n28514), .Z(n28517) );
  XNOR U28496 ( .A(n28514), .B(n28359), .Z(n28516) );
  IV U28497 ( .A(p_input[135]), .Z(n28359) );
  XOR U28498 ( .A(n28518), .B(n28519), .Z(n28514) );
  AND U28499 ( .A(n28520), .B(n28521), .Z(n28519) );
  XNOR U28500 ( .A(p_input[150]), .B(n28518), .Z(n28521) );
  XNOR U28501 ( .A(n28518), .B(n28368), .Z(n28520) );
  IV U28502 ( .A(p_input[134]), .Z(n28368) );
  XOR U28503 ( .A(n28522), .B(n28523), .Z(n28518) );
  AND U28504 ( .A(n28524), .B(n28525), .Z(n28523) );
  XNOR U28505 ( .A(p_input[149]), .B(n28522), .Z(n28525) );
  XNOR U28506 ( .A(n28522), .B(n28377), .Z(n28524) );
  IV U28507 ( .A(p_input[133]), .Z(n28377) );
  XOR U28508 ( .A(n28526), .B(n28527), .Z(n28522) );
  AND U28509 ( .A(n28528), .B(n28529), .Z(n28527) );
  XNOR U28510 ( .A(p_input[148]), .B(n28526), .Z(n28529) );
  XNOR U28511 ( .A(n28526), .B(n28386), .Z(n28528) );
  IV U28512 ( .A(p_input[132]), .Z(n28386) );
  XOR U28513 ( .A(n28530), .B(n28531), .Z(n28526) );
  AND U28514 ( .A(n28532), .B(n28533), .Z(n28531) );
  XNOR U28515 ( .A(p_input[147]), .B(n28530), .Z(n28533) );
  XNOR U28516 ( .A(n28530), .B(n28395), .Z(n28532) );
  IV U28517 ( .A(p_input[131]), .Z(n28395) );
  XOR U28518 ( .A(n28534), .B(n28535), .Z(n28530) );
  AND U28519 ( .A(n28536), .B(n28537), .Z(n28535) );
  XNOR U28520 ( .A(p_input[146]), .B(n28534), .Z(n28537) );
  XNOR U28521 ( .A(n28534), .B(n28404), .Z(n28536) );
  IV U28522 ( .A(p_input[130]), .Z(n28404) );
  XNOR U28523 ( .A(n28538), .B(n28539), .Z(n28534) );
  AND U28524 ( .A(n28540), .B(n28541), .Z(n28539) );
  XOR U28525 ( .A(p_input[145]), .B(n28538), .Z(n28541) );
  XNOR U28526 ( .A(p_input[129]), .B(n28538), .Z(n28540) );
  AND U28527 ( .A(p_input[144]), .B(n28542), .Z(n28538) );
  IV U28528 ( .A(p_input[128]), .Z(n28542) );
  XOR U28529 ( .A(n28543), .B(n28544), .Z(n27658) );
  AND U28530 ( .A(n836), .B(n28545), .Z(n28544) );
  XNOR U28531 ( .A(n28546), .B(n28543), .Z(n28545) );
  XOR U28532 ( .A(n28547), .B(n28548), .Z(n836) );
  AND U28533 ( .A(n28549), .B(n28550), .Z(n28548) );
  XNOR U28534 ( .A(n27670), .B(n28547), .Z(n28550) );
  AND U28535 ( .A(n28551), .B(n28552), .Z(n27670) );
  XOR U28536 ( .A(n28547), .B(n27669), .Z(n28549) );
  AND U28537 ( .A(n28553), .B(n28554), .Z(n27669) );
  XOR U28538 ( .A(n28555), .B(n28556), .Z(n28547) );
  AND U28539 ( .A(n28557), .B(n28558), .Z(n28556) );
  XOR U28540 ( .A(n28555), .B(n27682), .Z(n28558) );
  XOR U28541 ( .A(n28559), .B(n28560), .Z(n27682) );
  AND U28542 ( .A(n587), .B(n28561), .Z(n28560) );
  XOR U28543 ( .A(n28562), .B(n28559), .Z(n28561) );
  XNOR U28544 ( .A(n27679), .B(n28555), .Z(n28557) );
  XOR U28545 ( .A(n28563), .B(n28564), .Z(n27679) );
  AND U28546 ( .A(n584), .B(n28565), .Z(n28564) );
  XOR U28547 ( .A(n28566), .B(n28563), .Z(n28565) );
  XOR U28548 ( .A(n28567), .B(n28568), .Z(n28555) );
  AND U28549 ( .A(n28569), .B(n28570), .Z(n28568) );
  XOR U28550 ( .A(n28567), .B(n27694), .Z(n28570) );
  XOR U28551 ( .A(n28571), .B(n28572), .Z(n27694) );
  AND U28552 ( .A(n587), .B(n28573), .Z(n28572) );
  XOR U28553 ( .A(n28574), .B(n28571), .Z(n28573) );
  XNOR U28554 ( .A(n27691), .B(n28567), .Z(n28569) );
  XOR U28555 ( .A(n28575), .B(n28576), .Z(n27691) );
  AND U28556 ( .A(n584), .B(n28577), .Z(n28576) );
  XOR U28557 ( .A(n28578), .B(n28575), .Z(n28577) );
  XOR U28558 ( .A(n28579), .B(n28580), .Z(n28567) );
  AND U28559 ( .A(n28581), .B(n28582), .Z(n28580) );
  XOR U28560 ( .A(n28579), .B(n27706), .Z(n28582) );
  XOR U28561 ( .A(n28583), .B(n28584), .Z(n27706) );
  AND U28562 ( .A(n587), .B(n28585), .Z(n28584) );
  XOR U28563 ( .A(n28586), .B(n28583), .Z(n28585) );
  XNOR U28564 ( .A(n27703), .B(n28579), .Z(n28581) );
  XOR U28565 ( .A(n28587), .B(n28588), .Z(n27703) );
  AND U28566 ( .A(n584), .B(n28589), .Z(n28588) );
  XOR U28567 ( .A(n28590), .B(n28587), .Z(n28589) );
  XOR U28568 ( .A(n28591), .B(n28592), .Z(n28579) );
  AND U28569 ( .A(n28593), .B(n28594), .Z(n28592) );
  XOR U28570 ( .A(n28591), .B(n27718), .Z(n28594) );
  XOR U28571 ( .A(n28595), .B(n28596), .Z(n27718) );
  AND U28572 ( .A(n587), .B(n28597), .Z(n28596) );
  XOR U28573 ( .A(n28598), .B(n28595), .Z(n28597) );
  XNOR U28574 ( .A(n27715), .B(n28591), .Z(n28593) );
  XOR U28575 ( .A(n28599), .B(n28600), .Z(n27715) );
  AND U28576 ( .A(n584), .B(n28601), .Z(n28600) );
  XOR U28577 ( .A(n28602), .B(n28599), .Z(n28601) );
  XOR U28578 ( .A(n28603), .B(n28604), .Z(n28591) );
  AND U28579 ( .A(n28605), .B(n28606), .Z(n28604) );
  XOR U28580 ( .A(n28603), .B(n27730), .Z(n28606) );
  XOR U28581 ( .A(n28607), .B(n28608), .Z(n27730) );
  AND U28582 ( .A(n587), .B(n28609), .Z(n28608) );
  XOR U28583 ( .A(n28610), .B(n28607), .Z(n28609) );
  XNOR U28584 ( .A(n27727), .B(n28603), .Z(n28605) );
  XOR U28585 ( .A(n28611), .B(n28612), .Z(n27727) );
  AND U28586 ( .A(n584), .B(n28613), .Z(n28612) );
  XOR U28587 ( .A(n28614), .B(n28611), .Z(n28613) );
  XOR U28588 ( .A(n28615), .B(n28616), .Z(n28603) );
  AND U28589 ( .A(n28617), .B(n28618), .Z(n28616) );
  XOR U28590 ( .A(n28615), .B(n27742), .Z(n28618) );
  XOR U28591 ( .A(n28619), .B(n28620), .Z(n27742) );
  AND U28592 ( .A(n587), .B(n28621), .Z(n28620) );
  XOR U28593 ( .A(n28622), .B(n28619), .Z(n28621) );
  XNOR U28594 ( .A(n27739), .B(n28615), .Z(n28617) );
  XOR U28595 ( .A(n28623), .B(n28624), .Z(n27739) );
  AND U28596 ( .A(n584), .B(n28625), .Z(n28624) );
  XOR U28597 ( .A(n28626), .B(n28623), .Z(n28625) );
  XOR U28598 ( .A(n28627), .B(n28628), .Z(n28615) );
  AND U28599 ( .A(n28629), .B(n28630), .Z(n28628) );
  XOR U28600 ( .A(n28627), .B(n27754), .Z(n28630) );
  XOR U28601 ( .A(n28631), .B(n28632), .Z(n27754) );
  AND U28602 ( .A(n587), .B(n28633), .Z(n28632) );
  XOR U28603 ( .A(n28634), .B(n28631), .Z(n28633) );
  XNOR U28604 ( .A(n27751), .B(n28627), .Z(n28629) );
  XOR U28605 ( .A(n28635), .B(n28636), .Z(n27751) );
  AND U28606 ( .A(n584), .B(n28637), .Z(n28636) );
  XOR U28607 ( .A(n28638), .B(n28635), .Z(n28637) );
  XOR U28608 ( .A(n28639), .B(n28640), .Z(n28627) );
  AND U28609 ( .A(n28641), .B(n28642), .Z(n28640) );
  XOR U28610 ( .A(n28639), .B(n27766), .Z(n28642) );
  XOR U28611 ( .A(n28643), .B(n28644), .Z(n27766) );
  AND U28612 ( .A(n587), .B(n28645), .Z(n28644) );
  XOR U28613 ( .A(n28646), .B(n28643), .Z(n28645) );
  XNOR U28614 ( .A(n27763), .B(n28639), .Z(n28641) );
  XOR U28615 ( .A(n28647), .B(n28648), .Z(n27763) );
  AND U28616 ( .A(n584), .B(n28649), .Z(n28648) );
  XOR U28617 ( .A(n28650), .B(n28647), .Z(n28649) );
  XOR U28618 ( .A(n28651), .B(n28652), .Z(n28639) );
  AND U28619 ( .A(n28653), .B(n28654), .Z(n28652) );
  XOR U28620 ( .A(n28651), .B(n27778), .Z(n28654) );
  XOR U28621 ( .A(n28655), .B(n28656), .Z(n27778) );
  AND U28622 ( .A(n587), .B(n28657), .Z(n28656) );
  XOR U28623 ( .A(n28658), .B(n28655), .Z(n28657) );
  XNOR U28624 ( .A(n27775), .B(n28651), .Z(n28653) );
  XOR U28625 ( .A(n28659), .B(n28660), .Z(n27775) );
  AND U28626 ( .A(n584), .B(n28661), .Z(n28660) );
  XOR U28627 ( .A(n28662), .B(n28659), .Z(n28661) );
  XOR U28628 ( .A(n28663), .B(n28664), .Z(n28651) );
  AND U28629 ( .A(n28665), .B(n28666), .Z(n28664) );
  XOR U28630 ( .A(n28663), .B(n27790), .Z(n28666) );
  XOR U28631 ( .A(n28667), .B(n28668), .Z(n27790) );
  AND U28632 ( .A(n587), .B(n28669), .Z(n28668) );
  XOR U28633 ( .A(n28670), .B(n28667), .Z(n28669) );
  XNOR U28634 ( .A(n27787), .B(n28663), .Z(n28665) );
  XOR U28635 ( .A(n28671), .B(n28672), .Z(n27787) );
  AND U28636 ( .A(n584), .B(n28673), .Z(n28672) );
  XOR U28637 ( .A(n28674), .B(n28671), .Z(n28673) );
  XOR U28638 ( .A(n28675), .B(n28676), .Z(n28663) );
  AND U28639 ( .A(n28677), .B(n28678), .Z(n28676) );
  XOR U28640 ( .A(n28675), .B(n27802), .Z(n28678) );
  XOR U28641 ( .A(n28679), .B(n28680), .Z(n27802) );
  AND U28642 ( .A(n587), .B(n28681), .Z(n28680) );
  XOR U28643 ( .A(n28682), .B(n28679), .Z(n28681) );
  XNOR U28644 ( .A(n27799), .B(n28675), .Z(n28677) );
  XOR U28645 ( .A(n28683), .B(n28684), .Z(n27799) );
  AND U28646 ( .A(n584), .B(n28685), .Z(n28684) );
  XOR U28647 ( .A(n28686), .B(n28683), .Z(n28685) );
  XOR U28648 ( .A(n28687), .B(n28688), .Z(n28675) );
  AND U28649 ( .A(n28689), .B(n28690), .Z(n28688) );
  XOR U28650 ( .A(n28687), .B(n27814), .Z(n28690) );
  XOR U28651 ( .A(n28691), .B(n28692), .Z(n27814) );
  AND U28652 ( .A(n587), .B(n28693), .Z(n28692) );
  XOR U28653 ( .A(n28694), .B(n28691), .Z(n28693) );
  XNOR U28654 ( .A(n27811), .B(n28687), .Z(n28689) );
  XOR U28655 ( .A(n28695), .B(n28696), .Z(n27811) );
  AND U28656 ( .A(n584), .B(n28697), .Z(n28696) );
  XOR U28657 ( .A(n28698), .B(n28695), .Z(n28697) );
  XOR U28658 ( .A(n28699), .B(n28700), .Z(n28687) );
  AND U28659 ( .A(n28701), .B(n28702), .Z(n28700) );
  XOR U28660 ( .A(n28699), .B(n27826), .Z(n28702) );
  XOR U28661 ( .A(n28703), .B(n28704), .Z(n27826) );
  AND U28662 ( .A(n587), .B(n28705), .Z(n28704) );
  XOR U28663 ( .A(n28706), .B(n28703), .Z(n28705) );
  XNOR U28664 ( .A(n27823), .B(n28699), .Z(n28701) );
  XOR U28665 ( .A(n28707), .B(n28708), .Z(n27823) );
  AND U28666 ( .A(n584), .B(n28709), .Z(n28708) );
  XOR U28667 ( .A(n28710), .B(n28707), .Z(n28709) );
  XOR U28668 ( .A(n28711), .B(n28712), .Z(n28699) );
  AND U28669 ( .A(n28713), .B(n28714), .Z(n28712) );
  XNOR U28670 ( .A(n28715), .B(n27839), .Z(n28714) );
  XOR U28671 ( .A(n28716), .B(n28717), .Z(n27839) );
  AND U28672 ( .A(n587), .B(n28718), .Z(n28717) );
  XOR U28673 ( .A(n28716), .B(n28719), .Z(n28718) );
  XNOR U28674 ( .A(n27836), .B(n28711), .Z(n28713) );
  XOR U28675 ( .A(n28720), .B(n28721), .Z(n27836) );
  AND U28676 ( .A(n584), .B(n28722), .Z(n28721) );
  XOR U28677 ( .A(n28720), .B(n28723), .Z(n28722) );
  IV U28678 ( .A(n28715), .Z(n28711) );
  AND U28679 ( .A(n28543), .B(n28546), .Z(n28715) );
  XNOR U28680 ( .A(n28724), .B(n28725), .Z(n28546) );
  AND U28681 ( .A(n587), .B(n28726), .Z(n28725) );
  XNOR U28682 ( .A(n28727), .B(n28724), .Z(n28726) );
  XOR U28683 ( .A(n28728), .B(n28729), .Z(n587) );
  AND U28684 ( .A(n28730), .B(n28731), .Z(n28729) );
  XNOR U28685 ( .A(n28551), .B(n28728), .Z(n28731) );
  AND U28686 ( .A(p_input[127]), .B(p_input[111]), .Z(n28551) );
  XOR U28687 ( .A(n28728), .B(n28552), .Z(n28730) );
  AND U28688 ( .A(p_input[95]), .B(p_input[79]), .Z(n28552) );
  XOR U28689 ( .A(n28732), .B(n28733), .Z(n28728) );
  AND U28690 ( .A(n28734), .B(n28735), .Z(n28733) );
  XOR U28691 ( .A(n28732), .B(n28562), .Z(n28735) );
  XNOR U28692 ( .A(p_input[110]), .B(n28736), .Z(n28562) );
  AND U28693 ( .A(n1059), .B(n28737), .Z(n28736) );
  XOR U28694 ( .A(p_input[126]), .B(p_input[110]), .Z(n28737) );
  XNOR U28695 ( .A(n28559), .B(n28732), .Z(n28734) );
  XOR U28696 ( .A(n28738), .B(n28739), .Z(n28559) );
  AND U28697 ( .A(n1057), .B(n28740), .Z(n28739) );
  XOR U28698 ( .A(p_input[94]), .B(p_input[78]), .Z(n28740) );
  XOR U28699 ( .A(n28741), .B(n28742), .Z(n28732) );
  AND U28700 ( .A(n28743), .B(n28744), .Z(n28742) );
  XOR U28701 ( .A(n28741), .B(n28574), .Z(n28744) );
  XNOR U28702 ( .A(p_input[109]), .B(n28745), .Z(n28574) );
  AND U28703 ( .A(n1059), .B(n28746), .Z(n28745) );
  XOR U28704 ( .A(p_input[125]), .B(p_input[109]), .Z(n28746) );
  XNOR U28705 ( .A(n28571), .B(n28741), .Z(n28743) );
  XOR U28706 ( .A(n28747), .B(n28748), .Z(n28571) );
  AND U28707 ( .A(n1057), .B(n28749), .Z(n28748) );
  XOR U28708 ( .A(p_input[93]), .B(p_input[77]), .Z(n28749) );
  XOR U28709 ( .A(n28750), .B(n28751), .Z(n28741) );
  AND U28710 ( .A(n28752), .B(n28753), .Z(n28751) );
  XOR U28711 ( .A(n28750), .B(n28586), .Z(n28753) );
  XNOR U28712 ( .A(p_input[108]), .B(n28754), .Z(n28586) );
  AND U28713 ( .A(n1059), .B(n28755), .Z(n28754) );
  XOR U28714 ( .A(p_input[124]), .B(p_input[108]), .Z(n28755) );
  XNOR U28715 ( .A(n28583), .B(n28750), .Z(n28752) );
  XOR U28716 ( .A(n28756), .B(n28757), .Z(n28583) );
  AND U28717 ( .A(n1057), .B(n28758), .Z(n28757) );
  XOR U28718 ( .A(p_input[92]), .B(p_input[76]), .Z(n28758) );
  XOR U28719 ( .A(n28759), .B(n28760), .Z(n28750) );
  AND U28720 ( .A(n28761), .B(n28762), .Z(n28760) );
  XOR U28721 ( .A(n28759), .B(n28598), .Z(n28762) );
  XNOR U28722 ( .A(p_input[107]), .B(n28763), .Z(n28598) );
  AND U28723 ( .A(n1059), .B(n28764), .Z(n28763) );
  XOR U28724 ( .A(p_input[123]), .B(p_input[107]), .Z(n28764) );
  XNOR U28725 ( .A(n28595), .B(n28759), .Z(n28761) );
  XOR U28726 ( .A(n28765), .B(n28766), .Z(n28595) );
  AND U28727 ( .A(n1057), .B(n28767), .Z(n28766) );
  XOR U28728 ( .A(p_input[91]), .B(p_input[75]), .Z(n28767) );
  XOR U28729 ( .A(n28768), .B(n28769), .Z(n28759) );
  AND U28730 ( .A(n28770), .B(n28771), .Z(n28769) );
  XOR U28731 ( .A(n28768), .B(n28610), .Z(n28771) );
  XNOR U28732 ( .A(p_input[106]), .B(n28772), .Z(n28610) );
  AND U28733 ( .A(n1059), .B(n28773), .Z(n28772) );
  XOR U28734 ( .A(p_input[122]), .B(p_input[106]), .Z(n28773) );
  XNOR U28735 ( .A(n28607), .B(n28768), .Z(n28770) );
  XOR U28736 ( .A(n28774), .B(n28775), .Z(n28607) );
  AND U28737 ( .A(n1057), .B(n28776), .Z(n28775) );
  XOR U28738 ( .A(p_input[90]), .B(p_input[74]), .Z(n28776) );
  XOR U28739 ( .A(n28777), .B(n28778), .Z(n28768) );
  AND U28740 ( .A(n28779), .B(n28780), .Z(n28778) );
  XOR U28741 ( .A(n28777), .B(n28622), .Z(n28780) );
  XNOR U28742 ( .A(p_input[105]), .B(n28781), .Z(n28622) );
  AND U28743 ( .A(n1059), .B(n28782), .Z(n28781) );
  XOR U28744 ( .A(p_input[121]), .B(p_input[105]), .Z(n28782) );
  XNOR U28745 ( .A(n28619), .B(n28777), .Z(n28779) );
  XOR U28746 ( .A(n28783), .B(n28784), .Z(n28619) );
  AND U28747 ( .A(n1057), .B(n28785), .Z(n28784) );
  XOR U28748 ( .A(p_input[89]), .B(p_input[73]), .Z(n28785) );
  XOR U28749 ( .A(n28786), .B(n28787), .Z(n28777) );
  AND U28750 ( .A(n28788), .B(n28789), .Z(n28787) );
  XOR U28751 ( .A(n28786), .B(n28634), .Z(n28789) );
  XNOR U28752 ( .A(p_input[104]), .B(n28790), .Z(n28634) );
  AND U28753 ( .A(n1059), .B(n28791), .Z(n28790) );
  XOR U28754 ( .A(p_input[120]), .B(p_input[104]), .Z(n28791) );
  XNOR U28755 ( .A(n28631), .B(n28786), .Z(n28788) );
  XOR U28756 ( .A(n28792), .B(n28793), .Z(n28631) );
  AND U28757 ( .A(n1057), .B(n28794), .Z(n28793) );
  XOR U28758 ( .A(p_input[88]), .B(p_input[72]), .Z(n28794) );
  XOR U28759 ( .A(n28795), .B(n28796), .Z(n28786) );
  AND U28760 ( .A(n28797), .B(n28798), .Z(n28796) );
  XOR U28761 ( .A(n28795), .B(n28646), .Z(n28798) );
  XNOR U28762 ( .A(p_input[103]), .B(n28799), .Z(n28646) );
  AND U28763 ( .A(n1059), .B(n28800), .Z(n28799) );
  XOR U28764 ( .A(p_input[119]), .B(p_input[103]), .Z(n28800) );
  XNOR U28765 ( .A(n28643), .B(n28795), .Z(n28797) );
  XOR U28766 ( .A(n28801), .B(n28802), .Z(n28643) );
  AND U28767 ( .A(n1057), .B(n28803), .Z(n28802) );
  XOR U28768 ( .A(p_input[87]), .B(p_input[71]), .Z(n28803) );
  XOR U28769 ( .A(n28804), .B(n28805), .Z(n28795) );
  AND U28770 ( .A(n28806), .B(n28807), .Z(n28805) );
  XOR U28771 ( .A(n28804), .B(n28658), .Z(n28807) );
  XNOR U28772 ( .A(p_input[102]), .B(n28808), .Z(n28658) );
  AND U28773 ( .A(n1059), .B(n28809), .Z(n28808) );
  XOR U28774 ( .A(p_input[118]), .B(p_input[102]), .Z(n28809) );
  XNOR U28775 ( .A(n28655), .B(n28804), .Z(n28806) );
  XOR U28776 ( .A(n28810), .B(n28811), .Z(n28655) );
  AND U28777 ( .A(n1057), .B(n28812), .Z(n28811) );
  XOR U28778 ( .A(p_input[86]), .B(p_input[70]), .Z(n28812) );
  XOR U28779 ( .A(n28813), .B(n28814), .Z(n28804) );
  AND U28780 ( .A(n28815), .B(n28816), .Z(n28814) );
  XOR U28781 ( .A(n28813), .B(n28670), .Z(n28816) );
  XNOR U28782 ( .A(p_input[101]), .B(n28817), .Z(n28670) );
  AND U28783 ( .A(n1059), .B(n28818), .Z(n28817) );
  XOR U28784 ( .A(p_input[117]), .B(p_input[101]), .Z(n28818) );
  XNOR U28785 ( .A(n28667), .B(n28813), .Z(n28815) );
  XOR U28786 ( .A(n28819), .B(n28820), .Z(n28667) );
  AND U28787 ( .A(n1057), .B(n28821), .Z(n28820) );
  XOR U28788 ( .A(p_input[85]), .B(p_input[69]), .Z(n28821) );
  XOR U28789 ( .A(n28822), .B(n28823), .Z(n28813) );
  AND U28790 ( .A(n28824), .B(n28825), .Z(n28823) );
  XOR U28791 ( .A(n28822), .B(n28682), .Z(n28825) );
  XNOR U28792 ( .A(p_input[100]), .B(n28826), .Z(n28682) );
  AND U28793 ( .A(n1059), .B(n28827), .Z(n28826) );
  XOR U28794 ( .A(p_input[116]), .B(p_input[100]), .Z(n28827) );
  XNOR U28795 ( .A(n28679), .B(n28822), .Z(n28824) );
  XOR U28796 ( .A(n28828), .B(n28829), .Z(n28679) );
  AND U28797 ( .A(n1057), .B(n28830), .Z(n28829) );
  XOR U28798 ( .A(p_input[84]), .B(p_input[68]), .Z(n28830) );
  XOR U28799 ( .A(n28831), .B(n28832), .Z(n28822) );
  AND U28800 ( .A(n28833), .B(n28834), .Z(n28832) );
  XOR U28801 ( .A(n28831), .B(n28694), .Z(n28834) );
  XNOR U28802 ( .A(p_input[99]), .B(n28835), .Z(n28694) );
  AND U28803 ( .A(n1059), .B(n28836), .Z(n28835) );
  XOR U28804 ( .A(p_input[99]), .B(p_input[115]), .Z(n28836) );
  XNOR U28805 ( .A(n28691), .B(n28831), .Z(n28833) );
  XOR U28806 ( .A(n28837), .B(n28838), .Z(n28691) );
  AND U28807 ( .A(n1057), .B(n28839), .Z(n28838) );
  XOR U28808 ( .A(p_input[83]), .B(p_input[67]), .Z(n28839) );
  XOR U28809 ( .A(n28840), .B(n28841), .Z(n28831) );
  AND U28810 ( .A(n28842), .B(n28843), .Z(n28841) );
  XOR U28811 ( .A(n28840), .B(n28706), .Z(n28843) );
  XNOR U28812 ( .A(p_input[98]), .B(n28844), .Z(n28706) );
  AND U28813 ( .A(n1059), .B(n28845), .Z(n28844) );
  XOR U28814 ( .A(p_input[98]), .B(p_input[114]), .Z(n28845) );
  XNOR U28815 ( .A(n28703), .B(n28840), .Z(n28842) );
  XOR U28816 ( .A(n28846), .B(n28847), .Z(n28703) );
  AND U28817 ( .A(n1057), .B(n28848), .Z(n28847) );
  XOR U28818 ( .A(p_input[82]), .B(p_input[66]), .Z(n28848) );
  XOR U28819 ( .A(n28849), .B(n28850), .Z(n28840) );
  AND U28820 ( .A(n28851), .B(n28852), .Z(n28850) );
  XNOR U28821 ( .A(n28853), .B(n28719), .Z(n28852) );
  XNOR U28822 ( .A(p_input[97]), .B(n28854), .Z(n28719) );
  AND U28823 ( .A(n1059), .B(n28855), .Z(n28854) );
  XNOR U28824 ( .A(n28856), .B(p_input[113]), .Z(n28855) );
  IV U28825 ( .A(p_input[97]), .Z(n28856) );
  XNOR U28826 ( .A(n28716), .B(n28849), .Z(n28851) );
  XNOR U28827 ( .A(p_input[65]), .B(n28857), .Z(n28716) );
  AND U28828 ( .A(n1057), .B(n28858), .Z(n28857) );
  XOR U28829 ( .A(p_input[81]), .B(p_input[65]), .Z(n28858) );
  IV U28830 ( .A(n28853), .Z(n28849) );
  AND U28831 ( .A(n28724), .B(n28727), .Z(n28853) );
  XOR U28832 ( .A(p_input[96]), .B(n28859), .Z(n28727) );
  AND U28833 ( .A(n1059), .B(n28860), .Z(n28859) );
  XOR U28834 ( .A(p_input[96]), .B(p_input[112]), .Z(n28860) );
  XOR U28835 ( .A(n28861), .B(n28862), .Z(n1059) );
  AND U28836 ( .A(n28863), .B(n28864), .Z(n28862) );
  XNOR U28837 ( .A(p_input[127]), .B(n28861), .Z(n28864) );
  XOR U28838 ( .A(n28861), .B(p_input[111]), .Z(n28863) );
  XOR U28839 ( .A(n28865), .B(n28866), .Z(n28861) );
  AND U28840 ( .A(n28867), .B(n28868), .Z(n28866) );
  XNOR U28841 ( .A(p_input[126]), .B(n28865), .Z(n28868) );
  XOR U28842 ( .A(n28865), .B(p_input[110]), .Z(n28867) );
  XOR U28843 ( .A(n28869), .B(n28870), .Z(n28865) );
  AND U28844 ( .A(n28871), .B(n28872), .Z(n28870) );
  XNOR U28845 ( .A(p_input[125]), .B(n28869), .Z(n28872) );
  XOR U28846 ( .A(n28869), .B(p_input[109]), .Z(n28871) );
  XOR U28847 ( .A(n28873), .B(n28874), .Z(n28869) );
  AND U28848 ( .A(n28875), .B(n28876), .Z(n28874) );
  XNOR U28849 ( .A(p_input[124]), .B(n28873), .Z(n28876) );
  XOR U28850 ( .A(n28873), .B(p_input[108]), .Z(n28875) );
  XOR U28851 ( .A(n28877), .B(n28878), .Z(n28873) );
  AND U28852 ( .A(n28879), .B(n28880), .Z(n28878) );
  XNOR U28853 ( .A(p_input[123]), .B(n28877), .Z(n28880) );
  XOR U28854 ( .A(n28877), .B(p_input[107]), .Z(n28879) );
  XOR U28855 ( .A(n28881), .B(n28882), .Z(n28877) );
  AND U28856 ( .A(n28883), .B(n28884), .Z(n28882) );
  XNOR U28857 ( .A(p_input[122]), .B(n28881), .Z(n28884) );
  XOR U28858 ( .A(n28881), .B(p_input[106]), .Z(n28883) );
  XOR U28859 ( .A(n28885), .B(n28886), .Z(n28881) );
  AND U28860 ( .A(n28887), .B(n28888), .Z(n28886) );
  XNOR U28861 ( .A(p_input[121]), .B(n28885), .Z(n28888) );
  XOR U28862 ( .A(n28885), .B(p_input[105]), .Z(n28887) );
  XOR U28863 ( .A(n28889), .B(n28890), .Z(n28885) );
  AND U28864 ( .A(n28891), .B(n28892), .Z(n28890) );
  XNOR U28865 ( .A(p_input[120]), .B(n28889), .Z(n28892) );
  XOR U28866 ( .A(n28889), .B(p_input[104]), .Z(n28891) );
  XOR U28867 ( .A(n28893), .B(n28894), .Z(n28889) );
  AND U28868 ( .A(n28895), .B(n28896), .Z(n28894) );
  XNOR U28869 ( .A(p_input[119]), .B(n28893), .Z(n28896) );
  XOR U28870 ( .A(n28893), .B(p_input[103]), .Z(n28895) );
  XOR U28871 ( .A(n28897), .B(n28898), .Z(n28893) );
  AND U28872 ( .A(n28899), .B(n28900), .Z(n28898) );
  XNOR U28873 ( .A(p_input[118]), .B(n28897), .Z(n28900) );
  XOR U28874 ( .A(n28897), .B(p_input[102]), .Z(n28899) );
  XOR U28875 ( .A(n28901), .B(n28902), .Z(n28897) );
  AND U28876 ( .A(n28903), .B(n28904), .Z(n28902) );
  XNOR U28877 ( .A(p_input[117]), .B(n28901), .Z(n28904) );
  XOR U28878 ( .A(n28901), .B(p_input[101]), .Z(n28903) );
  XOR U28879 ( .A(n28905), .B(n28906), .Z(n28901) );
  AND U28880 ( .A(n28907), .B(n28908), .Z(n28906) );
  XNOR U28881 ( .A(p_input[116]), .B(n28905), .Z(n28908) );
  XOR U28882 ( .A(n28905), .B(p_input[100]), .Z(n28907) );
  XOR U28883 ( .A(n28909), .B(n28910), .Z(n28905) );
  AND U28884 ( .A(n28911), .B(n28912), .Z(n28910) );
  XNOR U28885 ( .A(p_input[115]), .B(n28909), .Z(n28912) );
  XOR U28886 ( .A(n28909), .B(p_input[99]), .Z(n28911) );
  XOR U28887 ( .A(n28913), .B(n28914), .Z(n28909) );
  AND U28888 ( .A(n28915), .B(n28916), .Z(n28914) );
  XNOR U28889 ( .A(p_input[114]), .B(n28913), .Z(n28916) );
  XOR U28890 ( .A(n28913), .B(p_input[98]), .Z(n28915) );
  XNOR U28891 ( .A(n28917), .B(n28918), .Z(n28913) );
  AND U28892 ( .A(n28919), .B(n28920), .Z(n28918) );
  XOR U28893 ( .A(p_input[113]), .B(n28917), .Z(n28920) );
  XNOR U28894 ( .A(p_input[97]), .B(n28917), .Z(n28919) );
  AND U28895 ( .A(p_input[112]), .B(n28921), .Z(n28917) );
  IV U28896 ( .A(p_input[96]), .Z(n28921) );
  XNOR U28897 ( .A(p_input[64]), .B(n28922), .Z(n28724) );
  AND U28898 ( .A(n1057), .B(n28923), .Z(n28922) );
  XOR U28899 ( .A(p_input[80]), .B(p_input[64]), .Z(n28923) );
  XOR U28900 ( .A(n28924), .B(n28925), .Z(n1057) );
  AND U28901 ( .A(n28926), .B(n28927), .Z(n28925) );
  XNOR U28902 ( .A(p_input[95]), .B(n28924), .Z(n28927) );
  XOR U28903 ( .A(n28924), .B(p_input[79]), .Z(n28926) );
  XOR U28904 ( .A(n28928), .B(n28929), .Z(n28924) );
  AND U28905 ( .A(n28930), .B(n28931), .Z(n28929) );
  XNOR U28906 ( .A(p_input[94]), .B(n28928), .Z(n28931) );
  XNOR U28907 ( .A(n28928), .B(n28738), .Z(n28930) );
  IV U28908 ( .A(p_input[78]), .Z(n28738) );
  XOR U28909 ( .A(n28932), .B(n28933), .Z(n28928) );
  AND U28910 ( .A(n28934), .B(n28935), .Z(n28933) );
  XNOR U28911 ( .A(p_input[93]), .B(n28932), .Z(n28935) );
  XNOR U28912 ( .A(n28932), .B(n28747), .Z(n28934) );
  IV U28913 ( .A(p_input[77]), .Z(n28747) );
  XOR U28914 ( .A(n28936), .B(n28937), .Z(n28932) );
  AND U28915 ( .A(n28938), .B(n28939), .Z(n28937) );
  XNOR U28916 ( .A(p_input[92]), .B(n28936), .Z(n28939) );
  XNOR U28917 ( .A(n28936), .B(n28756), .Z(n28938) );
  IV U28918 ( .A(p_input[76]), .Z(n28756) );
  XOR U28919 ( .A(n28940), .B(n28941), .Z(n28936) );
  AND U28920 ( .A(n28942), .B(n28943), .Z(n28941) );
  XNOR U28921 ( .A(p_input[91]), .B(n28940), .Z(n28943) );
  XNOR U28922 ( .A(n28940), .B(n28765), .Z(n28942) );
  IV U28923 ( .A(p_input[75]), .Z(n28765) );
  XOR U28924 ( .A(n28944), .B(n28945), .Z(n28940) );
  AND U28925 ( .A(n28946), .B(n28947), .Z(n28945) );
  XNOR U28926 ( .A(p_input[90]), .B(n28944), .Z(n28947) );
  XNOR U28927 ( .A(n28944), .B(n28774), .Z(n28946) );
  IV U28928 ( .A(p_input[74]), .Z(n28774) );
  XOR U28929 ( .A(n28948), .B(n28949), .Z(n28944) );
  AND U28930 ( .A(n28950), .B(n28951), .Z(n28949) );
  XNOR U28931 ( .A(p_input[89]), .B(n28948), .Z(n28951) );
  XNOR U28932 ( .A(n28948), .B(n28783), .Z(n28950) );
  IV U28933 ( .A(p_input[73]), .Z(n28783) );
  XOR U28934 ( .A(n28952), .B(n28953), .Z(n28948) );
  AND U28935 ( .A(n28954), .B(n28955), .Z(n28953) );
  XNOR U28936 ( .A(p_input[88]), .B(n28952), .Z(n28955) );
  XNOR U28937 ( .A(n28952), .B(n28792), .Z(n28954) );
  IV U28938 ( .A(p_input[72]), .Z(n28792) );
  XOR U28939 ( .A(n28956), .B(n28957), .Z(n28952) );
  AND U28940 ( .A(n28958), .B(n28959), .Z(n28957) );
  XNOR U28941 ( .A(p_input[87]), .B(n28956), .Z(n28959) );
  XNOR U28942 ( .A(n28956), .B(n28801), .Z(n28958) );
  IV U28943 ( .A(p_input[71]), .Z(n28801) );
  XOR U28944 ( .A(n28960), .B(n28961), .Z(n28956) );
  AND U28945 ( .A(n28962), .B(n28963), .Z(n28961) );
  XNOR U28946 ( .A(p_input[86]), .B(n28960), .Z(n28963) );
  XNOR U28947 ( .A(n28960), .B(n28810), .Z(n28962) );
  IV U28948 ( .A(p_input[70]), .Z(n28810) );
  XOR U28949 ( .A(n28964), .B(n28965), .Z(n28960) );
  AND U28950 ( .A(n28966), .B(n28967), .Z(n28965) );
  XNOR U28951 ( .A(p_input[85]), .B(n28964), .Z(n28967) );
  XNOR U28952 ( .A(n28964), .B(n28819), .Z(n28966) );
  IV U28953 ( .A(p_input[69]), .Z(n28819) );
  XOR U28954 ( .A(n28968), .B(n28969), .Z(n28964) );
  AND U28955 ( .A(n28970), .B(n28971), .Z(n28969) );
  XNOR U28956 ( .A(p_input[84]), .B(n28968), .Z(n28971) );
  XNOR U28957 ( .A(n28968), .B(n28828), .Z(n28970) );
  IV U28958 ( .A(p_input[68]), .Z(n28828) );
  XOR U28959 ( .A(n28972), .B(n28973), .Z(n28968) );
  AND U28960 ( .A(n28974), .B(n28975), .Z(n28973) );
  XNOR U28961 ( .A(p_input[83]), .B(n28972), .Z(n28975) );
  XNOR U28962 ( .A(n28972), .B(n28837), .Z(n28974) );
  IV U28963 ( .A(p_input[67]), .Z(n28837) );
  XOR U28964 ( .A(n28976), .B(n28977), .Z(n28972) );
  AND U28965 ( .A(n28978), .B(n28979), .Z(n28977) );
  XNOR U28966 ( .A(p_input[82]), .B(n28976), .Z(n28979) );
  XNOR U28967 ( .A(n28976), .B(n28846), .Z(n28978) );
  IV U28968 ( .A(p_input[66]), .Z(n28846) );
  XNOR U28969 ( .A(n28980), .B(n28981), .Z(n28976) );
  AND U28970 ( .A(n28982), .B(n28983), .Z(n28981) );
  XOR U28971 ( .A(p_input[81]), .B(n28980), .Z(n28983) );
  XNOR U28972 ( .A(p_input[65]), .B(n28980), .Z(n28982) );
  AND U28973 ( .A(p_input[80]), .B(n28984), .Z(n28980) );
  IV U28974 ( .A(p_input[64]), .Z(n28984) );
  XOR U28975 ( .A(n28985), .B(n28986), .Z(n28543) );
  AND U28976 ( .A(n584), .B(n28987), .Z(n28986) );
  XNOR U28977 ( .A(n28988), .B(n28985), .Z(n28987) );
  XOR U28978 ( .A(n28989), .B(n28990), .Z(n584) );
  AND U28979 ( .A(n28991), .B(n28992), .Z(n28990) );
  XNOR U28980 ( .A(n28554), .B(n28989), .Z(n28992) );
  AND U28981 ( .A(p_input[63]), .B(p_input[47]), .Z(n28554) );
  XOR U28982 ( .A(n28989), .B(n28553), .Z(n28991) );
  AND U28983 ( .A(p_input[15]), .B(p_input[31]), .Z(n28553) );
  XOR U28984 ( .A(n28993), .B(n28994), .Z(n28989) );
  AND U28985 ( .A(n28995), .B(n28996), .Z(n28994) );
  XOR U28986 ( .A(n28993), .B(n28566), .Z(n28996) );
  XNOR U28987 ( .A(p_input[46]), .B(n28997), .Z(n28566) );
  AND U28988 ( .A(n1067), .B(n28998), .Z(n28997) );
  XOR U28989 ( .A(p_input[62]), .B(p_input[46]), .Z(n28998) );
  XNOR U28990 ( .A(n28563), .B(n28993), .Z(n28995) );
  XOR U28991 ( .A(n28999), .B(n29000), .Z(n28563) );
  AND U28992 ( .A(n1064), .B(n29001), .Z(n29000) );
  XOR U28993 ( .A(p_input[30]), .B(p_input[14]), .Z(n29001) );
  XOR U28994 ( .A(n29002), .B(n29003), .Z(n28993) );
  AND U28995 ( .A(n29004), .B(n29005), .Z(n29003) );
  XOR U28996 ( .A(n29002), .B(n28578), .Z(n29005) );
  XNOR U28997 ( .A(p_input[45]), .B(n29006), .Z(n28578) );
  AND U28998 ( .A(n1067), .B(n29007), .Z(n29006) );
  XOR U28999 ( .A(p_input[61]), .B(p_input[45]), .Z(n29007) );
  XNOR U29000 ( .A(n28575), .B(n29002), .Z(n29004) );
  XOR U29001 ( .A(n29008), .B(n29009), .Z(n28575) );
  AND U29002 ( .A(n1064), .B(n29010), .Z(n29009) );
  XOR U29003 ( .A(p_input[29]), .B(p_input[13]), .Z(n29010) );
  XOR U29004 ( .A(n29011), .B(n29012), .Z(n29002) );
  AND U29005 ( .A(n29013), .B(n29014), .Z(n29012) );
  XOR U29006 ( .A(n29011), .B(n28590), .Z(n29014) );
  XNOR U29007 ( .A(p_input[44]), .B(n29015), .Z(n28590) );
  AND U29008 ( .A(n1067), .B(n29016), .Z(n29015) );
  XOR U29009 ( .A(p_input[60]), .B(p_input[44]), .Z(n29016) );
  XNOR U29010 ( .A(n28587), .B(n29011), .Z(n29013) );
  XOR U29011 ( .A(n29017), .B(n29018), .Z(n28587) );
  AND U29012 ( .A(n1064), .B(n29019), .Z(n29018) );
  XOR U29013 ( .A(p_input[28]), .B(p_input[12]), .Z(n29019) );
  XOR U29014 ( .A(n29020), .B(n29021), .Z(n29011) );
  AND U29015 ( .A(n29022), .B(n29023), .Z(n29021) );
  XOR U29016 ( .A(n29020), .B(n28602), .Z(n29023) );
  XNOR U29017 ( .A(p_input[43]), .B(n29024), .Z(n28602) );
  AND U29018 ( .A(n1067), .B(n29025), .Z(n29024) );
  XOR U29019 ( .A(p_input[59]), .B(p_input[43]), .Z(n29025) );
  XNOR U29020 ( .A(n28599), .B(n29020), .Z(n29022) );
  XOR U29021 ( .A(n29026), .B(n29027), .Z(n28599) );
  AND U29022 ( .A(n1064), .B(n29028), .Z(n29027) );
  XOR U29023 ( .A(p_input[27]), .B(p_input[11]), .Z(n29028) );
  XOR U29024 ( .A(n29029), .B(n29030), .Z(n29020) );
  AND U29025 ( .A(n29031), .B(n29032), .Z(n29030) );
  XOR U29026 ( .A(n29029), .B(n28614), .Z(n29032) );
  XNOR U29027 ( .A(p_input[42]), .B(n29033), .Z(n28614) );
  AND U29028 ( .A(n1067), .B(n29034), .Z(n29033) );
  XOR U29029 ( .A(p_input[58]), .B(p_input[42]), .Z(n29034) );
  XNOR U29030 ( .A(n28611), .B(n29029), .Z(n29031) );
  XOR U29031 ( .A(n29035), .B(n29036), .Z(n28611) );
  AND U29032 ( .A(n1064), .B(n29037), .Z(n29036) );
  XOR U29033 ( .A(p_input[26]), .B(p_input[10]), .Z(n29037) );
  XOR U29034 ( .A(n29038), .B(n29039), .Z(n29029) );
  AND U29035 ( .A(n29040), .B(n29041), .Z(n29039) );
  XOR U29036 ( .A(n29038), .B(n28626), .Z(n29041) );
  XNOR U29037 ( .A(p_input[41]), .B(n29042), .Z(n28626) );
  AND U29038 ( .A(n1067), .B(n29043), .Z(n29042) );
  XOR U29039 ( .A(p_input[57]), .B(p_input[41]), .Z(n29043) );
  XNOR U29040 ( .A(n28623), .B(n29038), .Z(n29040) );
  XOR U29041 ( .A(n29044), .B(n29045), .Z(n28623) );
  AND U29042 ( .A(n1064), .B(n29046), .Z(n29045) );
  XOR U29043 ( .A(p_input[9]), .B(p_input[25]), .Z(n29046) );
  XOR U29044 ( .A(n29047), .B(n29048), .Z(n29038) );
  AND U29045 ( .A(n29049), .B(n29050), .Z(n29048) );
  XOR U29046 ( .A(n29047), .B(n28638), .Z(n29050) );
  XNOR U29047 ( .A(p_input[40]), .B(n29051), .Z(n28638) );
  AND U29048 ( .A(n1067), .B(n29052), .Z(n29051) );
  XOR U29049 ( .A(p_input[56]), .B(p_input[40]), .Z(n29052) );
  XNOR U29050 ( .A(n28635), .B(n29047), .Z(n29049) );
  XOR U29051 ( .A(n29053), .B(n29054), .Z(n28635) );
  AND U29052 ( .A(n1064), .B(n29055), .Z(n29054) );
  XOR U29053 ( .A(p_input[8]), .B(p_input[24]), .Z(n29055) );
  XOR U29054 ( .A(n29056), .B(n29057), .Z(n29047) );
  AND U29055 ( .A(n29058), .B(n29059), .Z(n29057) );
  XOR U29056 ( .A(n29056), .B(n28650), .Z(n29059) );
  XNOR U29057 ( .A(p_input[39]), .B(n29060), .Z(n28650) );
  AND U29058 ( .A(n1067), .B(n29061), .Z(n29060) );
  XOR U29059 ( .A(p_input[55]), .B(p_input[39]), .Z(n29061) );
  XNOR U29060 ( .A(n28647), .B(n29056), .Z(n29058) );
  XOR U29061 ( .A(n29062), .B(n29063), .Z(n28647) );
  AND U29062 ( .A(n1064), .B(n29064), .Z(n29063) );
  XOR U29063 ( .A(p_input[7]), .B(p_input[23]), .Z(n29064) );
  XOR U29064 ( .A(n29065), .B(n29066), .Z(n29056) );
  AND U29065 ( .A(n29067), .B(n29068), .Z(n29066) );
  XOR U29066 ( .A(n29065), .B(n28662), .Z(n29068) );
  XNOR U29067 ( .A(p_input[38]), .B(n29069), .Z(n28662) );
  AND U29068 ( .A(n1067), .B(n29070), .Z(n29069) );
  XOR U29069 ( .A(p_input[54]), .B(p_input[38]), .Z(n29070) );
  XNOR U29070 ( .A(n28659), .B(n29065), .Z(n29067) );
  XOR U29071 ( .A(n29071), .B(n29072), .Z(n28659) );
  AND U29072 ( .A(n1064), .B(n29073), .Z(n29072) );
  XOR U29073 ( .A(p_input[6]), .B(p_input[22]), .Z(n29073) );
  XOR U29074 ( .A(n29074), .B(n29075), .Z(n29065) );
  AND U29075 ( .A(n29076), .B(n29077), .Z(n29075) );
  XOR U29076 ( .A(n29074), .B(n28674), .Z(n29077) );
  XNOR U29077 ( .A(p_input[37]), .B(n29078), .Z(n28674) );
  AND U29078 ( .A(n1067), .B(n29079), .Z(n29078) );
  XOR U29079 ( .A(p_input[53]), .B(p_input[37]), .Z(n29079) );
  XNOR U29080 ( .A(n28671), .B(n29074), .Z(n29076) );
  XOR U29081 ( .A(n29080), .B(n29081), .Z(n28671) );
  AND U29082 ( .A(n1064), .B(n29082), .Z(n29081) );
  XOR U29083 ( .A(p_input[5]), .B(p_input[21]), .Z(n29082) );
  XOR U29084 ( .A(n29083), .B(n29084), .Z(n29074) );
  AND U29085 ( .A(n29085), .B(n29086), .Z(n29084) );
  XOR U29086 ( .A(n29083), .B(n28686), .Z(n29086) );
  XNOR U29087 ( .A(p_input[36]), .B(n29087), .Z(n28686) );
  AND U29088 ( .A(n1067), .B(n29088), .Z(n29087) );
  XOR U29089 ( .A(p_input[52]), .B(p_input[36]), .Z(n29088) );
  XNOR U29090 ( .A(n28683), .B(n29083), .Z(n29085) );
  XOR U29091 ( .A(n29089), .B(n29090), .Z(n28683) );
  AND U29092 ( .A(n1064), .B(n29091), .Z(n29090) );
  XOR U29093 ( .A(p_input[4]), .B(p_input[20]), .Z(n29091) );
  XOR U29094 ( .A(n29092), .B(n29093), .Z(n29083) );
  AND U29095 ( .A(n29094), .B(n29095), .Z(n29093) );
  XOR U29096 ( .A(n29092), .B(n28698), .Z(n29095) );
  XNOR U29097 ( .A(p_input[35]), .B(n29096), .Z(n28698) );
  AND U29098 ( .A(n1067), .B(n29097), .Z(n29096) );
  XOR U29099 ( .A(p_input[51]), .B(p_input[35]), .Z(n29097) );
  XNOR U29100 ( .A(n28695), .B(n29092), .Z(n29094) );
  XOR U29101 ( .A(n29098), .B(n29099), .Z(n28695) );
  AND U29102 ( .A(n1064), .B(n29100), .Z(n29099) );
  XOR U29103 ( .A(p_input[3]), .B(p_input[19]), .Z(n29100) );
  XOR U29104 ( .A(n29101), .B(n29102), .Z(n29092) );
  AND U29105 ( .A(n29103), .B(n29104), .Z(n29102) );
  XOR U29106 ( .A(n29101), .B(n28710), .Z(n29104) );
  XNOR U29107 ( .A(p_input[34]), .B(n29105), .Z(n28710) );
  AND U29108 ( .A(n1067), .B(n29106), .Z(n29105) );
  XOR U29109 ( .A(p_input[50]), .B(p_input[34]), .Z(n29106) );
  XNOR U29110 ( .A(n28707), .B(n29101), .Z(n29103) );
  XOR U29111 ( .A(n29107), .B(n29108), .Z(n28707) );
  AND U29112 ( .A(n1064), .B(n29109), .Z(n29108) );
  XOR U29113 ( .A(p_input[2]), .B(p_input[18]), .Z(n29109) );
  XOR U29114 ( .A(n29110), .B(n29111), .Z(n29101) );
  AND U29115 ( .A(n29112), .B(n29113), .Z(n29111) );
  XNOR U29116 ( .A(n29114), .B(n28723), .Z(n29113) );
  XNOR U29117 ( .A(p_input[33]), .B(n29115), .Z(n28723) );
  AND U29118 ( .A(n1067), .B(n29116), .Z(n29115) );
  XNOR U29119 ( .A(p_input[49]), .B(n29117), .Z(n29116) );
  IV U29120 ( .A(p_input[33]), .Z(n29117) );
  XNOR U29121 ( .A(n28720), .B(n29110), .Z(n29112) );
  XNOR U29122 ( .A(p_input[1]), .B(n29118), .Z(n28720) );
  AND U29123 ( .A(n1064), .B(n29119), .Z(n29118) );
  XOR U29124 ( .A(p_input[1]), .B(p_input[17]), .Z(n29119) );
  IV U29125 ( .A(n29114), .Z(n29110) );
  AND U29126 ( .A(n28985), .B(n28988), .Z(n29114) );
  XOR U29127 ( .A(p_input[32]), .B(n29120), .Z(n28988) );
  AND U29128 ( .A(n1067), .B(n29121), .Z(n29120) );
  XOR U29129 ( .A(p_input[48]), .B(p_input[32]), .Z(n29121) );
  XOR U29130 ( .A(n29122), .B(n29123), .Z(n1067) );
  AND U29131 ( .A(n29124), .B(n29125), .Z(n29123) );
  XNOR U29132 ( .A(p_input[63]), .B(n29122), .Z(n29125) );
  XOR U29133 ( .A(n29122), .B(p_input[47]), .Z(n29124) );
  XOR U29134 ( .A(n29126), .B(n29127), .Z(n29122) );
  AND U29135 ( .A(n29128), .B(n29129), .Z(n29127) );
  XNOR U29136 ( .A(p_input[62]), .B(n29126), .Z(n29129) );
  XOR U29137 ( .A(n29126), .B(p_input[46]), .Z(n29128) );
  XOR U29138 ( .A(n29130), .B(n29131), .Z(n29126) );
  AND U29139 ( .A(n29132), .B(n29133), .Z(n29131) );
  XNOR U29140 ( .A(p_input[61]), .B(n29130), .Z(n29133) );
  XOR U29141 ( .A(n29130), .B(p_input[45]), .Z(n29132) );
  XOR U29142 ( .A(n29134), .B(n29135), .Z(n29130) );
  AND U29143 ( .A(n29136), .B(n29137), .Z(n29135) );
  XNOR U29144 ( .A(p_input[60]), .B(n29134), .Z(n29137) );
  XOR U29145 ( .A(n29134), .B(p_input[44]), .Z(n29136) );
  XOR U29146 ( .A(n29138), .B(n29139), .Z(n29134) );
  AND U29147 ( .A(n29140), .B(n29141), .Z(n29139) );
  XNOR U29148 ( .A(p_input[59]), .B(n29138), .Z(n29141) );
  XOR U29149 ( .A(n29138), .B(p_input[43]), .Z(n29140) );
  XOR U29150 ( .A(n29142), .B(n29143), .Z(n29138) );
  AND U29151 ( .A(n29144), .B(n29145), .Z(n29143) );
  XNOR U29152 ( .A(p_input[58]), .B(n29142), .Z(n29145) );
  XOR U29153 ( .A(n29142), .B(p_input[42]), .Z(n29144) );
  XOR U29154 ( .A(n29146), .B(n29147), .Z(n29142) );
  AND U29155 ( .A(n29148), .B(n29149), .Z(n29147) );
  XNOR U29156 ( .A(p_input[57]), .B(n29146), .Z(n29149) );
  XOR U29157 ( .A(n29146), .B(p_input[41]), .Z(n29148) );
  XOR U29158 ( .A(n29150), .B(n29151), .Z(n29146) );
  AND U29159 ( .A(n29152), .B(n29153), .Z(n29151) );
  XNOR U29160 ( .A(p_input[56]), .B(n29150), .Z(n29153) );
  XOR U29161 ( .A(n29150), .B(p_input[40]), .Z(n29152) );
  XOR U29162 ( .A(n29154), .B(n29155), .Z(n29150) );
  AND U29163 ( .A(n29156), .B(n29157), .Z(n29155) );
  XNOR U29164 ( .A(p_input[55]), .B(n29154), .Z(n29157) );
  XOR U29165 ( .A(n29154), .B(p_input[39]), .Z(n29156) );
  XOR U29166 ( .A(n29158), .B(n29159), .Z(n29154) );
  AND U29167 ( .A(n29160), .B(n29161), .Z(n29159) );
  XNOR U29168 ( .A(p_input[54]), .B(n29158), .Z(n29161) );
  XOR U29169 ( .A(n29158), .B(p_input[38]), .Z(n29160) );
  XOR U29170 ( .A(n29162), .B(n29163), .Z(n29158) );
  AND U29171 ( .A(n29164), .B(n29165), .Z(n29163) );
  XNOR U29172 ( .A(p_input[53]), .B(n29162), .Z(n29165) );
  XOR U29173 ( .A(n29162), .B(p_input[37]), .Z(n29164) );
  XOR U29174 ( .A(n29166), .B(n29167), .Z(n29162) );
  AND U29175 ( .A(n29168), .B(n29169), .Z(n29167) );
  XNOR U29176 ( .A(p_input[52]), .B(n29166), .Z(n29169) );
  XOR U29177 ( .A(n29166), .B(p_input[36]), .Z(n29168) );
  XOR U29178 ( .A(n29170), .B(n29171), .Z(n29166) );
  AND U29179 ( .A(n29172), .B(n29173), .Z(n29171) );
  XNOR U29180 ( .A(p_input[51]), .B(n29170), .Z(n29173) );
  XOR U29181 ( .A(n29170), .B(p_input[35]), .Z(n29172) );
  XOR U29182 ( .A(n29174), .B(n29175), .Z(n29170) );
  AND U29183 ( .A(n29176), .B(n29177), .Z(n29175) );
  XNOR U29184 ( .A(p_input[50]), .B(n29174), .Z(n29177) );
  XOR U29185 ( .A(n29174), .B(p_input[34]), .Z(n29176) );
  XNOR U29186 ( .A(n29178), .B(n29179), .Z(n29174) );
  AND U29187 ( .A(n29180), .B(n29181), .Z(n29179) );
  XOR U29188 ( .A(p_input[49]), .B(n29178), .Z(n29181) );
  XNOR U29189 ( .A(p_input[33]), .B(n29178), .Z(n29180) );
  AND U29190 ( .A(p_input[48]), .B(n29182), .Z(n29178) );
  IV U29191 ( .A(p_input[32]), .Z(n29182) );
  XNOR U29192 ( .A(p_input[0]), .B(n29183), .Z(n28985) );
  AND U29193 ( .A(n1064), .B(n29184), .Z(n29183) );
  XOR U29194 ( .A(p_input[16]), .B(p_input[0]), .Z(n29184) );
  XOR U29195 ( .A(n29185), .B(n29186), .Z(n1064) );
  AND U29196 ( .A(n29187), .B(n29188), .Z(n29186) );
  XNOR U29197 ( .A(p_input[31]), .B(n29185), .Z(n29188) );
  XOR U29198 ( .A(n29185), .B(p_input[15]), .Z(n29187) );
  XOR U29199 ( .A(n29189), .B(n29190), .Z(n29185) );
  AND U29200 ( .A(n29191), .B(n29192), .Z(n29190) );
  XNOR U29201 ( .A(p_input[30]), .B(n29189), .Z(n29192) );
  XNOR U29202 ( .A(n29189), .B(n28999), .Z(n29191) );
  IV U29203 ( .A(p_input[14]), .Z(n28999) );
  XOR U29204 ( .A(n29193), .B(n29194), .Z(n29189) );
  AND U29205 ( .A(n29195), .B(n29196), .Z(n29194) );
  XNOR U29206 ( .A(p_input[29]), .B(n29193), .Z(n29196) );
  XNOR U29207 ( .A(n29193), .B(n29008), .Z(n29195) );
  IV U29208 ( .A(p_input[13]), .Z(n29008) );
  XOR U29209 ( .A(n29197), .B(n29198), .Z(n29193) );
  AND U29210 ( .A(n29199), .B(n29200), .Z(n29198) );
  XNOR U29211 ( .A(p_input[28]), .B(n29197), .Z(n29200) );
  XNOR U29212 ( .A(n29197), .B(n29017), .Z(n29199) );
  IV U29213 ( .A(p_input[12]), .Z(n29017) );
  XOR U29214 ( .A(n29201), .B(n29202), .Z(n29197) );
  AND U29215 ( .A(n29203), .B(n29204), .Z(n29202) );
  XNOR U29216 ( .A(p_input[27]), .B(n29201), .Z(n29204) );
  XNOR U29217 ( .A(n29201), .B(n29026), .Z(n29203) );
  IV U29218 ( .A(p_input[11]), .Z(n29026) );
  XOR U29219 ( .A(n29205), .B(n29206), .Z(n29201) );
  AND U29220 ( .A(n29207), .B(n29208), .Z(n29206) );
  XNOR U29221 ( .A(p_input[26]), .B(n29205), .Z(n29208) );
  XNOR U29222 ( .A(n29205), .B(n29035), .Z(n29207) );
  IV U29223 ( .A(p_input[10]), .Z(n29035) );
  XOR U29224 ( .A(n29209), .B(n29210), .Z(n29205) );
  AND U29225 ( .A(n29211), .B(n29212), .Z(n29210) );
  XNOR U29226 ( .A(p_input[25]), .B(n29209), .Z(n29212) );
  XNOR U29227 ( .A(n29209), .B(n29044), .Z(n29211) );
  IV U29228 ( .A(p_input[9]), .Z(n29044) );
  XOR U29229 ( .A(n29213), .B(n29214), .Z(n29209) );
  AND U29230 ( .A(n29215), .B(n29216), .Z(n29214) );
  XNOR U29231 ( .A(p_input[24]), .B(n29213), .Z(n29216) );
  XNOR U29232 ( .A(n29213), .B(n29053), .Z(n29215) );
  IV U29233 ( .A(p_input[8]), .Z(n29053) );
  XOR U29234 ( .A(n29217), .B(n29218), .Z(n29213) );
  AND U29235 ( .A(n29219), .B(n29220), .Z(n29218) );
  XNOR U29236 ( .A(p_input[23]), .B(n29217), .Z(n29220) );
  XNOR U29237 ( .A(n29217), .B(n29062), .Z(n29219) );
  IV U29238 ( .A(p_input[7]), .Z(n29062) );
  XOR U29239 ( .A(n29221), .B(n29222), .Z(n29217) );
  AND U29240 ( .A(n29223), .B(n29224), .Z(n29222) );
  XNOR U29241 ( .A(p_input[22]), .B(n29221), .Z(n29224) );
  XNOR U29242 ( .A(n29221), .B(n29071), .Z(n29223) );
  IV U29243 ( .A(p_input[6]), .Z(n29071) );
  XOR U29244 ( .A(n29225), .B(n29226), .Z(n29221) );
  AND U29245 ( .A(n29227), .B(n29228), .Z(n29226) );
  XNOR U29246 ( .A(p_input[21]), .B(n29225), .Z(n29228) );
  XNOR U29247 ( .A(n29225), .B(n29080), .Z(n29227) );
  IV U29248 ( .A(p_input[5]), .Z(n29080) );
  XOR U29249 ( .A(n29229), .B(n29230), .Z(n29225) );
  AND U29250 ( .A(n29231), .B(n29232), .Z(n29230) );
  XNOR U29251 ( .A(p_input[20]), .B(n29229), .Z(n29232) );
  XNOR U29252 ( .A(n29229), .B(n29089), .Z(n29231) );
  IV U29253 ( .A(p_input[4]), .Z(n29089) );
  XOR U29254 ( .A(n29233), .B(n29234), .Z(n29229) );
  AND U29255 ( .A(n29235), .B(n29236), .Z(n29234) );
  XNOR U29256 ( .A(p_input[19]), .B(n29233), .Z(n29236) );
  XNOR U29257 ( .A(n29233), .B(n29098), .Z(n29235) );
  IV U29258 ( .A(p_input[3]), .Z(n29098) );
  XOR U29259 ( .A(n29237), .B(n29238), .Z(n29233) );
  AND U29260 ( .A(n29239), .B(n29240), .Z(n29238) );
  XNOR U29261 ( .A(p_input[18]), .B(n29237), .Z(n29240) );
  XNOR U29262 ( .A(n29237), .B(n29107), .Z(n29239) );
  IV U29263 ( .A(p_input[2]), .Z(n29107) );
  XNOR U29264 ( .A(n29241), .B(n29242), .Z(n29237) );
  AND U29265 ( .A(n29243), .B(n29244), .Z(n29242) );
  XOR U29266 ( .A(p_input[17]), .B(n29241), .Z(n29244) );
  XNOR U29267 ( .A(p_input[1]), .B(n29241), .Z(n29243) );
  AND U29268 ( .A(p_input[16]), .B(n29245), .Z(n29241) );
  IV U29269 ( .A(p_input[0]), .Z(n29245) );
endmodule

