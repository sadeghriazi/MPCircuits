
module knn_comb_BMR_W16_K3_N4 ( p_input, o );
  input [79:0] p_input;
  output [47:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953;
  assign \knn_comb_/min_val_out[0][0]  = p_input[48];
  assign \knn_comb_/min_val_out[0][1]  = p_input[49];
  assign \knn_comb_/min_val_out[0][2]  = p_input[50];
  assign \knn_comb_/min_val_out[0][3]  = p_input[51];
  assign \knn_comb_/min_val_out[0][4]  = p_input[52];
  assign \knn_comb_/min_val_out[0][5]  = p_input[53];
  assign \knn_comb_/min_val_out[0][6]  = p_input[54];
  assign \knn_comb_/min_val_out[0][7]  = p_input[55];
  assign \knn_comb_/min_val_out[0][8]  = p_input[56];
  assign \knn_comb_/min_val_out[0][9]  = p_input[57];
  assign \knn_comb_/min_val_out[0][10]  = p_input[58];
  assign \knn_comb_/min_val_out[0][11]  = p_input[59];
  assign \knn_comb_/min_val_out[0][12]  = p_input[60];
  assign \knn_comb_/min_val_out[0][13]  = p_input[61];
  assign \knn_comb_/min_val_out[0][14]  = p_input[62];
  assign \knn_comb_/min_val_out[0][15]  = p_input[63];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][0]  = p_input[16];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][1]  = p_input[17];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][2]  = p_input[18];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][3]  = p_input[19];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][4]  = p_input[20];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][5]  = p_input[21];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][6]  = p_input[22];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][7]  = p_input[23];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][8]  = p_input[24];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][9]  = p_input[25];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][10]  = p_input[26];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][11]  = p_input[27];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][12]  = p_input[28];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][13]  = p_input[29];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][14]  = p_input[30];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][15]  = p_input[31];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[32];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[33];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[34];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[35];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[36];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[37];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[38];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[39];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[40];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[41];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[42];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[43];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[44];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[45];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[46];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[47];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(n3), .B(n4), .Z(n1) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[8]) );
  AND U4 ( .A(n3), .B(n7), .Z(n5) );
  XOR U5 ( .A(n8), .B(n9), .Z(o[7]) );
  AND U6 ( .A(n3), .B(n10), .Z(n8) );
  XOR U7 ( .A(n11), .B(n12), .Z(o[6]) );
  AND U8 ( .A(n3), .B(n13), .Z(n11) );
  XOR U9 ( .A(n14), .B(n15), .Z(o[5]) );
  AND U10 ( .A(n3), .B(n16), .Z(n14) );
  XOR U11 ( .A(n17), .B(n18), .Z(o[4]) );
  AND U12 ( .A(n3), .B(n19), .Z(n17) );
  XOR U13 ( .A(n20), .B(n21), .Z(o[47]) );
  XOR U14 ( .A(n22), .B(n23), .Z(o[46]) );
  XOR U15 ( .A(n24), .B(n25), .Z(o[45]) );
  XOR U16 ( .A(n26), .B(n27), .Z(o[44]) );
  XOR U17 ( .A(n28), .B(n29), .Z(o[43]) );
  XOR U18 ( .A(n30), .B(n31), .Z(o[42]) );
  XOR U19 ( .A(n32), .B(n33), .Z(o[41]) );
  XOR U20 ( .A(n34), .B(n35), .Z(o[40]) );
  XOR U21 ( .A(n36), .B(n37), .Z(o[3]) );
  AND U22 ( .A(n3), .B(n38), .Z(n36) );
  XOR U23 ( .A(n39), .B(n40), .Z(o[39]) );
  XOR U24 ( .A(n41), .B(n42), .Z(o[38]) );
  XOR U25 ( .A(n43), .B(n44), .Z(o[37]) );
  XOR U26 ( .A(n45), .B(n46), .Z(o[36]) );
  XOR U27 ( .A(n47), .B(n48), .Z(o[35]) );
  XOR U28 ( .A(n49), .B(n50), .Z(o[34]) );
  XOR U29 ( .A(n51), .B(n52), .Z(o[33]) );
  XOR U30 ( .A(n53), .B(n54), .Z(o[32]) );
  XOR U31 ( .A(n55), .B(n56), .Z(o[31]) );
  AND U32 ( .A(n57), .B(n58), .Z(n55) );
  XOR U33 ( .A(n59), .B(n60), .Z(o[30]) );
  AND U34 ( .A(n57), .B(n61), .Z(n59) );
  XOR U35 ( .A(n62), .B(n63), .Z(o[2]) );
  AND U36 ( .A(n3), .B(n64), .Z(n62) );
  XOR U37 ( .A(n65), .B(n66), .Z(o[29]) );
  AND U38 ( .A(n57), .B(n67), .Z(n65) );
  XOR U39 ( .A(n68), .B(n69), .Z(o[28]) );
  AND U40 ( .A(n57), .B(n70), .Z(n68) );
  XOR U41 ( .A(n71), .B(n72), .Z(o[27]) );
  AND U42 ( .A(n57), .B(n73), .Z(n71) );
  XOR U43 ( .A(n74), .B(n75), .Z(o[26]) );
  AND U44 ( .A(n57), .B(n76), .Z(n74) );
  XOR U45 ( .A(n77), .B(n78), .Z(o[25]) );
  AND U46 ( .A(n57), .B(n4), .Z(n77) );
  XOR U47 ( .A(n2), .B(n78), .Z(n4) );
  XOR U48 ( .A(n79), .B(n32), .Z(n78) );
  AND U49 ( .A(n80), .B(n81), .Z(n32) );
  XNOR U50 ( .A(n82), .B(n33), .Z(n81) );
  XOR U51 ( .A(n83), .B(n84), .Z(n33) );
  AND U52 ( .A(n85), .B(n86), .Z(n84) );
  XOR U53 ( .A(p_input[9]), .B(n83), .Z(n86) );
  XOR U54 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n87), .Z(n83) );
  AND U55 ( .A(n88), .B(n89), .Z(n87) );
  IV U56 ( .A(n79), .Z(n82) );
  XOR U57 ( .A(n90), .B(n91), .Z(n79) );
  AND U58 ( .A(n92), .B(n93), .Z(n91) );
  XOR U59 ( .A(n94), .B(n95), .Z(n2) );
  AND U60 ( .A(n96), .B(n93), .Z(n95) );
  XNOR U61 ( .A(n97), .B(n90), .Z(n93) );
  XNOR U62 ( .A(n98), .B(n99), .Z(n90) );
  AND U63 ( .A(n100), .B(n89), .Z(n99) );
  XNOR U64 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n98), .Z(
        n89) );
  XNOR U65 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .B(n101), .Z(
        n98) );
  AND U66 ( .A(n102), .B(n103), .Z(n101) );
  IV U67 ( .A(n97), .Z(n94) );
  XNOR U68 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n104), .Z(n97) );
  AND U69 ( .A(n105), .B(n103), .Z(n104) );
  XOR U70 ( .A(\knn_comb_/min_val_out[0][9] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n103) );
  XOR U71 ( .A(n106), .B(n107), .Z(o[24]) );
  AND U72 ( .A(n57), .B(n7), .Z(n106) );
  XOR U73 ( .A(n6), .B(n107), .Z(n7) );
  XOR U74 ( .A(n108), .B(n34), .Z(n107) );
  AND U75 ( .A(n80), .B(n109), .Z(n34) );
  XNOR U76 ( .A(n110), .B(n35), .Z(n109) );
  XOR U77 ( .A(n111), .B(n112), .Z(n35) );
  AND U78 ( .A(n85), .B(n113), .Z(n112) );
  XOR U79 ( .A(p_input[8]), .B(n111), .Z(n113) );
  XOR U80 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n114), .Z(
        n111) );
  AND U81 ( .A(n88), .B(n115), .Z(n114) );
  IV U82 ( .A(n108), .Z(n110) );
  XOR U83 ( .A(n116), .B(n117), .Z(n108) );
  AND U84 ( .A(n92), .B(n118), .Z(n117) );
  XOR U85 ( .A(n119), .B(n120), .Z(n6) );
  AND U86 ( .A(n96), .B(n118), .Z(n120) );
  XNOR U87 ( .A(n121), .B(n116), .Z(n118) );
  XNOR U88 ( .A(n122), .B(n123), .Z(n116) );
  AND U89 ( .A(n100), .B(n115), .Z(n123) );
  XNOR U90 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n122), .Z(
        n115) );
  XNOR U91 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n124), .Z(
        n122) );
  AND U92 ( .A(n102), .B(n125), .Z(n124) );
  IV U93 ( .A(n121), .Z(n119) );
  XNOR U94 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n126), .Z(n121) );
  AND U95 ( .A(n105), .B(n125), .Z(n126) );
  XOR U96 ( .A(\knn_comb_/min_val_out[0][8] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n125) );
  XOR U97 ( .A(n127), .B(n128), .Z(o[23]) );
  AND U98 ( .A(n57), .B(n10), .Z(n127) );
  XOR U99 ( .A(n9), .B(n128), .Z(n10) );
  XOR U100 ( .A(n129), .B(n39), .Z(n128) );
  AND U101 ( .A(n80), .B(n130), .Z(n39) );
  XNOR U102 ( .A(n131), .B(n40), .Z(n130) );
  XOR U103 ( .A(n132), .B(n133), .Z(n40) );
  AND U104 ( .A(n85), .B(n134), .Z(n133) );
  XOR U105 ( .A(p_input[7]), .B(n132), .Z(n134) );
  XOR U106 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n135), .Z(
        n132) );
  AND U107 ( .A(n88), .B(n136), .Z(n135) );
  IV U108 ( .A(n129), .Z(n131) );
  XOR U109 ( .A(n137), .B(n138), .Z(n129) );
  AND U110 ( .A(n92), .B(n139), .Z(n138) );
  XOR U111 ( .A(n140), .B(n141), .Z(n9) );
  AND U112 ( .A(n96), .B(n139), .Z(n141) );
  XNOR U113 ( .A(n142), .B(n137), .Z(n139) );
  XNOR U114 ( .A(n143), .B(n144), .Z(n137) );
  AND U115 ( .A(n100), .B(n136), .Z(n144) );
  XNOR U116 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n143), .Z(
        n136) );
  XNOR U117 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(n145), .Z(
        n143) );
  AND U118 ( .A(n102), .B(n146), .Z(n145) );
  IV U119 ( .A(n142), .Z(n140) );
  XNOR U120 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n147), .Z(n142) );
  AND U121 ( .A(n105), .B(n146), .Z(n147) );
  XOR U122 ( .A(\knn_comb_/min_val_out[0][7] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n146) );
  XOR U123 ( .A(n148), .B(n149), .Z(o[22]) );
  AND U124 ( .A(n57), .B(n13), .Z(n148) );
  XOR U125 ( .A(n12), .B(n149), .Z(n13) );
  XOR U126 ( .A(n150), .B(n41), .Z(n149) );
  AND U127 ( .A(n80), .B(n151), .Z(n41) );
  XNOR U128 ( .A(n152), .B(n42), .Z(n151) );
  XOR U129 ( .A(n153), .B(n154), .Z(n42) );
  AND U130 ( .A(n85), .B(n155), .Z(n154) );
  XOR U131 ( .A(p_input[6]), .B(n153), .Z(n155) );
  XOR U132 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n156), .Z(
        n153) );
  AND U133 ( .A(n88), .B(n157), .Z(n156) );
  IV U134 ( .A(n150), .Z(n152) );
  XOR U135 ( .A(n158), .B(n159), .Z(n150) );
  AND U136 ( .A(n92), .B(n160), .Z(n159) );
  XOR U137 ( .A(n161), .B(n162), .Z(n12) );
  AND U138 ( .A(n96), .B(n160), .Z(n162) );
  XNOR U139 ( .A(n163), .B(n158), .Z(n160) );
  XNOR U140 ( .A(n164), .B(n165), .Z(n158) );
  AND U141 ( .A(n100), .B(n157), .Z(n165) );
  XNOR U142 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n164), .Z(
        n157) );
  XNOR U143 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(n166), .Z(
        n164) );
  AND U144 ( .A(n102), .B(n167), .Z(n166) );
  IV U145 ( .A(n163), .Z(n161) );
  XNOR U146 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n168), .Z(n163) );
  AND U147 ( .A(n105), .B(n167), .Z(n168) );
  XOR U148 ( .A(\knn_comb_/min_val_out[0][6] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n167) );
  XOR U149 ( .A(n169), .B(n170), .Z(o[21]) );
  AND U150 ( .A(n57), .B(n16), .Z(n169) );
  XOR U151 ( .A(n15), .B(n170), .Z(n16) );
  XOR U152 ( .A(n171), .B(n43), .Z(n170) );
  AND U153 ( .A(n80), .B(n172), .Z(n43) );
  XNOR U154 ( .A(n173), .B(n44), .Z(n172) );
  XOR U155 ( .A(n174), .B(n175), .Z(n44) );
  AND U156 ( .A(n85), .B(n176), .Z(n175) );
  XOR U157 ( .A(p_input[5]), .B(n174), .Z(n176) );
  XOR U158 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n177), .Z(
        n174) );
  AND U159 ( .A(n88), .B(n178), .Z(n177) );
  IV U160 ( .A(n171), .Z(n173) );
  XOR U161 ( .A(n179), .B(n180), .Z(n171) );
  AND U162 ( .A(n92), .B(n181), .Z(n180) );
  XOR U163 ( .A(n182), .B(n183), .Z(n15) );
  AND U164 ( .A(n96), .B(n181), .Z(n183) );
  XNOR U165 ( .A(n184), .B(n179), .Z(n181) );
  XNOR U166 ( .A(n185), .B(n186), .Z(n179) );
  AND U167 ( .A(n100), .B(n178), .Z(n186) );
  XNOR U168 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n185), .Z(
        n178) );
  XNOR U169 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n187), .Z(
        n185) );
  AND U170 ( .A(n102), .B(n188), .Z(n187) );
  IV U171 ( .A(n184), .Z(n182) );
  XNOR U172 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n189), .Z(n184) );
  AND U173 ( .A(n105), .B(n188), .Z(n189) );
  XOR U174 ( .A(\knn_comb_/min_val_out[0][5] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n188) );
  XOR U175 ( .A(n190), .B(n191), .Z(o[20]) );
  AND U176 ( .A(n57), .B(n19), .Z(n190) );
  XOR U177 ( .A(n18), .B(n191), .Z(n19) );
  XOR U178 ( .A(n192), .B(n45), .Z(n191) );
  AND U179 ( .A(n80), .B(n193), .Z(n45) );
  XNOR U180 ( .A(n194), .B(n46), .Z(n193) );
  XOR U181 ( .A(n195), .B(n196), .Z(n46) );
  AND U182 ( .A(n85), .B(n197), .Z(n196) );
  XOR U183 ( .A(p_input[4]), .B(n195), .Z(n197) );
  XOR U184 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n198), .Z(
        n195) );
  AND U185 ( .A(n88), .B(n199), .Z(n198) );
  IV U186 ( .A(n192), .Z(n194) );
  XOR U187 ( .A(n200), .B(n201), .Z(n192) );
  AND U188 ( .A(n92), .B(n202), .Z(n201) );
  XOR U189 ( .A(n203), .B(n204), .Z(n18) );
  AND U190 ( .A(n96), .B(n202), .Z(n204) );
  XNOR U191 ( .A(n205), .B(n200), .Z(n202) );
  XNOR U192 ( .A(n206), .B(n207), .Z(n200) );
  AND U193 ( .A(n100), .B(n199), .Z(n207) );
  XNOR U194 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n206), .Z(
        n199) );
  XNOR U195 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n208), .Z(
        n206) );
  AND U196 ( .A(n102), .B(n209), .Z(n208) );
  IV U197 ( .A(n205), .Z(n203) );
  XNOR U198 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n210), .Z(n205) );
  AND U199 ( .A(n105), .B(n209), .Z(n210) );
  XOR U200 ( .A(\knn_comb_/min_val_out[0][4] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n209) );
  XOR U201 ( .A(n211), .B(n212), .Z(o[1]) );
  AND U202 ( .A(n3), .B(n213), .Z(n211) );
  XOR U203 ( .A(n214), .B(n215), .Z(o[19]) );
  AND U204 ( .A(n57), .B(n38), .Z(n214) );
  XOR U205 ( .A(n37), .B(n215), .Z(n38) );
  XOR U206 ( .A(n216), .B(n47), .Z(n215) );
  AND U207 ( .A(n80), .B(n217), .Z(n47) );
  XNOR U208 ( .A(n218), .B(n48), .Z(n217) );
  XOR U209 ( .A(n219), .B(n220), .Z(n48) );
  AND U210 ( .A(n85), .B(n221), .Z(n220) );
  XOR U211 ( .A(p_input[3]), .B(n219), .Z(n221) );
  XOR U212 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n222), .Z(
        n219) );
  AND U213 ( .A(n88), .B(n223), .Z(n222) );
  IV U214 ( .A(n216), .Z(n218) );
  XOR U215 ( .A(n224), .B(n225), .Z(n216) );
  AND U216 ( .A(n92), .B(n226), .Z(n225) );
  XOR U217 ( .A(n227), .B(n228), .Z(n37) );
  AND U218 ( .A(n96), .B(n226), .Z(n228) );
  XNOR U219 ( .A(n229), .B(n224), .Z(n226) );
  XNOR U220 ( .A(n230), .B(n231), .Z(n224) );
  AND U221 ( .A(n100), .B(n223), .Z(n231) );
  XNOR U222 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n230), .Z(
        n223) );
  XNOR U223 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(n232), .Z(
        n230) );
  AND U224 ( .A(n102), .B(n233), .Z(n232) );
  IV U225 ( .A(n229), .Z(n227) );
  XNOR U226 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n234), .Z(n229) );
  AND U227 ( .A(n105), .B(n233), .Z(n234) );
  XOR U228 ( .A(\knn_comb_/min_val_out[0][3] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n233) );
  XOR U229 ( .A(n235), .B(n236), .Z(o[18]) );
  AND U230 ( .A(n57), .B(n64), .Z(n235) );
  XOR U231 ( .A(n63), .B(n236), .Z(n64) );
  XOR U232 ( .A(n237), .B(n49), .Z(n236) );
  AND U233 ( .A(n80), .B(n238), .Z(n49) );
  XOR U234 ( .A(n50), .B(n237), .Z(n238) );
  XOR U235 ( .A(n239), .B(n240), .Z(n50) );
  AND U236 ( .A(n85), .B(n241), .Z(n240) );
  XOR U237 ( .A(p_input[2]), .B(n239), .Z(n241) );
  XOR U238 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n242), .Z(
        n239) );
  AND U239 ( .A(n88), .B(n243), .Z(n242) );
  XOR U240 ( .A(n244), .B(n245), .Z(n237) );
  AND U241 ( .A(n92), .B(n246), .Z(n245) );
  XOR U242 ( .A(n247), .B(n248), .Z(n63) );
  AND U243 ( .A(n96), .B(n246), .Z(n248) );
  XNOR U244 ( .A(n249), .B(n247), .Z(n246) );
  IV U245 ( .A(n244), .Z(n249) );
  XOR U246 ( .A(n250), .B(n251), .Z(n244) );
  AND U247 ( .A(n100), .B(n243), .Z(n251) );
  XOR U248 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n250), .Z(
        n243) );
  XOR U249 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(n252), .Z(
        n250) );
  AND U250 ( .A(n102), .B(n253), .Z(n252) );
  XOR U251 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n254), .Z(n247) );
  AND U252 ( .A(n105), .B(n253), .Z(n254) );
  XOR U253 ( .A(\knn_comb_/min_val_out[0][2] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n253) );
  XOR U254 ( .A(n255), .B(n256), .Z(o[17]) );
  AND U255 ( .A(n57), .B(n213), .Z(n255) );
  XOR U256 ( .A(n212), .B(n256), .Z(n213) );
  XOR U257 ( .A(n257), .B(n51), .Z(n256) );
  AND U258 ( .A(n80), .B(n258), .Z(n51) );
  XOR U259 ( .A(n52), .B(n257), .Z(n258) );
  XOR U260 ( .A(n259), .B(n260), .Z(n52) );
  AND U261 ( .A(n85), .B(n261), .Z(n260) );
  XOR U262 ( .A(p_input[1]), .B(n259), .Z(n261) );
  XOR U263 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n262), .Z(
        n259) );
  AND U264 ( .A(n88), .B(n263), .Z(n262) );
  XOR U265 ( .A(n264), .B(n265), .Z(n257) );
  AND U266 ( .A(n92), .B(n266), .Z(n265) );
  XOR U267 ( .A(n267), .B(n268), .Z(n212) );
  AND U268 ( .A(n96), .B(n266), .Z(n268) );
  XNOR U269 ( .A(n269), .B(n267), .Z(n266) );
  IV U270 ( .A(n264), .Z(n269) );
  XOR U271 ( .A(n270), .B(n271), .Z(n264) );
  AND U272 ( .A(n100), .B(n263), .Z(n271) );
  XOR U273 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n270), .Z(
        n263) );
  XOR U274 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(n272), .Z(
        n270) );
  AND U275 ( .A(n102), .B(n273), .Z(n272) );
  XOR U276 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n274), .Z(n267) );
  AND U277 ( .A(n105), .B(n273), .Z(n274) );
  XOR U278 ( .A(\knn_comb_/min_val_out[0][1] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n273) );
  XOR U279 ( .A(n275), .B(n276), .Z(o[16]) );
  AND U280 ( .A(n57), .B(n277), .Z(n275) );
  XOR U281 ( .A(n278), .B(n279), .Z(n57) );
  MUX U282 ( .IN0(n280), .IN1(n281), .SEL(n278), .F(n279) );
  XNOR U283 ( .A(n282), .B(n283), .Z(n278) );
  XOR U284 ( .A(n284), .B(n285), .Z(o[15]) );
  AND U285 ( .A(n3), .B(n58), .Z(n284) );
  XOR U286 ( .A(n56), .B(n285), .Z(n58) );
  XOR U287 ( .A(n286), .B(n287), .Z(n285) );
  AND U288 ( .A(n96), .B(n288), .Z(n287) );
  XOR U289 ( .A(n289), .B(n20), .Z(n56) );
  AND U290 ( .A(n80), .B(n290), .Z(n20) );
  XOR U291 ( .A(n21), .B(n289), .Z(n290) );
  XOR U292 ( .A(n291), .B(n292), .Z(n21) );
  AND U293 ( .A(n85), .B(n293), .Z(n292) );
  XOR U294 ( .A(p_input[15]), .B(n291), .Z(n293) );
  XOR U295 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n294), .Z(
        n291) );
  AND U296 ( .A(n88), .B(n295), .Z(n294) );
  XOR U297 ( .A(n296), .B(n297), .Z(n289) );
  AND U298 ( .A(n92), .B(n288), .Z(n297) );
  XNOR U299 ( .A(n298), .B(n286), .Z(n288) );
  XOR U300 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n299), .Z(n286) );
  AND U301 ( .A(n105), .B(n300), .Z(n299) );
  IV U302 ( .A(n296), .Z(n298) );
  XOR U303 ( .A(n301), .B(n302), .Z(n296) );
  AND U304 ( .A(n100), .B(n295), .Z(n302) );
  XOR U305 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n301), .Z(
        n295) );
  XOR U306 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n303), .Z(
        n301) );
  AND U307 ( .A(n102), .B(n300), .Z(n303) );
  XOR U308 ( .A(n304), .B(n305), .Z(n300) );
  IV U309 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n305) );
  IV U310 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n304) );
  XOR U311 ( .A(n306), .B(n307), .Z(o[14]) );
  AND U312 ( .A(n3), .B(n61), .Z(n306) );
  XOR U313 ( .A(n60), .B(n307), .Z(n61) );
  XOR U314 ( .A(n308), .B(n309), .Z(n307) );
  AND U315 ( .A(n96), .B(n310), .Z(n309) );
  XOR U316 ( .A(n311), .B(n22), .Z(n60) );
  AND U317 ( .A(n80), .B(n312), .Z(n22) );
  XOR U318 ( .A(n23), .B(n311), .Z(n312) );
  XOR U319 ( .A(n313), .B(n314), .Z(n23) );
  AND U320 ( .A(n85), .B(n315), .Z(n314) );
  XOR U321 ( .A(p_input[14]), .B(n313), .Z(n315) );
  XOR U322 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n316), .Z(
        n313) );
  AND U323 ( .A(n88), .B(n317), .Z(n316) );
  XOR U324 ( .A(n318), .B(n319), .Z(n311) );
  AND U325 ( .A(n92), .B(n310), .Z(n319) );
  XNOR U326 ( .A(n320), .B(n308), .Z(n310) );
  XOR U327 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n321), .Z(n308) );
  AND U328 ( .A(n105), .B(n322), .Z(n321) );
  IV U329 ( .A(n318), .Z(n320) );
  XOR U330 ( .A(n323), .B(n324), .Z(n318) );
  AND U331 ( .A(n100), .B(n317), .Z(n324) );
  XOR U332 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n323), .Z(
        n317) );
  XOR U333 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n325), .Z(
        n323) );
  AND U334 ( .A(n102), .B(n322), .Z(n325) );
  XOR U335 ( .A(n326), .B(n327), .Z(n322) );
  IV U336 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n327) );
  IV U337 ( .A(\knn_comb_/min_val_out[0][14] ), .Z(n326) );
  XOR U338 ( .A(n328), .B(n329), .Z(o[13]) );
  AND U339 ( .A(n3), .B(n67), .Z(n328) );
  XOR U340 ( .A(n66), .B(n329), .Z(n67) );
  XOR U341 ( .A(n330), .B(n331), .Z(n329) );
  AND U342 ( .A(n96), .B(n332), .Z(n331) );
  XOR U343 ( .A(n333), .B(n24), .Z(n66) );
  AND U344 ( .A(n80), .B(n334), .Z(n24) );
  XOR U345 ( .A(n25), .B(n333), .Z(n334) );
  XOR U346 ( .A(n335), .B(n336), .Z(n25) );
  AND U347 ( .A(n85), .B(n337), .Z(n336) );
  XOR U348 ( .A(p_input[13]), .B(n335), .Z(n337) );
  XOR U349 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n338), .Z(
        n335) );
  AND U350 ( .A(n88), .B(n339), .Z(n338) );
  XOR U351 ( .A(n340), .B(n341), .Z(n333) );
  AND U352 ( .A(n92), .B(n332), .Z(n341) );
  XNOR U353 ( .A(n342), .B(n330), .Z(n332) );
  XOR U354 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n343), .Z(n330) );
  AND U355 ( .A(n105), .B(n344), .Z(n343) );
  IV U356 ( .A(n340), .Z(n342) );
  XOR U357 ( .A(n345), .B(n346), .Z(n340) );
  AND U358 ( .A(n100), .B(n339), .Z(n346) );
  XOR U359 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n345), .Z(
        n339) );
  XOR U360 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(n347), .Z(
        n345) );
  AND U361 ( .A(n102), .B(n344), .Z(n347) );
  XOR U362 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n344) );
  XOR U363 ( .A(n348), .B(n349), .Z(o[12]) );
  AND U364 ( .A(n3), .B(n70), .Z(n348) );
  XOR U365 ( .A(n69), .B(n349), .Z(n70) );
  XOR U366 ( .A(n350), .B(n351), .Z(n349) );
  AND U367 ( .A(n96), .B(n352), .Z(n351) );
  XOR U368 ( .A(n353), .B(n26), .Z(n69) );
  AND U369 ( .A(n80), .B(n354), .Z(n26) );
  XOR U370 ( .A(n27), .B(n353), .Z(n354) );
  XOR U371 ( .A(n355), .B(n356), .Z(n27) );
  AND U372 ( .A(n85), .B(n357), .Z(n356) );
  XOR U373 ( .A(p_input[12]), .B(n355), .Z(n357) );
  XOR U374 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n358), .Z(
        n355) );
  AND U375 ( .A(n88), .B(n359), .Z(n358) );
  XOR U376 ( .A(n360), .B(n361), .Z(n353) );
  AND U377 ( .A(n92), .B(n352), .Z(n361) );
  XNOR U378 ( .A(n362), .B(n350), .Z(n352) );
  XOR U379 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n363), .Z(n350) );
  AND U380 ( .A(n105), .B(n364), .Z(n363) );
  IV U381 ( .A(n360), .Z(n362) );
  XOR U382 ( .A(n365), .B(n366), .Z(n360) );
  AND U383 ( .A(n100), .B(n359), .Z(n366) );
  XOR U384 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n365), .Z(
        n359) );
  XOR U385 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n367), .Z(
        n365) );
  AND U386 ( .A(n102), .B(n364), .Z(n367) );
  XOR U387 ( .A(\knn_comb_/min_val_out[0][12] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n364) );
  XOR U388 ( .A(n368), .B(n369), .Z(o[11]) );
  AND U389 ( .A(n3), .B(n73), .Z(n368) );
  XOR U390 ( .A(n72), .B(n369), .Z(n73) );
  XOR U391 ( .A(n370), .B(n371), .Z(n369) );
  AND U392 ( .A(n96), .B(n372), .Z(n371) );
  XOR U393 ( .A(n373), .B(n28), .Z(n72) );
  AND U394 ( .A(n80), .B(n374), .Z(n28) );
  XOR U395 ( .A(n29), .B(n373), .Z(n374) );
  XOR U396 ( .A(n375), .B(n376), .Z(n29) );
  AND U397 ( .A(n85), .B(n377), .Z(n376) );
  XOR U398 ( .A(p_input[11]), .B(n375), .Z(n377) );
  XOR U399 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n378), .Z(
        n375) );
  AND U400 ( .A(n88), .B(n379), .Z(n378) );
  XOR U401 ( .A(n380), .B(n381), .Z(n373) );
  AND U402 ( .A(n92), .B(n372), .Z(n381) );
  XNOR U403 ( .A(n382), .B(n370), .Z(n372) );
  XOR U404 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n383), .Z(n370) );
  AND U405 ( .A(n105), .B(n384), .Z(n383) );
  IV U406 ( .A(n380), .Z(n382) );
  XOR U407 ( .A(n385), .B(n386), .Z(n380) );
  AND U408 ( .A(n100), .B(n379), .Z(n386) );
  XOR U409 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n385), .Z(
        n379) );
  XOR U410 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n387), .Z(
        n385) );
  AND U411 ( .A(n102), .B(n384), .Z(n387) );
  XOR U412 ( .A(n388), .B(n389), .Z(n384) );
  IV U413 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n389) );
  IV U414 ( .A(\knn_comb_/min_val_out[0][11] ), .Z(n388) );
  XOR U415 ( .A(n390), .B(n391), .Z(o[10]) );
  AND U416 ( .A(n3), .B(n76), .Z(n390) );
  XOR U417 ( .A(n75), .B(n391), .Z(n76) );
  XOR U418 ( .A(n392), .B(n393), .Z(n391) );
  AND U419 ( .A(n96), .B(n394), .Z(n393) );
  XOR U420 ( .A(n395), .B(n30), .Z(n75) );
  AND U421 ( .A(n80), .B(n396), .Z(n30) );
  XOR U422 ( .A(n31), .B(n395), .Z(n396) );
  XOR U423 ( .A(n397), .B(n398), .Z(n31) );
  AND U424 ( .A(n85), .B(n399), .Z(n398) );
  XOR U425 ( .A(p_input[10]), .B(n397), .Z(n399) );
  XOR U426 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n400), .Z(
        n397) );
  AND U427 ( .A(n88), .B(n401), .Z(n400) );
  XOR U428 ( .A(n402), .B(n403), .Z(n395) );
  AND U429 ( .A(n92), .B(n394), .Z(n403) );
  XNOR U430 ( .A(n404), .B(n392), .Z(n394) );
  XOR U431 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n405), .Z(n392) );
  AND U432 ( .A(n105), .B(n406), .Z(n405) );
  IV U433 ( .A(n402), .Z(n404) );
  XOR U434 ( .A(n407), .B(n408), .Z(n402) );
  AND U435 ( .A(n100), .B(n401), .Z(n408) );
  XOR U436 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n407), .Z(
        n401) );
  XOR U437 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(n409), .Z(
        n407) );
  AND U438 ( .A(n102), .B(n406), .Z(n409) );
  XOR U439 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n406) );
  XOR U440 ( .A(n410), .B(n411), .Z(o[0]) );
  AND U441 ( .A(n3), .B(n277), .Z(n410) );
  XOR U442 ( .A(n276), .B(n411), .Z(n277) );
  XOR U443 ( .A(n412), .B(n413), .Z(n411) );
  AND U444 ( .A(n96), .B(n414), .Z(n413) );
  XOR U445 ( .A(n415), .B(n53), .Z(n276) );
  AND U446 ( .A(n80), .B(n416), .Z(n53) );
  XOR U447 ( .A(n54), .B(n415), .Z(n416) );
  XOR U448 ( .A(n417), .B(n418), .Z(n54) );
  AND U449 ( .A(n85), .B(n419), .Z(n418) );
  XOR U450 ( .A(p_input[0]), .B(n417), .Z(n419) );
  XOR U451 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n420), .Z(
        n417) );
  AND U452 ( .A(n88), .B(n421), .Z(n420) );
  XOR U453 ( .A(n422), .B(n423), .Z(n415) );
  AND U454 ( .A(n92), .B(n414), .Z(n423) );
  XNOR U455 ( .A(n424), .B(n412), .Z(n414) );
  XOR U456 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n425), .Z(n412) );
  AND U457 ( .A(n105), .B(n426), .Z(n425) );
  IV U458 ( .A(n422), .Z(n424) );
  XOR U459 ( .A(n427), .B(n428), .Z(n422) );
  AND U460 ( .A(n100), .B(n421), .Z(n428) );
  XOR U461 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n427), .Z(
        n421) );
  XOR U462 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(n429), .Z(
        n427) );
  AND U463 ( .A(n102), .B(n426), .Z(n429) );
  XOR U464 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n426) );
  XNOR U465 ( .A(n430), .B(n431), .Z(n3) );
  MUX U466 ( .IN0(n281), .IN1(n280), .SEL(n430), .F(n431) );
  AND U467 ( .A(n432), .B(n433), .Z(n280) );
  NOR U468 ( .A(n434), .B(n435), .Z(n281) );
  IV U469 ( .A(n436), .Z(n434) );
  XOR U470 ( .A(n282), .B(n283), .Z(n430) );
  AND U471 ( .A(n437), .B(n438), .Z(n283) );
  XNOR U472 ( .A(n282), .B(n439), .Z(n438) );
  XOR U473 ( .A(n440), .B(n441), .Z(n439) );
  AND U474 ( .A(n80), .B(n442), .Z(n441) );
  XNOR U475 ( .A(n443), .B(n444), .Z(n442) );
  XNOR U476 ( .A(n282), .B(n445), .Z(n437) );
  XOR U477 ( .A(n446), .B(n447), .Z(n445) );
  AND U478 ( .A(n96), .B(n448), .Z(n447) );
  XNOR U479 ( .A(n446), .B(n449), .Z(n448) );
  XOR U480 ( .A(n450), .B(n451), .Z(n282) );
  AND U481 ( .A(n452), .B(n453), .Z(n451) );
  XOR U482 ( .A(n454), .B(n450), .Z(n453) );
  XNOR U483 ( .A(n455), .B(n456), .Z(n454) );
  AND U484 ( .A(n80), .B(n457), .Z(n456) );
  XNOR U485 ( .A(n458), .B(n455), .Z(n457) );
  XNOR U486 ( .A(n450), .B(n459), .Z(n452) );
  XOR U487 ( .A(n460), .B(n461), .Z(n459) );
  AND U488 ( .A(n96), .B(n462), .Z(n461) );
  XOR U489 ( .A(n463), .B(n464), .Z(n450) );
  AND U490 ( .A(n465), .B(n466), .Z(n464) );
  XOR U491 ( .A(n463), .B(n467), .Z(n466) );
  XOR U492 ( .A(n468), .B(n469), .Z(n467) );
  AND U493 ( .A(n80), .B(n470), .Z(n469) );
  XOR U494 ( .A(n471), .B(n468), .Z(n470) );
  XNOR U495 ( .A(n472), .B(n463), .Z(n465) );
  XNOR U496 ( .A(n473), .B(n474), .Z(n472) );
  AND U497 ( .A(n96), .B(n475), .Z(n474) );
  AND U498 ( .A(n476), .B(n477), .Z(n463) );
  XNOR U499 ( .A(n478), .B(n479), .Z(n477) );
  AND U500 ( .A(n80), .B(n480), .Z(n479) );
  XNOR U501 ( .A(n481), .B(n478), .Z(n480) );
  XNOR U502 ( .A(n482), .B(n483), .Z(n80) );
  NOR U503 ( .A(n484), .B(n485), .Z(n483) );
  XNOR U504 ( .A(n482), .B(n435), .Z(n485) );
  NOR U505 ( .A(n432), .B(n433), .Z(n435) );
  NOR U506 ( .A(n482), .B(n436), .Z(n484) );
  AND U507 ( .A(n486), .B(n487), .Z(n436) );
  IV U508 ( .A(n488), .Z(n486) );
  XOR U509 ( .A(n489), .B(n490), .Z(n482) );
  AND U510 ( .A(n491), .B(n492), .Z(n490) );
  XNOR U511 ( .A(n489), .B(n444), .Z(n492) );
  XOR U512 ( .A(n493), .B(n494), .Z(n444) );
  AND U513 ( .A(n85), .B(n495), .Z(n494) );
  XOR U514 ( .A(n496), .B(n493), .Z(n495) );
  XNOR U515 ( .A(n443), .B(n489), .Z(n491) );
  IV U516 ( .A(n440), .Z(n443) );
  AND U517 ( .A(n497), .B(n449), .Z(n440) );
  XOR U518 ( .A(n498), .B(n499), .Z(n489) );
  AND U519 ( .A(n500), .B(n501), .Z(n499) );
  XOR U520 ( .A(n458), .B(n498), .Z(n501) );
  XOR U521 ( .A(n502), .B(n503), .Z(n458) );
  AND U522 ( .A(n85), .B(n504), .Z(n503) );
  XNOR U523 ( .A(n505), .B(n502), .Z(n504) );
  XOR U524 ( .A(n498), .B(n455), .Z(n500) );
  XOR U525 ( .A(n506), .B(n507), .Z(n455) );
  AND U526 ( .A(n92), .B(n462), .Z(n507) );
  XOR U527 ( .A(n506), .B(n508), .Z(n462) );
  XOR U528 ( .A(n509), .B(n510), .Z(n498) );
  AND U529 ( .A(n511), .B(n512), .Z(n510) );
  XOR U530 ( .A(n509), .B(n471), .Z(n512) );
  XOR U531 ( .A(n513), .B(n514), .Z(n471) );
  AND U532 ( .A(n85), .B(n515), .Z(n514) );
  XOR U533 ( .A(n516), .B(n513), .Z(n515) );
  XNOR U534 ( .A(n468), .B(n509), .Z(n511) );
  XNOR U535 ( .A(n517), .B(n518), .Z(n468) );
  AND U536 ( .A(n92), .B(n475), .Z(n518) );
  XOR U537 ( .A(n517), .B(n473), .Z(n475) );
  AND U538 ( .A(n478), .B(n481), .Z(n509) );
  XOR U539 ( .A(n519), .B(n520), .Z(n481) );
  AND U540 ( .A(n85), .B(n521), .Z(n520) );
  XNOR U541 ( .A(n522), .B(n519), .Z(n521) );
  XNOR U542 ( .A(n523), .B(n524), .Z(n85) );
  NOR U543 ( .A(n525), .B(n526), .Z(n524) );
  XNOR U544 ( .A(n523), .B(n488), .Z(n526) );
  NOR U545 ( .A(n527), .B(n528), .Z(n488) );
  NOR U546 ( .A(n523), .B(n487), .Z(n525) );
  AND U547 ( .A(n496), .B(n529), .Z(n487) );
  XOR U548 ( .A(n530), .B(n531), .Z(n523) );
  AND U549 ( .A(n532), .B(n533), .Z(n531) );
  XNOR U550 ( .A(n530), .B(n496), .Z(n533) );
  XNOR U551 ( .A(n534), .B(n535), .Z(n496) );
  XOR U552 ( .A(n536), .B(n529), .Z(n535) );
  AND U553 ( .A(n505), .B(n537), .Z(n529) );
  AND U554 ( .A(n538), .B(n539), .Z(n536) );
  XOR U555 ( .A(n540), .B(n534), .Z(n538) );
  XOR U556 ( .A(n493), .B(n530), .Z(n532) );
  AND U557 ( .A(n541), .B(n542), .Z(n493) );
  XOR U558 ( .A(n543), .B(n544), .Z(n530) );
  AND U559 ( .A(n545), .B(n546), .Z(n544) );
  XNOR U560 ( .A(n543), .B(n505), .Z(n546) );
  XOR U561 ( .A(n547), .B(n539), .Z(n505) );
  XNOR U562 ( .A(n548), .B(n534), .Z(n539) );
  XOR U563 ( .A(n549), .B(n550), .Z(n534) );
  AND U564 ( .A(n551), .B(n552), .Z(n550) );
  XOR U565 ( .A(n553), .B(n549), .Z(n551) );
  XNOR U566 ( .A(n554), .B(n555), .Z(n548) );
  AND U567 ( .A(n556), .B(n557), .Z(n555) );
  XOR U568 ( .A(n554), .B(n558), .Z(n556) );
  XNOR U569 ( .A(n540), .B(n537), .Z(n547) );
  AND U570 ( .A(n559), .B(n560), .Z(n537) );
  XOR U571 ( .A(n561), .B(n562), .Z(n540) );
  AND U572 ( .A(n563), .B(n564), .Z(n562) );
  XOR U573 ( .A(n561), .B(n565), .Z(n563) );
  XNOR U574 ( .A(n502), .B(n543), .Z(n545) );
  XNOR U575 ( .A(n566), .B(n567), .Z(n502) );
  AND U576 ( .A(n88), .B(n568), .Z(n567) );
  XOR U577 ( .A(n569), .B(n570), .Z(n543) );
  AND U578 ( .A(n571), .B(n572), .Z(n570) );
  XNOR U579 ( .A(n569), .B(n559), .Z(n572) );
  IV U580 ( .A(n516), .Z(n559) );
  XNOR U581 ( .A(n573), .B(n552), .Z(n516) );
  XNOR U582 ( .A(n574), .B(n558), .Z(n552) );
  XOR U583 ( .A(n575), .B(n576), .Z(n558) );
  NOR U584 ( .A(n577), .B(n578), .Z(n576) );
  XNOR U585 ( .A(n575), .B(n579), .Z(n577) );
  XNOR U586 ( .A(n557), .B(n549), .Z(n574) );
  XOR U587 ( .A(n580), .B(n581), .Z(n549) );
  AND U588 ( .A(n582), .B(n583), .Z(n581) );
  XOR U589 ( .A(n584), .B(n585), .Z(n582) );
  XNOR U590 ( .A(n586), .B(n554), .Z(n557) );
  XOR U591 ( .A(n587), .B(n588), .Z(n554) );
  NOR U592 ( .A(n589), .B(n590), .Z(n588) );
  XNOR U593 ( .A(n587), .B(n591), .Z(n589) );
  XNOR U594 ( .A(n592), .B(n593), .Z(n586) );
  NOR U595 ( .A(n594), .B(n595), .Z(n593) );
  XNOR U596 ( .A(n592), .B(n596), .Z(n594) );
  XNOR U597 ( .A(n553), .B(n560), .Z(n573) );
  AND U598 ( .A(n522), .B(n597), .Z(n560) );
  XOR U599 ( .A(n565), .B(n564), .Z(n553) );
  XNOR U600 ( .A(n598), .B(n561), .Z(n564) );
  XOR U601 ( .A(n599), .B(n600), .Z(n561) );
  AND U602 ( .A(n601), .B(n602), .Z(n600) );
  XOR U603 ( .A(n599), .B(n603), .Z(n601) );
  XNOR U604 ( .A(n604), .B(n605), .Z(n598) );
  NOR U605 ( .A(n606), .B(n607), .Z(n605) );
  XNOR U606 ( .A(n604), .B(n608), .Z(n606) );
  XOR U607 ( .A(n609), .B(n610), .Z(n565) );
  NOR U608 ( .A(n611), .B(n612), .Z(n610) );
  XNOR U609 ( .A(n609), .B(n613), .Z(n611) );
  XNOR U610 ( .A(n513), .B(n569), .Z(n571) );
  XNOR U611 ( .A(n614), .B(n615), .Z(n513) );
  AND U612 ( .A(n88), .B(n616), .Z(n615) );
  XNOR U613 ( .A(n617), .B(n618), .Z(n616) );
  NOR U614 ( .A(n519), .B(n522), .Z(n569) );
  XOR U615 ( .A(n619), .B(n597), .Z(n522) );
  XOR U616 ( .A(p_input[0]), .B(p_input[64]), .Z(n597) );
  XOR U617 ( .A(n585), .B(n583), .Z(n619) );
  XNOR U618 ( .A(n620), .B(n591), .Z(n583) );
  XNOR U619 ( .A(n579), .B(n578), .Z(n591) );
  XOR U620 ( .A(n621), .B(n575), .Z(n578) );
  XOR U621 ( .A(p_input[10]), .B(p_input[74]), .Z(n575) );
  XNOR U622 ( .A(p_input[11]), .B(p_input[75]), .Z(n621) );
  XOR U623 ( .A(p_input[12]), .B(p_input[76]), .Z(n579) );
  XNOR U624 ( .A(n590), .B(n584), .Z(n620) );
  IV U625 ( .A(n580), .Z(n584) );
  XOR U626 ( .A(p_input[1]), .B(p_input[65]), .Z(n580) );
  XOR U627 ( .A(n622), .B(n596), .Z(n590) );
  XOR U628 ( .A(p_input[15]), .B(p_input[79]), .Z(n596) );
  XOR U629 ( .A(n587), .B(n595), .Z(n622) );
  XOR U630 ( .A(n623), .B(n592), .Z(n595) );
  XOR U631 ( .A(p_input[13]), .B(p_input[77]), .Z(n592) );
  XNOR U632 ( .A(p_input[14]), .B(p_input[78]), .Z(n623) );
  XOR U633 ( .A(p_input[73]), .B(p_input[9]), .Z(n587) );
  XNOR U634 ( .A(n603), .B(n602), .Z(n585) );
  XNOR U635 ( .A(n624), .B(n608), .Z(n602) );
  XOR U636 ( .A(p_input[72]), .B(p_input[8]), .Z(n608) );
  XOR U637 ( .A(n599), .B(n607), .Z(n624) );
  XOR U638 ( .A(n625), .B(n604), .Z(n607) );
  XOR U639 ( .A(p_input[6]), .B(p_input[70]), .Z(n604) );
  XNOR U640 ( .A(p_input[71]), .B(p_input[7]), .Z(n625) );
  XOR U641 ( .A(p_input[2]), .B(p_input[66]), .Z(n599) );
  XNOR U642 ( .A(n613), .B(n612), .Z(n603) );
  XOR U643 ( .A(n626), .B(n609), .Z(n612) );
  XOR U644 ( .A(p_input[3]), .B(p_input[67]), .Z(n609) );
  XNOR U645 ( .A(p_input[4]), .B(p_input[68]), .Z(n626) );
  XOR U646 ( .A(p_input[5]), .B(p_input[69]), .Z(n613) );
  XOR U647 ( .A(n627), .B(n628), .Z(n519) );
  AND U648 ( .A(n88), .B(n629), .Z(n628) );
  XNOR U649 ( .A(n630), .B(n631), .Z(n88) );
  NOR U650 ( .A(n632), .B(n633), .Z(n631) );
  XOR U651 ( .A(n630), .B(n527), .Z(n633) );
  XNOR U652 ( .A(n634), .B(n635), .Z(n478) );
  AND U653 ( .A(n92), .B(n636), .Z(n635) );
  XOR U654 ( .A(n637), .B(n638), .Z(n92) );
  MUX U655 ( .IN0(n433), .IN1(n432), .SEL(n637), .F(n638) );
  XNOR U656 ( .A(n639), .B(n640), .Z(n637) );
  AND U657 ( .A(n641), .B(n642), .Z(n640) );
  XNOR U658 ( .A(n639), .B(n449), .Z(n642) );
  XOR U659 ( .A(n639), .B(n497), .Z(n641) );
  XOR U660 ( .A(n643), .B(n644), .Z(n639) );
  AND U661 ( .A(n645), .B(n646), .Z(n644) );
  XOR U662 ( .A(n643), .B(n508), .Z(n645) );
  IV U663 ( .A(n460), .Z(n508) );
  XOR U664 ( .A(n647), .B(n648), .Z(n476) );
  AND U665 ( .A(n96), .B(n636), .Z(n648) );
  XNOR U666 ( .A(n634), .B(n647), .Z(n636) );
  XNOR U667 ( .A(n649), .B(n650), .Z(n96) );
  MUX U668 ( .IN0(n432), .IN1(n433), .SEL(n649), .F(n650) );
  AND U669 ( .A(n651), .B(n652), .Z(n433) );
  AND U670 ( .A(n527), .B(n528), .Z(n432) );
  IV U671 ( .A(n653), .Z(n527) );
  XOR U672 ( .A(n654), .B(n655), .Z(n649) );
  AND U673 ( .A(n656), .B(n657), .Z(n655) );
  XNOR U674 ( .A(n449), .B(n654), .Z(n657) );
  XNOR U675 ( .A(n658), .B(n659), .Z(n449) );
  AND U676 ( .A(n100), .B(n660), .Z(n659) );
  XOR U677 ( .A(n661), .B(n658), .Z(n660) );
  IV U678 ( .A(n542), .Z(n661) );
  XNOR U679 ( .A(n446), .B(n654), .Z(n656) );
  IV U680 ( .A(n497), .Z(n446) );
  XOR U681 ( .A(n662), .B(n663), .Z(n497) );
  AND U682 ( .A(n105), .B(n664), .Z(n663) );
  XOR U683 ( .A(n665), .B(n662), .Z(n664) );
  XOR U684 ( .A(n643), .B(n666), .Z(n654) );
  AND U685 ( .A(n667), .B(n646), .Z(n666) );
  XNOR U686 ( .A(n506), .B(n643), .Z(n646) );
  XOR U687 ( .A(n668), .B(n669), .Z(n506) );
  AND U688 ( .A(n100), .B(n568), .Z(n669) );
  XOR U689 ( .A(n566), .B(n668), .Z(n568) );
  XNOR U690 ( .A(n460), .B(n643), .Z(n667) );
  XNOR U691 ( .A(n670), .B(n671), .Z(n460) );
  AND U692 ( .A(n105), .B(n672), .Z(n671) );
  XOR U693 ( .A(n673), .B(n674), .Z(n643) );
  AND U694 ( .A(n675), .B(n676), .Z(n674) );
  XNOR U695 ( .A(n673), .B(n517), .Z(n676) );
  XOR U696 ( .A(n618), .B(n677), .Z(n517) );
  AND U697 ( .A(n100), .B(n678), .Z(n677) );
  XOR U698 ( .A(n614), .B(n618), .Z(n678) );
  XNOR U699 ( .A(n679), .B(n673), .Z(n675) );
  IV U700 ( .A(n473), .Z(n679) );
  XOR U701 ( .A(n680), .B(n681), .Z(n473) );
  AND U702 ( .A(n105), .B(n682), .Z(n681) );
  AND U703 ( .A(n647), .B(n634), .Z(n673) );
  XNOR U704 ( .A(n683), .B(n684), .Z(n634) );
  AND U705 ( .A(n100), .B(n629), .Z(n684) );
  XNOR U706 ( .A(n627), .B(n683), .Z(n629) );
  XNOR U707 ( .A(n630), .B(n685), .Z(n100) );
  NOR U708 ( .A(n632), .B(n686), .Z(n685) );
  XNOR U709 ( .A(n630), .B(n653), .Z(n686) );
  NOR U710 ( .A(n651), .B(n652), .Z(n653) );
  NOR U711 ( .A(n630), .B(n528), .Z(n632) );
  AND U712 ( .A(n542), .B(n687), .Z(n528) );
  XOR U713 ( .A(n688), .B(n689), .Z(n630) );
  AND U714 ( .A(n690), .B(n691), .Z(n689) );
  XNOR U715 ( .A(n542), .B(n688), .Z(n691) );
  XNOR U716 ( .A(n692), .B(n693), .Z(n542) );
  XOR U717 ( .A(n694), .B(n687), .Z(n693) );
  AND U718 ( .A(n566), .B(n695), .Z(n687) );
  AND U719 ( .A(n696), .B(n697), .Z(n694) );
  XOR U720 ( .A(n698), .B(n692), .Z(n696) );
  XNOR U721 ( .A(n658), .B(n688), .Z(n690) );
  IV U722 ( .A(n541), .Z(n658) );
  AND U723 ( .A(n662), .B(n665), .Z(n541) );
  XOR U724 ( .A(n699), .B(n700), .Z(n688) );
  AND U725 ( .A(n701), .B(n702), .Z(n700) );
  XNOR U726 ( .A(n566), .B(n699), .Z(n702) );
  XOR U727 ( .A(n703), .B(n697), .Z(n566) );
  XNOR U728 ( .A(n704), .B(n692), .Z(n697) );
  XOR U729 ( .A(n705), .B(n706), .Z(n692) );
  AND U730 ( .A(n707), .B(n708), .Z(n706) );
  XOR U731 ( .A(n709), .B(n705), .Z(n707) );
  XNOR U732 ( .A(n710), .B(n711), .Z(n704) );
  AND U733 ( .A(n712), .B(n713), .Z(n711) );
  XOR U734 ( .A(n710), .B(n714), .Z(n712) );
  XNOR U735 ( .A(n698), .B(n695), .Z(n703) );
  AND U736 ( .A(n614), .B(n715), .Z(n695) );
  XOR U737 ( .A(n716), .B(n717), .Z(n698) );
  AND U738 ( .A(n718), .B(n719), .Z(n717) );
  XOR U739 ( .A(n716), .B(n720), .Z(n718) );
  XOR U740 ( .A(n699), .B(n668), .Z(n701) );
  XOR U741 ( .A(n721), .B(n722), .Z(n668) );
  AND U742 ( .A(n102), .B(n672), .Z(n722) );
  XOR U743 ( .A(n721), .B(n670), .Z(n672) );
  XOR U744 ( .A(n723), .B(n724), .Z(n699) );
  AND U745 ( .A(n725), .B(n726), .Z(n724) );
  XNOR U746 ( .A(n723), .B(n614), .Z(n726) );
  IV U747 ( .A(n617), .Z(n614) );
  XNOR U748 ( .A(n727), .B(n708), .Z(n617) );
  XNOR U749 ( .A(n728), .B(n714), .Z(n708) );
  XOR U750 ( .A(n729), .B(n730), .Z(n714) );
  NOR U751 ( .A(n731), .B(n732), .Z(n730) );
  XNOR U752 ( .A(n729), .B(n733), .Z(n731) );
  XNOR U753 ( .A(n713), .B(n705), .Z(n728) );
  XOR U754 ( .A(n734), .B(n735), .Z(n705) );
  AND U755 ( .A(n736), .B(n737), .Z(n735) );
  XNOR U756 ( .A(n734), .B(n738), .Z(n736) );
  XNOR U757 ( .A(n739), .B(n710), .Z(n713) );
  XOR U758 ( .A(n740), .B(n741), .Z(n710) );
  AND U759 ( .A(n742), .B(n743), .Z(n741) );
  XNOR U760 ( .A(n744), .B(n745), .Z(n742) );
  XNOR U761 ( .A(n746), .B(n747), .Z(n739) );
  NOR U762 ( .A(n748), .B(n749), .Z(n747) );
  XOR U763 ( .A(n746), .B(n750), .Z(n748) );
  XNOR U764 ( .A(n709), .B(n715), .Z(n727) );
  NOR U765 ( .A(n627), .B(n751), .Z(n715) );
  XOR U766 ( .A(n720), .B(n719), .Z(n709) );
  XNOR U767 ( .A(n752), .B(n716), .Z(n719) );
  XOR U768 ( .A(n753), .B(n754), .Z(n716) );
  AND U769 ( .A(n755), .B(n756), .Z(n754) );
  XOR U770 ( .A(n753), .B(n757), .Z(n755) );
  XNOR U771 ( .A(n758), .B(n759), .Z(n752) );
  NOR U772 ( .A(n760), .B(n761), .Z(n759) );
  XOR U773 ( .A(n758), .B(n762), .Z(n760) );
  XOR U774 ( .A(n763), .B(n764), .Z(n720) );
  NOR U775 ( .A(n765), .B(n766), .Z(n764) );
  XNOR U776 ( .A(n763), .B(n767), .Z(n765) );
  XOR U777 ( .A(n618), .B(n723), .Z(n725) );
  XOR U778 ( .A(n768), .B(n769), .Z(n618) );
  AND U779 ( .A(n102), .B(n682), .Z(n769) );
  XOR U780 ( .A(n768), .B(n680), .Z(n682) );
  AND U781 ( .A(n683), .B(n627), .Z(n723) );
  XOR U782 ( .A(n770), .B(n751), .Z(n627) );
  XNOR U783 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(
        p_input[64]), .Z(n751) );
  XOR U784 ( .A(n738), .B(n737), .Z(n770) );
  XNOR U785 ( .A(n771), .B(n745), .Z(n737) );
  XNOR U786 ( .A(n733), .B(n732), .Z(n745) );
  XOR U787 ( .A(n772), .B(n729), .Z(n732) );
  XOR U788 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(
        p_input[74]), .Z(n729) );
  XOR U789 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n773), .Z(
        n772) );
  XOR U790 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(
        p_input[76]), .Z(n733) );
  XNOR U791 ( .A(n743), .B(n734), .Z(n771) );
  XOR U792 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(p_input[65]), .Z(n734) );
  XOR U793 ( .A(n774), .B(n750), .Z(n743) );
  XNOR U794 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(
        p_input[79]), .Z(n750) );
  XOR U795 ( .A(n740), .B(n749), .Z(n774) );
  XOR U796 ( .A(n775), .B(n746), .Z(n749) );
  XOR U797 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(
        p_input[77]), .Z(n746) );
  XOR U798 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n776), .Z(
        n775) );
  IV U799 ( .A(n744), .Z(n740) );
  XNOR U800 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(
        p_input[73]), .Z(n744) );
  XNOR U801 ( .A(n757), .B(n756), .Z(n738) );
  XOR U802 ( .A(n777), .B(n762), .Z(n756) );
  XNOR U803 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(
        p_input[72]), .Z(n762) );
  XOR U804 ( .A(n753), .B(n761), .Z(n777) );
  XOR U805 ( .A(n778), .B(n758), .Z(n761) );
  XOR U806 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(p_input[70]), .Z(n758) );
  XNOR U807 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(
        p_input[71]), .Z(n778) );
  XOR U808 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(p_input[66]), .Z(n753) );
  XNOR U809 ( .A(n767), .B(n766), .Z(n757) );
  XOR U810 ( .A(n779), .B(n763), .Z(n766) );
  XOR U811 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(p_input[67]), .Z(n763) );
  XNOR U812 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(
        p_input[68]), .Z(n779) );
  XOR U813 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(p_input[69]), .Z(n767) );
  XNOR U814 ( .A(n780), .B(n781), .Z(n683) );
  AND U815 ( .A(n102), .B(n782), .Z(n781) );
  XNOR U816 ( .A(n783), .B(n784), .Z(n102) );
  MUX U817 ( .IN0(n651), .IN1(n652), .SEL(n783), .F(n784) );
  XOR U818 ( .A(n785), .B(n786), .Z(n783) );
  AND U819 ( .A(n787), .B(n788), .Z(n786) );
  XOR U820 ( .A(n785), .B(n662), .Z(n787) );
  XOR U821 ( .A(n789), .B(n790), .Z(n647) );
  AND U822 ( .A(n105), .B(n782), .Z(n790) );
  XOR U823 ( .A(n791), .B(n789), .Z(n782) );
  XNOR U824 ( .A(n792), .B(n793), .Z(n105) );
  MUX U825 ( .IN0(n651), .IN1(n652), .SEL(n792), .F(n793) );
  AND U826 ( .A(n662), .B(n794), .Z(n652) );
  AND U827 ( .A(n665), .B(n795), .Z(n651) );
  XOR U828 ( .A(n785), .B(n796), .Z(n792) );
  AND U829 ( .A(n797), .B(n788), .Z(n796) );
  XNOR U830 ( .A(n665), .B(n785), .Z(n788) );
  XNOR U831 ( .A(n798), .B(n799), .Z(n665) );
  XOR U832 ( .A(n800), .B(n795), .Z(n799) );
  AND U833 ( .A(n721), .B(n801), .Z(n795) );
  AND U834 ( .A(n802), .B(n803), .Z(n800) );
  XOR U835 ( .A(n804), .B(n798), .Z(n802) );
  XNOR U836 ( .A(n805), .B(n785), .Z(n797) );
  IV U837 ( .A(n662), .Z(n805) );
  XNOR U838 ( .A(n806), .B(n807), .Z(n662) );
  XOR U839 ( .A(n808), .B(n794), .Z(n807) );
  AND U840 ( .A(n670), .B(n809), .Z(n794) );
  AND U841 ( .A(n810), .B(n811), .Z(n808) );
  XNOR U842 ( .A(n806), .B(n812), .Z(n810) );
  XOR U843 ( .A(n813), .B(n814), .Z(n785) );
  AND U844 ( .A(n815), .B(n816), .Z(n814) );
  XNOR U845 ( .A(n721), .B(n813), .Z(n816) );
  XOR U846 ( .A(n817), .B(n803), .Z(n721) );
  XNOR U847 ( .A(n818), .B(n798), .Z(n803) );
  XOR U848 ( .A(n819), .B(n820), .Z(n798) );
  AND U849 ( .A(n821), .B(n822), .Z(n820) );
  XOR U850 ( .A(n823), .B(n819), .Z(n821) );
  XNOR U851 ( .A(n824), .B(n825), .Z(n818) );
  AND U852 ( .A(n826), .B(n827), .Z(n825) );
  XOR U853 ( .A(n824), .B(n828), .Z(n826) );
  XNOR U854 ( .A(n804), .B(n801), .Z(n817) );
  AND U855 ( .A(n768), .B(n829), .Z(n801) );
  XOR U856 ( .A(n830), .B(n831), .Z(n804) );
  AND U857 ( .A(n832), .B(n833), .Z(n831) );
  XOR U858 ( .A(n830), .B(n834), .Z(n832) );
  XOR U859 ( .A(n813), .B(n670), .Z(n815) );
  XNOR U860 ( .A(n835), .B(n812), .Z(n670) );
  XNOR U861 ( .A(n836), .B(n837), .Z(n812) );
  AND U862 ( .A(n838), .B(n839), .Z(n837) );
  XOR U863 ( .A(n836), .B(n840), .Z(n838) );
  XNOR U864 ( .A(n811), .B(n809), .Z(n835) );
  AND U865 ( .A(n680), .B(n841), .Z(n809) );
  XNOR U866 ( .A(n842), .B(n806), .Z(n811) );
  XOR U867 ( .A(n843), .B(n844), .Z(n806) );
  AND U868 ( .A(n845), .B(n846), .Z(n844) );
  XOR U869 ( .A(n843), .B(n847), .Z(n845) );
  XNOR U870 ( .A(n848), .B(n849), .Z(n842) );
  AND U871 ( .A(n850), .B(n851), .Z(n849) );
  XNOR U872 ( .A(n848), .B(n852), .Z(n850) );
  XOR U873 ( .A(n853), .B(n854), .Z(n813) );
  AND U874 ( .A(n855), .B(n856), .Z(n854) );
  XNOR U875 ( .A(n853), .B(n768), .Z(n856) );
  XOR U876 ( .A(n857), .B(n822), .Z(n768) );
  XNOR U877 ( .A(n858), .B(n828), .Z(n822) );
  XOR U878 ( .A(n859), .B(n860), .Z(n828) );
  NOR U879 ( .A(n861), .B(n862), .Z(n860) );
  XNOR U880 ( .A(n859), .B(n863), .Z(n861) );
  XNOR U881 ( .A(n827), .B(n819), .Z(n858) );
  XOR U882 ( .A(n864), .B(n865), .Z(n819) );
  AND U883 ( .A(n866), .B(n867), .Z(n865) );
  XNOR U884 ( .A(n864), .B(n868), .Z(n866) );
  XNOR U885 ( .A(n869), .B(n824), .Z(n827) );
  XOR U886 ( .A(n870), .B(n871), .Z(n824) );
  AND U887 ( .A(n872), .B(n873), .Z(n871) );
  XOR U888 ( .A(n870), .B(n874), .Z(n872) );
  XNOR U889 ( .A(n875), .B(n876), .Z(n869) );
  NOR U890 ( .A(n877), .B(n878), .Z(n876) );
  XOR U891 ( .A(n875), .B(n879), .Z(n877) );
  XNOR U892 ( .A(n823), .B(n829), .Z(n857) );
  AND U893 ( .A(n791), .B(n880), .Z(n829) );
  IV U894 ( .A(n780), .Z(n791) );
  XOR U895 ( .A(n834), .B(n833), .Z(n823) );
  XNOR U896 ( .A(n881), .B(n830), .Z(n833) );
  XOR U897 ( .A(n882), .B(n883), .Z(n830) );
  AND U898 ( .A(n884), .B(n885), .Z(n883) );
  XOR U899 ( .A(n882), .B(n886), .Z(n884) );
  XNOR U900 ( .A(n887), .B(n888), .Z(n881) );
  NOR U901 ( .A(n889), .B(n890), .Z(n888) );
  XNOR U902 ( .A(n887), .B(n891), .Z(n889) );
  XOR U903 ( .A(n892), .B(n893), .Z(n834) );
  NOR U904 ( .A(n894), .B(n895), .Z(n893) );
  XNOR U905 ( .A(n892), .B(n896), .Z(n894) );
  XNOR U906 ( .A(n897), .B(n853), .Z(n855) );
  IV U907 ( .A(n680), .Z(n897) );
  XOR U908 ( .A(n898), .B(n847), .Z(n680) );
  XOR U909 ( .A(n840), .B(n839), .Z(n847) );
  XNOR U910 ( .A(n899), .B(n836), .Z(n839) );
  XOR U911 ( .A(n900), .B(n901), .Z(n836) );
  AND U912 ( .A(n902), .B(n903), .Z(n901) );
  XOR U913 ( .A(n900), .B(n904), .Z(n902) );
  XNOR U914 ( .A(n905), .B(n906), .Z(n899) );
  NOR U915 ( .A(n907), .B(n908), .Z(n906) );
  XNOR U916 ( .A(n905), .B(n909), .Z(n907) );
  XOR U917 ( .A(n910), .B(n911), .Z(n840) );
  NOR U918 ( .A(n912), .B(n913), .Z(n911) );
  XNOR U919 ( .A(n910), .B(n914), .Z(n912) );
  XNOR U920 ( .A(n846), .B(n841), .Z(n898) );
  AND U921 ( .A(n789), .B(n915), .Z(n841) );
  XOR U922 ( .A(n916), .B(n852), .Z(n846) );
  XNOR U923 ( .A(n917), .B(n918), .Z(n852) );
  NOR U924 ( .A(n919), .B(n920), .Z(n918) );
  XNOR U925 ( .A(n917), .B(n921), .Z(n919) );
  XNOR U926 ( .A(n851), .B(n843), .Z(n916) );
  XOR U927 ( .A(n922), .B(n923), .Z(n843) );
  AND U928 ( .A(n924), .B(n925), .Z(n923) );
  XOR U929 ( .A(n922), .B(n926), .Z(n924) );
  XNOR U930 ( .A(n927), .B(n848), .Z(n851) );
  XOR U931 ( .A(n928), .B(n929), .Z(n848) );
  AND U932 ( .A(n930), .B(n931), .Z(n929) );
  XOR U933 ( .A(n928), .B(n932), .Z(n930) );
  XNOR U934 ( .A(n933), .B(n934), .Z(n927) );
  NOR U935 ( .A(n935), .B(n936), .Z(n934) );
  XOR U936 ( .A(n933), .B(n937), .Z(n935) );
  AND U937 ( .A(n789), .B(n780), .Z(n853) );
  XNOR U938 ( .A(n938), .B(n880), .Z(n780) );
  XOR U939 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(p_input[64]), .Z(n880) );
  XOR U940 ( .A(n868), .B(n867), .Z(n938) );
  XNOR U941 ( .A(n939), .B(n874), .Z(n867) );
  XNOR U942 ( .A(n863), .B(n862), .Z(n874) );
  XOR U943 ( .A(n940), .B(n859), .Z(n862) );
  XOR U944 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(
        p_input[74]), .Z(n859) );
  XOR U945 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n773), .Z(
        n940) );
  XOR U946 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(
        p_input[76]), .Z(n863) );
  XNOR U947 ( .A(n873), .B(n864), .Z(n939) );
  XOR U948 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(p_input[65]), .Z(n864) );
  XOR U949 ( .A(n941), .B(n879), .Z(n873) );
  XNOR U950 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(
        p_input[79]), .Z(n879) );
  XOR U951 ( .A(n870), .B(n878), .Z(n941) );
  XOR U952 ( .A(n942), .B(n875), .Z(n878) );
  XOR U953 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(
        p_input[77]), .Z(n875) );
  XOR U954 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n776), .Z(
        n942) );
  XOR U955 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .B(p_input[73]), .Z(n870) );
  XNOR U956 ( .A(n886), .B(n885), .Z(n868) );
  XNOR U957 ( .A(n943), .B(n891), .Z(n885) );
  XOR U958 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(p_input[72]), .Z(n891) );
  XOR U959 ( .A(n882), .B(n890), .Z(n943) );
  XOR U960 ( .A(n944), .B(n887), .Z(n890) );
  XOR U961 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(p_input[70]), .Z(n887) );
  XNOR U962 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(
        p_input[71]), .Z(n944) );
  XOR U963 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(p_input[66]), .Z(n882) );
  XNOR U964 ( .A(n896), .B(n895), .Z(n886) );
  XOR U965 ( .A(n945), .B(n892), .Z(n895) );
  XOR U966 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(p_input[67]), .Z(n892) );
  XNOR U967 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(
        p_input[68]), .Z(n945) );
  XOR U968 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(p_input[69]), .Z(n896) );
  XOR U969 ( .A(n946), .B(n926), .Z(n789) );
  XOR U970 ( .A(n904), .B(n903), .Z(n926) );
  XNOR U971 ( .A(n947), .B(n909), .Z(n903) );
  XOR U972 ( .A(\knn_comb_/min_val_out[0][8] ), .B(p_input[72]), .Z(n909) );
  XOR U973 ( .A(n900), .B(n908), .Z(n947) );
  XOR U974 ( .A(n948), .B(n905), .Z(n908) );
  XOR U975 ( .A(\knn_comb_/min_val_out[0][6] ), .B(p_input[70]), .Z(n905) );
  XNOR U976 ( .A(\knn_comb_/min_val_out[0][7] ), .B(p_input[71]), .Z(n948) );
  XOR U977 ( .A(\knn_comb_/min_val_out[0][2] ), .B(p_input[66]), .Z(n900) );
  XNOR U978 ( .A(n914), .B(n913), .Z(n904) );
  XOR U979 ( .A(n949), .B(n910), .Z(n913) );
  XOR U980 ( .A(\knn_comb_/min_val_out[0][3] ), .B(p_input[67]), .Z(n910) );
  XNOR U981 ( .A(\knn_comb_/min_val_out[0][4] ), .B(p_input[68]), .Z(n949) );
  XOR U982 ( .A(\knn_comb_/min_val_out[0][5] ), .B(p_input[69]), .Z(n914) );
  XNOR U983 ( .A(n925), .B(n915), .Z(n946) );
  XOR U984 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[64]), .Z(n915) );
  XNOR U985 ( .A(n950), .B(n932), .Z(n925) );
  XNOR U986 ( .A(n921), .B(n920), .Z(n932) );
  XOR U987 ( .A(n951), .B(n917), .Z(n920) );
  XOR U988 ( .A(\knn_comb_/min_val_out[0][10] ), .B(p_input[74]), .Z(n917) );
  XOR U989 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n773), .Z(n951) );
  IV U990 ( .A(p_input[75]), .Z(n773) );
  XOR U991 ( .A(\knn_comb_/min_val_out[0][12] ), .B(p_input[76]), .Z(n921) );
  XNOR U992 ( .A(n931), .B(n922), .Z(n950) );
  XOR U993 ( .A(\knn_comb_/min_val_out[0][1] ), .B(p_input[65]), .Z(n922) );
  XOR U994 ( .A(n952), .B(n937), .Z(n931) );
  XNOR U995 ( .A(\knn_comb_/min_val_out[0][15] ), .B(p_input[79]), .Z(n937) );
  XOR U996 ( .A(n928), .B(n936), .Z(n952) );
  XOR U997 ( .A(n953), .B(n933), .Z(n936) );
  XOR U998 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[77]), .Z(n933) );
  XOR U999 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n776), .Z(n953) );
  IV U1000 ( .A(p_input[78]), .Z(n776) );
  XOR U1001 ( .A(\knn_comb_/min_val_out[0][9] ), .B(p_input[73]), .Z(n928) );
endmodule

