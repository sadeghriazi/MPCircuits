
module auction_BMR_N3_W32 ( p_input, o );
  input [255:0] p_input;
  output [34:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613;

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(o[2]), .B(n3), .Z(n1) );
  XOR U3 ( .A(n2), .B(n4), .Z(n3) );
  XOR U4 ( .A(n5), .B(n6), .Z(o[8]) );
  AND U5 ( .A(o[2]), .B(n7), .Z(n5) );
  XOR U6 ( .A(n8), .B(n9), .Z(n7) );
  XOR U7 ( .A(n10), .B(n11), .Z(o[7]) );
  AND U8 ( .A(o[2]), .B(n12), .Z(n10) );
  XOR U9 ( .A(n13), .B(n14), .Z(n12) );
  XOR U10 ( .A(n15), .B(n16), .Z(o[6]) );
  AND U11 ( .A(o[2]), .B(n17), .Z(n15) );
  XOR U12 ( .A(n18), .B(n19), .Z(n17) );
  XOR U13 ( .A(n20), .B(n21), .Z(o[5]) );
  AND U14 ( .A(o[2]), .B(n22), .Z(n20) );
  XOR U15 ( .A(n23), .B(n24), .Z(n22) );
  XOR U16 ( .A(n25), .B(n26), .Z(o[4]) );
  AND U17 ( .A(o[2]), .B(n27), .Z(n25) );
  XOR U18 ( .A(n28), .B(n29), .Z(n27) );
  XNOR U19 ( .A(n30), .B(n31), .Z(o[3]) );
  AND U20 ( .A(o[2]), .B(n32), .Z(n30) );
  XNOR U21 ( .A(n33), .B(n31), .Z(n32) );
  XNOR U22 ( .A(n34), .B(n35), .Z(o[34]) );
  AND U23 ( .A(o[2]), .B(n36), .Z(n34) );
  XOR U24 ( .A(n37), .B(n35), .Z(n36) );
  XOR U25 ( .A(n38), .B(n39), .Z(o[33]) );
  AND U26 ( .A(o[2]), .B(n40), .Z(n38) );
  XOR U27 ( .A(n41), .B(n42), .Z(n40) );
  XOR U28 ( .A(n43), .B(n44), .Z(o[32]) );
  AND U29 ( .A(o[2]), .B(n45), .Z(n43) );
  XOR U30 ( .A(n46), .B(n47), .Z(n45) );
  XOR U31 ( .A(n48), .B(n49), .Z(o[31]) );
  AND U32 ( .A(o[2]), .B(n50), .Z(n48) );
  XOR U33 ( .A(n51), .B(n52), .Z(n50) );
  XOR U34 ( .A(n53), .B(n54), .Z(o[30]) );
  AND U35 ( .A(o[2]), .B(n55), .Z(n53) );
  XOR U36 ( .A(n56), .B(n57), .Z(n55) );
  XOR U37 ( .A(n58), .B(n59), .Z(o[29]) );
  AND U38 ( .A(o[2]), .B(n60), .Z(n58) );
  XOR U39 ( .A(n61), .B(n62), .Z(n60) );
  XOR U40 ( .A(n63), .B(n64), .Z(o[28]) );
  AND U41 ( .A(o[2]), .B(n65), .Z(n63) );
  XOR U42 ( .A(n66), .B(n67), .Z(n65) );
  XOR U43 ( .A(n68), .B(n69), .Z(o[27]) );
  AND U44 ( .A(o[2]), .B(n70), .Z(n68) );
  XOR U45 ( .A(n71), .B(n72), .Z(n70) );
  XOR U46 ( .A(n73), .B(n74), .Z(o[26]) );
  AND U47 ( .A(o[2]), .B(n75), .Z(n73) );
  XOR U48 ( .A(n76), .B(n77), .Z(n75) );
  XOR U49 ( .A(n78), .B(n79), .Z(o[25]) );
  AND U50 ( .A(o[2]), .B(n80), .Z(n78) );
  XOR U51 ( .A(n81), .B(n82), .Z(n80) );
  XOR U52 ( .A(n83), .B(n84), .Z(o[24]) );
  AND U53 ( .A(o[2]), .B(n85), .Z(n83) );
  XOR U54 ( .A(n86), .B(n87), .Z(n85) );
  XOR U55 ( .A(n88), .B(n89), .Z(o[23]) );
  AND U56 ( .A(o[2]), .B(n90), .Z(n88) );
  XOR U57 ( .A(n91), .B(n92), .Z(n90) );
  XOR U58 ( .A(n93), .B(n94), .Z(o[22]) );
  AND U59 ( .A(o[2]), .B(n95), .Z(n93) );
  XOR U60 ( .A(n96), .B(n97), .Z(n95) );
  XOR U61 ( .A(n98), .B(n99), .Z(o[21]) );
  AND U62 ( .A(o[2]), .B(n100), .Z(n98) );
  XOR U63 ( .A(n101), .B(n102), .Z(n100) );
  XOR U64 ( .A(n103), .B(n104), .Z(o[20]) );
  AND U65 ( .A(o[2]), .B(n105), .Z(n103) );
  XOR U66 ( .A(n106), .B(n107), .Z(n105) );
  XOR U67 ( .A(n108), .B(n109), .Z(o[19]) );
  AND U68 ( .A(o[2]), .B(n110), .Z(n108) );
  XOR U69 ( .A(n111), .B(n112), .Z(n110) );
  XOR U70 ( .A(n113), .B(n114), .Z(o[18]) );
  AND U71 ( .A(o[2]), .B(n115), .Z(n113) );
  XOR U72 ( .A(n116), .B(n117), .Z(n115) );
  XOR U73 ( .A(n118), .B(n119), .Z(o[17]) );
  AND U74 ( .A(o[2]), .B(n120), .Z(n118) );
  XOR U75 ( .A(n121), .B(n122), .Z(n120) );
  XOR U76 ( .A(n123), .B(n124), .Z(o[16]) );
  AND U77 ( .A(o[2]), .B(n125), .Z(n123) );
  XOR U78 ( .A(n126), .B(n127), .Z(n125) );
  XOR U79 ( .A(n128), .B(n129), .Z(o[15]) );
  AND U80 ( .A(o[2]), .B(n130), .Z(n128) );
  XOR U81 ( .A(n131), .B(n132), .Z(n130) );
  XOR U82 ( .A(n133), .B(n134), .Z(o[14]) );
  AND U83 ( .A(o[2]), .B(n135), .Z(n133) );
  XOR U84 ( .A(n136), .B(n137), .Z(n135) );
  XOR U85 ( .A(n138), .B(n139), .Z(o[13]) );
  AND U86 ( .A(o[2]), .B(n140), .Z(n138) );
  XOR U87 ( .A(n141), .B(n142), .Z(n140) );
  XOR U88 ( .A(n143), .B(n144), .Z(o[12]) );
  AND U89 ( .A(o[2]), .B(n145), .Z(n143) );
  XOR U90 ( .A(n146), .B(n147), .Z(n145) );
  XOR U91 ( .A(n148), .B(n149), .Z(o[11]) );
  AND U92 ( .A(o[2]), .B(n150), .Z(n148) );
  XOR U93 ( .A(n151), .B(n152), .Z(n150) );
  XOR U94 ( .A(n153), .B(n154), .Z(o[10]) );
  AND U95 ( .A(o[2]), .B(n155), .Z(n153) );
  XOR U96 ( .A(n156), .B(n157), .Z(n155) );
  XOR U97 ( .A(n158), .B(n159), .Z(o[0]) );
  AND U98 ( .A(o[1]), .B(n160), .Z(n159) );
  XNOR U99 ( .A(n158), .B(n161), .Z(n160) );
  XNOR U100 ( .A(n162), .B(n163), .Z(n161) );
  AND U101 ( .A(o[2]), .B(n164), .Z(n162) );
  XOR U102 ( .A(n163), .B(n165), .Z(n164) );
  XOR U103 ( .A(n166), .B(n167), .Z(o[1]) );
  AND U104 ( .A(o[2]), .B(n168), .Z(n167) );
  XOR U105 ( .A(n166), .B(n169), .Z(n168) );
  XOR U106 ( .A(n170), .B(n171), .Z(n158) );
  AND U107 ( .A(o[2]), .B(n172), .Z(n171) );
  XOR U108 ( .A(n170), .B(n173), .Z(n172) );
  XOR U109 ( .A(n174), .B(n175), .Z(o[2]) );
  AND U110 ( .A(n176), .B(n177), .Z(n175) );
  XOR U111 ( .A(n174), .B(n37), .Z(n177) );
  XNOR U112 ( .A(n178), .B(n179), .Z(n37) );
  AND U113 ( .A(n180), .B(n169), .Z(n179) );
  AND U114 ( .A(n178), .B(n181), .Z(n180) );
  XNOR U115 ( .A(n35), .B(n174), .Z(n176) );
  XOR U116 ( .A(n182), .B(n183), .Z(n35) );
  AND U117 ( .A(n184), .B(n166), .Z(n183) );
  NOR U118 ( .A(n182), .B(n185), .Z(n184) );
  XOR U119 ( .A(n186), .B(n187), .Z(n174) );
  AND U120 ( .A(n188), .B(n189), .Z(n187) );
  XOR U121 ( .A(n186), .B(n41), .Z(n189) );
  XOR U122 ( .A(n190), .B(n191), .Z(n41) );
  AND U123 ( .A(n169), .B(n192), .Z(n191) );
  XOR U124 ( .A(n193), .B(n190), .Z(n192) );
  XNOR U125 ( .A(n42), .B(n186), .Z(n188) );
  IV U126 ( .A(n39), .Z(n42) );
  XNOR U127 ( .A(n194), .B(n195), .Z(n39) );
  AND U128 ( .A(n166), .B(n196), .Z(n195) );
  XOR U129 ( .A(n197), .B(n194), .Z(n196) );
  XOR U130 ( .A(n198), .B(n199), .Z(n186) );
  AND U131 ( .A(n200), .B(n201), .Z(n199) );
  XOR U132 ( .A(n198), .B(n46), .Z(n201) );
  XOR U133 ( .A(n202), .B(n203), .Z(n46) );
  AND U134 ( .A(n169), .B(n204), .Z(n203) );
  XOR U135 ( .A(n205), .B(n202), .Z(n204) );
  XNOR U136 ( .A(n47), .B(n198), .Z(n200) );
  IV U137 ( .A(n44), .Z(n47) );
  XNOR U138 ( .A(n206), .B(n207), .Z(n44) );
  AND U139 ( .A(n166), .B(n208), .Z(n207) );
  XOR U140 ( .A(n209), .B(n206), .Z(n208) );
  XOR U141 ( .A(n210), .B(n211), .Z(n198) );
  AND U142 ( .A(n212), .B(n213), .Z(n211) );
  XOR U143 ( .A(n210), .B(n51), .Z(n213) );
  XOR U144 ( .A(n214), .B(n215), .Z(n51) );
  AND U145 ( .A(n169), .B(n216), .Z(n215) );
  XOR U146 ( .A(n217), .B(n214), .Z(n216) );
  XNOR U147 ( .A(n52), .B(n210), .Z(n212) );
  IV U148 ( .A(n49), .Z(n52) );
  XNOR U149 ( .A(n218), .B(n219), .Z(n49) );
  AND U150 ( .A(n166), .B(n220), .Z(n219) );
  XOR U151 ( .A(n221), .B(n218), .Z(n220) );
  XOR U152 ( .A(n222), .B(n223), .Z(n210) );
  AND U153 ( .A(n224), .B(n225), .Z(n223) );
  XOR U154 ( .A(n222), .B(n56), .Z(n225) );
  XOR U155 ( .A(n226), .B(n227), .Z(n56) );
  AND U156 ( .A(n169), .B(n228), .Z(n227) );
  XOR U157 ( .A(n229), .B(n226), .Z(n228) );
  XNOR U158 ( .A(n57), .B(n222), .Z(n224) );
  IV U159 ( .A(n54), .Z(n57) );
  XNOR U160 ( .A(n230), .B(n231), .Z(n54) );
  AND U161 ( .A(n166), .B(n232), .Z(n231) );
  XOR U162 ( .A(n233), .B(n230), .Z(n232) );
  XOR U163 ( .A(n234), .B(n235), .Z(n222) );
  AND U164 ( .A(n236), .B(n237), .Z(n235) );
  XOR U165 ( .A(n234), .B(n61), .Z(n237) );
  XOR U166 ( .A(n238), .B(n239), .Z(n61) );
  AND U167 ( .A(n169), .B(n240), .Z(n239) );
  XOR U168 ( .A(n241), .B(n238), .Z(n240) );
  XNOR U169 ( .A(n62), .B(n234), .Z(n236) );
  IV U170 ( .A(n59), .Z(n62) );
  XNOR U171 ( .A(n242), .B(n243), .Z(n59) );
  AND U172 ( .A(n166), .B(n244), .Z(n243) );
  XOR U173 ( .A(n245), .B(n242), .Z(n244) );
  XOR U174 ( .A(n246), .B(n247), .Z(n234) );
  AND U175 ( .A(n248), .B(n249), .Z(n247) );
  XOR U176 ( .A(n246), .B(n66), .Z(n249) );
  XOR U177 ( .A(n250), .B(n251), .Z(n66) );
  AND U178 ( .A(n169), .B(n252), .Z(n251) );
  XOR U179 ( .A(n253), .B(n250), .Z(n252) );
  XNOR U180 ( .A(n67), .B(n246), .Z(n248) );
  IV U181 ( .A(n64), .Z(n67) );
  XNOR U182 ( .A(n254), .B(n255), .Z(n64) );
  AND U183 ( .A(n166), .B(n256), .Z(n255) );
  XOR U184 ( .A(n257), .B(n254), .Z(n256) );
  XOR U185 ( .A(n258), .B(n259), .Z(n246) );
  AND U186 ( .A(n260), .B(n261), .Z(n259) );
  XOR U187 ( .A(n258), .B(n71), .Z(n261) );
  XOR U188 ( .A(n262), .B(n263), .Z(n71) );
  AND U189 ( .A(n169), .B(n264), .Z(n263) );
  XOR U190 ( .A(n265), .B(n262), .Z(n264) );
  XNOR U191 ( .A(n72), .B(n258), .Z(n260) );
  IV U192 ( .A(n69), .Z(n72) );
  XNOR U193 ( .A(n266), .B(n267), .Z(n69) );
  AND U194 ( .A(n166), .B(n268), .Z(n267) );
  XOR U195 ( .A(n269), .B(n266), .Z(n268) );
  XOR U196 ( .A(n270), .B(n271), .Z(n258) );
  AND U197 ( .A(n272), .B(n273), .Z(n271) );
  XOR U198 ( .A(n270), .B(n76), .Z(n273) );
  XOR U199 ( .A(n274), .B(n275), .Z(n76) );
  AND U200 ( .A(n169), .B(n276), .Z(n275) );
  XOR U201 ( .A(n277), .B(n274), .Z(n276) );
  XNOR U202 ( .A(n77), .B(n270), .Z(n272) );
  IV U203 ( .A(n74), .Z(n77) );
  XNOR U204 ( .A(n278), .B(n279), .Z(n74) );
  AND U205 ( .A(n166), .B(n280), .Z(n279) );
  XOR U206 ( .A(n281), .B(n278), .Z(n280) );
  XOR U207 ( .A(n282), .B(n283), .Z(n270) );
  AND U208 ( .A(n284), .B(n285), .Z(n283) );
  XOR U209 ( .A(n282), .B(n81), .Z(n285) );
  XOR U210 ( .A(n286), .B(n287), .Z(n81) );
  AND U211 ( .A(n169), .B(n288), .Z(n287) );
  XOR U212 ( .A(n289), .B(n286), .Z(n288) );
  XNOR U213 ( .A(n82), .B(n282), .Z(n284) );
  IV U214 ( .A(n79), .Z(n82) );
  XNOR U215 ( .A(n290), .B(n291), .Z(n79) );
  AND U216 ( .A(n166), .B(n292), .Z(n291) );
  XOR U217 ( .A(n293), .B(n290), .Z(n292) );
  XOR U218 ( .A(n294), .B(n295), .Z(n282) );
  AND U219 ( .A(n296), .B(n297), .Z(n295) );
  XOR U220 ( .A(n294), .B(n86), .Z(n297) );
  XOR U221 ( .A(n298), .B(n299), .Z(n86) );
  AND U222 ( .A(n169), .B(n300), .Z(n299) );
  XOR U223 ( .A(n301), .B(n298), .Z(n300) );
  XNOR U224 ( .A(n87), .B(n294), .Z(n296) );
  IV U225 ( .A(n84), .Z(n87) );
  XNOR U226 ( .A(n302), .B(n303), .Z(n84) );
  AND U227 ( .A(n166), .B(n304), .Z(n303) );
  XOR U228 ( .A(n305), .B(n302), .Z(n304) );
  XOR U229 ( .A(n306), .B(n307), .Z(n294) );
  AND U230 ( .A(n308), .B(n309), .Z(n307) );
  XOR U231 ( .A(n306), .B(n91), .Z(n309) );
  XOR U232 ( .A(n310), .B(n311), .Z(n91) );
  AND U233 ( .A(n169), .B(n312), .Z(n311) );
  XOR U234 ( .A(n313), .B(n310), .Z(n312) );
  XNOR U235 ( .A(n92), .B(n306), .Z(n308) );
  IV U236 ( .A(n89), .Z(n92) );
  XNOR U237 ( .A(n314), .B(n315), .Z(n89) );
  AND U238 ( .A(n166), .B(n316), .Z(n315) );
  XOR U239 ( .A(n317), .B(n314), .Z(n316) );
  XOR U240 ( .A(n318), .B(n319), .Z(n306) );
  AND U241 ( .A(n320), .B(n321), .Z(n319) );
  XOR U242 ( .A(n318), .B(n96), .Z(n321) );
  XOR U243 ( .A(n322), .B(n323), .Z(n96) );
  AND U244 ( .A(n169), .B(n324), .Z(n323) );
  XOR U245 ( .A(n325), .B(n322), .Z(n324) );
  XNOR U246 ( .A(n97), .B(n318), .Z(n320) );
  IV U247 ( .A(n94), .Z(n97) );
  XNOR U248 ( .A(n326), .B(n327), .Z(n94) );
  AND U249 ( .A(n166), .B(n328), .Z(n327) );
  XOR U250 ( .A(n329), .B(n326), .Z(n328) );
  XOR U251 ( .A(n330), .B(n331), .Z(n318) );
  AND U252 ( .A(n332), .B(n333), .Z(n331) );
  XOR U253 ( .A(n330), .B(n101), .Z(n333) );
  XOR U254 ( .A(n334), .B(n335), .Z(n101) );
  AND U255 ( .A(n169), .B(n336), .Z(n335) );
  XOR U256 ( .A(n337), .B(n334), .Z(n336) );
  XNOR U257 ( .A(n102), .B(n330), .Z(n332) );
  IV U258 ( .A(n99), .Z(n102) );
  XNOR U259 ( .A(n338), .B(n339), .Z(n99) );
  AND U260 ( .A(n166), .B(n340), .Z(n339) );
  XOR U261 ( .A(n341), .B(n338), .Z(n340) );
  XOR U262 ( .A(n342), .B(n343), .Z(n330) );
  AND U263 ( .A(n344), .B(n345), .Z(n343) );
  XOR U264 ( .A(n342), .B(n106), .Z(n345) );
  XOR U265 ( .A(n346), .B(n347), .Z(n106) );
  AND U266 ( .A(n169), .B(n348), .Z(n347) );
  XOR U267 ( .A(n349), .B(n346), .Z(n348) );
  XNOR U268 ( .A(n107), .B(n342), .Z(n344) );
  IV U269 ( .A(n104), .Z(n107) );
  XNOR U270 ( .A(n350), .B(n351), .Z(n104) );
  AND U271 ( .A(n166), .B(n352), .Z(n351) );
  XOR U272 ( .A(n353), .B(n350), .Z(n352) );
  XOR U273 ( .A(n354), .B(n355), .Z(n342) );
  AND U274 ( .A(n356), .B(n357), .Z(n355) );
  XOR U275 ( .A(n354), .B(n111), .Z(n357) );
  XOR U276 ( .A(n358), .B(n359), .Z(n111) );
  AND U277 ( .A(n169), .B(n360), .Z(n359) );
  XOR U278 ( .A(n361), .B(n358), .Z(n360) );
  XNOR U279 ( .A(n112), .B(n354), .Z(n356) );
  IV U280 ( .A(n109), .Z(n112) );
  XNOR U281 ( .A(n362), .B(n363), .Z(n109) );
  AND U282 ( .A(n166), .B(n364), .Z(n363) );
  XOR U283 ( .A(n365), .B(n362), .Z(n364) );
  XOR U284 ( .A(n366), .B(n367), .Z(n354) );
  AND U285 ( .A(n368), .B(n369), .Z(n367) );
  XOR U286 ( .A(n366), .B(n116), .Z(n369) );
  XOR U287 ( .A(n370), .B(n371), .Z(n116) );
  AND U288 ( .A(n169), .B(n372), .Z(n371) );
  XOR U289 ( .A(n373), .B(n370), .Z(n372) );
  XNOR U290 ( .A(n117), .B(n366), .Z(n368) );
  IV U291 ( .A(n114), .Z(n117) );
  XNOR U292 ( .A(n374), .B(n375), .Z(n114) );
  AND U293 ( .A(n166), .B(n376), .Z(n375) );
  XOR U294 ( .A(n377), .B(n374), .Z(n376) );
  XOR U295 ( .A(n378), .B(n379), .Z(n366) );
  AND U296 ( .A(n380), .B(n381), .Z(n379) );
  XOR U297 ( .A(n378), .B(n121), .Z(n381) );
  XOR U298 ( .A(n382), .B(n383), .Z(n121) );
  AND U299 ( .A(n169), .B(n384), .Z(n383) );
  XOR U300 ( .A(n385), .B(n382), .Z(n384) );
  XNOR U301 ( .A(n122), .B(n378), .Z(n380) );
  IV U302 ( .A(n119), .Z(n122) );
  XNOR U303 ( .A(n386), .B(n387), .Z(n119) );
  AND U304 ( .A(n166), .B(n388), .Z(n387) );
  XOR U305 ( .A(n389), .B(n386), .Z(n388) );
  XOR U306 ( .A(n390), .B(n391), .Z(n378) );
  AND U307 ( .A(n392), .B(n393), .Z(n391) );
  XOR U308 ( .A(n390), .B(n126), .Z(n393) );
  XOR U309 ( .A(n394), .B(n395), .Z(n126) );
  AND U310 ( .A(n169), .B(n396), .Z(n395) );
  XOR U311 ( .A(n397), .B(n394), .Z(n396) );
  XNOR U312 ( .A(n127), .B(n390), .Z(n392) );
  IV U313 ( .A(n124), .Z(n127) );
  XNOR U314 ( .A(n398), .B(n399), .Z(n124) );
  AND U315 ( .A(n166), .B(n400), .Z(n399) );
  XOR U316 ( .A(n401), .B(n398), .Z(n400) );
  XOR U317 ( .A(n402), .B(n403), .Z(n390) );
  AND U318 ( .A(n404), .B(n405), .Z(n403) );
  XOR U319 ( .A(n402), .B(n131), .Z(n405) );
  XOR U320 ( .A(n406), .B(n407), .Z(n131) );
  AND U321 ( .A(n169), .B(n408), .Z(n407) );
  XOR U322 ( .A(n409), .B(n406), .Z(n408) );
  XNOR U323 ( .A(n132), .B(n402), .Z(n404) );
  IV U324 ( .A(n129), .Z(n132) );
  XNOR U325 ( .A(n410), .B(n411), .Z(n129) );
  AND U326 ( .A(n166), .B(n412), .Z(n411) );
  XOR U327 ( .A(n413), .B(n410), .Z(n412) );
  XOR U328 ( .A(n414), .B(n415), .Z(n402) );
  AND U329 ( .A(n416), .B(n417), .Z(n415) );
  XOR U330 ( .A(n414), .B(n136), .Z(n417) );
  XOR U331 ( .A(n418), .B(n419), .Z(n136) );
  AND U332 ( .A(n169), .B(n420), .Z(n419) );
  XOR U333 ( .A(n421), .B(n418), .Z(n420) );
  XNOR U334 ( .A(n137), .B(n414), .Z(n416) );
  IV U335 ( .A(n134), .Z(n137) );
  XNOR U336 ( .A(n422), .B(n423), .Z(n134) );
  AND U337 ( .A(n166), .B(n424), .Z(n423) );
  XOR U338 ( .A(n425), .B(n422), .Z(n424) );
  XOR U339 ( .A(n426), .B(n427), .Z(n414) );
  AND U340 ( .A(n428), .B(n429), .Z(n427) );
  XOR U341 ( .A(n426), .B(n141), .Z(n429) );
  XOR U342 ( .A(n430), .B(n431), .Z(n141) );
  AND U343 ( .A(n169), .B(n432), .Z(n431) );
  XOR U344 ( .A(n433), .B(n430), .Z(n432) );
  XNOR U345 ( .A(n142), .B(n426), .Z(n428) );
  IV U346 ( .A(n139), .Z(n142) );
  XNOR U347 ( .A(n434), .B(n435), .Z(n139) );
  AND U348 ( .A(n166), .B(n436), .Z(n435) );
  XOR U349 ( .A(n437), .B(n434), .Z(n436) );
  XOR U350 ( .A(n438), .B(n439), .Z(n426) );
  AND U351 ( .A(n440), .B(n441), .Z(n439) );
  XOR U352 ( .A(n438), .B(n146), .Z(n441) );
  XOR U353 ( .A(n442), .B(n443), .Z(n146) );
  AND U354 ( .A(n169), .B(n444), .Z(n443) );
  XOR U355 ( .A(n445), .B(n442), .Z(n444) );
  XNOR U356 ( .A(n147), .B(n438), .Z(n440) );
  IV U357 ( .A(n144), .Z(n147) );
  XNOR U358 ( .A(n446), .B(n447), .Z(n144) );
  AND U359 ( .A(n166), .B(n448), .Z(n447) );
  XOR U360 ( .A(n449), .B(n446), .Z(n448) );
  XOR U361 ( .A(n450), .B(n451), .Z(n438) );
  AND U362 ( .A(n452), .B(n453), .Z(n451) );
  XOR U363 ( .A(n450), .B(n151), .Z(n453) );
  XOR U364 ( .A(n454), .B(n455), .Z(n151) );
  AND U365 ( .A(n169), .B(n456), .Z(n455) );
  XOR U366 ( .A(n457), .B(n454), .Z(n456) );
  XNOR U367 ( .A(n152), .B(n450), .Z(n452) );
  IV U368 ( .A(n149), .Z(n152) );
  XNOR U369 ( .A(n458), .B(n459), .Z(n149) );
  AND U370 ( .A(n166), .B(n460), .Z(n459) );
  XOR U371 ( .A(n461), .B(n458), .Z(n460) );
  XOR U372 ( .A(n462), .B(n463), .Z(n450) );
  AND U373 ( .A(n464), .B(n465), .Z(n463) );
  XOR U374 ( .A(n462), .B(n156), .Z(n465) );
  XOR U375 ( .A(n466), .B(n467), .Z(n156) );
  AND U376 ( .A(n169), .B(n468), .Z(n467) );
  XOR U377 ( .A(n469), .B(n466), .Z(n468) );
  XNOR U378 ( .A(n157), .B(n462), .Z(n464) );
  IV U379 ( .A(n154), .Z(n157) );
  XNOR U380 ( .A(n470), .B(n471), .Z(n154) );
  AND U381 ( .A(n166), .B(n472), .Z(n471) );
  XOR U382 ( .A(n473), .B(n470), .Z(n472) );
  XOR U383 ( .A(n474), .B(n475), .Z(n462) );
  AND U384 ( .A(n476), .B(n477), .Z(n475) );
  XOR U385 ( .A(n4), .B(n474), .Z(n477) );
  XOR U386 ( .A(n478), .B(n479), .Z(n4) );
  AND U387 ( .A(n169), .B(n480), .Z(n479) );
  XOR U388 ( .A(n478), .B(n481), .Z(n480) );
  XNOR U389 ( .A(n474), .B(n2), .Z(n476) );
  XOR U390 ( .A(n482), .B(n483), .Z(n2) );
  AND U391 ( .A(n166), .B(n484), .Z(n483) );
  XOR U392 ( .A(n482), .B(n485), .Z(n484) );
  XOR U393 ( .A(n486), .B(n487), .Z(n474) );
  AND U394 ( .A(n488), .B(n489), .Z(n487) );
  XOR U395 ( .A(n486), .B(n8), .Z(n489) );
  XOR U396 ( .A(n490), .B(n491), .Z(n8) );
  AND U397 ( .A(n169), .B(n492), .Z(n491) );
  XOR U398 ( .A(n493), .B(n490), .Z(n492) );
  XNOR U399 ( .A(n9), .B(n486), .Z(n488) );
  IV U400 ( .A(n6), .Z(n9) );
  XNOR U401 ( .A(n494), .B(n495), .Z(n6) );
  AND U402 ( .A(n166), .B(n496), .Z(n495) );
  XOR U403 ( .A(n497), .B(n494), .Z(n496) );
  XOR U404 ( .A(n498), .B(n499), .Z(n486) );
  AND U405 ( .A(n500), .B(n501), .Z(n499) );
  XOR U406 ( .A(n498), .B(n13), .Z(n501) );
  XOR U407 ( .A(n502), .B(n503), .Z(n13) );
  AND U408 ( .A(n169), .B(n504), .Z(n503) );
  XOR U409 ( .A(n505), .B(n502), .Z(n504) );
  XNOR U410 ( .A(n14), .B(n498), .Z(n500) );
  IV U411 ( .A(n11), .Z(n14) );
  XNOR U412 ( .A(n506), .B(n507), .Z(n11) );
  AND U413 ( .A(n166), .B(n508), .Z(n507) );
  XOR U414 ( .A(n509), .B(n506), .Z(n508) );
  XOR U415 ( .A(n510), .B(n511), .Z(n498) );
  AND U416 ( .A(n512), .B(n513), .Z(n511) );
  XOR U417 ( .A(n510), .B(n18), .Z(n513) );
  XOR U418 ( .A(n514), .B(n515), .Z(n18) );
  AND U419 ( .A(n169), .B(n516), .Z(n515) );
  XOR U420 ( .A(n517), .B(n514), .Z(n516) );
  XNOR U421 ( .A(n19), .B(n510), .Z(n512) );
  IV U422 ( .A(n16), .Z(n19) );
  XNOR U423 ( .A(n518), .B(n519), .Z(n16) );
  AND U424 ( .A(n166), .B(n520), .Z(n519) );
  XOR U425 ( .A(n521), .B(n518), .Z(n520) );
  XOR U426 ( .A(n522), .B(n523), .Z(n510) );
  AND U427 ( .A(n524), .B(n525), .Z(n523) );
  XOR U428 ( .A(n522), .B(n23), .Z(n525) );
  XOR U429 ( .A(n526), .B(n527), .Z(n23) );
  AND U430 ( .A(n169), .B(n528), .Z(n527) );
  XOR U431 ( .A(n529), .B(n526), .Z(n528) );
  XNOR U432 ( .A(n24), .B(n522), .Z(n524) );
  IV U433 ( .A(n21), .Z(n24) );
  XNOR U434 ( .A(n530), .B(n531), .Z(n21) );
  AND U435 ( .A(n166), .B(n532), .Z(n531) );
  XOR U436 ( .A(n533), .B(n530), .Z(n532) );
  XNOR U437 ( .A(n534), .B(n535), .Z(n522) );
  AND U438 ( .A(n536), .B(n537), .Z(n535) );
  XNOR U439 ( .A(n534), .B(n28), .Z(n537) );
  XOR U440 ( .A(n538), .B(n539), .Z(n28) );
  AND U441 ( .A(n169), .B(n540), .Z(n539) );
  XOR U442 ( .A(n541), .B(n538), .Z(n540) );
  XOR U443 ( .A(n29), .B(n534), .Z(n536) );
  IV U444 ( .A(n26), .Z(n29) );
  XNOR U445 ( .A(n542), .B(n543), .Z(n26) );
  AND U446 ( .A(n166), .B(n544), .Z(n543) );
  XOR U447 ( .A(n545), .B(n542), .Z(n544) );
  AND U448 ( .A(n31), .B(n33), .Z(n534) );
  XNOR U449 ( .A(n546), .B(n547), .Z(n33) );
  AND U450 ( .A(n169), .B(n548), .Z(n547) );
  XNOR U451 ( .A(n549), .B(n546), .Z(n548) );
  XOR U452 ( .A(n550), .B(n551), .Z(n169) );
  AND U453 ( .A(n552), .B(n553), .Z(n551) );
  XOR U454 ( .A(n181), .B(n550), .Z(n553) );
  IV U455 ( .A(n554), .Z(n181) );
  AND U456 ( .A(p_input[255]), .B(p_input[223]), .Z(n554) );
  XOR U457 ( .A(n550), .B(n178), .Z(n552) );
  AND U458 ( .A(p_input[159]), .B(p_input[191]), .Z(n178) );
  XOR U459 ( .A(n555), .B(n556), .Z(n550) );
  AND U460 ( .A(n557), .B(n558), .Z(n556) );
  XOR U461 ( .A(n555), .B(n193), .Z(n558) );
  XNOR U462 ( .A(p_input[222]), .B(n559), .Z(n193) );
  AND U463 ( .A(n165), .B(n560), .Z(n559) );
  XOR U464 ( .A(p_input[254]), .B(p_input[222]), .Z(n560) );
  XNOR U465 ( .A(n190), .B(n555), .Z(n557) );
  XOR U466 ( .A(n561), .B(n562), .Z(n190) );
  AND U467 ( .A(n163), .B(n563), .Z(n562) );
  XOR U468 ( .A(p_input[190]), .B(p_input[158]), .Z(n563) );
  XOR U469 ( .A(n564), .B(n565), .Z(n555) );
  AND U470 ( .A(n566), .B(n567), .Z(n565) );
  XOR U471 ( .A(n564), .B(n205), .Z(n567) );
  XNOR U472 ( .A(p_input[221]), .B(n568), .Z(n205) );
  AND U473 ( .A(n165), .B(n569), .Z(n568) );
  XOR U474 ( .A(p_input[253]), .B(p_input[221]), .Z(n569) );
  XNOR U475 ( .A(n202), .B(n564), .Z(n566) );
  XOR U476 ( .A(n570), .B(n571), .Z(n202) );
  AND U477 ( .A(n163), .B(n572), .Z(n571) );
  XOR U478 ( .A(p_input[189]), .B(p_input[157]), .Z(n572) );
  XOR U479 ( .A(n573), .B(n574), .Z(n564) );
  AND U480 ( .A(n575), .B(n576), .Z(n574) );
  XOR U481 ( .A(n573), .B(n217), .Z(n576) );
  XNOR U482 ( .A(p_input[220]), .B(n577), .Z(n217) );
  AND U483 ( .A(n165), .B(n578), .Z(n577) );
  XOR U484 ( .A(p_input[252]), .B(p_input[220]), .Z(n578) );
  XNOR U485 ( .A(n214), .B(n573), .Z(n575) );
  XOR U486 ( .A(n579), .B(n580), .Z(n214) );
  AND U487 ( .A(n163), .B(n581), .Z(n580) );
  XOR U488 ( .A(p_input[188]), .B(p_input[156]), .Z(n581) );
  XOR U489 ( .A(n582), .B(n583), .Z(n573) );
  AND U490 ( .A(n584), .B(n585), .Z(n583) );
  XOR U491 ( .A(n582), .B(n229), .Z(n585) );
  XNOR U492 ( .A(p_input[219]), .B(n586), .Z(n229) );
  AND U493 ( .A(n165), .B(n587), .Z(n586) );
  XOR U494 ( .A(p_input[251]), .B(p_input[219]), .Z(n587) );
  XNOR U495 ( .A(n226), .B(n582), .Z(n584) );
  XOR U496 ( .A(n588), .B(n589), .Z(n226) );
  AND U497 ( .A(n163), .B(n590), .Z(n589) );
  XOR U498 ( .A(p_input[187]), .B(p_input[155]), .Z(n590) );
  XOR U499 ( .A(n591), .B(n592), .Z(n582) );
  AND U500 ( .A(n593), .B(n594), .Z(n592) );
  XOR U501 ( .A(n591), .B(n241), .Z(n594) );
  XNOR U502 ( .A(p_input[218]), .B(n595), .Z(n241) );
  AND U503 ( .A(n165), .B(n596), .Z(n595) );
  XOR U504 ( .A(p_input[250]), .B(p_input[218]), .Z(n596) );
  XNOR U505 ( .A(n238), .B(n591), .Z(n593) );
  XOR U506 ( .A(n597), .B(n598), .Z(n238) );
  AND U507 ( .A(n163), .B(n599), .Z(n598) );
  XOR U508 ( .A(p_input[186]), .B(p_input[154]), .Z(n599) );
  XOR U509 ( .A(n600), .B(n601), .Z(n591) );
  AND U510 ( .A(n602), .B(n603), .Z(n601) );
  XOR U511 ( .A(n600), .B(n253), .Z(n603) );
  XNOR U512 ( .A(p_input[217]), .B(n604), .Z(n253) );
  AND U513 ( .A(n165), .B(n605), .Z(n604) );
  XOR U514 ( .A(p_input[249]), .B(p_input[217]), .Z(n605) );
  XNOR U515 ( .A(n250), .B(n600), .Z(n602) );
  XOR U516 ( .A(n606), .B(n607), .Z(n250) );
  AND U517 ( .A(n163), .B(n608), .Z(n607) );
  XOR U518 ( .A(p_input[185]), .B(p_input[153]), .Z(n608) );
  XOR U519 ( .A(n609), .B(n610), .Z(n600) );
  AND U520 ( .A(n611), .B(n612), .Z(n610) );
  XOR U521 ( .A(n609), .B(n265), .Z(n612) );
  XNOR U522 ( .A(p_input[216]), .B(n613), .Z(n265) );
  AND U523 ( .A(n165), .B(n614), .Z(n613) );
  XOR U524 ( .A(p_input[248]), .B(p_input[216]), .Z(n614) );
  XNOR U525 ( .A(n262), .B(n609), .Z(n611) );
  XOR U526 ( .A(n615), .B(n616), .Z(n262) );
  AND U527 ( .A(n163), .B(n617), .Z(n616) );
  XOR U528 ( .A(p_input[184]), .B(p_input[152]), .Z(n617) );
  XOR U529 ( .A(n618), .B(n619), .Z(n609) );
  AND U530 ( .A(n620), .B(n621), .Z(n619) );
  XOR U531 ( .A(n618), .B(n277), .Z(n621) );
  XNOR U532 ( .A(p_input[215]), .B(n622), .Z(n277) );
  AND U533 ( .A(n165), .B(n623), .Z(n622) );
  XOR U534 ( .A(p_input[247]), .B(p_input[215]), .Z(n623) );
  XNOR U535 ( .A(n274), .B(n618), .Z(n620) );
  XOR U536 ( .A(n624), .B(n625), .Z(n274) );
  AND U537 ( .A(n163), .B(n626), .Z(n625) );
  XOR U538 ( .A(p_input[183]), .B(p_input[151]), .Z(n626) );
  XOR U539 ( .A(n627), .B(n628), .Z(n618) );
  AND U540 ( .A(n629), .B(n630), .Z(n628) );
  XOR U541 ( .A(n627), .B(n289), .Z(n630) );
  XNOR U542 ( .A(p_input[214]), .B(n631), .Z(n289) );
  AND U543 ( .A(n165), .B(n632), .Z(n631) );
  XOR U544 ( .A(p_input[246]), .B(p_input[214]), .Z(n632) );
  XNOR U545 ( .A(n286), .B(n627), .Z(n629) );
  XOR U546 ( .A(n633), .B(n634), .Z(n286) );
  AND U547 ( .A(n163), .B(n635), .Z(n634) );
  XOR U548 ( .A(p_input[182]), .B(p_input[150]), .Z(n635) );
  XOR U549 ( .A(n636), .B(n637), .Z(n627) );
  AND U550 ( .A(n638), .B(n639), .Z(n637) );
  XOR U551 ( .A(n636), .B(n301), .Z(n639) );
  XNOR U552 ( .A(p_input[213]), .B(n640), .Z(n301) );
  AND U553 ( .A(n165), .B(n641), .Z(n640) );
  XOR U554 ( .A(p_input[245]), .B(p_input[213]), .Z(n641) );
  XNOR U555 ( .A(n298), .B(n636), .Z(n638) );
  XOR U556 ( .A(n642), .B(n643), .Z(n298) );
  AND U557 ( .A(n163), .B(n644), .Z(n643) );
  XOR U558 ( .A(p_input[181]), .B(p_input[149]), .Z(n644) );
  XOR U559 ( .A(n645), .B(n646), .Z(n636) );
  AND U560 ( .A(n647), .B(n648), .Z(n646) );
  XOR U561 ( .A(n645), .B(n313), .Z(n648) );
  XNOR U562 ( .A(p_input[212]), .B(n649), .Z(n313) );
  AND U563 ( .A(n165), .B(n650), .Z(n649) );
  XOR U564 ( .A(p_input[244]), .B(p_input[212]), .Z(n650) );
  XNOR U565 ( .A(n310), .B(n645), .Z(n647) );
  XOR U566 ( .A(n651), .B(n652), .Z(n310) );
  AND U567 ( .A(n163), .B(n653), .Z(n652) );
  XOR U568 ( .A(p_input[180]), .B(p_input[148]), .Z(n653) );
  XOR U569 ( .A(n654), .B(n655), .Z(n645) );
  AND U570 ( .A(n656), .B(n657), .Z(n655) );
  XOR U571 ( .A(n654), .B(n325), .Z(n657) );
  XNOR U572 ( .A(p_input[211]), .B(n658), .Z(n325) );
  AND U573 ( .A(n165), .B(n659), .Z(n658) );
  XOR U574 ( .A(p_input[243]), .B(p_input[211]), .Z(n659) );
  XNOR U575 ( .A(n322), .B(n654), .Z(n656) );
  XOR U576 ( .A(n660), .B(n661), .Z(n322) );
  AND U577 ( .A(n163), .B(n662), .Z(n661) );
  XOR U578 ( .A(p_input[179]), .B(p_input[147]), .Z(n662) );
  XOR U579 ( .A(n663), .B(n664), .Z(n654) );
  AND U580 ( .A(n665), .B(n666), .Z(n664) );
  XOR U581 ( .A(n663), .B(n337), .Z(n666) );
  XNOR U582 ( .A(p_input[210]), .B(n667), .Z(n337) );
  AND U583 ( .A(n165), .B(n668), .Z(n667) );
  XOR U584 ( .A(p_input[242]), .B(p_input[210]), .Z(n668) );
  XNOR U585 ( .A(n334), .B(n663), .Z(n665) );
  XOR U586 ( .A(n669), .B(n670), .Z(n334) );
  AND U587 ( .A(n163), .B(n671), .Z(n670) );
  XOR U588 ( .A(p_input[178]), .B(p_input[146]), .Z(n671) );
  XOR U589 ( .A(n672), .B(n673), .Z(n663) );
  AND U590 ( .A(n674), .B(n675), .Z(n673) );
  XOR U591 ( .A(n672), .B(n349), .Z(n675) );
  XNOR U592 ( .A(p_input[209]), .B(n676), .Z(n349) );
  AND U593 ( .A(n165), .B(n677), .Z(n676) );
  XOR U594 ( .A(p_input[241]), .B(p_input[209]), .Z(n677) );
  XNOR U595 ( .A(n346), .B(n672), .Z(n674) );
  XOR U596 ( .A(n678), .B(n679), .Z(n346) );
  AND U597 ( .A(n163), .B(n680), .Z(n679) );
  XOR U598 ( .A(p_input[177]), .B(p_input[145]), .Z(n680) );
  XOR U599 ( .A(n681), .B(n682), .Z(n672) );
  AND U600 ( .A(n683), .B(n684), .Z(n682) );
  XOR U601 ( .A(n681), .B(n361), .Z(n684) );
  XNOR U602 ( .A(p_input[208]), .B(n685), .Z(n361) );
  AND U603 ( .A(n165), .B(n686), .Z(n685) );
  XOR U604 ( .A(p_input[240]), .B(p_input[208]), .Z(n686) );
  XNOR U605 ( .A(n358), .B(n681), .Z(n683) );
  XOR U606 ( .A(n687), .B(n688), .Z(n358) );
  AND U607 ( .A(n163), .B(n689), .Z(n688) );
  XOR U608 ( .A(p_input[176]), .B(p_input[144]), .Z(n689) );
  XOR U609 ( .A(n690), .B(n691), .Z(n681) );
  AND U610 ( .A(n692), .B(n693), .Z(n691) );
  XOR U611 ( .A(n690), .B(n373), .Z(n693) );
  XNOR U612 ( .A(p_input[207]), .B(n694), .Z(n373) );
  AND U613 ( .A(n165), .B(n695), .Z(n694) );
  XOR U614 ( .A(p_input[239]), .B(p_input[207]), .Z(n695) );
  XNOR U615 ( .A(n370), .B(n690), .Z(n692) );
  XOR U616 ( .A(n696), .B(n697), .Z(n370) );
  AND U617 ( .A(n163), .B(n698), .Z(n697) );
  XOR U618 ( .A(p_input[175]), .B(p_input[143]), .Z(n698) );
  XOR U619 ( .A(n699), .B(n700), .Z(n690) );
  AND U620 ( .A(n701), .B(n702), .Z(n700) );
  XOR U621 ( .A(n699), .B(n385), .Z(n702) );
  XNOR U622 ( .A(p_input[206]), .B(n703), .Z(n385) );
  AND U623 ( .A(n165), .B(n704), .Z(n703) );
  XOR U624 ( .A(p_input[238]), .B(p_input[206]), .Z(n704) );
  XNOR U625 ( .A(n382), .B(n699), .Z(n701) );
  XOR U626 ( .A(n705), .B(n706), .Z(n382) );
  AND U627 ( .A(n163), .B(n707), .Z(n706) );
  XOR U628 ( .A(p_input[174]), .B(p_input[142]), .Z(n707) );
  XOR U629 ( .A(n708), .B(n709), .Z(n699) );
  AND U630 ( .A(n710), .B(n711), .Z(n709) );
  XOR U631 ( .A(n708), .B(n397), .Z(n711) );
  XNOR U632 ( .A(p_input[205]), .B(n712), .Z(n397) );
  AND U633 ( .A(n165), .B(n713), .Z(n712) );
  XOR U634 ( .A(p_input[237]), .B(p_input[205]), .Z(n713) );
  XNOR U635 ( .A(n394), .B(n708), .Z(n710) );
  XOR U636 ( .A(n714), .B(n715), .Z(n394) );
  AND U637 ( .A(n163), .B(n716), .Z(n715) );
  XOR U638 ( .A(p_input[173]), .B(p_input[141]), .Z(n716) );
  XOR U639 ( .A(n717), .B(n718), .Z(n708) );
  AND U640 ( .A(n719), .B(n720), .Z(n718) );
  XOR U641 ( .A(n717), .B(n409), .Z(n720) );
  XNOR U642 ( .A(p_input[204]), .B(n721), .Z(n409) );
  AND U643 ( .A(n165), .B(n722), .Z(n721) );
  XOR U644 ( .A(p_input[236]), .B(p_input[204]), .Z(n722) );
  XNOR U645 ( .A(n406), .B(n717), .Z(n719) );
  XOR U646 ( .A(n723), .B(n724), .Z(n406) );
  AND U647 ( .A(n163), .B(n725), .Z(n724) );
  XOR U648 ( .A(p_input[172]), .B(p_input[140]), .Z(n725) );
  XOR U649 ( .A(n726), .B(n727), .Z(n717) );
  AND U650 ( .A(n728), .B(n729), .Z(n727) );
  XOR U651 ( .A(n726), .B(n421), .Z(n729) );
  XNOR U652 ( .A(p_input[203]), .B(n730), .Z(n421) );
  AND U653 ( .A(n165), .B(n731), .Z(n730) );
  XOR U654 ( .A(p_input[235]), .B(p_input[203]), .Z(n731) );
  XNOR U655 ( .A(n418), .B(n726), .Z(n728) );
  XOR U656 ( .A(n732), .B(n733), .Z(n418) );
  AND U657 ( .A(n163), .B(n734), .Z(n733) );
  XOR U658 ( .A(p_input[171]), .B(p_input[139]), .Z(n734) );
  XOR U659 ( .A(n735), .B(n736), .Z(n726) );
  AND U660 ( .A(n737), .B(n738), .Z(n736) );
  XOR U661 ( .A(n735), .B(n433), .Z(n738) );
  XNOR U662 ( .A(p_input[202]), .B(n739), .Z(n433) );
  AND U663 ( .A(n165), .B(n740), .Z(n739) );
  XOR U664 ( .A(p_input[234]), .B(p_input[202]), .Z(n740) );
  XNOR U665 ( .A(n430), .B(n735), .Z(n737) );
  XOR U666 ( .A(n741), .B(n742), .Z(n430) );
  AND U667 ( .A(n163), .B(n743), .Z(n742) );
  XOR U668 ( .A(p_input[170]), .B(p_input[138]), .Z(n743) );
  XOR U669 ( .A(n744), .B(n745), .Z(n735) );
  AND U670 ( .A(n746), .B(n747), .Z(n745) );
  XOR U671 ( .A(n744), .B(n445), .Z(n747) );
  XNOR U672 ( .A(p_input[201]), .B(n748), .Z(n445) );
  AND U673 ( .A(n165), .B(n749), .Z(n748) );
  XOR U674 ( .A(p_input[233]), .B(p_input[201]), .Z(n749) );
  XNOR U675 ( .A(n442), .B(n744), .Z(n746) );
  XOR U676 ( .A(n750), .B(n751), .Z(n442) );
  AND U677 ( .A(n163), .B(n752), .Z(n751) );
  XOR U678 ( .A(p_input[169]), .B(p_input[137]), .Z(n752) );
  XOR U679 ( .A(n753), .B(n754), .Z(n744) );
  AND U680 ( .A(n755), .B(n756), .Z(n754) );
  XOR U681 ( .A(n753), .B(n457), .Z(n756) );
  XNOR U682 ( .A(p_input[200]), .B(n757), .Z(n457) );
  AND U683 ( .A(n165), .B(n758), .Z(n757) );
  XOR U684 ( .A(p_input[232]), .B(p_input[200]), .Z(n758) );
  XNOR U685 ( .A(n454), .B(n753), .Z(n755) );
  XOR U686 ( .A(n759), .B(n760), .Z(n454) );
  AND U687 ( .A(n163), .B(n761), .Z(n760) );
  XOR U688 ( .A(p_input[168]), .B(p_input[136]), .Z(n761) );
  XOR U689 ( .A(n762), .B(n763), .Z(n753) );
  AND U690 ( .A(n764), .B(n765), .Z(n763) );
  XOR U691 ( .A(n762), .B(n469), .Z(n765) );
  XNOR U692 ( .A(p_input[199]), .B(n766), .Z(n469) );
  AND U693 ( .A(n165), .B(n767), .Z(n766) );
  XOR U694 ( .A(p_input[231]), .B(p_input[199]), .Z(n767) );
  XNOR U695 ( .A(n466), .B(n762), .Z(n764) );
  XOR U696 ( .A(n768), .B(n769), .Z(n466) );
  AND U697 ( .A(n163), .B(n770), .Z(n769) );
  XOR U698 ( .A(p_input[167]), .B(p_input[135]), .Z(n770) );
  XOR U699 ( .A(n771), .B(n772), .Z(n762) );
  AND U700 ( .A(n773), .B(n774), .Z(n772) );
  XOR U701 ( .A(n481), .B(n771), .Z(n774) );
  XNOR U702 ( .A(p_input[198]), .B(n775), .Z(n481) );
  AND U703 ( .A(n165), .B(n776), .Z(n775) );
  XOR U704 ( .A(p_input[230]), .B(p_input[198]), .Z(n776) );
  XNOR U705 ( .A(n771), .B(n478), .Z(n773) );
  XOR U706 ( .A(n777), .B(n778), .Z(n478) );
  AND U707 ( .A(n163), .B(n779), .Z(n778) );
  XOR U708 ( .A(p_input[166]), .B(p_input[134]), .Z(n779) );
  XOR U709 ( .A(n780), .B(n781), .Z(n771) );
  AND U710 ( .A(n782), .B(n783), .Z(n781) );
  XOR U711 ( .A(n780), .B(n493), .Z(n783) );
  XNOR U712 ( .A(p_input[197]), .B(n784), .Z(n493) );
  AND U713 ( .A(n165), .B(n785), .Z(n784) );
  XOR U714 ( .A(p_input[229]), .B(p_input[197]), .Z(n785) );
  XNOR U715 ( .A(n490), .B(n780), .Z(n782) );
  XOR U716 ( .A(n786), .B(n787), .Z(n490) );
  AND U717 ( .A(n163), .B(n788), .Z(n787) );
  XOR U718 ( .A(p_input[165]), .B(p_input[133]), .Z(n788) );
  XOR U719 ( .A(n789), .B(n790), .Z(n780) );
  AND U720 ( .A(n791), .B(n792), .Z(n790) );
  XOR U721 ( .A(n789), .B(n505), .Z(n792) );
  XNOR U722 ( .A(p_input[196]), .B(n793), .Z(n505) );
  AND U723 ( .A(n165), .B(n794), .Z(n793) );
  XOR U724 ( .A(p_input[228]), .B(p_input[196]), .Z(n794) );
  XNOR U725 ( .A(n502), .B(n789), .Z(n791) );
  XOR U726 ( .A(n795), .B(n796), .Z(n502) );
  AND U727 ( .A(n163), .B(n797), .Z(n796) );
  XOR U728 ( .A(p_input[164]), .B(p_input[132]), .Z(n797) );
  XOR U729 ( .A(n798), .B(n799), .Z(n789) );
  AND U730 ( .A(n800), .B(n801), .Z(n799) );
  XOR U731 ( .A(n798), .B(n517), .Z(n801) );
  XNOR U732 ( .A(p_input[195]), .B(n802), .Z(n517) );
  AND U733 ( .A(n165), .B(n803), .Z(n802) );
  XOR U734 ( .A(p_input[227]), .B(p_input[195]), .Z(n803) );
  XNOR U735 ( .A(n514), .B(n798), .Z(n800) );
  XOR U736 ( .A(n804), .B(n805), .Z(n514) );
  AND U737 ( .A(n163), .B(n806), .Z(n805) );
  XOR U738 ( .A(p_input[163]), .B(p_input[131]), .Z(n806) );
  XOR U739 ( .A(n807), .B(n808), .Z(n798) );
  AND U740 ( .A(n809), .B(n810), .Z(n808) );
  XOR U741 ( .A(n807), .B(n529), .Z(n810) );
  XNOR U742 ( .A(p_input[194]), .B(n811), .Z(n529) );
  AND U743 ( .A(n165), .B(n812), .Z(n811) );
  XOR U744 ( .A(p_input[226]), .B(p_input[194]), .Z(n812) );
  XNOR U745 ( .A(n526), .B(n807), .Z(n809) );
  XOR U746 ( .A(n813), .B(n814), .Z(n526) );
  AND U747 ( .A(n163), .B(n815), .Z(n814) );
  XOR U748 ( .A(p_input[162]), .B(p_input[130]), .Z(n815) );
  XOR U749 ( .A(n816), .B(n817), .Z(n807) );
  AND U750 ( .A(n818), .B(n819), .Z(n817) );
  XNOR U751 ( .A(n820), .B(n541), .Z(n819) );
  XNOR U752 ( .A(p_input[193]), .B(n821), .Z(n541) );
  AND U753 ( .A(n165), .B(n822), .Z(n821) );
  XNOR U754 ( .A(p_input[225]), .B(n823), .Z(n822) );
  IV U755 ( .A(p_input[193]), .Z(n823) );
  XNOR U756 ( .A(n538), .B(n816), .Z(n818) );
  XNOR U757 ( .A(p_input[129]), .B(n824), .Z(n538) );
  AND U758 ( .A(n163), .B(n825), .Z(n824) );
  XOR U759 ( .A(p_input[161]), .B(p_input[129]), .Z(n825) );
  IV U760 ( .A(n820), .Z(n816) );
  AND U761 ( .A(n546), .B(n549), .Z(n820) );
  XOR U762 ( .A(p_input[192]), .B(n826), .Z(n549) );
  AND U763 ( .A(n165), .B(n827), .Z(n826) );
  XOR U764 ( .A(p_input[224]), .B(p_input[192]), .Z(n827) );
  XOR U765 ( .A(n828), .B(n829), .Z(n165) );
  AND U766 ( .A(n830), .B(n831), .Z(n829) );
  XNOR U767 ( .A(p_input[255]), .B(n828), .Z(n831) );
  XOR U768 ( .A(n828), .B(p_input[223]), .Z(n830) );
  XOR U769 ( .A(n832), .B(n833), .Z(n828) );
  AND U770 ( .A(n834), .B(n835), .Z(n833) );
  XNOR U771 ( .A(p_input[254]), .B(n832), .Z(n835) );
  XOR U772 ( .A(n832), .B(p_input[222]), .Z(n834) );
  XOR U773 ( .A(n836), .B(n837), .Z(n832) );
  AND U774 ( .A(n838), .B(n839), .Z(n837) );
  XNOR U775 ( .A(p_input[253]), .B(n836), .Z(n839) );
  XOR U776 ( .A(n836), .B(p_input[221]), .Z(n838) );
  XOR U777 ( .A(n840), .B(n841), .Z(n836) );
  AND U778 ( .A(n842), .B(n843), .Z(n841) );
  XNOR U779 ( .A(p_input[252]), .B(n840), .Z(n843) );
  XOR U780 ( .A(n840), .B(p_input[220]), .Z(n842) );
  XOR U781 ( .A(n844), .B(n845), .Z(n840) );
  AND U782 ( .A(n846), .B(n847), .Z(n845) );
  XNOR U783 ( .A(p_input[251]), .B(n844), .Z(n847) );
  XOR U784 ( .A(n844), .B(p_input[219]), .Z(n846) );
  XOR U785 ( .A(n848), .B(n849), .Z(n844) );
  AND U786 ( .A(n850), .B(n851), .Z(n849) );
  XNOR U787 ( .A(p_input[250]), .B(n848), .Z(n851) );
  XOR U788 ( .A(n848), .B(p_input[218]), .Z(n850) );
  XOR U789 ( .A(n852), .B(n853), .Z(n848) );
  AND U790 ( .A(n854), .B(n855), .Z(n853) );
  XNOR U791 ( .A(p_input[249]), .B(n852), .Z(n855) );
  XOR U792 ( .A(n852), .B(p_input[217]), .Z(n854) );
  XOR U793 ( .A(n856), .B(n857), .Z(n852) );
  AND U794 ( .A(n858), .B(n859), .Z(n857) );
  XNOR U795 ( .A(p_input[248]), .B(n856), .Z(n859) );
  XOR U796 ( .A(n856), .B(p_input[216]), .Z(n858) );
  XOR U797 ( .A(n860), .B(n861), .Z(n856) );
  AND U798 ( .A(n862), .B(n863), .Z(n861) );
  XNOR U799 ( .A(p_input[247]), .B(n860), .Z(n863) );
  XOR U800 ( .A(n860), .B(p_input[215]), .Z(n862) );
  XOR U801 ( .A(n864), .B(n865), .Z(n860) );
  AND U802 ( .A(n866), .B(n867), .Z(n865) );
  XNOR U803 ( .A(p_input[246]), .B(n864), .Z(n867) );
  XOR U804 ( .A(n864), .B(p_input[214]), .Z(n866) );
  XOR U805 ( .A(n868), .B(n869), .Z(n864) );
  AND U806 ( .A(n870), .B(n871), .Z(n869) );
  XNOR U807 ( .A(p_input[245]), .B(n868), .Z(n871) );
  XOR U808 ( .A(n868), .B(p_input[213]), .Z(n870) );
  XOR U809 ( .A(n872), .B(n873), .Z(n868) );
  AND U810 ( .A(n874), .B(n875), .Z(n873) );
  XNOR U811 ( .A(p_input[244]), .B(n872), .Z(n875) );
  XOR U812 ( .A(n872), .B(p_input[212]), .Z(n874) );
  XOR U813 ( .A(n876), .B(n877), .Z(n872) );
  AND U814 ( .A(n878), .B(n879), .Z(n877) );
  XNOR U815 ( .A(p_input[243]), .B(n876), .Z(n879) );
  XOR U816 ( .A(n876), .B(p_input[211]), .Z(n878) );
  XOR U817 ( .A(n880), .B(n881), .Z(n876) );
  AND U818 ( .A(n882), .B(n883), .Z(n881) );
  XNOR U819 ( .A(p_input[242]), .B(n880), .Z(n883) );
  XOR U820 ( .A(n880), .B(p_input[210]), .Z(n882) );
  XOR U821 ( .A(n884), .B(n885), .Z(n880) );
  AND U822 ( .A(n886), .B(n887), .Z(n885) );
  XNOR U823 ( .A(p_input[241]), .B(n884), .Z(n887) );
  XOR U824 ( .A(n884), .B(p_input[209]), .Z(n886) );
  XOR U825 ( .A(n888), .B(n889), .Z(n884) );
  AND U826 ( .A(n890), .B(n891), .Z(n889) );
  XNOR U827 ( .A(p_input[240]), .B(n888), .Z(n891) );
  XOR U828 ( .A(n888), .B(p_input[208]), .Z(n890) );
  XOR U829 ( .A(n892), .B(n893), .Z(n888) );
  AND U830 ( .A(n894), .B(n895), .Z(n893) );
  XNOR U831 ( .A(p_input[239]), .B(n892), .Z(n895) );
  XOR U832 ( .A(n892), .B(p_input[207]), .Z(n894) );
  XOR U833 ( .A(n896), .B(n897), .Z(n892) );
  AND U834 ( .A(n898), .B(n899), .Z(n897) );
  XNOR U835 ( .A(p_input[238]), .B(n896), .Z(n899) );
  XOR U836 ( .A(n896), .B(p_input[206]), .Z(n898) );
  XOR U837 ( .A(n900), .B(n901), .Z(n896) );
  AND U838 ( .A(n902), .B(n903), .Z(n901) );
  XNOR U839 ( .A(p_input[237]), .B(n900), .Z(n903) );
  XOR U840 ( .A(n900), .B(p_input[205]), .Z(n902) );
  XOR U841 ( .A(n904), .B(n905), .Z(n900) );
  AND U842 ( .A(n906), .B(n907), .Z(n905) );
  XNOR U843 ( .A(p_input[236]), .B(n904), .Z(n907) );
  XOR U844 ( .A(n904), .B(p_input[204]), .Z(n906) );
  XOR U845 ( .A(n908), .B(n909), .Z(n904) );
  AND U846 ( .A(n910), .B(n911), .Z(n909) );
  XNOR U847 ( .A(p_input[235]), .B(n908), .Z(n911) );
  XOR U848 ( .A(n908), .B(p_input[203]), .Z(n910) );
  XOR U849 ( .A(n912), .B(n913), .Z(n908) );
  AND U850 ( .A(n914), .B(n915), .Z(n913) );
  XNOR U851 ( .A(p_input[234]), .B(n912), .Z(n915) );
  XOR U852 ( .A(n912), .B(p_input[202]), .Z(n914) );
  XOR U853 ( .A(n916), .B(n917), .Z(n912) );
  AND U854 ( .A(n918), .B(n919), .Z(n917) );
  XNOR U855 ( .A(p_input[233]), .B(n916), .Z(n919) );
  XOR U856 ( .A(n916), .B(p_input[201]), .Z(n918) );
  XOR U857 ( .A(n920), .B(n921), .Z(n916) );
  AND U858 ( .A(n922), .B(n923), .Z(n921) );
  XNOR U859 ( .A(p_input[232]), .B(n920), .Z(n923) );
  XOR U860 ( .A(n920), .B(p_input[200]), .Z(n922) );
  XOR U861 ( .A(n924), .B(n925), .Z(n920) );
  AND U862 ( .A(n926), .B(n927), .Z(n925) );
  XNOR U863 ( .A(p_input[231]), .B(n924), .Z(n927) );
  XOR U864 ( .A(n924), .B(p_input[199]), .Z(n926) );
  XOR U865 ( .A(n928), .B(n929), .Z(n924) );
  AND U866 ( .A(n930), .B(n931), .Z(n929) );
  XNOR U867 ( .A(p_input[230]), .B(n928), .Z(n931) );
  XOR U868 ( .A(n928), .B(p_input[198]), .Z(n930) );
  XOR U869 ( .A(n932), .B(n933), .Z(n928) );
  AND U870 ( .A(n934), .B(n935), .Z(n933) );
  XNOR U871 ( .A(p_input[229]), .B(n932), .Z(n935) );
  XOR U872 ( .A(n932), .B(p_input[197]), .Z(n934) );
  XOR U873 ( .A(n936), .B(n937), .Z(n932) );
  AND U874 ( .A(n938), .B(n939), .Z(n937) );
  XNOR U875 ( .A(p_input[228]), .B(n936), .Z(n939) );
  XOR U876 ( .A(n936), .B(p_input[196]), .Z(n938) );
  XOR U877 ( .A(n940), .B(n941), .Z(n936) );
  AND U878 ( .A(n942), .B(n943), .Z(n941) );
  XNOR U879 ( .A(p_input[227]), .B(n940), .Z(n943) );
  XOR U880 ( .A(n940), .B(p_input[195]), .Z(n942) );
  XOR U881 ( .A(n944), .B(n945), .Z(n940) );
  AND U882 ( .A(n946), .B(n947), .Z(n945) );
  XNOR U883 ( .A(p_input[226]), .B(n944), .Z(n947) );
  XOR U884 ( .A(n944), .B(p_input[194]), .Z(n946) );
  XNOR U885 ( .A(n948), .B(n949), .Z(n944) );
  AND U886 ( .A(n950), .B(n951), .Z(n949) );
  XOR U887 ( .A(p_input[225]), .B(n948), .Z(n951) );
  XNOR U888 ( .A(p_input[193]), .B(n948), .Z(n950) );
  AND U889 ( .A(p_input[224]), .B(n952), .Z(n948) );
  IV U890 ( .A(p_input[192]), .Z(n952) );
  XNOR U891 ( .A(p_input[128]), .B(n953), .Z(n546) );
  AND U892 ( .A(n163), .B(n954), .Z(n953) );
  XOR U893 ( .A(p_input[160]), .B(p_input[128]), .Z(n954) );
  XOR U894 ( .A(n955), .B(n956), .Z(n163) );
  AND U895 ( .A(n957), .B(n958), .Z(n956) );
  XNOR U896 ( .A(p_input[191]), .B(n955), .Z(n958) );
  XOR U897 ( .A(n955), .B(p_input[159]), .Z(n957) );
  XOR U898 ( .A(n959), .B(n960), .Z(n955) );
  AND U899 ( .A(n961), .B(n962), .Z(n960) );
  XNOR U900 ( .A(p_input[190]), .B(n959), .Z(n962) );
  XNOR U901 ( .A(n959), .B(n561), .Z(n961) );
  IV U902 ( .A(p_input[158]), .Z(n561) );
  XOR U903 ( .A(n963), .B(n964), .Z(n959) );
  AND U904 ( .A(n965), .B(n966), .Z(n964) );
  XNOR U905 ( .A(p_input[189]), .B(n963), .Z(n966) );
  XNOR U906 ( .A(n963), .B(n570), .Z(n965) );
  IV U907 ( .A(p_input[157]), .Z(n570) );
  XOR U908 ( .A(n967), .B(n968), .Z(n963) );
  AND U909 ( .A(n969), .B(n970), .Z(n968) );
  XNOR U910 ( .A(p_input[188]), .B(n967), .Z(n970) );
  XNOR U911 ( .A(n967), .B(n579), .Z(n969) );
  IV U912 ( .A(p_input[156]), .Z(n579) );
  XOR U913 ( .A(n971), .B(n972), .Z(n967) );
  AND U914 ( .A(n973), .B(n974), .Z(n972) );
  XNOR U915 ( .A(p_input[187]), .B(n971), .Z(n974) );
  XNOR U916 ( .A(n971), .B(n588), .Z(n973) );
  IV U917 ( .A(p_input[155]), .Z(n588) );
  XOR U918 ( .A(n975), .B(n976), .Z(n971) );
  AND U919 ( .A(n977), .B(n978), .Z(n976) );
  XNOR U920 ( .A(p_input[186]), .B(n975), .Z(n978) );
  XNOR U921 ( .A(n975), .B(n597), .Z(n977) );
  IV U922 ( .A(p_input[154]), .Z(n597) );
  XOR U923 ( .A(n979), .B(n980), .Z(n975) );
  AND U924 ( .A(n981), .B(n982), .Z(n980) );
  XNOR U925 ( .A(p_input[185]), .B(n979), .Z(n982) );
  XNOR U926 ( .A(n979), .B(n606), .Z(n981) );
  IV U927 ( .A(p_input[153]), .Z(n606) );
  XOR U928 ( .A(n983), .B(n984), .Z(n979) );
  AND U929 ( .A(n985), .B(n986), .Z(n984) );
  XNOR U930 ( .A(p_input[184]), .B(n983), .Z(n986) );
  XNOR U931 ( .A(n983), .B(n615), .Z(n985) );
  IV U932 ( .A(p_input[152]), .Z(n615) );
  XOR U933 ( .A(n987), .B(n988), .Z(n983) );
  AND U934 ( .A(n989), .B(n990), .Z(n988) );
  XNOR U935 ( .A(p_input[183]), .B(n987), .Z(n990) );
  XNOR U936 ( .A(n987), .B(n624), .Z(n989) );
  IV U937 ( .A(p_input[151]), .Z(n624) );
  XOR U938 ( .A(n991), .B(n992), .Z(n987) );
  AND U939 ( .A(n993), .B(n994), .Z(n992) );
  XNOR U940 ( .A(p_input[182]), .B(n991), .Z(n994) );
  XNOR U941 ( .A(n991), .B(n633), .Z(n993) );
  IV U942 ( .A(p_input[150]), .Z(n633) );
  XOR U943 ( .A(n995), .B(n996), .Z(n991) );
  AND U944 ( .A(n997), .B(n998), .Z(n996) );
  XNOR U945 ( .A(p_input[181]), .B(n995), .Z(n998) );
  XNOR U946 ( .A(n995), .B(n642), .Z(n997) );
  IV U947 ( .A(p_input[149]), .Z(n642) );
  XOR U948 ( .A(n999), .B(n1000), .Z(n995) );
  AND U949 ( .A(n1001), .B(n1002), .Z(n1000) );
  XNOR U950 ( .A(p_input[180]), .B(n999), .Z(n1002) );
  XNOR U951 ( .A(n999), .B(n651), .Z(n1001) );
  IV U952 ( .A(p_input[148]), .Z(n651) );
  XOR U953 ( .A(n1003), .B(n1004), .Z(n999) );
  AND U954 ( .A(n1005), .B(n1006), .Z(n1004) );
  XNOR U955 ( .A(p_input[179]), .B(n1003), .Z(n1006) );
  XNOR U956 ( .A(n1003), .B(n660), .Z(n1005) );
  IV U957 ( .A(p_input[147]), .Z(n660) );
  XOR U958 ( .A(n1007), .B(n1008), .Z(n1003) );
  AND U959 ( .A(n1009), .B(n1010), .Z(n1008) );
  XNOR U960 ( .A(p_input[178]), .B(n1007), .Z(n1010) );
  XNOR U961 ( .A(n1007), .B(n669), .Z(n1009) );
  IV U962 ( .A(p_input[146]), .Z(n669) );
  XOR U963 ( .A(n1011), .B(n1012), .Z(n1007) );
  AND U964 ( .A(n1013), .B(n1014), .Z(n1012) );
  XNOR U965 ( .A(p_input[177]), .B(n1011), .Z(n1014) );
  XNOR U966 ( .A(n1011), .B(n678), .Z(n1013) );
  IV U967 ( .A(p_input[145]), .Z(n678) );
  XOR U968 ( .A(n1015), .B(n1016), .Z(n1011) );
  AND U969 ( .A(n1017), .B(n1018), .Z(n1016) );
  XNOR U970 ( .A(p_input[176]), .B(n1015), .Z(n1018) );
  XNOR U971 ( .A(n1015), .B(n687), .Z(n1017) );
  IV U972 ( .A(p_input[144]), .Z(n687) );
  XOR U973 ( .A(n1019), .B(n1020), .Z(n1015) );
  AND U974 ( .A(n1021), .B(n1022), .Z(n1020) );
  XNOR U975 ( .A(p_input[175]), .B(n1019), .Z(n1022) );
  XNOR U976 ( .A(n1019), .B(n696), .Z(n1021) );
  IV U977 ( .A(p_input[143]), .Z(n696) );
  XOR U978 ( .A(n1023), .B(n1024), .Z(n1019) );
  AND U979 ( .A(n1025), .B(n1026), .Z(n1024) );
  XNOR U980 ( .A(p_input[174]), .B(n1023), .Z(n1026) );
  XNOR U981 ( .A(n1023), .B(n705), .Z(n1025) );
  IV U982 ( .A(p_input[142]), .Z(n705) );
  XOR U983 ( .A(n1027), .B(n1028), .Z(n1023) );
  AND U984 ( .A(n1029), .B(n1030), .Z(n1028) );
  XNOR U985 ( .A(p_input[173]), .B(n1027), .Z(n1030) );
  XNOR U986 ( .A(n1027), .B(n714), .Z(n1029) );
  IV U987 ( .A(p_input[141]), .Z(n714) );
  XOR U988 ( .A(n1031), .B(n1032), .Z(n1027) );
  AND U989 ( .A(n1033), .B(n1034), .Z(n1032) );
  XNOR U990 ( .A(p_input[172]), .B(n1031), .Z(n1034) );
  XNOR U991 ( .A(n1031), .B(n723), .Z(n1033) );
  IV U992 ( .A(p_input[140]), .Z(n723) );
  XOR U993 ( .A(n1035), .B(n1036), .Z(n1031) );
  AND U994 ( .A(n1037), .B(n1038), .Z(n1036) );
  XNOR U995 ( .A(p_input[171]), .B(n1035), .Z(n1038) );
  XNOR U996 ( .A(n1035), .B(n732), .Z(n1037) );
  IV U997 ( .A(p_input[139]), .Z(n732) );
  XOR U998 ( .A(n1039), .B(n1040), .Z(n1035) );
  AND U999 ( .A(n1041), .B(n1042), .Z(n1040) );
  XNOR U1000 ( .A(p_input[170]), .B(n1039), .Z(n1042) );
  XNOR U1001 ( .A(n1039), .B(n741), .Z(n1041) );
  IV U1002 ( .A(p_input[138]), .Z(n741) );
  XOR U1003 ( .A(n1043), .B(n1044), .Z(n1039) );
  AND U1004 ( .A(n1045), .B(n1046), .Z(n1044) );
  XNOR U1005 ( .A(p_input[169]), .B(n1043), .Z(n1046) );
  XNOR U1006 ( .A(n1043), .B(n750), .Z(n1045) );
  IV U1007 ( .A(p_input[137]), .Z(n750) );
  XOR U1008 ( .A(n1047), .B(n1048), .Z(n1043) );
  AND U1009 ( .A(n1049), .B(n1050), .Z(n1048) );
  XNOR U1010 ( .A(p_input[168]), .B(n1047), .Z(n1050) );
  XNOR U1011 ( .A(n1047), .B(n759), .Z(n1049) );
  IV U1012 ( .A(p_input[136]), .Z(n759) );
  XOR U1013 ( .A(n1051), .B(n1052), .Z(n1047) );
  AND U1014 ( .A(n1053), .B(n1054), .Z(n1052) );
  XNOR U1015 ( .A(p_input[167]), .B(n1051), .Z(n1054) );
  XNOR U1016 ( .A(n1051), .B(n768), .Z(n1053) );
  IV U1017 ( .A(p_input[135]), .Z(n768) );
  XOR U1018 ( .A(n1055), .B(n1056), .Z(n1051) );
  AND U1019 ( .A(n1057), .B(n1058), .Z(n1056) );
  XNOR U1020 ( .A(p_input[166]), .B(n1055), .Z(n1058) );
  XNOR U1021 ( .A(n1055), .B(n777), .Z(n1057) );
  IV U1022 ( .A(p_input[134]), .Z(n777) );
  XOR U1023 ( .A(n1059), .B(n1060), .Z(n1055) );
  AND U1024 ( .A(n1061), .B(n1062), .Z(n1060) );
  XNOR U1025 ( .A(p_input[165]), .B(n1059), .Z(n1062) );
  XNOR U1026 ( .A(n1059), .B(n786), .Z(n1061) );
  IV U1027 ( .A(p_input[133]), .Z(n786) );
  XOR U1028 ( .A(n1063), .B(n1064), .Z(n1059) );
  AND U1029 ( .A(n1065), .B(n1066), .Z(n1064) );
  XNOR U1030 ( .A(p_input[164]), .B(n1063), .Z(n1066) );
  XNOR U1031 ( .A(n1063), .B(n795), .Z(n1065) );
  IV U1032 ( .A(p_input[132]), .Z(n795) );
  XOR U1033 ( .A(n1067), .B(n1068), .Z(n1063) );
  AND U1034 ( .A(n1069), .B(n1070), .Z(n1068) );
  XNOR U1035 ( .A(p_input[163]), .B(n1067), .Z(n1070) );
  XNOR U1036 ( .A(n1067), .B(n804), .Z(n1069) );
  IV U1037 ( .A(p_input[131]), .Z(n804) );
  XOR U1038 ( .A(n1071), .B(n1072), .Z(n1067) );
  AND U1039 ( .A(n1073), .B(n1074), .Z(n1072) );
  XNOR U1040 ( .A(p_input[162]), .B(n1071), .Z(n1074) );
  XNOR U1041 ( .A(n1071), .B(n813), .Z(n1073) );
  IV U1042 ( .A(p_input[130]), .Z(n813) );
  XNOR U1043 ( .A(n1075), .B(n1076), .Z(n1071) );
  AND U1044 ( .A(n1077), .B(n1078), .Z(n1076) );
  XOR U1045 ( .A(p_input[161]), .B(n1075), .Z(n1078) );
  XNOR U1046 ( .A(p_input[129]), .B(n1075), .Z(n1077) );
  AND U1047 ( .A(p_input[160]), .B(n1079), .Z(n1075) );
  IV U1048 ( .A(p_input[128]), .Z(n1079) );
  XOR U1049 ( .A(n1080), .B(n1081), .Z(n31) );
  AND U1050 ( .A(n166), .B(n1082), .Z(n1081) );
  XNOR U1051 ( .A(n1083), .B(n1080), .Z(n1082) );
  XOR U1052 ( .A(n1084), .B(n1085), .Z(n166) );
  AND U1053 ( .A(n1086), .B(n1087), .Z(n1085) );
  XNOR U1054 ( .A(n185), .B(n1084), .Z(n1087) );
  AND U1055 ( .A(p_input[95]), .B(p_input[127]), .Z(n185) );
  XNOR U1056 ( .A(n1084), .B(n182), .Z(n1086) );
  IV U1057 ( .A(n1088), .Z(n182) );
  AND U1058 ( .A(p_input[31]), .B(p_input[63]), .Z(n1088) );
  XOR U1059 ( .A(n1089), .B(n1090), .Z(n1084) );
  AND U1060 ( .A(n1091), .B(n1092), .Z(n1090) );
  XOR U1061 ( .A(n1089), .B(n197), .Z(n1092) );
  XNOR U1062 ( .A(p_input[94]), .B(n1093), .Z(n197) );
  AND U1063 ( .A(n173), .B(n1094), .Z(n1093) );
  XOR U1064 ( .A(p_input[94]), .B(p_input[126]), .Z(n1094) );
  XNOR U1065 ( .A(n194), .B(n1089), .Z(n1091) );
  XOR U1066 ( .A(n1095), .B(n1096), .Z(n194) );
  AND U1067 ( .A(n170), .B(n1097), .Z(n1096) );
  XOR U1068 ( .A(p_input[62]), .B(p_input[30]), .Z(n1097) );
  XOR U1069 ( .A(n1098), .B(n1099), .Z(n1089) );
  AND U1070 ( .A(n1100), .B(n1101), .Z(n1099) );
  XOR U1071 ( .A(n1098), .B(n209), .Z(n1101) );
  XNOR U1072 ( .A(p_input[93]), .B(n1102), .Z(n209) );
  AND U1073 ( .A(n173), .B(n1103), .Z(n1102) );
  XOR U1074 ( .A(p_input[93]), .B(p_input[125]), .Z(n1103) );
  XNOR U1075 ( .A(n206), .B(n1098), .Z(n1100) );
  XOR U1076 ( .A(n1104), .B(n1105), .Z(n206) );
  AND U1077 ( .A(n170), .B(n1106), .Z(n1105) );
  XOR U1078 ( .A(p_input[61]), .B(p_input[29]), .Z(n1106) );
  XOR U1079 ( .A(n1107), .B(n1108), .Z(n1098) );
  AND U1080 ( .A(n1109), .B(n1110), .Z(n1108) );
  XOR U1081 ( .A(n1107), .B(n221), .Z(n1110) );
  XNOR U1082 ( .A(p_input[92]), .B(n1111), .Z(n221) );
  AND U1083 ( .A(n173), .B(n1112), .Z(n1111) );
  XOR U1084 ( .A(p_input[92]), .B(p_input[124]), .Z(n1112) );
  XNOR U1085 ( .A(n218), .B(n1107), .Z(n1109) );
  XOR U1086 ( .A(n1113), .B(n1114), .Z(n218) );
  AND U1087 ( .A(n170), .B(n1115), .Z(n1114) );
  XOR U1088 ( .A(p_input[60]), .B(p_input[28]), .Z(n1115) );
  XOR U1089 ( .A(n1116), .B(n1117), .Z(n1107) );
  AND U1090 ( .A(n1118), .B(n1119), .Z(n1117) );
  XOR U1091 ( .A(n1116), .B(n233), .Z(n1119) );
  XNOR U1092 ( .A(p_input[91]), .B(n1120), .Z(n233) );
  AND U1093 ( .A(n173), .B(n1121), .Z(n1120) );
  XOR U1094 ( .A(p_input[91]), .B(p_input[123]), .Z(n1121) );
  XNOR U1095 ( .A(n230), .B(n1116), .Z(n1118) );
  XOR U1096 ( .A(n1122), .B(n1123), .Z(n230) );
  AND U1097 ( .A(n170), .B(n1124), .Z(n1123) );
  XOR U1098 ( .A(p_input[59]), .B(p_input[27]), .Z(n1124) );
  XOR U1099 ( .A(n1125), .B(n1126), .Z(n1116) );
  AND U1100 ( .A(n1127), .B(n1128), .Z(n1126) );
  XOR U1101 ( .A(n1125), .B(n245), .Z(n1128) );
  XNOR U1102 ( .A(p_input[90]), .B(n1129), .Z(n245) );
  AND U1103 ( .A(n173), .B(n1130), .Z(n1129) );
  XOR U1104 ( .A(p_input[90]), .B(p_input[122]), .Z(n1130) );
  XNOR U1105 ( .A(n242), .B(n1125), .Z(n1127) );
  XOR U1106 ( .A(n1131), .B(n1132), .Z(n242) );
  AND U1107 ( .A(n170), .B(n1133), .Z(n1132) );
  XOR U1108 ( .A(p_input[58]), .B(p_input[26]), .Z(n1133) );
  XOR U1109 ( .A(n1134), .B(n1135), .Z(n1125) );
  AND U1110 ( .A(n1136), .B(n1137), .Z(n1135) );
  XOR U1111 ( .A(n1134), .B(n257), .Z(n1137) );
  XNOR U1112 ( .A(p_input[89]), .B(n1138), .Z(n257) );
  AND U1113 ( .A(n173), .B(n1139), .Z(n1138) );
  XOR U1114 ( .A(p_input[89]), .B(p_input[121]), .Z(n1139) );
  XNOR U1115 ( .A(n254), .B(n1134), .Z(n1136) );
  XOR U1116 ( .A(n1140), .B(n1141), .Z(n254) );
  AND U1117 ( .A(n170), .B(n1142), .Z(n1141) );
  XOR U1118 ( .A(p_input[57]), .B(p_input[25]), .Z(n1142) );
  XOR U1119 ( .A(n1143), .B(n1144), .Z(n1134) );
  AND U1120 ( .A(n1145), .B(n1146), .Z(n1144) );
  XOR U1121 ( .A(n1143), .B(n269), .Z(n1146) );
  XNOR U1122 ( .A(p_input[88]), .B(n1147), .Z(n269) );
  AND U1123 ( .A(n173), .B(n1148), .Z(n1147) );
  XOR U1124 ( .A(p_input[88]), .B(p_input[120]), .Z(n1148) );
  XNOR U1125 ( .A(n266), .B(n1143), .Z(n1145) );
  XOR U1126 ( .A(n1149), .B(n1150), .Z(n266) );
  AND U1127 ( .A(n170), .B(n1151), .Z(n1150) );
  XOR U1128 ( .A(p_input[56]), .B(p_input[24]), .Z(n1151) );
  XOR U1129 ( .A(n1152), .B(n1153), .Z(n1143) );
  AND U1130 ( .A(n1154), .B(n1155), .Z(n1153) );
  XOR U1131 ( .A(n1152), .B(n281), .Z(n1155) );
  XNOR U1132 ( .A(p_input[87]), .B(n1156), .Z(n281) );
  AND U1133 ( .A(n173), .B(n1157), .Z(n1156) );
  XOR U1134 ( .A(p_input[87]), .B(p_input[119]), .Z(n1157) );
  XNOR U1135 ( .A(n278), .B(n1152), .Z(n1154) );
  XOR U1136 ( .A(n1158), .B(n1159), .Z(n278) );
  AND U1137 ( .A(n170), .B(n1160), .Z(n1159) );
  XOR U1138 ( .A(p_input[55]), .B(p_input[23]), .Z(n1160) );
  XOR U1139 ( .A(n1161), .B(n1162), .Z(n1152) );
  AND U1140 ( .A(n1163), .B(n1164), .Z(n1162) );
  XOR U1141 ( .A(n1161), .B(n293), .Z(n1164) );
  XNOR U1142 ( .A(p_input[86]), .B(n1165), .Z(n293) );
  AND U1143 ( .A(n173), .B(n1166), .Z(n1165) );
  XOR U1144 ( .A(p_input[86]), .B(p_input[118]), .Z(n1166) );
  XNOR U1145 ( .A(n290), .B(n1161), .Z(n1163) );
  XOR U1146 ( .A(n1167), .B(n1168), .Z(n290) );
  AND U1147 ( .A(n170), .B(n1169), .Z(n1168) );
  XOR U1148 ( .A(p_input[54]), .B(p_input[22]), .Z(n1169) );
  XOR U1149 ( .A(n1170), .B(n1171), .Z(n1161) );
  AND U1150 ( .A(n1172), .B(n1173), .Z(n1171) );
  XOR U1151 ( .A(n1170), .B(n305), .Z(n1173) );
  XNOR U1152 ( .A(p_input[85]), .B(n1174), .Z(n305) );
  AND U1153 ( .A(n173), .B(n1175), .Z(n1174) );
  XOR U1154 ( .A(p_input[85]), .B(p_input[117]), .Z(n1175) );
  XNOR U1155 ( .A(n302), .B(n1170), .Z(n1172) );
  XOR U1156 ( .A(n1176), .B(n1177), .Z(n302) );
  AND U1157 ( .A(n170), .B(n1178), .Z(n1177) );
  XOR U1158 ( .A(p_input[53]), .B(p_input[21]), .Z(n1178) );
  XOR U1159 ( .A(n1179), .B(n1180), .Z(n1170) );
  AND U1160 ( .A(n1181), .B(n1182), .Z(n1180) );
  XOR U1161 ( .A(n1179), .B(n317), .Z(n1182) );
  XNOR U1162 ( .A(p_input[84]), .B(n1183), .Z(n317) );
  AND U1163 ( .A(n173), .B(n1184), .Z(n1183) );
  XOR U1164 ( .A(p_input[84]), .B(p_input[116]), .Z(n1184) );
  XNOR U1165 ( .A(n314), .B(n1179), .Z(n1181) );
  XOR U1166 ( .A(n1185), .B(n1186), .Z(n314) );
  AND U1167 ( .A(n170), .B(n1187), .Z(n1186) );
  XOR U1168 ( .A(p_input[52]), .B(p_input[20]), .Z(n1187) );
  XOR U1169 ( .A(n1188), .B(n1189), .Z(n1179) );
  AND U1170 ( .A(n1190), .B(n1191), .Z(n1189) );
  XOR U1171 ( .A(n1188), .B(n329), .Z(n1191) );
  XNOR U1172 ( .A(p_input[83]), .B(n1192), .Z(n329) );
  AND U1173 ( .A(n173), .B(n1193), .Z(n1192) );
  XOR U1174 ( .A(p_input[83]), .B(p_input[115]), .Z(n1193) );
  XNOR U1175 ( .A(n326), .B(n1188), .Z(n1190) );
  XOR U1176 ( .A(n1194), .B(n1195), .Z(n326) );
  AND U1177 ( .A(n170), .B(n1196), .Z(n1195) );
  XOR U1178 ( .A(p_input[51]), .B(p_input[19]), .Z(n1196) );
  XOR U1179 ( .A(n1197), .B(n1198), .Z(n1188) );
  AND U1180 ( .A(n1199), .B(n1200), .Z(n1198) );
  XOR U1181 ( .A(n1197), .B(n341), .Z(n1200) );
  XNOR U1182 ( .A(p_input[82]), .B(n1201), .Z(n341) );
  AND U1183 ( .A(n173), .B(n1202), .Z(n1201) );
  XOR U1184 ( .A(p_input[82]), .B(p_input[114]), .Z(n1202) );
  XNOR U1185 ( .A(n338), .B(n1197), .Z(n1199) );
  XOR U1186 ( .A(n1203), .B(n1204), .Z(n338) );
  AND U1187 ( .A(n170), .B(n1205), .Z(n1204) );
  XOR U1188 ( .A(p_input[50]), .B(p_input[18]), .Z(n1205) );
  XOR U1189 ( .A(n1206), .B(n1207), .Z(n1197) );
  AND U1190 ( .A(n1208), .B(n1209), .Z(n1207) );
  XOR U1191 ( .A(n1206), .B(n353), .Z(n1209) );
  XNOR U1192 ( .A(p_input[81]), .B(n1210), .Z(n353) );
  AND U1193 ( .A(n173), .B(n1211), .Z(n1210) );
  XOR U1194 ( .A(p_input[81]), .B(p_input[113]), .Z(n1211) );
  XNOR U1195 ( .A(n350), .B(n1206), .Z(n1208) );
  XOR U1196 ( .A(n1212), .B(n1213), .Z(n350) );
  AND U1197 ( .A(n170), .B(n1214), .Z(n1213) );
  XOR U1198 ( .A(p_input[49]), .B(p_input[17]), .Z(n1214) );
  XOR U1199 ( .A(n1215), .B(n1216), .Z(n1206) );
  AND U1200 ( .A(n1217), .B(n1218), .Z(n1216) );
  XOR U1201 ( .A(n1215), .B(n365), .Z(n1218) );
  XNOR U1202 ( .A(p_input[80]), .B(n1219), .Z(n365) );
  AND U1203 ( .A(n173), .B(n1220), .Z(n1219) );
  XOR U1204 ( .A(p_input[80]), .B(p_input[112]), .Z(n1220) );
  XNOR U1205 ( .A(n362), .B(n1215), .Z(n1217) );
  XOR U1206 ( .A(n1221), .B(n1222), .Z(n362) );
  AND U1207 ( .A(n170), .B(n1223), .Z(n1222) );
  XOR U1208 ( .A(p_input[48]), .B(p_input[16]), .Z(n1223) );
  XOR U1209 ( .A(n1224), .B(n1225), .Z(n1215) );
  AND U1210 ( .A(n1226), .B(n1227), .Z(n1225) );
  XOR U1211 ( .A(n1224), .B(n377), .Z(n1227) );
  XNOR U1212 ( .A(p_input[79]), .B(n1228), .Z(n377) );
  AND U1213 ( .A(n173), .B(n1229), .Z(n1228) );
  XOR U1214 ( .A(p_input[79]), .B(p_input[111]), .Z(n1229) );
  XNOR U1215 ( .A(n374), .B(n1224), .Z(n1226) );
  XOR U1216 ( .A(n1230), .B(n1231), .Z(n374) );
  AND U1217 ( .A(n170), .B(n1232), .Z(n1231) );
  XOR U1218 ( .A(p_input[47]), .B(p_input[15]), .Z(n1232) );
  XOR U1219 ( .A(n1233), .B(n1234), .Z(n1224) );
  AND U1220 ( .A(n1235), .B(n1236), .Z(n1234) );
  XOR U1221 ( .A(n1233), .B(n389), .Z(n1236) );
  XNOR U1222 ( .A(p_input[78]), .B(n1237), .Z(n389) );
  AND U1223 ( .A(n173), .B(n1238), .Z(n1237) );
  XOR U1224 ( .A(p_input[78]), .B(p_input[110]), .Z(n1238) );
  XNOR U1225 ( .A(n386), .B(n1233), .Z(n1235) );
  XOR U1226 ( .A(n1239), .B(n1240), .Z(n386) );
  AND U1227 ( .A(n170), .B(n1241), .Z(n1240) );
  XOR U1228 ( .A(p_input[46]), .B(p_input[14]), .Z(n1241) );
  XOR U1229 ( .A(n1242), .B(n1243), .Z(n1233) );
  AND U1230 ( .A(n1244), .B(n1245), .Z(n1243) );
  XOR U1231 ( .A(n1242), .B(n401), .Z(n1245) );
  XNOR U1232 ( .A(p_input[77]), .B(n1246), .Z(n401) );
  AND U1233 ( .A(n173), .B(n1247), .Z(n1246) );
  XOR U1234 ( .A(p_input[77]), .B(p_input[109]), .Z(n1247) );
  XNOR U1235 ( .A(n398), .B(n1242), .Z(n1244) );
  XOR U1236 ( .A(n1248), .B(n1249), .Z(n398) );
  AND U1237 ( .A(n170), .B(n1250), .Z(n1249) );
  XOR U1238 ( .A(p_input[45]), .B(p_input[13]), .Z(n1250) );
  XOR U1239 ( .A(n1251), .B(n1252), .Z(n1242) );
  AND U1240 ( .A(n1253), .B(n1254), .Z(n1252) );
  XOR U1241 ( .A(n1251), .B(n413), .Z(n1254) );
  XNOR U1242 ( .A(p_input[76]), .B(n1255), .Z(n413) );
  AND U1243 ( .A(n173), .B(n1256), .Z(n1255) );
  XOR U1244 ( .A(p_input[76]), .B(p_input[108]), .Z(n1256) );
  XNOR U1245 ( .A(n410), .B(n1251), .Z(n1253) );
  XOR U1246 ( .A(n1257), .B(n1258), .Z(n410) );
  AND U1247 ( .A(n170), .B(n1259), .Z(n1258) );
  XOR U1248 ( .A(p_input[44]), .B(p_input[12]), .Z(n1259) );
  XOR U1249 ( .A(n1260), .B(n1261), .Z(n1251) );
  AND U1250 ( .A(n1262), .B(n1263), .Z(n1261) );
  XOR U1251 ( .A(n1260), .B(n425), .Z(n1263) );
  XNOR U1252 ( .A(p_input[75]), .B(n1264), .Z(n425) );
  AND U1253 ( .A(n173), .B(n1265), .Z(n1264) );
  XOR U1254 ( .A(p_input[75]), .B(p_input[107]), .Z(n1265) );
  XNOR U1255 ( .A(n422), .B(n1260), .Z(n1262) );
  XOR U1256 ( .A(n1266), .B(n1267), .Z(n422) );
  AND U1257 ( .A(n170), .B(n1268), .Z(n1267) );
  XOR U1258 ( .A(p_input[43]), .B(p_input[11]), .Z(n1268) );
  XOR U1259 ( .A(n1269), .B(n1270), .Z(n1260) );
  AND U1260 ( .A(n1271), .B(n1272), .Z(n1270) );
  XOR U1261 ( .A(n1269), .B(n437), .Z(n1272) );
  XNOR U1262 ( .A(p_input[74]), .B(n1273), .Z(n437) );
  AND U1263 ( .A(n173), .B(n1274), .Z(n1273) );
  XOR U1264 ( .A(p_input[74]), .B(p_input[106]), .Z(n1274) );
  XNOR U1265 ( .A(n434), .B(n1269), .Z(n1271) );
  XOR U1266 ( .A(n1275), .B(n1276), .Z(n434) );
  AND U1267 ( .A(n170), .B(n1277), .Z(n1276) );
  XOR U1268 ( .A(p_input[42]), .B(p_input[10]), .Z(n1277) );
  XOR U1269 ( .A(n1278), .B(n1279), .Z(n1269) );
  AND U1270 ( .A(n1280), .B(n1281), .Z(n1279) );
  XOR U1271 ( .A(n1278), .B(n449), .Z(n1281) );
  XNOR U1272 ( .A(p_input[73]), .B(n1282), .Z(n449) );
  AND U1273 ( .A(n173), .B(n1283), .Z(n1282) );
  XOR U1274 ( .A(p_input[73]), .B(p_input[105]), .Z(n1283) );
  XNOR U1275 ( .A(n446), .B(n1278), .Z(n1280) );
  XOR U1276 ( .A(n1284), .B(n1285), .Z(n446) );
  AND U1277 ( .A(n170), .B(n1286), .Z(n1285) );
  XOR U1278 ( .A(p_input[9]), .B(p_input[41]), .Z(n1286) );
  XOR U1279 ( .A(n1287), .B(n1288), .Z(n1278) );
  AND U1280 ( .A(n1289), .B(n1290), .Z(n1288) );
  XOR U1281 ( .A(n1287), .B(n461), .Z(n1290) );
  XNOR U1282 ( .A(p_input[72]), .B(n1291), .Z(n461) );
  AND U1283 ( .A(n173), .B(n1292), .Z(n1291) );
  XOR U1284 ( .A(p_input[72]), .B(p_input[104]), .Z(n1292) );
  XNOR U1285 ( .A(n458), .B(n1287), .Z(n1289) );
  XOR U1286 ( .A(n1293), .B(n1294), .Z(n458) );
  AND U1287 ( .A(n170), .B(n1295), .Z(n1294) );
  XOR U1288 ( .A(p_input[8]), .B(p_input[40]), .Z(n1295) );
  XOR U1289 ( .A(n1296), .B(n1297), .Z(n1287) );
  AND U1290 ( .A(n1298), .B(n1299), .Z(n1297) );
  XOR U1291 ( .A(n1296), .B(n473), .Z(n1299) );
  XNOR U1292 ( .A(p_input[71]), .B(n1300), .Z(n473) );
  AND U1293 ( .A(n173), .B(n1301), .Z(n1300) );
  XOR U1294 ( .A(p_input[71]), .B(p_input[103]), .Z(n1301) );
  XNOR U1295 ( .A(n470), .B(n1296), .Z(n1298) );
  XOR U1296 ( .A(n1302), .B(n1303), .Z(n470) );
  AND U1297 ( .A(n170), .B(n1304), .Z(n1303) );
  XOR U1298 ( .A(p_input[7]), .B(p_input[39]), .Z(n1304) );
  XOR U1299 ( .A(n1305), .B(n1306), .Z(n1296) );
  AND U1300 ( .A(n1307), .B(n1308), .Z(n1306) );
  XOR U1301 ( .A(n485), .B(n1305), .Z(n1308) );
  XNOR U1302 ( .A(p_input[70]), .B(n1309), .Z(n485) );
  AND U1303 ( .A(n173), .B(n1310), .Z(n1309) );
  XOR U1304 ( .A(p_input[70]), .B(p_input[102]), .Z(n1310) );
  XNOR U1305 ( .A(n1305), .B(n482), .Z(n1307) );
  XOR U1306 ( .A(n1311), .B(n1312), .Z(n482) );
  AND U1307 ( .A(n170), .B(n1313), .Z(n1312) );
  XOR U1308 ( .A(p_input[6]), .B(p_input[38]), .Z(n1313) );
  XOR U1309 ( .A(n1314), .B(n1315), .Z(n1305) );
  AND U1310 ( .A(n1316), .B(n1317), .Z(n1315) );
  XOR U1311 ( .A(n1314), .B(n497), .Z(n1317) );
  XNOR U1312 ( .A(p_input[69]), .B(n1318), .Z(n497) );
  AND U1313 ( .A(n173), .B(n1319), .Z(n1318) );
  XOR U1314 ( .A(p_input[69]), .B(p_input[101]), .Z(n1319) );
  XNOR U1315 ( .A(n494), .B(n1314), .Z(n1316) );
  XOR U1316 ( .A(n1320), .B(n1321), .Z(n494) );
  AND U1317 ( .A(n170), .B(n1322), .Z(n1321) );
  XOR U1318 ( .A(p_input[5]), .B(p_input[37]), .Z(n1322) );
  XOR U1319 ( .A(n1323), .B(n1324), .Z(n1314) );
  AND U1320 ( .A(n1325), .B(n1326), .Z(n1324) );
  XOR U1321 ( .A(n1323), .B(n509), .Z(n1326) );
  XNOR U1322 ( .A(p_input[68]), .B(n1327), .Z(n509) );
  AND U1323 ( .A(n173), .B(n1328), .Z(n1327) );
  XOR U1324 ( .A(p_input[68]), .B(p_input[100]), .Z(n1328) );
  XNOR U1325 ( .A(n506), .B(n1323), .Z(n1325) );
  XOR U1326 ( .A(n1329), .B(n1330), .Z(n506) );
  AND U1327 ( .A(n170), .B(n1331), .Z(n1330) );
  XOR U1328 ( .A(p_input[4]), .B(p_input[36]), .Z(n1331) );
  XOR U1329 ( .A(n1332), .B(n1333), .Z(n1323) );
  AND U1330 ( .A(n1334), .B(n1335), .Z(n1333) );
  XOR U1331 ( .A(n1332), .B(n521), .Z(n1335) );
  XNOR U1332 ( .A(p_input[67]), .B(n1336), .Z(n521) );
  AND U1333 ( .A(n173), .B(n1337), .Z(n1336) );
  XOR U1334 ( .A(p_input[99]), .B(p_input[67]), .Z(n1337) );
  XNOR U1335 ( .A(n518), .B(n1332), .Z(n1334) );
  XOR U1336 ( .A(n1338), .B(n1339), .Z(n518) );
  AND U1337 ( .A(n170), .B(n1340), .Z(n1339) );
  XOR U1338 ( .A(p_input[3]), .B(p_input[35]), .Z(n1340) );
  XOR U1339 ( .A(n1341), .B(n1342), .Z(n1332) );
  AND U1340 ( .A(n1343), .B(n1344), .Z(n1342) );
  XOR U1341 ( .A(n1341), .B(n533), .Z(n1344) );
  XNOR U1342 ( .A(p_input[66]), .B(n1345), .Z(n533) );
  AND U1343 ( .A(n173), .B(n1346), .Z(n1345) );
  XOR U1344 ( .A(p_input[98]), .B(p_input[66]), .Z(n1346) );
  XNOR U1345 ( .A(n530), .B(n1341), .Z(n1343) );
  XOR U1346 ( .A(n1347), .B(n1348), .Z(n530) );
  AND U1347 ( .A(n170), .B(n1349), .Z(n1348) );
  XOR U1348 ( .A(p_input[34]), .B(p_input[2]), .Z(n1349) );
  XOR U1349 ( .A(n1350), .B(n1351), .Z(n1341) );
  AND U1350 ( .A(n1352), .B(n1353), .Z(n1351) );
  XNOR U1351 ( .A(n1354), .B(n545), .Z(n1353) );
  XNOR U1352 ( .A(p_input[65]), .B(n1355), .Z(n545) );
  AND U1353 ( .A(n173), .B(n1356), .Z(n1355) );
  XNOR U1354 ( .A(p_input[97]), .B(n1357), .Z(n1356) );
  IV U1355 ( .A(p_input[65]), .Z(n1357) );
  XNOR U1356 ( .A(n542), .B(n1350), .Z(n1352) );
  XNOR U1357 ( .A(p_input[1]), .B(n1358), .Z(n542) );
  AND U1358 ( .A(n170), .B(n1359), .Z(n1358) );
  XOR U1359 ( .A(p_input[33]), .B(p_input[1]), .Z(n1359) );
  IV U1360 ( .A(n1354), .Z(n1350) );
  AND U1361 ( .A(n1080), .B(n1083), .Z(n1354) );
  XOR U1362 ( .A(p_input[64]), .B(n1360), .Z(n1083) );
  AND U1363 ( .A(n173), .B(n1361), .Z(n1360) );
  XOR U1364 ( .A(p_input[96]), .B(p_input[64]), .Z(n1361) );
  XOR U1365 ( .A(n1362), .B(n1363), .Z(n173) );
  AND U1366 ( .A(n1364), .B(n1365), .Z(n1363) );
  XNOR U1367 ( .A(p_input[127]), .B(n1362), .Z(n1365) );
  XOR U1368 ( .A(n1362), .B(p_input[95]), .Z(n1364) );
  XOR U1369 ( .A(n1366), .B(n1367), .Z(n1362) );
  AND U1370 ( .A(n1368), .B(n1369), .Z(n1367) );
  XNOR U1371 ( .A(p_input[126]), .B(n1366), .Z(n1369) );
  XOR U1372 ( .A(n1366), .B(p_input[94]), .Z(n1368) );
  XOR U1373 ( .A(n1370), .B(n1371), .Z(n1366) );
  AND U1374 ( .A(n1372), .B(n1373), .Z(n1371) );
  XNOR U1375 ( .A(p_input[125]), .B(n1370), .Z(n1373) );
  XOR U1376 ( .A(n1370), .B(p_input[93]), .Z(n1372) );
  XOR U1377 ( .A(n1374), .B(n1375), .Z(n1370) );
  AND U1378 ( .A(n1376), .B(n1377), .Z(n1375) );
  XNOR U1379 ( .A(p_input[124]), .B(n1374), .Z(n1377) );
  XOR U1380 ( .A(n1374), .B(p_input[92]), .Z(n1376) );
  XOR U1381 ( .A(n1378), .B(n1379), .Z(n1374) );
  AND U1382 ( .A(n1380), .B(n1381), .Z(n1379) );
  XNOR U1383 ( .A(p_input[123]), .B(n1378), .Z(n1381) );
  XOR U1384 ( .A(n1378), .B(p_input[91]), .Z(n1380) );
  XOR U1385 ( .A(n1382), .B(n1383), .Z(n1378) );
  AND U1386 ( .A(n1384), .B(n1385), .Z(n1383) );
  XNOR U1387 ( .A(p_input[122]), .B(n1382), .Z(n1385) );
  XOR U1388 ( .A(n1382), .B(p_input[90]), .Z(n1384) );
  XOR U1389 ( .A(n1386), .B(n1387), .Z(n1382) );
  AND U1390 ( .A(n1388), .B(n1389), .Z(n1387) );
  XNOR U1391 ( .A(p_input[121]), .B(n1386), .Z(n1389) );
  XOR U1392 ( .A(n1386), .B(p_input[89]), .Z(n1388) );
  XOR U1393 ( .A(n1390), .B(n1391), .Z(n1386) );
  AND U1394 ( .A(n1392), .B(n1393), .Z(n1391) );
  XNOR U1395 ( .A(p_input[120]), .B(n1390), .Z(n1393) );
  XOR U1396 ( .A(n1390), .B(p_input[88]), .Z(n1392) );
  XOR U1397 ( .A(n1394), .B(n1395), .Z(n1390) );
  AND U1398 ( .A(n1396), .B(n1397), .Z(n1395) );
  XNOR U1399 ( .A(p_input[119]), .B(n1394), .Z(n1397) );
  XOR U1400 ( .A(n1394), .B(p_input[87]), .Z(n1396) );
  XOR U1401 ( .A(n1398), .B(n1399), .Z(n1394) );
  AND U1402 ( .A(n1400), .B(n1401), .Z(n1399) );
  XNOR U1403 ( .A(p_input[118]), .B(n1398), .Z(n1401) );
  XOR U1404 ( .A(n1398), .B(p_input[86]), .Z(n1400) );
  XOR U1405 ( .A(n1402), .B(n1403), .Z(n1398) );
  AND U1406 ( .A(n1404), .B(n1405), .Z(n1403) );
  XNOR U1407 ( .A(p_input[117]), .B(n1402), .Z(n1405) );
  XOR U1408 ( .A(n1402), .B(p_input[85]), .Z(n1404) );
  XOR U1409 ( .A(n1406), .B(n1407), .Z(n1402) );
  AND U1410 ( .A(n1408), .B(n1409), .Z(n1407) );
  XNOR U1411 ( .A(p_input[116]), .B(n1406), .Z(n1409) );
  XOR U1412 ( .A(n1406), .B(p_input[84]), .Z(n1408) );
  XOR U1413 ( .A(n1410), .B(n1411), .Z(n1406) );
  AND U1414 ( .A(n1412), .B(n1413), .Z(n1411) );
  XNOR U1415 ( .A(p_input[115]), .B(n1410), .Z(n1413) );
  XOR U1416 ( .A(n1410), .B(p_input[83]), .Z(n1412) );
  XOR U1417 ( .A(n1414), .B(n1415), .Z(n1410) );
  AND U1418 ( .A(n1416), .B(n1417), .Z(n1415) );
  XNOR U1419 ( .A(p_input[114]), .B(n1414), .Z(n1417) );
  XOR U1420 ( .A(n1414), .B(p_input[82]), .Z(n1416) );
  XOR U1421 ( .A(n1418), .B(n1419), .Z(n1414) );
  AND U1422 ( .A(n1420), .B(n1421), .Z(n1419) );
  XNOR U1423 ( .A(p_input[113]), .B(n1418), .Z(n1421) );
  XOR U1424 ( .A(n1418), .B(p_input[81]), .Z(n1420) );
  XOR U1425 ( .A(n1422), .B(n1423), .Z(n1418) );
  AND U1426 ( .A(n1424), .B(n1425), .Z(n1423) );
  XNOR U1427 ( .A(p_input[112]), .B(n1422), .Z(n1425) );
  XOR U1428 ( .A(n1422), .B(p_input[80]), .Z(n1424) );
  XOR U1429 ( .A(n1426), .B(n1427), .Z(n1422) );
  AND U1430 ( .A(n1428), .B(n1429), .Z(n1427) );
  XNOR U1431 ( .A(p_input[111]), .B(n1426), .Z(n1429) );
  XOR U1432 ( .A(n1426), .B(p_input[79]), .Z(n1428) );
  XOR U1433 ( .A(n1430), .B(n1431), .Z(n1426) );
  AND U1434 ( .A(n1432), .B(n1433), .Z(n1431) );
  XNOR U1435 ( .A(p_input[110]), .B(n1430), .Z(n1433) );
  XOR U1436 ( .A(n1430), .B(p_input[78]), .Z(n1432) );
  XOR U1437 ( .A(n1434), .B(n1435), .Z(n1430) );
  AND U1438 ( .A(n1436), .B(n1437), .Z(n1435) );
  XNOR U1439 ( .A(p_input[109]), .B(n1434), .Z(n1437) );
  XOR U1440 ( .A(n1434), .B(p_input[77]), .Z(n1436) );
  XOR U1441 ( .A(n1438), .B(n1439), .Z(n1434) );
  AND U1442 ( .A(n1440), .B(n1441), .Z(n1439) );
  XNOR U1443 ( .A(p_input[108]), .B(n1438), .Z(n1441) );
  XOR U1444 ( .A(n1438), .B(p_input[76]), .Z(n1440) );
  XOR U1445 ( .A(n1442), .B(n1443), .Z(n1438) );
  AND U1446 ( .A(n1444), .B(n1445), .Z(n1443) );
  XNOR U1447 ( .A(p_input[107]), .B(n1442), .Z(n1445) );
  XOR U1448 ( .A(n1442), .B(p_input[75]), .Z(n1444) );
  XOR U1449 ( .A(n1446), .B(n1447), .Z(n1442) );
  AND U1450 ( .A(n1448), .B(n1449), .Z(n1447) );
  XNOR U1451 ( .A(p_input[106]), .B(n1446), .Z(n1449) );
  XOR U1452 ( .A(n1446), .B(p_input[74]), .Z(n1448) );
  XOR U1453 ( .A(n1450), .B(n1451), .Z(n1446) );
  AND U1454 ( .A(n1452), .B(n1453), .Z(n1451) );
  XNOR U1455 ( .A(p_input[105]), .B(n1450), .Z(n1453) );
  XOR U1456 ( .A(n1450), .B(p_input[73]), .Z(n1452) );
  XOR U1457 ( .A(n1454), .B(n1455), .Z(n1450) );
  AND U1458 ( .A(n1456), .B(n1457), .Z(n1455) );
  XNOR U1459 ( .A(p_input[104]), .B(n1454), .Z(n1457) );
  XOR U1460 ( .A(n1454), .B(p_input[72]), .Z(n1456) );
  XOR U1461 ( .A(n1458), .B(n1459), .Z(n1454) );
  AND U1462 ( .A(n1460), .B(n1461), .Z(n1459) );
  XNOR U1463 ( .A(p_input[103]), .B(n1458), .Z(n1461) );
  XOR U1464 ( .A(n1458), .B(p_input[71]), .Z(n1460) );
  XOR U1465 ( .A(n1462), .B(n1463), .Z(n1458) );
  AND U1466 ( .A(n1464), .B(n1465), .Z(n1463) );
  XNOR U1467 ( .A(p_input[102]), .B(n1462), .Z(n1465) );
  XOR U1468 ( .A(n1462), .B(p_input[70]), .Z(n1464) );
  XOR U1469 ( .A(n1466), .B(n1467), .Z(n1462) );
  AND U1470 ( .A(n1468), .B(n1469), .Z(n1467) );
  XNOR U1471 ( .A(p_input[101]), .B(n1466), .Z(n1469) );
  XOR U1472 ( .A(n1466), .B(p_input[69]), .Z(n1468) );
  XOR U1473 ( .A(n1470), .B(n1471), .Z(n1466) );
  AND U1474 ( .A(n1472), .B(n1473), .Z(n1471) );
  XNOR U1475 ( .A(p_input[100]), .B(n1470), .Z(n1473) );
  XOR U1476 ( .A(n1470), .B(p_input[68]), .Z(n1472) );
  XOR U1477 ( .A(n1474), .B(n1475), .Z(n1470) );
  AND U1478 ( .A(n1476), .B(n1477), .Z(n1475) );
  XNOR U1479 ( .A(p_input[99]), .B(n1474), .Z(n1477) );
  XOR U1480 ( .A(n1474), .B(p_input[67]), .Z(n1476) );
  XOR U1481 ( .A(n1478), .B(n1479), .Z(n1474) );
  AND U1482 ( .A(n1480), .B(n1481), .Z(n1479) );
  XNOR U1483 ( .A(p_input[98]), .B(n1478), .Z(n1481) );
  XOR U1484 ( .A(n1478), .B(p_input[66]), .Z(n1480) );
  XNOR U1485 ( .A(n1482), .B(n1483), .Z(n1478) );
  AND U1486 ( .A(n1484), .B(n1485), .Z(n1483) );
  XOR U1487 ( .A(p_input[97]), .B(n1482), .Z(n1485) );
  XNOR U1488 ( .A(p_input[65]), .B(n1482), .Z(n1484) );
  AND U1489 ( .A(p_input[96]), .B(n1486), .Z(n1482) );
  IV U1490 ( .A(p_input[64]), .Z(n1486) );
  XNOR U1491 ( .A(p_input[0]), .B(n1487), .Z(n1080) );
  AND U1492 ( .A(n170), .B(n1488), .Z(n1487) );
  XOR U1493 ( .A(p_input[32]), .B(p_input[0]), .Z(n1488) );
  XOR U1494 ( .A(n1489), .B(n1490), .Z(n170) );
  AND U1495 ( .A(n1491), .B(n1492), .Z(n1490) );
  XNOR U1496 ( .A(p_input[63]), .B(n1489), .Z(n1492) );
  XOR U1497 ( .A(n1489), .B(p_input[31]), .Z(n1491) );
  XOR U1498 ( .A(n1493), .B(n1494), .Z(n1489) );
  AND U1499 ( .A(n1495), .B(n1496), .Z(n1494) );
  XNOR U1500 ( .A(p_input[62]), .B(n1493), .Z(n1496) );
  XNOR U1501 ( .A(n1493), .B(n1095), .Z(n1495) );
  IV U1502 ( .A(p_input[30]), .Z(n1095) );
  XOR U1503 ( .A(n1497), .B(n1498), .Z(n1493) );
  AND U1504 ( .A(n1499), .B(n1500), .Z(n1498) );
  XNOR U1505 ( .A(p_input[61]), .B(n1497), .Z(n1500) );
  XNOR U1506 ( .A(n1497), .B(n1104), .Z(n1499) );
  IV U1507 ( .A(p_input[29]), .Z(n1104) );
  XOR U1508 ( .A(n1501), .B(n1502), .Z(n1497) );
  AND U1509 ( .A(n1503), .B(n1504), .Z(n1502) );
  XNOR U1510 ( .A(p_input[60]), .B(n1501), .Z(n1504) );
  XNOR U1511 ( .A(n1501), .B(n1113), .Z(n1503) );
  IV U1512 ( .A(p_input[28]), .Z(n1113) );
  XOR U1513 ( .A(n1505), .B(n1506), .Z(n1501) );
  AND U1514 ( .A(n1507), .B(n1508), .Z(n1506) );
  XNOR U1515 ( .A(p_input[59]), .B(n1505), .Z(n1508) );
  XNOR U1516 ( .A(n1505), .B(n1122), .Z(n1507) );
  IV U1517 ( .A(p_input[27]), .Z(n1122) );
  XOR U1518 ( .A(n1509), .B(n1510), .Z(n1505) );
  AND U1519 ( .A(n1511), .B(n1512), .Z(n1510) );
  XNOR U1520 ( .A(p_input[58]), .B(n1509), .Z(n1512) );
  XNOR U1521 ( .A(n1509), .B(n1131), .Z(n1511) );
  IV U1522 ( .A(p_input[26]), .Z(n1131) );
  XOR U1523 ( .A(n1513), .B(n1514), .Z(n1509) );
  AND U1524 ( .A(n1515), .B(n1516), .Z(n1514) );
  XNOR U1525 ( .A(p_input[57]), .B(n1513), .Z(n1516) );
  XNOR U1526 ( .A(n1513), .B(n1140), .Z(n1515) );
  IV U1527 ( .A(p_input[25]), .Z(n1140) );
  XOR U1528 ( .A(n1517), .B(n1518), .Z(n1513) );
  AND U1529 ( .A(n1519), .B(n1520), .Z(n1518) );
  XNOR U1530 ( .A(p_input[56]), .B(n1517), .Z(n1520) );
  XNOR U1531 ( .A(n1517), .B(n1149), .Z(n1519) );
  IV U1532 ( .A(p_input[24]), .Z(n1149) );
  XOR U1533 ( .A(n1521), .B(n1522), .Z(n1517) );
  AND U1534 ( .A(n1523), .B(n1524), .Z(n1522) );
  XNOR U1535 ( .A(p_input[55]), .B(n1521), .Z(n1524) );
  XNOR U1536 ( .A(n1521), .B(n1158), .Z(n1523) );
  IV U1537 ( .A(p_input[23]), .Z(n1158) );
  XOR U1538 ( .A(n1525), .B(n1526), .Z(n1521) );
  AND U1539 ( .A(n1527), .B(n1528), .Z(n1526) );
  XNOR U1540 ( .A(p_input[54]), .B(n1525), .Z(n1528) );
  XNOR U1541 ( .A(n1525), .B(n1167), .Z(n1527) );
  IV U1542 ( .A(p_input[22]), .Z(n1167) );
  XOR U1543 ( .A(n1529), .B(n1530), .Z(n1525) );
  AND U1544 ( .A(n1531), .B(n1532), .Z(n1530) );
  XNOR U1545 ( .A(p_input[53]), .B(n1529), .Z(n1532) );
  XNOR U1546 ( .A(n1529), .B(n1176), .Z(n1531) );
  IV U1547 ( .A(p_input[21]), .Z(n1176) );
  XOR U1548 ( .A(n1533), .B(n1534), .Z(n1529) );
  AND U1549 ( .A(n1535), .B(n1536), .Z(n1534) );
  XNOR U1550 ( .A(p_input[52]), .B(n1533), .Z(n1536) );
  XNOR U1551 ( .A(n1533), .B(n1185), .Z(n1535) );
  IV U1552 ( .A(p_input[20]), .Z(n1185) );
  XOR U1553 ( .A(n1537), .B(n1538), .Z(n1533) );
  AND U1554 ( .A(n1539), .B(n1540), .Z(n1538) );
  XNOR U1555 ( .A(p_input[51]), .B(n1537), .Z(n1540) );
  XNOR U1556 ( .A(n1537), .B(n1194), .Z(n1539) );
  IV U1557 ( .A(p_input[19]), .Z(n1194) );
  XOR U1558 ( .A(n1541), .B(n1542), .Z(n1537) );
  AND U1559 ( .A(n1543), .B(n1544), .Z(n1542) );
  XNOR U1560 ( .A(p_input[50]), .B(n1541), .Z(n1544) );
  XNOR U1561 ( .A(n1541), .B(n1203), .Z(n1543) );
  IV U1562 ( .A(p_input[18]), .Z(n1203) );
  XOR U1563 ( .A(n1545), .B(n1546), .Z(n1541) );
  AND U1564 ( .A(n1547), .B(n1548), .Z(n1546) );
  XNOR U1565 ( .A(p_input[49]), .B(n1545), .Z(n1548) );
  XNOR U1566 ( .A(n1545), .B(n1212), .Z(n1547) );
  IV U1567 ( .A(p_input[17]), .Z(n1212) );
  XOR U1568 ( .A(n1549), .B(n1550), .Z(n1545) );
  AND U1569 ( .A(n1551), .B(n1552), .Z(n1550) );
  XNOR U1570 ( .A(p_input[48]), .B(n1549), .Z(n1552) );
  XNOR U1571 ( .A(n1549), .B(n1221), .Z(n1551) );
  IV U1572 ( .A(p_input[16]), .Z(n1221) );
  XOR U1573 ( .A(n1553), .B(n1554), .Z(n1549) );
  AND U1574 ( .A(n1555), .B(n1556), .Z(n1554) );
  XNOR U1575 ( .A(p_input[47]), .B(n1553), .Z(n1556) );
  XNOR U1576 ( .A(n1553), .B(n1230), .Z(n1555) );
  IV U1577 ( .A(p_input[15]), .Z(n1230) );
  XOR U1578 ( .A(n1557), .B(n1558), .Z(n1553) );
  AND U1579 ( .A(n1559), .B(n1560), .Z(n1558) );
  XNOR U1580 ( .A(p_input[46]), .B(n1557), .Z(n1560) );
  XNOR U1581 ( .A(n1557), .B(n1239), .Z(n1559) );
  IV U1582 ( .A(p_input[14]), .Z(n1239) );
  XOR U1583 ( .A(n1561), .B(n1562), .Z(n1557) );
  AND U1584 ( .A(n1563), .B(n1564), .Z(n1562) );
  XNOR U1585 ( .A(p_input[45]), .B(n1561), .Z(n1564) );
  XNOR U1586 ( .A(n1561), .B(n1248), .Z(n1563) );
  IV U1587 ( .A(p_input[13]), .Z(n1248) );
  XOR U1588 ( .A(n1565), .B(n1566), .Z(n1561) );
  AND U1589 ( .A(n1567), .B(n1568), .Z(n1566) );
  XNOR U1590 ( .A(p_input[44]), .B(n1565), .Z(n1568) );
  XNOR U1591 ( .A(n1565), .B(n1257), .Z(n1567) );
  IV U1592 ( .A(p_input[12]), .Z(n1257) );
  XOR U1593 ( .A(n1569), .B(n1570), .Z(n1565) );
  AND U1594 ( .A(n1571), .B(n1572), .Z(n1570) );
  XNOR U1595 ( .A(p_input[43]), .B(n1569), .Z(n1572) );
  XNOR U1596 ( .A(n1569), .B(n1266), .Z(n1571) );
  IV U1597 ( .A(p_input[11]), .Z(n1266) );
  XOR U1598 ( .A(n1573), .B(n1574), .Z(n1569) );
  AND U1599 ( .A(n1575), .B(n1576), .Z(n1574) );
  XNOR U1600 ( .A(p_input[42]), .B(n1573), .Z(n1576) );
  XNOR U1601 ( .A(n1573), .B(n1275), .Z(n1575) );
  IV U1602 ( .A(p_input[10]), .Z(n1275) );
  XOR U1603 ( .A(n1577), .B(n1578), .Z(n1573) );
  AND U1604 ( .A(n1579), .B(n1580), .Z(n1578) );
  XNOR U1605 ( .A(p_input[41]), .B(n1577), .Z(n1580) );
  XNOR U1606 ( .A(n1577), .B(n1284), .Z(n1579) );
  IV U1607 ( .A(p_input[9]), .Z(n1284) );
  XOR U1608 ( .A(n1581), .B(n1582), .Z(n1577) );
  AND U1609 ( .A(n1583), .B(n1584), .Z(n1582) );
  XNOR U1610 ( .A(p_input[40]), .B(n1581), .Z(n1584) );
  XNOR U1611 ( .A(n1581), .B(n1293), .Z(n1583) );
  IV U1612 ( .A(p_input[8]), .Z(n1293) );
  XOR U1613 ( .A(n1585), .B(n1586), .Z(n1581) );
  AND U1614 ( .A(n1587), .B(n1588), .Z(n1586) );
  XNOR U1615 ( .A(p_input[39]), .B(n1585), .Z(n1588) );
  XNOR U1616 ( .A(n1585), .B(n1302), .Z(n1587) );
  IV U1617 ( .A(p_input[7]), .Z(n1302) );
  XOR U1618 ( .A(n1589), .B(n1590), .Z(n1585) );
  AND U1619 ( .A(n1591), .B(n1592), .Z(n1590) );
  XNOR U1620 ( .A(p_input[38]), .B(n1589), .Z(n1592) );
  XNOR U1621 ( .A(n1589), .B(n1311), .Z(n1591) );
  IV U1622 ( .A(p_input[6]), .Z(n1311) );
  XOR U1623 ( .A(n1593), .B(n1594), .Z(n1589) );
  AND U1624 ( .A(n1595), .B(n1596), .Z(n1594) );
  XNOR U1625 ( .A(p_input[37]), .B(n1593), .Z(n1596) );
  XNOR U1626 ( .A(n1593), .B(n1320), .Z(n1595) );
  IV U1627 ( .A(p_input[5]), .Z(n1320) );
  XOR U1628 ( .A(n1597), .B(n1598), .Z(n1593) );
  AND U1629 ( .A(n1599), .B(n1600), .Z(n1598) );
  XNOR U1630 ( .A(p_input[36]), .B(n1597), .Z(n1600) );
  XNOR U1631 ( .A(n1597), .B(n1329), .Z(n1599) );
  IV U1632 ( .A(p_input[4]), .Z(n1329) );
  XOR U1633 ( .A(n1601), .B(n1602), .Z(n1597) );
  AND U1634 ( .A(n1603), .B(n1604), .Z(n1602) );
  XNOR U1635 ( .A(p_input[35]), .B(n1601), .Z(n1604) );
  XNOR U1636 ( .A(n1601), .B(n1338), .Z(n1603) );
  IV U1637 ( .A(p_input[3]), .Z(n1338) );
  XOR U1638 ( .A(n1605), .B(n1606), .Z(n1601) );
  AND U1639 ( .A(n1607), .B(n1608), .Z(n1606) );
  XNOR U1640 ( .A(p_input[34]), .B(n1605), .Z(n1608) );
  XNOR U1641 ( .A(n1605), .B(n1347), .Z(n1607) );
  IV U1642 ( .A(p_input[2]), .Z(n1347) );
  XNOR U1643 ( .A(n1609), .B(n1610), .Z(n1605) );
  AND U1644 ( .A(n1611), .B(n1612), .Z(n1610) );
  XOR U1645 ( .A(p_input[33]), .B(n1609), .Z(n1612) );
  XNOR U1646 ( .A(p_input[1]), .B(n1609), .Z(n1611) );
  AND U1647 ( .A(p_input[32]), .B(n1613), .Z(n1609) );
  IV U1648 ( .A(p_input[0]), .Z(n1613) );
endmodule

